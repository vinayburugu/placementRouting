magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 37 3 38 4 
<< m1 >>
rect 38 3 39 4 
<< m1 >>
rect 39 3 40 4 
<< m1 >>
rect 40 3 41 4 
<< m1 >>
rect 41 3 42 4 
<< m1 >>
rect 42 3 43 4 
<< m1 >>
rect 43 3 44 4 
<< m1 >>
rect 44 3 45 4 
<< m1 >>
rect 45 3 46 4 
<< m1 >>
rect 46 3 47 4 
<< m1 >>
rect 47 3 48 4 
<< m1 >>
rect 48 3 49 4 
<< m1 >>
rect 49 3 50 4 
<< m1 >>
rect 50 3 51 4 
<< m1 >>
rect 51 3 52 4 
<< m1 >>
rect 52 3 53 4 
<< m1 >>
rect 53 3 54 4 
<< m1 >>
rect 54 3 55 4 
<< m1 >>
rect 55 3 56 4 
<< m1 >>
rect 56 3 57 4 
<< m1 >>
rect 57 3 58 4 
<< m1 >>
rect 58 3 59 4 
<< m1 >>
rect 59 3 60 4 
<< m1 >>
rect 60 3 61 4 
<< m1 >>
rect 61 3 62 4 
<< m1 >>
rect 62 3 63 4 
<< m1 >>
rect 63 3 64 4 
<< m1 >>
rect 64 3 65 4 
<< m1 >>
rect 65 3 66 4 
<< m1 >>
rect 66 3 67 4 
<< m1 >>
rect 67 3 68 4 
<< m1 >>
rect 68 3 69 4 
<< m1 >>
rect 69 3 70 4 
<< m1 >>
rect 70 3 71 4 
<< m1 >>
rect 71 3 72 4 
<< m1 >>
rect 72 3 73 4 
<< m1 >>
rect 73 3 74 4 
<< m1 >>
rect 74 3 75 4 
<< m1 >>
rect 75 3 76 4 
<< m1 >>
rect 76 3 77 4 
<< m1 >>
rect 77 3 78 4 
<< m1 >>
rect 78 3 79 4 
<< m1 >>
rect 79 3 80 4 
<< m1 >>
rect 80 3 81 4 
<< m1 >>
rect 81 3 82 4 
<< m1 >>
rect 82 3 83 4 
<< m1 >>
rect 83 3 84 4 
<< m1 >>
rect 84 3 85 4 
<< m1 >>
rect 85 3 86 4 
<< m1 >>
rect 86 3 87 4 
<< m1 >>
rect 87 3 88 4 
<< m1 >>
rect 88 3 89 4 
<< m1 >>
rect 89 3 90 4 
<< m1 >>
rect 90 3 91 4 
<< m1 >>
rect 91 3 92 4 
<< m1 >>
rect 92 3 93 4 
<< m1 >>
rect 93 3 94 4 
<< m1 >>
rect 94 3 95 4 
<< m1 >>
rect 95 3 96 4 
<< m1 >>
rect 96 3 97 4 
<< m1 >>
rect 97 3 98 4 
<< m1 >>
rect 98 3 99 4 
<< m1 >>
rect 99 3 100 4 
<< m1 >>
rect 100 3 101 4 
<< m1 >>
rect 101 3 102 4 
<< m1 >>
rect 102 3 103 4 
<< m1 >>
rect 103 3 104 4 
<< m1 >>
rect 104 3 105 4 
<< m1 >>
rect 105 3 106 4 
<< m1 >>
rect 106 3 107 4 
<< m1 >>
rect 107 3 108 4 
<< m1 >>
rect 108 3 109 4 
<< m1 >>
rect 109 3 110 4 
<< m1 >>
rect 110 3 111 4 
<< m1 >>
rect 111 3 112 4 
<< m1 >>
rect 112 3 113 4 
<< m1 >>
rect 113 3 114 4 
<< m1 >>
rect 114 3 115 4 
<< m1 >>
rect 115 3 116 4 
<< m1 >>
rect 116 3 117 4 
<< m1 >>
rect 117 3 118 4 
<< m1 >>
rect 118 3 119 4 
<< m1 >>
rect 119 3 120 4 
<< m1 >>
rect 120 3 121 4 
<< m1 >>
rect 121 3 122 4 
<< m1 >>
rect 122 3 123 4 
<< m1 >>
rect 123 3 124 4 
<< m1 >>
rect 124 3 125 4 
<< m1 >>
rect 125 3 126 4 
<< m1 >>
rect 126 3 127 4 
<< m1 >>
rect 127 3 128 4 
<< m1 >>
rect 128 3 129 4 
<< m1 >>
rect 129 3 130 4 
<< m1 >>
rect 130 3 131 4 
<< m1 >>
rect 131 3 132 4 
<< m1 >>
rect 132 3 133 4 
<< m1 >>
rect 133 3 134 4 
<< m1 >>
rect 134 3 135 4 
<< m1 >>
rect 135 3 136 4 
<< m1 >>
rect 136 3 137 4 
<< m1 >>
rect 137 3 138 4 
<< m1 >>
rect 138 3 139 4 
<< m1 >>
rect 139 3 140 4 
<< m1 >>
rect 140 3 141 4 
<< m1 >>
rect 141 3 142 4 
<< m1 >>
rect 142 3 143 4 
<< m1 >>
rect 143 3 144 4 
<< m1 >>
rect 144 3 145 4 
<< m1 >>
rect 145 3 146 4 
<< m1 >>
rect 146 3 147 4 
<< m1 >>
rect 147 3 148 4 
<< m1 >>
rect 148 3 149 4 
<< m1 >>
rect 149 3 150 4 
<< m1 >>
rect 150 3 151 4 
<< m1 >>
rect 151 3 152 4 
<< m1 >>
rect 152 3 153 4 
<< m1 >>
rect 153 3 154 4 
<< m1 >>
rect 154 3 155 4 
<< m1 >>
rect 155 3 156 4 
<< m1 >>
rect 156 3 157 4 
<< m1 >>
rect 157 3 158 4 
<< m1 >>
rect 158 3 159 4 
<< m1 >>
rect 159 3 160 4 
<< m1 >>
rect 160 3 161 4 
<< m1 >>
rect 161 3 162 4 
<< m1 >>
rect 162 3 163 4 
<< m1 >>
rect 163 3 164 4 
<< m1 >>
rect 164 3 165 4 
<< m1 >>
rect 165 3 166 4 
<< m1 >>
rect 166 3 167 4 
<< m1 >>
rect 167 3 168 4 
<< m1 >>
rect 168 3 169 4 
<< m1 >>
rect 169 3 170 4 
<< m1 >>
rect 170 3 171 4 
<< m1 >>
rect 171 3 172 4 
<< m1 >>
rect 172 3 173 4 
<< m1 >>
rect 173 3 174 4 
<< m1 >>
rect 174 3 175 4 
<< m1 >>
rect 175 3 176 4 
<< m1 >>
rect 176 3 177 4 
<< m1 >>
rect 177 3 178 4 
<< m1 >>
rect 178 3 179 4 
<< m1 >>
rect 179 3 180 4 
<< m1 >>
rect 180 3 181 4 
<< m1 >>
rect 181 3 182 4 
<< m1 >>
rect 182 3 183 4 
<< m1 >>
rect 183 3 184 4 
<< m1 >>
rect 184 3 185 4 
<< m1 >>
rect 185 3 186 4 
<< m1 >>
rect 186 3 187 4 
<< m1 >>
rect 187 3 188 4 
<< m1 >>
rect 188 3 189 4 
<< m1 >>
rect 189 3 190 4 
<< m1 >>
rect 190 3 191 4 
<< m1 >>
rect 191 3 192 4 
<< m1 >>
rect 192 3 193 4 
<< m1 >>
rect 193 3 194 4 
<< m1 >>
rect 194 3 195 4 
<< m1 >>
rect 195 3 196 4 
<< m1 >>
rect 196 3 197 4 
<< m1 >>
rect 197 3 198 4 
<< m1 >>
rect 198 3 199 4 
<< m1 >>
rect 199 3 200 4 
<< m1 >>
rect 200 3 201 4 
<< m1 >>
rect 201 3 202 4 
<< m1 >>
rect 37 4 38 5 
<< m1 >>
rect 201 4 202 5 
<< m1 >>
rect 37 5 38 6 
<< m1 >>
rect 49 5 50 6 
<< m2 >>
rect 49 5 50 6 
<< m2c >>
rect 49 5 50 6 
<< m1 >>
rect 49 5 50 6 
<< m2 >>
rect 49 5 50 6 
<< m1 >>
rect 50 5 51 6 
<< m1 >>
rect 51 5 52 6 
<< m1 >>
rect 52 5 53 6 
<< m1 >>
rect 53 5 54 6 
<< m1 >>
rect 54 5 55 6 
<< m1 >>
rect 55 5 56 6 
<< m1 >>
rect 56 5 57 6 
<< m2 >>
rect 56 5 57 6 
<< m2c >>
rect 56 5 57 6 
<< m1 >>
rect 56 5 57 6 
<< m2 >>
rect 56 5 57 6 
<< m2 >>
rect 57 5 58 6 
<< m1 >>
rect 58 5 59 6 
<< m2 >>
rect 58 5 59 6 
<< m1 >>
rect 59 5 60 6 
<< m2 >>
rect 59 5 60 6 
<< m1 >>
rect 60 5 61 6 
<< m2 >>
rect 60 5 61 6 
<< m1 >>
rect 61 5 62 6 
<< m2 >>
rect 61 5 62 6 
<< m1 >>
rect 62 5 63 6 
<< m2 >>
rect 62 5 63 6 
<< m1 >>
rect 63 5 64 6 
<< m2 >>
rect 63 5 64 6 
<< m1 >>
rect 64 5 65 6 
<< m2 >>
rect 64 5 65 6 
<< m1 >>
rect 65 5 66 6 
<< m2 >>
rect 65 5 66 6 
<< m1 >>
rect 66 5 67 6 
<< m2 >>
rect 66 5 67 6 
<< m1 >>
rect 67 5 68 6 
<< m2 >>
rect 67 5 68 6 
<< m1 >>
rect 68 5 69 6 
<< m2 >>
rect 68 5 69 6 
<< m1 >>
rect 69 5 70 6 
<< m2 >>
rect 69 5 70 6 
<< m1 >>
rect 70 5 71 6 
<< m2 >>
rect 70 5 71 6 
<< m1 >>
rect 71 5 72 6 
<< m2 >>
rect 71 5 72 6 
<< m1 >>
rect 72 5 73 6 
<< m2 >>
rect 72 5 73 6 
<< m1 >>
rect 73 5 74 6 
<< m2 >>
rect 73 5 74 6 
<< m1 >>
rect 74 5 75 6 
<< m2 >>
rect 74 5 75 6 
<< m1 >>
rect 75 5 76 6 
<< m2 >>
rect 75 5 76 6 
<< m1 >>
rect 76 5 77 6 
<< m2 >>
rect 76 5 77 6 
<< m1 >>
rect 77 5 78 6 
<< m2 >>
rect 77 5 78 6 
<< m1 >>
rect 78 5 79 6 
<< m2 >>
rect 78 5 79 6 
<< m1 >>
rect 79 5 80 6 
<< m2 >>
rect 79 5 80 6 
<< m1 >>
rect 80 5 81 6 
<< m2 >>
rect 80 5 81 6 
<< m1 >>
rect 81 5 82 6 
<< m2 >>
rect 81 5 82 6 
<< m1 >>
rect 82 5 83 6 
<< m2 >>
rect 82 5 83 6 
<< m1 >>
rect 83 5 84 6 
<< m2 >>
rect 83 5 84 6 
<< m1 >>
rect 84 5 85 6 
<< m2 >>
rect 84 5 85 6 
<< m1 >>
rect 85 5 86 6 
<< m2 >>
rect 85 5 86 6 
<< m1 >>
rect 86 5 87 6 
<< m2 >>
rect 86 5 87 6 
<< m1 >>
rect 87 5 88 6 
<< m2 >>
rect 87 5 88 6 
<< m1 >>
rect 88 5 89 6 
<< m2 >>
rect 88 5 89 6 
<< m1 >>
rect 89 5 90 6 
<< m2 >>
rect 89 5 90 6 
<< m1 >>
rect 90 5 91 6 
<< m2 >>
rect 90 5 91 6 
<< m1 >>
rect 91 5 92 6 
<< m2 >>
rect 91 5 92 6 
<< m1 >>
rect 92 5 93 6 
<< m2 >>
rect 92 5 93 6 
<< m1 >>
rect 93 5 94 6 
<< m2 >>
rect 93 5 94 6 
<< m1 >>
rect 94 5 95 6 
<< m2 >>
rect 94 5 95 6 
<< m1 >>
rect 95 5 96 6 
<< m2 >>
rect 95 5 96 6 
<< m1 >>
rect 96 5 97 6 
<< m2 >>
rect 96 5 97 6 
<< m1 >>
rect 97 5 98 6 
<< m2 >>
rect 97 5 98 6 
<< m1 >>
rect 98 5 99 6 
<< m2 >>
rect 98 5 99 6 
<< m1 >>
rect 99 5 100 6 
<< m2 >>
rect 99 5 100 6 
<< m1 >>
rect 100 5 101 6 
<< m2 >>
rect 100 5 101 6 
<< m1 >>
rect 101 5 102 6 
<< m2 >>
rect 101 5 102 6 
<< m1 >>
rect 102 5 103 6 
<< m2 >>
rect 102 5 103 6 
<< m1 >>
rect 103 5 104 6 
<< m2 >>
rect 103 5 104 6 
<< m1 >>
rect 104 5 105 6 
<< m2 >>
rect 104 5 105 6 
<< m1 >>
rect 105 5 106 6 
<< m2 >>
rect 105 5 106 6 
<< m1 >>
rect 106 5 107 6 
<< m2 >>
rect 106 5 107 6 
<< m1 >>
rect 107 5 108 6 
<< m2 >>
rect 107 5 108 6 
<< m1 >>
rect 108 5 109 6 
<< m2 >>
rect 108 5 109 6 
<< m1 >>
rect 109 5 110 6 
<< m2 >>
rect 109 5 110 6 
<< m1 >>
rect 110 5 111 6 
<< m2 >>
rect 110 5 111 6 
<< m1 >>
rect 111 5 112 6 
<< m2 >>
rect 111 5 112 6 
<< m1 >>
rect 112 5 113 6 
<< m2 >>
rect 112 5 113 6 
<< m1 >>
rect 113 5 114 6 
<< m2 >>
rect 113 5 114 6 
<< m1 >>
rect 114 5 115 6 
<< m2 >>
rect 114 5 115 6 
<< m1 >>
rect 115 5 116 6 
<< m2 >>
rect 115 5 116 6 
<< m1 >>
rect 116 5 117 6 
<< m2 >>
rect 116 5 117 6 
<< m1 >>
rect 117 5 118 6 
<< m2 >>
rect 117 5 118 6 
<< m1 >>
rect 118 5 119 6 
<< m2 >>
rect 118 5 119 6 
<< m1 >>
rect 119 5 120 6 
<< m2 >>
rect 119 5 120 6 
<< m1 >>
rect 120 5 121 6 
<< m2 >>
rect 120 5 121 6 
<< m1 >>
rect 121 5 122 6 
<< m2 >>
rect 121 5 122 6 
<< m1 >>
rect 122 5 123 6 
<< m2 >>
rect 122 5 123 6 
<< m1 >>
rect 123 5 124 6 
<< m2 >>
rect 123 5 124 6 
<< m1 >>
rect 124 5 125 6 
<< m2 >>
rect 124 5 125 6 
<< m1 >>
rect 125 5 126 6 
<< m2 >>
rect 125 5 126 6 
<< m1 >>
rect 126 5 127 6 
<< m2 >>
rect 126 5 127 6 
<< m1 >>
rect 127 5 128 6 
<< m2 >>
rect 127 5 128 6 
<< m1 >>
rect 128 5 129 6 
<< m2 >>
rect 128 5 129 6 
<< m1 >>
rect 129 5 130 6 
<< m2 >>
rect 129 5 130 6 
<< m1 >>
rect 130 5 131 6 
<< m2 >>
rect 130 5 131 6 
<< m1 >>
rect 131 5 132 6 
<< m1 >>
rect 132 5 133 6 
<< m1 >>
rect 133 5 134 6 
<< m1 >>
rect 134 5 135 6 
<< m1 >>
rect 135 5 136 6 
<< m1 >>
rect 136 5 137 6 
<< m1 >>
rect 137 5 138 6 
<< m1 >>
rect 138 5 139 6 
<< m1 >>
rect 139 5 140 6 
<< m1 >>
rect 140 5 141 6 
<< m1 >>
rect 141 5 142 6 
<< m1 >>
rect 142 5 143 6 
<< m1 >>
rect 143 5 144 6 
<< m1 >>
rect 144 5 145 6 
<< m1 >>
rect 145 5 146 6 
<< m1 >>
rect 146 5 147 6 
<< m2 >>
rect 146 5 147 6 
<< m1 >>
rect 147 5 148 6 
<< m2 >>
rect 147 5 148 6 
<< m1 >>
rect 148 5 149 6 
<< m2 >>
rect 148 5 149 6 
<< m1 >>
rect 149 5 150 6 
<< m2 >>
rect 149 5 150 6 
<< m1 >>
rect 150 5 151 6 
<< m2 >>
rect 150 5 151 6 
<< m1 >>
rect 151 5 152 6 
<< m2 >>
rect 151 5 152 6 
<< m1 >>
rect 152 5 153 6 
<< m2 >>
rect 152 5 153 6 
<< m1 >>
rect 153 5 154 6 
<< m2 >>
rect 153 5 154 6 
<< m1 >>
rect 154 5 155 6 
<< m2 >>
rect 154 5 155 6 
<< m1 >>
rect 155 5 156 6 
<< m2 >>
rect 155 5 156 6 
<< m1 >>
rect 156 5 157 6 
<< m2 >>
rect 156 5 157 6 
<< m1 >>
rect 157 5 158 6 
<< m2 >>
rect 157 5 158 6 
<< m1 >>
rect 158 5 159 6 
<< m2 >>
rect 158 5 159 6 
<< m1 >>
rect 159 5 160 6 
<< m2 >>
rect 159 5 160 6 
<< m1 >>
rect 160 5 161 6 
<< m2 >>
rect 160 5 161 6 
<< m1 >>
rect 161 5 162 6 
<< m2 >>
rect 161 5 162 6 
<< m1 >>
rect 162 5 163 6 
<< m2 >>
rect 162 5 163 6 
<< m1 >>
rect 163 5 164 6 
<< m2 >>
rect 163 5 164 6 
<< m1 >>
rect 164 5 165 6 
<< m2 >>
rect 164 5 165 6 
<< m1 >>
rect 165 5 166 6 
<< m2 >>
rect 165 5 166 6 
<< m1 >>
rect 166 5 167 6 
<< m2 >>
rect 166 5 167 6 
<< m1 >>
rect 167 5 168 6 
<< m2 >>
rect 167 5 168 6 
<< m1 >>
rect 168 5 169 6 
<< m2 >>
rect 168 5 169 6 
<< m1 >>
rect 169 5 170 6 
<< m2 >>
rect 169 5 170 6 
<< m1 >>
rect 170 5 171 6 
<< m2 >>
rect 170 5 171 6 
<< m1 >>
rect 171 5 172 6 
<< m2 >>
rect 171 5 172 6 
<< m1 >>
rect 172 5 173 6 
<< m2 >>
rect 172 5 173 6 
<< m1 >>
rect 173 5 174 6 
<< m2 >>
rect 173 5 174 6 
<< m1 >>
rect 174 5 175 6 
<< m2 >>
rect 174 5 175 6 
<< m1 >>
rect 175 5 176 6 
<< m2 >>
rect 175 5 176 6 
<< m1 >>
rect 176 5 177 6 
<< m2 >>
rect 176 5 177 6 
<< m1 >>
rect 177 5 178 6 
<< m2 >>
rect 177 5 178 6 
<< m1 >>
rect 178 5 179 6 
<< m2 >>
rect 178 5 179 6 
<< m1 >>
rect 179 5 180 6 
<< m2 >>
rect 179 5 180 6 
<< m1 >>
rect 180 5 181 6 
<< m2 >>
rect 180 5 181 6 
<< m1 >>
rect 181 5 182 6 
<< m2 >>
rect 181 5 182 6 
<< m1 >>
rect 182 5 183 6 
<< m2 >>
rect 182 5 183 6 
<< m1 >>
rect 183 5 184 6 
<< m2 >>
rect 183 5 184 6 
<< m1 >>
rect 184 5 185 6 
<< m2 >>
rect 184 5 185 6 
<< m1 >>
rect 185 5 186 6 
<< m2 >>
rect 185 5 186 6 
<< m1 >>
rect 186 5 187 6 
<< m2 >>
rect 186 5 187 6 
<< m1 >>
rect 187 5 188 6 
<< m2 >>
rect 187 5 188 6 
<< m1 >>
rect 188 5 189 6 
<< m2 >>
rect 188 5 189 6 
<< m1 >>
rect 189 5 190 6 
<< m2 >>
rect 189 5 190 6 
<< m1 >>
rect 190 5 191 6 
<< m2 >>
rect 190 5 191 6 
<< m1 >>
rect 191 5 192 6 
<< m2 >>
rect 191 5 192 6 
<< m1 >>
rect 192 5 193 6 
<< m2 >>
rect 192 5 193 6 
<< m1 >>
rect 193 5 194 6 
<< m2 >>
rect 193 5 194 6 
<< m1 >>
rect 194 5 195 6 
<< m2 >>
rect 194 5 195 6 
<< m1 >>
rect 195 5 196 6 
<< m2 >>
rect 195 5 196 6 
<< m1 >>
rect 196 5 197 6 
<< m2 >>
rect 196 5 197 6 
<< m1 >>
rect 197 5 198 6 
<< m1 >>
rect 198 5 199 6 
<< m1 >>
rect 199 5 200 6 
<< m2 >>
rect 199 5 200 6 
<< m2c >>
rect 199 5 200 6 
<< m1 >>
rect 199 5 200 6 
<< m2 >>
rect 199 5 200 6 
<< m1 >>
rect 201 5 202 6 
<< m2 >>
rect 201 5 202 6 
<< m2c >>
rect 201 5 202 6 
<< m1 >>
rect 201 5 202 6 
<< m2 >>
rect 201 5 202 6 
<< m1 >>
rect 37 6 38 7 
<< m2 >>
rect 49 6 50 7 
<< m1 >>
rect 58 6 59 7 
<< m2 >>
rect 130 6 131 7 
<< m2 >>
rect 146 6 147 7 
<< m2 >>
rect 196 6 197 7 
<< m2 >>
rect 199 6 200 7 
<< m2 >>
rect 201 6 202 7 
<< m1 >>
rect 37 7 38 8 
<< m1 >>
rect 40 7 41 8 
<< m1 >>
rect 41 7 42 8 
<< m1 >>
rect 42 7 43 8 
<< m1 >>
rect 43 7 44 8 
<< m1 >>
rect 44 7 45 8 
<< m1 >>
rect 45 7 46 8 
<< m1 >>
rect 46 7 47 8 
<< m1 >>
rect 47 7 48 8 
<< m1 >>
rect 48 7 49 8 
<< m1 >>
rect 49 7 50 8 
<< m2 >>
rect 49 7 50 8 
<< m1 >>
rect 50 7 51 8 
<< m1 >>
rect 51 7 52 8 
<< m1 >>
rect 52 7 53 8 
<< m1 >>
rect 53 7 54 8 
<< m1 >>
rect 54 7 55 8 
<< m1 >>
rect 55 7 56 8 
<< m1 >>
rect 56 7 57 8 
<< m2 >>
rect 56 7 57 8 
<< m2c >>
rect 56 7 57 8 
<< m1 >>
rect 56 7 57 8 
<< m2 >>
rect 56 7 57 8 
<< m2 >>
rect 57 7 58 8 
<< m1 >>
rect 58 7 59 8 
<< m2 >>
rect 58 7 59 8 
<< m2 >>
rect 59 7 60 8 
<< m1 >>
rect 60 7 61 8 
<< m2 >>
rect 60 7 61 8 
<< m1 >>
rect 61 7 62 8 
<< m2 >>
rect 61 7 62 8 
<< m1 >>
rect 62 7 63 8 
<< m2 >>
rect 62 7 63 8 
<< m1 >>
rect 63 7 64 8 
<< m2 >>
rect 63 7 64 8 
<< m1 >>
rect 64 7 65 8 
<< m2 >>
rect 64 7 65 8 
<< m1 >>
rect 65 7 66 8 
<< m2 >>
rect 65 7 66 8 
<< m1 >>
rect 66 7 67 8 
<< m2 >>
rect 66 7 67 8 
<< m1 >>
rect 67 7 68 8 
<< m2 >>
rect 67 7 68 8 
<< m1 >>
rect 68 7 69 8 
<< m2 >>
rect 68 7 69 8 
<< m1 >>
rect 69 7 70 8 
<< m2 >>
rect 69 7 70 8 
<< m1 >>
rect 70 7 71 8 
<< m2 >>
rect 70 7 71 8 
<< m1 >>
rect 71 7 72 8 
<< m2 >>
rect 71 7 72 8 
<< m1 >>
rect 72 7 73 8 
<< m2 >>
rect 72 7 73 8 
<< m1 >>
rect 73 7 74 8 
<< m2 >>
rect 73 7 74 8 
<< m1 >>
rect 74 7 75 8 
<< m2 >>
rect 74 7 75 8 
<< m1 >>
rect 75 7 76 8 
<< m2 >>
rect 75 7 76 8 
<< m1 >>
rect 76 7 77 8 
<< m2 >>
rect 76 7 77 8 
<< m1 >>
rect 77 7 78 8 
<< m2 >>
rect 77 7 78 8 
<< m1 >>
rect 78 7 79 8 
<< m2 >>
rect 78 7 79 8 
<< m1 >>
rect 79 7 80 8 
<< m2 >>
rect 79 7 80 8 
<< m1 >>
rect 80 7 81 8 
<< m2 >>
rect 80 7 81 8 
<< m1 >>
rect 81 7 82 8 
<< m2 >>
rect 81 7 82 8 
<< m1 >>
rect 82 7 83 8 
<< m2 >>
rect 82 7 83 8 
<< m1 >>
rect 83 7 84 8 
<< m2 >>
rect 83 7 84 8 
<< m1 >>
rect 84 7 85 8 
<< m2 >>
rect 84 7 85 8 
<< m1 >>
rect 85 7 86 8 
<< m2 >>
rect 85 7 86 8 
<< m1 >>
rect 86 7 87 8 
<< m2 >>
rect 86 7 87 8 
<< m1 >>
rect 87 7 88 8 
<< m2 >>
rect 87 7 88 8 
<< m1 >>
rect 88 7 89 8 
<< m2 >>
rect 88 7 89 8 
<< m1 >>
rect 89 7 90 8 
<< m2 >>
rect 89 7 90 8 
<< m1 >>
rect 90 7 91 8 
<< m2 >>
rect 90 7 91 8 
<< m1 >>
rect 91 7 92 8 
<< m2 >>
rect 91 7 92 8 
<< m1 >>
rect 92 7 93 8 
<< m2 >>
rect 92 7 93 8 
<< m1 >>
rect 93 7 94 8 
<< m2 >>
rect 93 7 94 8 
<< m1 >>
rect 94 7 95 8 
<< m2 >>
rect 94 7 95 8 
<< m1 >>
rect 95 7 96 8 
<< m2 >>
rect 95 7 96 8 
<< m1 >>
rect 96 7 97 8 
<< m2 >>
rect 96 7 97 8 
<< m1 >>
rect 97 7 98 8 
<< m2 >>
rect 97 7 98 8 
<< m1 >>
rect 98 7 99 8 
<< m2 >>
rect 98 7 99 8 
<< m1 >>
rect 99 7 100 8 
<< m2 >>
rect 99 7 100 8 
<< m1 >>
rect 100 7 101 8 
<< m2 >>
rect 100 7 101 8 
<< m1 >>
rect 101 7 102 8 
<< m2 >>
rect 101 7 102 8 
<< m1 >>
rect 102 7 103 8 
<< m2 >>
rect 102 7 103 8 
<< m1 >>
rect 103 7 104 8 
<< m2 >>
rect 103 7 104 8 
<< m1 >>
rect 104 7 105 8 
<< m2 >>
rect 104 7 105 8 
<< m1 >>
rect 105 7 106 8 
<< m2 >>
rect 105 7 106 8 
<< m1 >>
rect 106 7 107 8 
<< m2 >>
rect 106 7 107 8 
<< m1 >>
rect 107 7 108 8 
<< m2 >>
rect 107 7 108 8 
<< m1 >>
rect 108 7 109 8 
<< m2 >>
rect 108 7 109 8 
<< m1 >>
rect 109 7 110 8 
<< m2 >>
rect 109 7 110 8 
<< m1 >>
rect 110 7 111 8 
<< m2 >>
rect 110 7 111 8 
<< m1 >>
rect 111 7 112 8 
<< m2 >>
rect 111 7 112 8 
<< m1 >>
rect 112 7 113 8 
<< m2 >>
rect 112 7 113 8 
<< m1 >>
rect 113 7 114 8 
<< m2 >>
rect 113 7 114 8 
<< m1 >>
rect 114 7 115 8 
<< m2 >>
rect 114 7 115 8 
<< m1 >>
rect 115 7 116 8 
<< m2 >>
rect 115 7 116 8 
<< m1 >>
rect 116 7 117 8 
<< m2 >>
rect 116 7 117 8 
<< m1 >>
rect 117 7 118 8 
<< m2 >>
rect 117 7 118 8 
<< m1 >>
rect 118 7 119 8 
<< m2 >>
rect 118 7 119 8 
<< m1 >>
rect 119 7 120 8 
<< m2 >>
rect 119 7 120 8 
<< m1 >>
rect 120 7 121 8 
<< m2 >>
rect 120 7 121 8 
<< m1 >>
rect 121 7 122 8 
<< m2 >>
rect 121 7 122 8 
<< m1 >>
rect 122 7 123 8 
<< m2 >>
rect 122 7 123 8 
<< m1 >>
rect 123 7 124 8 
<< m2 >>
rect 123 7 124 8 
<< m1 >>
rect 124 7 125 8 
<< m2 >>
rect 124 7 125 8 
<< m1 >>
rect 125 7 126 8 
<< m2 >>
rect 125 7 126 8 
<< m1 >>
rect 126 7 127 8 
<< m2 >>
rect 126 7 127 8 
<< m1 >>
rect 127 7 128 8 
<< m2 >>
rect 127 7 128 8 
<< m1 >>
rect 128 7 129 8 
<< m2 >>
rect 128 7 129 8 
<< m1 >>
rect 129 7 130 8 
<< m1 >>
rect 130 7 131 8 
<< m2 >>
rect 130 7 131 8 
<< m1 >>
rect 131 7 132 8 
<< m1 >>
rect 132 7 133 8 
<< m1 >>
rect 133 7 134 8 
<< m1 >>
rect 134 7 135 8 
<< m1 >>
rect 135 7 136 8 
<< m1 >>
rect 136 7 137 8 
<< m1 >>
rect 137 7 138 8 
<< m1 >>
rect 138 7 139 8 
<< m1 >>
rect 139 7 140 8 
<< m1 >>
rect 140 7 141 8 
<< m1 >>
rect 141 7 142 8 
<< m1 >>
rect 142 7 143 8 
<< m1 >>
rect 143 7 144 8 
<< m1 >>
rect 144 7 145 8 
<< m1 >>
rect 145 7 146 8 
<< m1 >>
rect 146 7 147 8 
<< m2 >>
rect 146 7 147 8 
<< m1 >>
rect 147 7 148 8 
<< m1 >>
rect 148 7 149 8 
<< m2 >>
rect 148 7 149 8 
<< m2c >>
rect 148 7 149 8 
<< m1 >>
rect 148 7 149 8 
<< m2 >>
rect 148 7 149 8 
<< m2 >>
rect 149 7 150 8 
<< m1 >>
rect 150 7 151 8 
<< m2 >>
rect 150 7 151 8 
<< m1 >>
rect 151 7 152 8 
<< m2 >>
rect 151 7 152 8 
<< m1 >>
rect 152 7 153 8 
<< m2 >>
rect 152 7 153 8 
<< m1 >>
rect 153 7 154 8 
<< m2 >>
rect 153 7 154 8 
<< m1 >>
rect 154 7 155 8 
<< m2 >>
rect 154 7 155 8 
<< m1 >>
rect 155 7 156 8 
<< m2 >>
rect 155 7 156 8 
<< m1 >>
rect 156 7 157 8 
<< m2 >>
rect 156 7 157 8 
<< m1 >>
rect 157 7 158 8 
<< m2 >>
rect 157 7 158 8 
<< m1 >>
rect 158 7 159 8 
<< m2 >>
rect 158 7 159 8 
<< m1 >>
rect 159 7 160 8 
<< m1 >>
rect 160 7 161 8 
<< m1 >>
rect 161 7 162 8 
<< m1 >>
rect 162 7 163 8 
<< m1 >>
rect 163 7 164 8 
<< m1 >>
rect 164 7 165 8 
<< m1 >>
rect 165 7 166 8 
<< m1 >>
rect 166 7 167 8 
<< m1 >>
rect 167 7 168 8 
<< m1 >>
rect 168 7 169 8 
<< m1 >>
rect 169 7 170 8 
<< m1 >>
rect 170 7 171 8 
<< m1 >>
rect 171 7 172 8 
<< m1 >>
rect 172 7 173 8 
<< m1 >>
rect 173 7 174 8 
<< m1 >>
rect 174 7 175 8 
<< m1 >>
rect 175 7 176 8 
<< m1 >>
rect 176 7 177 8 
<< m1 >>
rect 177 7 178 8 
<< m1 >>
rect 178 7 179 8 
<< m1 >>
rect 179 7 180 8 
<< m1 >>
rect 180 7 181 8 
<< m1 >>
rect 181 7 182 8 
<< m1 >>
rect 182 7 183 8 
<< m1 >>
rect 183 7 184 8 
<< m1 >>
rect 184 7 185 8 
<< m1 >>
rect 185 7 186 8 
<< m1 >>
rect 186 7 187 8 
<< m1 >>
rect 187 7 188 8 
<< m1 >>
rect 188 7 189 8 
<< m1 >>
rect 189 7 190 8 
<< m1 >>
rect 190 7 191 8 
<< m1 >>
rect 191 7 192 8 
<< m1 >>
rect 192 7 193 8 
<< m1 >>
rect 193 7 194 8 
<< m1 >>
rect 194 7 195 8 
<< m1 >>
rect 195 7 196 8 
<< m1 >>
rect 196 7 197 8 
<< m2 >>
rect 196 7 197 8 
<< m1 >>
rect 197 7 198 8 
<< m1 >>
rect 198 7 199 8 
<< m1 >>
rect 199 7 200 8 
<< m2 >>
rect 199 7 200 8 
<< m1 >>
rect 200 7 201 8 
<< m1 >>
rect 201 7 202 8 
<< m2 >>
rect 201 7 202 8 
<< m1 >>
rect 202 7 203 8 
<< m1 >>
rect 203 7 204 8 
<< m1 >>
rect 204 7 205 8 
<< m1 >>
rect 205 7 206 8 
<< m1 >>
rect 206 7 207 8 
<< m1 >>
rect 207 7 208 8 
<< m1 >>
rect 208 7 209 8 
<< m1 >>
rect 209 7 210 8 
<< m1 >>
rect 210 7 211 8 
<< m1 >>
rect 211 7 212 8 
<< m1 >>
rect 212 7 213 8 
<< m1 >>
rect 213 7 214 8 
<< m1 >>
rect 214 7 215 8 
<< m1 >>
rect 37 8 38 9 
<< m1 >>
rect 40 8 41 9 
<< m2 >>
rect 49 8 50 9 
<< m1 >>
rect 58 8 59 9 
<< m1 >>
rect 60 8 61 9 
<< m2 >>
rect 128 8 129 9 
<< m2 >>
rect 130 8 131 9 
<< m2 >>
rect 146 8 147 9 
<< m1 >>
rect 150 8 151 9 
<< m2 >>
rect 158 8 159 9 
<< m2 >>
rect 196 8 197 9 
<< m2 >>
rect 199 8 200 9 
<< m2 >>
rect 201 8 202 9 
<< m1 >>
rect 214 8 215 9 
<< m1 >>
rect 37 9 38 10 
<< m1 >>
rect 40 9 41 10 
<< m1 >>
rect 49 9 50 10 
<< m2 >>
rect 49 9 50 10 
<< m2c >>
rect 49 9 50 10 
<< m1 >>
rect 49 9 50 10 
<< m2 >>
rect 49 9 50 10 
<< m1 >>
rect 58 9 59 10 
<< m1 >>
rect 60 9 61 10 
<< m2 >>
rect 69 9 70 10 
<< m2 >>
rect 70 9 71 10 
<< m2 >>
rect 71 9 72 10 
<< m2 >>
rect 72 9 73 10 
<< m2 >>
rect 73 9 74 10 
<< m1 >>
rect 128 9 129 10 
<< m2 >>
rect 128 9 129 10 
<< m2c >>
rect 128 9 129 10 
<< m1 >>
rect 128 9 129 10 
<< m2 >>
rect 128 9 129 10 
<< m1 >>
rect 130 9 131 10 
<< m2 >>
rect 130 9 131 10 
<< m2c >>
rect 130 9 131 10 
<< m1 >>
rect 130 9 131 10 
<< m2 >>
rect 130 9 131 10 
<< m1 >>
rect 146 9 147 10 
<< m2 >>
rect 146 9 147 10 
<< m2c >>
rect 146 9 147 10 
<< m1 >>
rect 146 9 147 10 
<< m2 >>
rect 146 9 147 10 
<< m1 >>
rect 150 9 151 10 
<< m2 >>
rect 158 9 159 10 
<< m1 >>
rect 159 9 160 10 
<< m2 >>
rect 159 9 160 10 
<< m2c >>
rect 159 9 160 10 
<< m1 >>
rect 159 9 160 10 
<< m2 >>
rect 159 9 160 10 
<< m1 >>
rect 160 9 161 10 
<< m1 >>
rect 161 9 162 10 
<< m1 >>
rect 162 9 163 10 
<< m1 >>
rect 163 9 164 10 
<< m1 >>
rect 175 9 176 10 
<< m1 >>
rect 176 9 177 10 
<< m1 >>
rect 177 9 178 10 
<< m1 >>
rect 178 9 179 10 
<< m1 >>
rect 179 9 180 10 
<< m1 >>
rect 180 9 181 10 
<< m1 >>
rect 181 9 182 10 
<< m1 >>
rect 182 9 183 10 
<< m1 >>
rect 183 9 184 10 
<< m1 >>
rect 184 9 185 10 
<< m1 >>
rect 185 9 186 10 
<< m1 >>
rect 186 9 187 10 
<< m1 >>
rect 187 9 188 10 
<< m1 >>
rect 188 9 189 10 
<< m1 >>
rect 189 9 190 10 
<< m1 >>
rect 190 9 191 10 
<< m1 >>
rect 196 9 197 10 
<< m2 >>
rect 196 9 197 10 
<< m2c >>
rect 196 9 197 10 
<< m1 >>
rect 196 9 197 10 
<< m2 >>
rect 196 9 197 10 
<< m1 >>
rect 199 9 200 10 
<< m2 >>
rect 199 9 200 10 
<< m2c >>
rect 199 9 200 10 
<< m1 >>
rect 199 9 200 10 
<< m2 >>
rect 199 9 200 10 
<< m1 >>
rect 201 9 202 10 
<< m2 >>
rect 201 9 202 10 
<< m2c >>
rect 201 9 202 10 
<< m1 >>
rect 201 9 202 10 
<< m2 >>
rect 201 9 202 10 
<< m1 >>
rect 214 9 215 10 
<< m1 >>
rect 37 10 38 11 
<< m1 >>
rect 40 10 41 11 
<< m1 >>
rect 49 10 50 11 
<< m1 >>
rect 58 10 59 11 
<< m1 >>
rect 60 10 61 11 
<< m1 >>
rect 67 10 68 11 
<< m1 >>
rect 68 10 69 11 
<< m2 >>
rect 68 10 69 11 
<< m2c >>
rect 68 10 69 11 
<< m1 >>
rect 68 10 69 11 
<< m2 >>
rect 68 10 69 11 
<< m2 >>
rect 69 10 70 11 
<< m1 >>
rect 70 10 71 11 
<< m1 >>
rect 71 10 72 11 
<< m1 >>
rect 72 10 73 11 
<< m1 >>
rect 73 10 74 11 
<< m2 >>
rect 73 10 74 11 
<< m1 >>
rect 118 10 119 11 
<< m1 >>
rect 119 10 120 11 
<< m1 >>
rect 120 10 121 11 
<< m1 >>
rect 121 10 122 11 
<< m1 >>
rect 128 10 129 11 
<< m1 >>
rect 130 10 131 11 
<< m1 >>
rect 146 10 147 11 
<< m1 >>
rect 150 10 151 11 
<< m1 >>
rect 154 10 155 11 
<< m1 >>
rect 155 10 156 11 
<< m1 >>
rect 156 10 157 11 
<< m1 >>
rect 157 10 158 11 
<< m1 >>
rect 163 10 164 11 
<< m1 >>
rect 175 10 176 11 
<< m2 >>
rect 181 10 182 11 
<< m2 >>
rect 182 10 183 11 
<< m2 >>
rect 183 10 184 11 
<< m2 >>
rect 184 10 185 11 
<< m2 >>
rect 185 10 186 11 
<< m2 >>
rect 186 10 187 11 
<< m2 >>
rect 187 10 188 11 
<< m2 >>
rect 188 10 189 11 
<< m2 >>
rect 189 10 190 11 
<< m1 >>
rect 190 10 191 11 
<< m2 >>
rect 190 10 191 11 
<< m2 >>
rect 191 10 192 11 
<< m1 >>
rect 192 10 193 11 
<< m2 >>
rect 192 10 193 11 
<< m2c >>
rect 192 10 193 11 
<< m1 >>
rect 192 10 193 11 
<< m2 >>
rect 192 10 193 11 
<< m1 >>
rect 193 10 194 11 
<< m1 >>
rect 196 10 197 11 
<< m1 >>
rect 199 10 200 11 
<< m1 >>
rect 201 10 202 11 
<< m1 >>
rect 214 10 215 11 
<< m1 >>
rect 37 11 38 12 
<< m1 >>
rect 40 11 41 12 
<< m1 >>
rect 49 11 50 12 
<< m1 >>
rect 58 11 59 12 
<< m1 >>
rect 60 11 61 12 
<< m1 >>
rect 67 11 68 12 
<< m1 >>
rect 70 11 71 12 
<< m1 >>
rect 73 11 74 12 
<< m2 >>
rect 73 11 74 12 
<< m1 >>
rect 118 11 119 12 
<< m1 >>
rect 121 11 122 12 
<< m1 >>
rect 128 11 129 12 
<< m2 >>
rect 129 11 130 12 
<< m1 >>
rect 130 11 131 12 
<< m2 >>
rect 130 11 131 12 
<< m2c >>
rect 130 11 131 12 
<< m1 >>
rect 130 11 131 12 
<< m2 >>
rect 130 11 131 12 
<< m1 >>
rect 146 11 147 12 
<< m1 >>
rect 150 11 151 12 
<< m1 >>
rect 154 11 155 12 
<< m1 >>
rect 157 11 158 12 
<< m1 >>
rect 163 11 164 12 
<< m1 >>
rect 175 11 176 12 
<< m1 >>
rect 181 11 182 12 
<< m2 >>
rect 181 11 182 12 
<< m2c >>
rect 181 11 182 12 
<< m1 >>
rect 181 11 182 12 
<< m2 >>
rect 181 11 182 12 
<< m1 >>
rect 190 11 191 12 
<< m1 >>
rect 193 11 194 12 
<< m1 >>
rect 196 11 197 12 
<< m1 >>
rect 199 11 200 12 
<< m1 >>
rect 201 11 202 12 
<< m1 >>
rect 214 11 215 12 
<< pdiffusion >>
rect 12 12 13 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< pdiffusion >>
rect 30 12 31 13 
<< pdiffusion >>
rect 31 12 32 13 
<< pdiffusion >>
rect 32 12 33 13 
<< pdiffusion >>
rect 33 12 34 13 
<< pdiffusion >>
rect 34 12 35 13 
<< pdiffusion >>
rect 35 12 36 13 
<< m1 >>
rect 37 12 38 13 
<< m1 >>
rect 40 12 41 13 
<< pdiffusion >>
rect 48 12 49 13 
<< m1 >>
rect 49 12 50 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< pdiffusion >>
rect 51 12 52 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< m1 >>
rect 58 12 59 13 
<< m1 >>
rect 60 12 61 13 
<< pdiffusion >>
rect 66 12 67 13 
<< m1 >>
rect 67 12 68 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< m1 >>
rect 70 12 71 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< m1 >>
rect 73 12 74 13 
<< m2 >>
rect 73 12 74 13 
<< pdiffusion >>
rect 84 12 85 13 
<< pdiffusion >>
rect 85 12 86 13 
<< pdiffusion >>
rect 86 12 87 13 
<< pdiffusion >>
rect 87 12 88 13 
<< pdiffusion >>
rect 88 12 89 13 
<< pdiffusion >>
rect 89 12 90 13 
<< pdiffusion >>
rect 102 12 103 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< m1 >>
rect 118 12 119 13 
<< pdiffusion >>
rect 120 12 121 13 
<< m1 >>
rect 121 12 122 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< m1 >>
rect 128 12 129 13 
<< m2 >>
rect 129 12 130 13 
<< pdiffusion >>
rect 138 12 139 13 
<< pdiffusion >>
rect 139 12 140 13 
<< pdiffusion >>
rect 140 12 141 13 
<< pdiffusion >>
rect 141 12 142 13 
<< pdiffusion >>
rect 142 12 143 13 
<< pdiffusion >>
rect 143 12 144 13 
<< m1 >>
rect 146 12 147 13 
<< m1 >>
rect 150 12 151 13 
<< m1 >>
rect 154 12 155 13 
<< pdiffusion >>
rect 156 12 157 13 
<< m1 >>
rect 157 12 158 13 
<< pdiffusion >>
rect 157 12 158 13 
<< pdiffusion >>
rect 158 12 159 13 
<< pdiffusion >>
rect 159 12 160 13 
<< pdiffusion >>
rect 160 12 161 13 
<< pdiffusion >>
rect 161 12 162 13 
<< m1 >>
rect 163 12 164 13 
<< pdiffusion >>
rect 174 12 175 13 
<< m1 >>
rect 175 12 176 13 
<< pdiffusion >>
rect 175 12 176 13 
<< pdiffusion >>
rect 176 12 177 13 
<< pdiffusion >>
rect 177 12 178 13 
<< pdiffusion >>
rect 178 12 179 13 
<< pdiffusion >>
rect 179 12 180 13 
<< m1 >>
rect 181 12 182 13 
<< m1 >>
rect 190 12 191 13 
<< pdiffusion >>
rect 192 12 193 13 
<< m1 >>
rect 193 12 194 13 
<< pdiffusion >>
rect 193 12 194 13 
<< pdiffusion >>
rect 194 12 195 13 
<< pdiffusion >>
rect 195 12 196 13 
<< m1 >>
rect 196 12 197 13 
<< pdiffusion >>
rect 196 12 197 13 
<< pdiffusion >>
rect 197 12 198 13 
<< m1 >>
rect 199 12 200 13 
<< m1 >>
rect 201 12 202 13 
<< pdiffusion >>
rect 210 12 211 13 
<< pdiffusion >>
rect 211 12 212 13 
<< pdiffusion >>
rect 212 12 213 13 
<< pdiffusion >>
rect 213 12 214 13 
<< m1 >>
rect 214 12 215 13 
<< pdiffusion >>
rect 214 12 215 13 
<< pdiffusion >>
rect 215 12 216 13 
<< pdiffusion >>
rect 228 12 229 13 
<< pdiffusion >>
rect 229 12 230 13 
<< pdiffusion >>
rect 230 12 231 13 
<< pdiffusion >>
rect 231 12 232 13 
<< pdiffusion >>
rect 232 12 233 13 
<< pdiffusion >>
rect 233 12 234 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< pdiffusion >>
rect 30 13 31 14 
<< pdiffusion >>
rect 31 13 32 14 
<< pdiffusion >>
rect 32 13 33 14 
<< pdiffusion >>
rect 33 13 34 14 
<< pdiffusion >>
rect 34 13 35 14 
<< pdiffusion >>
rect 35 13 36 14 
<< m1 >>
rect 37 13 38 14 
<< m1 >>
rect 40 13 41 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< m1 >>
rect 58 13 59 14 
<< m1 >>
rect 60 13 61 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< m1 >>
rect 73 13 74 14 
<< m2 >>
rect 73 13 74 14 
<< pdiffusion >>
rect 84 13 85 14 
<< pdiffusion >>
rect 85 13 86 14 
<< pdiffusion >>
rect 86 13 87 14 
<< pdiffusion >>
rect 87 13 88 14 
<< pdiffusion >>
rect 88 13 89 14 
<< pdiffusion >>
rect 89 13 90 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< m1 >>
rect 118 13 119 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< m1 >>
rect 128 13 129 14 
<< m2 >>
rect 129 13 130 14 
<< pdiffusion >>
rect 138 13 139 14 
<< pdiffusion >>
rect 139 13 140 14 
<< pdiffusion >>
rect 140 13 141 14 
<< pdiffusion >>
rect 141 13 142 14 
<< pdiffusion >>
rect 142 13 143 14 
<< pdiffusion >>
rect 143 13 144 14 
<< m1 >>
rect 146 13 147 14 
<< m1 >>
rect 150 13 151 14 
<< m1 >>
rect 154 13 155 14 
<< pdiffusion >>
rect 156 13 157 14 
<< pdiffusion >>
rect 157 13 158 14 
<< pdiffusion >>
rect 158 13 159 14 
<< pdiffusion >>
rect 159 13 160 14 
<< pdiffusion >>
rect 160 13 161 14 
<< pdiffusion >>
rect 161 13 162 14 
<< m1 >>
rect 163 13 164 14 
<< pdiffusion >>
rect 174 13 175 14 
<< pdiffusion >>
rect 175 13 176 14 
<< pdiffusion >>
rect 176 13 177 14 
<< pdiffusion >>
rect 177 13 178 14 
<< pdiffusion >>
rect 178 13 179 14 
<< pdiffusion >>
rect 179 13 180 14 
<< m1 >>
rect 181 13 182 14 
<< m1 >>
rect 190 13 191 14 
<< pdiffusion >>
rect 192 13 193 14 
<< pdiffusion >>
rect 193 13 194 14 
<< pdiffusion >>
rect 194 13 195 14 
<< pdiffusion >>
rect 195 13 196 14 
<< pdiffusion >>
rect 196 13 197 14 
<< pdiffusion >>
rect 197 13 198 14 
<< m1 >>
rect 199 13 200 14 
<< m1 >>
rect 201 13 202 14 
<< pdiffusion >>
rect 210 13 211 14 
<< pdiffusion >>
rect 211 13 212 14 
<< pdiffusion >>
rect 212 13 213 14 
<< pdiffusion >>
rect 213 13 214 14 
<< pdiffusion >>
rect 214 13 215 14 
<< pdiffusion >>
rect 215 13 216 14 
<< pdiffusion >>
rect 228 13 229 14 
<< pdiffusion >>
rect 229 13 230 14 
<< pdiffusion >>
rect 230 13 231 14 
<< pdiffusion >>
rect 231 13 232 14 
<< pdiffusion >>
rect 232 13 233 14 
<< pdiffusion >>
rect 233 13 234 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< pdiffusion >>
rect 30 14 31 15 
<< pdiffusion >>
rect 31 14 32 15 
<< pdiffusion >>
rect 32 14 33 15 
<< pdiffusion >>
rect 33 14 34 15 
<< pdiffusion >>
rect 34 14 35 15 
<< pdiffusion >>
rect 35 14 36 15 
<< m1 >>
rect 37 14 38 15 
<< m1 >>
rect 40 14 41 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< m1 >>
rect 58 14 59 15 
<< m1 >>
rect 60 14 61 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< m1 >>
rect 73 14 74 15 
<< m2 >>
rect 73 14 74 15 
<< pdiffusion >>
rect 84 14 85 15 
<< pdiffusion >>
rect 85 14 86 15 
<< pdiffusion >>
rect 86 14 87 15 
<< pdiffusion >>
rect 87 14 88 15 
<< pdiffusion >>
rect 88 14 89 15 
<< pdiffusion >>
rect 89 14 90 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< m1 >>
rect 118 14 119 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< m1 >>
rect 128 14 129 15 
<< m2 >>
rect 129 14 130 15 
<< pdiffusion >>
rect 138 14 139 15 
<< pdiffusion >>
rect 139 14 140 15 
<< pdiffusion >>
rect 140 14 141 15 
<< pdiffusion >>
rect 141 14 142 15 
<< pdiffusion >>
rect 142 14 143 15 
<< pdiffusion >>
rect 143 14 144 15 
<< m1 >>
rect 146 14 147 15 
<< m1 >>
rect 150 14 151 15 
<< m1 >>
rect 154 14 155 15 
<< pdiffusion >>
rect 156 14 157 15 
<< pdiffusion >>
rect 157 14 158 15 
<< pdiffusion >>
rect 158 14 159 15 
<< pdiffusion >>
rect 159 14 160 15 
<< pdiffusion >>
rect 160 14 161 15 
<< pdiffusion >>
rect 161 14 162 15 
<< m1 >>
rect 163 14 164 15 
<< pdiffusion >>
rect 174 14 175 15 
<< pdiffusion >>
rect 175 14 176 15 
<< pdiffusion >>
rect 176 14 177 15 
<< pdiffusion >>
rect 177 14 178 15 
<< pdiffusion >>
rect 178 14 179 15 
<< pdiffusion >>
rect 179 14 180 15 
<< m1 >>
rect 181 14 182 15 
<< m1 >>
rect 190 14 191 15 
<< pdiffusion >>
rect 192 14 193 15 
<< pdiffusion >>
rect 193 14 194 15 
<< pdiffusion >>
rect 194 14 195 15 
<< pdiffusion >>
rect 195 14 196 15 
<< pdiffusion >>
rect 196 14 197 15 
<< pdiffusion >>
rect 197 14 198 15 
<< m1 >>
rect 199 14 200 15 
<< m1 >>
rect 201 14 202 15 
<< pdiffusion >>
rect 210 14 211 15 
<< pdiffusion >>
rect 211 14 212 15 
<< pdiffusion >>
rect 212 14 213 15 
<< pdiffusion >>
rect 213 14 214 15 
<< pdiffusion >>
rect 214 14 215 15 
<< pdiffusion >>
rect 215 14 216 15 
<< pdiffusion >>
rect 228 14 229 15 
<< pdiffusion >>
rect 229 14 230 15 
<< pdiffusion >>
rect 230 14 231 15 
<< pdiffusion >>
rect 231 14 232 15 
<< pdiffusion >>
rect 232 14 233 15 
<< pdiffusion >>
rect 233 14 234 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< pdiffusion >>
rect 30 15 31 16 
<< pdiffusion >>
rect 31 15 32 16 
<< pdiffusion >>
rect 32 15 33 16 
<< pdiffusion >>
rect 33 15 34 16 
<< pdiffusion >>
rect 34 15 35 16 
<< pdiffusion >>
rect 35 15 36 16 
<< m1 >>
rect 37 15 38 16 
<< m1 >>
rect 40 15 41 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< m1 >>
rect 58 15 59 16 
<< m1 >>
rect 60 15 61 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< m1 >>
rect 73 15 74 16 
<< m2 >>
rect 73 15 74 16 
<< pdiffusion >>
rect 84 15 85 16 
<< pdiffusion >>
rect 85 15 86 16 
<< pdiffusion >>
rect 86 15 87 16 
<< pdiffusion >>
rect 87 15 88 16 
<< pdiffusion >>
rect 88 15 89 16 
<< pdiffusion >>
rect 89 15 90 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< m1 >>
rect 118 15 119 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< m1 >>
rect 128 15 129 16 
<< m2 >>
rect 129 15 130 16 
<< pdiffusion >>
rect 138 15 139 16 
<< pdiffusion >>
rect 139 15 140 16 
<< pdiffusion >>
rect 140 15 141 16 
<< pdiffusion >>
rect 141 15 142 16 
<< pdiffusion >>
rect 142 15 143 16 
<< pdiffusion >>
rect 143 15 144 16 
<< m1 >>
rect 146 15 147 16 
<< m1 >>
rect 150 15 151 16 
<< m1 >>
rect 154 15 155 16 
<< pdiffusion >>
rect 156 15 157 16 
<< pdiffusion >>
rect 157 15 158 16 
<< pdiffusion >>
rect 158 15 159 16 
<< pdiffusion >>
rect 159 15 160 16 
<< pdiffusion >>
rect 160 15 161 16 
<< pdiffusion >>
rect 161 15 162 16 
<< m1 >>
rect 163 15 164 16 
<< pdiffusion >>
rect 174 15 175 16 
<< pdiffusion >>
rect 175 15 176 16 
<< pdiffusion >>
rect 176 15 177 16 
<< pdiffusion >>
rect 177 15 178 16 
<< pdiffusion >>
rect 178 15 179 16 
<< pdiffusion >>
rect 179 15 180 16 
<< m1 >>
rect 181 15 182 16 
<< m1 >>
rect 190 15 191 16 
<< pdiffusion >>
rect 192 15 193 16 
<< pdiffusion >>
rect 193 15 194 16 
<< pdiffusion >>
rect 194 15 195 16 
<< pdiffusion >>
rect 195 15 196 16 
<< pdiffusion >>
rect 196 15 197 16 
<< pdiffusion >>
rect 197 15 198 16 
<< m1 >>
rect 199 15 200 16 
<< m1 >>
rect 201 15 202 16 
<< pdiffusion >>
rect 210 15 211 16 
<< pdiffusion >>
rect 211 15 212 16 
<< pdiffusion >>
rect 212 15 213 16 
<< pdiffusion >>
rect 213 15 214 16 
<< pdiffusion >>
rect 214 15 215 16 
<< pdiffusion >>
rect 215 15 216 16 
<< pdiffusion >>
rect 228 15 229 16 
<< pdiffusion >>
rect 229 15 230 16 
<< pdiffusion >>
rect 230 15 231 16 
<< pdiffusion >>
rect 231 15 232 16 
<< pdiffusion >>
rect 232 15 233 16 
<< pdiffusion >>
rect 233 15 234 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< pdiffusion >>
rect 30 16 31 17 
<< pdiffusion >>
rect 31 16 32 17 
<< pdiffusion >>
rect 32 16 33 17 
<< pdiffusion >>
rect 33 16 34 17 
<< pdiffusion >>
rect 34 16 35 17 
<< pdiffusion >>
rect 35 16 36 17 
<< m1 >>
rect 37 16 38 17 
<< m1 >>
rect 40 16 41 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< m1 >>
rect 58 16 59 17 
<< m1 >>
rect 60 16 61 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< m1 >>
rect 73 16 74 17 
<< m2 >>
rect 73 16 74 17 
<< pdiffusion >>
rect 84 16 85 17 
<< pdiffusion >>
rect 85 16 86 17 
<< pdiffusion >>
rect 86 16 87 17 
<< pdiffusion >>
rect 87 16 88 17 
<< pdiffusion >>
rect 88 16 89 17 
<< pdiffusion >>
rect 89 16 90 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< m1 >>
rect 118 16 119 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< m1 >>
rect 128 16 129 17 
<< m2 >>
rect 129 16 130 17 
<< pdiffusion >>
rect 138 16 139 17 
<< pdiffusion >>
rect 139 16 140 17 
<< pdiffusion >>
rect 140 16 141 17 
<< pdiffusion >>
rect 141 16 142 17 
<< pdiffusion >>
rect 142 16 143 17 
<< pdiffusion >>
rect 143 16 144 17 
<< m1 >>
rect 146 16 147 17 
<< m1 >>
rect 150 16 151 17 
<< m1 >>
rect 154 16 155 17 
<< pdiffusion >>
rect 156 16 157 17 
<< pdiffusion >>
rect 157 16 158 17 
<< pdiffusion >>
rect 158 16 159 17 
<< pdiffusion >>
rect 159 16 160 17 
<< pdiffusion >>
rect 160 16 161 17 
<< pdiffusion >>
rect 161 16 162 17 
<< m1 >>
rect 163 16 164 17 
<< pdiffusion >>
rect 174 16 175 17 
<< pdiffusion >>
rect 175 16 176 17 
<< pdiffusion >>
rect 176 16 177 17 
<< pdiffusion >>
rect 177 16 178 17 
<< pdiffusion >>
rect 178 16 179 17 
<< pdiffusion >>
rect 179 16 180 17 
<< m1 >>
rect 181 16 182 17 
<< m1 >>
rect 190 16 191 17 
<< pdiffusion >>
rect 192 16 193 17 
<< pdiffusion >>
rect 193 16 194 17 
<< pdiffusion >>
rect 194 16 195 17 
<< pdiffusion >>
rect 195 16 196 17 
<< pdiffusion >>
rect 196 16 197 17 
<< pdiffusion >>
rect 197 16 198 17 
<< m1 >>
rect 199 16 200 17 
<< m1 >>
rect 201 16 202 17 
<< pdiffusion >>
rect 210 16 211 17 
<< pdiffusion >>
rect 211 16 212 17 
<< pdiffusion >>
rect 212 16 213 17 
<< pdiffusion >>
rect 213 16 214 17 
<< pdiffusion >>
rect 214 16 215 17 
<< pdiffusion >>
rect 215 16 216 17 
<< pdiffusion >>
rect 228 16 229 17 
<< pdiffusion >>
rect 229 16 230 17 
<< pdiffusion >>
rect 230 16 231 17 
<< pdiffusion >>
rect 231 16 232 17 
<< pdiffusion >>
rect 232 16 233 17 
<< pdiffusion >>
rect 233 16 234 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< pdiffusion >>
rect 30 17 31 18 
<< m1 >>
rect 31 17 32 18 
<< pdiffusion >>
rect 31 17 32 18 
<< pdiffusion >>
rect 32 17 33 18 
<< pdiffusion >>
rect 33 17 34 18 
<< pdiffusion >>
rect 34 17 35 18 
<< pdiffusion >>
rect 35 17 36 18 
<< m1 >>
rect 37 17 38 18 
<< m1 >>
rect 40 17 41 18 
<< pdiffusion >>
rect 48 17 49 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< m1 >>
rect 58 17 59 18 
<< m1 >>
rect 60 17 61 18 
<< pdiffusion >>
rect 66 17 67 18 
<< m1 >>
rect 67 17 68 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< m1 >>
rect 73 17 74 18 
<< m2 >>
rect 73 17 74 18 
<< pdiffusion >>
rect 84 17 85 18 
<< pdiffusion >>
rect 85 17 86 18 
<< pdiffusion >>
rect 86 17 87 18 
<< pdiffusion >>
rect 87 17 88 18 
<< m1 >>
rect 88 17 89 18 
<< pdiffusion >>
rect 88 17 89 18 
<< pdiffusion >>
rect 89 17 90 18 
<< pdiffusion >>
rect 102 17 103 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< m1 >>
rect 118 17 119 18 
<< pdiffusion >>
rect 120 17 121 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< m1 >>
rect 128 17 129 18 
<< m2 >>
rect 129 17 130 18 
<< pdiffusion >>
rect 138 17 139 18 
<< m1 >>
rect 139 17 140 18 
<< pdiffusion >>
rect 139 17 140 18 
<< pdiffusion >>
rect 140 17 141 18 
<< pdiffusion >>
rect 141 17 142 18 
<< pdiffusion >>
rect 142 17 143 18 
<< pdiffusion >>
rect 143 17 144 18 
<< m1 >>
rect 146 17 147 18 
<< m1 >>
rect 150 17 151 18 
<< m1 >>
rect 154 17 155 18 
<< pdiffusion >>
rect 156 17 157 18 
<< pdiffusion >>
rect 157 17 158 18 
<< pdiffusion >>
rect 158 17 159 18 
<< pdiffusion >>
rect 159 17 160 18 
<< pdiffusion >>
rect 160 17 161 18 
<< pdiffusion >>
rect 161 17 162 18 
<< m1 >>
rect 163 17 164 18 
<< pdiffusion >>
rect 174 17 175 18 
<< pdiffusion >>
rect 175 17 176 18 
<< pdiffusion >>
rect 176 17 177 18 
<< pdiffusion >>
rect 177 17 178 18 
<< pdiffusion >>
rect 178 17 179 18 
<< pdiffusion >>
rect 179 17 180 18 
<< m1 >>
rect 181 17 182 18 
<< m1 >>
rect 190 17 191 18 
<< pdiffusion >>
rect 192 17 193 18 
<< pdiffusion >>
rect 193 17 194 18 
<< pdiffusion >>
rect 194 17 195 18 
<< pdiffusion >>
rect 195 17 196 18 
<< m1 >>
rect 196 17 197 18 
<< pdiffusion >>
rect 196 17 197 18 
<< pdiffusion >>
rect 197 17 198 18 
<< m1 >>
rect 199 17 200 18 
<< m1 >>
rect 201 17 202 18 
<< pdiffusion >>
rect 210 17 211 18 
<< pdiffusion >>
rect 211 17 212 18 
<< pdiffusion >>
rect 212 17 213 18 
<< pdiffusion >>
rect 213 17 214 18 
<< pdiffusion >>
rect 214 17 215 18 
<< pdiffusion >>
rect 215 17 216 18 
<< pdiffusion >>
rect 228 17 229 18 
<< m1 >>
rect 229 17 230 18 
<< pdiffusion >>
rect 229 17 230 18 
<< pdiffusion >>
rect 230 17 231 18 
<< pdiffusion >>
rect 231 17 232 18 
<< m1 >>
rect 232 17 233 18 
<< pdiffusion >>
rect 232 17 233 18 
<< pdiffusion >>
rect 233 17 234 18 
<< m1 >>
rect 31 18 32 19 
<< m1 >>
rect 37 18 38 19 
<< m1 >>
rect 40 18 41 19 
<< m1 >>
rect 58 18 59 19 
<< m1 >>
rect 60 18 61 19 
<< m1 >>
rect 67 18 68 19 
<< m1 >>
rect 73 18 74 19 
<< m2 >>
rect 73 18 74 19 
<< m1 >>
rect 88 18 89 19 
<< m1 >>
rect 118 18 119 19 
<< m1 >>
rect 128 18 129 19 
<< m2 >>
rect 129 18 130 19 
<< m1 >>
rect 139 18 140 19 
<< m1 >>
rect 146 18 147 19 
<< m1 >>
rect 150 18 151 19 
<< m1 >>
rect 154 18 155 19 
<< m1 >>
rect 163 18 164 19 
<< m1 >>
rect 181 18 182 19 
<< m1 >>
rect 190 18 191 19 
<< m1 >>
rect 196 18 197 19 
<< m1 >>
rect 199 18 200 19 
<< m1 >>
rect 201 18 202 19 
<< m1 >>
rect 229 18 230 19 
<< m1 >>
rect 232 18 233 19 
<< m1 >>
rect 28 19 29 20 
<< m1 >>
rect 29 19 30 20 
<< m1 >>
rect 30 19 31 20 
<< m1 >>
rect 31 19 32 20 
<< m1 >>
rect 37 19 38 20 
<< m1 >>
rect 40 19 41 20 
<< m1 >>
rect 58 19 59 20 
<< m1 >>
rect 60 19 61 20 
<< m1 >>
rect 67 19 68 20 
<< m1 >>
rect 73 19 74 20 
<< m2 >>
rect 73 19 74 20 
<< m1 >>
rect 88 19 89 20 
<< m1 >>
rect 118 19 119 20 
<< m1 >>
rect 126 19 127 20 
<< m2 >>
rect 126 19 127 20 
<< m2c >>
rect 126 19 127 20 
<< m1 >>
rect 126 19 127 20 
<< m2 >>
rect 126 19 127 20 
<< m2 >>
rect 127 19 128 20 
<< m1 >>
rect 128 19 129 20 
<< m2 >>
rect 128 19 129 20 
<< m2 >>
rect 129 19 130 20 
<< m1 >>
rect 139 19 140 20 
<< m1 >>
rect 146 19 147 20 
<< m1 >>
rect 150 19 151 20 
<< m1 >>
rect 154 19 155 20 
<< m1 >>
rect 163 19 164 20 
<< m1 >>
rect 181 19 182 20 
<< m1 >>
rect 190 19 191 20 
<< m1 >>
rect 196 19 197 20 
<< m1 >>
rect 199 19 200 20 
<< m1 >>
rect 201 19 202 20 
<< m1 >>
rect 229 19 230 20 
<< m1 >>
rect 232 19 233 20 
<< m1 >>
rect 28 20 29 21 
<< m1 >>
rect 37 20 38 21 
<< m1 >>
rect 40 20 41 21 
<< m1 >>
rect 58 20 59 21 
<< m1 >>
rect 60 20 61 21 
<< m1 >>
rect 67 20 68 21 
<< m1 >>
rect 73 20 74 21 
<< m2 >>
rect 73 20 74 21 
<< m1 >>
rect 88 20 89 21 
<< m1 >>
rect 118 20 119 21 
<< m1 >>
rect 126 20 127 21 
<< m1 >>
rect 128 20 129 21 
<< m1 >>
rect 139 20 140 21 
<< m2 >>
rect 140 20 141 21 
<< m1 >>
rect 141 20 142 21 
<< m2 >>
rect 141 20 142 21 
<< m2c >>
rect 141 20 142 21 
<< m1 >>
rect 141 20 142 21 
<< m2 >>
rect 141 20 142 21 
<< m1 >>
rect 142 20 143 21 
<< m1 >>
rect 143 20 144 21 
<< m1 >>
rect 144 20 145 21 
<< m1 >>
rect 145 20 146 21 
<< m1 >>
rect 146 20 147 21 
<< m1 >>
rect 150 20 151 21 
<< m1 >>
rect 154 20 155 21 
<< m1 >>
rect 163 20 164 21 
<< m2 >>
rect 163 20 164 21 
<< m2c >>
rect 163 20 164 21 
<< m1 >>
rect 163 20 164 21 
<< m2 >>
rect 163 20 164 21 
<< m1 >>
rect 176 20 177 21 
<< m2 >>
rect 176 20 177 21 
<< m2c >>
rect 176 20 177 21 
<< m1 >>
rect 176 20 177 21 
<< m2 >>
rect 176 20 177 21 
<< m1 >>
rect 177 20 178 21 
<< m1 >>
rect 178 20 179 21 
<< m1 >>
rect 179 20 180 21 
<< m1 >>
rect 180 20 181 21 
<< m1 >>
rect 181 20 182 21 
<< m1 >>
rect 190 20 191 21 
<< m1 >>
rect 196 20 197 21 
<< m1 >>
rect 199 20 200 21 
<< m1 >>
rect 201 20 202 21 
<< m1 >>
rect 229 20 230 21 
<< m1 >>
rect 232 20 233 21 
<< m1 >>
rect 28 21 29 22 
<< m1 >>
rect 37 21 38 22 
<< m1 >>
rect 40 21 41 22 
<< m1 >>
rect 58 21 59 22 
<< m1 >>
rect 60 21 61 22 
<< m1 >>
rect 67 21 68 22 
<< m1 >>
rect 73 21 74 22 
<< m2 >>
rect 73 21 74 22 
<< m1 >>
rect 86 21 87 22 
<< m2 >>
rect 86 21 87 22 
<< m2c >>
rect 86 21 87 22 
<< m1 >>
rect 86 21 87 22 
<< m2 >>
rect 86 21 87 22 
<< m2 >>
rect 87 21 88 22 
<< m1 >>
rect 88 21 89 22 
<< m2 >>
rect 88 21 89 22 
<< m2 >>
rect 89 21 90 22 
<< m1 >>
rect 90 21 91 22 
<< m2 >>
rect 90 21 91 22 
<< m2c >>
rect 90 21 91 22 
<< m1 >>
rect 90 21 91 22 
<< m2 >>
rect 90 21 91 22 
<< m1 >>
rect 91 21 92 22 
<< m1 >>
rect 92 21 93 22 
<< m1 >>
rect 93 21 94 22 
<< m1 >>
rect 94 21 95 22 
<< m1 >>
rect 95 21 96 22 
<< m1 >>
rect 96 21 97 22 
<< m1 >>
rect 97 21 98 22 
<< m1 >>
rect 98 21 99 22 
<< m1 >>
rect 99 21 100 22 
<< m1 >>
rect 100 21 101 22 
<< m1 >>
rect 101 21 102 22 
<< m1 >>
rect 102 21 103 22 
<< m1 >>
rect 118 21 119 22 
<< m1 >>
rect 119 21 120 22 
<< m1 >>
rect 120 21 121 22 
<< m1 >>
rect 126 21 127 22 
<< m1 >>
rect 128 21 129 22 
<< m1 >>
rect 139 21 140 22 
<< m2 >>
rect 140 21 141 22 
<< m1 >>
rect 150 21 151 22 
<< m1 >>
rect 154 21 155 22 
<< m2 >>
rect 163 21 164 22 
<< m2 >>
rect 176 21 177 22 
<< m1 >>
rect 190 21 191 22 
<< m1 >>
rect 196 21 197 22 
<< m1 >>
rect 199 21 200 22 
<< m1 >>
rect 201 21 202 22 
<< m1 >>
rect 229 21 230 22 
<< m1 >>
rect 232 21 233 22 
<< m1 >>
rect 28 22 29 23 
<< m1 >>
rect 37 22 38 23 
<< m1 >>
rect 40 22 41 23 
<< m1 >>
rect 58 22 59 23 
<< m1 >>
rect 60 22 61 23 
<< m1 >>
rect 67 22 68 23 
<< m1 >>
rect 73 22 74 23 
<< m2 >>
rect 73 22 74 23 
<< m1 >>
rect 85 22 86 23 
<< m1 >>
rect 86 22 87 23 
<< m1 >>
rect 88 22 89 23 
<< m1 >>
rect 102 22 103 23 
<< m1 >>
rect 120 22 121 23 
<< m1 >>
rect 121 22 122 23 
<< m1 >>
rect 122 22 123 23 
<< m1 >>
rect 123 22 124 23 
<< m1 >>
rect 124 22 125 23 
<< m1 >>
rect 125 22 126 23 
<< m1 >>
rect 126 22 127 23 
<< m1 >>
rect 128 22 129 23 
<< m1 >>
rect 139 22 140 23 
<< m2 >>
rect 140 22 141 23 
<< m1 >>
rect 150 22 151 23 
<< m1 >>
rect 152 22 153 23 
<< m2 >>
rect 152 22 153 23 
<< m2c >>
rect 152 22 153 23 
<< m1 >>
rect 152 22 153 23 
<< m2 >>
rect 152 22 153 23 
<< m2 >>
rect 153 22 154 23 
<< m1 >>
rect 154 22 155 23 
<< m2 >>
rect 154 22 155 23 
<< m2 >>
rect 155 22 156 23 
<< m1 >>
rect 156 22 157 23 
<< m2 >>
rect 156 22 157 23 
<< m2c >>
rect 156 22 157 23 
<< m1 >>
rect 156 22 157 23 
<< m2 >>
rect 156 22 157 23 
<< m1 >>
rect 157 22 158 23 
<< m1 >>
rect 158 22 159 23 
<< m1 >>
rect 159 22 160 23 
<< m1 >>
rect 160 22 161 23 
<< m1 >>
rect 161 22 162 23 
<< m1 >>
rect 162 22 163 23 
<< m1 >>
rect 163 22 164 23 
<< m2 >>
rect 163 22 164 23 
<< m1 >>
rect 164 22 165 23 
<< m1 >>
rect 165 22 166 23 
<< m1 >>
rect 166 22 167 23 
<< m1 >>
rect 167 22 168 23 
<< m1 >>
rect 168 22 169 23 
<< m1 >>
rect 169 22 170 23 
<< m1 >>
rect 170 22 171 23 
<< m1 >>
rect 171 22 172 23 
<< m1 >>
rect 172 22 173 23 
<< m1 >>
rect 173 22 174 23 
<< m1 >>
rect 174 22 175 23 
<< m1 >>
rect 175 22 176 23 
<< m1 >>
rect 176 22 177 23 
<< m2 >>
rect 176 22 177 23 
<< m1 >>
rect 177 22 178 23 
<< m1 >>
rect 178 22 179 23 
<< m1 >>
rect 179 22 180 23 
<< m1 >>
rect 180 22 181 23 
<< m1 >>
rect 181 22 182 23 
<< m1 >>
rect 182 22 183 23 
<< m1 >>
rect 183 22 184 23 
<< m1 >>
rect 184 22 185 23 
<< m1 >>
rect 185 22 186 23 
<< m1 >>
rect 186 22 187 23 
<< m1 >>
rect 187 22 188 23 
<< m1 >>
rect 188 22 189 23 
<< m2 >>
rect 188 22 189 23 
<< m2c >>
rect 188 22 189 23 
<< m1 >>
rect 188 22 189 23 
<< m2 >>
rect 188 22 189 23 
<< m2 >>
rect 189 22 190 23 
<< m1 >>
rect 190 22 191 23 
<< m2 >>
rect 190 22 191 23 
<< m2 >>
rect 191 22 192 23 
<< m1 >>
rect 192 22 193 23 
<< m2 >>
rect 192 22 193 23 
<< m2c >>
rect 192 22 193 23 
<< m1 >>
rect 192 22 193 23 
<< m2 >>
rect 192 22 193 23 
<< m1 >>
rect 193 22 194 23 
<< m1 >>
rect 194 22 195 23 
<< m1 >>
rect 195 22 196 23 
<< m1 >>
rect 196 22 197 23 
<< m1 >>
rect 199 22 200 23 
<< m1 >>
rect 201 22 202 23 
<< m1 >>
rect 229 22 230 23 
<< m1 >>
rect 232 22 233 23 
<< m1 >>
rect 28 23 29 24 
<< m1 >>
rect 37 23 38 24 
<< m1 >>
rect 40 23 41 24 
<< m1 >>
rect 58 23 59 24 
<< m1 >>
rect 60 23 61 24 
<< m1 >>
rect 67 23 68 24 
<< m1 >>
rect 73 23 74 24 
<< m2 >>
rect 73 23 74 24 
<< m1 >>
rect 85 23 86 24 
<< m1 >>
rect 88 23 89 24 
<< m2 >>
rect 88 23 89 24 
<< m2c >>
rect 88 23 89 24 
<< m1 >>
rect 88 23 89 24 
<< m2 >>
rect 88 23 89 24 
<< m1 >>
rect 102 23 103 24 
<< m1 >>
rect 103 23 104 24 
<< m1 >>
rect 104 23 105 24 
<< m1 >>
rect 105 23 106 24 
<< m1 >>
rect 106 23 107 24 
<< m1 >>
rect 107 23 108 24 
<< m1 >>
rect 108 23 109 24 
<< m1 >>
rect 109 23 110 24 
<< m1 >>
rect 110 23 111 24 
<< m1 >>
rect 111 23 112 24 
<< m1 >>
rect 112 23 113 24 
<< m1 >>
rect 113 23 114 24 
<< m1 >>
rect 114 23 115 24 
<< m1 >>
rect 115 23 116 24 
<< m1 >>
rect 116 23 117 24 
<< m1 >>
rect 117 23 118 24 
<< m1 >>
rect 118 23 119 24 
<< m2 >>
rect 118 23 119 24 
<< m2c >>
rect 118 23 119 24 
<< m1 >>
rect 118 23 119 24 
<< m2 >>
rect 118 23 119 24 
<< m1 >>
rect 128 23 129 24 
<< m2 >>
rect 128 23 129 24 
<< m2c >>
rect 128 23 129 24 
<< m1 >>
rect 128 23 129 24 
<< m2 >>
rect 128 23 129 24 
<< m1 >>
rect 139 23 140 24 
<< m2 >>
rect 140 23 141 24 
<< m1 >>
rect 150 23 151 24 
<< m1 >>
rect 152 23 153 24 
<< m1 >>
rect 154 23 155 24 
<< m2 >>
rect 163 23 164 24 
<< m2 >>
rect 165 23 166 24 
<< m2 >>
rect 166 23 167 24 
<< m2 >>
rect 167 23 168 24 
<< m2 >>
rect 168 23 169 24 
<< m2 >>
rect 169 23 170 24 
<< m2 >>
rect 170 23 171 24 
<< m2 >>
rect 171 23 172 24 
<< m2 >>
rect 172 23 173 24 
<< m2 >>
rect 173 23 174 24 
<< m2 >>
rect 174 23 175 24 
<< m2 >>
rect 175 23 176 24 
<< m2 >>
rect 176 23 177 24 
<< m1 >>
rect 190 23 191 24 
<< m2 >>
rect 194 23 195 24 
<< m2 >>
rect 195 23 196 24 
<< m2 >>
rect 196 23 197 24 
<< m2 >>
rect 197 23 198 24 
<< m1 >>
rect 198 23 199 24 
<< m2 >>
rect 198 23 199 24 
<< m2c >>
rect 198 23 199 24 
<< m1 >>
rect 198 23 199 24 
<< m2 >>
rect 198 23 199 24 
<< m1 >>
rect 199 23 200 24 
<< m1 >>
rect 201 23 202 24 
<< m2 >>
rect 201 23 202 24 
<< m2c >>
rect 201 23 202 24 
<< m1 >>
rect 201 23 202 24 
<< m2 >>
rect 201 23 202 24 
<< m1 >>
rect 229 23 230 24 
<< m1 >>
rect 230 23 231 24 
<< m2 >>
rect 230 23 231 24 
<< m2c >>
rect 230 23 231 24 
<< m1 >>
rect 230 23 231 24 
<< m2 >>
rect 230 23 231 24 
<< m2 >>
rect 231 23 232 24 
<< m1 >>
rect 232 23 233 24 
<< m2 >>
rect 232 23 233 24 
<< m2 >>
rect 233 23 234 24 
<< m1 >>
rect 28 24 29 25 
<< m1 >>
rect 37 24 38 25 
<< m1 >>
rect 40 24 41 25 
<< m1 >>
rect 58 24 59 25 
<< m1 >>
rect 60 24 61 25 
<< m1 >>
rect 67 24 68 25 
<< m1 >>
rect 73 24 74 25 
<< m2 >>
rect 73 24 74 25 
<< m1 >>
rect 85 24 86 25 
<< m2 >>
rect 88 24 89 25 
<< m2 >>
rect 118 24 119 25 
<< m2 >>
rect 128 24 129 25 
<< m2 >>
rect 136 24 137 25 
<< m2 >>
rect 137 24 138 25 
<< m2 >>
rect 138 24 139 25 
<< m1 >>
rect 139 24 140 25 
<< m2 >>
rect 139 24 140 25 
<< m2 >>
rect 140 24 141 25 
<< m1 >>
rect 150 24 151 25 
<< m2 >>
rect 150 24 151 25 
<< m2c >>
rect 150 24 151 25 
<< m1 >>
rect 150 24 151 25 
<< m2 >>
rect 150 24 151 25 
<< m1 >>
rect 152 24 153 25 
<< m1 >>
rect 154 24 155 25 
<< m1 >>
rect 163 24 164 25 
<< m2 >>
rect 163 24 164 25 
<< m2c >>
rect 163 24 164 25 
<< m1 >>
rect 163 24 164 25 
<< m2 >>
rect 163 24 164 25 
<< m1 >>
rect 165 24 166 25 
<< m2 >>
rect 165 24 166 25 
<< m2c >>
rect 165 24 166 25 
<< m1 >>
rect 165 24 166 25 
<< m2 >>
rect 165 24 166 25 
<< m1 >>
rect 190 24 191 25 
<< m1 >>
rect 194 24 195 25 
<< m2 >>
rect 194 24 195 25 
<< m2c >>
rect 194 24 195 25 
<< m1 >>
rect 194 24 195 25 
<< m2 >>
rect 194 24 195 25 
<< m2 >>
rect 201 24 202 25 
<< m1 >>
rect 232 24 233 25 
<< m2 >>
rect 233 24 234 25 
<< m1 >>
rect 28 25 29 26 
<< m1 >>
rect 37 25 38 26 
<< m1 >>
rect 40 25 41 26 
<< m1 >>
rect 58 25 59 26 
<< m1 >>
rect 60 25 61 26 
<< m1 >>
rect 67 25 68 26 
<< m1 >>
rect 73 25 74 26 
<< m2 >>
rect 73 25 74 26 
<< m1 >>
rect 85 25 86 26 
<< m1 >>
rect 88 25 89 26 
<< m2 >>
rect 88 25 89 26 
<< m1 >>
rect 89 25 90 26 
<< m1 >>
rect 90 25 91 26 
<< m1 >>
rect 91 25 92 26 
<< m1 >>
rect 92 25 93 26 
<< m1 >>
rect 93 25 94 26 
<< m1 >>
rect 94 25 95 26 
<< m1 >>
rect 95 25 96 26 
<< m1 >>
rect 96 25 97 26 
<< m1 >>
rect 97 25 98 26 
<< m1 >>
rect 98 25 99 26 
<< m1 >>
rect 99 25 100 26 
<< m1 >>
rect 100 25 101 26 
<< m1 >>
rect 101 25 102 26 
<< m1 >>
rect 102 25 103 26 
<< m1 >>
rect 103 25 104 26 
<< m1 >>
rect 104 25 105 26 
<< m1 >>
rect 105 25 106 26 
<< m1 >>
rect 106 25 107 26 
<< m1 >>
rect 107 25 108 26 
<< m1 >>
rect 108 25 109 26 
<< m1 >>
rect 109 25 110 26 
<< m1 >>
rect 110 25 111 26 
<< m1 >>
rect 111 25 112 26 
<< m1 >>
rect 112 25 113 26 
<< m1 >>
rect 113 25 114 26 
<< m1 >>
rect 114 25 115 26 
<< m1 >>
rect 115 25 116 26 
<< m1 >>
rect 116 25 117 26 
<< m1 >>
rect 117 25 118 26 
<< m1 >>
rect 118 25 119 26 
<< m2 >>
rect 118 25 119 26 
<< m1 >>
rect 119 25 120 26 
<< m1 >>
rect 120 25 121 26 
<< m1 >>
rect 121 25 122 26 
<< m1 >>
rect 122 25 123 26 
<< m1 >>
rect 123 25 124 26 
<< m1 >>
rect 124 25 125 26 
<< m1 >>
rect 125 25 126 26 
<< m1 >>
rect 126 25 127 26 
<< m1 >>
rect 127 25 128 26 
<< m1 >>
rect 128 25 129 26 
<< m2 >>
rect 128 25 129 26 
<< m1 >>
rect 129 25 130 26 
<< m1 >>
rect 130 25 131 26 
<< m1 >>
rect 131 25 132 26 
<< m1 >>
rect 132 25 133 26 
<< m1 >>
rect 133 25 134 26 
<< m1 >>
rect 134 25 135 26 
<< m1 >>
rect 135 25 136 26 
<< m1 >>
rect 136 25 137 26 
<< m2 >>
rect 136 25 137 26 
<< m1 >>
rect 137 25 138 26 
<< m1 >>
rect 138 25 139 26 
<< m1 >>
rect 139 25 140 26 
<< m2 >>
rect 150 25 151 26 
<< m1 >>
rect 152 25 153 26 
<< m1 >>
rect 154 25 155 26 
<< m1 >>
rect 155 25 156 26 
<< m1 >>
rect 156 25 157 26 
<< m1 >>
rect 157 25 158 26 
<< m1 >>
rect 158 25 159 26 
<< m1 >>
rect 159 25 160 26 
<< m1 >>
rect 160 25 161 26 
<< m1 >>
rect 163 25 164 26 
<< m1 >>
rect 165 25 166 26 
<< m1 >>
rect 167 25 168 26 
<< m1 >>
rect 168 25 169 26 
<< m1 >>
rect 169 25 170 26 
<< m1 >>
rect 170 25 171 26 
<< m1 >>
rect 171 25 172 26 
<< m1 >>
rect 172 25 173 26 
<< m1 >>
rect 173 25 174 26 
<< m1 >>
rect 174 25 175 26 
<< m1 >>
rect 175 25 176 26 
<< m1 >>
rect 176 25 177 26 
<< m1 >>
rect 177 25 178 26 
<< m1 >>
rect 178 25 179 26 
<< m1 >>
rect 190 25 191 26 
<< m1 >>
rect 192 25 193 26 
<< m1 >>
rect 193 25 194 26 
<< m1 >>
rect 194 25 195 26 
<< m1 >>
rect 199 25 200 26 
<< m1 >>
rect 200 25 201 26 
<< m1 >>
rect 201 25 202 26 
<< m2 >>
rect 201 25 202 26 
<< m1 >>
rect 202 25 203 26 
<< m1 >>
rect 203 25 204 26 
<< m1 >>
rect 204 25 205 26 
<< m1 >>
rect 205 25 206 26 
<< m1 >>
rect 206 25 207 26 
<< m1 >>
rect 207 25 208 26 
<< m1 >>
rect 208 25 209 26 
<< m1 >>
rect 209 25 210 26 
<< m1 >>
rect 210 25 211 26 
<< m1 >>
rect 211 25 212 26 
<< m1 >>
rect 212 25 213 26 
<< m1 >>
rect 213 25 214 26 
<< m1 >>
rect 214 25 215 26 
<< m1 >>
rect 215 25 216 26 
<< m1 >>
rect 216 25 217 26 
<< m1 >>
rect 217 25 218 26 
<< m1 >>
rect 218 25 219 26 
<< m1 >>
rect 219 25 220 26 
<< m1 >>
rect 220 25 221 26 
<< m1 >>
rect 221 25 222 26 
<< m1 >>
rect 222 25 223 26 
<< m1 >>
rect 223 25 224 26 
<< m1 >>
rect 224 25 225 26 
<< m1 >>
rect 225 25 226 26 
<< m1 >>
rect 226 25 227 26 
<< m1 >>
rect 227 25 228 26 
<< m1 >>
rect 228 25 229 26 
<< m1 >>
rect 229 25 230 26 
<< m1 >>
rect 230 25 231 26 
<< m1 >>
rect 231 25 232 26 
<< m1 >>
rect 232 25 233 26 
<< m2 >>
rect 233 25 234 26 
<< m1 >>
rect 28 26 29 27 
<< m1 >>
rect 37 26 38 27 
<< m1 >>
rect 40 26 41 27 
<< m1 >>
rect 58 26 59 27 
<< m1 >>
rect 60 26 61 27 
<< m1 >>
rect 67 26 68 27 
<< m1 >>
rect 73 26 74 27 
<< m2 >>
rect 73 26 74 27 
<< m1 >>
rect 85 26 86 27 
<< m1 >>
rect 88 26 89 27 
<< m2 >>
rect 88 26 89 27 
<< m2 >>
rect 118 26 119 27 
<< m2 >>
rect 128 26 129 27 
<< m2 >>
rect 136 26 137 27 
<< m2 >>
rect 146 26 147 27 
<< m2 >>
rect 147 26 148 27 
<< m2 >>
rect 148 26 149 27 
<< m2 >>
rect 149 26 150 27 
<< m2 >>
rect 150 26 151 27 
<< m2 >>
rect 151 26 152 27 
<< m1 >>
rect 152 26 153 27 
<< m2 >>
rect 152 26 153 27 
<< m2c >>
rect 152 26 153 27 
<< m1 >>
rect 152 26 153 27 
<< m2 >>
rect 152 26 153 27 
<< m1 >>
rect 160 26 161 27 
<< m1 >>
rect 163 26 164 27 
<< m2 >>
rect 163 26 164 27 
<< m2c >>
rect 163 26 164 27 
<< m1 >>
rect 163 26 164 27 
<< m2 >>
rect 163 26 164 27 
<< m2 >>
rect 164 26 165 27 
<< m1 >>
rect 165 26 166 27 
<< m2 >>
rect 165 26 166 27 
<< m2 >>
rect 166 26 167 27 
<< m1 >>
rect 167 26 168 27 
<< m2 >>
rect 167 26 168 27 
<< m2c >>
rect 167 26 168 27 
<< m1 >>
rect 167 26 168 27 
<< m2 >>
rect 167 26 168 27 
<< m1 >>
rect 178 26 179 27 
<< m1 >>
rect 190 26 191 27 
<< m1 >>
rect 192 26 193 27 
<< m1 >>
rect 199 26 200 27 
<< m2 >>
rect 201 26 202 27 
<< m2 >>
rect 233 26 234 27 
<< m1 >>
rect 234 26 235 27 
<< m2 >>
rect 234 26 235 27 
<< m2c >>
rect 234 26 235 27 
<< m1 >>
rect 234 26 235 27 
<< m2 >>
rect 234 26 235 27 
<< m1 >>
rect 235 26 236 27 
<< m1 >>
rect 236 26 237 27 
<< m1 >>
rect 237 26 238 27 
<< m1 >>
rect 238 26 239 27 
<< m1 >>
rect 239 26 240 27 
<< m1 >>
rect 240 26 241 27 
<< m1 >>
rect 241 26 242 27 
<< m1 >>
rect 242 26 243 27 
<< m1 >>
rect 243 26 244 27 
<< m1 >>
rect 244 26 245 27 
<< m1 >>
rect 28 27 29 28 
<< m1 >>
rect 37 27 38 28 
<< m1 >>
rect 40 27 41 28 
<< m1 >>
rect 58 27 59 28 
<< m1 >>
rect 60 27 61 28 
<< m1 >>
rect 67 27 68 28 
<< m1 >>
rect 73 27 74 28 
<< m2 >>
rect 73 27 74 28 
<< m1 >>
rect 85 27 86 28 
<< m1 >>
rect 88 27 89 28 
<< m2 >>
rect 88 27 89 28 
<< m2 >>
rect 89 27 90 28 
<< m1 >>
rect 90 27 91 28 
<< m2 >>
rect 90 27 91 28 
<< m2c >>
rect 90 27 91 28 
<< m1 >>
rect 90 27 91 28 
<< m2 >>
rect 90 27 91 28 
<< m1 >>
rect 91 27 92 28 
<< m1 >>
rect 103 27 104 28 
<< m1 >>
rect 104 27 105 28 
<< m1 >>
rect 105 27 106 28 
<< m1 >>
rect 106 27 107 28 
<< m1 >>
rect 107 27 108 28 
<< m1 >>
rect 108 27 109 28 
<< m1 >>
rect 109 27 110 28 
<< m1 >>
rect 110 27 111 28 
<< m1 >>
rect 111 27 112 28 
<< m1 >>
rect 112 27 113 28 
<< m1 >>
rect 113 27 114 28 
<< m1 >>
rect 114 27 115 28 
<< m1 >>
rect 115 27 116 28 
<< m1 >>
rect 116 27 117 28 
<< m1 >>
rect 117 27 118 28 
<< m1 >>
rect 118 27 119 28 
<< m2 >>
rect 118 27 119 28 
<< m2 >>
rect 128 27 129 28 
<< m2 >>
rect 136 27 137 28 
<< m1 >>
rect 139 27 140 28 
<< m1 >>
rect 140 27 141 28 
<< m1 >>
rect 141 27 142 28 
<< m1 >>
rect 142 27 143 28 
<< m1 >>
rect 143 27 144 28 
<< m1 >>
rect 144 27 145 28 
<< m1 >>
rect 145 27 146 28 
<< m1 >>
rect 146 27 147 28 
<< m2 >>
rect 146 27 147 28 
<< m1 >>
rect 147 27 148 28 
<< m1 >>
rect 148 27 149 28 
<< m1 >>
rect 149 27 150 28 
<< m1 >>
rect 150 27 151 28 
<< m2 >>
rect 151 27 152 28 
<< m1 >>
rect 160 27 161 28 
<< m1 >>
rect 165 27 166 28 
<< m1 >>
rect 178 27 179 28 
<< m1 >>
rect 190 27 191 28 
<< m1 >>
rect 192 27 193 28 
<< m1 >>
rect 199 27 200 28 
<< m1 >>
rect 201 27 202 28 
<< m2 >>
rect 201 27 202 28 
<< m2c >>
rect 201 27 202 28 
<< m1 >>
rect 201 27 202 28 
<< m2 >>
rect 201 27 202 28 
<< m1 >>
rect 202 27 203 28 
<< m1 >>
rect 203 27 204 28 
<< m1 >>
rect 244 27 245 28 
<< m1 >>
rect 16 28 17 29 
<< m1 >>
rect 17 28 18 29 
<< m1 >>
rect 18 28 19 29 
<< m1 >>
rect 19 28 20 29 
<< m1 >>
rect 20 28 21 29 
<< m1 >>
rect 21 28 22 29 
<< m1 >>
rect 22 28 23 29 
<< m1 >>
rect 23 28 24 29 
<< m1 >>
rect 24 28 25 29 
<< m1 >>
rect 25 28 26 29 
<< m1 >>
rect 26 28 27 29 
<< m1 >>
rect 28 28 29 29 
<< m1 >>
rect 37 28 38 29 
<< m1 >>
rect 40 28 41 29 
<< m1 >>
rect 44 28 45 29 
<< m1 >>
rect 45 28 46 29 
<< m1 >>
rect 46 28 47 29 
<< m1 >>
rect 47 28 48 29 
<< m1 >>
rect 48 28 49 29 
<< m1 >>
rect 49 28 50 29 
<< m1 >>
rect 58 28 59 29 
<< m1 >>
rect 60 28 61 29 
<< m1 >>
rect 67 28 68 29 
<< m1 >>
rect 73 28 74 29 
<< m2 >>
rect 73 28 74 29 
<< m1 >>
rect 85 28 86 29 
<< m1 >>
rect 88 28 89 29 
<< m1 >>
rect 91 28 92 29 
<< m1 >>
rect 103 28 104 29 
<< m1 >>
rect 118 28 119 29 
<< m2 >>
rect 118 28 119 29 
<< m1 >>
rect 124 28 125 29 
<< m1 >>
rect 125 28 126 29 
<< m1 >>
rect 126 28 127 29 
<< m1 >>
rect 127 28 128 29 
<< m1 >>
rect 128 28 129 29 
<< m2 >>
rect 128 28 129 29 
<< m1 >>
rect 129 28 130 29 
<< m1 >>
rect 130 28 131 29 
<< m1 >>
rect 131 28 132 29 
<< m1 >>
rect 132 28 133 29 
<< m1 >>
rect 133 28 134 29 
<< m1 >>
rect 134 28 135 29 
<< m1 >>
rect 135 28 136 29 
<< m1 >>
rect 136 28 137 29 
<< m2 >>
rect 136 28 137 29 
<< m1 >>
rect 139 28 140 29 
<< m2 >>
rect 146 28 147 29 
<< m1 >>
rect 150 28 151 29 
<< m2 >>
rect 151 28 152 29 
<< m1 >>
rect 160 28 161 29 
<< m1 >>
rect 165 28 166 29 
<< m1 >>
rect 178 28 179 29 
<< m2 >>
rect 189 28 190 29 
<< m1 >>
rect 190 28 191 29 
<< m2 >>
rect 190 28 191 29 
<< m2 >>
rect 191 28 192 29 
<< m1 >>
rect 192 28 193 29 
<< m2 >>
rect 192 28 193 29 
<< m2c >>
rect 192 28 193 29 
<< m1 >>
rect 192 28 193 29 
<< m2 >>
rect 192 28 193 29 
<< m1 >>
rect 199 28 200 29 
<< m1 >>
rect 203 28 204 29 
<< m1 >>
rect 214 28 215 29 
<< m1 >>
rect 215 28 216 29 
<< m1 >>
rect 216 28 217 29 
<< m1 >>
rect 217 28 218 29 
<< m1 >>
rect 218 28 219 29 
<< m1 >>
rect 219 28 220 29 
<< m1 >>
rect 220 28 221 29 
<< m1 >>
rect 221 28 222 29 
<< m1 >>
rect 222 28 223 29 
<< m1 >>
rect 223 28 224 29 
<< m1 >>
rect 224 28 225 29 
<< m1 >>
rect 225 28 226 29 
<< m1 >>
rect 226 28 227 29 
<< m1 >>
rect 244 28 245 29 
<< m1 >>
rect 16 29 17 30 
<< m1 >>
rect 26 29 27 30 
<< m1 >>
rect 28 29 29 30 
<< m1 >>
rect 37 29 38 30 
<< m1 >>
rect 40 29 41 30 
<< m1 >>
rect 44 29 45 30 
<< m1 >>
rect 49 29 50 30 
<< m1 >>
rect 58 29 59 30 
<< m1 >>
rect 60 29 61 30 
<< m1 >>
rect 67 29 68 30 
<< m1 >>
rect 73 29 74 30 
<< m2 >>
rect 73 29 74 30 
<< m1 >>
rect 85 29 86 30 
<< m1 >>
rect 88 29 89 30 
<< m1 >>
rect 91 29 92 30 
<< m1 >>
rect 103 29 104 30 
<< m1 >>
rect 118 29 119 30 
<< m2 >>
rect 118 29 119 30 
<< m1 >>
rect 124 29 125 30 
<< m2 >>
rect 128 29 129 30 
<< m1 >>
rect 136 29 137 30 
<< m2 >>
rect 136 29 137 30 
<< m1 >>
rect 139 29 140 30 
<< m1 >>
rect 146 29 147 30 
<< m2 >>
rect 146 29 147 30 
<< m2c >>
rect 146 29 147 30 
<< m1 >>
rect 146 29 147 30 
<< m2 >>
rect 146 29 147 30 
<< m1 >>
rect 148 29 149 30 
<< m2 >>
rect 148 29 149 30 
<< m2c >>
rect 148 29 149 30 
<< m1 >>
rect 148 29 149 30 
<< m2 >>
rect 148 29 149 30 
<< m2 >>
rect 149 29 150 30 
<< m1 >>
rect 150 29 151 30 
<< m2 >>
rect 150 29 151 30 
<< m2 >>
rect 151 29 152 30 
<< m1 >>
rect 160 29 161 30 
<< m1 >>
rect 165 29 166 30 
<< m1 >>
rect 178 29 179 30 
<< m2 >>
rect 189 29 190 30 
<< m1 >>
rect 190 29 191 30 
<< m1 >>
rect 199 29 200 30 
<< m1 >>
rect 203 29 204 30 
<< m1 >>
rect 214 29 215 30 
<< m1 >>
rect 226 29 227 30 
<< m1 >>
rect 244 29 245 30 
<< pdiffusion >>
rect 12 30 13 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< pdiffusion >>
rect 15 30 16 31 
<< m1 >>
rect 16 30 17 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< m1 >>
rect 26 30 27 31 
<< m1 >>
rect 28 30 29 31 
<< pdiffusion >>
rect 30 30 31 31 
<< pdiffusion >>
rect 31 30 32 31 
<< pdiffusion >>
rect 32 30 33 31 
<< pdiffusion >>
rect 33 30 34 31 
<< pdiffusion >>
rect 34 30 35 31 
<< pdiffusion >>
rect 35 30 36 31 
<< m1 >>
rect 37 30 38 31 
<< m1 >>
rect 40 30 41 31 
<< m1 >>
rect 44 30 45 31 
<< pdiffusion >>
rect 48 30 49 31 
<< m1 >>
rect 49 30 50 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 58 30 59 31 
<< m1 >>
rect 60 30 61 31 
<< m1 >>
rect 67 30 68 31 
<< m1 >>
rect 73 30 74 31 
<< m2 >>
rect 73 30 74 31 
<< pdiffusion >>
rect 84 30 85 31 
<< m1 >>
rect 85 30 86 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< m1 >>
rect 88 30 89 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< m1 >>
rect 91 30 92 31 
<< pdiffusion >>
rect 102 30 103 31 
<< m1 >>
rect 103 30 104 31 
<< pdiffusion >>
rect 103 30 104 31 
<< pdiffusion >>
rect 104 30 105 31 
<< pdiffusion >>
rect 105 30 106 31 
<< pdiffusion >>
rect 106 30 107 31 
<< pdiffusion >>
rect 107 30 108 31 
<< m1 >>
rect 118 30 119 31 
<< m2 >>
rect 118 30 119 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< m1 >>
rect 124 30 125 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< m1 >>
rect 128 30 129 31 
<< m2 >>
rect 128 30 129 31 
<< m2c >>
rect 128 30 129 31 
<< m1 >>
rect 128 30 129 31 
<< m2 >>
rect 128 30 129 31 
<< m1 >>
rect 136 30 137 31 
<< m2 >>
rect 136 30 137 31 
<< pdiffusion >>
rect 138 30 139 31 
<< m1 >>
rect 139 30 140 31 
<< pdiffusion >>
rect 139 30 140 31 
<< pdiffusion >>
rect 140 30 141 31 
<< pdiffusion >>
rect 141 30 142 31 
<< pdiffusion >>
rect 142 30 143 31 
<< pdiffusion >>
rect 143 30 144 31 
<< m1 >>
rect 146 30 147 31 
<< m1 >>
rect 148 30 149 31 
<< m1 >>
rect 150 30 151 31 
<< pdiffusion >>
rect 156 30 157 31 
<< pdiffusion >>
rect 157 30 158 31 
<< pdiffusion >>
rect 158 30 159 31 
<< pdiffusion >>
rect 159 30 160 31 
<< m1 >>
rect 160 30 161 31 
<< pdiffusion >>
rect 160 30 161 31 
<< pdiffusion >>
rect 161 30 162 31 
<< m1 >>
rect 165 30 166 31 
<< pdiffusion >>
rect 174 30 175 31 
<< pdiffusion >>
rect 175 30 176 31 
<< pdiffusion >>
rect 176 30 177 31 
<< pdiffusion >>
rect 177 30 178 31 
<< m1 >>
rect 178 30 179 31 
<< pdiffusion >>
rect 178 30 179 31 
<< pdiffusion >>
rect 179 30 180 31 
<< m2 >>
rect 189 30 190 31 
<< m1 >>
rect 190 30 191 31 
<< pdiffusion >>
rect 192 30 193 31 
<< pdiffusion >>
rect 193 30 194 31 
<< pdiffusion >>
rect 194 30 195 31 
<< pdiffusion >>
rect 195 30 196 31 
<< pdiffusion >>
rect 196 30 197 31 
<< pdiffusion >>
rect 197 30 198 31 
<< m1 >>
rect 199 30 200 31 
<< m1 >>
rect 203 30 204 31 
<< pdiffusion >>
rect 210 30 211 31 
<< pdiffusion >>
rect 211 30 212 31 
<< pdiffusion >>
rect 212 30 213 31 
<< pdiffusion >>
rect 213 30 214 31 
<< m1 >>
rect 214 30 215 31 
<< pdiffusion >>
rect 214 30 215 31 
<< pdiffusion >>
rect 215 30 216 31 
<< m1 >>
rect 226 30 227 31 
<< pdiffusion >>
rect 228 30 229 31 
<< pdiffusion >>
rect 229 30 230 31 
<< pdiffusion >>
rect 230 30 231 31 
<< pdiffusion >>
rect 231 30 232 31 
<< pdiffusion >>
rect 232 30 233 31 
<< pdiffusion >>
rect 233 30 234 31 
<< m1 >>
rect 244 30 245 31 
<< pdiffusion >>
rect 246 30 247 31 
<< pdiffusion >>
rect 247 30 248 31 
<< pdiffusion >>
rect 248 30 249 31 
<< pdiffusion >>
rect 249 30 250 31 
<< pdiffusion >>
rect 250 30 251 31 
<< pdiffusion >>
rect 251 30 252 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< m1 >>
rect 26 31 27 32 
<< m1 >>
rect 28 31 29 32 
<< pdiffusion >>
rect 30 31 31 32 
<< pdiffusion >>
rect 31 31 32 32 
<< pdiffusion >>
rect 32 31 33 32 
<< pdiffusion >>
rect 33 31 34 32 
<< pdiffusion >>
rect 34 31 35 32 
<< pdiffusion >>
rect 35 31 36 32 
<< m1 >>
rect 37 31 38 32 
<< m1 >>
rect 40 31 41 32 
<< m1 >>
rect 44 31 45 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 58 31 59 32 
<< m1 >>
rect 60 31 61 32 
<< m1 >>
rect 67 31 68 32 
<< m1 >>
rect 73 31 74 32 
<< m2 >>
rect 73 31 74 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< m1 >>
rect 91 31 92 32 
<< pdiffusion >>
rect 102 31 103 32 
<< pdiffusion >>
rect 103 31 104 32 
<< pdiffusion >>
rect 104 31 105 32 
<< pdiffusion >>
rect 105 31 106 32 
<< pdiffusion >>
rect 106 31 107 32 
<< pdiffusion >>
rect 107 31 108 32 
<< m1 >>
rect 118 31 119 32 
<< m2 >>
rect 118 31 119 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< m1 >>
rect 128 31 129 32 
<< m1 >>
rect 136 31 137 32 
<< m2 >>
rect 136 31 137 32 
<< pdiffusion >>
rect 138 31 139 32 
<< pdiffusion >>
rect 139 31 140 32 
<< pdiffusion >>
rect 140 31 141 32 
<< pdiffusion >>
rect 141 31 142 32 
<< pdiffusion >>
rect 142 31 143 32 
<< pdiffusion >>
rect 143 31 144 32 
<< m1 >>
rect 146 31 147 32 
<< m1 >>
rect 148 31 149 32 
<< m1 >>
rect 150 31 151 32 
<< pdiffusion >>
rect 156 31 157 32 
<< pdiffusion >>
rect 157 31 158 32 
<< pdiffusion >>
rect 158 31 159 32 
<< pdiffusion >>
rect 159 31 160 32 
<< pdiffusion >>
rect 160 31 161 32 
<< pdiffusion >>
rect 161 31 162 32 
<< m1 >>
rect 165 31 166 32 
<< pdiffusion >>
rect 174 31 175 32 
<< pdiffusion >>
rect 175 31 176 32 
<< pdiffusion >>
rect 176 31 177 32 
<< pdiffusion >>
rect 177 31 178 32 
<< pdiffusion >>
rect 178 31 179 32 
<< pdiffusion >>
rect 179 31 180 32 
<< m2 >>
rect 189 31 190 32 
<< m1 >>
rect 190 31 191 32 
<< pdiffusion >>
rect 192 31 193 32 
<< pdiffusion >>
rect 193 31 194 32 
<< pdiffusion >>
rect 194 31 195 32 
<< pdiffusion >>
rect 195 31 196 32 
<< pdiffusion >>
rect 196 31 197 32 
<< pdiffusion >>
rect 197 31 198 32 
<< m1 >>
rect 199 31 200 32 
<< m1 >>
rect 203 31 204 32 
<< pdiffusion >>
rect 210 31 211 32 
<< pdiffusion >>
rect 211 31 212 32 
<< pdiffusion >>
rect 212 31 213 32 
<< pdiffusion >>
rect 213 31 214 32 
<< pdiffusion >>
rect 214 31 215 32 
<< pdiffusion >>
rect 215 31 216 32 
<< m1 >>
rect 226 31 227 32 
<< pdiffusion >>
rect 228 31 229 32 
<< pdiffusion >>
rect 229 31 230 32 
<< pdiffusion >>
rect 230 31 231 32 
<< pdiffusion >>
rect 231 31 232 32 
<< pdiffusion >>
rect 232 31 233 32 
<< pdiffusion >>
rect 233 31 234 32 
<< m1 >>
rect 244 31 245 32 
<< pdiffusion >>
rect 246 31 247 32 
<< pdiffusion >>
rect 247 31 248 32 
<< pdiffusion >>
rect 248 31 249 32 
<< pdiffusion >>
rect 249 31 250 32 
<< pdiffusion >>
rect 250 31 251 32 
<< pdiffusion >>
rect 251 31 252 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< m1 >>
rect 26 32 27 33 
<< m1 >>
rect 28 32 29 33 
<< pdiffusion >>
rect 30 32 31 33 
<< pdiffusion >>
rect 31 32 32 33 
<< pdiffusion >>
rect 32 32 33 33 
<< pdiffusion >>
rect 33 32 34 33 
<< pdiffusion >>
rect 34 32 35 33 
<< pdiffusion >>
rect 35 32 36 33 
<< m1 >>
rect 37 32 38 33 
<< m1 >>
rect 40 32 41 33 
<< m1 >>
rect 44 32 45 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 58 32 59 33 
<< m1 >>
rect 60 32 61 33 
<< m1 >>
rect 67 32 68 33 
<< m1 >>
rect 73 32 74 33 
<< m2 >>
rect 73 32 74 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< m1 >>
rect 91 32 92 33 
<< pdiffusion >>
rect 102 32 103 33 
<< pdiffusion >>
rect 103 32 104 33 
<< pdiffusion >>
rect 104 32 105 33 
<< pdiffusion >>
rect 105 32 106 33 
<< pdiffusion >>
rect 106 32 107 33 
<< pdiffusion >>
rect 107 32 108 33 
<< m1 >>
rect 118 32 119 33 
<< m2 >>
rect 118 32 119 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< m1 >>
rect 128 32 129 33 
<< m1 >>
rect 136 32 137 33 
<< m2 >>
rect 136 32 137 33 
<< pdiffusion >>
rect 138 32 139 33 
<< pdiffusion >>
rect 139 32 140 33 
<< pdiffusion >>
rect 140 32 141 33 
<< pdiffusion >>
rect 141 32 142 33 
<< pdiffusion >>
rect 142 32 143 33 
<< pdiffusion >>
rect 143 32 144 33 
<< m1 >>
rect 146 32 147 33 
<< m1 >>
rect 148 32 149 33 
<< m1 >>
rect 150 32 151 33 
<< pdiffusion >>
rect 156 32 157 33 
<< pdiffusion >>
rect 157 32 158 33 
<< pdiffusion >>
rect 158 32 159 33 
<< pdiffusion >>
rect 159 32 160 33 
<< pdiffusion >>
rect 160 32 161 33 
<< pdiffusion >>
rect 161 32 162 33 
<< m1 >>
rect 165 32 166 33 
<< pdiffusion >>
rect 174 32 175 33 
<< pdiffusion >>
rect 175 32 176 33 
<< pdiffusion >>
rect 176 32 177 33 
<< pdiffusion >>
rect 177 32 178 33 
<< pdiffusion >>
rect 178 32 179 33 
<< pdiffusion >>
rect 179 32 180 33 
<< m2 >>
rect 189 32 190 33 
<< m1 >>
rect 190 32 191 33 
<< pdiffusion >>
rect 192 32 193 33 
<< pdiffusion >>
rect 193 32 194 33 
<< pdiffusion >>
rect 194 32 195 33 
<< pdiffusion >>
rect 195 32 196 33 
<< pdiffusion >>
rect 196 32 197 33 
<< pdiffusion >>
rect 197 32 198 33 
<< m1 >>
rect 199 32 200 33 
<< m1 >>
rect 203 32 204 33 
<< pdiffusion >>
rect 210 32 211 33 
<< pdiffusion >>
rect 211 32 212 33 
<< pdiffusion >>
rect 212 32 213 33 
<< pdiffusion >>
rect 213 32 214 33 
<< pdiffusion >>
rect 214 32 215 33 
<< pdiffusion >>
rect 215 32 216 33 
<< m1 >>
rect 226 32 227 33 
<< pdiffusion >>
rect 228 32 229 33 
<< pdiffusion >>
rect 229 32 230 33 
<< pdiffusion >>
rect 230 32 231 33 
<< pdiffusion >>
rect 231 32 232 33 
<< pdiffusion >>
rect 232 32 233 33 
<< pdiffusion >>
rect 233 32 234 33 
<< m1 >>
rect 244 32 245 33 
<< pdiffusion >>
rect 246 32 247 33 
<< pdiffusion >>
rect 247 32 248 33 
<< pdiffusion >>
rect 248 32 249 33 
<< pdiffusion >>
rect 249 32 250 33 
<< pdiffusion >>
rect 250 32 251 33 
<< pdiffusion >>
rect 251 32 252 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< m1 >>
rect 26 33 27 34 
<< m1 >>
rect 28 33 29 34 
<< pdiffusion >>
rect 30 33 31 34 
<< pdiffusion >>
rect 31 33 32 34 
<< pdiffusion >>
rect 32 33 33 34 
<< pdiffusion >>
rect 33 33 34 34 
<< pdiffusion >>
rect 34 33 35 34 
<< pdiffusion >>
rect 35 33 36 34 
<< m1 >>
rect 37 33 38 34 
<< m1 >>
rect 40 33 41 34 
<< m1 >>
rect 44 33 45 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 58 33 59 34 
<< m1 >>
rect 60 33 61 34 
<< m1 >>
rect 67 33 68 34 
<< m1 >>
rect 73 33 74 34 
<< m2 >>
rect 73 33 74 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< m1 >>
rect 91 33 92 34 
<< pdiffusion >>
rect 102 33 103 34 
<< pdiffusion >>
rect 103 33 104 34 
<< pdiffusion >>
rect 104 33 105 34 
<< pdiffusion >>
rect 105 33 106 34 
<< pdiffusion >>
rect 106 33 107 34 
<< pdiffusion >>
rect 107 33 108 34 
<< m1 >>
rect 118 33 119 34 
<< m2 >>
rect 118 33 119 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< m1 >>
rect 128 33 129 34 
<< m1 >>
rect 136 33 137 34 
<< m2 >>
rect 136 33 137 34 
<< pdiffusion >>
rect 138 33 139 34 
<< pdiffusion >>
rect 139 33 140 34 
<< pdiffusion >>
rect 140 33 141 34 
<< pdiffusion >>
rect 141 33 142 34 
<< pdiffusion >>
rect 142 33 143 34 
<< pdiffusion >>
rect 143 33 144 34 
<< m1 >>
rect 146 33 147 34 
<< m1 >>
rect 148 33 149 34 
<< m1 >>
rect 150 33 151 34 
<< pdiffusion >>
rect 156 33 157 34 
<< pdiffusion >>
rect 157 33 158 34 
<< pdiffusion >>
rect 158 33 159 34 
<< pdiffusion >>
rect 159 33 160 34 
<< pdiffusion >>
rect 160 33 161 34 
<< pdiffusion >>
rect 161 33 162 34 
<< m1 >>
rect 165 33 166 34 
<< pdiffusion >>
rect 174 33 175 34 
<< pdiffusion >>
rect 175 33 176 34 
<< pdiffusion >>
rect 176 33 177 34 
<< pdiffusion >>
rect 177 33 178 34 
<< pdiffusion >>
rect 178 33 179 34 
<< pdiffusion >>
rect 179 33 180 34 
<< m2 >>
rect 189 33 190 34 
<< m1 >>
rect 190 33 191 34 
<< pdiffusion >>
rect 192 33 193 34 
<< pdiffusion >>
rect 193 33 194 34 
<< pdiffusion >>
rect 194 33 195 34 
<< pdiffusion >>
rect 195 33 196 34 
<< pdiffusion >>
rect 196 33 197 34 
<< pdiffusion >>
rect 197 33 198 34 
<< m1 >>
rect 199 33 200 34 
<< m1 >>
rect 203 33 204 34 
<< pdiffusion >>
rect 210 33 211 34 
<< pdiffusion >>
rect 211 33 212 34 
<< pdiffusion >>
rect 212 33 213 34 
<< pdiffusion >>
rect 213 33 214 34 
<< pdiffusion >>
rect 214 33 215 34 
<< pdiffusion >>
rect 215 33 216 34 
<< m1 >>
rect 226 33 227 34 
<< pdiffusion >>
rect 228 33 229 34 
<< pdiffusion >>
rect 229 33 230 34 
<< pdiffusion >>
rect 230 33 231 34 
<< pdiffusion >>
rect 231 33 232 34 
<< pdiffusion >>
rect 232 33 233 34 
<< pdiffusion >>
rect 233 33 234 34 
<< m1 >>
rect 244 33 245 34 
<< pdiffusion >>
rect 246 33 247 34 
<< pdiffusion >>
rect 247 33 248 34 
<< pdiffusion >>
rect 248 33 249 34 
<< pdiffusion >>
rect 249 33 250 34 
<< pdiffusion >>
rect 250 33 251 34 
<< pdiffusion >>
rect 251 33 252 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< m1 >>
rect 26 34 27 35 
<< m1 >>
rect 28 34 29 35 
<< pdiffusion >>
rect 30 34 31 35 
<< pdiffusion >>
rect 31 34 32 35 
<< pdiffusion >>
rect 32 34 33 35 
<< pdiffusion >>
rect 33 34 34 35 
<< pdiffusion >>
rect 34 34 35 35 
<< pdiffusion >>
rect 35 34 36 35 
<< m1 >>
rect 37 34 38 35 
<< m1 >>
rect 40 34 41 35 
<< m1 >>
rect 44 34 45 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 58 34 59 35 
<< m1 >>
rect 60 34 61 35 
<< m1 >>
rect 67 34 68 35 
<< m1 >>
rect 73 34 74 35 
<< m2 >>
rect 73 34 74 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< m1 >>
rect 91 34 92 35 
<< pdiffusion >>
rect 102 34 103 35 
<< pdiffusion >>
rect 103 34 104 35 
<< pdiffusion >>
rect 104 34 105 35 
<< pdiffusion >>
rect 105 34 106 35 
<< pdiffusion >>
rect 106 34 107 35 
<< pdiffusion >>
rect 107 34 108 35 
<< m1 >>
rect 118 34 119 35 
<< m2 >>
rect 118 34 119 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< m1 >>
rect 128 34 129 35 
<< m1 >>
rect 136 34 137 35 
<< m2 >>
rect 136 34 137 35 
<< pdiffusion >>
rect 138 34 139 35 
<< pdiffusion >>
rect 139 34 140 35 
<< pdiffusion >>
rect 140 34 141 35 
<< pdiffusion >>
rect 141 34 142 35 
<< pdiffusion >>
rect 142 34 143 35 
<< pdiffusion >>
rect 143 34 144 35 
<< m1 >>
rect 146 34 147 35 
<< m1 >>
rect 148 34 149 35 
<< m1 >>
rect 150 34 151 35 
<< pdiffusion >>
rect 156 34 157 35 
<< pdiffusion >>
rect 157 34 158 35 
<< pdiffusion >>
rect 158 34 159 35 
<< pdiffusion >>
rect 159 34 160 35 
<< pdiffusion >>
rect 160 34 161 35 
<< pdiffusion >>
rect 161 34 162 35 
<< m1 >>
rect 165 34 166 35 
<< pdiffusion >>
rect 174 34 175 35 
<< pdiffusion >>
rect 175 34 176 35 
<< pdiffusion >>
rect 176 34 177 35 
<< pdiffusion >>
rect 177 34 178 35 
<< pdiffusion >>
rect 178 34 179 35 
<< pdiffusion >>
rect 179 34 180 35 
<< m2 >>
rect 189 34 190 35 
<< m1 >>
rect 190 34 191 35 
<< pdiffusion >>
rect 192 34 193 35 
<< pdiffusion >>
rect 193 34 194 35 
<< pdiffusion >>
rect 194 34 195 35 
<< pdiffusion >>
rect 195 34 196 35 
<< pdiffusion >>
rect 196 34 197 35 
<< pdiffusion >>
rect 197 34 198 35 
<< m1 >>
rect 199 34 200 35 
<< m1 >>
rect 203 34 204 35 
<< pdiffusion >>
rect 210 34 211 35 
<< pdiffusion >>
rect 211 34 212 35 
<< pdiffusion >>
rect 212 34 213 35 
<< pdiffusion >>
rect 213 34 214 35 
<< pdiffusion >>
rect 214 34 215 35 
<< pdiffusion >>
rect 215 34 216 35 
<< m1 >>
rect 226 34 227 35 
<< pdiffusion >>
rect 228 34 229 35 
<< pdiffusion >>
rect 229 34 230 35 
<< pdiffusion >>
rect 230 34 231 35 
<< pdiffusion >>
rect 231 34 232 35 
<< pdiffusion >>
rect 232 34 233 35 
<< pdiffusion >>
rect 233 34 234 35 
<< m1 >>
rect 244 34 245 35 
<< pdiffusion >>
rect 246 34 247 35 
<< pdiffusion >>
rect 247 34 248 35 
<< pdiffusion >>
rect 248 34 249 35 
<< pdiffusion >>
rect 249 34 250 35 
<< pdiffusion >>
rect 250 34 251 35 
<< pdiffusion >>
rect 251 34 252 35 
<< pdiffusion >>
rect 12 35 13 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< m1 >>
rect 26 35 27 36 
<< m1 >>
rect 28 35 29 36 
<< pdiffusion >>
rect 30 35 31 36 
<< m1 >>
rect 31 35 32 36 
<< pdiffusion >>
rect 31 35 32 36 
<< pdiffusion >>
rect 32 35 33 36 
<< pdiffusion >>
rect 33 35 34 36 
<< pdiffusion >>
rect 34 35 35 36 
<< pdiffusion >>
rect 35 35 36 36 
<< m1 >>
rect 37 35 38 36 
<< m1 >>
rect 40 35 41 36 
<< m1 >>
rect 44 35 45 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 58 35 59 36 
<< m1 >>
rect 60 35 61 36 
<< m1 >>
rect 67 35 68 36 
<< m1 >>
rect 73 35 74 36 
<< m2 >>
rect 73 35 74 36 
<< pdiffusion >>
rect 84 35 85 36 
<< m1 >>
rect 85 35 86 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< m1 >>
rect 91 35 92 36 
<< pdiffusion >>
rect 102 35 103 36 
<< m1 >>
rect 103 35 104 36 
<< pdiffusion >>
rect 103 35 104 36 
<< pdiffusion >>
rect 104 35 105 36 
<< pdiffusion >>
rect 105 35 106 36 
<< pdiffusion >>
rect 106 35 107 36 
<< pdiffusion >>
rect 107 35 108 36 
<< m1 >>
rect 118 35 119 36 
<< m2 >>
rect 118 35 119 36 
<< pdiffusion >>
rect 120 35 121 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< m1 >>
rect 124 35 125 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< m1 >>
rect 128 35 129 36 
<< m1 >>
rect 136 35 137 36 
<< m2 >>
rect 136 35 137 36 
<< pdiffusion >>
rect 138 35 139 36 
<< pdiffusion >>
rect 139 35 140 36 
<< pdiffusion >>
rect 140 35 141 36 
<< pdiffusion >>
rect 141 35 142 36 
<< m1 >>
rect 142 35 143 36 
<< pdiffusion >>
rect 142 35 143 36 
<< pdiffusion >>
rect 143 35 144 36 
<< m1 >>
rect 146 35 147 36 
<< m1 >>
rect 148 35 149 36 
<< m1 >>
rect 150 35 151 36 
<< pdiffusion >>
rect 156 35 157 36 
<< pdiffusion >>
rect 157 35 158 36 
<< pdiffusion >>
rect 158 35 159 36 
<< pdiffusion >>
rect 159 35 160 36 
<< m1 >>
rect 160 35 161 36 
<< pdiffusion >>
rect 160 35 161 36 
<< pdiffusion >>
rect 161 35 162 36 
<< m1 >>
rect 165 35 166 36 
<< pdiffusion >>
rect 174 35 175 36 
<< pdiffusion >>
rect 175 35 176 36 
<< pdiffusion >>
rect 176 35 177 36 
<< pdiffusion >>
rect 177 35 178 36 
<< m1 >>
rect 178 35 179 36 
<< pdiffusion >>
rect 178 35 179 36 
<< pdiffusion >>
rect 179 35 180 36 
<< m2 >>
rect 189 35 190 36 
<< m1 >>
rect 190 35 191 36 
<< pdiffusion >>
rect 192 35 193 36 
<< pdiffusion >>
rect 193 35 194 36 
<< pdiffusion >>
rect 194 35 195 36 
<< pdiffusion >>
rect 195 35 196 36 
<< m1 >>
rect 196 35 197 36 
<< pdiffusion >>
rect 196 35 197 36 
<< pdiffusion >>
rect 197 35 198 36 
<< m1 >>
rect 199 35 200 36 
<< m1 >>
rect 203 35 204 36 
<< pdiffusion >>
rect 210 35 211 36 
<< pdiffusion >>
rect 211 35 212 36 
<< pdiffusion >>
rect 212 35 213 36 
<< pdiffusion >>
rect 213 35 214 36 
<< pdiffusion >>
rect 214 35 215 36 
<< pdiffusion >>
rect 215 35 216 36 
<< m1 >>
rect 226 35 227 36 
<< pdiffusion >>
rect 228 35 229 36 
<< pdiffusion >>
rect 229 35 230 36 
<< pdiffusion >>
rect 230 35 231 36 
<< pdiffusion >>
rect 231 35 232 36 
<< m1 >>
rect 232 35 233 36 
<< pdiffusion >>
rect 232 35 233 36 
<< pdiffusion >>
rect 233 35 234 36 
<< m1 >>
rect 244 35 245 36 
<< pdiffusion >>
rect 246 35 247 36 
<< pdiffusion >>
rect 247 35 248 36 
<< pdiffusion >>
rect 248 35 249 36 
<< pdiffusion >>
rect 249 35 250 36 
<< pdiffusion >>
rect 250 35 251 36 
<< pdiffusion >>
rect 251 35 252 36 
<< m1 >>
rect 26 36 27 37 
<< m1 >>
rect 28 36 29 37 
<< m1 >>
rect 31 36 32 37 
<< m1 >>
rect 37 36 38 37 
<< m2 >>
rect 37 36 38 37 
<< m2c >>
rect 37 36 38 37 
<< m1 >>
rect 37 36 38 37 
<< m2 >>
rect 37 36 38 37 
<< m1 >>
rect 40 36 41 37 
<< m2 >>
rect 40 36 41 37 
<< m2c >>
rect 40 36 41 37 
<< m1 >>
rect 40 36 41 37 
<< m2 >>
rect 40 36 41 37 
<< m1 >>
rect 44 36 45 37 
<< m1 >>
rect 58 36 59 37 
<< m1 >>
rect 60 36 61 37 
<< m1 >>
rect 67 36 68 37 
<< m1 >>
rect 73 36 74 37 
<< m2 >>
rect 73 36 74 37 
<< m1 >>
rect 85 36 86 37 
<< m1 >>
rect 91 36 92 37 
<< m1 >>
rect 103 36 104 37 
<< m1 >>
rect 118 36 119 37 
<< m2 >>
rect 118 36 119 37 
<< m1 >>
rect 124 36 125 37 
<< m1 >>
rect 128 36 129 37 
<< m1 >>
rect 136 36 137 37 
<< m2 >>
rect 136 36 137 37 
<< m1 >>
rect 142 36 143 37 
<< m1 >>
rect 146 36 147 37 
<< m1 >>
rect 148 36 149 37 
<< m1 >>
rect 150 36 151 37 
<< m1 >>
rect 160 36 161 37 
<< m1 >>
rect 165 36 166 37 
<< m1 >>
rect 178 36 179 37 
<< m2 >>
rect 189 36 190 37 
<< m1 >>
rect 190 36 191 37 
<< m1 >>
rect 196 36 197 37 
<< m1 >>
rect 199 36 200 37 
<< m1 >>
rect 203 36 204 37 
<< m1 >>
rect 226 36 227 37 
<< m1 >>
rect 232 36 233 37 
<< m1 >>
rect 244 36 245 37 
<< m1 >>
rect 26 37 27 38 
<< m1 >>
rect 28 37 29 38 
<< m1 >>
rect 31 37 32 38 
<< m2 >>
rect 37 37 38 38 
<< m2 >>
rect 40 37 41 38 
<< m1 >>
rect 44 37 45 38 
<< m1 >>
rect 58 37 59 38 
<< m1 >>
rect 60 37 61 38 
<< m1 >>
rect 67 37 68 38 
<< m1 >>
rect 73 37 74 38 
<< m2 >>
rect 73 37 74 38 
<< m1 >>
rect 74 37 75 38 
<< m1 >>
rect 75 37 76 38 
<< m1 >>
rect 76 37 77 38 
<< m1 >>
rect 77 37 78 38 
<< m1 >>
rect 78 37 79 38 
<< m1 >>
rect 79 37 80 38 
<< m1 >>
rect 80 37 81 38 
<< m1 >>
rect 81 37 82 38 
<< m1 >>
rect 82 37 83 38 
<< m1 >>
rect 83 37 84 38 
<< m1 >>
rect 84 37 85 38 
<< m1 >>
rect 85 37 86 38 
<< m1 >>
rect 91 37 92 38 
<< m1 >>
rect 103 37 104 38 
<< m1 >>
rect 118 37 119 38 
<< m2 >>
rect 118 37 119 38 
<< m1 >>
rect 124 37 125 38 
<< m1 >>
rect 128 37 129 38 
<< m1 >>
rect 136 37 137 38 
<< m2 >>
rect 136 37 137 38 
<< m1 >>
rect 142 37 143 38 
<< m1 >>
rect 146 37 147 38 
<< m1 >>
rect 148 37 149 38 
<< m1 >>
rect 150 37 151 38 
<< m1 >>
rect 160 37 161 38 
<< m1 >>
rect 161 37 162 38 
<< m1 >>
rect 162 37 163 38 
<< m1 >>
rect 163 37 164 38 
<< m1 >>
rect 165 37 166 38 
<< m1 >>
rect 178 37 179 38 
<< m2 >>
rect 189 37 190 38 
<< m1 >>
rect 190 37 191 38 
<< m1 >>
rect 196 37 197 38 
<< m1 >>
rect 199 37 200 38 
<< m1 >>
rect 203 37 204 38 
<< m1 >>
rect 226 37 227 38 
<< m1 >>
rect 232 37 233 38 
<< m1 >>
rect 244 37 245 38 
<< m1 >>
rect 26 38 27 39 
<< m1 >>
rect 28 38 29 39 
<< m1 >>
rect 31 38 32 39 
<< m1 >>
rect 32 38 33 39 
<< m1 >>
rect 33 38 34 39 
<< m1 >>
rect 34 38 35 39 
<< m1 >>
rect 35 38 36 39 
<< m1 >>
rect 36 38 37 39 
<< m1 >>
rect 37 38 38 39 
<< m2 >>
rect 37 38 38 39 
<< m1 >>
rect 38 38 39 39 
<< m1 >>
rect 39 38 40 39 
<< m1 >>
rect 40 38 41 39 
<< m2 >>
rect 40 38 41 39 
<< m1 >>
rect 41 38 42 39 
<< m1 >>
rect 42 38 43 39 
<< m2 >>
rect 42 38 43 39 
<< m2c >>
rect 42 38 43 39 
<< m1 >>
rect 42 38 43 39 
<< m2 >>
rect 42 38 43 39 
<< m2 >>
rect 43 38 44 39 
<< m1 >>
rect 44 38 45 39 
<< m1 >>
rect 58 38 59 39 
<< m1 >>
rect 60 38 61 39 
<< m1 >>
rect 67 38 68 39 
<< m2 >>
rect 73 38 74 39 
<< m1 >>
rect 91 38 92 39 
<< m1 >>
rect 103 38 104 39 
<< m1 >>
rect 118 38 119 39 
<< m2 >>
rect 118 38 119 39 
<< m1 >>
rect 124 38 125 39 
<< m1 >>
rect 128 38 129 39 
<< m1 >>
rect 136 38 137 39 
<< m2 >>
rect 136 38 137 39 
<< m1 >>
rect 137 38 138 39 
<< m1 >>
rect 138 38 139 39 
<< m2 >>
rect 138 38 139 39 
<< m2c >>
rect 138 38 139 39 
<< m1 >>
rect 138 38 139 39 
<< m2 >>
rect 138 38 139 39 
<< m1 >>
rect 142 38 143 39 
<< m1 >>
rect 146 38 147 39 
<< m1 >>
rect 148 38 149 39 
<< m1 >>
rect 150 38 151 39 
<< m1 >>
rect 163 38 164 39 
<< m1 >>
rect 165 38 166 39 
<< m1 >>
rect 178 38 179 39 
<< m1 >>
rect 186 38 187 39 
<< m1 >>
rect 187 38 188 39 
<< m1 >>
rect 188 38 189 39 
<< m2 >>
rect 188 38 189 39 
<< m2c >>
rect 188 38 189 39 
<< m1 >>
rect 188 38 189 39 
<< m2 >>
rect 188 38 189 39 
<< m2 >>
rect 189 38 190 39 
<< m1 >>
rect 190 38 191 39 
<< m1 >>
rect 196 38 197 39 
<< m1 >>
rect 199 38 200 39 
<< m1 >>
rect 203 38 204 39 
<< m2 >>
rect 203 38 204 39 
<< m2c >>
rect 203 38 204 39 
<< m1 >>
rect 203 38 204 39 
<< m2 >>
rect 203 38 204 39 
<< m1 >>
rect 226 38 227 39 
<< m1 >>
rect 227 38 228 39 
<< m1 >>
rect 228 38 229 39 
<< m2 >>
rect 228 38 229 39 
<< m2c >>
rect 228 38 229 39 
<< m1 >>
rect 228 38 229 39 
<< m2 >>
rect 228 38 229 39 
<< m1 >>
rect 232 38 233 39 
<< m1 >>
rect 244 38 245 39 
<< m1 >>
rect 26 39 27 40 
<< m1 >>
rect 28 39 29 40 
<< m2 >>
rect 37 39 38 40 
<< m2 >>
rect 40 39 41 40 
<< m2 >>
rect 43 39 44 40 
<< m1 >>
rect 44 39 45 40 
<< m1 >>
rect 58 39 59 40 
<< m1 >>
rect 60 39 61 40 
<< m1 >>
rect 67 39 68 40 
<< m1 >>
rect 73 39 74 40 
<< m2 >>
rect 73 39 74 40 
<< m2c >>
rect 73 39 74 40 
<< m1 >>
rect 73 39 74 40 
<< m2 >>
rect 73 39 74 40 
<< m1 >>
rect 91 39 92 40 
<< m2 >>
rect 91 39 92 40 
<< m2c >>
rect 91 39 92 40 
<< m1 >>
rect 91 39 92 40 
<< m2 >>
rect 91 39 92 40 
<< m1 >>
rect 103 39 104 40 
<< m1 >>
rect 118 39 119 40 
<< m2 >>
rect 118 39 119 40 
<< m1 >>
rect 124 39 125 40 
<< m1 >>
rect 128 39 129 40 
<< m2 >>
rect 136 39 137 40 
<< m2 >>
rect 138 39 139 40 
<< m1 >>
rect 142 39 143 40 
<< m1 >>
rect 146 39 147 40 
<< m2 >>
rect 146 39 147 40 
<< m2c >>
rect 146 39 147 40 
<< m1 >>
rect 146 39 147 40 
<< m2 >>
rect 146 39 147 40 
<< m1 >>
rect 148 39 149 40 
<< m2 >>
rect 148 39 149 40 
<< m2c >>
rect 148 39 149 40 
<< m1 >>
rect 148 39 149 40 
<< m2 >>
rect 148 39 149 40 
<< m1 >>
rect 150 39 151 40 
<< m2 >>
rect 150 39 151 40 
<< m2c >>
rect 150 39 151 40 
<< m1 >>
rect 150 39 151 40 
<< m2 >>
rect 150 39 151 40 
<< m1 >>
rect 163 39 164 40 
<< m1 >>
rect 165 39 166 40 
<< m1 >>
rect 178 39 179 40 
<< m1 >>
rect 186 39 187 40 
<< m1 >>
rect 190 39 191 40 
<< m1 >>
rect 196 39 197 40 
<< m1 >>
rect 199 39 200 40 
<< m2 >>
rect 203 39 204 40 
<< m2 >>
rect 228 39 229 40 
<< m1 >>
rect 232 39 233 40 
<< m1 >>
rect 244 39 245 40 
<< m1 >>
rect 26 40 27 41 
<< m1 >>
rect 28 40 29 41 
<< m1 >>
rect 37 40 38 41 
<< m2 >>
rect 37 40 38 41 
<< m2c >>
rect 37 40 38 41 
<< m1 >>
rect 37 40 38 41 
<< m2 >>
rect 37 40 38 41 
<< m1 >>
rect 40 40 41 41 
<< m2 >>
rect 40 40 41 41 
<< m2c >>
rect 40 40 41 41 
<< m1 >>
rect 40 40 41 41 
<< m2 >>
rect 40 40 41 41 
<< m2 >>
rect 43 40 44 41 
<< m1 >>
rect 44 40 45 41 
<< m1 >>
rect 58 40 59 41 
<< m1 >>
rect 60 40 61 41 
<< m1 >>
rect 67 40 68 41 
<< m1 >>
rect 73 40 74 41 
<< m2 >>
rect 91 40 92 41 
<< m2 >>
rect 92 40 93 41 
<< m2 >>
rect 93 40 94 41 
<< m2 >>
rect 94 40 95 41 
<< m2 >>
rect 95 40 96 41 
<< m2 >>
rect 96 40 97 41 
<< m2 >>
rect 97 40 98 41 
<< m2 >>
rect 98 40 99 41 
<< m2 >>
rect 99 40 100 41 
<< m2 >>
rect 100 40 101 41 
<< m2 >>
rect 101 40 102 41 
<< m2 >>
rect 102 40 103 41 
<< m1 >>
rect 103 40 104 41 
<< m2 >>
rect 103 40 104 41 
<< m2 >>
rect 104 40 105 41 
<< m1 >>
rect 105 40 106 41 
<< m2 >>
rect 105 40 106 41 
<< m2c >>
rect 105 40 106 41 
<< m1 >>
rect 105 40 106 41 
<< m2 >>
rect 105 40 106 41 
<< m1 >>
rect 106 40 107 41 
<< m1 >>
rect 107 40 108 41 
<< m1 >>
rect 108 40 109 41 
<< m1 >>
rect 118 40 119 41 
<< m2 >>
rect 118 40 119 41 
<< m1 >>
rect 124 40 125 41 
<< m1 >>
rect 128 40 129 41 
<< m1 >>
rect 136 40 137 41 
<< m2 >>
rect 136 40 137 41 
<< m1 >>
rect 137 40 138 41 
<< m1 >>
rect 138 40 139 41 
<< m2 >>
rect 138 40 139 41 
<< m1 >>
rect 139 40 140 41 
<< m1 >>
rect 140 40 141 41 
<< m1 >>
rect 141 40 142 41 
<< m1 >>
rect 142 40 143 41 
<< m2 >>
rect 146 40 147 41 
<< m2 >>
rect 148 40 149 41 
<< m2 >>
rect 150 40 151 41 
<< m1 >>
rect 163 40 164 41 
<< m1 >>
rect 165 40 166 41 
<< m1 >>
rect 178 40 179 41 
<< m1 >>
rect 186 40 187 41 
<< m1 >>
rect 190 40 191 41 
<< m2 >>
rect 190 40 191 41 
<< m1 >>
rect 191 40 192 41 
<< m2 >>
rect 191 40 192 41 
<< m1 >>
rect 192 40 193 41 
<< m2 >>
rect 192 40 193 41 
<< m1 >>
rect 193 40 194 41 
<< m2 >>
rect 193 40 194 41 
<< m1 >>
rect 194 40 195 41 
<< m2 >>
rect 194 40 195 41 
<< m1 >>
rect 195 40 196 41 
<< m2 >>
rect 195 40 196 41 
<< m1 >>
rect 196 40 197 41 
<< m2 >>
rect 196 40 197 41 
<< m2 >>
rect 197 40 198 41 
<< m2 >>
rect 198 40 199 41 
<< m1 >>
rect 199 40 200 41 
<< m2 >>
rect 199 40 200 41 
<< m2 >>
rect 200 40 201 41 
<< m1 >>
rect 201 40 202 41 
<< m2 >>
rect 201 40 202 41 
<< m2c >>
rect 201 40 202 41 
<< m1 >>
rect 201 40 202 41 
<< m2 >>
rect 201 40 202 41 
<< m1 >>
rect 202 40 203 41 
<< m1 >>
rect 203 40 204 41 
<< m2 >>
rect 203 40 204 41 
<< m1 >>
rect 204 40 205 41 
<< m1 >>
rect 205 40 206 41 
<< m1 >>
rect 206 40 207 41 
<< m1 >>
rect 207 40 208 41 
<< m1 >>
rect 208 40 209 41 
<< m1 >>
rect 209 40 210 41 
<< m1 >>
rect 210 40 211 41 
<< m1 >>
rect 211 40 212 41 
<< m1 >>
rect 212 40 213 41 
<< m1 >>
rect 213 40 214 41 
<< m1 >>
rect 214 40 215 41 
<< m1 >>
rect 215 40 216 41 
<< m1 >>
rect 216 40 217 41 
<< m1 >>
rect 217 40 218 41 
<< m1 >>
rect 218 40 219 41 
<< m1 >>
rect 219 40 220 41 
<< m1 >>
rect 220 40 221 41 
<< m1 >>
rect 221 40 222 41 
<< m1 >>
rect 222 40 223 41 
<< m1 >>
rect 223 40 224 41 
<< m1 >>
rect 224 40 225 41 
<< m1 >>
rect 225 40 226 41 
<< m1 >>
rect 226 40 227 41 
<< m1 >>
rect 227 40 228 41 
<< m1 >>
rect 228 40 229 41 
<< m2 >>
rect 228 40 229 41 
<< m1 >>
rect 229 40 230 41 
<< m1 >>
rect 230 40 231 41 
<< m1 >>
rect 231 40 232 41 
<< m1 >>
rect 232 40 233 41 
<< m1 >>
rect 244 40 245 41 
<< m1 >>
rect 26 41 27 42 
<< m1 >>
rect 28 41 29 42 
<< m1 >>
rect 37 41 38 42 
<< m1 >>
rect 40 41 41 42 
<< m2 >>
rect 43 41 44 42 
<< m1 >>
rect 44 41 45 42 
<< m1 >>
rect 58 41 59 42 
<< m1 >>
rect 60 41 61 42 
<< m1 >>
rect 67 41 68 42 
<< m1 >>
rect 68 41 69 42 
<< m1 >>
rect 69 41 70 42 
<< m1 >>
rect 70 41 71 42 
<< m1 >>
rect 71 41 72 42 
<< m2 >>
rect 71 41 72 42 
<< m2c >>
rect 71 41 72 42 
<< m1 >>
rect 71 41 72 42 
<< m2 >>
rect 71 41 72 42 
<< m2 >>
rect 72 41 73 42 
<< m1 >>
rect 73 41 74 42 
<< m2 >>
rect 73 41 74 42 
<< m2 >>
rect 74 41 75 42 
<< m1 >>
rect 75 41 76 42 
<< m2 >>
rect 75 41 76 42 
<< m1 >>
rect 76 41 77 42 
<< m2 >>
rect 76 41 77 42 
<< m1 >>
rect 77 41 78 42 
<< m2 >>
rect 77 41 78 42 
<< m1 >>
rect 78 41 79 42 
<< m2 >>
rect 78 41 79 42 
<< m1 >>
rect 79 41 80 42 
<< m2 >>
rect 79 41 80 42 
<< m1 >>
rect 80 41 81 42 
<< m2 >>
rect 80 41 81 42 
<< m1 >>
rect 81 41 82 42 
<< m2 >>
rect 81 41 82 42 
<< m1 >>
rect 82 41 83 42 
<< m2 >>
rect 82 41 83 42 
<< m1 >>
rect 83 41 84 42 
<< m2 >>
rect 83 41 84 42 
<< m1 >>
rect 84 41 85 42 
<< m2 >>
rect 84 41 85 42 
<< m1 >>
rect 85 41 86 42 
<< m2 >>
rect 85 41 86 42 
<< m1 >>
rect 86 41 87 42 
<< m2 >>
rect 86 41 87 42 
<< m1 >>
rect 87 41 88 42 
<< m2 >>
rect 87 41 88 42 
<< m1 >>
rect 88 41 89 42 
<< m1 >>
rect 89 41 90 42 
<< m1 >>
rect 90 41 91 42 
<< m1 >>
rect 91 41 92 42 
<< m1 >>
rect 92 41 93 42 
<< m1 >>
rect 93 41 94 42 
<< m1 >>
rect 94 41 95 42 
<< m1 >>
rect 95 41 96 42 
<< m1 >>
rect 96 41 97 42 
<< m1 >>
rect 97 41 98 42 
<< m1 >>
rect 98 41 99 42 
<< m1 >>
rect 99 41 100 42 
<< m1 >>
rect 100 41 101 42 
<< m1 >>
rect 101 41 102 42 
<< m1 >>
rect 102 41 103 42 
<< m1 >>
rect 103 41 104 42 
<< m1 >>
rect 108 41 109 42 
<< m2 >>
rect 108 41 109 42 
<< m2c >>
rect 108 41 109 42 
<< m1 >>
rect 108 41 109 42 
<< m2 >>
rect 108 41 109 42 
<< m1 >>
rect 118 41 119 42 
<< m2 >>
rect 118 41 119 42 
<< m1 >>
rect 119 41 120 42 
<< m1 >>
rect 120 41 121 42 
<< m1 >>
rect 121 41 122 42 
<< m1 >>
rect 122 41 123 42 
<< m2 >>
rect 122 41 123 42 
<< m2c >>
rect 122 41 123 42 
<< m1 >>
rect 122 41 123 42 
<< m2 >>
rect 122 41 123 42 
<< m2 >>
rect 123 41 124 42 
<< m1 >>
rect 124 41 125 42 
<< m2 >>
rect 124 41 125 42 
<< m2 >>
rect 125 41 126 42 
<< m1 >>
rect 128 41 129 42 
<< m1 >>
rect 136 41 137 42 
<< m2 >>
rect 136 41 137 42 
<< m2 >>
rect 138 41 139 42 
<< m2 >>
rect 139 41 140 42 
<< m2 >>
rect 140 41 141 42 
<< m2 >>
rect 141 41 142 42 
<< m2 >>
rect 142 41 143 42 
<< m2 >>
rect 143 41 144 42 
<< m1 >>
rect 144 41 145 42 
<< m2 >>
rect 144 41 145 42 
<< m2c >>
rect 144 41 145 42 
<< m1 >>
rect 144 41 145 42 
<< m2 >>
rect 144 41 145 42 
<< m1 >>
rect 145 41 146 42 
<< m1 >>
rect 146 41 147 42 
<< m2 >>
rect 146 41 147 42 
<< m1 >>
rect 147 41 148 42 
<< m1 >>
rect 148 41 149 42 
<< m2 >>
rect 148 41 149 42 
<< m1 >>
rect 149 41 150 42 
<< m1 >>
rect 150 41 151 42 
<< m2 >>
rect 150 41 151 42 
<< m1 >>
rect 151 41 152 42 
<< m1 >>
rect 152 41 153 42 
<< m1 >>
rect 153 41 154 42 
<< m1 >>
rect 154 41 155 42 
<< m1 >>
rect 163 41 164 42 
<< m1 >>
rect 165 41 166 42 
<< m1 >>
rect 178 41 179 42 
<< m1 >>
rect 186 41 187 42 
<< m2 >>
rect 190 41 191 42 
<< m1 >>
rect 199 41 200 42 
<< m2 >>
rect 203 41 204 42 
<< m2 >>
rect 228 41 229 42 
<< m2 >>
rect 229 41 230 42 
<< m2 >>
rect 230 41 231 42 
<< m2 >>
rect 231 41 232 42 
<< m2 >>
rect 232 41 233 42 
<< m1 >>
rect 244 41 245 42 
<< m1 >>
rect 26 42 27 43 
<< m1 >>
rect 28 42 29 43 
<< m1 >>
rect 37 42 38 43 
<< m1 >>
rect 40 42 41 43 
<< m2 >>
rect 43 42 44 43 
<< m1 >>
rect 44 42 45 43 
<< m1 >>
rect 58 42 59 43 
<< m1 >>
rect 60 42 61 43 
<< m1 >>
rect 73 42 74 43 
<< m1 >>
rect 75 42 76 43 
<< m2 >>
rect 87 42 88 43 
<< m2 >>
rect 108 42 109 43 
<< m2 >>
rect 109 42 110 43 
<< m2 >>
rect 118 42 119 43 
<< m1 >>
rect 124 42 125 43 
<< m2 >>
rect 125 42 126 43 
<< m1 >>
rect 128 42 129 43 
<< m2 >>
rect 128 42 129 43 
<< m2c >>
rect 128 42 129 43 
<< m1 >>
rect 128 42 129 43 
<< m2 >>
rect 128 42 129 43 
<< m1 >>
rect 136 42 137 43 
<< m2 >>
rect 136 42 137 43 
<< m2 >>
rect 146 42 147 43 
<< m2 >>
rect 148 42 149 43 
<< m2 >>
rect 150 42 151 43 
<< m1 >>
rect 154 42 155 43 
<< m1 >>
rect 163 42 164 43 
<< m1 >>
rect 165 42 166 43 
<< m1 >>
rect 178 42 179 43 
<< m1 >>
rect 186 42 187 43 
<< m2 >>
rect 190 42 191 43 
<< m1 >>
rect 199 42 200 43 
<< m2 >>
rect 203 42 204 43 
<< m1 >>
rect 232 42 233 43 
<< m2 >>
rect 232 42 233 43 
<< m1 >>
rect 244 42 245 43 
<< m1 >>
rect 26 43 27 44 
<< m1 >>
rect 28 43 29 44 
<< m1 >>
rect 37 43 38 44 
<< m1 >>
rect 40 43 41 44 
<< m2 >>
rect 43 43 44 44 
<< m1 >>
rect 44 43 45 44 
<< m1 >>
rect 58 43 59 44 
<< m1 >>
rect 60 43 61 44 
<< m1 >>
rect 73 43 74 44 
<< m1 >>
rect 75 43 76 44 
<< m2 >>
rect 76 43 77 44 
<< m1 >>
rect 77 43 78 44 
<< m2 >>
rect 77 43 78 44 
<< m2c >>
rect 77 43 78 44 
<< m1 >>
rect 77 43 78 44 
<< m2 >>
rect 77 43 78 44 
<< m1 >>
rect 78 43 79 44 
<< m1 >>
rect 79 43 80 44 
<< m1 >>
rect 80 43 81 44 
<< m1 >>
rect 81 43 82 44 
<< m1 >>
rect 82 43 83 44 
<< m1 >>
rect 83 43 84 44 
<< m1 >>
rect 84 43 85 44 
<< m1 >>
rect 85 43 86 44 
<< m1 >>
rect 86 43 87 44 
<< m1 >>
rect 87 43 88 44 
<< m2 >>
rect 87 43 88 44 
<< m1 >>
rect 88 43 89 44 
<< m1 >>
rect 89 43 90 44 
<< m2 >>
rect 89 43 90 44 
<< m2c >>
rect 89 43 90 44 
<< m1 >>
rect 89 43 90 44 
<< m2 >>
rect 89 43 90 44 
<< m2 >>
rect 90 43 91 44 
<< m1 >>
rect 91 43 92 44 
<< m2 >>
rect 91 43 92 44 
<< m1 >>
rect 92 43 93 44 
<< m2 >>
rect 92 43 93 44 
<< m1 >>
rect 93 43 94 44 
<< m2 >>
rect 93 43 94 44 
<< m1 >>
rect 94 43 95 44 
<< m2 >>
rect 94 43 95 44 
<< m1 >>
rect 95 43 96 44 
<< m2 >>
rect 95 43 96 44 
<< m1 >>
rect 96 43 97 44 
<< m2 >>
rect 96 43 97 44 
<< m1 >>
rect 97 43 98 44 
<< m2 >>
rect 97 43 98 44 
<< m1 >>
rect 98 43 99 44 
<< m2 >>
rect 98 43 99 44 
<< m1 >>
rect 99 43 100 44 
<< m2 >>
rect 99 43 100 44 
<< m1 >>
rect 100 43 101 44 
<< m2 >>
rect 100 43 101 44 
<< m1 >>
rect 101 43 102 44 
<< m2 >>
rect 101 43 102 44 
<< m1 >>
rect 102 43 103 44 
<< m2 >>
rect 102 43 103 44 
<< m1 >>
rect 103 43 104 44 
<< m2 >>
rect 103 43 104 44 
<< m1 >>
rect 104 43 105 44 
<< m2 >>
rect 104 43 105 44 
<< m1 >>
rect 105 43 106 44 
<< m2 >>
rect 105 43 106 44 
<< m1 >>
rect 106 43 107 44 
<< m2 >>
rect 106 43 107 44 
<< m1 >>
rect 107 43 108 44 
<< m1 >>
rect 108 43 109 44 
<< m1 >>
rect 109 43 110 44 
<< m2 >>
rect 109 43 110 44 
<< m1 >>
rect 110 43 111 44 
<< m1 >>
rect 111 43 112 44 
<< m1 >>
rect 112 43 113 44 
<< m1 >>
rect 113 43 114 44 
<< m1 >>
rect 114 43 115 44 
<< m1 >>
rect 115 43 116 44 
<< m1 >>
rect 116 43 117 44 
<< m1 >>
rect 117 43 118 44 
<< m1 >>
rect 118 43 119 44 
<< m2 >>
rect 118 43 119 44 
<< m1 >>
rect 119 43 120 44 
<< m1 >>
rect 120 43 121 44 
<< m1 >>
rect 121 43 122 44 
<< m1 >>
rect 122 43 123 44 
<< m1 >>
rect 123 43 124 44 
<< m1 >>
rect 124 43 125 44 
<< m2 >>
rect 125 43 126 44 
<< m2 >>
rect 128 43 129 44 
<< m2 >>
rect 130 43 131 44 
<< m2 >>
rect 131 43 132 44 
<< m2 >>
rect 132 43 133 44 
<< m2 >>
rect 133 43 134 44 
<< m2 >>
rect 134 43 135 44 
<< m2 >>
rect 135 43 136 44 
<< m1 >>
rect 136 43 137 44 
<< m2 >>
rect 136 43 137 44 
<< m2 >>
rect 137 43 138 44 
<< m1 >>
rect 138 43 139 44 
<< m2 >>
rect 138 43 139 44 
<< m2c >>
rect 138 43 139 44 
<< m1 >>
rect 138 43 139 44 
<< m2 >>
rect 138 43 139 44 
<< m1 >>
rect 139 43 140 44 
<< m1 >>
rect 140 43 141 44 
<< m2 >>
rect 140 43 141 44 
<< m2c >>
rect 140 43 141 44 
<< m1 >>
rect 140 43 141 44 
<< m2 >>
rect 140 43 141 44 
<< m2 >>
rect 141 43 142 44 
<< m1 >>
rect 142 43 143 44 
<< m2 >>
rect 142 43 143 44 
<< m1 >>
rect 143 43 144 44 
<< m2 >>
rect 143 43 144 44 
<< m1 >>
rect 144 43 145 44 
<< m2 >>
rect 144 43 145 44 
<< m1 >>
rect 145 43 146 44 
<< m2 >>
rect 145 43 146 44 
<< m1 >>
rect 146 43 147 44 
<< m2 >>
rect 146 43 147 44 
<< m1 >>
rect 147 43 148 44 
<< m1 >>
rect 148 43 149 44 
<< m2 >>
rect 148 43 149 44 
<< m2c >>
rect 148 43 149 44 
<< m1 >>
rect 148 43 149 44 
<< m2 >>
rect 148 43 149 44 
<< m1 >>
rect 150 43 151 44 
<< m2 >>
rect 150 43 151 44 
<< m2c >>
rect 150 43 151 44 
<< m1 >>
rect 150 43 151 44 
<< m2 >>
rect 150 43 151 44 
<< m1 >>
rect 152 43 153 44 
<< m2 >>
rect 152 43 153 44 
<< m2c >>
rect 152 43 153 44 
<< m1 >>
rect 152 43 153 44 
<< m2 >>
rect 152 43 153 44 
<< m2 >>
rect 153 43 154 44 
<< m1 >>
rect 154 43 155 44 
<< m2 >>
rect 154 43 155 44 
<< m2 >>
rect 155 43 156 44 
<< m1 >>
rect 156 43 157 44 
<< m2 >>
rect 156 43 157 44 
<< m2c >>
rect 156 43 157 44 
<< m1 >>
rect 156 43 157 44 
<< m2 >>
rect 156 43 157 44 
<< m1 >>
rect 157 43 158 44 
<< m1 >>
rect 158 43 159 44 
<< m1 >>
rect 159 43 160 44 
<< m1 >>
rect 160 43 161 44 
<< m1 >>
rect 161 43 162 44 
<< m2 >>
rect 161 43 162 44 
<< m2c >>
rect 161 43 162 44 
<< m1 >>
rect 161 43 162 44 
<< m2 >>
rect 161 43 162 44 
<< m2 >>
rect 162 43 163 44 
<< m1 >>
rect 163 43 164 44 
<< m2 >>
rect 163 43 164 44 
<< m2 >>
rect 164 43 165 44 
<< m1 >>
rect 165 43 166 44 
<< m2 >>
rect 165 43 166 44 
<< m2 >>
rect 166 43 167 44 
<< m1 >>
rect 167 43 168 44 
<< m2 >>
rect 167 43 168 44 
<< m2c >>
rect 167 43 168 44 
<< m1 >>
rect 167 43 168 44 
<< m2 >>
rect 167 43 168 44 
<< m1 >>
rect 168 43 169 44 
<< m1 >>
rect 169 43 170 44 
<< m1 >>
rect 170 43 171 44 
<< m2 >>
rect 170 43 171 44 
<< m2c >>
rect 170 43 171 44 
<< m1 >>
rect 170 43 171 44 
<< m2 >>
rect 170 43 171 44 
<< m2 >>
rect 171 43 172 44 
<< m1 >>
rect 172 43 173 44 
<< m2 >>
rect 172 43 173 44 
<< m1 >>
rect 173 43 174 44 
<< m2 >>
rect 173 43 174 44 
<< m1 >>
rect 174 43 175 44 
<< m2 >>
rect 174 43 175 44 
<< m1 >>
rect 175 43 176 44 
<< m2 >>
rect 175 43 176 44 
<< m1 >>
rect 176 43 177 44 
<< m2 >>
rect 176 43 177 44 
<< m1 >>
rect 177 43 178 44 
<< m2 >>
rect 177 43 178 44 
<< m1 >>
rect 178 43 179 44 
<< m2 >>
rect 178 43 179 44 
<< m2 >>
rect 179 43 180 44 
<< m1 >>
rect 186 43 187 44 
<< m1 >>
rect 190 43 191 44 
<< m2 >>
rect 190 43 191 44 
<< m1 >>
rect 191 43 192 44 
<< m1 >>
rect 192 43 193 44 
<< m1 >>
rect 193 43 194 44 
<< m1 >>
rect 194 43 195 44 
<< m1 >>
rect 195 43 196 44 
<< m1 >>
rect 196 43 197 44 
<< m1 >>
rect 197 43 198 44 
<< m2 >>
rect 197 43 198 44 
<< m2c >>
rect 197 43 198 44 
<< m1 >>
rect 197 43 198 44 
<< m2 >>
rect 197 43 198 44 
<< m2 >>
rect 198 43 199 44 
<< m1 >>
rect 199 43 200 44 
<< m2 >>
rect 199 43 200 44 
<< m2 >>
rect 200 43 201 44 
<< m1 >>
rect 201 43 202 44 
<< m2 >>
rect 201 43 202 44 
<< m2c >>
rect 201 43 202 44 
<< m1 >>
rect 201 43 202 44 
<< m2 >>
rect 201 43 202 44 
<< m1 >>
rect 202 43 203 44 
<< m1 >>
rect 203 43 204 44 
<< m2 >>
rect 203 43 204 44 
<< m1 >>
rect 204 43 205 44 
<< m1 >>
rect 205 43 206 44 
<< m1 >>
rect 206 43 207 44 
<< m1 >>
rect 207 43 208 44 
<< m1 >>
rect 208 43 209 44 
<< m1 >>
rect 209 43 210 44 
<< m1 >>
rect 210 43 211 44 
<< m1 >>
rect 211 43 212 44 
<< m1 >>
rect 212 43 213 44 
<< m1 >>
rect 213 43 214 44 
<< m1 >>
rect 214 43 215 44 
<< m1 >>
rect 232 43 233 44 
<< m2 >>
rect 232 43 233 44 
<< m2c >>
rect 232 43 233 44 
<< m1 >>
rect 232 43 233 44 
<< m2 >>
rect 232 43 233 44 
<< m2 >>
rect 243 43 244 44 
<< m1 >>
rect 244 43 245 44 
<< m2 >>
rect 244 43 245 44 
<< m1 >>
rect 245 43 246 44 
<< m2 >>
rect 245 43 246 44 
<< m1 >>
rect 246 43 247 44 
<< m2 >>
rect 246 43 247 44 
<< m1 >>
rect 247 43 248 44 
<< m2 >>
rect 247 43 248 44 
<< m1 >>
rect 248 43 249 44 
<< m2 >>
rect 248 43 249 44 
<< m1 >>
rect 249 43 250 44 
<< m2 >>
rect 249 43 250 44 
<< m1 >>
rect 250 43 251 44 
<< m2 >>
rect 250 43 251 44 
<< m1 >>
rect 251 43 252 44 
<< m2 >>
rect 251 43 252 44 
<< m1 >>
rect 252 43 253 44 
<< m2 >>
rect 252 43 253 44 
<< m1 >>
rect 253 43 254 44 
<< m2 >>
rect 253 43 254 44 
<< m1 >>
rect 254 43 255 44 
<< m2 >>
rect 254 43 255 44 
<< m2 >>
rect 255 43 256 44 
<< m1 >>
rect 256 43 257 44 
<< m2 >>
rect 256 43 257 44 
<< m2c >>
rect 256 43 257 44 
<< m1 >>
rect 256 43 257 44 
<< m2 >>
rect 256 43 257 44 
<< m1 >>
rect 26 44 27 45 
<< m1 >>
rect 28 44 29 45 
<< m2 >>
rect 28 44 29 45 
<< m2c >>
rect 28 44 29 45 
<< m1 >>
rect 28 44 29 45 
<< m2 >>
rect 28 44 29 45 
<< m1 >>
rect 37 44 38 45 
<< m1 >>
rect 40 44 41 45 
<< m2 >>
rect 43 44 44 45 
<< m1 >>
rect 44 44 45 45 
<< m1 >>
rect 58 44 59 45 
<< m1 >>
rect 60 44 61 45 
<< m1 >>
rect 73 44 74 45 
<< m1 >>
rect 75 44 76 45 
<< m2 >>
rect 76 44 77 45 
<< m2 >>
rect 87 44 88 45 
<< m1 >>
rect 91 44 92 45 
<< m2 >>
rect 106 44 107 45 
<< m2 >>
rect 109 44 110 45 
<< m2 >>
rect 118 44 119 45 
<< m2 >>
rect 125 44 126 45 
<< m1 >>
rect 126 44 127 45 
<< m2 >>
rect 126 44 127 45 
<< m2c >>
rect 126 44 127 45 
<< m1 >>
rect 126 44 127 45 
<< m2 >>
rect 126 44 127 45 
<< m1 >>
rect 127 44 128 45 
<< m1 >>
rect 128 44 129 45 
<< m2 >>
rect 128 44 129 45 
<< m1 >>
rect 129 44 130 45 
<< m1 >>
rect 130 44 131 45 
<< m2 >>
rect 130 44 131 45 
<< m1 >>
rect 131 44 132 45 
<< m1 >>
rect 132 44 133 45 
<< m1 >>
rect 133 44 134 45 
<< m1 >>
rect 134 44 135 45 
<< m1 >>
rect 136 44 137 45 
<< m2 >>
rect 137 44 138 45 
<< m1 >>
rect 142 44 143 45 
<< m1 >>
rect 150 44 151 45 
<< m1 >>
rect 152 44 153 45 
<< m1 >>
rect 154 44 155 45 
<< m1 >>
rect 163 44 164 45 
<< m1 >>
rect 165 44 166 45 
<< m1 >>
rect 172 44 173 45 
<< m2 >>
rect 179 44 180 45 
<< m1 >>
rect 186 44 187 45 
<< m1 >>
rect 190 44 191 45 
<< m2 >>
rect 190 44 191 45 
<< m1 >>
rect 199 44 200 45 
<< m2 >>
rect 203 44 204 45 
<< m1 >>
rect 214 44 215 45 
<< m2 >>
rect 232 44 233 45 
<< m2 >>
rect 243 44 244 45 
<< m1 >>
rect 254 44 255 45 
<< m1 >>
rect 256 44 257 45 
<< m1 >>
rect 26 45 27 46 
<< m2 >>
rect 28 45 29 46 
<< m1 >>
rect 37 45 38 46 
<< m1 >>
rect 40 45 41 46 
<< m2 >>
rect 43 45 44 46 
<< m1 >>
rect 44 45 45 46 
<< m1 >>
rect 58 45 59 46 
<< m1 >>
rect 60 45 61 46 
<< m1 >>
rect 73 45 74 46 
<< m1 >>
rect 75 45 76 46 
<< m2 >>
rect 76 45 77 46 
<< m1 >>
rect 87 45 88 46 
<< m2 >>
rect 87 45 88 46 
<< m2c >>
rect 87 45 88 46 
<< m1 >>
rect 87 45 88 46 
<< m2 >>
rect 87 45 88 46 
<< m1 >>
rect 88 45 89 46 
<< m1 >>
rect 89 45 90 46 
<< m1 >>
rect 91 45 92 46 
<< m1 >>
rect 106 45 107 46 
<< m2 >>
rect 106 45 107 46 
<< m2c >>
rect 106 45 107 46 
<< m1 >>
rect 106 45 107 46 
<< m2 >>
rect 106 45 107 46 
<< m2 >>
rect 109 45 110 46 
<< m2 >>
rect 118 45 119 46 
<< m2 >>
rect 128 45 129 46 
<< m2 >>
rect 130 45 131 46 
<< m1 >>
rect 134 45 135 46 
<< m1 >>
rect 136 45 137 46 
<< m2 >>
rect 137 45 138 46 
<< m1 >>
rect 142 45 143 46 
<< m1 >>
rect 148 45 149 46 
<< m2 >>
rect 148 45 149 46 
<< m2c >>
rect 148 45 149 46 
<< m1 >>
rect 148 45 149 46 
<< m2 >>
rect 148 45 149 46 
<< m2 >>
rect 149 45 150 46 
<< m1 >>
rect 150 45 151 46 
<< m2 >>
rect 150 45 151 46 
<< m2 >>
rect 151 45 152 46 
<< m1 >>
rect 152 45 153 46 
<< m2 >>
rect 152 45 153 46 
<< m2c >>
rect 152 45 153 46 
<< m1 >>
rect 152 45 153 46 
<< m2 >>
rect 152 45 153 46 
<< m1 >>
rect 154 45 155 46 
<< m1 >>
rect 163 45 164 46 
<< m1 >>
rect 165 45 166 46 
<< m1 >>
rect 172 45 173 46 
<< m1 >>
rect 175 45 176 46 
<< m1 >>
rect 176 45 177 46 
<< m1 >>
rect 177 45 178 46 
<< m1 >>
rect 178 45 179 46 
<< m1 >>
rect 179 45 180 46 
<< m2 >>
rect 179 45 180 46 
<< m1 >>
rect 180 45 181 46 
<< m1 >>
rect 181 45 182 46 
<< m1 >>
rect 186 45 187 46 
<< m1 >>
rect 190 45 191 46 
<< m2 >>
rect 190 45 191 46 
<< m1 >>
rect 199 45 200 46 
<< m2 >>
rect 203 45 204 46 
<< m1 >>
rect 204 45 205 46 
<< m2 >>
rect 204 45 205 46 
<< m2c >>
rect 204 45 205 46 
<< m1 >>
rect 204 45 205 46 
<< m2 >>
rect 204 45 205 46 
<< m1 >>
rect 214 45 215 46 
<< m1 >>
rect 229 45 230 46 
<< m1 >>
rect 230 45 231 46 
<< m1 >>
rect 231 45 232 46 
<< m1 >>
rect 232 45 233 46 
<< m2 >>
rect 232 45 233 46 
<< m1 >>
rect 233 45 234 46 
<< m1 >>
rect 234 45 235 46 
<< m1 >>
rect 235 45 236 46 
<< m1 >>
rect 236 45 237 46 
<< m1 >>
rect 237 45 238 46 
<< m1 >>
rect 238 45 239 46 
<< m1 >>
rect 239 45 240 46 
<< m1 >>
rect 240 45 241 46 
<< m1 >>
rect 241 45 242 46 
<< m1 >>
rect 242 45 243 46 
<< m1 >>
rect 243 45 244 46 
<< m2 >>
rect 243 45 244 46 
<< m1 >>
rect 254 45 255 46 
<< m1 >>
rect 256 45 257 46 
<< m1 >>
rect 26 46 27 47 
<< m1 >>
rect 28 46 29 47 
<< m2 >>
rect 28 46 29 47 
<< m1 >>
rect 29 46 30 47 
<< m1 >>
rect 30 46 31 47 
<< m1 >>
rect 31 46 32 47 
<< m1 >>
rect 37 46 38 47 
<< m1 >>
rect 40 46 41 47 
<< m2 >>
rect 43 46 44 47 
<< m1 >>
rect 44 46 45 47 
<< m1 >>
rect 46 46 47 47 
<< m1 >>
rect 47 46 48 47 
<< m1 >>
rect 48 46 49 47 
<< m1 >>
rect 49 46 50 47 
<< m1 >>
rect 58 46 59 47 
<< m1 >>
rect 60 46 61 47 
<< m1 >>
rect 73 46 74 47 
<< m1 >>
rect 75 46 76 47 
<< m2 >>
rect 76 46 77 47 
<< m1 >>
rect 82 46 83 47 
<< m1 >>
rect 83 46 84 47 
<< m1 >>
rect 84 46 85 47 
<< m1 >>
rect 85 46 86 47 
<< m1 >>
rect 89 46 90 47 
<< m2 >>
rect 89 46 90 47 
<< m2c >>
rect 89 46 90 47 
<< m1 >>
rect 89 46 90 47 
<< m2 >>
rect 89 46 90 47 
<< m2 >>
rect 90 46 91 47 
<< m1 >>
rect 91 46 92 47 
<< m2 >>
rect 91 46 92 47 
<< m2 >>
rect 92 46 93 47 
<< m1 >>
rect 106 46 107 47 
<< m1 >>
rect 109 46 110 47 
<< m2 >>
rect 109 46 110 47 
<< m1 >>
rect 110 46 111 47 
<< m1 >>
rect 111 46 112 47 
<< m1 >>
rect 112 46 113 47 
<< m1 >>
rect 113 46 114 47 
<< m1 >>
rect 114 46 115 47 
<< m1 >>
rect 115 46 116 47 
<< m1 >>
rect 116 46 117 47 
<< m1 >>
rect 117 46 118 47 
<< m1 >>
rect 118 46 119 47 
<< m2 >>
rect 118 46 119 47 
<< m1 >>
rect 119 46 120 47 
<< m1 >>
rect 120 46 121 47 
<< m1 >>
rect 121 46 122 47 
<< m1 >>
rect 124 46 125 47 
<< m1 >>
rect 125 46 126 47 
<< m1 >>
rect 126 46 127 47 
<< m1 >>
rect 127 46 128 47 
<< m1 >>
rect 128 46 129 47 
<< m2 >>
rect 128 46 129 47 
<< m1 >>
rect 129 46 130 47 
<< m1 >>
rect 130 46 131 47 
<< m2 >>
rect 130 46 131 47 
<< m2c >>
rect 130 46 131 47 
<< m1 >>
rect 130 46 131 47 
<< m2 >>
rect 130 46 131 47 
<< m1 >>
rect 132 46 133 47 
<< m2 >>
rect 132 46 133 47 
<< m2c >>
rect 132 46 133 47 
<< m1 >>
rect 132 46 133 47 
<< m2 >>
rect 132 46 133 47 
<< m2 >>
rect 133 46 134 47 
<< m1 >>
rect 134 46 135 47 
<< m2 >>
rect 134 46 135 47 
<< m2 >>
rect 135 46 136 47 
<< m1 >>
rect 136 46 137 47 
<< m2 >>
rect 136 46 137 47 
<< m2 >>
rect 137 46 138 47 
<< m1 >>
rect 142 46 143 47 
<< m1 >>
rect 148 46 149 47 
<< m1 >>
rect 150 46 151 47 
<< m1 >>
rect 154 46 155 47 
<< m1 >>
rect 163 46 164 47 
<< m1 >>
rect 165 46 166 47 
<< m1 >>
rect 172 46 173 47 
<< m1 >>
rect 175 46 176 47 
<< m2 >>
rect 179 46 180 47 
<< m2 >>
rect 180 46 181 47 
<< m1 >>
rect 181 46 182 47 
<< m2 >>
rect 181 46 182 47 
<< m2 >>
rect 182 46 183 47 
<< m1 >>
rect 186 46 187 47 
<< m1 >>
rect 190 46 191 47 
<< m2 >>
rect 190 46 191 47 
<< m1 >>
rect 196 46 197 47 
<< m1 >>
rect 197 46 198 47 
<< m2 >>
rect 197 46 198 47 
<< m2c >>
rect 197 46 198 47 
<< m1 >>
rect 197 46 198 47 
<< m2 >>
rect 197 46 198 47 
<< m2 >>
rect 198 46 199 47 
<< m1 >>
rect 199 46 200 47 
<< m2 >>
rect 199 46 200 47 
<< m2 >>
rect 200 46 201 47 
<< m1 >>
rect 201 46 202 47 
<< m2 >>
rect 201 46 202 47 
<< m2c >>
rect 201 46 202 47 
<< m1 >>
rect 201 46 202 47 
<< m2 >>
rect 201 46 202 47 
<< m1 >>
rect 202 46 203 47 
<< m1 >>
rect 204 46 205 47 
<< m1 >>
rect 214 46 215 47 
<< m1 >>
rect 229 46 230 47 
<< m2 >>
rect 232 46 233 47 
<< m1 >>
rect 243 46 244 47 
<< m2 >>
rect 243 46 244 47 
<< m1 >>
rect 254 46 255 47 
<< m1 >>
rect 256 46 257 47 
<< m1 >>
rect 26 47 27 48 
<< m1 >>
rect 28 47 29 48 
<< m2 >>
rect 28 47 29 48 
<< m1 >>
rect 31 47 32 48 
<< m1 >>
rect 37 47 38 48 
<< m1 >>
rect 40 47 41 48 
<< m2 >>
rect 43 47 44 48 
<< m1 >>
rect 44 47 45 48 
<< m1 >>
rect 46 47 47 48 
<< m1 >>
rect 49 47 50 48 
<< m1 >>
rect 58 47 59 48 
<< m1 >>
rect 60 47 61 48 
<< m1 >>
rect 73 47 74 48 
<< m1 >>
rect 75 47 76 48 
<< m2 >>
rect 76 47 77 48 
<< m1 >>
rect 82 47 83 48 
<< m1 >>
rect 85 47 86 48 
<< m1 >>
rect 91 47 92 48 
<< m2 >>
rect 92 47 93 48 
<< m1 >>
rect 106 47 107 48 
<< m1 >>
rect 109 47 110 48 
<< m2 >>
rect 109 47 110 48 
<< m2 >>
rect 118 47 119 48 
<< m1 >>
rect 121 47 122 48 
<< m1 >>
rect 124 47 125 48 
<< m2 >>
rect 128 47 129 48 
<< m1 >>
rect 132 47 133 48 
<< m1 >>
rect 134 47 135 48 
<< m1 >>
rect 136 47 137 48 
<< m1 >>
rect 142 47 143 48 
<< m1 >>
rect 148 47 149 48 
<< m1 >>
rect 150 47 151 48 
<< m1 >>
rect 154 47 155 48 
<< m1 >>
rect 163 47 164 48 
<< m1 >>
rect 165 47 166 48 
<< m1 >>
rect 172 47 173 48 
<< m1 >>
rect 175 47 176 48 
<< m1 >>
rect 181 47 182 48 
<< m2 >>
rect 182 47 183 48 
<< m1 >>
rect 186 47 187 48 
<< m1 >>
rect 190 47 191 48 
<< m2 >>
rect 190 47 191 48 
<< m1 >>
rect 196 47 197 48 
<< m1 >>
rect 199 47 200 48 
<< m1 >>
rect 202 47 203 48 
<< m1 >>
rect 204 47 205 48 
<< m1 >>
rect 214 47 215 48 
<< m1 >>
rect 229 47 230 48 
<< m1 >>
rect 232 47 233 48 
<< m2 >>
rect 232 47 233 48 
<< m1 >>
rect 243 47 244 48 
<< m2 >>
rect 243 47 244 48 
<< m1 >>
rect 254 47 255 48 
<< m1 >>
rect 256 47 257 48 
<< pdiffusion >>
rect 12 48 13 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< m1 >>
rect 26 48 27 49 
<< m1 >>
rect 28 48 29 49 
<< m2 >>
rect 28 48 29 49 
<< pdiffusion >>
rect 30 48 31 49 
<< m1 >>
rect 31 48 32 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< m1 >>
rect 37 48 38 49 
<< m1 >>
rect 40 48 41 49 
<< m2 >>
rect 43 48 44 49 
<< m1 >>
rect 44 48 45 49 
<< m1 >>
rect 46 48 47 49 
<< pdiffusion >>
rect 48 48 49 49 
<< m1 >>
rect 49 48 50 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 58 48 59 49 
<< m1 >>
rect 60 48 61 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< m1 >>
rect 73 48 74 49 
<< m1 >>
rect 75 48 76 49 
<< m2 >>
rect 76 48 77 49 
<< m1 >>
rect 82 48 83 49 
<< pdiffusion >>
rect 84 48 85 49 
<< m1 >>
rect 85 48 86 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< m2 >>
rect 92 48 93 49 
<< pdiffusion >>
rect 102 48 103 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< m1 >>
rect 106 48 107 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< m1 >>
rect 109 48 110 49 
<< m2 >>
rect 109 48 110 49 
<< m2 >>
rect 110 48 111 49 
<< m1 >>
rect 111 48 112 49 
<< m2 >>
rect 111 48 112 49 
<< m2c >>
rect 111 48 112 49 
<< m1 >>
rect 111 48 112 49 
<< m2 >>
rect 111 48 112 49 
<< m1 >>
rect 112 48 113 49 
<< m1 >>
rect 113 48 114 49 
<< m1 >>
rect 118 48 119 49 
<< m2 >>
rect 118 48 119 49 
<< m2c >>
rect 118 48 119 49 
<< m1 >>
rect 118 48 119 49 
<< m2 >>
rect 118 48 119 49 
<< pdiffusion >>
rect 120 48 121 49 
<< m1 >>
rect 121 48 122 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< m1 >>
rect 124 48 125 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< m1 >>
rect 128 48 129 49 
<< m2 >>
rect 128 48 129 49 
<< m2c >>
rect 128 48 129 49 
<< m1 >>
rect 128 48 129 49 
<< m2 >>
rect 128 48 129 49 
<< m1 >>
rect 132 48 133 49 
<< m1 >>
rect 134 48 135 49 
<< m1 >>
rect 136 48 137 49 
<< pdiffusion >>
rect 138 48 139 49 
<< pdiffusion >>
rect 139 48 140 49 
<< pdiffusion >>
rect 140 48 141 49 
<< pdiffusion >>
rect 141 48 142 49 
<< m1 >>
rect 142 48 143 49 
<< pdiffusion >>
rect 142 48 143 49 
<< pdiffusion >>
rect 143 48 144 49 
<< m1 >>
rect 148 48 149 49 
<< m1 >>
rect 150 48 151 49 
<< m1 >>
rect 154 48 155 49 
<< pdiffusion >>
rect 156 48 157 49 
<< pdiffusion >>
rect 157 48 158 49 
<< pdiffusion >>
rect 158 48 159 49 
<< pdiffusion >>
rect 159 48 160 49 
<< pdiffusion >>
rect 160 48 161 49 
<< pdiffusion >>
rect 161 48 162 49 
<< m1 >>
rect 163 48 164 49 
<< m1 >>
rect 165 48 166 49 
<< m1 >>
rect 172 48 173 49 
<< pdiffusion >>
rect 174 48 175 49 
<< m1 >>
rect 175 48 176 49 
<< pdiffusion >>
rect 175 48 176 49 
<< pdiffusion >>
rect 176 48 177 49 
<< pdiffusion >>
rect 177 48 178 49 
<< pdiffusion >>
rect 178 48 179 49 
<< pdiffusion >>
rect 179 48 180 49 
<< m1 >>
rect 181 48 182 49 
<< m2 >>
rect 182 48 183 49 
<< m1 >>
rect 186 48 187 49 
<< m1 >>
rect 190 48 191 49 
<< m2 >>
rect 190 48 191 49 
<< pdiffusion >>
rect 192 48 193 49 
<< pdiffusion >>
rect 193 48 194 49 
<< pdiffusion >>
rect 194 48 195 49 
<< pdiffusion >>
rect 195 48 196 49 
<< m1 >>
rect 196 48 197 49 
<< pdiffusion >>
rect 196 48 197 49 
<< pdiffusion >>
rect 197 48 198 49 
<< m1 >>
rect 199 48 200 49 
<< m1 >>
rect 202 48 203 49 
<< m1 >>
rect 204 48 205 49 
<< pdiffusion >>
rect 210 48 211 49 
<< pdiffusion >>
rect 211 48 212 49 
<< pdiffusion >>
rect 212 48 213 49 
<< pdiffusion >>
rect 213 48 214 49 
<< m1 >>
rect 214 48 215 49 
<< pdiffusion >>
rect 214 48 215 49 
<< pdiffusion >>
rect 215 48 216 49 
<< pdiffusion >>
rect 228 48 229 49 
<< m1 >>
rect 229 48 230 49 
<< pdiffusion >>
rect 229 48 230 49 
<< pdiffusion >>
rect 230 48 231 49 
<< m1 >>
rect 231 48 232 49 
<< m2 >>
rect 231 48 232 49 
<< m2c >>
rect 231 48 232 49 
<< m1 >>
rect 231 48 232 49 
<< m2 >>
rect 231 48 232 49 
<< pdiffusion >>
rect 231 48 232 49 
<< m1 >>
rect 232 48 233 49 
<< pdiffusion >>
rect 232 48 233 49 
<< pdiffusion >>
rect 233 48 234 49 
<< m1 >>
rect 243 48 244 49 
<< m2 >>
rect 243 48 244 49 
<< pdiffusion >>
rect 246 48 247 49 
<< pdiffusion >>
rect 247 48 248 49 
<< pdiffusion >>
rect 248 48 249 49 
<< pdiffusion >>
rect 249 48 250 49 
<< pdiffusion >>
rect 250 48 251 49 
<< pdiffusion >>
rect 251 48 252 49 
<< m1 >>
rect 254 48 255 49 
<< m1 >>
rect 256 48 257 49 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< m1 >>
rect 26 49 27 50 
<< m1 >>
rect 28 49 29 50 
<< m2 >>
rect 28 49 29 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< m1 >>
rect 37 49 38 50 
<< m1 >>
rect 40 49 41 50 
<< m2 >>
rect 43 49 44 50 
<< m1 >>
rect 44 49 45 50 
<< m1 >>
rect 46 49 47 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 58 49 59 50 
<< m1 >>
rect 60 49 61 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< m1 >>
rect 73 49 74 50 
<< m1 >>
rect 75 49 76 50 
<< m2 >>
rect 76 49 77 50 
<< m1 >>
rect 82 49 83 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< m2 >>
rect 92 49 93 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< m1 >>
rect 109 49 110 50 
<< m1 >>
rect 113 49 114 50 
<< m1 >>
rect 118 49 119 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< m1 >>
rect 128 49 129 50 
<< m1 >>
rect 132 49 133 50 
<< m1 >>
rect 134 49 135 50 
<< m1 >>
rect 136 49 137 50 
<< pdiffusion >>
rect 138 49 139 50 
<< pdiffusion >>
rect 139 49 140 50 
<< pdiffusion >>
rect 140 49 141 50 
<< pdiffusion >>
rect 141 49 142 50 
<< pdiffusion >>
rect 142 49 143 50 
<< pdiffusion >>
rect 143 49 144 50 
<< m1 >>
rect 148 49 149 50 
<< m1 >>
rect 150 49 151 50 
<< m1 >>
rect 154 49 155 50 
<< pdiffusion >>
rect 156 49 157 50 
<< pdiffusion >>
rect 157 49 158 50 
<< pdiffusion >>
rect 158 49 159 50 
<< pdiffusion >>
rect 159 49 160 50 
<< pdiffusion >>
rect 160 49 161 50 
<< pdiffusion >>
rect 161 49 162 50 
<< m1 >>
rect 163 49 164 50 
<< m1 >>
rect 165 49 166 50 
<< m1 >>
rect 172 49 173 50 
<< pdiffusion >>
rect 174 49 175 50 
<< pdiffusion >>
rect 175 49 176 50 
<< pdiffusion >>
rect 176 49 177 50 
<< pdiffusion >>
rect 177 49 178 50 
<< pdiffusion >>
rect 178 49 179 50 
<< pdiffusion >>
rect 179 49 180 50 
<< m1 >>
rect 181 49 182 50 
<< m2 >>
rect 182 49 183 50 
<< m1 >>
rect 186 49 187 50 
<< m1 >>
rect 190 49 191 50 
<< m2 >>
rect 190 49 191 50 
<< pdiffusion >>
rect 192 49 193 50 
<< pdiffusion >>
rect 193 49 194 50 
<< pdiffusion >>
rect 194 49 195 50 
<< pdiffusion >>
rect 195 49 196 50 
<< pdiffusion >>
rect 196 49 197 50 
<< pdiffusion >>
rect 197 49 198 50 
<< m1 >>
rect 199 49 200 50 
<< m1 >>
rect 202 49 203 50 
<< m1 >>
rect 204 49 205 50 
<< pdiffusion >>
rect 210 49 211 50 
<< pdiffusion >>
rect 211 49 212 50 
<< pdiffusion >>
rect 212 49 213 50 
<< pdiffusion >>
rect 213 49 214 50 
<< pdiffusion >>
rect 214 49 215 50 
<< pdiffusion >>
rect 215 49 216 50 
<< pdiffusion >>
rect 228 49 229 50 
<< pdiffusion >>
rect 229 49 230 50 
<< pdiffusion >>
rect 230 49 231 50 
<< pdiffusion >>
rect 231 49 232 50 
<< pdiffusion >>
rect 232 49 233 50 
<< pdiffusion >>
rect 233 49 234 50 
<< m1 >>
rect 243 49 244 50 
<< m2 >>
rect 243 49 244 50 
<< pdiffusion >>
rect 246 49 247 50 
<< pdiffusion >>
rect 247 49 248 50 
<< pdiffusion >>
rect 248 49 249 50 
<< pdiffusion >>
rect 249 49 250 50 
<< pdiffusion >>
rect 250 49 251 50 
<< pdiffusion >>
rect 251 49 252 50 
<< m1 >>
rect 254 49 255 50 
<< m1 >>
rect 256 49 257 50 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< m1 >>
rect 26 50 27 51 
<< m1 >>
rect 28 50 29 51 
<< m2 >>
rect 28 50 29 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< m1 >>
rect 37 50 38 51 
<< m1 >>
rect 40 50 41 51 
<< m2 >>
rect 43 50 44 51 
<< m1 >>
rect 44 50 45 51 
<< m1 >>
rect 46 50 47 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 58 50 59 51 
<< m1 >>
rect 60 50 61 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< m1 >>
rect 73 50 74 51 
<< m1 >>
rect 75 50 76 51 
<< m2 >>
rect 76 50 77 51 
<< m1 >>
rect 82 50 83 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< m2 >>
rect 92 50 93 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< m1 >>
rect 109 50 110 51 
<< m1 >>
rect 113 50 114 51 
<< m1 >>
rect 118 50 119 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< m1 >>
rect 128 50 129 51 
<< m1 >>
rect 132 50 133 51 
<< m1 >>
rect 134 50 135 51 
<< m1 >>
rect 136 50 137 51 
<< pdiffusion >>
rect 138 50 139 51 
<< pdiffusion >>
rect 139 50 140 51 
<< pdiffusion >>
rect 140 50 141 51 
<< pdiffusion >>
rect 141 50 142 51 
<< pdiffusion >>
rect 142 50 143 51 
<< pdiffusion >>
rect 143 50 144 51 
<< m1 >>
rect 148 50 149 51 
<< m1 >>
rect 150 50 151 51 
<< m1 >>
rect 154 50 155 51 
<< pdiffusion >>
rect 156 50 157 51 
<< pdiffusion >>
rect 157 50 158 51 
<< pdiffusion >>
rect 158 50 159 51 
<< pdiffusion >>
rect 159 50 160 51 
<< pdiffusion >>
rect 160 50 161 51 
<< pdiffusion >>
rect 161 50 162 51 
<< m1 >>
rect 163 50 164 51 
<< m1 >>
rect 165 50 166 51 
<< m1 >>
rect 172 50 173 51 
<< pdiffusion >>
rect 174 50 175 51 
<< pdiffusion >>
rect 175 50 176 51 
<< pdiffusion >>
rect 176 50 177 51 
<< pdiffusion >>
rect 177 50 178 51 
<< pdiffusion >>
rect 178 50 179 51 
<< pdiffusion >>
rect 179 50 180 51 
<< m1 >>
rect 181 50 182 51 
<< m2 >>
rect 182 50 183 51 
<< m1 >>
rect 186 50 187 51 
<< m1 >>
rect 190 50 191 51 
<< m2 >>
rect 190 50 191 51 
<< pdiffusion >>
rect 192 50 193 51 
<< pdiffusion >>
rect 193 50 194 51 
<< pdiffusion >>
rect 194 50 195 51 
<< pdiffusion >>
rect 195 50 196 51 
<< pdiffusion >>
rect 196 50 197 51 
<< pdiffusion >>
rect 197 50 198 51 
<< m1 >>
rect 199 50 200 51 
<< m1 >>
rect 202 50 203 51 
<< m1 >>
rect 204 50 205 51 
<< pdiffusion >>
rect 210 50 211 51 
<< pdiffusion >>
rect 211 50 212 51 
<< pdiffusion >>
rect 212 50 213 51 
<< pdiffusion >>
rect 213 50 214 51 
<< pdiffusion >>
rect 214 50 215 51 
<< pdiffusion >>
rect 215 50 216 51 
<< pdiffusion >>
rect 228 50 229 51 
<< pdiffusion >>
rect 229 50 230 51 
<< pdiffusion >>
rect 230 50 231 51 
<< pdiffusion >>
rect 231 50 232 51 
<< pdiffusion >>
rect 232 50 233 51 
<< pdiffusion >>
rect 233 50 234 51 
<< m1 >>
rect 243 50 244 51 
<< m2 >>
rect 243 50 244 51 
<< pdiffusion >>
rect 246 50 247 51 
<< pdiffusion >>
rect 247 50 248 51 
<< pdiffusion >>
rect 248 50 249 51 
<< pdiffusion >>
rect 249 50 250 51 
<< pdiffusion >>
rect 250 50 251 51 
<< pdiffusion >>
rect 251 50 252 51 
<< m1 >>
rect 254 50 255 51 
<< m1 >>
rect 256 50 257 51 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< m1 >>
rect 26 51 27 52 
<< m1 >>
rect 28 51 29 52 
<< m2 >>
rect 28 51 29 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< m1 >>
rect 37 51 38 52 
<< m1 >>
rect 40 51 41 52 
<< m2 >>
rect 43 51 44 52 
<< m1 >>
rect 44 51 45 52 
<< m1 >>
rect 46 51 47 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 58 51 59 52 
<< m1 >>
rect 60 51 61 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< m1 >>
rect 73 51 74 52 
<< m1 >>
rect 75 51 76 52 
<< m2 >>
rect 76 51 77 52 
<< m1 >>
rect 82 51 83 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< m2 >>
rect 92 51 93 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< m1 >>
rect 109 51 110 52 
<< m1 >>
rect 113 51 114 52 
<< m1 >>
rect 118 51 119 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< m1 >>
rect 128 51 129 52 
<< m1 >>
rect 132 51 133 52 
<< m1 >>
rect 134 51 135 52 
<< m1 >>
rect 136 51 137 52 
<< pdiffusion >>
rect 138 51 139 52 
<< pdiffusion >>
rect 139 51 140 52 
<< pdiffusion >>
rect 140 51 141 52 
<< pdiffusion >>
rect 141 51 142 52 
<< pdiffusion >>
rect 142 51 143 52 
<< pdiffusion >>
rect 143 51 144 52 
<< m1 >>
rect 148 51 149 52 
<< m1 >>
rect 150 51 151 52 
<< m1 >>
rect 154 51 155 52 
<< pdiffusion >>
rect 156 51 157 52 
<< pdiffusion >>
rect 157 51 158 52 
<< pdiffusion >>
rect 158 51 159 52 
<< pdiffusion >>
rect 159 51 160 52 
<< pdiffusion >>
rect 160 51 161 52 
<< pdiffusion >>
rect 161 51 162 52 
<< m1 >>
rect 163 51 164 52 
<< m1 >>
rect 165 51 166 52 
<< m1 >>
rect 172 51 173 52 
<< pdiffusion >>
rect 174 51 175 52 
<< pdiffusion >>
rect 175 51 176 52 
<< pdiffusion >>
rect 176 51 177 52 
<< pdiffusion >>
rect 177 51 178 52 
<< pdiffusion >>
rect 178 51 179 52 
<< pdiffusion >>
rect 179 51 180 52 
<< m1 >>
rect 181 51 182 52 
<< m2 >>
rect 182 51 183 52 
<< m1 >>
rect 186 51 187 52 
<< m1 >>
rect 190 51 191 52 
<< m2 >>
rect 190 51 191 52 
<< pdiffusion >>
rect 192 51 193 52 
<< pdiffusion >>
rect 193 51 194 52 
<< pdiffusion >>
rect 194 51 195 52 
<< pdiffusion >>
rect 195 51 196 52 
<< pdiffusion >>
rect 196 51 197 52 
<< pdiffusion >>
rect 197 51 198 52 
<< m1 >>
rect 199 51 200 52 
<< m1 >>
rect 202 51 203 52 
<< m1 >>
rect 204 51 205 52 
<< pdiffusion >>
rect 210 51 211 52 
<< pdiffusion >>
rect 211 51 212 52 
<< pdiffusion >>
rect 212 51 213 52 
<< pdiffusion >>
rect 213 51 214 52 
<< pdiffusion >>
rect 214 51 215 52 
<< pdiffusion >>
rect 215 51 216 52 
<< pdiffusion >>
rect 228 51 229 52 
<< pdiffusion >>
rect 229 51 230 52 
<< pdiffusion >>
rect 230 51 231 52 
<< pdiffusion >>
rect 231 51 232 52 
<< pdiffusion >>
rect 232 51 233 52 
<< pdiffusion >>
rect 233 51 234 52 
<< m1 >>
rect 243 51 244 52 
<< m2 >>
rect 243 51 244 52 
<< pdiffusion >>
rect 246 51 247 52 
<< pdiffusion >>
rect 247 51 248 52 
<< pdiffusion >>
rect 248 51 249 52 
<< pdiffusion >>
rect 249 51 250 52 
<< pdiffusion >>
rect 250 51 251 52 
<< pdiffusion >>
rect 251 51 252 52 
<< m1 >>
rect 254 51 255 52 
<< m1 >>
rect 256 51 257 52 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< m1 >>
rect 26 52 27 53 
<< m1 >>
rect 28 52 29 53 
<< m2 >>
rect 28 52 29 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< m1 >>
rect 37 52 38 53 
<< m1 >>
rect 40 52 41 53 
<< m2 >>
rect 43 52 44 53 
<< m1 >>
rect 44 52 45 53 
<< m1 >>
rect 46 52 47 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 58 52 59 53 
<< m1 >>
rect 60 52 61 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< m1 >>
rect 73 52 74 53 
<< m1 >>
rect 75 52 76 53 
<< m2 >>
rect 76 52 77 53 
<< m1 >>
rect 82 52 83 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< m2 >>
rect 92 52 93 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< m1 >>
rect 109 52 110 53 
<< m1 >>
rect 113 52 114 53 
<< m1 >>
rect 118 52 119 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< m1 >>
rect 128 52 129 53 
<< m1 >>
rect 132 52 133 53 
<< m1 >>
rect 134 52 135 53 
<< m1 >>
rect 136 52 137 53 
<< pdiffusion >>
rect 138 52 139 53 
<< pdiffusion >>
rect 139 52 140 53 
<< pdiffusion >>
rect 140 52 141 53 
<< pdiffusion >>
rect 141 52 142 53 
<< pdiffusion >>
rect 142 52 143 53 
<< pdiffusion >>
rect 143 52 144 53 
<< m1 >>
rect 148 52 149 53 
<< m1 >>
rect 150 52 151 53 
<< m1 >>
rect 154 52 155 53 
<< pdiffusion >>
rect 156 52 157 53 
<< pdiffusion >>
rect 157 52 158 53 
<< pdiffusion >>
rect 158 52 159 53 
<< pdiffusion >>
rect 159 52 160 53 
<< pdiffusion >>
rect 160 52 161 53 
<< pdiffusion >>
rect 161 52 162 53 
<< m1 >>
rect 163 52 164 53 
<< m1 >>
rect 165 52 166 53 
<< m1 >>
rect 172 52 173 53 
<< pdiffusion >>
rect 174 52 175 53 
<< pdiffusion >>
rect 175 52 176 53 
<< pdiffusion >>
rect 176 52 177 53 
<< pdiffusion >>
rect 177 52 178 53 
<< pdiffusion >>
rect 178 52 179 53 
<< pdiffusion >>
rect 179 52 180 53 
<< m1 >>
rect 181 52 182 53 
<< m2 >>
rect 182 52 183 53 
<< m1 >>
rect 186 52 187 53 
<< m1 >>
rect 190 52 191 53 
<< m2 >>
rect 190 52 191 53 
<< pdiffusion >>
rect 192 52 193 53 
<< pdiffusion >>
rect 193 52 194 53 
<< pdiffusion >>
rect 194 52 195 53 
<< pdiffusion >>
rect 195 52 196 53 
<< pdiffusion >>
rect 196 52 197 53 
<< pdiffusion >>
rect 197 52 198 53 
<< m1 >>
rect 199 52 200 53 
<< m1 >>
rect 202 52 203 53 
<< m1 >>
rect 204 52 205 53 
<< pdiffusion >>
rect 210 52 211 53 
<< pdiffusion >>
rect 211 52 212 53 
<< pdiffusion >>
rect 212 52 213 53 
<< pdiffusion >>
rect 213 52 214 53 
<< pdiffusion >>
rect 214 52 215 53 
<< pdiffusion >>
rect 215 52 216 53 
<< pdiffusion >>
rect 228 52 229 53 
<< pdiffusion >>
rect 229 52 230 53 
<< pdiffusion >>
rect 230 52 231 53 
<< pdiffusion >>
rect 231 52 232 53 
<< pdiffusion >>
rect 232 52 233 53 
<< pdiffusion >>
rect 233 52 234 53 
<< m1 >>
rect 243 52 244 53 
<< m2 >>
rect 243 52 244 53 
<< pdiffusion >>
rect 246 52 247 53 
<< pdiffusion >>
rect 247 52 248 53 
<< pdiffusion >>
rect 248 52 249 53 
<< pdiffusion >>
rect 249 52 250 53 
<< pdiffusion >>
rect 250 52 251 53 
<< pdiffusion >>
rect 251 52 252 53 
<< m1 >>
rect 254 52 255 53 
<< m1 >>
rect 256 52 257 53 
<< pdiffusion >>
rect 12 53 13 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< m1 >>
rect 26 53 27 54 
<< m1 >>
rect 28 53 29 54 
<< m2 >>
rect 28 53 29 54 
<< pdiffusion >>
rect 30 53 31 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< m1 >>
rect 37 53 38 54 
<< m1 >>
rect 40 53 41 54 
<< m2 >>
rect 43 53 44 54 
<< m1 >>
rect 44 53 45 54 
<< m1 >>
rect 46 53 47 54 
<< pdiffusion >>
rect 48 53 49 54 
<< m1 >>
rect 49 53 50 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 58 53 59 54 
<< m1 >>
rect 60 53 61 54 
<< pdiffusion >>
rect 66 53 67 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< m1 >>
rect 73 53 74 54 
<< m1 >>
rect 75 53 76 54 
<< m2 >>
rect 76 53 77 54 
<< m1 >>
rect 82 53 83 54 
<< pdiffusion >>
rect 84 53 85 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< m1 >>
rect 88 53 89 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< m2 >>
rect 92 53 93 54 
<< pdiffusion >>
rect 102 53 103 54 
<< m1 >>
rect 103 53 104 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< m1 >>
rect 106 53 107 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< m1 >>
rect 109 53 110 54 
<< m1 >>
rect 113 53 114 54 
<< m1 >>
rect 118 53 119 54 
<< pdiffusion >>
rect 120 53 121 54 
<< m1 >>
rect 121 53 122 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< m1 >>
rect 124 53 125 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< m1 >>
rect 128 53 129 54 
<< m1 >>
rect 129 53 130 54 
<< m1 >>
rect 130 53 131 54 
<< m2 >>
rect 130 53 131 54 
<< m2c >>
rect 130 53 131 54 
<< m1 >>
rect 130 53 131 54 
<< m2 >>
rect 130 53 131 54 
<< m2 >>
rect 131 53 132 54 
<< m1 >>
rect 132 53 133 54 
<< m2 >>
rect 132 53 133 54 
<< m2 >>
rect 133 53 134 54 
<< m1 >>
rect 134 53 135 54 
<< m2 >>
rect 134 53 135 54 
<< m2 >>
rect 135 53 136 54 
<< m1 >>
rect 136 53 137 54 
<< m2 >>
rect 136 53 137 54 
<< pdiffusion >>
rect 138 53 139 54 
<< m1 >>
rect 139 53 140 54 
<< pdiffusion >>
rect 139 53 140 54 
<< pdiffusion >>
rect 140 53 141 54 
<< pdiffusion >>
rect 141 53 142 54 
<< pdiffusion >>
rect 142 53 143 54 
<< pdiffusion >>
rect 143 53 144 54 
<< m1 >>
rect 148 53 149 54 
<< m1 >>
rect 150 53 151 54 
<< m1 >>
rect 154 53 155 54 
<< pdiffusion >>
rect 156 53 157 54 
<< pdiffusion >>
rect 157 53 158 54 
<< pdiffusion >>
rect 158 53 159 54 
<< pdiffusion >>
rect 159 53 160 54 
<< pdiffusion >>
rect 160 53 161 54 
<< pdiffusion >>
rect 161 53 162 54 
<< m1 >>
rect 163 53 164 54 
<< m1 >>
rect 165 53 166 54 
<< m1 >>
rect 172 53 173 54 
<< pdiffusion >>
rect 174 53 175 54 
<< pdiffusion >>
rect 175 53 176 54 
<< pdiffusion >>
rect 176 53 177 54 
<< pdiffusion >>
rect 177 53 178 54 
<< pdiffusion >>
rect 178 53 179 54 
<< pdiffusion >>
rect 179 53 180 54 
<< m1 >>
rect 181 53 182 54 
<< m2 >>
rect 182 53 183 54 
<< m1 >>
rect 186 53 187 54 
<< m1 >>
rect 190 53 191 54 
<< m2 >>
rect 190 53 191 54 
<< pdiffusion >>
rect 192 53 193 54 
<< pdiffusion >>
rect 193 53 194 54 
<< pdiffusion >>
rect 194 53 195 54 
<< pdiffusion >>
rect 195 53 196 54 
<< m1 >>
rect 196 53 197 54 
<< pdiffusion >>
rect 196 53 197 54 
<< pdiffusion >>
rect 197 53 198 54 
<< m1 >>
rect 199 53 200 54 
<< m1 >>
rect 202 53 203 54 
<< m1 >>
rect 204 53 205 54 
<< pdiffusion >>
rect 210 53 211 54 
<< pdiffusion >>
rect 211 53 212 54 
<< pdiffusion >>
rect 212 53 213 54 
<< pdiffusion >>
rect 213 53 214 54 
<< pdiffusion >>
rect 214 53 215 54 
<< pdiffusion >>
rect 215 53 216 54 
<< pdiffusion >>
rect 228 53 229 54 
<< pdiffusion >>
rect 229 53 230 54 
<< pdiffusion >>
rect 230 53 231 54 
<< pdiffusion >>
rect 231 53 232 54 
<< m1 >>
rect 232 53 233 54 
<< pdiffusion >>
rect 232 53 233 54 
<< pdiffusion >>
rect 233 53 234 54 
<< m1 >>
rect 243 53 244 54 
<< m2 >>
rect 243 53 244 54 
<< pdiffusion >>
rect 246 53 247 54 
<< pdiffusion >>
rect 247 53 248 54 
<< pdiffusion >>
rect 248 53 249 54 
<< pdiffusion >>
rect 249 53 250 54 
<< m1 >>
rect 250 53 251 54 
<< pdiffusion >>
rect 250 53 251 54 
<< pdiffusion >>
rect 251 53 252 54 
<< m1 >>
rect 254 53 255 54 
<< m1 >>
rect 256 53 257 54 
<< m1 >>
rect 26 54 27 55 
<< m1 >>
rect 28 54 29 55 
<< m2 >>
rect 28 54 29 55 
<< m1 >>
rect 37 54 38 55 
<< m1 >>
rect 40 54 41 55 
<< m2 >>
rect 43 54 44 55 
<< m1 >>
rect 44 54 45 55 
<< m1 >>
rect 46 54 47 55 
<< m1 >>
rect 49 54 50 55 
<< m1 >>
rect 58 54 59 55 
<< m1 >>
rect 60 54 61 55 
<< m1 >>
rect 73 54 74 55 
<< m1 >>
rect 75 54 76 55 
<< m2 >>
rect 76 54 77 55 
<< m1 >>
rect 82 54 83 55 
<< m1 >>
rect 88 54 89 55 
<< m1 >>
rect 91 54 92 55 
<< m2 >>
rect 92 54 93 55 
<< m1 >>
rect 103 54 104 55 
<< m1 >>
rect 106 54 107 55 
<< m1 >>
rect 109 54 110 55 
<< m1 >>
rect 113 54 114 55 
<< m1 >>
rect 118 54 119 55 
<< m1 >>
rect 121 54 122 55 
<< m1 >>
rect 124 54 125 55 
<< m1 >>
rect 132 54 133 55 
<< m1 >>
rect 134 54 135 55 
<< m1 >>
rect 136 54 137 55 
<< m2 >>
rect 136 54 137 55 
<< m1 >>
rect 139 54 140 55 
<< m1 >>
rect 148 54 149 55 
<< m1 >>
rect 150 54 151 55 
<< m1 >>
rect 154 54 155 55 
<< m1 >>
rect 163 54 164 55 
<< m1 >>
rect 165 54 166 55 
<< m1 >>
rect 172 54 173 55 
<< m1 >>
rect 181 54 182 55 
<< m2 >>
rect 182 54 183 55 
<< m1 >>
rect 183 54 184 55 
<< m2 >>
rect 183 54 184 55 
<< m2c >>
rect 183 54 184 55 
<< m1 >>
rect 183 54 184 55 
<< m2 >>
rect 183 54 184 55 
<< m1 >>
rect 186 54 187 55 
<< m1 >>
rect 190 54 191 55 
<< m2 >>
rect 190 54 191 55 
<< m1 >>
rect 196 54 197 55 
<< m1 >>
rect 199 54 200 55 
<< m1 >>
rect 202 54 203 55 
<< m1 >>
rect 204 54 205 55 
<< m1 >>
rect 232 54 233 55 
<< m1 >>
rect 235 54 236 55 
<< m1 >>
rect 236 54 237 55 
<< m1 >>
rect 237 54 238 55 
<< m1 >>
rect 238 54 239 55 
<< m1 >>
rect 239 54 240 55 
<< m1 >>
rect 240 54 241 55 
<< m1 >>
rect 241 54 242 55 
<< m2 >>
rect 241 54 242 55 
<< m2c >>
rect 241 54 242 55 
<< m1 >>
rect 241 54 242 55 
<< m2 >>
rect 241 54 242 55 
<< m2 >>
rect 242 54 243 55 
<< m1 >>
rect 243 54 244 55 
<< m2 >>
rect 243 54 244 55 
<< m1 >>
rect 250 54 251 55 
<< m1 >>
rect 254 54 255 55 
<< m1 >>
rect 256 54 257 55 
<< m1 >>
rect 26 55 27 56 
<< m1 >>
rect 28 55 29 56 
<< m2 >>
rect 28 55 29 56 
<< m1 >>
rect 37 55 38 56 
<< m1 >>
rect 40 55 41 56 
<< m2 >>
rect 43 55 44 56 
<< m1 >>
rect 44 55 45 56 
<< m1 >>
rect 46 55 47 56 
<< m1 >>
rect 49 55 50 56 
<< m1 >>
rect 58 55 59 56 
<< m1 >>
rect 60 55 61 56 
<< m1 >>
rect 71 55 72 56 
<< m2 >>
rect 71 55 72 56 
<< m2c >>
rect 71 55 72 56 
<< m1 >>
rect 71 55 72 56 
<< m2 >>
rect 71 55 72 56 
<< m2 >>
rect 72 55 73 56 
<< m1 >>
rect 73 55 74 56 
<< m2 >>
rect 73 55 74 56 
<< m2 >>
rect 74 55 75 56 
<< m1 >>
rect 75 55 76 56 
<< m2 >>
rect 75 55 76 56 
<< m2 >>
rect 76 55 77 56 
<< m1 >>
rect 82 55 83 56 
<< m1 >>
rect 88 55 89 56 
<< m1 >>
rect 89 55 90 56 
<< m1 >>
rect 90 55 91 56 
<< m1 >>
rect 91 55 92 56 
<< m2 >>
rect 92 55 93 56 
<< m1 >>
rect 93 55 94 56 
<< m2 >>
rect 93 55 94 56 
<< m2c >>
rect 93 55 94 56 
<< m1 >>
rect 93 55 94 56 
<< m2 >>
rect 93 55 94 56 
<< m1 >>
rect 94 55 95 56 
<< m1 >>
rect 95 55 96 56 
<< m1 >>
rect 96 55 97 56 
<< m1 >>
rect 97 55 98 56 
<< m1 >>
rect 98 55 99 56 
<< m1 >>
rect 99 55 100 56 
<< m1 >>
rect 100 55 101 56 
<< m1 >>
rect 101 55 102 56 
<< m1 >>
rect 102 55 103 56 
<< m1 >>
rect 103 55 104 56 
<< m1 >>
rect 106 55 107 56 
<< m1 >>
rect 109 55 110 56 
<< m1 >>
rect 113 55 114 56 
<< m1 >>
rect 118 55 119 56 
<< m1 >>
rect 121 55 122 56 
<< m1 >>
rect 124 55 125 56 
<< m2 >>
rect 125 55 126 56 
<< m1 >>
rect 126 55 127 56 
<< m2 >>
rect 126 55 127 56 
<< m2c >>
rect 126 55 127 56 
<< m1 >>
rect 126 55 127 56 
<< m2 >>
rect 126 55 127 56 
<< m1 >>
rect 127 55 128 56 
<< m1 >>
rect 128 55 129 56 
<< m1 >>
rect 129 55 130 56 
<< m1 >>
rect 130 55 131 56 
<< m1 >>
rect 131 55 132 56 
<< m1 >>
rect 132 55 133 56 
<< m1 >>
rect 134 55 135 56 
<< m1 >>
rect 136 55 137 56 
<< m2 >>
rect 136 55 137 56 
<< m1 >>
rect 137 55 138 56 
<< m1 >>
rect 138 55 139 56 
<< m1 >>
rect 139 55 140 56 
<< m1 >>
rect 148 55 149 56 
<< m1 >>
rect 150 55 151 56 
<< m1 >>
rect 154 55 155 56 
<< m1 >>
rect 163 55 164 56 
<< m1 >>
rect 165 55 166 56 
<< m1 >>
rect 172 55 173 56 
<< m1 >>
rect 181 55 182 56 
<< m1 >>
rect 183 55 184 56 
<< m1 >>
rect 186 55 187 56 
<< m1 >>
rect 190 55 191 56 
<< m2 >>
rect 190 55 191 56 
<< m1 >>
rect 196 55 197 56 
<< m1 >>
rect 197 55 198 56 
<< m2 >>
rect 197 55 198 56 
<< m2c >>
rect 197 55 198 56 
<< m1 >>
rect 197 55 198 56 
<< m2 >>
rect 197 55 198 56 
<< m2 >>
rect 198 55 199 56 
<< m1 >>
rect 199 55 200 56 
<< m2 >>
rect 199 55 200 56 
<< m2 >>
rect 200 55 201 56 
<< m1 >>
rect 202 55 203 56 
<< m1 >>
rect 204 55 205 56 
<< m1 >>
rect 232 55 233 56 
<< m1 >>
rect 233 55 234 56 
<< m1 >>
rect 234 55 235 56 
<< m1 >>
rect 235 55 236 56 
<< m1 >>
rect 243 55 244 56 
<< m1 >>
rect 250 55 251 56 
<< m1 >>
rect 254 55 255 56 
<< m1 >>
rect 256 55 257 56 
<< m1 >>
rect 26 56 27 57 
<< m1 >>
rect 28 56 29 57 
<< m2 >>
rect 28 56 29 57 
<< m1 >>
rect 37 56 38 57 
<< m1 >>
rect 40 56 41 57 
<< m2 >>
rect 43 56 44 57 
<< m1 >>
rect 44 56 45 57 
<< m1 >>
rect 46 56 47 57 
<< m1 >>
rect 49 56 50 57 
<< m1 >>
rect 50 56 51 57 
<< m1 >>
rect 51 56 52 57 
<< m1 >>
rect 52 56 53 57 
<< m1 >>
rect 53 56 54 57 
<< m1 >>
rect 54 56 55 57 
<< m1 >>
rect 55 56 56 57 
<< m1 >>
rect 56 56 57 57 
<< m1 >>
rect 57 56 58 57 
<< m1 >>
rect 58 56 59 57 
<< m1 >>
rect 60 56 61 57 
<< m2 >>
rect 60 56 61 57 
<< m2c >>
rect 60 56 61 57 
<< m1 >>
rect 60 56 61 57 
<< m2 >>
rect 60 56 61 57 
<< m1 >>
rect 71 56 72 57 
<< m1 >>
rect 73 56 74 57 
<< m1 >>
rect 75 56 76 57 
<< m1 >>
rect 82 56 83 57 
<< m1 >>
rect 106 56 107 57 
<< m1 >>
rect 109 56 110 57 
<< m1 >>
rect 113 56 114 57 
<< m1 >>
rect 118 56 119 57 
<< m1 >>
rect 121 56 122 57 
<< m1 >>
rect 122 56 123 57 
<< m2 >>
rect 122 56 123 57 
<< m2c >>
rect 122 56 123 57 
<< m1 >>
rect 122 56 123 57 
<< m2 >>
rect 122 56 123 57 
<< m2 >>
rect 123 56 124 57 
<< m1 >>
rect 124 56 125 57 
<< m2 >>
rect 124 56 125 57 
<< m2 >>
rect 125 56 126 57 
<< m1 >>
rect 134 56 135 57 
<< m2 >>
rect 136 56 137 57 
<< m1 >>
rect 148 56 149 57 
<< m1 >>
rect 150 56 151 57 
<< m1 >>
rect 154 56 155 57 
<< m1 >>
rect 163 56 164 57 
<< m1 >>
rect 165 56 166 57 
<< m1 >>
rect 172 56 173 57 
<< m1 >>
rect 181 56 182 57 
<< m2 >>
rect 181 56 182 57 
<< m2c >>
rect 181 56 182 57 
<< m1 >>
rect 181 56 182 57 
<< m2 >>
rect 181 56 182 57 
<< m1 >>
rect 183 56 184 57 
<< m2 >>
rect 183 56 184 57 
<< m2c >>
rect 183 56 184 57 
<< m1 >>
rect 183 56 184 57 
<< m2 >>
rect 183 56 184 57 
<< m1 >>
rect 186 56 187 57 
<< m2 >>
rect 186 56 187 57 
<< m2c >>
rect 186 56 187 57 
<< m1 >>
rect 186 56 187 57 
<< m2 >>
rect 186 56 187 57 
<< m1 >>
rect 190 56 191 57 
<< m2 >>
rect 190 56 191 57 
<< m1 >>
rect 199 56 200 57 
<< m2 >>
rect 200 56 201 57 
<< m1 >>
rect 202 56 203 57 
<< m1 >>
rect 204 56 205 57 
<< m1 >>
rect 243 56 244 57 
<< m2 >>
rect 243 56 244 57 
<< m2c >>
rect 243 56 244 57 
<< m1 >>
rect 243 56 244 57 
<< m2 >>
rect 243 56 244 57 
<< m1 >>
rect 250 56 251 57 
<< m1 >>
rect 254 56 255 57 
<< m2 >>
rect 254 56 255 57 
<< m2c >>
rect 254 56 255 57 
<< m1 >>
rect 254 56 255 57 
<< m2 >>
rect 254 56 255 57 
<< m1 >>
rect 256 56 257 57 
<< m1 >>
rect 26 57 27 58 
<< m1 >>
rect 28 57 29 58 
<< m2 >>
rect 28 57 29 58 
<< m1 >>
rect 37 57 38 58 
<< m1 >>
rect 40 57 41 58 
<< m2 >>
rect 43 57 44 58 
<< m1 >>
rect 44 57 45 58 
<< m1 >>
rect 46 57 47 58 
<< m2 >>
rect 60 57 61 58 
<< m1 >>
rect 71 57 72 58 
<< m1 >>
rect 73 57 74 58 
<< m1 >>
rect 75 57 76 58 
<< m2 >>
rect 76 57 77 58 
<< m1 >>
rect 77 57 78 58 
<< m2 >>
rect 77 57 78 58 
<< m2c >>
rect 77 57 78 58 
<< m1 >>
rect 77 57 78 58 
<< m2 >>
rect 77 57 78 58 
<< m1 >>
rect 78 57 79 58 
<< m1 >>
rect 79 57 80 58 
<< m1 >>
rect 80 57 81 58 
<< m1 >>
rect 81 57 82 58 
<< m1 >>
rect 82 57 83 58 
<< m1 >>
rect 106 57 107 58 
<< m1 >>
rect 109 57 110 58 
<< m1 >>
rect 113 57 114 58 
<< m2 >>
rect 113 57 114 58 
<< m2c >>
rect 113 57 114 58 
<< m1 >>
rect 113 57 114 58 
<< m2 >>
rect 113 57 114 58 
<< m1 >>
rect 118 57 119 58 
<< m1 >>
rect 119 57 120 58 
<< m2 >>
rect 119 57 120 58 
<< m2c >>
rect 119 57 120 58 
<< m1 >>
rect 119 57 120 58 
<< m2 >>
rect 119 57 120 58 
<< m2 >>
rect 120 57 121 58 
<< m1 >>
rect 124 57 125 58 
<< m1 >>
rect 134 57 135 58 
<< m1 >>
rect 136 57 137 58 
<< m2 >>
rect 136 57 137 58 
<< m2c >>
rect 136 57 137 58 
<< m1 >>
rect 136 57 137 58 
<< m2 >>
rect 136 57 137 58 
<< m1 >>
rect 148 57 149 58 
<< m1 >>
rect 150 57 151 58 
<< m1 >>
rect 154 57 155 58 
<< m1 >>
rect 163 57 164 58 
<< m1 >>
rect 165 57 166 58 
<< m1 >>
rect 172 57 173 58 
<< m2 >>
rect 181 57 182 58 
<< m2 >>
rect 183 57 184 58 
<< m2 >>
rect 186 57 187 58 
<< m1 >>
rect 190 57 191 58 
<< m2 >>
rect 190 57 191 58 
<< m1 >>
rect 199 57 200 58 
<< m2 >>
rect 200 57 201 58 
<< m1 >>
rect 202 57 203 58 
<< m1 >>
rect 204 57 205 58 
<< m2 >>
rect 243 57 244 58 
<< m1 >>
rect 250 57 251 58 
<< m2 >>
rect 254 57 255 58 
<< m1 >>
rect 256 57 257 58 
<< m1 >>
rect 26 58 27 59 
<< m1 >>
rect 28 58 29 59 
<< m2 >>
rect 28 58 29 59 
<< m1 >>
rect 37 58 38 59 
<< m1 >>
rect 40 58 41 59 
<< m2 >>
rect 43 58 44 59 
<< m1 >>
rect 44 58 45 59 
<< m1 >>
rect 46 58 47 59 
<< m1 >>
rect 49 58 50 59 
<< m1 >>
rect 50 58 51 59 
<< m1 >>
rect 51 58 52 59 
<< m1 >>
rect 52 58 53 59 
<< m1 >>
rect 53 58 54 59 
<< m1 >>
rect 54 58 55 59 
<< m1 >>
rect 55 58 56 59 
<< m1 >>
rect 56 58 57 59 
<< m1 >>
rect 57 58 58 59 
<< m1 >>
rect 58 58 59 59 
<< m1 >>
rect 59 58 60 59 
<< m1 >>
rect 60 58 61 59 
<< m2 >>
rect 60 58 61 59 
<< m1 >>
rect 61 58 62 59 
<< m1 >>
rect 62 58 63 59 
<< m1 >>
rect 63 58 64 59 
<< m1 >>
rect 64 58 65 59 
<< m2 >>
rect 64 58 65 59 
<< m2c >>
rect 64 58 65 59 
<< m1 >>
rect 64 58 65 59 
<< m2 >>
rect 64 58 65 59 
<< m2 >>
rect 65 58 66 59 
<< m1 >>
rect 66 58 67 59 
<< m2 >>
rect 66 58 67 59 
<< m1 >>
rect 67 58 68 59 
<< m2 >>
rect 67 58 68 59 
<< m1 >>
rect 68 58 69 59 
<< m2 >>
rect 68 58 69 59 
<< m1 >>
rect 69 58 70 59 
<< m2 >>
rect 69 58 70 59 
<< m1 >>
rect 70 58 71 59 
<< m2 >>
rect 70 58 71 59 
<< m1 >>
rect 71 58 72 59 
<< m2 >>
rect 71 58 72 59 
<< m2 >>
rect 72 58 73 59 
<< m1 >>
rect 73 58 74 59 
<< m2 >>
rect 73 58 74 59 
<< m2 >>
rect 74 58 75 59 
<< m1 >>
rect 75 58 76 59 
<< m2 >>
rect 75 58 76 59 
<< m2 >>
rect 76 58 77 59 
<< m1 >>
rect 106 58 107 59 
<< m1 >>
rect 109 58 110 59 
<< m2 >>
rect 113 58 114 59 
<< m2 >>
rect 120 58 121 59 
<< m1 >>
rect 124 58 125 59 
<< m1 >>
rect 134 58 135 59 
<< m1 >>
rect 136 58 137 59 
<< m1 >>
rect 148 58 149 59 
<< m1 >>
rect 150 58 151 59 
<< m1 >>
rect 154 58 155 59 
<< m1 >>
rect 163 58 164 59 
<< m1 >>
rect 165 58 166 59 
<< m1 >>
rect 172 58 173 59 
<< m2 >>
rect 173 58 174 59 
<< m1 >>
rect 174 58 175 59 
<< m2 >>
rect 174 58 175 59 
<< m2c >>
rect 174 58 175 59 
<< m1 >>
rect 174 58 175 59 
<< m2 >>
rect 174 58 175 59 
<< m1 >>
rect 175 58 176 59 
<< m1 >>
rect 176 58 177 59 
<< m1 >>
rect 177 58 178 59 
<< m1 >>
rect 178 58 179 59 
<< m1 >>
rect 179 58 180 59 
<< m1 >>
rect 180 58 181 59 
<< m1 >>
rect 181 58 182 59 
<< m2 >>
rect 181 58 182 59 
<< m1 >>
rect 182 58 183 59 
<< m1 >>
rect 183 58 184 59 
<< m2 >>
rect 183 58 184 59 
<< m1 >>
rect 184 58 185 59 
<< m1 >>
rect 185 58 186 59 
<< m1 >>
rect 186 58 187 59 
<< m2 >>
rect 186 58 187 59 
<< m1 >>
rect 187 58 188 59 
<< m1 >>
rect 188 58 189 59 
<< m1 >>
rect 189 58 190 59 
<< m1 >>
rect 190 58 191 59 
<< m2 >>
rect 190 58 191 59 
<< m1 >>
rect 199 58 200 59 
<< m2 >>
rect 200 58 201 59 
<< m1 >>
rect 202 58 203 59 
<< m1 >>
rect 204 58 205 59 
<< m2 >>
rect 243 58 244 59 
<< m1 >>
rect 244 58 245 59 
<< m2 >>
rect 244 58 245 59 
<< m1 >>
rect 245 58 246 59 
<< m2 >>
rect 245 58 246 59 
<< m1 >>
rect 246 58 247 59 
<< m2 >>
rect 246 58 247 59 
<< m1 >>
rect 247 58 248 59 
<< m2 >>
rect 247 58 248 59 
<< m1 >>
rect 248 58 249 59 
<< m2 >>
rect 248 58 249 59 
<< m1 >>
rect 249 58 250 59 
<< m2 >>
rect 249 58 250 59 
<< m1 >>
rect 250 58 251 59 
<< m2 >>
rect 250 58 251 59 
<< m2 >>
rect 251 58 252 59 
<< m1 >>
rect 252 58 253 59 
<< m2 >>
rect 252 58 253 59 
<< m2c >>
rect 252 58 253 59 
<< m1 >>
rect 252 58 253 59 
<< m2 >>
rect 252 58 253 59 
<< m1 >>
rect 253 58 254 59 
<< m2 >>
rect 254 58 255 59 
<< m1 >>
rect 256 58 257 59 
<< m1 >>
rect 26 59 27 60 
<< m1 >>
rect 28 59 29 60 
<< m2 >>
rect 28 59 29 60 
<< m1 >>
rect 37 59 38 60 
<< m1 >>
rect 40 59 41 60 
<< m2 >>
rect 43 59 44 60 
<< m1 >>
rect 44 59 45 60 
<< m1 >>
rect 46 59 47 60 
<< m1 >>
rect 49 59 50 60 
<< m2 >>
rect 60 59 61 60 
<< m1 >>
rect 66 59 67 60 
<< m1 >>
rect 73 59 74 60 
<< m1 >>
rect 75 59 76 60 
<< m1 >>
rect 77 59 78 60 
<< m2 >>
rect 77 59 78 60 
<< m2c >>
rect 77 59 78 60 
<< m1 >>
rect 77 59 78 60 
<< m2 >>
rect 77 59 78 60 
<< m1 >>
rect 78 59 79 60 
<< m1 >>
rect 79 59 80 60 
<< m1 >>
rect 80 59 81 60 
<< m1 >>
rect 81 59 82 60 
<< m1 >>
rect 82 59 83 60 
<< m1 >>
rect 83 59 84 60 
<< m1 >>
rect 84 59 85 60 
<< m1 >>
rect 85 59 86 60 
<< m1 >>
rect 86 59 87 60 
<< m1 >>
rect 87 59 88 60 
<< m1 >>
rect 88 59 89 60 
<< m1 >>
rect 89 59 90 60 
<< m1 >>
rect 90 59 91 60 
<< m1 >>
rect 91 59 92 60 
<< m1 >>
rect 92 59 93 60 
<< m1 >>
rect 93 59 94 60 
<< m1 >>
rect 94 59 95 60 
<< m1 >>
rect 95 59 96 60 
<< m1 >>
rect 96 59 97 60 
<< m1 >>
rect 97 59 98 60 
<< m1 >>
rect 98 59 99 60 
<< m1 >>
rect 99 59 100 60 
<< m1 >>
rect 100 59 101 60 
<< m1 >>
rect 101 59 102 60 
<< m1 >>
rect 102 59 103 60 
<< m1 >>
rect 103 59 104 60 
<< m1 >>
rect 104 59 105 60 
<< m2 >>
rect 104 59 105 60 
<< m2c >>
rect 104 59 105 60 
<< m1 >>
rect 104 59 105 60 
<< m2 >>
rect 104 59 105 60 
<< m2 >>
rect 105 59 106 60 
<< m1 >>
rect 106 59 107 60 
<< m2 >>
rect 106 59 107 60 
<< m2 >>
rect 107 59 108 60 
<< m2 >>
rect 108 59 109 60 
<< m1 >>
rect 109 59 110 60 
<< m2 >>
rect 109 59 110 60 
<< m2 >>
rect 110 59 111 60 
<< m1 >>
rect 111 59 112 60 
<< m2 >>
rect 111 59 112 60 
<< m2c >>
rect 111 59 112 60 
<< m1 >>
rect 111 59 112 60 
<< m2 >>
rect 111 59 112 60 
<< m1 >>
rect 112 59 113 60 
<< m1 >>
rect 113 59 114 60 
<< m2 >>
rect 113 59 114 60 
<< m1 >>
rect 114 59 115 60 
<< m1 >>
rect 115 59 116 60 
<< m1 >>
rect 116 59 117 60 
<< m1 >>
rect 117 59 118 60 
<< m1 >>
rect 118 59 119 60 
<< m1 >>
rect 119 59 120 60 
<< m1 >>
rect 120 59 121 60 
<< m2 >>
rect 120 59 121 60 
<< m1 >>
rect 121 59 122 60 
<< m1 >>
rect 122 59 123 60 
<< m1 >>
rect 123 59 124 60 
<< m1 >>
rect 124 59 125 60 
<< m1 >>
rect 134 59 135 60 
<< m1 >>
rect 136 59 137 60 
<< m2 >>
rect 136 59 137 60 
<< m2c >>
rect 136 59 137 60 
<< m1 >>
rect 136 59 137 60 
<< m2 >>
rect 136 59 137 60 
<< m1 >>
rect 148 59 149 60 
<< m2 >>
rect 148 59 149 60 
<< m2c >>
rect 148 59 149 60 
<< m1 >>
rect 148 59 149 60 
<< m2 >>
rect 148 59 149 60 
<< m1 >>
rect 150 59 151 60 
<< m2 >>
rect 150 59 151 60 
<< m2c >>
rect 150 59 151 60 
<< m1 >>
rect 150 59 151 60 
<< m2 >>
rect 150 59 151 60 
<< m1 >>
rect 154 59 155 60 
<< m1 >>
rect 163 59 164 60 
<< m2 >>
rect 163 59 164 60 
<< m2c >>
rect 163 59 164 60 
<< m1 >>
rect 163 59 164 60 
<< m2 >>
rect 163 59 164 60 
<< m1 >>
rect 165 59 166 60 
<< m2 >>
rect 165 59 166 60 
<< m2c >>
rect 165 59 166 60 
<< m1 >>
rect 165 59 166 60 
<< m2 >>
rect 165 59 166 60 
<< m1 >>
rect 172 59 173 60 
<< m2 >>
rect 173 59 174 60 
<< m2 >>
rect 181 59 182 60 
<< m2 >>
rect 183 59 184 60 
<< m2 >>
rect 186 59 187 60 
<< m2 >>
rect 190 59 191 60 
<< m1 >>
rect 199 59 200 60 
<< m2 >>
rect 200 59 201 60 
<< m1 >>
rect 202 59 203 60 
<< m1 >>
rect 204 59 205 60 
<< m1 >>
rect 244 59 245 60 
<< m1 >>
rect 253 59 254 60 
<< m2 >>
rect 254 59 255 60 
<< m1 >>
rect 256 59 257 60 
<< m1 >>
rect 26 60 27 61 
<< m1 >>
rect 28 60 29 61 
<< m2 >>
rect 28 60 29 61 
<< m1 >>
rect 37 60 38 61 
<< m1 >>
rect 40 60 41 61 
<< m2 >>
rect 43 60 44 61 
<< m1 >>
rect 44 60 45 61 
<< m2 >>
rect 44 60 45 61 
<< m2 >>
rect 45 60 46 61 
<< m1 >>
rect 46 60 47 61 
<< m2 >>
rect 46 60 47 61 
<< m2 >>
rect 47 60 48 61 
<< m2 >>
rect 48 60 49 61 
<< m1 >>
rect 49 60 50 61 
<< m2 >>
rect 49 60 50 61 
<< m2 >>
rect 50 60 51 61 
<< m1 >>
rect 51 60 52 61 
<< m2 >>
rect 51 60 52 61 
<< m2c >>
rect 51 60 52 61 
<< m1 >>
rect 51 60 52 61 
<< m2 >>
rect 51 60 52 61 
<< m1 >>
rect 52 60 53 61 
<< m1 >>
rect 53 60 54 61 
<< m1 >>
rect 54 60 55 61 
<< m1 >>
rect 55 60 56 61 
<< m1 >>
rect 56 60 57 61 
<< m1 >>
rect 57 60 58 61 
<< m1 >>
rect 58 60 59 61 
<< m1 >>
rect 59 60 60 61 
<< m1 >>
rect 60 60 61 61 
<< m2 >>
rect 60 60 61 61 
<< m1 >>
rect 61 60 62 61 
<< m1 >>
rect 62 60 63 61 
<< m1 >>
rect 63 60 64 61 
<< m1 >>
rect 64 60 65 61 
<< m2 >>
rect 64 60 65 61 
<< m2c >>
rect 64 60 65 61 
<< m1 >>
rect 64 60 65 61 
<< m2 >>
rect 64 60 65 61 
<< m2 >>
rect 65 60 66 61 
<< m1 >>
rect 66 60 67 61 
<< m2 >>
rect 66 60 67 61 
<< m2 >>
rect 67 60 68 61 
<< m1 >>
rect 68 60 69 61 
<< m2 >>
rect 68 60 69 61 
<< m2c >>
rect 68 60 69 61 
<< m1 >>
rect 68 60 69 61 
<< m2 >>
rect 68 60 69 61 
<< m1 >>
rect 69 60 70 61 
<< m1 >>
rect 70 60 71 61 
<< m1 >>
rect 71 60 72 61 
<< m2 >>
rect 71 60 72 61 
<< m2c >>
rect 71 60 72 61 
<< m1 >>
rect 71 60 72 61 
<< m2 >>
rect 71 60 72 61 
<< m2 >>
rect 72 60 73 61 
<< m1 >>
rect 73 60 74 61 
<< m2 >>
rect 73 60 74 61 
<< m2 >>
rect 74 60 75 61 
<< m1 >>
rect 75 60 76 61 
<< m2 >>
rect 75 60 76 61 
<< m2 >>
rect 76 60 77 61 
<< m2 >>
rect 77 60 78 61 
<< m1 >>
rect 106 60 107 61 
<< m1 >>
rect 109 60 110 61 
<< m2 >>
rect 113 60 114 61 
<< m2 >>
rect 120 60 121 61 
<< m2 >>
rect 121 60 122 61 
<< m2 >>
rect 122 60 123 61 
<< m2 >>
rect 123 60 124 61 
<< m2 >>
rect 124 60 125 61 
<< m1 >>
rect 134 60 135 61 
<< m2 >>
rect 136 60 137 61 
<< m2 >>
rect 138 60 139 61 
<< m2 >>
rect 139 60 140 61 
<< m2 >>
rect 140 60 141 61 
<< m2 >>
rect 141 60 142 61 
<< m2 >>
rect 142 60 143 61 
<< m2 >>
rect 143 60 144 61 
<< m2 >>
rect 144 60 145 61 
<< m2 >>
rect 145 60 146 61 
<< m2 >>
rect 146 60 147 61 
<< m2 >>
rect 147 60 148 61 
<< m2 >>
rect 148 60 149 61 
<< m2 >>
rect 150 60 151 61 
<< m1 >>
rect 154 60 155 61 
<< m2 >>
rect 163 60 164 61 
<< m2 >>
rect 165 60 166 61 
<< m1 >>
rect 172 60 173 61 
<< m2 >>
rect 173 60 174 61 
<< m1 >>
rect 181 60 182 61 
<< m2 >>
rect 181 60 182 61 
<< m2c >>
rect 181 60 182 61 
<< m1 >>
rect 181 60 182 61 
<< m2 >>
rect 181 60 182 61 
<< m1 >>
rect 183 60 184 61 
<< m2 >>
rect 183 60 184 61 
<< m2c >>
rect 183 60 184 61 
<< m1 >>
rect 183 60 184 61 
<< m2 >>
rect 183 60 184 61 
<< m1 >>
rect 186 60 187 61 
<< m2 >>
rect 186 60 187 61 
<< m2c >>
rect 186 60 187 61 
<< m1 >>
rect 186 60 187 61 
<< m2 >>
rect 186 60 187 61 
<< m1 >>
rect 190 60 191 61 
<< m2 >>
rect 190 60 191 61 
<< m2c >>
rect 190 60 191 61 
<< m1 >>
rect 190 60 191 61 
<< m2 >>
rect 190 60 191 61 
<< m1 >>
rect 199 60 200 61 
<< m2 >>
rect 200 60 201 61 
<< m1 >>
rect 202 60 203 61 
<< m1 >>
rect 204 60 205 61 
<< m1 >>
rect 205 60 206 61 
<< m1 >>
rect 206 60 207 61 
<< m1 >>
rect 207 60 208 61 
<< m1 >>
rect 208 60 209 61 
<< m1 >>
rect 209 60 210 61 
<< m1 >>
rect 210 60 211 61 
<< m1 >>
rect 211 60 212 61 
<< m1 >>
rect 212 60 213 61 
<< m1 >>
rect 213 60 214 61 
<< m1 >>
rect 214 60 215 61 
<< m1 >>
rect 215 60 216 61 
<< m1 >>
rect 216 60 217 61 
<< m1 >>
rect 217 60 218 61 
<< m1 >>
rect 218 60 219 61 
<< m1 >>
rect 219 60 220 61 
<< m1 >>
rect 220 60 221 61 
<< m1 >>
rect 221 60 222 61 
<< m1 >>
rect 222 60 223 61 
<< m1 >>
rect 223 60 224 61 
<< m1 >>
rect 224 60 225 61 
<< m1 >>
rect 225 60 226 61 
<< m1 >>
rect 226 60 227 61 
<< m1 >>
rect 227 60 228 61 
<< m1 >>
rect 228 60 229 61 
<< m1 >>
rect 229 60 230 61 
<< m1 >>
rect 230 60 231 61 
<< m1 >>
rect 231 60 232 61 
<< m1 >>
rect 232 60 233 61 
<< m1 >>
rect 233 60 234 61 
<< m1 >>
rect 234 60 235 61 
<< m1 >>
rect 235 60 236 61 
<< m1 >>
rect 236 60 237 61 
<< m1 >>
rect 237 60 238 61 
<< m1 >>
rect 238 60 239 61 
<< m1 >>
rect 239 60 240 61 
<< m1 >>
rect 240 60 241 61 
<< m1 >>
rect 241 60 242 61 
<< m1 >>
rect 242 60 243 61 
<< m2 >>
rect 242 60 243 61 
<< m2c >>
rect 242 60 243 61 
<< m1 >>
rect 242 60 243 61 
<< m2 >>
rect 242 60 243 61 
<< m2 >>
rect 243 60 244 61 
<< m1 >>
rect 244 60 245 61 
<< m1 >>
rect 253 60 254 61 
<< m2 >>
rect 254 60 255 61 
<< m1 >>
rect 256 60 257 61 
<< m1 >>
rect 26 61 27 62 
<< m1 >>
rect 28 61 29 62 
<< m2 >>
rect 28 61 29 62 
<< m1 >>
rect 37 61 38 62 
<< m1 >>
rect 40 61 41 62 
<< m1 >>
rect 44 61 45 62 
<< m1 >>
rect 46 61 47 62 
<< m1 >>
rect 49 61 50 62 
<< m2 >>
rect 60 61 61 62 
<< m1 >>
rect 66 61 67 62 
<< m1 >>
rect 73 61 74 62 
<< m1 >>
rect 75 61 76 62 
<< m1 >>
rect 77 61 78 62 
<< m1 >>
rect 78 61 79 62 
<< m1 >>
rect 79 61 80 62 
<< m1 >>
rect 80 61 81 62 
<< m1 >>
rect 81 61 82 62 
<< m1 >>
rect 82 61 83 62 
<< m1 >>
rect 83 61 84 62 
<< m1 >>
rect 84 61 85 62 
<< m1 >>
rect 85 61 86 62 
<< m1 >>
rect 86 61 87 62 
<< m1 >>
rect 87 61 88 62 
<< m1 >>
rect 88 61 89 62 
<< m1 >>
rect 89 61 90 62 
<< m1 >>
rect 90 61 91 62 
<< m1 >>
rect 91 61 92 62 
<< m1 >>
rect 92 61 93 62 
<< m1 >>
rect 93 61 94 62 
<< m1 >>
rect 94 61 95 62 
<< m1 >>
rect 95 61 96 62 
<< m1 >>
rect 96 61 97 62 
<< m1 >>
rect 97 61 98 62 
<< m1 >>
rect 98 61 99 62 
<< m1 >>
rect 99 61 100 62 
<< m1 >>
rect 100 61 101 62 
<< m1 >>
rect 101 61 102 62 
<< m1 >>
rect 102 61 103 62 
<< m1 >>
rect 103 61 104 62 
<< m1 >>
rect 104 61 105 62 
<< m2 >>
rect 104 61 105 62 
<< m2c >>
rect 104 61 105 62 
<< m1 >>
rect 104 61 105 62 
<< m2 >>
rect 104 61 105 62 
<< m2 >>
rect 105 61 106 62 
<< m1 >>
rect 106 61 107 62 
<< m2 >>
rect 106 61 107 62 
<< m2 >>
rect 107 61 108 62 
<< m1 >>
rect 108 61 109 62 
<< m2 >>
rect 108 61 109 62 
<< m2c >>
rect 108 61 109 62 
<< m1 >>
rect 108 61 109 62 
<< m2 >>
rect 108 61 109 62 
<< m1 >>
rect 109 61 110 62 
<< m1 >>
rect 113 61 114 62 
<< m2 >>
rect 113 61 114 62 
<< m2c >>
rect 113 61 114 62 
<< m1 >>
rect 113 61 114 62 
<< m2 >>
rect 113 61 114 62 
<< m1 >>
rect 124 61 125 62 
<< m2 >>
rect 124 61 125 62 
<< m2c >>
rect 124 61 125 62 
<< m1 >>
rect 124 61 125 62 
<< m2 >>
rect 124 61 125 62 
<< m1 >>
rect 134 61 135 62 
<< m1 >>
rect 135 61 136 62 
<< m1 >>
rect 136 61 137 62 
<< m2 >>
rect 136 61 137 62 
<< m1 >>
rect 137 61 138 62 
<< m1 >>
rect 138 61 139 62 
<< m2 >>
rect 138 61 139 62 
<< m1 >>
rect 139 61 140 62 
<< m1 >>
rect 140 61 141 62 
<< m1 >>
rect 141 61 142 62 
<< m1 >>
rect 142 61 143 62 
<< m1 >>
rect 143 61 144 62 
<< m1 >>
rect 144 61 145 62 
<< m1 >>
rect 145 61 146 62 
<< m1 >>
rect 146 61 147 62 
<< m1 >>
rect 147 61 148 62 
<< m1 >>
rect 148 61 149 62 
<< m1 >>
rect 149 61 150 62 
<< m1 >>
rect 150 61 151 62 
<< m2 >>
rect 150 61 151 62 
<< m1 >>
rect 151 61 152 62 
<< m1 >>
rect 152 61 153 62 
<< m2 >>
rect 152 61 153 62 
<< m2c >>
rect 152 61 153 62 
<< m1 >>
rect 152 61 153 62 
<< m2 >>
rect 152 61 153 62 
<< m2 >>
rect 153 61 154 62 
<< m1 >>
rect 154 61 155 62 
<< m2 >>
rect 154 61 155 62 
<< m2 >>
rect 155 61 156 62 
<< m1 >>
rect 156 61 157 62 
<< m2 >>
rect 156 61 157 62 
<< m2c >>
rect 156 61 157 62 
<< m1 >>
rect 156 61 157 62 
<< m2 >>
rect 156 61 157 62 
<< m1 >>
rect 157 61 158 62 
<< m1 >>
rect 158 61 159 62 
<< m1 >>
rect 159 61 160 62 
<< m1 >>
rect 160 61 161 62 
<< m1 >>
rect 161 61 162 62 
<< m1 >>
rect 162 61 163 62 
<< m1 >>
rect 163 61 164 62 
<< m2 >>
rect 163 61 164 62 
<< m1 >>
rect 164 61 165 62 
<< m1 >>
rect 165 61 166 62 
<< m2 >>
rect 165 61 166 62 
<< m1 >>
rect 166 61 167 62 
<< m1 >>
rect 167 61 168 62 
<< m1 >>
rect 168 61 169 62 
<< m1 >>
rect 169 61 170 62 
<< m1 >>
rect 170 61 171 62 
<< m1 >>
rect 172 61 173 62 
<< m2 >>
rect 173 61 174 62 
<< m1 >>
rect 181 61 182 62 
<< m1 >>
rect 183 61 184 62 
<< m1 >>
rect 186 61 187 62 
<< m1 >>
rect 190 61 191 62 
<< m1 >>
rect 199 61 200 62 
<< m2 >>
rect 200 61 201 62 
<< m1 >>
rect 202 61 203 62 
<< m2 >>
rect 243 61 244 62 
<< m1 >>
rect 244 61 245 62 
<< m1 >>
rect 253 61 254 62 
<< m2 >>
rect 254 61 255 62 
<< m1 >>
rect 256 61 257 62 
<< m1 >>
rect 26 62 27 63 
<< m1 >>
rect 28 62 29 63 
<< m2 >>
rect 28 62 29 63 
<< m1 >>
rect 37 62 38 63 
<< m1 >>
rect 40 62 41 63 
<< m1 >>
rect 44 62 45 63 
<< m1 >>
rect 46 62 47 63 
<< m1 >>
rect 49 62 50 63 
<< m2 >>
rect 60 62 61 63 
<< m1 >>
rect 66 62 67 63 
<< m1 >>
rect 73 62 74 63 
<< m2 >>
rect 73 62 74 63 
<< m2c >>
rect 73 62 74 63 
<< m1 >>
rect 73 62 74 63 
<< m2 >>
rect 73 62 74 63 
<< m1 >>
rect 75 62 76 63 
<< m2 >>
rect 75 62 76 63 
<< m2c >>
rect 75 62 76 63 
<< m1 >>
rect 75 62 76 63 
<< m2 >>
rect 75 62 76 63 
<< m1 >>
rect 77 62 78 63 
<< m2 >>
rect 77 62 78 63 
<< m2c >>
rect 77 62 78 63 
<< m1 >>
rect 77 62 78 63 
<< m2 >>
rect 77 62 78 63 
<< m1 >>
rect 106 62 107 63 
<< m2 >>
rect 113 62 114 63 
<< m1 >>
rect 124 62 125 63 
<< m2 >>
rect 136 62 137 63 
<< m2 >>
rect 138 62 139 63 
<< m2 >>
rect 150 62 151 63 
<< m1 >>
rect 154 62 155 63 
<< m2 >>
rect 163 62 164 63 
<< m2 >>
rect 165 62 166 63 
<< m1 >>
rect 170 62 171 63 
<< m1 >>
rect 172 62 173 63 
<< m2 >>
rect 173 62 174 63 
<< m1 >>
rect 181 62 182 63 
<< m1 >>
rect 183 62 184 63 
<< m1 >>
rect 186 62 187 63 
<< m1 >>
rect 190 62 191 63 
<< m1 >>
rect 199 62 200 63 
<< m2 >>
rect 200 62 201 63 
<< m1 >>
rect 202 62 203 63 
<< m2 >>
rect 243 62 244 63 
<< m1 >>
rect 244 62 245 63 
<< m1 >>
rect 253 62 254 63 
<< m2 >>
rect 254 62 255 63 
<< m1 >>
rect 256 62 257 63 
<< m1 >>
rect 26 63 27 64 
<< m1 >>
rect 28 63 29 64 
<< m2 >>
rect 28 63 29 64 
<< m1 >>
rect 37 63 38 64 
<< m1 >>
rect 40 63 41 64 
<< m1 >>
rect 44 63 45 64 
<< m1 >>
rect 46 63 47 64 
<< m1 >>
rect 49 63 50 64 
<< m2 >>
rect 56 63 57 64 
<< m1 >>
rect 57 63 58 64 
<< m2 >>
rect 57 63 58 64 
<< m2c >>
rect 57 63 58 64 
<< m1 >>
rect 57 63 58 64 
<< m2 >>
rect 57 63 58 64 
<< m1 >>
rect 58 63 59 64 
<< m1 >>
rect 59 63 60 64 
<< m1 >>
rect 60 63 61 64 
<< m2 >>
rect 60 63 61 64 
<< m1 >>
rect 61 63 62 64 
<< m1 >>
rect 62 63 63 64 
<< m1 >>
rect 63 63 64 64 
<< m1 >>
rect 64 63 65 64 
<< m1 >>
rect 65 63 66 64 
<< m1 >>
rect 66 63 67 64 
<< m2 >>
rect 73 63 74 64 
<< m2 >>
rect 75 63 76 64 
<< m2 >>
rect 77 63 78 64 
<< m2 >>
rect 105 63 106 64 
<< m1 >>
rect 106 63 107 64 
<< m2 >>
rect 106 63 107 64 
<< m1 >>
rect 107 63 108 64 
<< m2 >>
rect 107 63 108 64 
<< m1 >>
rect 108 63 109 64 
<< m2 >>
rect 108 63 109 64 
<< m1 >>
rect 109 63 110 64 
<< m2 >>
rect 109 63 110 64 
<< m1 >>
rect 110 63 111 64 
<< m1 >>
rect 111 63 112 64 
<< m1 >>
rect 112 63 113 64 
<< m1 >>
rect 113 63 114 64 
<< m2 >>
rect 113 63 114 64 
<< m1 >>
rect 114 63 115 64 
<< m1 >>
rect 115 63 116 64 
<< m1 >>
rect 116 63 117 64 
<< m1 >>
rect 117 63 118 64 
<< m1 >>
rect 118 63 119 64 
<< m1 >>
rect 124 63 125 64 
<< m1 >>
rect 136 63 137 64 
<< m2 >>
rect 136 63 137 64 
<< m1 >>
rect 137 63 138 64 
<< m1 >>
rect 138 63 139 64 
<< m2 >>
rect 138 63 139 64 
<< m2c >>
rect 138 63 139 64 
<< m1 >>
rect 138 63 139 64 
<< m2 >>
rect 138 63 139 64 
<< m1 >>
rect 150 63 151 64 
<< m2 >>
rect 150 63 151 64 
<< m2c >>
rect 150 63 151 64 
<< m1 >>
rect 150 63 151 64 
<< m2 >>
rect 150 63 151 64 
<< m1 >>
rect 154 63 155 64 
<< m1 >>
rect 163 63 164 64 
<< m2 >>
rect 163 63 164 64 
<< m2c >>
rect 163 63 164 64 
<< m1 >>
rect 163 63 164 64 
<< m2 >>
rect 163 63 164 64 
<< m1 >>
rect 165 63 166 64 
<< m2 >>
rect 165 63 166 64 
<< m2c >>
rect 165 63 166 64 
<< m1 >>
rect 165 63 166 64 
<< m2 >>
rect 165 63 166 64 
<< m1 >>
rect 168 63 169 64 
<< m2 >>
rect 168 63 169 64 
<< m2c >>
rect 168 63 169 64 
<< m1 >>
rect 168 63 169 64 
<< m2 >>
rect 168 63 169 64 
<< m2 >>
rect 169 63 170 64 
<< m1 >>
rect 170 63 171 64 
<< m2 >>
rect 170 63 171 64 
<< m2 >>
rect 171 63 172 64 
<< m1 >>
rect 172 63 173 64 
<< m2 >>
rect 172 63 173 64 
<< m2 >>
rect 173 63 174 64 
<< m1 >>
rect 175 63 176 64 
<< m1 >>
rect 176 63 177 64 
<< m1 >>
rect 177 63 178 64 
<< m1 >>
rect 178 63 179 64 
<< m1 >>
rect 179 63 180 64 
<< m2 >>
rect 179 63 180 64 
<< m2c >>
rect 179 63 180 64 
<< m1 >>
rect 179 63 180 64 
<< m2 >>
rect 179 63 180 64 
<< m2 >>
rect 180 63 181 64 
<< m1 >>
rect 181 63 182 64 
<< m2 >>
rect 181 63 182 64 
<< m2 >>
rect 182 63 183 64 
<< m1 >>
rect 183 63 184 64 
<< m2 >>
rect 183 63 184 64 
<< m2c >>
rect 183 63 184 64 
<< m1 >>
rect 183 63 184 64 
<< m2 >>
rect 183 63 184 64 
<< m1 >>
rect 186 63 187 64 
<< m1 >>
rect 190 63 191 64 
<< m1 >>
rect 199 63 200 64 
<< m2 >>
rect 200 63 201 64 
<< m1 >>
rect 202 63 203 64 
<< m2 >>
rect 243 63 244 64 
<< m1 >>
rect 244 63 245 64 
<< m1 >>
rect 253 63 254 64 
<< m2 >>
rect 254 63 255 64 
<< m1 >>
rect 256 63 257 64 
<< m1 >>
rect 26 64 27 65 
<< m1 >>
rect 28 64 29 65 
<< m2 >>
rect 28 64 29 65 
<< m1 >>
rect 37 64 38 65 
<< m1 >>
rect 40 64 41 65 
<< m1 >>
rect 44 64 45 65 
<< m1 >>
rect 46 64 47 65 
<< m1 >>
rect 49 64 50 65 
<< m1 >>
rect 52 64 53 65 
<< m1 >>
rect 53 64 54 65 
<< m1 >>
rect 54 64 55 65 
<< m1 >>
rect 55 64 56 65 
<< m2 >>
rect 56 64 57 65 
<< m2 >>
rect 60 64 61 65 
<< m1 >>
rect 70 64 71 65 
<< m1 >>
rect 71 64 72 65 
<< m1 >>
rect 72 64 73 65 
<< m1 >>
rect 73 64 74 65 
<< m2 >>
rect 73 64 74 65 
<< m1 >>
rect 74 64 75 65 
<< m1 >>
rect 75 64 76 65 
<< m2 >>
rect 75 64 76 65 
<< m1 >>
rect 76 64 77 65 
<< m1 >>
rect 77 64 78 65 
<< m2 >>
rect 77 64 78 65 
<< m1 >>
rect 78 64 79 65 
<< m1 >>
rect 79 64 80 65 
<< m1 >>
rect 80 64 81 65 
<< m1 >>
rect 81 64 82 65 
<< m1 >>
rect 82 64 83 65 
<< m1 >>
rect 103 64 104 65 
<< m1 >>
rect 104 64 105 65 
<< m2 >>
rect 104 64 105 65 
<< m2c >>
rect 104 64 105 65 
<< m1 >>
rect 104 64 105 65 
<< m2 >>
rect 104 64 105 65 
<< m2 >>
rect 105 64 106 65 
<< m2 >>
rect 109 64 110 65 
<< m2 >>
rect 113 64 114 65 
<< m1 >>
rect 118 64 119 65 
<< m1 >>
rect 124 64 125 65 
<< m1 >>
rect 136 64 137 65 
<< m2 >>
rect 136 64 137 65 
<< m1 >>
rect 150 64 151 65 
<< m1 >>
rect 151 64 152 65 
<< m1 >>
rect 152 64 153 65 
<< m2 >>
rect 152 64 153 65 
<< m2c >>
rect 152 64 153 65 
<< m1 >>
rect 152 64 153 65 
<< m2 >>
rect 152 64 153 65 
<< m2 >>
rect 153 64 154 65 
<< m1 >>
rect 154 64 155 65 
<< m2 >>
rect 154 64 155 65 
<< m2 >>
rect 155 64 156 65 
<< m1 >>
rect 156 64 157 65 
<< m2 >>
rect 156 64 157 65 
<< m2c >>
rect 156 64 157 65 
<< m1 >>
rect 156 64 157 65 
<< m2 >>
rect 156 64 157 65 
<< m1 >>
rect 157 64 158 65 
<< m1 >>
rect 163 64 164 65 
<< m1 >>
rect 165 64 166 65 
<< m1 >>
rect 168 64 169 65 
<< m1 >>
rect 170 64 171 65 
<< m1 >>
rect 172 64 173 65 
<< m1 >>
rect 175 64 176 65 
<< m1 >>
rect 181 64 182 65 
<< m1 >>
rect 186 64 187 65 
<< m1 >>
rect 190 64 191 65 
<< m1 >>
rect 199 64 200 65 
<< m2 >>
rect 200 64 201 65 
<< m1 >>
rect 202 64 203 65 
<< m2 >>
rect 243 64 244 65 
<< m1 >>
rect 244 64 245 65 
<< m1 >>
rect 253 64 254 65 
<< m2 >>
rect 254 64 255 65 
<< m1 >>
rect 256 64 257 65 
<< m1 >>
rect 26 65 27 66 
<< m1 >>
rect 28 65 29 66 
<< m2 >>
rect 28 65 29 66 
<< m1 >>
rect 37 65 38 66 
<< m1 >>
rect 40 65 41 66 
<< m1 >>
rect 44 65 45 66 
<< m1 >>
rect 46 65 47 66 
<< m1 >>
rect 49 65 50 66 
<< m1 >>
rect 52 65 53 66 
<< m1 >>
rect 55 65 56 66 
<< m2 >>
rect 56 65 57 66 
<< m1 >>
rect 60 65 61 66 
<< m2 >>
rect 60 65 61 66 
<< m2c >>
rect 60 65 61 66 
<< m1 >>
rect 60 65 61 66 
<< m2 >>
rect 60 65 61 66 
<< m1 >>
rect 70 65 71 66 
<< m2 >>
rect 73 65 74 66 
<< m2 >>
rect 75 65 76 66 
<< m2 >>
rect 77 65 78 66 
<< m1 >>
rect 82 65 83 66 
<< m1 >>
rect 103 65 104 66 
<< m1 >>
rect 109 65 110 66 
<< m2 >>
rect 109 65 110 66 
<< m2c >>
rect 109 65 110 66 
<< m1 >>
rect 109 65 110 66 
<< m2 >>
rect 109 65 110 66 
<< m1 >>
rect 113 65 114 66 
<< m2 >>
rect 113 65 114 66 
<< m2c >>
rect 113 65 114 66 
<< m1 >>
rect 113 65 114 66 
<< m2 >>
rect 113 65 114 66 
<< m1 >>
rect 118 65 119 66 
<< m1 >>
rect 124 65 125 66 
<< m1 >>
rect 136 65 137 66 
<< m2 >>
rect 136 65 137 66 
<< m1 >>
rect 154 65 155 66 
<< m1 >>
rect 157 65 158 66 
<< m1 >>
rect 163 65 164 66 
<< m1 >>
rect 165 65 166 66 
<< m2 >>
rect 166 65 167 66 
<< m1 >>
rect 167 65 168 66 
<< m2 >>
rect 167 65 168 66 
<< m2c >>
rect 167 65 168 66 
<< m1 >>
rect 167 65 168 66 
<< m2 >>
rect 167 65 168 66 
<< m1 >>
rect 168 65 169 66 
<< m1 >>
rect 170 65 171 66 
<< m1 >>
rect 172 65 173 66 
<< m1 >>
rect 175 65 176 66 
<< m1 >>
rect 181 65 182 66 
<< m1 >>
rect 186 65 187 66 
<< m1 >>
rect 190 65 191 66 
<< m1 >>
rect 199 65 200 66 
<< m2 >>
rect 200 65 201 66 
<< m1 >>
rect 202 65 203 66 
<< m2 >>
rect 243 65 244 66 
<< m1 >>
rect 244 65 245 66 
<< m1 >>
rect 253 65 254 66 
<< m2 >>
rect 254 65 255 66 
<< m1 >>
rect 256 65 257 66 
<< pdiffusion >>
rect 12 66 13 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< m1 >>
rect 26 66 27 67 
<< m1 >>
rect 28 66 29 67 
<< m2 >>
rect 28 66 29 67 
<< pdiffusion >>
rect 30 66 31 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< m1 >>
rect 37 66 38 67 
<< m1 >>
rect 40 66 41 67 
<< m1 >>
rect 44 66 45 67 
<< m1 >>
rect 46 66 47 67 
<< pdiffusion >>
rect 48 66 49 67 
<< m1 >>
rect 49 66 50 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< m1 >>
rect 52 66 53 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 55 66 56 67 
<< m2 >>
rect 56 66 57 67 
<< m1 >>
rect 60 66 61 67 
<< pdiffusion >>
rect 66 66 67 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< m1 >>
rect 70 66 71 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< m1 >>
rect 73 66 74 67 
<< m2 >>
rect 73 66 74 67 
<< m2c >>
rect 73 66 74 67 
<< m1 >>
rect 73 66 74 67 
<< m2 >>
rect 73 66 74 67 
<< m1 >>
rect 75 66 76 67 
<< m2 >>
rect 75 66 76 67 
<< m2c >>
rect 75 66 76 67 
<< m1 >>
rect 75 66 76 67 
<< m2 >>
rect 75 66 76 67 
<< m1 >>
rect 77 66 78 67 
<< m2 >>
rect 77 66 78 67 
<< m2c >>
rect 77 66 78 67 
<< m1 >>
rect 77 66 78 67 
<< m2 >>
rect 77 66 78 67 
<< m1 >>
rect 82 66 83 67 
<< pdiffusion >>
rect 84 66 85 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< pdiffusion >>
rect 102 66 103 67 
<< m1 >>
rect 103 66 104 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< m1 >>
rect 109 66 110 67 
<< m1 >>
rect 113 66 114 67 
<< m1 >>
rect 118 66 119 67 
<< pdiffusion >>
rect 120 66 121 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< m1 >>
rect 124 66 125 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< m1 >>
rect 136 66 137 67 
<< m2 >>
rect 136 66 137 67 
<< pdiffusion >>
rect 138 66 139 67 
<< pdiffusion >>
rect 139 66 140 67 
<< pdiffusion >>
rect 140 66 141 67 
<< pdiffusion >>
rect 141 66 142 67 
<< pdiffusion >>
rect 142 66 143 67 
<< pdiffusion >>
rect 143 66 144 67 
<< m1 >>
rect 154 66 155 67 
<< pdiffusion >>
rect 156 66 157 67 
<< m1 >>
rect 157 66 158 67 
<< pdiffusion >>
rect 157 66 158 67 
<< pdiffusion >>
rect 158 66 159 67 
<< pdiffusion >>
rect 159 66 160 67 
<< pdiffusion >>
rect 160 66 161 67 
<< pdiffusion >>
rect 161 66 162 67 
<< m1 >>
rect 163 66 164 67 
<< m1 >>
rect 165 66 166 67 
<< m2 >>
rect 166 66 167 67 
<< m1 >>
rect 170 66 171 67 
<< m1 >>
rect 172 66 173 67 
<< pdiffusion >>
rect 174 66 175 67 
<< m1 >>
rect 175 66 176 67 
<< pdiffusion >>
rect 175 66 176 67 
<< pdiffusion >>
rect 176 66 177 67 
<< pdiffusion >>
rect 177 66 178 67 
<< pdiffusion >>
rect 178 66 179 67 
<< pdiffusion >>
rect 179 66 180 67 
<< m1 >>
rect 181 66 182 67 
<< m1 >>
rect 186 66 187 67 
<< m1 >>
rect 190 66 191 67 
<< pdiffusion >>
rect 192 66 193 67 
<< pdiffusion >>
rect 193 66 194 67 
<< pdiffusion >>
rect 194 66 195 67 
<< pdiffusion >>
rect 195 66 196 67 
<< pdiffusion >>
rect 196 66 197 67 
<< pdiffusion >>
rect 197 66 198 67 
<< m1 >>
rect 199 66 200 67 
<< m2 >>
rect 200 66 201 67 
<< m1 >>
rect 202 66 203 67 
<< pdiffusion >>
rect 210 66 211 67 
<< pdiffusion >>
rect 211 66 212 67 
<< pdiffusion >>
rect 212 66 213 67 
<< pdiffusion >>
rect 213 66 214 67 
<< pdiffusion >>
rect 214 66 215 67 
<< pdiffusion >>
rect 215 66 216 67 
<< pdiffusion >>
rect 228 66 229 67 
<< pdiffusion >>
rect 229 66 230 67 
<< pdiffusion >>
rect 230 66 231 67 
<< pdiffusion >>
rect 231 66 232 67 
<< pdiffusion >>
rect 232 66 233 67 
<< pdiffusion >>
rect 233 66 234 67 
<< m2 >>
rect 243 66 244 67 
<< m1 >>
rect 244 66 245 67 
<< pdiffusion >>
rect 246 66 247 67 
<< pdiffusion >>
rect 247 66 248 67 
<< pdiffusion >>
rect 248 66 249 67 
<< pdiffusion >>
rect 249 66 250 67 
<< pdiffusion >>
rect 250 66 251 67 
<< pdiffusion >>
rect 251 66 252 67 
<< m1 >>
rect 253 66 254 67 
<< m2 >>
rect 254 66 255 67 
<< m1 >>
rect 256 66 257 67 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< m1 >>
rect 26 67 27 68 
<< m1 >>
rect 28 67 29 68 
<< m2 >>
rect 28 67 29 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< m1 >>
rect 37 67 38 68 
<< m1 >>
rect 40 67 41 68 
<< m1 >>
rect 44 67 45 68 
<< m1 >>
rect 46 67 47 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 55 67 56 68 
<< m2 >>
rect 56 67 57 68 
<< m1 >>
rect 60 67 61 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< m1 >>
rect 73 67 74 68 
<< m1 >>
rect 75 67 76 68 
<< m1 >>
rect 77 67 78 68 
<< m1 >>
rect 82 67 83 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< m1 >>
rect 109 67 110 68 
<< m2 >>
rect 110 67 111 68 
<< m1 >>
rect 111 67 112 68 
<< m2 >>
rect 111 67 112 68 
<< m2c >>
rect 111 67 112 68 
<< m1 >>
rect 111 67 112 68 
<< m2 >>
rect 111 67 112 68 
<< m1 >>
rect 112 67 113 68 
<< m1 >>
rect 113 67 114 68 
<< m1 >>
rect 118 67 119 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< m1 >>
rect 136 67 137 68 
<< m2 >>
rect 136 67 137 68 
<< pdiffusion >>
rect 138 67 139 68 
<< pdiffusion >>
rect 139 67 140 68 
<< pdiffusion >>
rect 140 67 141 68 
<< pdiffusion >>
rect 141 67 142 68 
<< pdiffusion >>
rect 142 67 143 68 
<< pdiffusion >>
rect 143 67 144 68 
<< m1 >>
rect 154 67 155 68 
<< pdiffusion >>
rect 156 67 157 68 
<< pdiffusion >>
rect 157 67 158 68 
<< pdiffusion >>
rect 158 67 159 68 
<< pdiffusion >>
rect 159 67 160 68 
<< pdiffusion >>
rect 160 67 161 68 
<< pdiffusion >>
rect 161 67 162 68 
<< m1 >>
rect 163 67 164 68 
<< m1 >>
rect 165 67 166 68 
<< m2 >>
rect 166 67 167 68 
<< m1 >>
rect 170 67 171 68 
<< m1 >>
rect 172 67 173 68 
<< pdiffusion >>
rect 174 67 175 68 
<< pdiffusion >>
rect 175 67 176 68 
<< pdiffusion >>
rect 176 67 177 68 
<< pdiffusion >>
rect 177 67 178 68 
<< pdiffusion >>
rect 178 67 179 68 
<< pdiffusion >>
rect 179 67 180 68 
<< m1 >>
rect 181 67 182 68 
<< m1 >>
rect 186 67 187 68 
<< m1 >>
rect 190 67 191 68 
<< pdiffusion >>
rect 192 67 193 68 
<< pdiffusion >>
rect 193 67 194 68 
<< pdiffusion >>
rect 194 67 195 68 
<< pdiffusion >>
rect 195 67 196 68 
<< pdiffusion >>
rect 196 67 197 68 
<< pdiffusion >>
rect 197 67 198 68 
<< m1 >>
rect 199 67 200 68 
<< m2 >>
rect 200 67 201 68 
<< m1 >>
rect 202 67 203 68 
<< pdiffusion >>
rect 210 67 211 68 
<< pdiffusion >>
rect 211 67 212 68 
<< pdiffusion >>
rect 212 67 213 68 
<< pdiffusion >>
rect 213 67 214 68 
<< pdiffusion >>
rect 214 67 215 68 
<< pdiffusion >>
rect 215 67 216 68 
<< pdiffusion >>
rect 228 67 229 68 
<< pdiffusion >>
rect 229 67 230 68 
<< pdiffusion >>
rect 230 67 231 68 
<< pdiffusion >>
rect 231 67 232 68 
<< pdiffusion >>
rect 232 67 233 68 
<< pdiffusion >>
rect 233 67 234 68 
<< m2 >>
rect 243 67 244 68 
<< m1 >>
rect 244 67 245 68 
<< pdiffusion >>
rect 246 67 247 68 
<< pdiffusion >>
rect 247 67 248 68 
<< pdiffusion >>
rect 248 67 249 68 
<< pdiffusion >>
rect 249 67 250 68 
<< pdiffusion >>
rect 250 67 251 68 
<< pdiffusion >>
rect 251 67 252 68 
<< m1 >>
rect 253 67 254 68 
<< m2 >>
rect 254 67 255 68 
<< m1 >>
rect 256 67 257 68 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< m1 >>
rect 26 68 27 69 
<< m1 >>
rect 28 68 29 69 
<< m2 >>
rect 28 68 29 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< m1 >>
rect 37 68 38 69 
<< m1 >>
rect 40 68 41 69 
<< m1 >>
rect 44 68 45 69 
<< m1 >>
rect 46 68 47 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 55 68 56 69 
<< m2 >>
rect 56 68 57 69 
<< m1 >>
rect 60 68 61 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< m1 >>
rect 73 68 74 69 
<< m1 >>
rect 75 68 76 69 
<< m1 >>
rect 77 68 78 69 
<< m1 >>
rect 82 68 83 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< m1 >>
rect 109 68 110 69 
<< m2 >>
rect 110 68 111 69 
<< m1 >>
rect 118 68 119 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< m1 >>
rect 136 68 137 69 
<< m2 >>
rect 136 68 137 69 
<< pdiffusion >>
rect 138 68 139 69 
<< pdiffusion >>
rect 139 68 140 69 
<< pdiffusion >>
rect 140 68 141 69 
<< pdiffusion >>
rect 141 68 142 69 
<< pdiffusion >>
rect 142 68 143 69 
<< pdiffusion >>
rect 143 68 144 69 
<< m1 >>
rect 154 68 155 69 
<< pdiffusion >>
rect 156 68 157 69 
<< pdiffusion >>
rect 157 68 158 69 
<< pdiffusion >>
rect 158 68 159 69 
<< pdiffusion >>
rect 159 68 160 69 
<< pdiffusion >>
rect 160 68 161 69 
<< pdiffusion >>
rect 161 68 162 69 
<< m1 >>
rect 163 68 164 69 
<< m1 >>
rect 165 68 166 69 
<< m2 >>
rect 166 68 167 69 
<< m1 >>
rect 170 68 171 69 
<< m1 >>
rect 172 68 173 69 
<< pdiffusion >>
rect 174 68 175 69 
<< pdiffusion >>
rect 175 68 176 69 
<< pdiffusion >>
rect 176 68 177 69 
<< pdiffusion >>
rect 177 68 178 69 
<< pdiffusion >>
rect 178 68 179 69 
<< pdiffusion >>
rect 179 68 180 69 
<< m1 >>
rect 181 68 182 69 
<< m1 >>
rect 186 68 187 69 
<< m1 >>
rect 190 68 191 69 
<< pdiffusion >>
rect 192 68 193 69 
<< pdiffusion >>
rect 193 68 194 69 
<< pdiffusion >>
rect 194 68 195 69 
<< pdiffusion >>
rect 195 68 196 69 
<< pdiffusion >>
rect 196 68 197 69 
<< pdiffusion >>
rect 197 68 198 69 
<< m1 >>
rect 199 68 200 69 
<< m2 >>
rect 200 68 201 69 
<< m1 >>
rect 202 68 203 69 
<< pdiffusion >>
rect 210 68 211 69 
<< pdiffusion >>
rect 211 68 212 69 
<< pdiffusion >>
rect 212 68 213 69 
<< pdiffusion >>
rect 213 68 214 69 
<< pdiffusion >>
rect 214 68 215 69 
<< pdiffusion >>
rect 215 68 216 69 
<< pdiffusion >>
rect 228 68 229 69 
<< pdiffusion >>
rect 229 68 230 69 
<< pdiffusion >>
rect 230 68 231 69 
<< pdiffusion >>
rect 231 68 232 69 
<< pdiffusion >>
rect 232 68 233 69 
<< pdiffusion >>
rect 233 68 234 69 
<< m2 >>
rect 243 68 244 69 
<< m1 >>
rect 244 68 245 69 
<< pdiffusion >>
rect 246 68 247 69 
<< pdiffusion >>
rect 247 68 248 69 
<< pdiffusion >>
rect 248 68 249 69 
<< pdiffusion >>
rect 249 68 250 69 
<< pdiffusion >>
rect 250 68 251 69 
<< pdiffusion >>
rect 251 68 252 69 
<< m1 >>
rect 253 68 254 69 
<< m2 >>
rect 254 68 255 69 
<< m1 >>
rect 256 68 257 69 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< m1 >>
rect 26 69 27 70 
<< m1 >>
rect 28 69 29 70 
<< m2 >>
rect 28 69 29 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< m1 >>
rect 37 69 38 70 
<< m1 >>
rect 40 69 41 70 
<< m1 >>
rect 44 69 45 70 
<< m1 >>
rect 46 69 47 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 55 69 56 70 
<< m2 >>
rect 56 69 57 70 
<< m1 >>
rect 60 69 61 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< m1 >>
rect 73 69 74 70 
<< m1 >>
rect 75 69 76 70 
<< m1 >>
rect 77 69 78 70 
<< m1 >>
rect 82 69 83 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< m1 >>
rect 109 69 110 70 
<< m2 >>
rect 110 69 111 70 
<< m1 >>
rect 118 69 119 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< m1 >>
rect 136 69 137 70 
<< m2 >>
rect 136 69 137 70 
<< pdiffusion >>
rect 138 69 139 70 
<< pdiffusion >>
rect 139 69 140 70 
<< pdiffusion >>
rect 140 69 141 70 
<< pdiffusion >>
rect 141 69 142 70 
<< pdiffusion >>
rect 142 69 143 70 
<< pdiffusion >>
rect 143 69 144 70 
<< m1 >>
rect 154 69 155 70 
<< pdiffusion >>
rect 156 69 157 70 
<< pdiffusion >>
rect 157 69 158 70 
<< pdiffusion >>
rect 158 69 159 70 
<< pdiffusion >>
rect 159 69 160 70 
<< pdiffusion >>
rect 160 69 161 70 
<< pdiffusion >>
rect 161 69 162 70 
<< m1 >>
rect 163 69 164 70 
<< m1 >>
rect 165 69 166 70 
<< m2 >>
rect 166 69 167 70 
<< m1 >>
rect 170 69 171 70 
<< m1 >>
rect 172 69 173 70 
<< pdiffusion >>
rect 174 69 175 70 
<< pdiffusion >>
rect 175 69 176 70 
<< pdiffusion >>
rect 176 69 177 70 
<< pdiffusion >>
rect 177 69 178 70 
<< pdiffusion >>
rect 178 69 179 70 
<< pdiffusion >>
rect 179 69 180 70 
<< m1 >>
rect 181 69 182 70 
<< m1 >>
rect 186 69 187 70 
<< m1 >>
rect 190 69 191 70 
<< pdiffusion >>
rect 192 69 193 70 
<< pdiffusion >>
rect 193 69 194 70 
<< pdiffusion >>
rect 194 69 195 70 
<< pdiffusion >>
rect 195 69 196 70 
<< pdiffusion >>
rect 196 69 197 70 
<< pdiffusion >>
rect 197 69 198 70 
<< m1 >>
rect 199 69 200 70 
<< m2 >>
rect 200 69 201 70 
<< m1 >>
rect 202 69 203 70 
<< pdiffusion >>
rect 210 69 211 70 
<< pdiffusion >>
rect 211 69 212 70 
<< pdiffusion >>
rect 212 69 213 70 
<< pdiffusion >>
rect 213 69 214 70 
<< pdiffusion >>
rect 214 69 215 70 
<< pdiffusion >>
rect 215 69 216 70 
<< pdiffusion >>
rect 228 69 229 70 
<< pdiffusion >>
rect 229 69 230 70 
<< pdiffusion >>
rect 230 69 231 70 
<< pdiffusion >>
rect 231 69 232 70 
<< pdiffusion >>
rect 232 69 233 70 
<< pdiffusion >>
rect 233 69 234 70 
<< m2 >>
rect 243 69 244 70 
<< m1 >>
rect 244 69 245 70 
<< pdiffusion >>
rect 246 69 247 70 
<< pdiffusion >>
rect 247 69 248 70 
<< pdiffusion >>
rect 248 69 249 70 
<< pdiffusion >>
rect 249 69 250 70 
<< pdiffusion >>
rect 250 69 251 70 
<< pdiffusion >>
rect 251 69 252 70 
<< m1 >>
rect 253 69 254 70 
<< m2 >>
rect 254 69 255 70 
<< m1 >>
rect 256 69 257 70 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< m1 >>
rect 26 70 27 71 
<< m1 >>
rect 28 70 29 71 
<< m2 >>
rect 28 70 29 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< m1 >>
rect 37 70 38 71 
<< m1 >>
rect 40 70 41 71 
<< m1 >>
rect 44 70 45 71 
<< m1 >>
rect 46 70 47 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 55 70 56 71 
<< m2 >>
rect 56 70 57 71 
<< m1 >>
rect 60 70 61 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< m1 >>
rect 73 70 74 71 
<< m1 >>
rect 75 70 76 71 
<< m1 >>
rect 77 70 78 71 
<< m1 >>
rect 82 70 83 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< m1 >>
rect 109 70 110 71 
<< m2 >>
rect 110 70 111 71 
<< m1 >>
rect 118 70 119 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< m1 >>
rect 136 70 137 71 
<< m2 >>
rect 136 70 137 71 
<< pdiffusion >>
rect 138 70 139 71 
<< pdiffusion >>
rect 139 70 140 71 
<< pdiffusion >>
rect 140 70 141 71 
<< pdiffusion >>
rect 141 70 142 71 
<< pdiffusion >>
rect 142 70 143 71 
<< pdiffusion >>
rect 143 70 144 71 
<< m1 >>
rect 154 70 155 71 
<< pdiffusion >>
rect 156 70 157 71 
<< pdiffusion >>
rect 157 70 158 71 
<< pdiffusion >>
rect 158 70 159 71 
<< pdiffusion >>
rect 159 70 160 71 
<< pdiffusion >>
rect 160 70 161 71 
<< pdiffusion >>
rect 161 70 162 71 
<< m1 >>
rect 163 70 164 71 
<< m1 >>
rect 165 70 166 71 
<< m2 >>
rect 166 70 167 71 
<< m1 >>
rect 170 70 171 71 
<< m1 >>
rect 172 70 173 71 
<< pdiffusion >>
rect 174 70 175 71 
<< pdiffusion >>
rect 175 70 176 71 
<< pdiffusion >>
rect 176 70 177 71 
<< pdiffusion >>
rect 177 70 178 71 
<< pdiffusion >>
rect 178 70 179 71 
<< pdiffusion >>
rect 179 70 180 71 
<< m1 >>
rect 181 70 182 71 
<< m1 >>
rect 186 70 187 71 
<< m1 >>
rect 190 70 191 71 
<< pdiffusion >>
rect 192 70 193 71 
<< pdiffusion >>
rect 193 70 194 71 
<< pdiffusion >>
rect 194 70 195 71 
<< pdiffusion >>
rect 195 70 196 71 
<< pdiffusion >>
rect 196 70 197 71 
<< pdiffusion >>
rect 197 70 198 71 
<< m1 >>
rect 199 70 200 71 
<< m2 >>
rect 200 70 201 71 
<< m1 >>
rect 202 70 203 71 
<< pdiffusion >>
rect 210 70 211 71 
<< pdiffusion >>
rect 211 70 212 71 
<< pdiffusion >>
rect 212 70 213 71 
<< pdiffusion >>
rect 213 70 214 71 
<< pdiffusion >>
rect 214 70 215 71 
<< pdiffusion >>
rect 215 70 216 71 
<< pdiffusion >>
rect 228 70 229 71 
<< pdiffusion >>
rect 229 70 230 71 
<< pdiffusion >>
rect 230 70 231 71 
<< pdiffusion >>
rect 231 70 232 71 
<< pdiffusion >>
rect 232 70 233 71 
<< pdiffusion >>
rect 233 70 234 71 
<< m2 >>
rect 243 70 244 71 
<< m1 >>
rect 244 70 245 71 
<< pdiffusion >>
rect 246 70 247 71 
<< pdiffusion >>
rect 247 70 248 71 
<< pdiffusion >>
rect 248 70 249 71 
<< pdiffusion >>
rect 249 70 250 71 
<< pdiffusion >>
rect 250 70 251 71 
<< pdiffusion >>
rect 251 70 252 71 
<< m1 >>
rect 253 70 254 71 
<< m2 >>
rect 254 70 255 71 
<< m1 >>
rect 256 70 257 71 
<< pdiffusion >>
rect 12 71 13 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< m1 >>
rect 16 71 17 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< m1 >>
rect 26 71 27 72 
<< m2 >>
rect 26 71 27 72 
<< m2c >>
rect 26 71 27 72 
<< m1 >>
rect 26 71 27 72 
<< m2 >>
rect 26 71 27 72 
<< m1 >>
rect 28 71 29 72 
<< m2 >>
rect 28 71 29 72 
<< pdiffusion >>
rect 30 71 31 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< m1 >>
rect 37 71 38 72 
<< m1 >>
rect 40 71 41 72 
<< m1 >>
rect 44 71 45 72 
<< m1 >>
rect 46 71 47 72 
<< pdiffusion >>
rect 48 71 49 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< m1 >>
rect 52 71 53 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 55 71 56 72 
<< m2 >>
rect 56 71 57 72 
<< m1 >>
rect 60 71 61 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< m1 >>
rect 73 71 74 72 
<< m1 >>
rect 75 71 76 72 
<< m1 >>
rect 77 71 78 72 
<< m1 >>
rect 82 71 83 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< m1 >>
rect 88 71 89 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< pdiffusion >>
rect 102 71 103 72 
<< m1 >>
rect 103 71 104 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< m1 >>
rect 106 71 107 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< m1 >>
rect 109 71 110 72 
<< m2 >>
rect 110 71 111 72 
<< m1 >>
rect 118 71 119 72 
<< pdiffusion >>
rect 120 71 121 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< m1 >>
rect 124 71 125 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< m1 >>
rect 136 71 137 72 
<< m2 >>
rect 136 71 137 72 
<< pdiffusion >>
rect 138 71 139 72 
<< pdiffusion >>
rect 139 71 140 72 
<< pdiffusion >>
rect 140 71 141 72 
<< pdiffusion >>
rect 141 71 142 72 
<< m1 >>
rect 142 71 143 72 
<< pdiffusion >>
rect 142 71 143 72 
<< pdiffusion >>
rect 143 71 144 72 
<< m1 >>
rect 154 71 155 72 
<< pdiffusion >>
rect 156 71 157 72 
<< m1 >>
rect 157 71 158 72 
<< pdiffusion >>
rect 157 71 158 72 
<< pdiffusion >>
rect 158 71 159 72 
<< pdiffusion >>
rect 159 71 160 72 
<< pdiffusion >>
rect 160 71 161 72 
<< pdiffusion >>
rect 161 71 162 72 
<< m1 >>
rect 163 71 164 72 
<< m1 >>
rect 165 71 166 72 
<< m2 >>
rect 166 71 167 72 
<< m1 >>
rect 170 71 171 72 
<< m1 >>
rect 172 71 173 72 
<< pdiffusion >>
rect 174 71 175 72 
<< m1 >>
rect 175 71 176 72 
<< pdiffusion >>
rect 175 71 176 72 
<< pdiffusion >>
rect 176 71 177 72 
<< pdiffusion >>
rect 177 71 178 72 
<< pdiffusion >>
rect 178 71 179 72 
<< pdiffusion >>
rect 179 71 180 72 
<< m1 >>
rect 181 71 182 72 
<< m1 >>
rect 186 71 187 72 
<< m1 >>
rect 190 71 191 72 
<< pdiffusion >>
rect 192 71 193 72 
<< pdiffusion >>
rect 193 71 194 72 
<< pdiffusion >>
rect 194 71 195 72 
<< pdiffusion >>
rect 195 71 196 72 
<< pdiffusion >>
rect 196 71 197 72 
<< pdiffusion >>
rect 197 71 198 72 
<< m1 >>
rect 199 71 200 72 
<< m2 >>
rect 200 71 201 72 
<< m1 >>
rect 202 71 203 72 
<< pdiffusion >>
rect 210 71 211 72 
<< m1 >>
rect 211 71 212 72 
<< pdiffusion >>
rect 211 71 212 72 
<< pdiffusion >>
rect 212 71 213 72 
<< pdiffusion >>
rect 213 71 214 72 
<< pdiffusion >>
rect 214 71 215 72 
<< pdiffusion >>
rect 215 71 216 72 
<< pdiffusion >>
rect 228 71 229 72 
<< pdiffusion >>
rect 229 71 230 72 
<< pdiffusion >>
rect 230 71 231 72 
<< pdiffusion >>
rect 231 71 232 72 
<< m1 >>
rect 232 71 233 72 
<< pdiffusion >>
rect 232 71 233 72 
<< pdiffusion >>
rect 233 71 234 72 
<< m2 >>
rect 243 71 244 72 
<< m1 >>
rect 244 71 245 72 
<< pdiffusion >>
rect 246 71 247 72 
<< pdiffusion >>
rect 247 71 248 72 
<< pdiffusion >>
rect 248 71 249 72 
<< pdiffusion >>
rect 249 71 250 72 
<< pdiffusion >>
rect 250 71 251 72 
<< pdiffusion >>
rect 251 71 252 72 
<< m1 >>
rect 253 71 254 72 
<< m2 >>
rect 254 71 255 72 
<< m1 >>
rect 256 71 257 72 
<< m1 >>
rect 16 72 17 73 
<< m2 >>
rect 26 72 27 73 
<< m1 >>
rect 28 72 29 73 
<< m2 >>
rect 28 72 29 73 
<< m1 >>
rect 37 72 38 73 
<< m1 >>
rect 40 72 41 73 
<< m1 >>
rect 44 72 45 73 
<< m1 >>
rect 46 72 47 73 
<< m1 >>
rect 52 72 53 73 
<< m1 >>
rect 55 72 56 73 
<< m2 >>
rect 56 72 57 73 
<< m1 >>
rect 60 72 61 73 
<< m1 >>
rect 73 72 74 73 
<< m1 >>
rect 75 72 76 73 
<< m1 >>
rect 77 72 78 73 
<< m1 >>
rect 82 72 83 73 
<< m1 >>
rect 88 72 89 73 
<< m1 >>
rect 103 72 104 73 
<< m1 >>
rect 106 72 107 73 
<< m1 >>
rect 109 72 110 73 
<< m2 >>
rect 110 72 111 73 
<< m1 >>
rect 118 72 119 73 
<< m1 >>
rect 124 72 125 73 
<< m1 >>
rect 136 72 137 73 
<< m2 >>
rect 136 72 137 73 
<< m1 >>
rect 142 72 143 73 
<< m1 >>
rect 154 72 155 73 
<< m1 >>
rect 157 72 158 73 
<< m1 >>
rect 163 72 164 73 
<< m1 >>
rect 165 72 166 73 
<< m2 >>
rect 166 72 167 73 
<< m1 >>
rect 170 72 171 73 
<< m1 >>
rect 172 72 173 73 
<< m1 >>
rect 175 72 176 73 
<< m1 >>
rect 181 72 182 73 
<< m1 >>
rect 186 72 187 73 
<< m1 >>
rect 190 72 191 73 
<< m1 >>
rect 199 72 200 73 
<< m2 >>
rect 200 72 201 73 
<< m1 >>
rect 202 72 203 73 
<< m1 >>
rect 211 72 212 73 
<< m1 >>
rect 232 72 233 73 
<< m2 >>
rect 243 72 244 73 
<< m1 >>
rect 244 72 245 73 
<< m1 >>
rect 253 72 254 73 
<< m2 >>
rect 254 72 255 73 
<< m1 >>
rect 256 72 257 73 
<< m1 >>
rect 16 73 17 74 
<< m1 >>
rect 17 73 18 74 
<< m1 >>
rect 18 73 19 74 
<< m1 >>
rect 19 73 20 74 
<< m1 >>
rect 20 73 21 74 
<< m1 >>
rect 21 73 22 74 
<< m1 >>
rect 22 73 23 74 
<< m1 >>
rect 23 73 24 74 
<< m1 >>
rect 24 73 25 74 
<< m1 >>
rect 25 73 26 74 
<< m1 >>
rect 26 73 27 74 
<< m2 >>
rect 26 73 27 74 
<< m1 >>
rect 27 73 28 74 
<< m1 >>
rect 28 73 29 74 
<< m2 >>
rect 28 73 29 74 
<< m1 >>
rect 37 73 38 74 
<< m1 >>
rect 40 73 41 74 
<< m1 >>
rect 44 73 45 74 
<< m1 >>
rect 46 73 47 74 
<< m1 >>
rect 52 73 53 74 
<< m1 >>
rect 53 73 54 74 
<< m2 >>
rect 53 73 54 74 
<< m2c >>
rect 53 73 54 74 
<< m1 >>
rect 53 73 54 74 
<< m2 >>
rect 53 73 54 74 
<< m2 >>
rect 54 73 55 74 
<< m1 >>
rect 55 73 56 74 
<< m2 >>
rect 55 73 56 74 
<< m2 >>
rect 56 73 57 74 
<< m1 >>
rect 60 73 61 74 
<< m1 >>
rect 73 73 74 74 
<< m1 >>
rect 75 73 76 74 
<< m1 >>
rect 77 73 78 74 
<< m1 >>
rect 82 73 83 74 
<< m1 >>
rect 88 73 89 74 
<< m1 >>
rect 103 73 104 74 
<< m1 >>
rect 106 73 107 74 
<< m1 >>
rect 109 73 110 74 
<< m2 >>
rect 110 73 111 74 
<< m1 >>
rect 118 73 119 74 
<< m1 >>
rect 124 73 125 74 
<< m1 >>
rect 125 73 126 74 
<< m1 >>
rect 126 73 127 74 
<< m1 >>
rect 127 73 128 74 
<< m1 >>
rect 128 73 129 74 
<< m1 >>
rect 129 73 130 74 
<< m1 >>
rect 130 73 131 74 
<< m1 >>
rect 131 73 132 74 
<< m1 >>
rect 132 73 133 74 
<< m1 >>
rect 133 73 134 74 
<< m1 >>
rect 134 73 135 74 
<< m1 >>
rect 135 73 136 74 
<< m1 >>
rect 136 73 137 74 
<< m2 >>
rect 136 73 137 74 
<< m1 >>
rect 142 73 143 74 
<< m1 >>
rect 152 73 153 74 
<< m2 >>
rect 152 73 153 74 
<< m2c >>
rect 152 73 153 74 
<< m1 >>
rect 152 73 153 74 
<< m2 >>
rect 152 73 153 74 
<< m2 >>
rect 153 73 154 74 
<< m1 >>
rect 154 73 155 74 
<< m2 >>
rect 154 73 155 74 
<< m2 >>
rect 155 73 156 74 
<< m1 >>
rect 156 73 157 74 
<< m2 >>
rect 156 73 157 74 
<< m2c >>
rect 156 73 157 74 
<< m1 >>
rect 156 73 157 74 
<< m2 >>
rect 156 73 157 74 
<< m1 >>
rect 157 73 158 74 
<< m1 >>
rect 161 73 162 74 
<< m2 >>
rect 161 73 162 74 
<< m2c >>
rect 161 73 162 74 
<< m1 >>
rect 161 73 162 74 
<< m2 >>
rect 161 73 162 74 
<< m2 >>
rect 162 73 163 74 
<< m1 >>
rect 163 73 164 74 
<< m2 >>
rect 163 73 164 74 
<< m2 >>
rect 164 73 165 74 
<< m1 >>
rect 165 73 166 74 
<< m2 >>
rect 165 73 166 74 
<< m2 >>
rect 166 73 167 74 
<< m1 >>
rect 170 73 171 74 
<< m2 >>
rect 170 73 171 74 
<< m2c >>
rect 170 73 171 74 
<< m1 >>
rect 170 73 171 74 
<< m2 >>
rect 170 73 171 74 
<< m2 >>
rect 171 73 172 74 
<< m1 >>
rect 172 73 173 74 
<< m2 >>
rect 172 73 173 74 
<< m2 >>
rect 173 73 174 74 
<< m1 >>
rect 174 73 175 74 
<< m2 >>
rect 174 73 175 74 
<< m2c >>
rect 174 73 175 74 
<< m1 >>
rect 174 73 175 74 
<< m2 >>
rect 174 73 175 74 
<< m1 >>
rect 175 73 176 74 
<< m1 >>
rect 181 73 182 74 
<< m1 >>
rect 186 73 187 74 
<< m1 >>
rect 190 73 191 74 
<< m1 >>
rect 199 73 200 74 
<< m2 >>
rect 200 73 201 74 
<< m1 >>
rect 202 73 203 74 
<< m1 >>
rect 211 73 212 74 
<< m1 >>
rect 232 73 233 74 
<< m2 >>
rect 243 73 244 74 
<< m1 >>
rect 244 73 245 74 
<< m1 >>
rect 253 73 254 74 
<< m2 >>
rect 254 73 255 74 
<< m1 >>
rect 256 73 257 74 
<< m2 >>
rect 26 74 27 75 
<< m2 >>
rect 28 74 29 75 
<< m1 >>
rect 37 74 38 75 
<< m1 >>
rect 40 74 41 75 
<< m1 >>
rect 44 74 45 75 
<< m1 >>
rect 46 74 47 75 
<< m1 >>
rect 55 74 56 75 
<< m1 >>
rect 60 74 61 75 
<< m1 >>
rect 68 74 69 75 
<< m2 >>
rect 68 74 69 75 
<< m2c >>
rect 68 74 69 75 
<< m1 >>
rect 68 74 69 75 
<< m2 >>
rect 68 74 69 75 
<< m1 >>
rect 69 74 70 75 
<< m1 >>
rect 70 74 71 75 
<< m1 >>
rect 71 74 72 75 
<< m2 >>
rect 71 74 72 75 
<< m2c >>
rect 71 74 72 75 
<< m1 >>
rect 71 74 72 75 
<< m2 >>
rect 71 74 72 75 
<< m2 >>
rect 72 74 73 75 
<< m1 >>
rect 73 74 74 75 
<< m2 >>
rect 73 74 74 75 
<< m2 >>
rect 74 74 75 75 
<< m1 >>
rect 75 74 76 75 
<< m2 >>
rect 75 74 76 75 
<< m2c >>
rect 75 74 76 75 
<< m1 >>
rect 75 74 76 75 
<< m2 >>
rect 75 74 76 75 
<< m1 >>
rect 77 74 78 75 
<< m2 >>
rect 77 74 78 75 
<< m2c >>
rect 77 74 78 75 
<< m1 >>
rect 77 74 78 75 
<< m2 >>
rect 77 74 78 75 
<< m1 >>
rect 82 74 83 75 
<< m1 >>
rect 88 74 89 75 
<< m1 >>
rect 103 74 104 75 
<< m1 >>
rect 104 74 105 75 
<< m2 >>
rect 104 74 105 75 
<< m2c >>
rect 104 74 105 75 
<< m1 >>
rect 104 74 105 75 
<< m2 >>
rect 104 74 105 75 
<< m2 >>
rect 105 74 106 75 
<< m1 >>
rect 106 74 107 75 
<< m2 >>
rect 106 74 107 75 
<< m2 >>
rect 107 74 108 75 
<< m2 >>
rect 108 74 109 75 
<< m1 >>
rect 109 74 110 75 
<< m2 >>
rect 109 74 110 75 
<< m2 >>
rect 110 74 111 75 
<< m1 >>
rect 118 74 119 75 
<< m2 >>
rect 136 74 137 75 
<< m2 >>
rect 137 74 138 75 
<< m1 >>
rect 138 74 139 75 
<< m2 >>
rect 138 74 139 75 
<< m1 >>
rect 142 74 143 75 
<< m1 >>
rect 152 74 153 75 
<< m1 >>
rect 154 74 155 75 
<< m1 >>
rect 161 74 162 75 
<< m1 >>
rect 163 74 164 75 
<< m1 >>
rect 165 74 166 75 
<< m1 >>
rect 172 74 173 75 
<< m1 >>
rect 181 74 182 75 
<< m1 >>
rect 186 74 187 75 
<< m1 >>
rect 190 74 191 75 
<< m1 >>
rect 199 74 200 75 
<< m2 >>
rect 200 74 201 75 
<< m1 >>
rect 202 74 203 75 
<< m1 >>
rect 211 74 212 75 
<< m1 >>
rect 232 74 233 75 
<< m2 >>
rect 243 74 244 75 
<< m1 >>
rect 244 74 245 75 
<< m1 >>
rect 253 74 254 75 
<< m2 >>
rect 254 74 255 75 
<< m1 >>
rect 256 74 257 75 
<< m2 >>
rect 26 75 27 76 
<< m1 >>
rect 28 75 29 76 
<< m2 >>
rect 28 75 29 76 
<< m2c >>
rect 28 75 29 76 
<< m1 >>
rect 28 75 29 76 
<< m2 >>
rect 28 75 29 76 
<< m1 >>
rect 37 75 38 76 
<< m1 >>
rect 40 75 41 76 
<< m1 >>
rect 44 75 45 76 
<< m1 >>
rect 46 75 47 76 
<< m1 >>
rect 55 75 56 76 
<< m1 >>
rect 60 75 61 76 
<< m2 >>
rect 68 75 69 76 
<< m1 >>
rect 73 75 74 76 
<< m2 >>
rect 77 75 78 76 
<< m1 >>
rect 82 75 83 76 
<< m1 >>
rect 88 75 89 76 
<< m1 >>
rect 106 75 107 76 
<< m1 >>
rect 109 75 110 76 
<< m1 >>
rect 118 75 119 76 
<< m1 >>
rect 138 75 139 76 
<< m2 >>
rect 138 75 139 76 
<< m2c >>
rect 138 75 139 76 
<< m1 >>
rect 138 75 139 76 
<< m2 >>
rect 138 75 139 76 
<< m1 >>
rect 142 75 143 76 
<< m2 >>
rect 142 75 143 76 
<< m2c >>
rect 142 75 143 76 
<< m1 >>
rect 142 75 143 76 
<< m2 >>
rect 142 75 143 76 
<< m1 >>
rect 152 75 153 76 
<< m2 >>
rect 152 75 153 76 
<< m2c >>
rect 152 75 153 76 
<< m1 >>
rect 152 75 153 76 
<< m2 >>
rect 152 75 153 76 
<< m1 >>
rect 154 75 155 76 
<< m2 >>
rect 154 75 155 76 
<< m2c >>
rect 154 75 155 76 
<< m1 >>
rect 154 75 155 76 
<< m2 >>
rect 154 75 155 76 
<< m1 >>
rect 161 75 162 76 
<< m2 >>
rect 161 75 162 76 
<< m2c >>
rect 161 75 162 76 
<< m1 >>
rect 161 75 162 76 
<< m2 >>
rect 161 75 162 76 
<< m1 >>
rect 163 75 164 76 
<< m2 >>
rect 163 75 164 76 
<< m2c >>
rect 163 75 164 76 
<< m1 >>
rect 163 75 164 76 
<< m2 >>
rect 163 75 164 76 
<< m1 >>
rect 165 75 166 76 
<< m2 >>
rect 165 75 166 76 
<< m2c >>
rect 165 75 166 76 
<< m1 >>
rect 165 75 166 76 
<< m2 >>
rect 165 75 166 76 
<< m1 >>
rect 172 75 173 76 
<< m1 >>
rect 181 75 182 76 
<< m1 >>
rect 186 75 187 76 
<< m1 >>
rect 190 75 191 76 
<< m1 >>
rect 199 75 200 76 
<< m2 >>
rect 200 75 201 76 
<< m1 >>
rect 202 75 203 76 
<< m1 >>
rect 211 75 212 76 
<< m1 >>
rect 232 75 233 76 
<< m2 >>
rect 243 75 244 76 
<< m1 >>
rect 244 75 245 76 
<< m1 >>
rect 253 75 254 76 
<< m2 >>
rect 254 75 255 76 
<< m1 >>
rect 256 75 257 76 
<< m1 >>
rect 13 76 14 77 
<< m1 >>
rect 14 76 15 77 
<< m1 >>
rect 15 76 16 77 
<< m1 >>
rect 16 76 17 77 
<< m1 >>
rect 17 76 18 77 
<< m1 >>
rect 18 76 19 77 
<< m1 >>
rect 19 76 20 77 
<< m1 >>
rect 20 76 21 77 
<< m1 >>
rect 21 76 22 77 
<< m1 >>
rect 22 76 23 77 
<< m1 >>
rect 23 76 24 77 
<< m1 >>
rect 24 76 25 77 
<< m1 >>
rect 25 76 26 77 
<< m1 >>
rect 26 76 27 77 
<< m2 >>
rect 26 76 27 77 
<< m1 >>
rect 27 76 28 77 
<< m1 >>
rect 28 76 29 77 
<< m1 >>
rect 37 76 38 77 
<< m1 >>
rect 40 76 41 77 
<< m1 >>
rect 44 76 45 77 
<< m1 >>
rect 46 76 47 77 
<< m1 >>
rect 55 76 56 77 
<< m1 >>
rect 60 76 61 77 
<< m1 >>
rect 64 76 65 77 
<< m1 >>
rect 65 76 66 77 
<< m1 >>
rect 66 76 67 77 
<< m1 >>
rect 67 76 68 77 
<< m1 >>
rect 68 76 69 77 
<< m2 >>
rect 68 76 69 77 
<< m1 >>
rect 69 76 70 77 
<< m1 >>
rect 70 76 71 77 
<< m1 >>
rect 71 76 72 77 
<< m2 >>
rect 71 76 72 77 
<< m2c >>
rect 71 76 72 77 
<< m1 >>
rect 71 76 72 77 
<< m2 >>
rect 71 76 72 77 
<< m2 >>
rect 72 76 73 77 
<< m1 >>
rect 73 76 74 77 
<< m2 >>
rect 73 76 74 77 
<< m2 >>
rect 74 76 75 77 
<< m1 >>
rect 75 76 76 77 
<< m2 >>
rect 75 76 76 77 
<< m2c >>
rect 75 76 76 77 
<< m1 >>
rect 75 76 76 77 
<< m2 >>
rect 75 76 76 77 
<< m1 >>
rect 76 76 77 77 
<< m1 >>
rect 77 76 78 77 
<< m2 >>
rect 77 76 78 77 
<< m1 >>
rect 78 76 79 77 
<< m1 >>
rect 79 76 80 77 
<< m1 >>
rect 80 76 81 77 
<< m2 >>
rect 80 76 81 77 
<< m2c >>
rect 80 76 81 77 
<< m1 >>
rect 80 76 81 77 
<< m2 >>
rect 80 76 81 77 
<< m2 >>
rect 81 76 82 77 
<< m1 >>
rect 82 76 83 77 
<< m2 >>
rect 82 76 83 77 
<< m2 >>
rect 83 76 84 77 
<< m1 >>
rect 84 76 85 77 
<< m2 >>
rect 84 76 85 77 
<< m2c >>
rect 84 76 85 77 
<< m1 >>
rect 84 76 85 77 
<< m2 >>
rect 84 76 85 77 
<< m1 >>
rect 85 76 86 77 
<< m1 >>
rect 86 76 87 77 
<< m1 >>
rect 87 76 88 77 
<< m1 >>
rect 88 76 89 77 
<< m1 >>
rect 106 76 107 77 
<< m1 >>
rect 109 76 110 77 
<< m1 >>
rect 118 76 119 77 
<< m2 >>
rect 138 76 139 77 
<< m2 >>
rect 142 76 143 77 
<< m2 >>
rect 152 76 153 77 
<< m2 >>
rect 154 76 155 77 
<< m2 >>
rect 161 76 162 77 
<< m2 >>
rect 163 76 164 77 
<< m2 >>
rect 165 76 166 77 
<< m1 >>
rect 172 76 173 77 
<< m1 >>
rect 181 76 182 77 
<< m1 >>
rect 186 76 187 77 
<< m1 >>
rect 190 76 191 77 
<< m1 >>
rect 199 76 200 77 
<< m2 >>
rect 200 76 201 77 
<< m1 >>
rect 202 76 203 77 
<< m1 >>
rect 211 76 212 77 
<< m1 >>
rect 212 76 213 77 
<< m1 >>
rect 213 76 214 77 
<< m1 >>
rect 214 76 215 77 
<< m1 >>
rect 215 76 216 77 
<< m1 >>
rect 216 76 217 77 
<< m1 >>
rect 217 76 218 77 
<< m1 >>
rect 218 76 219 77 
<< m1 >>
rect 219 76 220 77 
<< m1 >>
rect 220 76 221 77 
<< m1 >>
rect 221 76 222 77 
<< m1 >>
rect 222 76 223 77 
<< m1 >>
rect 223 76 224 77 
<< m1 >>
rect 224 76 225 77 
<< m1 >>
rect 225 76 226 77 
<< m1 >>
rect 226 76 227 77 
<< m1 >>
rect 227 76 228 77 
<< m1 >>
rect 228 76 229 77 
<< m1 >>
rect 229 76 230 77 
<< m1 >>
rect 230 76 231 77 
<< m1 >>
rect 231 76 232 77 
<< m1 >>
rect 232 76 233 77 
<< m2 >>
rect 243 76 244 77 
<< m1 >>
rect 244 76 245 77 
<< m1 >>
rect 253 76 254 77 
<< m2 >>
rect 254 76 255 77 
<< m1 >>
rect 256 76 257 77 
<< m1 >>
rect 13 77 14 78 
<< m2 >>
rect 26 77 27 78 
<< m2 >>
rect 27 77 28 78 
<< m2 >>
rect 28 77 29 78 
<< m1 >>
rect 37 77 38 78 
<< m1 >>
rect 40 77 41 78 
<< m1 >>
rect 44 77 45 78 
<< m1 >>
rect 46 77 47 78 
<< m1 >>
rect 55 77 56 78 
<< m1 >>
rect 60 77 61 78 
<< m2 >>
rect 63 77 64 78 
<< m1 >>
rect 64 77 65 78 
<< m2 >>
rect 64 77 65 78 
<< m2 >>
rect 65 77 66 78 
<< m2 >>
rect 66 77 67 78 
<< m2 >>
rect 67 77 68 78 
<< m2 >>
rect 68 77 69 78 
<< m1 >>
rect 73 77 74 78 
<< m2 >>
rect 77 77 78 78 
<< m1 >>
rect 82 77 83 78 
<< m1 >>
rect 106 77 107 78 
<< m2 >>
rect 106 77 107 78 
<< m2c >>
rect 106 77 107 78 
<< m1 >>
rect 106 77 107 78 
<< m2 >>
rect 106 77 107 78 
<< m1 >>
rect 109 77 110 78 
<< m2 >>
rect 109 77 110 78 
<< m2c >>
rect 109 77 110 78 
<< m1 >>
rect 109 77 110 78 
<< m2 >>
rect 109 77 110 78 
<< m1 >>
rect 118 77 119 78 
<< m1 >>
rect 119 77 120 78 
<< m1 >>
rect 120 77 121 78 
<< m1 >>
rect 121 77 122 78 
<< m1 >>
rect 122 77 123 78 
<< m1 >>
rect 123 77 124 78 
<< m1 >>
rect 124 77 125 78 
<< m1 >>
rect 125 77 126 78 
<< m1 >>
rect 126 77 127 78 
<< m1 >>
rect 127 77 128 78 
<< m1 >>
rect 128 77 129 78 
<< m1 >>
rect 129 77 130 78 
<< m1 >>
rect 130 77 131 78 
<< m1 >>
rect 131 77 132 78 
<< m1 >>
rect 132 77 133 78 
<< m1 >>
rect 133 77 134 78 
<< m1 >>
rect 134 77 135 78 
<< m1 >>
rect 135 77 136 78 
<< m1 >>
rect 136 77 137 78 
<< m1 >>
rect 137 77 138 78 
<< m1 >>
rect 138 77 139 78 
<< m2 >>
rect 138 77 139 78 
<< m1 >>
rect 139 77 140 78 
<< m2 >>
rect 139 77 140 78 
<< m1 >>
rect 140 77 141 78 
<< m2 >>
rect 140 77 141 78 
<< m1 >>
rect 141 77 142 78 
<< m1 >>
rect 142 77 143 78 
<< m2 >>
rect 142 77 143 78 
<< m1 >>
rect 143 77 144 78 
<< m1 >>
rect 144 77 145 78 
<< m1 >>
rect 145 77 146 78 
<< m1 >>
rect 146 77 147 78 
<< m1 >>
rect 147 77 148 78 
<< m1 >>
rect 148 77 149 78 
<< m1 >>
rect 149 77 150 78 
<< m1 >>
rect 150 77 151 78 
<< m1 >>
rect 151 77 152 78 
<< m1 >>
rect 152 77 153 78 
<< m2 >>
rect 152 77 153 78 
<< m1 >>
rect 153 77 154 78 
<< m1 >>
rect 154 77 155 78 
<< m2 >>
rect 154 77 155 78 
<< m1 >>
rect 155 77 156 78 
<< m1 >>
rect 156 77 157 78 
<< m1 >>
rect 157 77 158 78 
<< m1 >>
rect 158 77 159 78 
<< m1 >>
rect 159 77 160 78 
<< m1 >>
rect 160 77 161 78 
<< m1 >>
rect 161 77 162 78 
<< m2 >>
rect 161 77 162 78 
<< m1 >>
rect 162 77 163 78 
<< m1 >>
rect 163 77 164 78 
<< m2 >>
rect 163 77 164 78 
<< m1 >>
rect 164 77 165 78 
<< m1 >>
rect 165 77 166 78 
<< m2 >>
rect 165 77 166 78 
<< m1 >>
rect 166 77 167 78 
<< m1 >>
rect 167 77 168 78 
<< m1 >>
rect 168 77 169 78 
<< m1 >>
rect 169 77 170 78 
<< m1 >>
rect 170 77 171 78 
<< m1 >>
rect 172 77 173 78 
<< m1 >>
rect 181 77 182 78 
<< m2 >>
rect 181 77 182 78 
<< m2c >>
rect 181 77 182 78 
<< m1 >>
rect 181 77 182 78 
<< m2 >>
rect 181 77 182 78 
<< m1 >>
rect 186 77 187 78 
<< m2 >>
rect 186 77 187 78 
<< m2c >>
rect 186 77 187 78 
<< m1 >>
rect 186 77 187 78 
<< m2 >>
rect 186 77 187 78 
<< m1 >>
rect 190 77 191 78 
<< m2 >>
rect 190 77 191 78 
<< m2c >>
rect 190 77 191 78 
<< m1 >>
rect 190 77 191 78 
<< m2 >>
rect 190 77 191 78 
<< m1 >>
rect 199 77 200 78 
<< m2 >>
rect 200 77 201 78 
<< m1 >>
rect 202 77 203 78 
<< m2 >>
rect 243 77 244 78 
<< m1 >>
rect 244 77 245 78 
<< m1 >>
rect 253 77 254 78 
<< m2 >>
rect 254 77 255 78 
<< m1 >>
rect 256 77 257 78 
<< m1 >>
rect 13 78 14 79 
<< m1 >>
rect 28 78 29 79 
<< m2 >>
rect 28 78 29 79 
<< m2c >>
rect 28 78 29 79 
<< m1 >>
rect 28 78 29 79 
<< m2 >>
rect 28 78 29 79 
<< m1 >>
rect 37 78 38 79 
<< m1 >>
rect 40 78 41 79 
<< m1 >>
rect 44 78 45 79 
<< m1 >>
rect 46 78 47 79 
<< m1 >>
rect 55 78 56 79 
<< m1 >>
rect 60 78 61 79 
<< m2 >>
rect 63 78 64 79 
<< m1 >>
rect 64 78 65 79 
<< m1 >>
rect 73 78 74 79 
<< m1 >>
rect 77 78 78 79 
<< m2 >>
rect 77 78 78 79 
<< m2c >>
rect 77 78 78 79 
<< m1 >>
rect 77 78 78 79 
<< m2 >>
rect 77 78 78 79 
<< m1 >>
rect 82 78 83 79 
<< m2 >>
rect 106 78 107 79 
<< m2 >>
rect 109 78 110 79 
<< m2 >>
rect 140 78 141 79 
<< m2 >>
rect 142 78 143 79 
<< m2 >>
rect 152 78 153 79 
<< m2 >>
rect 154 78 155 79 
<< m2 >>
rect 161 78 162 79 
<< m2 >>
rect 163 78 164 79 
<< m2 >>
rect 165 78 166 79 
<< m1 >>
rect 170 78 171 79 
<< m1 >>
rect 172 78 173 79 
<< m2 >>
rect 181 78 182 79 
<< m2 >>
rect 186 78 187 79 
<< m2 >>
rect 190 78 191 79 
<< m1 >>
rect 199 78 200 79 
<< m2 >>
rect 200 78 201 79 
<< m1 >>
rect 202 78 203 79 
<< m2 >>
rect 243 78 244 79 
<< m1 >>
rect 244 78 245 79 
<< m1 >>
rect 253 78 254 79 
<< m2 >>
rect 254 78 255 79 
<< m1 >>
rect 256 78 257 79 
<< m1 >>
rect 13 79 14 80 
<< m1 >>
rect 28 79 29 80 
<< m1 >>
rect 37 79 38 80 
<< m1 >>
rect 40 79 41 80 
<< m1 >>
rect 44 79 45 80 
<< m1 >>
rect 46 79 47 80 
<< m1 >>
rect 55 79 56 80 
<< m1 >>
rect 60 79 61 80 
<< m2 >>
rect 63 79 64 80 
<< m1 >>
rect 64 79 65 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m2c >>
rect 66 79 67 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m1 >>
rect 67 79 68 80 
<< m1 >>
rect 68 79 69 80 
<< m1 >>
rect 69 79 70 80 
<< m1 >>
rect 70 79 71 80 
<< m1 >>
rect 71 79 72 80 
<< m2 >>
rect 71 79 72 80 
<< m2c >>
rect 71 79 72 80 
<< m1 >>
rect 71 79 72 80 
<< m2 >>
rect 71 79 72 80 
<< m2 >>
rect 72 79 73 80 
<< m1 >>
rect 73 79 74 80 
<< m2 >>
rect 73 79 74 80 
<< m2 >>
rect 74 79 75 80 
<< m1 >>
rect 77 79 78 80 
<< m1 >>
rect 80 79 81 80 
<< m2 >>
rect 80 79 81 80 
<< m2c >>
rect 80 79 81 80 
<< m1 >>
rect 80 79 81 80 
<< m2 >>
rect 80 79 81 80 
<< m2 >>
rect 81 79 82 80 
<< m1 >>
rect 82 79 83 80 
<< m2 >>
rect 82 79 83 80 
<< m1 >>
rect 83 79 84 80 
<< m2 >>
rect 83 79 84 80 
<< m1 >>
rect 84 79 85 80 
<< m2 >>
rect 84 79 85 80 
<< m1 >>
rect 85 79 86 80 
<< m2 >>
rect 85 79 86 80 
<< m1 >>
rect 86 79 87 80 
<< m2 >>
rect 86 79 87 80 
<< m1 >>
rect 87 79 88 80 
<< m2 >>
rect 87 79 88 80 
<< m1 >>
rect 88 79 89 80 
<< m2 >>
rect 88 79 89 80 
<< m1 >>
rect 89 79 90 80 
<< m2 >>
rect 89 79 90 80 
<< m1 >>
rect 90 79 91 80 
<< m2 >>
rect 90 79 91 80 
<< m1 >>
rect 91 79 92 80 
<< m2 >>
rect 91 79 92 80 
<< m1 >>
rect 92 79 93 80 
<< m2 >>
rect 92 79 93 80 
<< m1 >>
rect 93 79 94 80 
<< m2 >>
rect 93 79 94 80 
<< m1 >>
rect 94 79 95 80 
<< m2 >>
rect 94 79 95 80 
<< m1 >>
rect 95 79 96 80 
<< m2 >>
rect 95 79 96 80 
<< m1 >>
rect 96 79 97 80 
<< m2 >>
rect 96 79 97 80 
<< m1 >>
rect 97 79 98 80 
<< m2 >>
rect 97 79 98 80 
<< m1 >>
rect 98 79 99 80 
<< m2 >>
rect 98 79 99 80 
<< m1 >>
rect 99 79 100 80 
<< m2 >>
rect 99 79 100 80 
<< m1 >>
rect 100 79 101 80 
<< m2 >>
rect 100 79 101 80 
<< m1 >>
rect 101 79 102 80 
<< m2 >>
rect 101 79 102 80 
<< m1 >>
rect 102 79 103 80 
<< m2 >>
rect 102 79 103 80 
<< m1 >>
rect 103 79 104 80 
<< m2 >>
rect 103 79 104 80 
<< m1 >>
rect 104 79 105 80 
<< m2 >>
rect 104 79 105 80 
<< m1 >>
rect 105 79 106 80 
<< m1 >>
rect 106 79 107 80 
<< m2 >>
rect 106 79 107 80 
<< m1 >>
rect 107 79 108 80 
<< m1 >>
rect 108 79 109 80 
<< m1 >>
rect 109 79 110 80 
<< m2 >>
rect 109 79 110 80 
<< m1 >>
rect 110 79 111 80 
<< m2 >>
rect 110 79 111 80 
<< m1 >>
rect 111 79 112 80 
<< m2 >>
rect 111 79 112 80 
<< m1 >>
rect 112 79 113 80 
<< m2 >>
rect 112 79 113 80 
<< m1 >>
rect 113 79 114 80 
<< m2 >>
rect 113 79 114 80 
<< m1 >>
rect 114 79 115 80 
<< m2 >>
rect 114 79 115 80 
<< m1 >>
rect 115 79 116 80 
<< m2 >>
rect 115 79 116 80 
<< m1 >>
rect 116 79 117 80 
<< m2 >>
rect 116 79 117 80 
<< m1 >>
rect 117 79 118 80 
<< m2 >>
rect 117 79 118 80 
<< m1 >>
rect 118 79 119 80 
<< m2 >>
rect 118 79 119 80 
<< m1 >>
rect 119 79 120 80 
<< m2 >>
rect 119 79 120 80 
<< m1 >>
rect 120 79 121 80 
<< m2 >>
rect 120 79 121 80 
<< m1 >>
rect 121 79 122 80 
<< m2 >>
rect 121 79 122 80 
<< m1 >>
rect 122 79 123 80 
<< m2 >>
rect 122 79 123 80 
<< m1 >>
rect 123 79 124 80 
<< m2 >>
rect 123 79 124 80 
<< m1 >>
rect 124 79 125 80 
<< m2 >>
rect 124 79 125 80 
<< m1 >>
rect 125 79 126 80 
<< m2 >>
rect 125 79 126 80 
<< m1 >>
rect 126 79 127 80 
<< m2 >>
rect 126 79 127 80 
<< m1 >>
rect 127 79 128 80 
<< m2 >>
rect 127 79 128 80 
<< m1 >>
rect 128 79 129 80 
<< m2 >>
rect 128 79 129 80 
<< m1 >>
rect 129 79 130 80 
<< m2 >>
rect 129 79 130 80 
<< m1 >>
rect 130 79 131 80 
<< m2 >>
rect 130 79 131 80 
<< m1 >>
rect 131 79 132 80 
<< m2 >>
rect 131 79 132 80 
<< m1 >>
rect 132 79 133 80 
<< m2 >>
rect 132 79 133 80 
<< m1 >>
rect 133 79 134 80 
<< m2 >>
rect 133 79 134 80 
<< m1 >>
rect 134 79 135 80 
<< m2 >>
rect 134 79 135 80 
<< m1 >>
rect 135 79 136 80 
<< m2 >>
rect 135 79 136 80 
<< m1 >>
rect 136 79 137 80 
<< m2 >>
rect 136 79 137 80 
<< m2 >>
rect 137 79 138 80 
<< m1 >>
rect 138 79 139 80 
<< m2 >>
rect 138 79 139 80 
<< m2c >>
rect 138 79 139 80 
<< m1 >>
rect 138 79 139 80 
<< m2 >>
rect 138 79 139 80 
<< m1 >>
rect 139 79 140 80 
<< m1 >>
rect 140 79 141 80 
<< m2 >>
rect 140 79 141 80 
<< m1 >>
rect 142 79 143 80 
<< m2 >>
rect 142 79 143 80 
<< m2c >>
rect 142 79 143 80 
<< m1 >>
rect 142 79 143 80 
<< m2 >>
rect 142 79 143 80 
<< m1 >>
rect 143 79 144 80 
<< m1 >>
rect 144 79 145 80 
<< m1 >>
rect 145 79 146 80 
<< m1 >>
rect 152 79 153 80 
<< m2 >>
rect 152 79 153 80 
<< m2c >>
rect 152 79 153 80 
<< m1 >>
rect 152 79 153 80 
<< m2 >>
rect 152 79 153 80 
<< m1 >>
rect 154 79 155 80 
<< m2 >>
rect 154 79 155 80 
<< m2c >>
rect 154 79 155 80 
<< m1 >>
rect 154 79 155 80 
<< m2 >>
rect 154 79 155 80 
<< m1 >>
rect 156 79 157 80 
<< m1 >>
rect 157 79 158 80 
<< m1 >>
rect 158 79 159 80 
<< m2 >>
rect 158 79 159 80 
<< m2c >>
rect 158 79 159 80 
<< m1 >>
rect 158 79 159 80 
<< m2 >>
rect 158 79 159 80 
<< m2 >>
rect 159 79 160 80 
<< m1 >>
rect 160 79 161 80 
<< m1 >>
rect 161 79 162 80 
<< m2 >>
rect 161 79 162 80 
<< m2c >>
rect 161 79 162 80 
<< m1 >>
rect 161 79 162 80 
<< m2 >>
rect 161 79 162 80 
<< m1 >>
rect 163 79 164 80 
<< m2 >>
rect 163 79 164 80 
<< m2c >>
rect 163 79 164 80 
<< m1 >>
rect 163 79 164 80 
<< m2 >>
rect 163 79 164 80 
<< m1 >>
rect 165 79 166 80 
<< m2 >>
rect 165 79 166 80 
<< m2c >>
rect 165 79 166 80 
<< m1 >>
rect 165 79 166 80 
<< m2 >>
rect 165 79 166 80 
<< m1 >>
rect 170 79 171 80 
<< m2 >>
rect 170 79 171 80 
<< m2c >>
rect 170 79 171 80 
<< m1 >>
rect 170 79 171 80 
<< m2 >>
rect 170 79 171 80 
<< m2 >>
rect 171 79 172 80 
<< m1 >>
rect 172 79 173 80 
<< m2 >>
rect 172 79 173 80 
<< m2 >>
rect 173 79 174 80 
<< m1 >>
rect 174 79 175 80 
<< m2 >>
rect 174 79 175 80 
<< m2c >>
rect 174 79 175 80 
<< m1 >>
rect 174 79 175 80 
<< m2 >>
rect 174 79 175 80 
<< m1 >>
rect 175 79 176 80 
<< m1 >>
rect 176 79 177 80 
<< m1 >>
rect 177 79 178 80 
<< m1 >>
rect 178 79 179 80 
<< m1 >>
rect 179 79 180 80 
<< m1 >>
rect 180 79 181 80 
<< m1 >>
rect 181 79 182 80 
<< m2 >>
rect 181 79 182 80 
<< m1 >>
rect 182 79 183 80 
<< m1 >>
rect 183 79 184 80 
<< m1 >>
rect 184 79 185 80 
<< m1 >>
rect 185 79 186 80 
<< m1 >>
rect 186 79 187 80 
<< m2 >>
rect 186 79 187 80 
<< m1 >>
rect 187 79 188 80 
<< m1 >>
rect 188 79 189 80 
<< m1 >>
rect 189 79 190 80 
<< m1 >>
rect 190 79 191 80 
<< m2 >>
rect 190 79 191 80 
<< m1 >>
rect 191 79 192 80 
<< m1 >>
rect 192 79 193 80 
<< m1 >>
rect 193 79 194 80 
<< m1 >>
rect 194 79 195 80 
<< m1 >>
rect 195 79 196 80 
<< m1 >>
rect 196 79 197 80 
<< m1 >>
rect 199 79 200 80 
<< m2 >>
rect 200 79 201 80 
<< m1 >>
rect 202 79 203 80 
<< m2 >>
rect 243 79 244 80 
<< m1 >>
rect 244 79 245 80 
<< m1 >>
rect 253 79 254 80 
<< m2 >>
rect 254 79 255 80 
<< m1 >>
rect 256 79 257 80 
<< m1 >>
rect 13 80 14 81 
<< m1 >>
rect 28 80 29 81 
<< m1 >>
rect 37 80 38 81 
<< m1 >>
rect 40 80 41 81 
<< m1 >>
rect 44 80 45 81 
<< m1 >>
rect 46 80 47 81 
<< m1 >>
rect 55 80 56 81 
<< m1 >>
rect 60 80 61 81 
<< m2 >>
rect 60 80 61 81 
<< m2c >>
rect 60 80 61 81 
<< m1 >>
rect 60 80 61 81 
<< m2 >>
rect 60 80 61 81 
<< m2 >>
rect 63 80 64 81 
<< m1 >>
rect 64 80 65 81 
<< m2 >>
rect 66 80 67 81 
<< m1 >>
rect 73 80 74 81 
<< m2 >>
rect 74 80 75 81 
<< m1 >>
rect 75 80 76 81 
<< m2 >>
rect 75 80 76 81 
<< m2c >>
rect 75 80 76 81 
<< m1 >>
rect 75 80 76 81 
<< m2 >>
rect 75 80 76 81 
<< m2 >>
rect 76 80 77 81 
<< m1 >>
rect 77 80 78 81 
<< m2 >>
rect 77 80 78 81 
<< m2 >>
rect 78 80 79 81 
<< m1 >>
rect 79 80 80 81 
<< m2 >>
rect 79 80 80 81 
<< m1 >>
rect 80 80 81 81 
<< m2 >>
rect 104 80 105 81 
<< m2 >>
rect 106 80 107 81 
<< m1 >>
rect 136 80 137 81 
<< m1 >>
rect 140 80 141 81 
<< m2 >>
rect 140 80 141 81 
<< m1 >>
rect 145 80 146 81 
<< m1 >>
rect 152 80 153 81 
<< m1 >>
rect 154 80 155 81 
<< m1 >>
rect 156 80 157 81 
<< m2 >>
rect 159 80 160 81 
<< m1 >>
rect 160 80 161 81 
<< m1 >>
rect 163 80 164 81 
<< m1 >>
rect 165 80 166 81 
<< m1 >>
rect 172 80 173 81 
<< m2 >>
rect 181 80 182 81 
<< m2 >>
rect 186 80 187 81 
<< m2 >>
rect 190 80 191 81 
<< m1 >>
rect 196 80 197 81 
<< m1 >>
rect 199 80 200 81 
<< m2 >>
rect 200 80 201 81 
<< m1 >>
rect 202 80 203 81 
<< m2 >>
rect 243 80 244 81 
<< m1 >>
rect 244 80 245 81 
<< m1 >>
rect 253 80 254 81 
<< m2 >>
rect 254 80 255 81 
<< m1 >>
rect 256 80 257 81 
<< m1 >>
rect 13 81 14 82 
<< m1 >>
rect 28 81 29 82 
<< m1 >>
rect 37 81 38 82 
<< m1 >>
rect 40 81 41 82 
<< m1 >>
rect 44 81 45 82 
<< m1 >>
rect 46 81 47 82 
<< m1 >>
rect 55 81 56 82 
<< m2 >>
rect 60 81 61 82 
<< m2 >>
rect 63 81 64 82 
<< m1 >>
rect 64 81 65 82 
<< m2 >>
rect 66 81 67 82 
<< m1 >>
rect 67 81 68 82 
<< m1 >>
rect 68 81 69 82 
<< m1 >>
rect 69 81 70 82 
<< m1 >>
rect 70 81 71 82 
<< m1 >>
rect 71 81 72 82 
<< m1 >>
rect 73 81 74 82 
<< m1 >>
rect 77 81 78 82 
<< m1 >>
rect 104 81 105 82 
<< m2 >>
rect 104 81 105 82 
<< m2c >>
rect 104 81 105 82 
<< m1 >>
rect 104 81 105 82 
<< m2 >>
rect 104 81 105 82 
<< m1 >>
rect 106 81 107 82 
<< m2 >>
rect 106 81 107 82 
<< m2c >>
rect 106 81 107 82 
<< m1 >>
rect 106 81 107 82 
<< m2 >>
rect 106 81 107 82 
<< m1 >>
rect 107 81 108 82 
<< m1 >>
rect 108 81 109 82 
<< m1 >>
rect 109 81 110 82 
<< m1 >>
rect 136 81 137 82 
<< m1 >>
rect 140 81 141 82 
<< m2 >>
rect 140 81 141 82 
<< m1 >>
rect 141 81 142 82 
<< m1 >>
rect 142 81 143 82 
<< m1 >>
rect 143 81 144 82 
<< m2 >>
rect 143 81 144 82 
<< m2c >>
rect 143 81 144 82 
<< m1 >>
rect 143 81 144 82 
<< m2 >>
rect 143 81 144 82 
<< m2 >>
rect 144 81 145 82 
<< m1 >>
rect 145 81 146 82 
<< m2 >>
rect 145 81 146 82 
<< m2 >>
rect 146 81 147 82 
<< m1 >>
rect 147 81 148 82 
<< m2 >>
rect 147 81 148 82 
<< m2c >>
rect 147 81 148 82 
<< m1 >>
rect 147 81 148 82 
<< m2 >>
rect 147 81 148 82 
<< m1 >>
rect 148 81 149 82 
<< m1 >>
rect 149 81 150 82 
<< m1 >>
rect 150 81 151 82 
<< m2 >>
rect 150 81 151 82 
<< m2c >>
rect 150 81 151 82 
<< m1 >>
rect 150 81 151 82 
<< m2 >>
rect 150 81 151 82 
<< m2 >>
rect 151 81 152 82 
<< m1 >>
rect 152 81 153 82 
<< m2 >>
rect 152 81 153 82 
<< m2 >>
rect 153 81 154 82 
<< m1 >>
rect 154 81 155 82 
<< m2 >>
rect 154 81 155 82 
<< m2 >>
rect 155 81 156 82 
<< m1 >>
rect 156 81 157 82 
<< m2 >>
rect 156 81 157 82 
<< m2c >>
rect 156 81 157 82 
<< m1 >>
rect 156 81 157 82 
<< m2 >>
rect 156 81 157 82 
<< m2 >>
rect 159 81 160 82 
<< m1 >>
rect 160 81 161 82 
<< m2 >>
rect 160 81 161 82 
<< m2 >>
rect 161 81 162 82 
<< m2 >>
rect 162 81 163 82 
<< m1 >>
rect 163 81 164 82 
<< m2 >>
rect 163 81 164 82 
<< m2 >>
rect 164 81 165 82 
<< m1 >>
rect 165 81 166 82 
<< m2 >>
rect 165 81 166 82 
<< m2 >>
rect 166 81 167 82 
<< m1 >>
rect 167 81 168 82 
<< m2 >>
rect 167 81 168 82 
<< m2c >>
rect 167 81 168 82 
<< m1 >>
rect 167 81 168 82 
<< m2 >>
rect 167 81 168 82 
<< m1 >>
rect 168 81 169 82 
<< m1 >>
rect 169 81 170 82 
<< m1 >>
rect 170 81 171 82 
<< m2 >>
rect 170 81 171 82 
<< m2c >>
rect 170 81 171 82 
<< m1 >>
rect 170 81 171 82 
<< m2 >>
rect 170 81 171 82 
<< m2 >>
rect 171 81 172 82 
<< m1 >>
rect 172 81 173 82 
<< m1 >>
rect 181 81 182 82 
<< m2 >>
rect 181 81 182 82 
<< m2c >>
rect 181 81 182 82 
<< m1 >>
rect 181 81 182 82 
<< m2 >>
rect 181 81 182 82 
<< m1 >>
rect 186 81 187 82 
<< m2 >>
rect 186 81 187 82 
<< m2c >>
rect 186 81 187 82 
<< m1 >>
rect 186 81 187 82 
<< m2 >>
rect 186 81 187 82 
<< m1 >>
rect 190 81 191 82 
<< m2 >>
rect 190 81 191 82 
<< m2c >>
rect 190 81 191 82 
<< m1 >>
rect 190 81 191 82 
<< m2 >>
rect 190 81 191 82 
<< m2 >>
rect 195 81 196 82 
<< m1 >>
rect 196 81 197 82 
<< m2 >>
rect 196 81 197 82 
<< m2 >>
rect 197 81 198 82 
<< m1 >>
rect 198 81 199 82 
<< m2 >>
rect 198 81 199 82 
<< m2c >>
rect 198 81 199 82 
<< m1 >>
rect 198 81 199 82 
<< m2 >>
rect 198 81 199 82 
<< m1 >>
rect 199 81 200 82 
<< m2 >>
rect 200 81 201 82 
<< m1 >>
rect 202 81 203 82 
<< m1 >>
rect 211 81 212 82 
<< m1 >>
rect 212 81 213 82 
<< m1 >>
rect 213 81 214 82 
<< m1 >>
rect 214 81 215 82 
<< m1 >>
rect 215 81 216 82 
<< m2 >>
rect 243 81 244 82 
<< m1 >>
rect 244 81 245 82 
<< m1 >>
rect 253 81 254 82 
<< m2 >>
rect 254 81 255 82 
<< m1 >>
rect 256 81 257 82 
<< m1 >>
rect 13 82 14 83 
<< m1 >>
rect 16 82 17 83 
<< m1 >>
rect 17 82 18 83 
<< m1 >>
rect 18 82 19 83 
<< m1 >>
rect 19 82 20 83 
<< m1 >>
rect 28 82 29 83 
<< m1 >>
rect 37 82 38 83 
<< m1 >>
rect 40 82 41 83 
<< m1 >>
rect 44 82 45 83 
<< m1 >>
rect 46 82 47 83 
<< m1 >>
rect 52 82 53 83 
<< m1 >>
rect 53 82 54 83 
<< m2 >>
rect 53 82 54 83 
<< m2c >>
rect 53 82 54 83 
<< m1 >>
rect 53 82 54 83 
<< m2 >>
rect 53 82 54 83 
<< m2 >>
rect 54 82 55 83 
<< m1 >>
rect 55 82 56 83 
<< m2 >>
rect 55 82 56 83 
<< m2 >>
rect 56 82 57 83 
<< m1 >>
rect 57 82 58 83 
<< m2 >>
rect 57 82 58 83 
<< m2c >>
rect 57 82 58 83 
<< m1 >>
rect 57 82 58 83 
<< m2 >>
rect 57 82 58 83 
<< m1 >>
rect 58 82 59 83 
<< m1 >>
rect 59 82 60 83 
<< m1 >>
rect 60 82 61 83 
<< m2 >>
rect 60 82 61 83 
<< m1 >>
rect 61 82 62 83 
<< m1 >>
rect 62 82 63 83 
<< m2 >>
rect 62 82 63 83 
<< m2c >>
rect 62 82 63 83 
<< m1 >>
rect 62 82 63 83 
<< m2 >>
rect 62 82 63 83 
<< m2 >>
rect 63 82 64 83 
<< m1 >>
rect 64 82 65 83 
<< m2 >>
rect 64 82 65 83 
<< m2 >>
rect 65 82 66 83 
<< m2 >>
rect 66 82 67 83 
<< m1 >>
rect 67 82 68 83 
<< m1 >>
rect 71 82 72 83 
<< m2 >>
rect 71 82 72 83 
<< m2c >>
rect 71 82 72 83 
<< m1 >>
rect 71 82 72 83 
<< m2 >>
rect 71 82 72 83 
<< m2 >>
rect 72 82 73 83 
<< m1 >>
rect 73 82 74 83 
<< m2 >>
rect 73 82 74 83 
<< m2 >>
rect 74 82 75 83 
<< m1 >>
rect 77 82 78 83 
<< m1 >>
rect 88 82 89 83 
<< m1 >>
rect 89 82 90 83 
<< m1 >>
rect 90 82 91 83 
<< m1 >>
rect 91 82 92 83 
<< m1 >>
rect 92 82 93 83 
<< m1 >>
rect 93 82 94 83 
<< m1 >>
rect 94 82 95 83 
<< m1 >>
rect 95 82 96 83 
<< m1 >>
rect 96 82 97 83 
<< m1 >>
rect 97 82 98 83 
<< m1 >>
rect 98 82 99 83 
<< m1 >>
rect 99 82 100 83 
<< m1 >>
rect 100 82 101 83 
<< m1 >>
rect 101 82 102 83 
<< m1 >>
rect 102 82 103 83 
<< m1 >>
rect 104 82 105 83 
<< m1 >>
rect 109 82 110 83 
<< m1 >>
rect 136 82 137 83 
<< m2 >>
rect 139 82 140 83 
<< m2 >>
rect 140 82 141 83 
<< m1 >>
rect 145 82 146 83 
<< m1 >>
rect 152 82 153 83 
<< m1 >>
rect 154 82 155 83 
<< m1 >>
rect 160 82 161 83 
<< m1 >>
rect 163 82 164 83 
<< m1 >>
rect 165 82 166 83 
<< m2 >>
rect 171 82 172 83 
<< m1 >>
rect 172 82 173 83 
<< m1 >>
rect 181 82 182 83 
<< m2 >>
rect 186 82 187 83 
<< m1 >>
rect 190 82 191 83 
<< m1 >>
rect 193 82 194 83 
<< m1 >>
rect 194 82 195 83 
<< m2 >>
rect 194 82 195 83 
<< m2c >>
rect 194 82 195 83 
<< m1 >>
rect 194 82 195 83 
<< m2 >>
rect 194 82 195 83 
<< m2 >>
rect 195 82 196 83 
<< m1 >>
rect 196 82 197 83 
<< m2 >>
rect 200 82 201 83 
<< m1 >>
rect 202 82 203 83 
<< m1 >>
rect 211 82 212 83 
<< m1 >>
rect 215 82 216 83 
<< m2 >>
rect 215 82 216 83 
<< m2c >>
rect 215 82 216 83 
<< m1 >>
rect 215 82 216 83 
<< m2 >>
rect 215 82 216 83 
<< m2 >>
rect 216 82 217 83 
<< m1 >>
rect 217 82 218 83 
<< m2 >>
rect 217 82 218 83 
<< m1 >>
rect 218 82 219 83 
<< m2 >>
rect 218 82 219 83 
<< m1 >>
rect 219 82 220 83 
<< m1 >>
rect 220 82 221 83 
<< m1 >>
rect 221 82 222 83 
<< m1 >>
rect 222 82 223 83 
<< m1 >>
rect 223 82 224 83 
<< m1 >>
rect 224 82 225 83 
<< m1 >>
rect 225 82 226 83 
<< m1 >>
rect 226 82 227 83 
<< m1 >>
rect 227 82 228 83 
<< m1 >>
rect 228 82 229 83 
<< m1 >>
rect 229 82 230 83 
<< m2 >>
rect 243 82 244 83 
<< m1 >>
rect 244 82 245 83 
<< m1 >>
rect 253 82 254 83 
<< m2 >>
rect 254 82 255 83 
<< m1 >>
rect 256 82 257 83 
<< m1 >>
rect 13 83 14 84 
<< m1 >>
rect 16 83 17 84 
<< m1 >>
rect 19 83 20 84 
<< m1 >>
rect 28 83 29 84 
<< m1 >>
rect 37 83 38 84 
<< m1 >>
rect 40 83 41 84 
<< m1 >>
rect 44 83 45 84 
<< m1 >>
rect 46 83 47 84 
<< m1 >>
rect 52 83 53 84 
<< m1 >>
rect 55 83 56 84 
<< m2 >>
rect 60 83 61 84 
<< m1 >>
rect 64 83 65 84 
<< m2 >>
rect 64 83 65 84 
<< m1 >>
rect 67 83 68 84 
<< m1 >>
rect 73 83 74 84 
<< m2 >>
rect 74 83 75 84 
<< m1 >>
rect 77 83 78 84 
<< m1 >>
rect 88 83 89 84 
<< m1 >>
rect 102 83 103 84 
<< m1 >>
rect 104 83 105 84 
<< m1 >>
rect 109 83 110 84 
<< m1 >>
rect 136 83 137 84 
<< m1 >>
rect 139 83 140 84 
<< m2 >>
rect 139 83 140 84 
<< m1 >>
rect 145 83 146 84 
<< m1 >>
rect 152 83 153 84 
<< m1 >>
rect 154 83 155 84 
<< m1 >>
rect 160 83 161 84 
<< m1 >>
rect 163 83 164 84 
<< m1 >>
rect 165 83 166 84 
<< m2 >>
rect 171 83 172 84 
<< m1 >>
rect 172 83 173 84 
<< m1 >>
rect 181 83 182 84 
<< m1 >>
rect 182 83 183 84 
<< m1 >>
rect 183 83 184 84 
<< m1 >>
rect 184 83 185 84 
<< m1 >>
rect 185 83 186 84 
<< m1 >>
rect 186 83 187 84 
<< m2 >>
rect 186 83 187 84 
<< m1 >>
rect 187 83 188 84 
<< m1 >>
rect 188 83 189 84 
<< m2 >>
rect 188 83 189 84 
<< m2c >>
rect 188 83 189 84 
<< m1 >>
rect 188 83 189 84 
<< m2 >>
rect 188 83 189 84 
<< m2 >>
rect 189 83 190 84 
<< m1 >>
rect 190 83 191 84 
<< m1 >>
rect 193 83 194 84 
<< m1 >>
rect 196 83 197 84 
<< m1 >>
rect 200 83 201 84 
<< m2 >>
rect 200 83 201 84 
<< m2c >>
rect 200 83 201 84 
<< m1 >>
rect 200 83 201 84 
<< m2 >>
rect 200 83 201 84 
<< m1 >>
rect 202 83 203 84 
<< m1 >>
rect 211 83 212 84 
<< m1 >>
rect 217 83 218 84 
<< m2 >>
rect 218 83 219 84 
<< m1 >>
rect 229 83 230 84 
<< m2 >>
rect 243 83 244 84 
<< m1 >>
rect 244 83 245 84 
<< m1 >>
rect 253 83 254 84 
<< m2 >>
rect 254 83 255 84 
<< m1 >>
rect 256 83 257 84 
<< pdiffusion >>
rect 12 84 13 85 
<< m1 >>
rect 13 84 14 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< m1 >>
rect 16 84 17 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< m1 >>
rect 19 84 20 85 
<< m1 >>
rect 28 84 29 85 
<< pdiffusion >>
rect 30 84 31 85 
<< pdiffusion >>
rect 31 84 32 85 
<< pdiffusion >>
rect 32 84 33 85 
<< pdiffusion >>
rect 33 84 34 85 
<< pdiffusion >>
rect 34 84 35 85 
<< pdiffusion >>
rect 35 84 36 85 
<< m1 >>
rect 37 84 38 85 
<< m1 >>
rect 40 84 41 85 
<< m1 >>
rect 44 84 45 85 
<< m1 >>
rect 46 84 47 85 
<< pdiffusion >>
rect 48 84 49 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< m1 >>
rect 52 84 53 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< m1 >>
rect 55 84 56 85 
<< m1 >>
rect 60 84 61 85 
<< m2 >>
rect 60 84 61 85 
<< m2c >>
rect 60 84 61 85 
<< m1 >>
rect 60 84 61 85 
<< m2 >>
rect 60 84 61 85 
<< m1 >>
rect 61 84 62 85 
<< m1 >>
rect 62 84 63 85 
<< m2 >>
rect 62 84 63 85 
<< m2c >>
rect 62 84 63 85 
<< m1 >>
rect 62 84 63 85 
<< m2 >>
rect 62 84 63 85 
<< m2 >>
rect 63 84 64 85 
<< m1 >>
rect 64 84 65 85 
<< m2 >>
rect 64 84 65 85 
<< pdiffusion >>
rect 66 84 67 85 
<< m1 >>
rect 67 84 68 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< m1 >>
rect 73 84 74 85 
<< m2 >>
rect 74 84 75 85 
<< m1 >>
rect 77 84 78 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< m1 >>
rect 88 84 89 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 102 84 103 85 
<< m1 >>
rect 104 84 105 85 
<< m1 >>
rect 109 84 110 85 
<< pdiffusion >>
rect 120 84 121 85 
<< pdiffusion >>
rect 121 84 122 85 
<< pdiffusion >>
rect 122 84 123 85 
<< pdiffusion >>
rect 123 84 124 85 
<< pdiffusion >>
rect 124 84 125 85 
<< pdiffusion >>
rect 125 84 126 85 
<< m1 >>
rect 136 84 137 85 
<< m1 >>
rect 138 84 139 85 
<< m2 >>
rect 138 84 139 85 
<< m2c >>
rect 138 84 139 85 
<< m1 >>
rect 138 84 139 85 
<< m2 >>
rect 138 84 139 85 
<< pdiffusion >>
rect 138 84 139 85 
<< m1 >>
rect 139 84 140 85 
<< pdiffusion >>
rect 139 84 140 85 
<< pdiffusion >>
rect 140 84 141 85 
<< pdiffusion >>
rect 141 84 142 85 
<< pdiffusion >>
rect 142 84 143 85 
<< pdiffusion >>
rect 143 84 144 85 
<< m1 >>
rect 145 84 146 85 
<< m1 >>
rect 152 84 153 85 
<< m1 >>
rect 154 84 155 85 
<< pdiffusion >>
rect 156 84 157 85 
<< pdiffusion >>
rect 157 84 158 85 
<< pdiffusion >>
rect 158 84 159 85 
<< pdiffusion >>
rect 159 84 160 85 
<< m1 >>
rect 160 84 161 85 
<< pdiffusion >>
rect 160 84 161 85 
<< pdiffusion >>
rect 161 84 162 85 
<< m1 >>
rect 163 84 164 85 
<< m1 >>
rect 165 84 166 85 
<< m2 >>
rect 171 84 172 85 
<< m1 >>
rect 172 84 173 85 
<< pdiffusion >>
rect 174 84 175 85 
<< pdiffusion >>
rect 175 84 176 85 
<< pdiffusion >>
rect 176 84 177 85 
<< pdiffusion >>
rect 177 84 178 85 
<< pdiffusion >>
rect 178 84 179 85 
<< pdiffusion >>
rect 179 84 180 85 
<< m2 >>
rect 186 84 187 85 
<< m2 >>
rect 189 84 190 85 
<< m1 >>
rect 190 84 191 85 
<< pdiffusion >>
rect 192 84 193 85 
<< m1 >>
rect 193 84 194 85 
<< pdiffusion >>
rect 193 84 194 85 
<< pdiffusion >>
rect 194 84 195 85 
<< pdiffusion >>
rect 195 84 196 85 
<< m1 >>
rect 196 84 197 85 
<< pdiffusion >>
rect 196 84 197 85 
<< pdiffusion >>
rect 197 84 198 85 
<< m1 >>
rect 200 84 201 85 
<< m1 >>
rect 202 84 203 85 
<< pdiffusion >>
rect 210 84 211 85 
<< m1 >>
rect 211 84 212 85 
<< pdiffusion >>
rect 211 84 212 85 
<< pdiffusion >>
rect 212 84 213 85 
<< pdiffusion >>
rect 213 84 214 85 
<< pdiffusion >>
rect 214 84 215 85 
<< pdiffusion >>
rect 215 84 216 85 
<< m1 >>
rect 217 84 218 85 
<< m2 >>
rect 218 84 219 85 
<< pdiffusion >>
rect 228 84 229 85 
<< m1 >>
rect 229 84 230 85 
<< pdiffusion >>
rect 229 84 230 85 
<< pdiffusion >>
rect 230 84 231 85 
<< pdiffusion >>
rect 231 84 232 85 
<< pdiffusion >>
rect 232 84 233 85 
<< pdiffusion >>
rect 233 84 234 85 
<< m2 >>
rect 243 84 244 85 
<< m1 >>
rect 244 84 245 85 
<< pdiffusion >>
rect 246 84 247 85 
<< pdiffusion >>
rect 247 84 248 85 
<< pdiffusion >>
rect 248 84 249 85 
<< pdiffusion >>
rect 249 84 250 85 
<< pdiffusion >>
rect 250 84 251 85 
<< pdiffusion >>
rect 251 84 252 85 
<< m1 >>
rect 253 84 254 85 
<< m2 >>
rect 254 84 255 85 
<< m1 >>
rect 256 84 257 85 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< m1 >>
rect 19 85 20 86 
<< m1 >>
rect 28 85 29 86 
<< pdiffusion >>
rect 30 85 31 86 
<< pdiffusion >>
rect 31 85 32 86 
<< pdiffusion >>
rect 32 85 33 86 
<< pdiffusion >>
rect 33 85 34 86 
<< pdiffusion >>
rect 34 85 35 86 
<< pdiffusion >>
rect 35 85 36 86 
<< m1 >>
rect 37 85 38 86 
<< m1 >>
rect 40 85 41 86 
<< m1 >>
rect 44 85 45 86 
<< m1 >>
rect 46 85 47 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< m1 >>
rect 55 85 56 86 
<< m1 >>
rect 64 85 65 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< m1 >>
rect 73 85 74 86 
<< m2 >>
rect 74 85 75 86 
<< m1 >>
rect 77 85 78 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 102 85 103 86 
<< m1 >>
rect 104 85 105 86 
<< m1 >>
rect 109 85 110 86 
<< pdiffusion >>
rect 120 85 121 86 
<< pdiffusion >>
rect 121 85 122 86 
<< pdiffusion >>
rect 122 85 123 86 
<< pdiffusion >>
rect 123 85 124 86 
<< pdiffusion >>
rect 124 85 125 86 
<< pdiffusion >>
rect 125 85 126 86 
<< m1 >>
rect 136 85 137 86 
<< pdiffusion >>
rect 138 85 139 86 
<< pdiffusion >>
rect 139 85 140 86 
<< pdiffusion >>
rect 140 85 141 86 
<< pdiffusion >>
rect 141 85 142 86 
<< pdiffusion >>
rect 142 85 143 86 
<< pdiffusion >>
rect 143 85 144 86 
<< m1 >>
rect 145 85 146 86 
<< m1 >>
rect 152 85 153 86 
<< m1 >>
rect 154 85 155 86 
<< pdiffusion >>
rect 156 85 157 86 
<< pdiffusion >>
rect 157 85 158 86 
<< pdiffusion >>
rect 158 85 159 86 
<< pdiffusion >>
rect 159 85 160 86 
<< pdiffusion >>
rect 160 85 161 86 
<< pdiffusion >>
rect 161 85 162 86 
<< m1 >>
rect 163 85 164 86 
<< m1 >>
rect 165 85 166 86 
<< m2 >>
rect 171 85 172 86 
<< m1 >>
rect 172 85 173 86 
<< pdiffusion >>
rect 174 85 175 86 
<< pdiffusion >>
rect 175 85 176 86 
<< pdiffusion >>
rect 176 85 177 86 
<< pdiffusion >>
rect 177 85 178 86 
<< pdiffusion >>
rect 178 85 179 86 
<< pdiffusion >>
rect 179 85 180 86 
<< m1 >>
rect 186 85 187 86 
<< m2 >>
rect 186 85 187 86 
<< m2c >>
rect 186 85 187 86 
<< m1 >>
rect 186 85 187 86 
<< m2 >>
rect 186 85 187 86 
<< m2 >>
rect 189 85 190 86 
<< m1 >>
rect 190 85 191 86 
<< pdiffusion >>
rect 192 85 193 86 
<< pdiffusion >>
rect 193 85 194 86 
<< pdiffusion >>
rect 194 85 195 86 
<< pdiffusion >>
rect 195 85 196 86 
<< pdiffusion >>
rect 196 85 197 86 
<< pdiffusion >>
rect 197 85 198 86 
<< m1 >>
rect 200 85 201 86 
<< m2 >>
rect 201 85 202 86 
<< m1 >>
rect 202 85 203 86 
<< m2 >>
rect 202 85 203 86 
<< m2c >>
rect 202 85 203 86 
<< m1 >>
rect 202 85 203 86 
<< m2 >>
rect 202 85 203 86 
<< pdiffusion >>
rect 210 85 211 86 
<< pdiffusion >>
rect 211 85 212 86 
<< pdiffusion >>
rect 212 85 213 86 
<< pdiffusion >>
rect 213 85 214 86 
<< pdiffusion >>
rect 214 85 215 86 
<< pdiffusion >>
rect 215 85 216 86 
<< m1 >>
rect 217 85 218 86 
<< m2 >>
rect 218 85 219 86 
<< pdiffusion >>
rect 228 85 229 86 
<< pdiffusion >>
rect 229 85 230 86 
<< pdiffusion >>
rect 230 85 231 86 
<< pdiffusion >>
rect 231 85 232 86 
<< pdiffusion >>
rect 232 85 233 86 
<< pdiffusion >>
rect 233 85 234 86 
<< m2 >>
rect 243 85 244 86 
<< m1 >>
rect 244 85 245 86 
<< pdiffusion >>
rect 246 85 247 86 
<< pdiffusion >>
rect 247 85 248 86 
<< pdiffusion >>
rect 248 85 249 86 
<< pdiffusion >>
rect 249 85 250 86 
<< pdiffusion >>
rect 250 85 251 86 
<< pdiffusion >>
rect 251 85 252 86 
<< m1 >>
rect 253 85 254 86 
<< m2 >>
rect 254 85 255 86 
<< m1 >>
rect 256 85 257 86 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< m1 >>
rect 19 86 20 87 
<< m1 >>
rect 28 86 29 87 
<< pdiffusion >>
rect 30 86 31 87 
<< pdiffusion >>
rect 31 86 32 87 
<< pdiffusion >>
rect 32 86 33 87 
<< pdiffusion >>
rect 33 86 34 87 
<< pdiffusion >>
rect 34 86 35 87 
<< pdiffusion >>
rect 35 86 36 87 
<< m1 >>
rect 37 86 38 87 
<< m1 >>
rect 40 86 41 87 
<< m1 >>
rect 44 86 45 87 
<< m1 >>
rect 46 86 47 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< m1 >>
rect 55 86 56 87 
<< m1 >>
rect 64 86 65 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< m1 >>
rect 73 86 74 87 
<< m2 >>
rect 74 86 75 87 
<< m1 >>
rect 77 86 78 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 102 86 103 87 
<< m1 >>
rect 104 86 105 87 
<< m1 >>
rect 109 86 110 87 
<< pdiffusion >>
rect 120 86 121 87 
<< pdiffusion >>
rect 121 86 122 87 
<< pdiffusion >>
rect 122 86 123 87 
<< pdiffusion >>
rect 123 86 124 87 
<< pdiffusion >>
rect 124 86 125 87 
<< pdiffusion >>
rect 125 86 126 87 
<< m1 >>
rect 136 86 137 87 
<< pdiffusion >>
rect 138 86 139 87 
<< pdiffusion >>
rect 139 86 140 87 
<< pdiffusion >>
rect 140 86 141 87 
<< pdiffusion >>
rect 141 86 142 87 
<< pdiffusion >>
rect 142 86 143 87 
<< pdiffusion >>
rect 143 86 144 87 
<< m1 >>
rect 145 86 146 87 
<< m1 >>
rect 152 86 153 87 
<< m1 >>
rect 154 86 155 87 
<< pdiffusion >>
rect 156 86 157 87 
<< pdiffusion >>
rect 157 86 158 87 
<< pdiffusion >>
rect 158 86 159 87 
<< pdiffusion >>
rect 159 86 160 87 
<< pdiffusion >>
rect 160 86 161 87 
<< pdiffusion >>
rect 161 86 162 87 
<< m1 >>
rect 163 86 164 87 
<< m1 >>
rect 165 86 166 87 
<< m2 >>
rect 171 86 172 87 
<< m1 >>
rect 172 86 173 87 
<< pdiffusion >>
rect 174 86 175 87 
<< pdiffusion >>
rect 175 86 176 87 
<< pdiffusion >>
rect 176 86 177 87 
<< pdiffusion >>
rect 177 86 178 87 
<< pdiffusion >>
rect 178 86 179 87 
<< pdiffusion >>
rect 179 86 180 87 
<< m1 >>
rect 186 86 187 87 
<< m2 >>
rect 189 86 190 87 
<< m1 >>
rect 190 86 191 87 
<< pdiffusion >>
rect 192 86 193 87 
<< pdiffusion >>
rect 193 86 194 87 
<< pdiffusion >>
rect 194 86 195 87 
<< pdiffusion >>
rect 195 86 196 87 
<< pdiffusion >>
rect 196 86 197 87 
<< pdiffusion >>
rect 197 86 198 87 
<< m1 >>
rect 200 86 201 87 
<< m2 >>
rect 201 86 202 87 
<< pdiffusion >>
rect 210 86 211 87 
<< pdiffusion >>
rect 211 86 212 87 
<< pdiffusion >>
rect 212 86 213 87 
<< pdiffusion >>
rect 213 86 214 87 
<< pdiffusion >>
rect 214 86 215 87 
<< pdiffusion >>
rect 215 86 216 87 
<< m1 >>
rect 217 86 218 87 
<< m2 >>
rect 218 86 219 87 
<< pdiffusion >>
rect 228 86 229 87 
<< pdiffusion >>
rect 229 86 230 87 
<< pdiffusion >>
rect 230 86 231 87 
<< pdiffusion >>
rect 231 86 232 87 
<< pdiffusion >>
rect 232 86 233 87 
<< pdiffusion >>
rect 233 86 234 87 
<< m2 >>
rect 243 86 244 87 
<< m1 >>
rect 244 86 245 87 
<< pdiffusion >>
rect 246 86 247 87 
<< pdiffusion >>
rect 247 86 248 87 
<< pdiffusion >>
rect 248 86 249 87 
<< pdiffusion >>
rect 249 86 250 87 
<< pdiffusion >>
rect 250 86 251 87 
<< pdiffusion >>
rect 251 86 252 87 
<< m1 >>
rect 253 86 254 87 
<< m2 >>
rect 254 86 255 87 
<< m1 >>
rect 256 86 257 87 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< m1 >>
rect 19 87 20 88 
<< m1 >>
rect 28 87 29 88 
<< pdiffusion >>
rect 30 87 31 88 
<< pdiffusion >>
rect 31 87 32 88 
<< pdiffusion >>
rect 32 87 33 88 
<< pdiffusion >>
rect 33 87 34 88 
<< pdiffusion >>
rect 34 87 35 88 
<< pdiffusion >>
rect 35 87 36 88 
<< m1 >>
rect 37 87 38 88 
<< m1 >>
rect 40 87 41 88 
<< m1 >>
rect 44 87 45 88 
<< m1 >>
rect 46 87 47 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< m1 >>
rect 55 87 56 88 
<< m1 >>
rect 64 87 65 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< m1 >>
rect 73 87 74 88 
<< m2 >>
rect 74 87 75 88 
<< m1 >>
rect 77 87 78 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 102 87 103 88 
<< m1 >>
rect 104 87 105 88 
<< m1 >>
rect 109 87 110 88 
<< pdiffusion >>
rect 120 87 121 88 
<< pdiffusion >>
rect 121 87 122 88 
<< pdiffusion >>
rect 122 87 123 88 
<< pdiffusion >>
rect 123 87 124 88 
<< pdiffusion >>
rect 124 87 125 88 
<< pdiffusion >>
rect 125 87 126 88 
<< m1 >>
rect 136 87 137 88 
<< pdiffusion >>
rect 138 87 139 88 
<< pdiffusion >>
rect 139 87 140 88 
<< pdiffusion >>
rect 140 87 141 88 
<< pdiffusion >>
rect 141 87 142 88 
<< pdiffusion >>
rect 142 87 143 88 
<< pdiffusion >>
rect 143 87 144 88 
<< m1 >>
rect 145 87 146 88 
<< m1 >>
rect 152 87 153 88 
<< m1 >>
rect 154 87 155 88 
<< pdiffusion >>
rect 156 87 157 88 
<< pdiffusion >>
rect 157 87 158 88 
<< pdiffusion >>
rect 158 87 159 88 
<< pdiffusion >>
rect 159 87 160 88 
<< pdiffusion >>
rect 160 87 161 88 
<< pdiffusion >>
rect 161 87 162 88 
<< m1 >>
rect 163 87 164 88 
<< m1 >>
rect 165 87 166 88 
<< m2 >>
rect 171 87 172 88 
<< m1 >>
rect 172 87 173 88 
<< pdiffusion >>
rect 174 87 175 88 
<< pdiffusion >>
rect 175 87 176 88 
<< pdiffusion >>
rect 176 87 177 88 
<< pdiffusion >>
rect 177 87 178 88 
<< pdiffusion >>
rect 178 87 179 88 
<< pdiffusion >>
rect 179 87 180 88 
<< m1 >>
rect 186 87 187 88 
<< m2 >>
rect 189 87 190 88 
<< m1 >>
rect 190 87 191 88 
<< pdiffusion >>
rect 192 87 193 88 
<< pdiffusion >>
rect 193 87 194 88 
<< pdiffusion >>
rect 194 87 195 88 
<< pdiffusion >>
rect 195 87 196 88 
<< pdiffusion >>
rect 196 87 197 88 
<< pdiffusion >>
rect 197 87 198 88 
<< m1 >>
rect 200 87 201 88 
<< m2 >>
rect 201 87 202 88 
<< pdiffusion >>
rect 210 87 211 88 
<< pdiffusion >>
rect 211 87 212 88 
<< pdiffusion >>
rect 212 87 213 88 
<< pdiffusion >>
rect 213 87 214 88 
<< pdiffusion >>
rect 214 87 215 88 
<< pdiffusion >>
rect 215 87 216 88 
<< m1 >>
rect 217 87 218 88 
<< m2 >>
rect 218 87 219 88 
<< pdiffusion >>
rect 228 87 229 88 
<< pdiffusion >>
rect 229 87 230 88 
<< pdiffusion >>
rect 230 87 231 88 
<< pdiffusion >>
rect 231 87 232 88 
<< pdiffusion >>
rect 232 87 233 88 
<< pdiffusion >>
rect 233 87 234 88 
<< m2 >>
rect 243 87 244 88 
<< m1 >>
rect 244 87 245 88 
<< pdiffusion >>
rect 246 87 247 88 
<< pdiffusion >>
rect 247 87 248 88 
<< pdiffusion >>
rect 248 87 249 88 
<< pdiffusion >>
rect 249 87 250 88 
<< pdiffusion >>
rect 250 87 251 88 
<< pdiffusion >>
rect 251 87 252 88 
<< m1 >>
rect 253 87 254 88 
<< m2 >>
rect 254 87 255 88 
<< m1 >>
rect 256 87 257 88 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< m1 >>
rect 19 88 20 89 
<< m1 >>
rect 28 88 29 89 
<< pdiffusion >>
rect 30 88 31 89 
<< pdiffusion >>
rect 31 88 32 89 
<< pdiffusion >>
rect 32 88 33 89 
<< pdiffusion >>
rect 33 88 34 89 
<< pdiffusion >>
rect 34 88 35 89 
<< pdiffusion >>
rect 35 88 36 89 
<< m1 >>
rect 37 88 38 89 
<< m1 >>
rect 40 88 41 89 
<< m1 >>
rect 44 88 45 89 
<< m1 >>
rect 46 88 47 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< m1 >>
rect 55 88 56 89 
<< m1 >>
rect 64 88 65 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< m1 >>
rect 73 88 74 89 
<< m2 >>
rect 74 88 75 89 
<< m1 >>
rect 77 88 78 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 102 88 103 89 
<< m1 >>
rect 104 88 105 89 
<< m1 >>
rect 109 88 110 89 
<< pdiffusion >>
rect 120 88 121 89 
<< pdiffusion >>
rect 121 88 122 89 
<< pdiffusion >>
rect 122 88 123 89 
<< pdiffusion >>
rect 123 88 124 89 
<< pdiffusion >>
rect 124 88 125 89 
<< pdiffusion >>
rect 125 88 126 89 
<< m1 >>
rect 136 88 137 89 
<< pdiffusion >>
rect 138 88 139 89 
<< pdiffusion >>
rect 139 88 140 89 
<< pdiffusion >>
rect 140 88 141 89 
<< pdiffusion >>
rect 141 88 142 89 
<< pdiffusion >>
rect 142 88 143 89 
<< pdiffusion >>
rect 143 88 144 89 
<< m1 >>
rect 145 88 146 89 
<< m1 >>
rect 152 88 153 89 
<< m1 >>
rect 154 88 155 89 
<< pdiffusion >>
rect 156 88 157 89 
<< pdiffusion >>
rect 157 88 158 89 
<< pdiffusion >>
rect 158 88 159 89 
<< pdiffusion >>
rect 159 88 160 89 
<< pdiffusion >>
rect 160 88 161 89 
<< pdiffusion >>
rect 161 88 162 89 
<< m1 >>
rect 163 88 164 89 
<< m1 >>
rect 165 88 166 89 
<< m2 >>
rect 171 88 172 89 
<< m1 >>
rect 172 88 173 89 
<< pdiffusion >>
rect 174 88 175 89 
<< pdiffusion >>
rect 175 88 176 89 
<< pdiffusion >>
rect 176 88 177 89 
<< pdiffusion >>
rect 177 88 178 89 
<< pdiffusion >>
rect 178 88 179 89 
<< pdiffusion >>
rect 179 88 180 89 
<< m1 >>
rect 186 88 187 89 
<< m2 >>
rect 189 88 190 89 
<< m1 >>
rect 190 88 191 89 
<< pdiffusion >>
rect 192 88 193 89 
<< pdiffusion >>
rect 193 88 194 89 
<< pdiffusion >>
rect 194 88 195 89 
<< pdiffusion >>
rect 195 88 196 89 
<< pdiffusion >>
rect 196 88 197 89 
<< pdiffusion >>
rect 197 88 198 89 
<< m1 >>
rect 200 88 201 89 
<< m2 >>
rect 201 88 202 89 
<< pdiffusion >>
rect 210 88 211 89 
<< pdiffusion >>
rect 211 88 212 89 
<< pdiffusion >>
rect 212 88 213 89 
<< pdiffusion >>
rect 213 88 214 89 
<< pdiffusion >>
rect 214 88 215 89 
<< pdiffusion >>
rect 215 88 216 89 
<< m1 >>
rect 217 88 218 89 
<< m2 >>
rect 218 88 219 89 
<< pdiffusion >>
rect 228 88 229 89 
<< pdiffusion >>
rect 229 88 230 89 
<< pdiffusion >>
rect 230 88 231 89 
<< pdiffusion >>
rect 231 88 232 89 
<< pdiffusion >>
rect 232 88 233 89 
<< pdiffusion >>
rect 233 88 234 89 
<< m2 >>
rect 243 88 244 89 
<< m1 >>
rect 244 88 245 89 
<< pdiffusion >>
rect 246 88 247 89 
<< pdiffusion >>
rect 247 88 248 89 
<< pdiffusion >>
rect 248 88 249 89 
<< pdiffusion >>
rect 249 88 250 89 
<< pdiffusion >>
rect 250 88 251 89 
<< pdiffusion >>
rect 251 88 252 89 
<< m1 >>
rect 253 88 254 89 
<< m2 >>
rect 254 88 255 89 
<< m1 >>
rect 256 88 257 89 
<< pdiffusion >>
rect 12 89 13 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< m1 >>
rect 19 89 20 90 
<< m1 >>
rect 28 89 29 90 
<< pdiffusion >>
rect 30 89 31 90 
<< pdiffusion >>
rect 31 89 32 90 
<< pdiffusion >>
rect 32 89 33 90 
<< pdiffusion >>
rect 33 89 34 90 
<< pdiffusion >>
rect 34 89 35 90 
<< pdiffusion >>
rect 35 89 36 90 
<< m1 >>
rect 37 89 38 90 
<< m1 >>
rect 40 89 41 90 
<< m1 >>
rect 44 89 45 90 
<< m1 >>
rect 46 89 47 90 
<< pdiffusion >>
rect 48 89 49 90 
<< m1 >>
rect 49 89 50 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< m1 >>
rect 55 89 56 90 
<< m1 >>
rect 64 89 65 90 
<< pdiffusion >>
rect 66 89 67 90 
<< m1 >>
rect 67 89 68 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< m1 >>
rect 73 89 74 90 
<< m2 >>
rect 74 89 75 90 
<< m1 >>
rect 77 89 78 90 
<< pdiffusion >>
rect 84 89 85 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 102 89 103 90 
<< m1 >>
rect 104 89 105 90 
<< m1 >>
rect 109 89 110 90 
<< pdiffusion >>
rect 120 89 121 90 
<< m1 >>
rect 121 89 122 90 
<< pdiffusion >>
rect 121 89 122 90 
<< pdiffusion >>
rect 122 89 123 90 
<< pdiffusion >>
rect 123 89 124 90 
<< m1 >>
rect 124 89 125 90 
<< pdiffusion >>
rect 124 89 125 90 
<< pdiffusion >>
rect 125 89 126 90 
<< m1 >>
rect 136 89 137 90 
<< pdiffusion >>
rect 138 89 139 90 
<< m1 >>
rect 139 89 140 90 
<< pdiffusion >>
rect 139 89 140 90 
<< pdiffusion >>
rect 140 89 141 90 
<< pdiffusion >>
rect 141 89 142 90 
<< m1 >>
rect 142 89 143 90 
<< pdiffusion >>
rect 142 89 143 90 
<< pdiffusion >>
rect 143 89 144 90 
<< m1 >>
rect 145 89 146 90 
<< m2 >>
rect 145 89 146 90 
<< m2c >>
rect 145 89 146 90 
<< m1 >>
rect 145 89 146 90 
<< m2 >>
rect 145 89 146 90 
<< m1 >>
rect 152 89 153 90 
<< m1 >>
rect 154 89 155 90 
<< pdiffusion >>
rect 156 89 157 90 
<< pdiffusion >>
rect 157 89 158 90 
<< pdiffusion >>
rect 158 89 159 90 
<< pdiffusion >>
rect 159 89 160 90 
<< pdiffusion >>
rect 160 89 161 90 
<< pdiffusion >>
rect 161 89 162 90 
<< m1 >>
rect 163 89 164 90 
<< m1 >>
rect 165 89 166 90 
<< m2 >>
rect 171 89 172 90 
<< m1 >>
rect 172 89 173 90 
<< pdiffusion >>
rect 174 89 175 90 
<< m1 >>
rect 175 89 176 90 
<< pdiffusion >>
rect 175 89 176 90 
<< pdiffusion >>
rect 176 89 177 90 
<< pdiffusion >>
rect 177 89 178 90 
<< m1 >>
rect 178 89 179 90 
<< pdiffusion >>
rect 178 89 179 90 
<< pdiffusion >>
rect 179 89 180 90 
<< m1 >>
rect 186 89 187 90 
<< m2 >>
rect 189 89 190 90 
<< m1 >>
rect 190 89 191 90 
<< pdiffusion >>
rect 192 89 193 90 
<< pdiffusion >>
rect 193 89 194 90 
<< pdiffusion >>
rect 194 89 195 90 
<< pdiffusion >>
rect 195 89 196 90 
<< pdiffusion >>
rect 196 89 197 90 
<< pdiffusion >>
rect 197 89 198 90 
<< m1 >>
rect 200 89 201 90 
<< m2 >>
rect 201 89 202 90 
<< pdiffusion >>
rect 210 89 211 90 
<< pdiffusion >>
rect 211 89 212 90 
<< pdiffusion >>
rect 212 89 213 90 
<< pdiffusion >>
rect 213 89 214 90 
<< m1 >>
rect 214 89 215 90 
<< pdiffusion >>
rect 214 89 215 90 
<< pdiffusion >>
rect 215 89 216 90 
<< m1 >>
rect 217 89 218 90 
<< m2 >>
rect 218 89 219 90 
<< pdiffusion >>
rect 228 89 229 90 
<< pdiffusion >>
rect 229 89 230 90 
<< pdiffusion >>
rect 230 89 231 90 
<< pdiffusion >>
rect 231 89 232 90 
<< pdiffusion >>
rect 232 89 233 90 
<< pdiffusion >>
rect 233 89 234 90 
<< m2 >>
rect 243 89 244 90 
<< m1 >>
rect 244 89 245 90 
<< pdiffusion >>
rect 246 89 247 90 
<< m1 >>
rect 247 89 248 90 
<< pdiffusion >>
rect 247 89 248 90 
<< pdiffusion >>
rect 248 89 249 90 
<< pdiffusion >>
rect 249 89 250 90 
<< pdiffusion >>
rect 250 89 251 90 
<< pdiffusion >>
rect 251 89 252 90 
<< m1 >>
rect 253 89 254 90 
<< m2 >>
rect 254 89 255 90 
<< m1 >>
rect 256 89 257 90 
<< m1 >>
rect 19 90 20 91 
<< m1 >>
rect 28 90 29 91 
<< m1 >>
rect 37 90 38 91 
<< m1 >>
rect 40 90 41 91 
<< m1 >>
rect 44 90 45 91 
<< m1 >>
rect 46 90 47 91 
<< m1 >>
rect 49 90 50 91 
<< m1 >>
rect 55 90 56 91 
<< m1 >>
rect 64 90 65 91 
<< m1 >>
rect 67 90 68 91 
<< m1 >>
rect 73 90 74 91 
<< m2 >>
rect 74 90 75 91 
<< m1 >>
rect 77 90 78 91 
<< m1 >>
rect 102 90 103 91 
<< m1 >>
rect 104 90 105 91 
<< m1 >>
rect 109 90 110 91 
<< m1 >>
rect 121 90 122 91 
<< m1 >>
rect 124 90 125 91 
<< m1 >>
rect 136 90 137 91 
<< m1 >>
rect 139 90 140 91 
<< m1 >>
rect 142 90 143 91 
<< m2 >>
rect 145 90 146 91 
<< m1 >>
rect 152 90 153 91 
<< m1 >>
rect 154 90 155 91 
<< m1 >>
rect 163 90 164 91 
<< m1 >>
rect 165 90 166 91 
<< m2 >>
rect 171 90 172 91 
<< m1 >>
rect 172 90 173 91 
<< m1 >>
rect 175 90 176 91 
<< m1 >>
rect 178 90 179 91 
<< m1 >>
rect 186 90 187 91 
<< m2 >>
rect 189 90 190 91 
<< m1 >>
rect 190 90 191 91 
<< m1 >>
rect 200 90 201 91 
<< m2 >>
rect 201 90 202 91 
<< m1 >>
rect 214 90 215 91 
<< m1 >>
rect 217 90 218 91 
<< m2 >>
rect 218 90 219 91 
<< m2 >>
rect 243 90 244 91 
<< m1 >>
rect 244 90 245 91 
<< m1 >>
rect 247 90 248 91 
<< m1 >>
rect 253 90 254 91 
<< m2 >>
rect 254 90 255 91 
<< m1 >>
rect 256 90 257 91 
<< m1 >>
rect 19 91 20 92 
<< m1 >>
rect 28 91 29 92 
<< m1 >>
rect 37 91 38 92 
<< m1 >>
rect 40 91 41 92 
<< m1 >>
rect 44 91 45 92 
<< m1 >>
rect 46 91 47 92 
<< m1 >>
rect 47 91 48 92 
<< m1 >>
rect 48 91 49 92 
<< m1 >>
rect 49 91 50 92 
<< m1 >>
rect 55 91 56 92 
<< m1 >>
rect 64 91 65 92 
<< m1 >>
rect 67 91 68 92 
<< m1 >>
rect 73 91 74 92 
<< m2 >>
rect 74 91 75 92 
<< m1 >>
rect 77 91 78 92 
<< m2 >>
rect 77 91 78 92 
<< m2c >>
rect 77 91 78 92 
<< m1 >>
rect 77 91 78 92 
<< m2 >>
rect 77 91 78 92 
<< m1 >>
rect 102 91 103 92 
<< m1 >>
rect 104 91 105 92 
<< m1 >>
rect 105 91 106 92 
<< m1 >>
rect 106 91 107 92 
<< m1 >>
rect 107 91 108 92 
<< m2 >>
rect 107 91 108 92 
<< m2c >>
rect 107 91 108 92 
<< m1 >>
rect 107 91 108 92 
<< m2 >>
rect 107 91 108 92 
<< m2 >>
rect 108 91 109 92 
<< m1 >>
rect 109 91 110 92 
<< m2 >>
rect 109 91 110 92 
<< m2 >>
rect 110 91 111 92 
<< m1 >>
rect 111 91 112 92 
<< m2 >>
rect 111 91 112 92 
<< m2c >>
rect 111 91 112 92 
<< m1 >>
rect 111 91 112 92 
<< m2 >>
rect 111 91 112 92 
<< m1 >>
rect 112 91 113 92 
<< m1 >>
rect 113 91 114 92 
<< m1 >>
rect 114 91 115 92 
<< m1 >>
rect 115 91 116 92 
<< m1 >>
rect 116 91 117 92 
<< m1 >>
rect 117 91 118 92 
<< m1 >>
rect 118 91 119 92 
<< m1 >>
rect 119 91 120 92 
<< m1 >>
rect 120 91 121 92 
<< m1 >>
rect 121 91 122 92 
<< m1 >>
rect 124 91 125 92 
<< m1 >>
rect 136 91 137 92 
<< m1 >>
rect 137 91 138 92 
<< m1 >>
rect 138 91 139 92 
<< m1 >>
rect 139 91 140 92 
<< m1 >>
rect 142 91 143 92 
<< m1 >>
rect 143 91 144 92 
<< m1 >>
rect 144 91 145 92 
<< m1 >>
rect 145 91 146 92 
<< m2 >>
rect 145 91 146 92 
<< m1 >>
rect 146 91 147 92 
<< m2 >>
rect 146 91 147 92 
<< m1 >>
rect 147 91 148 92 
<< m2 >>
rect 147 91 148 92 
<< m1 >>
rect 148 91 149 92 
<< m2 >>
rect 148 91 149 92 
<< m1 >>
rect 149 91 150 92 
<< m2 >>
rect 149 91 150 92 
<< m1 >>
rect 150 91 151 92 
<< m2 >>
rect 150 91 151 92 
<< m1 >>
rect 151 91 152 92 
<< m2 >>
rect 151 91 152 92 
<< m1 >>
rect 152 91 153 92 
<< m2 >>
rect 152 91 153 92 
<< m2 >>
rect 153 91 154 92 
<< m1 >>
rect 154 91 155 92 
<< m2 >>
rect 154 91 155 92 
<< m2 >>
rect 155 91 156 92 
<< m1 >>
rect 156 91 157 92 
<< m2 >>
rect 156 91 157 92 
<< m2c >>
rect 156 91 157 92 
<< m1 >>
rect 156 91 157 92 
<< m2 >>
rect 156 91 157 92 
<< m1 >>
rect 163 91 164 92 
<< m1 >>
rect 165 91 166 92 
<< m2 >>
rect 171 91 172 92 
<< m1 >>
rect 172 91 173 92 
<< m1 >>
rect 175 91 176 92 
<< m1 >>
rect 178 91 179 92 
<< m1 >>
rect 186 91 187 92 
<< m2 >>
rect 189 91 190 92 
<< m1 >>
rect 190 91 191 92 
<< m2 >>
rect 190 91 191 92 
<< m2 >>
rect 191 91 192 92 
<< m1 >>
rect 192 91 193 92 
<< m2 >>
rect 192 91 193 92 
<< m2c >>
rect 192 91 193 92 
<< m1 >>
rect 192 91 193 92 
<< m2 >>
rect 192 91 193 92 
<< m1 >>
rect 198 91 199 92 
<< m2 >>
rect 198 91 199 92 
<< m2c >>
rect 198 91 199 92 
<< m1 >>
rect 198 91 199 92 
<< m2 >>
rect 198 91 199 92 
<< m2 >>
rect 199 91 200 92 
<< m1 >>
rect 200 91 201 92 
<< m2 >>
rect 200 91 201 92 
<< m2 >>
rect 201 91 202 92 
<< m1 >>
rect 214 91 215 92 
<< m1 >>
rect 217 91 218 92 
<< m2 >>
rect 218 91 219 92 
<< m2 >>
rect 243 91 244 92 
<< m1 >>
rect 244 91 245 92 
<< m2 >>
rect 244 91 245 92 
<< m2 >>
rect 245 91 246 92 
<< m1 >>
rect 246 91 247 92 
<< m2 >>
rect 246 91 247 92 
<< m2c >>
rect 246 91 247 92 
<< m1 >>
rect 246 91 247 92 
<< m2 >>
rect 246 91 247 92 
<< m1 >>
rect 247 91 248 92 
<< m1 >>
rect 253 91 254 92 
<< m2 >>
rect 254 91 255 92 
<< m1 >>
rect 256 91 257 92 
<< m1 >>
rect 19 92 20 93 
<< m1 >>
rect 28 92 29 93 
<< m1 >>
rect 37 92 38 93 
<< m1 >>
rect 40 92 41 93 
<< m1 >>
rect 44 92 45 93 
<< m1 >>
rect 55 92 56 93 
<< m1 >>
rect 64 92 65 93 
<< m1 >>
rect 67 92 68 93 
<< m1 >>
rect 73 92 74 93 
<< m2 >>
rect 74 92 75 93 
<< m2 >>
rect 77 92 78 93 
<< m1 >>
rect 102 92 103 93 
<< m1 >>
rect 109 92 110 93 
<< m1 >>
rect 124 92 125 93 
<< m1 >>
rect 154 92 155 93 
<< m1 >>
rect 156 92 157 93 
<< m1 >>
rect 163 92 164 93 
<< m1 >>
rect 165 92 166 93 
<< m2 >>
rect 171 92 172 93 
<< m1 >>
rect 172 92 173 93 
<< m1 >>
rect 175 92 176 93 
<< m1 >>
rect 178 92 179 93 
<< m1 >>
rect 186 92 187 93 
<< m1 >>
rect 190 92 191 93 
<< m1 >>
rect 192 92 193 93 
<< m1 >>
rect 196 92 197 93 
<< m2 >>
rect 196 92 197 93 
<< m2c >>
rect 196 92 197 93 
<< m1 >>
rect 196 92 197 93 
<< m2 >>
rect 196 92 197 93 
<< m1 >>
rect 197 92 198 93 
<< m1 >>
rect 198 92 199 93 
<< m1 >>
rect 200 92 201 93 
<< m1 >>
rect 214 92 215 93 
<< m1 >>
rect 217 92 218 93 
<< m2 >>
rect 218 92 219 93 
<< m1 >>
rect 244 92 245 93 
<< m1 >>
rect 253 92 254 93 
<< m2 >>
rect 254 92 255 93 
<< m1 >>
rect 256 92 257 93 
<< m1 >>
rect 19 93 20 94 
<< m1 >>
rect 28 93 29 94 
<< m1 >>
rect 37 93 38 94 
<< m1 >>
rect 40 93 41 94 
<< m1 >>
rect 44 93 45 94 
<< m1 >>
rect 55 93 56 94 
<< m1 >>
rect 64 93 65 94 
<< m1 >>
rect 67 93 68 94 
<< m1 >>
rect 73 93 74 94 
<< m2 >>
rect 74 93 75 94 
<< m1 >>
rect 75 93 76 94 
<< m2 >>
rect 75 93 76 94 
<< m2c >>
rect 75 93 76 94 
<< m1 >>
rect 75 93 76 94 
<< m2 >>
rect 75 93 76 94 
<< m1 >>
rect 76 93 77 94 
<< m1 >>
rect 77 93 78 94 
<< m2 >>
rect 77 93 78 94 
<< m1 >>
rect 78 93 79 94 
<< m1 >>
rect 79 93 80 94 
<< m1 >>
rect 80 93 81 94 
<< m1 >>
rect 81 93 82 94 
<< m1 >>
rect 82 93 83 94 
<< m1 >>
rect 83 93 84 94 
<< m1 >>
rect 84 93 85 94 
<< m2 >>
rect 84 93 85 94 
<< m2c >>
rect 84 93 85 94 
<< m1 >>
rect 84 93 85 94 
<< m2 >>
rect 84 93 85 94 
<< m1 >>
rect 102 93 103 94 
<< m1 >>
rect 103 93 104 94 
<< m2 >>
rect 103 93 104 94 
<< m2c >>
rect 103 93 104 94 
<< m1 >>
rect 103 93 104 94 
<< m2 >>
rect 103 93 104 94 
<< m1 >>
rect 109 93 110 94 
<< m1 >>
rect 124 93 125 94 
<< m1 >>
rect 154 93 155 94 
<< m1 >>
rect 156 93 157 94 
<< m1 >>
rect 158 93 159 94 
<< m1 >>
rect 159 93 160 94 
<< m1 >>
rect 160 93 161 94 
<< m1 >>
rect 161 93 162 94 
<< m2 >>
rect 161 93 162 94 
<< m2c >>
rect 161 93 162 94 
<< m1 >>
rect 161 93 162 94 
<< m2 >>
rect 161 93 162 94 
<< m2 >>
rect 162 93 163 94 
<< m1 >>
rect 163 93 164 94 
<< m2 >>
rect 163 93 164 94 
<< m2 >>
rect 164 93 165 94 
<< m1 >>
rect 165 93 166 94 
<< m2 >>
rect 165 93 166 94 
<< m2 >>
rect 166 93 167 94 
<< m1 >>
rect 167 93 168 94 
<< m2 >>
rect 167 93 168 94 
<< m2c >>
rect 167 93 168 94 
<< m1 >>
rect 167 93 168 94 
<< m2 >>
rect 167 93 168 94 
<< m2 >>
rect 171 93 172 94 
<< m1 >>
rect 172 93 173 94 
<< m1 >>
rect 175 93 176 94 
<< m1 >>
rect 178 93 179 94 
<< m1 >>
rect 186 93 187 94 
<< m1 >>
rect 190 93 191 94 
<< m1 >>
rect 192 93 193 94 
<< m2 >>
rect 196 93 197 94 
<< m1 >>
rect 200 93 201 94 
<< m1 >>
rect 214 93 215 94 
<< m1 >>
rect 217 93 218 94 
<< m2 >>
rect 218 93 219 94 
<< m1 >>
rect 244 93 245 94 
<< m1 >>
rect 253 93 254 94 
<< m2 >>
rect 254 93 255 94 
<< m1 >>
rect 256 93 257 94 
<< m1 >>
rect 19 94 20 95 
<< m1 >>
rect 28 94 29 95 
<< m1 >>
rect 37 94 38 95 
<< m1 >>
rect 40 94 41 95 
<< m1 >>
rect 44 94 45 95 
<< m1 >>
rect 55 94 56 95 
<< m1 >>
rect 64 94 65 95 
<< m1 >>
rect 67 94 68 95 
<< m1 >>
rect 73 94 74 95 
<< m2 >>
rect 77 94 78 95 
<< m2 >>
rect 84 94 85 95 
<< m2 >>
rect 103 94 104 95 
<< m1 >>
rect 109 94 110 95 
<< m1 >>
rect 118 94 119 95 
<< m1 >>
rect 119 94 120 95 
<< m1 >>
rect 120 94 121 95 
<< m1 >>
rect 121 94 122 95 
<< m1 >>
rect 122 94 123 95 
<< m1 >>
rect 123 94 124 95 
<< m1 >>
rect 124 94 125 95 
<< m1 >>
rect 154 94 155 95 
<< m1 >>
rect 156 94 157 95 
<< m1 >>
rect 157 94 158 95 
<< m1 >>
rect 158 94 159 95 
<< m1 >>
rect 163 94 164 95 
<< m1 >>
rect 165 94 166 95 
<< m1 >>
rect 167 94 168 95 
<< m2 >>
rect 171 94 172 95 
<< m1 >>
rect 172 94 173 95 
<< m2 >>
rect 172 94 173 95 
<< m2 >>
rect 173 94 174 95 
<< m2 >>
rect 174 94 175 95 
<< m1 >>
rect 175 94 176 95 
<< m2 >>
rect 175 94 176 95 
<< m2 >>
rect 176 94 177 95 
<< m2 >>
rect 177 94 178 95 
<< m1 >>
rect 178 94 179 95 
<< m2 >>
rect 178 94 179 95 
<< m2 >>
rect 179 94 180 95 
<< m1 >>
rect 180 94 181 95 
<< m2 >>
rect 180 94 181 95 
<< m2c >>
rect 180 94 181 95 
<< m1 >>
rect 180 94 181 95 
<< m2 >>
rect 180 94 181 95 
<< m1 >>
rect 181 94 182 95 
<< m1 >>
rect 186 94 187 95 
<< m1 >>
rect 190 94 191 95 
<< m1 >>
rect 192 94 193 95 
<< m1 >>
rect 193 94 194 95 
<< m1 >>
rect 194 94 195 95 
<< m1 >>
rect 195 94 196 95 
<< m1 >>
rect 196 94 197 95 
<< m2 >>
rect 196 94 197 95 
<< m1 >>
rect 197 94 198 95 
<< m1 >>
rect 198 94 199 95 
<< m2 >>
rect 198 94 199 95 
<< m2c >>
rect 198 94 199 95 
<< m1 >>
rect 198 94 199 95 
<< m2 >>
rect 198 94 199 95 
<< m2 >>
rect 199 94 200 95 
<< m1 >>
rect 200 94 201 95 
<< m2 >>
rect 200 94 201 95 
<< m1 >>
rect 201 94 202 95 
<< m2 >>
rect 201 94 202 95 
<< m1 >>
rect 202 94 203 95 
<< m2 >>
rect 202 94 203 95 
<< m1 >>
rect 203 94 204 95 
<< m2 >>
rect 203 94 204 95 
<< m1 >>
rect 204 94 205 95 
<< m2 >>
rect 204 94 205 95 
<< m1 >>
rect 205 94 206 95 
<< m2 >>
rect 205 94 206 95 
<< m1 >>
rect 206 94 207 95 
<< m2 >>
rect 206 94 207 95 
<< m1 >>
rect 207 94 208 95 
<< m2 >>
rect 207 94 208 95 
<< m1 >>
rect 208 94 209 95 
<< m2 >>
rect 208 94 209 95 
<< m1 >>
rect 209 94 210 95 
<< m2 >>
rect 209 94 210 95 
<< m1 >>
rect 210 94 211 95 
<< m2 >>
rect 210 94 211 95 
<< m1 >>
rect 211 94 212 95 
<< m2 >>
rect 211 94 212 95 
<< m1 >>
rect 212 94 213 95 
<< m2 >>
rect 212 94 213 95 
<< m1 >>
rect 213 94 214 95 
<< m2 >>
rect 213 94 214 95 
<< m1 >>
rect 214 94 215 95 
<< m2 >>
rect 214 94 215 95 
<< m2 >>
rect 215 94 216 95 
<< m1 >>
rect 216 94 217 95 
<< m2 >>
rect 216 94 217 95 
<< m2c >>
rect 216 94 217 95 
<< m1 >>
rect 216 94 217 95 
<< m2 >>
rect 216 94 217 95 
<< m1 >>
rect 217 94 218 95 
<< m2 >>
rect 218 94 219 95 
<< m1 >>
rect 244 94 245 95 
<< m1 >>
rect 253 94 254 95 
<< m2 >>
rect 254 94 255 95 
<< m1 >>
rect 256 94 257 95 
<< m1 >>
rect 19 95 20 96 
<< m1 >>
rect 28 95 29 96 
<< m1 >>
rect 37 95 38 96 
<< m1 >>
rect 40 95 41 96 
<< m1 >>
rect 44 95 45 96 
<< m1 >>
rect 55 95 56 96 
<< m2 >>
rect 63 95 64 96 
<< m1 >>
rect 64 95 65 96 
<< m2 >>
rect 64 95 65 96 
<< m2 >>
rect 65 95 66 96 
<< m1 >>
rect 66 95 67 96 
<< m2 >>
rect 66 95 67 96 
<< m2c >>
rect 66 95 67 96 
<< m1 >>
rect 66 95 67 96 
<< m2 >>
rect 66 95 67 96 
<< m1 >>
rect 67 95 68 96 
<< m1 >>
rect 73 95 74 96 
<< m1 >>
rect 77 95 78 96 
<< m2 >>
rect 77 95 78 96 
<< m2c >>
rect 77 95 78 96 
<< m1 >>
rect 77 95 78 96 
<< m2 >>
rect 77 95 78 96 
<< m1 >>
rect 82 95 83 96 
<< m2 >>
rect 82 95 83 96 
<< m2c >>
rect 82 95 83 96 
<< m1 >>
rect 82 95 83 96 
<< m2 >>
rect 82 95 83 96 
<< m1 >>
rect 83 95 84 96 
<< m1 >>
rect 84 95 85 96 
<< m2 >>
rect 84 95 85 96 
<< m1 >>
rect 85 95 86 96 
<< m1 >>
rect 86 95 87 96 
<< m1 >>
rect 87 95 88 96 
<< m1 >>
rect 88 95 89 96 
<< m1 >>
rect 89 95 90 96 
<< m1 >>
rect 90 95 91 96 
<< m1 >>
rect 91 95 92 96 
<< m1 >>
rect 92 95 93 96 
<< m1 >>
rect 93 95 94 96 
<< m1 >>
rect 94 95 95 96 
<< m1 >>
rect 95 95 96 96 
<< m1 >>
rect 96 95 97 96 
<< m1 >>
rect 97 95 98 96 
<< m1 >>
rect 98 95 99 96 
<< m1 >>
rect 99 95 100 96 
<< m1 >>
rect 100 95 101 96 
<< m1 >>
rect 101 95 102 96 
<< m1 >>
rect 102 95 103 96 
<< m1 >>
rect 103 95 104 96 
<< m2 >>
rect 103 95 104 96 
<< m1 >>
rect 104 95 105 96 
<< m1 >>
rect 105 95 106 96 
<< m1 >>
rect 106 95 107 96 
<< m1 >>
rect 107 95 108 96 
<< m2 >>
rect 107 95 108 96 
<< m2c >>
rect 107 95 108 96 
<< m1 >>
rect 107 95 108 96 
<< m2 >>
rect 107 95 108 96 
<< m2 >>
rect 108 95 109 96 
<< m1 >>
rect 109 95 110 96 
<< m2 >>
rect 109 95 110 96 
<< m2 >>
rect 110 95 111 96 
<< m1 >>
rect 111 95 112 96 
<< m2 >>
rect 111 95 112 96 
<< m2c >>
rect 111 95 112 96 
<< m1 >>
rect 111 95 112 96 
<< m2 >>
rect 111 95 112 96 
<< m1 >>
rect 112 95 113 96 
<< m1 >>
rect 113 95 114 96 
<< m1 >>
rect 114 95 115 96 
<< m1 >>
rect 115 95 116 96 
<< m1 >>
rect 116 95 117 96 
<< m2 >>
rect 116 95 117 96 
<< m2c >>
rect 116 95 117 96 
<< m1 >>
rect 116 95 117 96 
<< m2 >>
rect 116 95 117 96 
<< m2 >>
rect 117 95 118 96 
<< m1 >>
rect 118 95 119 96 
<< m2 >>
rect 118 95 119 96 
<< m2 >>
rect 119 95 120 96 
<< m2 >>
rect 120 95 121 96 
<< m2 >>
rect 121 95 122 96 
<< m2 >>
rect 122 95 123 96 
<< m1 >>
rect 154 95 155 96 
<< m1 >>
rect 163 95 164 96 
<< m2 >>
rect 163 95 164 96 
<< m2c >>
rect 163 95 164 96 
<< m1 >>
rect 163 95 164 96 
<< m2 >>
rect 163 95 164 96 
<< m1 >>
rect 165 95 166 96 
<< m2 >>
rect 165 95 166 96 
<< m2c >>
rect 165 95 166 96 
<< m1 >>
rect 165 95 166 96 
<< m2 >>
rect 165 95 166 96 
<< m1 >>
rect 167 95 168 96 
<< m2 >>
rect 167 95 168 96 
<< m2c >>
rect 167 95 168 96 
<< m1 >>
rect 167 95 168 96 
<< m2 >>
rect 167 95 168 96 
<< m1 >>
rect 172 95 173 96 
<< m1 >>
rect 175 95 176 96 
<< m1 >>
rect 178 95 179 96 
<< m1 >>
rect 181 95 182 96 
<< m1 >>
rect 186 95 187 96 
<< m1 >>
rect 190 95 191 96 
<< m2 >>
rect 196 95 197 96 
<< m2 >>
rect 218 95 219 96 
<< m1 >>
rect 244 95 245 96 
<< m1 >>
rect 253 95 254 96 
<< m2 >>
rect 254 95 255 96 
<< m1 >>
rect 256 95 257 96 
<< m1 >>
rect 19 96 20 97 
<< m1 >>
rect 28 96 29 97 
<< m1 >>
rect 37 96 38 97 
<< m1 >>
rect 40 96 41 97 
<< m1 >>
rect 44 96 45 97 
<< m1 >>
rect 55 96 56 97 
<< m2 >>
rect 63 96 64 97 
<< m1 >>
rect 64 96 65 97 
<< m1 >>
rect 73 96 74 97 
<< m2 >>
rect 77 96 78 97 
<< m2 >>
rect 82 96 83 97 
<< m2 >>
rect 84 96 85 97 
<< m2 >>
rect 103 96 104 97 
<< m1 >>
rect 109 96 110 97 
<< m1 >>
rect 118 96 119 97 
<< m2 >>
rect 122 96 123 97 
<< m1 >>
rect 154 96 155 97 
<< m2 >>
rect 163 96 164 97 
<< m2 >>
rect 165 96 166 97 
<< m2 >>
rect 167 96 168 97 
<< m1 >>
rect 172 96 173 97 
<< m1 >>
rect 175 96 176 97 
<< m1 >>
rect 178 96 179 97 
<< m1 >>
rect 181 96 182 97 
<< m1 >>
rect 186 96 187 97 
<< m1 >>
rect 190 96 191 97 
<< m1 >>
rect 196 96 197 97 
<< m2 >>
rect 196 96 197 97 
<< m2c >>
rect 196 96 197 97 
<< m1 >>
rect 196 96 197 97 
<< m2 >>
rect 196 96 197 97 
<< m1 >>
rect 197 96 198 97 
<< m1 >>
rect 198 96 199 97 
<< m1 >>
rect 199 96 200 97 
<< m1 >>
rect 200 96 201 97 
<< m1 >>
rect 201 96 202 97 
<< m1 >>
rect 218 96 219 97 
<< m2 >>
rect 218 96 219 97 
<< m2c >>
rect 218 96 219 97 
<< m1 >>
rect 218 96 219 97 
<< m2 >>
rect 218 96 219 97 
<< m1 >>
rect 244 96 245 97 
<< m1 >>
rect 253 96 254 97 
<< m2 >>
rect 254 96 255 97 
<< m1 >>
rect 256 96 257 97 
<< m1 >>
rect 19 97 20 98 
<< m1 >>
rect 28 97 29 98 
<< m1 >>
rect 34 97 35 98 
<< m2 >>
rect 34 97 35 98 
<< m2c >>
rect 34 97 35 98 
<< m1 >>
rect 34 97 35 98 
<< m2 >>
rect 34 97 35 98 
<< m1 >>
rect 35 97 36 98 
<< m1 >>
rect 36 97 37 98 
<< m1 >>
rect 37 97 38 98 
<< m1 >>
rect 40 97 41 98 
<< m1 >>
rect 44 97 45 98 
<< m1 >>
rect 46 97 47 98 
<< m1 >>
rect 47 97 48 98 
<< m1 >>
rect 48 97 49 98 
<< m1 >>
rect 49 97 50 98 
<< m1 >>
rect 50 97 51 98 
<< m1 >>
rect 51 97 52 98 
<< m1 >>
rect 52 97 53 98 
<< m1 >>
rect 53 97 54 98 
<< m2 >>
rect 53 97 54 98 
<< m2c >>
rect 53 97 54 98 
<< m1 >>
rect 53 97 54 98 
<< m2 >>
rect 53 97 54 98 
<< m2 >>
rect 54 97 55 98 
<< m1 >>
rect 55 97 56 98 
<< m2 >>
rect 55 97 56 98 
<< m2 >>
rect 56 97 57 98 
<< m1 >>
rect 57 97 58 98 
<< m2 >>
rect 57 97 58 98 
<< m2c >>
rect 57 97 58 98 
<< m1 >>
rect 57 97 58 98 
<< m2 >>
rect 57 97 58 98 
<< m1 >>
rect 58 97 59 98 
<< m1 >>
rect 59 97 60 98 
<< m1 >>
rect 60 97 61 98 
<< m1 >>
rect 61 97 62 98 
<< m1 >>
rect 62 97 63 98 
<< m2 >>
rect 62 97 63 98 
<< m2c >>
rect 62 97 63 98 
<< m1 >>
rect 62 97 63 98 
<< m2 >>
rect 62 97 63 98 
<< m2 >>
rect 63 97 64 98 
<< m1 >>
rect 64 97 65 98 
<< m1 >>
rect 66 97 67 98 
<< m1 >>
rect 67 97 68 98 
<< m1 >>
rect 68 97 69 98 
<< m1 >>
rect 69 97 70 98 
<< m1 >>
rect 70 97 71 98 
<< m1 >>
rect 71 97 72 98 
<< m2 >>
rect 71 97 72 98 
<< m2c >>
rect 71 97 72 98 
<< m1 >>
rect 71 97 72 98 
<< m2 >>
rect 71 97 72 98 
<< m2 >>
rect 72 97 73 98 
<< m1 >>
rect 73 97 74 98 
<< m2 >>
rect 73 97 74 98 
<< m2 >>
rect 74 97 75 98 
<< m1 >>
rect 75 97 76 98 
<< m2 >>
rect 75 97 76 98 
<< m2c >>
rect 75 97 76 98 
<< m1 >>
rect 75 97 76 98 
<< m2 >>
rect 75 97 76 98 
<< m1 >>
rect 76 97 77 98 
<< m1 >>
rect 77 97 78 98 
<< m2 >>
rect 77 97 78 98 
<< m1 >>
rect 78 97 79 98 
<< m1 >>
rect 79 97 80 98 
<< m1 >>
rect 80 97 81 98 
<< m1 >>
rect 81 97 82 98 
<< m1 >>
rect 82 97 83 98 
<< m2 >>
rect 82 97 83 98 
<< m1 >>
rect 83 97 84 98 
<< m1 >>
rect 84 97 85 98 
<< m2 >>
rect 84 97 85 98 
<< m1 >>
rect 85 97 86 98 
<< m2 >>
rect 85 97 86 98 
<< m1 >>
rect 86 97 87 98 
<< m2 >>
rect 86 97 87 98 
<< m1 >>
rect 87 97 88 98 
<< m2 >>
rect 87 97 88 98 
<< m1 >>
rect 88 97 89 98 
<< m2 >>
rect 88 97 89 98 
<< m1 >>
rect 89 97 90 98 
<< m2 >>
rect 89 97 90 98 
<< m1 >>
rect 90 97 91 98 
<< m2 >>
rect 90 97 91 98 
<< m1 >>
rect 91 97 92 98 
<< m2 >>
rect 91 97 92 98 
<< m1 >>
rect 92 97 93 98 
<< m2 >>
rect 92 97 93 98 
<< m1 >>
rect 93 97 94 98 
<< m2 >>
rect 93 97 94 98 
<< m1 >>
rect 94 97 95 98 
<< m2 >>
rect 94 97 95 98 
<< m1 >>
rect 95 97 96 98 
<< m2 >>
rect 95 97 96 98 
<< m1 >>
rect 96 97 97 98 
<< m2 >>
rect 96 97 97 98 
<< m1 >>
rect 97 97 98 98 
<< m2 >>
rect 97 97 98 98 
<< m1 >>
rect 98 97 99 98 
<< m2 >>
rect 98 97 99 98 
<< m1 >>
rect 99 97 100 98 
<< m2 >>
rect 99 97 100 98 
<< m1 >>
rect 100 97 101 98 
<< m2 >>
rect 100 97 101 98 
<< m1 >>
rect 101 97 102 98 
<< m1 >>
rect 102 97 103 98 
<< m1 >>
rect 103 97 104 98 
<< m2 >>
rect 103 97 104 98 
<< m1 >>
rect 104 97 105 98 
<< m1 >>
rect 105 97 106 98 
<< m1 >>
rect 106 97 107 98 
<< m1 >>
rect 107 97 108 98 
<< m2 >>
rect 107 97 108 98 
<< m2c >>
rect 107 97 108 98 
<< m1 >>
rect 107 97 108 98 
<< m2 >>
rect 107 97 108 98 
<< m2 >>
rect 108 97 109 98 
<< m1 >>
rect 109 97 110 98 
<< m2 >>
rect 109 97 110 98 
<< m2 >>
rect 110 97 111 98 
<< m1 >>
rect 111 97 112 98 
<< m2 >>
rect 111 97 112 98 
<< m2c >>
rect 111 97 112 98 
<< m1 >>
rect 111 97 112 98 
<< m2 >>
rect 111 97 112 98 
<< m1 >>
rect 112 97 113 98 
<< m1 >>
rect 113 97 114 98 
<< m1 >>
rect 114 97 115 98 
<< m1 >>
rect 115 97 116 98 
<< m1 >>
rect 116 97 117 98 
<< m2 >>
rect 116 97 117 98 
<< m2c >>
rect 116 97 117 98 
<< m1 >>
rect 116 97 117 98 
<< m2 >>
rect 116 97 117 98 
<< m2 >>
rect 117 97 118 98 
<< m1 >>
rect 118 97 119 98 
<< m2 >>
rect 118 97 119 98 
<< m2 >>
rect 119 97 120 98 
<< m1 >>
rect 120 97 121 98 
<< m2 >>
rect 120 97 121 98 
<< m2c >>
rect 120 97 121 98 
<< m1 >>
rect 120 97 121 98 
<< m2 >>
rect 120 97 121 98 
<< m1 >>
rect 121 97 122 98 
<< m1 >>
rect 122 97 123 98 
<< m2 >>
rect 122 97 123 98 
<< m1 >>
rect 123 97 124 98 
<< m1 >>
rect 124 97 125 98 
<< m1 >>
rect 125 97 126 98 
<< m1 >>
rect 126 97 127 98 
<< m1 >>
rect 127 97 128 98 
<< m1 >>
rect 128 97 129 98 
<< m1 >>
rect 129 97 130 98 
<< m1 >>
rect 130 97 131 98 
<< m1 >>
rect 131 97 132 98 
<< m1 >>
rect 132 97 133 98 
<< m1 >>
rect 133 97 134 98 
<< m1 >>
rect 134 97 135 98 
<< m1 >>
rect 135 97 136 98 
<< m1 >>
rect 136 97 137 98 
<< m1 >>
rect 137 97 138 98 
<< m1 >>
rect 138 97 139 98 
<< m1 >>
rect 139 97 140 98 
<< m1 >>
rect 140 97 141 98 
<< m1 >>
rect 141 97 142 98 
<< m1 >>
rect 142 97 143 98 
<< m1 >>
rect 143 97 144 98 
<< m1 >>
rect 144 97 145 98 
<< m1 >>
rect 145 97 146 98 
<< m1 >>
rect 146 97 147 98 
<< m1 >>
rect 147 97 148 98 
<< m1 >>
rect 148 97 149 98 
<< m1 >>
rect 149 97 150 98 
<< m1 >>
rect 150 97 151 98 
<< m1 >>
rect 151 97 152 98 
<< m1 >>
rect 152 97 153 98 
<< m2 >>
rect 152 97 153 98 
<< m2c >>
rect 152 97 153 98 
<< m1 >>
rect 152 97 153 98 
<< m2 >>
rect 152 97 153 98 
<< m2 >>
rect 153 97 154 98 
<< m1 >>
rect 154 97 155 98 
<< m2 >>
rect 154 97 155 98 
<< m2 >>
rect 155 97 156 98 
<< m1 >>
rect 156 97 157 98 
<< m2 >>
rect 156 97 157 98 
<< m2c >>
rect 156 97 157 98 
<< m1 >>
rect 156 97 157 98 
<< m2 >>
rect 156 97 157 98 
<< m1 >>
rect 157 97 158 98 
<< m1 >>
rect 158 97 159 98 
<< m1 >>
rect 159 97 160 98 
<< m1 >>
rect 160 97 161 98 
<< m1 >>
rect 161 97 162 98 
<< m1 >>
rect 162 97 163 98 
<< m1 >>
rect 163 97 164 98 
<< m2 >>
rect 163 97 164 98 
<< m1 >>
rect 164 97 165 98 
<< m1 >>
rect 165 97 166 98 
<< m2 >>
rect 165 97 166 98 
<< m1 >>
rect 166 97 167 98 
<< m1 >>
rect 167 97 168 98 
<< m2 >>
rect 167 97 168 98 
<< m1 >>
rect 168 97 169 98 
<< m1 >>
rect 169 97 170 98 
<< m1 >>
rect 170 97 171 98 
<< m2 >>
rect 170 97 171 98 
<< m2c >>
rect 170 97 171 98 
<< m1 >>
rect 170 97 171 98 
<< m2 >>
rect 170 97 171 98 
<< m2 >>
rect 171 97 172 98 
<< m1 >>
rect 172 97 173 98 
<< m2 >>
rect 172 97 173 98 
<< m2 >>
rect 173 97 174 98 
<< m1 >>
rect 174 97 175 98 
<< m2 >>
rect 174 97 175 98 
<< m1 >>
rect 175 97 176 98 
<< m2 >>
rect 175 97 176 98 
<< m2 >>
rect 176 97 177 98 
<< m1 >>
rect 177 97 178 98 
<< m2 >>
rect 177 97 178 98 
<< m2c >>
rect 177 97 178 98 
<< m1 >>
rect 177 97 178 98 
<< m2 >>
rect 177 97 178 98 
<< m1 >>
rect 178 97 179 98 
<< m1 >>
rect 181 97 182 98 
<< m1 >>
rect 186 97 187 98 
<< m1 >>
rect 187 97 188 98 
<< m1 >>
rect 188 97 189 98 
<< m2 >>
rect 188 97 189 98 
<< m2c >>
rect 188 97 189 98 
<< m1 >>
rect 188 97 189 98 
<< m2 >>
rect 188 97 189 98 
<< m2 >>
rect 189 97 190 98 
<< m1 >>
rect 190 97 191 98 
<< m2 >>
rect 190 97 191 98 
<< m2 >>
rect 191 97 192 98 
<< m1 >>
rect 192 97 193 98 
<< m2 >>
rect 192 97 193 98 
<< m1 >>
rect 193 97 194 98 
<< m2 >>
rect 193 97 194 98 
<< m1 >>
rect 194 97 195 98 
<< m2 >>
rect 194 97 195 98 
<< m1 >>
rect 201 97 202 98 
<< m1 >>
rect 203 97 204 98 
<< m1 >>
rect 204 97 205 98 
<< m1 >>
rect 205 97 206 98 
<< m1 >>
rect 206 97 207 98 
<< m1 >>
rect 207 97 208 98 
<< m1 >>
rect 208 97 209 98 
<< m1 >>
rect 209 97 210 98 
<< m1 >>
rect 210 97 211 98 
<< m1 >>
rect 211 97 212 98 
<< m1 >>
rect 212 97 213 98 
<< m1 >>
rect 218 97 219 98 
<< m1 >>
rect 244 97 245 98 
<< m1 >>
rect 253 97 254 98 
<< m2 >>
rect 254 97 255 98 
<< m1 >>
rect 256 97 257 98 
<< m1 >>
rect 19 98 20 99 
<< m1 >>
rect 28 98 29 99 
<< m2 >>
rect 34 98 35 99 
<< m1 >>
rect 40 98 41 99 
<< m1 >>
rect 44 98 45 99 
<< m1 >>
rect 46 98 47 99 
<< m1 >>
rect 55 98 56 99 
<< m1 >>
rect 64 98 65 99 
<< m1 >>
rect 66 98 67 99 
<< m1 >>
rect 73 98 74 99 
<< m2 >>
rect 77 98 78 99 
<< m2 >>
rect 82 98 83 99 
<< m2 >>
rect 100 98 101 99 
<< m2 >>
rect 103 98 104 99 
<< m1 >>
rect 109 98 110 99 
<< m1 >>
rect 118 98 119 99 
<< m2 >>
rect 122 98 123 99 
<< m1 >>
rect 154 98 155 99 
<< m2 >>
rect 163 98 164 99 
<< m2 >>
rect 165 98 166 99 
<< m2 >>
rect 167 98 168 99 
<< m1 >>
rect 172 98 173 99 
<< m1 >>
rect 174 98 175 99 
<< m1 >>
rect 181 98 182 99 
<< m1 >>
rect 190 98 191 99 
<< m1 >>
rect 192 98 193 99 
<< m1 >>
rect 194 98 195 99 
<< m2 >>
rect 194 98 195 99 
<< m1 >>
rect 195 98 196 99 
<< m1 >>
rect 196 98 197 99 
<< m1 >>
rect 197 98 198 99 
<< m1 >>
rect 198 98 199 99 
<< m1 >>
rect 199 98 200 99 
<< m2 >>
rect 199 98 200 99 
<< m2c >>
rect 199 98 200 99 
<< m1 >>
rect 199 98 200 99 
<< m2 >>
rect 199 98 200 99 
<< m2 >>
rect 200 98 201 99 
<< m1 >>
rect 201 98 202 99 
<< m2 >>
rect 201 98 202 99 
<< m2 >>
rect 202 98 203 99 
<< m1 >>
rect 203 98 204 99 
<< m2 >>
rect 203 98 204 99 
<< m2c >>
rect 203 98 204 99 
<< m1 >>
rect 203 98 204 99 
<< m2 >>
rect 203 98 204 99 
<< m1 >>
rect 212 98 213 99 
<< m1 >>
rect 213 98 214 99 
<< m1 >>
rect 214 98 215 99 
<< m1 >>
rect 215 98 216 99 
<< m1 >>
rect 216 98 217 99 
<< m2 >>
rect 216 98 217 99 
<< m2c >>
rect 216 98 217 99 
<< m1 >>
rect 216 98 217 99 
<< m2 >>
rect 216 98 217 99 
<< m2 >>
rect 217 98 218 99 
<< m1 >>
rect 218 98 219 99 
<< m2 >>
rect 218 98 219 99 
<< m2 >>
rect 219 98 220 99 
<< m1 >>
rect 220 98 221 99 
<< m2 >>
rect 220 98 221 99 
<< m2c >>
rect 220 98 221 99 
<< m1 >>
rect 220 98 221 99 
<< m2 >>
rect 220 98 221 99 
<< m1 >>
rect 244 98 245 99 
<< m1 >>
rect 253 98 254 99 
<< m2 >>
rect 254 98 255 99 
<< m1 >>
rect 256 98 257 99 
<< m1 >>
rect 19 99 20 100 
<< m1 >>
rect 28 99 29 100 
<< m1 >>
rect 31 99 32 100 
<< m1 >>
rect 32 99 33 100 
<< m1 >>
rect 33 99 34 100 
<< m1 >>
rect 34 99 35 100 
<< m2 >>
rect 34 99 35 100 
<< m1 >>
rect 35 99 36 100 
<< m1 >>
rect 36 99 37 100 
<< m1 >>
rect 37 99 38 100 
<< m1 >>
rect 40 99 41 100 
<< m1 >>
rect 44 99 45 100 
<< m1 >>
rect 46 99 47 100 
<< m1 >>
rect 49 99 50 100 
<< m1 >>
rect 50 99 51 100 
<< m1 >>
rect 51 99 52 100 
<< m1 >>
rect 52 99 53 100 
<< m1 >>
rect 53 99 54 100 
<< m1 >>
rect 55 99 56 100 
<< m1 >>
rect 64 99 65 100 
<< m1 >>
rect 66 99 67 100 
<< m1 >>
rect 73 99 74 100 
<< m1 >>
rect 77 99 78 100 
<< m2 >>
rect 77 99 78 100 
<< m2c >>
rect 77 99 78 100 
<< m1 >>
rect 77 99 78 100 
<< m2 >>
rect 77 99 78 100 
<< m1 >>
rect 82 99 83 100 
<< m2 >>
rect 82 99 83 100 
<< m2c >>
rect 82 99 83 100 
<< m1 >>
rect 82 99 83 100 
<< m2 >>
rect 82 99 83 100 
<< m1 >>
rect 100 99 101 100 
<< m2 >>
rect 100 99 101 100 
<< m2c >>
rect 100 99 101 100 
<< m1 >>
rect 100 99 101 100 
<< m2 >>
rect 100 99 101 100 
<< m1 >>
rect 103 99 104 100 
<< m2 >>
rect 103 99 104 100 
<< m2c >>
rect 103 99 104 100 
<< m1 >>
rect 103 99 104 100 
<< m2 >>
rect 103 99 104 100 
<< m1 >>
rect 109 99 110 100 
<< m1 >>
rect 118 99 119 100 
<< m1 >>
rect 122 99 123 100 
<< m2 >>
rect 122 99 123 100 
<< m2c >>
rect 122 99 123 100 
<< m1 >>
rect 122 99 123 100 
<< m2 >>
rect 122 99 123 100 
<< m1 >>
rect 123 99 124 100 
<< m1 >>
rect 124 99 125 100 
<< m1 >>
rect 125 99 126 100 
<< m1 >>
rect 126 99 127 100 
<< m1 >>
rect 127 99 128 100 
<< m1 >>
rect 128 99 129 100 
<< m1 >>
rect 129 99 130 100 
<< m1 >>
rect 154 99 155 100 
<< m1 >>
rect 163 99 164 100 
<< m2 >>
rect 163 99 164 100 
<< m2c >>
rect 163 99 164 100 
<< m1 >>
rect 163 99 164 100 
<< m2 >>
rect 163 99 164 100 
<< m1 >>
rect 165 99 166 100 
<< m2 >>
rect 165 99 166 100 
<< m2c >>
rect 165 99 166 100 
<< m1 >>
rect 165 99 166 100 
<< m2 >>
rect 165 99 166 100 
<< m1 >>
rect 167 99 168 100 
<< m2 >>
rect 167 99 168 100 
<< m2c >>
rect 167 99 168 100 
<< m1 >>
rect 167 99 168 100 
<< m2 >>
rect 167 99 168 100 
<< m1 >>
rect 172 99 173 100 
<< m1 >>
rect 174 99 175 100 
<< m1 >>
rect 181 99 182 100 
<< m1 >>
rect 190 99 191 100 
<< m1 >>
rect 192 99 193 100 
<< m2 >>
rect 194 99 195 100 
<< m2 >>
rect 195 99 196 100 
<< m2 >>
rect 196 99 197 100 
<< m2 >>
rect 197 99 198 100 
<< m1 >>
rect 201 99 202 100 
<< m1 >>
rect 218 99 219 100 
<< m1 >>
rect 220 99 221 100 
<< m1 >>
rect 244 99 245 100 
<< m1 >>
rect 253 99 254 100 
<< m2 >>
rect 254 99 255 100 
<< m1 >>
rect 256 99 257 100 
<< m1 >>
rect 19 100 20 101 
<< m1 >>
rect 28 100 29 101 
<< m1 >>
rect 31 100 32 101 
<< m2 >>
rect 34 100 35 101 
<< m1 >>
rect 37 100 38 101 
<< m1 >>
rect 40 100 41 101 
<< m1 >>
rect 44 100 45 101 
<< m1 >>
rect 46 100 47 101 
<< m1 >>
rect 49 100 50 101 
<< m1 >>
rect 53 100 54 101 
<< m2 >>
rect 53 100 54 101 
<< m2c >>
rect 53 100 54 101 
<< m1 >>
rect 53 100 54 101 
<< m2 >>
rect 53 100 54 101 
<< m2 >>
rect 54 100 55 101 
<< m1 >>
rect 55 100 56 101 
<< m2 >>
rect 55 100 56 101 
<< m2 >>
rect 56 100 57 101 
<< m2 >>
rect 63 100 64 101 
<< m1 >>
rect 64 100 65 101 
<< m2 >>
rect 64 100 65 101 
<< m2 >>
rect 65 100 66 101 
<< m1 >>
rect 66 100 67 101 
<< m2 >>
rect 66 100 67 101 
<< m2c >>
rect 66 100 67 101 
<< m1 >>
rect 66 100 67 101 
<< m2 >>
rect 66 100 67 101 
<< m1 >>
rect 73 100 74 101 
<< m1 >>
rect 77 100 78 101 
<< m1 >>
rect 82 100 83 101 
<< m1 >>
rect 88 100 89 101 
<< m1 >>
rect 89 100 90 101 
<< m1 >>
rect 90 100 91 101 
<< m1 >>
rect 91 100 92 101 
<< m1 >>
rect 100 100 101 101 
<< m1 >>
rect 103 100 104 101 
<< m1 >>
rect 109 100 110 101 
<< m1 >>
rect 118 100 119 101 
<< m1 >>
rect 129 100 130 101 
<< m1 >>
rect 154 100 155 101 
<< m1 >>
rect 163 100 164 101 
<< m1 >>
rect 165 100 166 101 
<< m1 >>
rect 167 100 168 101 
<< m2 >>
rect 171 100 172 101 
<< m1 >>
rect 172 100 173 101 
<< m2 >>
rect 172 100 173 101 
<< m2 >>
rect 173 100 174 101 
<< m1 >>
rect 174 100 175 101 
<< m2 >>
rect 174 100 175 101 
<< m2c >>
rect 174 100 175 101 
<< m1 >>
rect 174 100 175 101 
<< m2 >>
rect 174 100 175 101 
<< m1 >>
rect 178 100 179 101 
<< m1 >>
rect 179 100 180 101 
<< m2 >>
rect 179 100 180 101 
<< m2c >>
rect 179 100 180 101 
<< m1 >>
rect 179 100 180 101 
<< m2 >>
rect 179 100 180 101 
<< m2 >>
rect 180 100 181 101 
<< m1 >>
rect 181 100 182 101 
<< m2 >>
rect 181 100 182 101 
<< m2 >>
rect 182 100 183 101 
<< m2 >>
rect 189 100 190 101 
<< m1 >>
rect 190 100 191 101 
<< m2 >>
rect 190 100 191 101 
<< m2 >>
rect 191 100 192 101 
<< m1 >>
rect 192 100 193 101 
<< m2 >>
rect 192 100 193 101 
<< m2c >>
rect 192 100 193 101 
<< m1 >>
rect 192 100 193 101 
<< m2 >>
rect 192 100 193 101 
<< m1 >>
rect 196 100 197 101 
<< m1 >>
rect 197 100 198 101 
<< m2 >>
rect 197 100 198 101 
<< m1 >>
rect 198 100 199 101 
<< m2 >>
rect 198 100 199 101 
<< m1 >>
rect 199 100 200 101 
<< m2 >>
rect 199 100 200 101 
<< m2 >>
rect 200 100 201 101 
<< m1 >>
rect 201 100 202 101 
<< m2 >>
rect 201 100 202 101 
<< m2 >>
rect 202 100 203 101 
<< m1 >>
rect 203 100 204 101 
<< m2 >>
rect 203 100 204 101 
<< m2c >>
rect 203 100 204 101 
<< m1 >>
rect 203 100 204 101 
<< m2 >>
rect 203 100 204 101 
<< m1 >>
rect 204 100 205 101 
<< m1 >>
rect 205 100 206 101 
<< m1 >>
rect 206 100 207 101 
<< m1 >>
rect 207 100 208 101 
<< m1 >>
rect 208 100 209 101 
<< m1 >>
rect 209 100 210 101 
<< m1 >>
rect 210 100 211 101 
<< m1 >>
rect 211 100 212 101 
<< m1 >>
rect 218 100 219 101 
<< m1 >>
rect 220 100 221 101 
<< m1 >>
rect 244 100 245 101 
<< m1 >>
rect 253 100 254 101 
<< m2 >>
rect 254 100 255 101 
<< m1 >>
rect 256 100 257 101 
<< m1 >>
rect 19 101 20 102 
<< m1 >>
rect 28 101 29 102 
<< m1 >>
rect 31 101 32 102 
<< m1 >>
rect 34 101 35 102 
<< m2 >>
rect 34 101 35 102 
<< m1 >>
rect 37 101 38 102 
<< m1 >>
rect 40 101 41 102 
<< m1 >>
rect 44 101 45 102 
<< m1 >>
rect 46 101 47 102 
<< m1 >>
rect 49 101 50 102 
<< m1 >>
rect 55 101 56 102 
<< m2 >>
rect 56 101 57 102 
<< m2 >>
rect 63 101 64 102 
<< m1 >>
rect 64 101 65 102 
<< m1 >>
rect 73 101 74 102 
<< m1 >>
rect 77 101 78 102 
<< m1 >>
rect 82 101 83 102 
<< m1 >>
rect 88 101 89 102 
<< m1 >>
rect 91 101 92 102 
<< m1 >>
rect 100 101 101 102 
<< m1 >>
rect 103 101 104 102 
<< m1 >>
rect 109 101 110 102 
<< m1 >>
rect 118 101 119 102 
<< m1 >>
rect 129 101 130 102 
<< m1 >>
rect 154 101 155 102 
<< m1 >>
rect 163 101 164 102 
<< m1 >>
rect 165 101 166 102 
<< m1 >>
rect 167 101 168 102 
<< m2 >>
rect 171 101 172 102 
<< m1 >>
rect 172 101 173 102 
<< m1 >>
rect 178 101 179 102 
<< m1 >>
rect 181 101 182 102 
<< m2 >>
rect 182 101 183 102 
<< m2 >>
rect 189 101 190 102 
<< m1 >>
rect 190 101 191 102 
<< m1 >>
rect 196 101 197 102 
<< m1 >>
rect 199 101 200 102 
<< m1 >>
rect 201 101 202 102 
<< m1 >>
rect 211 101 212 102 
<< m1 >>
rect 218 101 219 102 
<< m1 >>
rect 220 101 221 102 
<< m1 >>
rect 244 101 245 102 
<< m1 >>
rect 253 101 254 102 
<< m2 >>
rect 254 101 255 102 
<< m1 >>
rect 256 101 257 102 
<< pdiffusion >>
rect 12 102 13 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< m1 >>
rect 19 102 20 103 
<< m1 >>
rect 28 102 29 103 
<< pdiffusion >>
rect 30 102 31 103 
<< m1 >>
rect 31 102 32 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< m1 >>
rect 33 102 34 103 
<< m2 >>
rect 33 102 34 103 
<< m2c >>
rect 33 102 34 103 
<< m1 >>
rect 33 102 34 103 
<< m2 >>
rect 33 102 34 103 
<< pdiffusion >>
rect 33 102 34 103 
<< m1 >>
rect 34 102 35 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< m1 >>
rect 37 102 38 103 
<< m1 >>
rect 40 102 41 103 
<< m1 >>
rect 44 102 45 103 
<< m1 >>
rect 46 102 47 103 
<< pdiffusion >>
rect 48 102 49 103 
<< m1 >>
rect 49 102 50 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m1 >>
rect 55 102 56 103 
<< m2 >>
rect 56 102 57 103 
<< m2 >>
rect 63 102 64 103 
<< m1 >>
rect 64 102 65 103 
<< pdiffusion >>
rect 66 102 67 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< m1 >>
rect 73 102 74 103 
<< m1 >>
rect 77 102 78 103 
<< m1 >>
rect 82 102 83 103 
<< pdiffusion >>
rect 84 102 85 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< m1 >>
rect 88 102 89 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< m1 >>
rect 91 102 92 103 
<< m1 >>
rect 100 102 101 103 
<< pdiffusion >>
rect 102 102 103 103 
<< m1 >>
rect 103 102 104 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< m1 >>
rect 109 102 110 103 
<< m1 >>
rect 118 102 119 103 
<< pdiffusion >>
rect 120 102 121 103 
<< pdiffusion >>
rect 121 102 122 103 
<< pdiffusion >>
rect 122 102 123 103 
<< pdiffusion >>
rect 123 102 124 103 
<< pdiffusion >>
rect 124 102 125 103 
<< pdiffusion >>
rect 125 102 126 103 
<< m1 >>
rect 129 102 130 103 
<< pdiffusion >>
rect 138 102 139 103 
<< pdiffusion >>
rect 139 102 140 103 
<< pdiffusion >>
rect 140 102 141 103 
<< pdiffusion >>
rect 141 102 142 103 
<< pdiffusion >>
rect 142 102 143 103 
<< pdiffusion >>
rect 143 102 144 103 
<< m1 >>
rect 154 102 155 103 
<< pdiffusion >>
rect 156 102 157 103 
<< pdiffusion >>
rect 157 102 158 103 
<< pdiffusion >>
rect 158 102 159 103 
<< pdiffusion >>
rect 159 102 160 103 
<< pdiffusion >>
rect 160 102 161 103 
<< pdiffusion >>
rect 161 102 162 103 
<< m1 >>
rect 163 102 164 103 
<< m1 >>
rect 165 102 166 103 
<< m1 >>
rect 167 102 168 103 
<< m2 >>
rect 171 102 172 103 
<< m1 >>
rect 172 102 173 103 
<< pdiffusion >>
rect 174 102 175 103 
<< pdiffusion >>
rect 175 102 176 103 
<< pdiffusion >>
rect 176 102 177 103 
<< pdiffusion >>
rect 177 102 178 103 
<< m1 >>
rect 178 102 179 103 
<< pdiffusion >>
rect 178 102 179 103 
<< pdiffusion >>
rect 179 102 180 103 
<< m1 >>
rect 181 102 182 103 
<< m2 >>
rect 182 102 183 103 
<< m2 >>
rect 189 102 190 103 
<< m1 >>
rect 190 102 191 103 
<< pdiffusion >>
rect 192 102 193 103 
<< pdiffusion >>
rect 193 102 194 103 
<< pdiffusion >>
rect 194 102 195 103 
<< pdiffusion >>
rect 195 102 196 103 
<< m1 >>
rect 196 102 197 103 
<< pdiffusion >>
rect 196 102 197 103 
<< pdiffusion >>
rect 197 102 198 103 
<< m1 >>
rect 199 102 200 103 
<< m1 >>
rect 201 102 202 103 
<< pdiffusion >>
rect 210 102 211 103 
<< m1 >>
rect 211 102 212 103 
<< pdiffusion >>
rect 211 102 212 103 
<< pdiffusion >>
rect 212 102 213 103 
<< pdiffusion >>
rect 213 102 214 103 
<< pdiffusion >>
rect 214 102 215 103 
<< pdiffusion >>
rect 215 102 216 103 
<< m1 >>
rect 218 102 219 103 
<< m1 >>
rect 220 102 221 103 
<< pdiffusion >>
rect 228 102 229 103 
<< pdiffusion >>
rect 229 102 230 103 
<< pdiffusion >>
rect 230 102 231 103 
<< pdiffusion >>
rect 231 102 232 103 
<< pdiffusion >>
rect 232 102 233 103 
<< pdiffusion >>
rect 233 102 234 103 
<< m1 >>
rect 244 102 245 103 
<< pdiffusion >>
rect 246 102 247 103 
<< pdiffusion >>
rect 247 102 248 103 
<< pdiffusion >>
rect 248 102 249 103 
<< pdiffusion >>
rect 249 102 250 103 
<< pdiffusion >>
rect 250 102 251 103 
<< pdiffusion >>
rect 251 102 252 103 
<< m1 >>
rect 253 102 254 103 
<< m2 >>
rect 254 102 255 103 
<< m1 >>
rect 256 102 257 103 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< m1 >>
rect 19 103 20 104 
<< m1 >>
rect 28 103 29 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< m1 >>
rect 37 103 38 104 
<< m1 >>
rect 40 103 41 104 
<< m1 >>
rect 44 103 45 104 
<< m1 >>
rect 46 103 47 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m1 >>
rect 55 103 56 104 
<< m2 >>
rect 56 103 57 104 
<< m2 >>
rect 63 103 64 104 
<< m1 >>
rect 64 103 65 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< m1 >>
rect 73 103 74 104 
<< m1 >>
rect 77 103 78 104 
<< m1 >>
rect 82 103 83 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< m1 >>
rect 91 103 92 104 
<< m1 >>
rect 100 103 101 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< m1 >>
rect 109 103 110 104 
<< m1 >>
rect 118 103 119 104 
<< pdiffusion >>
rect 120 103 121 104 
<< pdiffusion >>
rect 121 103 122 104 
<< pdiffusion >>
rect 122 103 123 104 
<< pdiffusion >>
rect 123 103 124 104 
<< pdiffusion >>
rect 124 103 125 104 
<< pdiffusion >>
rect 125 103 126 104 
<< m1 >>
rect 129 103 130 104 
<< pdiffusion >>
rect 138 103 139 104 
<< pdiffusion >>
rect 139 103 140 104 
<< pdiffusion >>
rect 140 103 141 104 
<< pdiffusion >>
rect 141 103 142 104 
<< pdiffusion >>
rect 142 103 143 104 
<< pdiffusion >>
rect 143 103 144 104 
<< m1 >>
rect 154 103 155 104 
<< pdiffusion >>
rect 156 103 157 104 
<< pdiffusion >>
rect 157 103 158 104 
<< pdiffusion >>
rect 158 103 159 104 
<< pdiffusion >>
rect 159 103 160 104 
<< pdiffusion >>
rect 160 103 161 104 
<< pdiffusion >>
rect 161 103 162 104 
<< m1 >>
rect 163 103 164 104 
<< m1 >>
rect 165 103 166 104 
<< m1 >>
rect 167 103 168 104 
<< m2 >>
rect 171 103 172 104 
<< m1 >>
rect 172 103 173 104 
<< pdiffusion >>
rect 174 103 175 104 
<< pdiffusion >>
rect 175 103 176 104 
<< pdiffusion >>
rect 176 103 177 104 
<< pdiffusion >>
rect 177 103 178 104 
<< pdiffusion >>
rect 178 103 179 104 
<< pdiffusion >>
rect 179 103 180 104 
<< m1 >>
rect 181 103 182 104 
<< m2 >>
rect 182 103 183 104 
<< m2 >>
rect 189 103 190 104 
<< m1 >>
rect 190 103 191 104 
<< pdiffusion >>
rect 192 103 193 104 
<< pdiffusion >>
rect 193 103 194 104 
<< pdiffusion >>
rect 194 103 195 104 
<< pdiffusion >>
rect 195 103 196 104 
<< pdiffusion >>
rect 196 103 197 104 
<< pdiffusion >>
rect 197 103 198 104 
<< m1 >>
rect 199 103 200 104 
<< m1 >>
rect 201 103 202 104 
<< pdiffusion >>
rect 210 103 211 104 
<< pdiffusion >>
rect 211 103 212 104 
<< pdiffusion >>
rect 212 103 213 104 
<< pdiffusion >>
rect 213 103 214 104 
<< pdiffusion >>
rect 214 103 215 104 
<< pdiffusion >>
rect 215 103 216 104 
<< m1 >>
rect 218 103 219 104 
<< m1 >>
rect 220 103 221 104 
<< pdiffusion >>
rect 228 103 229 104 
<< pdiffusion >>
rect 229 103 230 104 
<< pdiffusion >>
rect 230 103 231 104 
<< pdiffusion >>
rect 231 103 232 104 
<< pdiffusion >>
rect 232 103 233 104 
<< pdiffusion >>
rect 233 103 234 104 
<< m1 >>
rect 244 103 245 104 
<< pdiffusion >>
rect 246 103 247 104 
<< pdiffusion >>
rect 247 103 248 104 
<< pdiffusion >>
rect 248 103 249 104 
<< pdiffusion >>
rect 249 103 250 104 
<< pdiffusion >>
rect 250 103 251 104 
<< pdiffusion >>
rect 251 103 252 104 
<< m1 >>
rect 253 103 254 104 
<< m2 >>
rect 254 103 255 104 
<< m1 >>
rect 256 103 257 104 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< m1 >>
rect 19 104 20 105 
<< m1 >>
rect 28 104 29 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< m1 >>
rect 37 104 38 105 
<< m1 >>
rect 40 104 41 105 
<< m1 >>
rect 44 104 45 105 
<< m1 >>
rect 46 104 47 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m1 >>
rect 55 104 56 105 
<< m2 >>
rect 56 104 57 105 
<< m2 >>
rect 63 104 64 105 
<< m1 >>
rect 64 104 65 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< m1 >>
rect 73 104 74 105 
<< m1 >>
rect 77 104 78 105 
<< m1 >>
rect 82 104 83 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< m1 >>
rect 91 104 92 105 
<< m1 >>
rect 100 104 101 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< m1 >>
rect 109 104 110 105 
<< m1 >>
rect 118 104 119 105 
<< pdiffusion >>
rect 120 104 121 105 
<< pdiffusion >>
rect 121 104 122 105 
<< pdiffusion >>
rect 122 104 123 105 
<< pdiffusion >>
rect 123 104 124 105 
<< pdiffusion >>
rect 124 104 125 105 
<< pdiffusion >>
rect 125 104 126 105 
<< m1 >>
rect 129 104 130 105 
<< pdiffusion >>
rect 138 104 139 105 
<< pdiffusion >>
rect 139 104 140 105 
<< pdiffusion >>
rect 140 104 141 105 
<< pdiffusion >>
rect 141 104 142 105 
<< pdiffusion >>
rect 142 104 143 105 
<< pdiffusion >>
rect 143 104 144 105 
<< m1 >>
rect 154 104 155 105 
<< pdiffusion >>
rect 156 104 157 105 
<< pdiffusion >>
rect 157 104 158 105 
<< pdiffusion >>
rect 158 104 159 105 
<< pdiffusion >>
rect 159 104 160 105 
<< pdiffusion >>
rect 160 104 161 105 
<< pdiffusion >>
rect 161 104 162 105 
<< m1 >>
rect 163 104 164 105 
<< m1 >>
rect 165 104 166 105 
<< m1 >>
rect 167 104 168 105 
<< m2 >>
rect 171 104 172 105 
<< m1 >>
rect 172 104 173 105 
<< pdiffusion >>
rect 174 104 175 105 
<< pdiffusion >>
rect 175 104 176 105 
<< pdiffusion >>
rect 176 104 177 105 
<< pdiffusion >>
rect 177 104 178 105 
<< pdiffusion >>
rect 178 104 179 105 
<< pdiffusion >>
rect 179 104 180 105 
<< m1 >>
rect 181 104 182 105 
<< m2 >>
rect 182 104 183 105 
<< m2 >>
rect 189 104 190 105 
<< m1 >>
rect 190 104 191 105 
<< pdiffusion >>
rect 192 104 193 105 
<< pdiffusion >>
rect 193 104 194 105 
<< pdiffusion >>
rect 194 104 195 105 
<< pdiffusion >>
rect 195 104 196 105 
<< pdiffusion >>
rect 196 104 197 105 
<< pdiffusion >>
rect 197 104 198 105 
<< m1 >>
rect 199 104 200 105 
<< m1 >>
rect 201 104 202 105 
<< pdiffusion >>
rect 210 104 211 105 
<< pdiffusion >>
rect 211 104 212 105 
<< pdiffusion >>
rect 212 104 213 105 
<< pdiffusion >>
rect 213 104 214 105 
<< pdiffusion >>
rect 214 104 215 105 
<< pdiffusion >>
rect 215 104 216 105 
<< m1 >>
rect 218 104 219 105 
<< m1 >>
rect 220 104 221 105 
<< pdiffusion >>
rect 228 104 229 105 
<< pdiffusion >>
rect 229 104 230 105 
<< pdiffusion >>
rect 230 104 231 105 
<< pdiffusion >>
rect 231 104 232 105 
<< pdiffusion >>
rect 232 104 233 105 
<< pdiffusion >>
rect 233 104 234 105 
<< m1 >>
rect 244 104 245 105 
<< pdiffusion >>
rect 246 104 247 105 
<< pdiffusion >>
rect 247 104 248 105 
<< pdiffusion >>
rect 248 104 249 105 
<< pdiffusion >>
rect 249 104 250 105 
<< pdiffusion >>
rect 250 104 251 105 
<< pdiffusion >>
rect 251 104 252 105 
<< m1 >>
rect 253 104 254 105 
<< m2 >>
rect 254 104 255 105 
<< m1 >>
rect 256 104 257 105 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< m1 >>
rect 19 105 20 106 
<< m1 >>
rect 28 105 29 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< m1 >>
rect 37 105 38 106 
<< m1 >>
rect 40 105 41 106 
<< m1 >>
rect 44 105 45 106 
<< m1 >>
rect 46 105 47 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m1 >>
rect 55 105 56 106 
<< m2 >>
rect 56 105 57 106 
<< m2 >>
rect 63 105 64 106 
<< m1 >>
rect 64 105 65 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< m1 >>
rect 73 105 74 106 
<< m1 >>
rect 77 105 78 106 
<< m1 >>
rect 82 105 83 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< m1 >>
rect 91 105 92 106 
<< m1 >>
rect 100 105 101 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< m1 >>
rect 109 105 110 106 
<< m1 >>
rect 118 105 119 106 
<< pdiffusion >>
rect 120 105 121 106 
<< pdiffusion >>
rect 121 105 122 106 
<< pdiffusion >>
rect 122 105 123 106 
<< pdiffusion >>
rect 123 105 124 106 
<< pdiffusion >>
rect 124 105 125 106 
<< pdiffusion >>
rect 125 105 126 106 
<< m1 >>
rect 129 105 130 106 
<< pdiffusion >>
rect 138 105 139 106 
<< pdiffusion >>
rect 139 105 140 106 
<< pdiffusion >>
rect 140 105 141 106 
<< pdiffusion >>
rect 141 105 142 106 
<< pdiffusion >>
rect 142 105 143 106 
<< pdiffusion >>
rect 143 105 144 106 
<< m1 >>
rect 154 105 155 106 
<< pdiffusion >>
rect 156 105 157 106 
<< pdiffusion >>
rect 157 105 158 106 
<< pdiffusion >>
rect 158 105 159 106 
<< pdiffusion >>
rect 159 105 160 106 
<< pdiffusion >>
rect 160 105 161 106 
<< pdiffusion >>
rect 161 105 162 106 
<< m1 >>
rect 163 105 164 106 
<< m1 >>
rect 165 105 166 106 
<< m1 >>
rect 167 105 168 106 
<< m2 >>
rect 171 105 172 106 
<< m1 >>
rect 172 105 173 106 
<< pdiffusion >>
rect 174 105 175 106 
<< pdiffusion >>
rect 175 105 176 106 
<< pdiffusion >>
rect 176 105 177 106 
<< pdiffusion >>
rect 177 105 178 106 
<< pdiffusion >>
rect 178 105 179 106 
<< pdiffusion >>
rect 179 105 180 106 
<< m1 >>
rect 181 105 182 106 
<< m2 >>
rect 182 105 183 106 
<< m2 >>
rect 189 105 190 106 
<< m1 >>
rect 190 105 191 106 
<< pdiffusion >>
rect 192 105 193 106 
<< pdiffusion >>
rect 193 105 194 106 
<< pdiffusion >>
rect 194 105 195 106 
<< pdiffusion >>
rect 195 105 196 106 
<< pdiffusion >>
rect 196 105 197 106 
<< pdiffusion >>
rect 197 105 198 106 
<< m1 >>
rect 199 105 200 106 
<< m1 >>
rect 201 105 202 106 
<< pdiffusion >>
rect 210 105 211 106 
<< pdiffusion >>
rect 211 105 212 106 
<< pdiffusion >>
rect 212 105 213 106 
<< pdiffusion >>
rect 213 105 214 106 
<< pdiffusion >>
rect 214 105 215 106 
<< pdiffusion >>
rect 215 105 216 106 
<< m1 >>
rect 218 105 219 106 
<< m1 >>
rect 220 105 221 106 
<< pdiffusion >>
rect 228 105 229 106 
<< pdiffusion >>
rect 229 105 230 106 
<< pdiffusion >>
rect 230 105 231 106 
<< pdiffusion >>
rect 231 105 232 106 
<< pdiffusion >>
rect 232 105 233 106 
<< pdiffusion >>
rect 233 105 234 106 
<< m1 >>
rect 244 105 245 106 
<< pdiffusion >>
rect 246 105 247 106 
<< pdiffusion >>
rect 247 105 248 106 
<< pdiffusion >>
rect 248 105 249 106 
<< pdiffusion >>
rect 249 105 250 106 
<< pdiffusion >>
rect 250 105 251 106 
<< pdiffusion >>
rect 251 105 252 106 
<< m1 >>
rect 253 105 254 106 
<< m2 >>
rect 254 105 255 106 
<< m1 >>
rect 256 105 257 106 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< m1 >>
rect 19 106 20 107 
<< m1 >>
rect 28 106 29 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< m1 >>
rect 37 106 38 107 
<< m1 >>
rect 40 106 41 107 
<< m1 >>
rect 44 106 45 107 
<< m1 >>
rect 46 106 47 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m1 >>
rect 55 106 56 107 
<< m2 >>
rect 56 106 57 107 
<< m2 >>
rect 63 106 64 107 
<< m1 >>
rect 64 106 65 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< m1 >>
rect 73 106 74 107 
<< m1 >>
rect 77 106 78 107 
<< m1 >>
rect 82 106 83 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< m1 >>
rect 91 106 92 107 
<< m1 >>
rect 100 106 101 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< m1 >>
rect 109 106 110 107 
<< m1 >>
rect 118 106 119 107 
<< pdiffusion >>
rect 120 106 121 107 
<< pdiffusion >>
rect 121 106 122 107 
<< pdiffusion >>
rect 122 106 123 107 
<< pdiffusion >>
rect 123 106 124 107 
<< pdiffusion >>
rect 124 106 125 107 
<< pdiffusion >>
rect 125 106 126 107 
<< m1 >>
rect 129 106 130 107 
<< pdiffusion >>
rect 138 106 139 107 
<< pdiffusion >>
rect 139 106 140 107 
<< pdiffusion >>
rect 140 106 141 107 
<< pdiffusion >>
rect 141 106 142 107 
<< pdiffusion >>
rect 142 106 143 107 
<< pdiffusion >>
rect 143 106 144 107 
<< m1 >>
rect 154 106 155 107 
<< pdiffusion >>
rect 156 106 157 107 
<< pdiffusion >>
rect 157 106 158 107 
<< pdiffusion >>
rect 158 106 159 107 
<< pdiffusion >>
rect 159 106 160 107 
<< pdiffusion >>
rect 160 106 161 107 
<< pdiffusion >>
rect 161 106 162 107 
<< m1 >>
rect 163 106 164 107 
<< m1 >>
rect 165 106 166 107 
<< m1 >>
rect 167 106 168 107 
<< m2 >>
rect 171 106 172 107 
<< m1 >>
rect 172 106 173 107 
<< pdiffusion >>
rect 174 106 175 107 
<< pdiffusion >>
rect 175 106 176 107 
<< pdiffusion >>
rect 176 106 177 107 
<< pdiffusion >>
rect 177 106 178 107 
<< pdiffusion >>
rect 178 106 179 107 
<< pdiffusion >>
rect 179 106 180 107 
<< m1 >>
rect 181 106 182 107 
<< m2 >>
rect 182 106 183 107 
<< m2 >>
rect 189 106 190 107 
<< m1 >>
rect 190 106 191 107 
<< pdiffusion >>
rect 192 106 193 107 
<< pdiffusion >>
rect 193 106 194 107 
<< pdiffusion >>
rect 194 106 195 107 
<< pdiffusion >>
rect 195 106 196 107 
<< pdiffusion >>
rect 196 106 197 107 
<< pdiffusion >>
rect 197 106 198 107 
<< m1 >>
rect 199 106 200 107 
<< m1 >>
rect 201 106 202 107 
<< pdiffusion >>
rect 210 106 211 107 
<< pdiffusion >>
rect 211 106 212 107 
<< pdiffusion >>
rect 212 106 213 107 
<< pdiffusion >>
rect 213 106 214 107 
<< pdiffusion >>
rect 214 106 215 107 
<< pdiffusion >>
rect 215 106 216 107 
<< m1 >>
rect 218 106 219 107 
<< m1 >>
rect 220 106 221 107 
<< pdiffusion >>
rect 228 106 229 107 
<< pdiffusion >>
rect 229 106 230 107 
<< pdiffusion >>
rect 230 106 231 107 
<< pdiffusion >>
rect 231 106 232 107 
<< pdiffusion >>
rect 232 106 233 107 
<< pdiffusion >>
rect 233 106 234 107 
<< m1 >>
rect 244 106 245 107 
<< pdiffusion >>
rect 246 106 247 107 
<< pdiffusion >>
rect 247 106 248 107 
<< pdiffusion >>
rect 248 106 249 107 
<< pdiffusion >>
rect 249 106 250 107 
<< pdiffusion >>
rect 250 106 251 107 
<< pdiffusion >>
rect 251 106 252 107 
<< m1 >>
rect 253 106 254 107 
<< m2 >>
rect 254 106 255 107 
<< m1 >>
rect 256 106 257 107 
<< pdiffusion >>
rect 12 107 13 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< m1 >>
rect 19 107 20 108 
<< m1 >>
rect 28 107 29 108 
<< pdiffusion >>
rect 30 107 31 108 
<< m1 >>
rect 31 107 32 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< m1 >>
rect 37 107 38 108 
<< m1 >>
rect 40 107 41 108 
<< m1 >>
rect 44 107 45 108 
<< m1 >>
rect 46 107 47 108 
<< pdiffusion >>
rect 48 107 49 108 
<< m1 >>
rect 49 107 50 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m1 >>
rect 55 107 56 108 
<< m2 >>
rect 56 107 57 108 
<< m1 >>
rect 59 107 60 108 
<< m1 >>
rect 60 107 61 108 
<< m1 >>
rect 61 107 62 108 
<< m1 >>
rect 62 107 63 108 
<< m2 >>
rect 62 107 63 108 
<< m2c >>
rect 62 107 63 108 
<< m1 >>
rect 62 107 63 108 
<< m2 >>
rect 62 107 63 108 
<< m2 >>
rect 63 107 64 108 
<< m1 >>
rect 64 107 65 108 
<< pdiffusion >>
rect 66 107 67 108 
<< m1 >>
rect 67 107 68 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< m1 >>
rect 73 107 74 108 
<< m1 >>
rect 77 107 78 108 
<< m1 >>
rect 82 107 83 108 
<< pdiffusion >>
rect 84 107 85 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< m1 >>
rect 91 107 92 108 
<< m1 >>
rect 100 107 101 108 
<< pdiffusion >>
rect 102 107 103 108 
<< m1 >>
rect 103 107 104 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< m1 >>
rect 109 107 110 108 
<< m1 >>
rect 118 107 119 108 
<< pdiffusion >>
rect 120 107 121 108 
<< pdiffusion >>
rect 121 107 122 108 
<< pdiffusion >>
rect 122 107 123 108 
<< pdiffusion >>
rect 123 107 124 108 
<< m1 >>
rect 124 107 125 108 
<< pdiffusion >>
rect 124 107 125 108 
<< pdiffusion >>
rect 125 107 126 108 
<< m1 >>
rect 129 107 130 108 
<< pdiffusion >>
rect 138 107 139 108 
<< pdiffusion >>
rect 139 107 140 108 
<< pdiffusion >>
rect 140 107 141 108 
<< pdiffusion >>
rect 141 107 142 108 
<< pdiffusion >>
rect 142 107 143 108 
<< pdiffusion >>
rect 143 107 144 108 
<< m1 >>
rect 154 107 155 108 
<< pdiffusion >>
rect 156 107 157 108 
<< pdiffusion >>
rect 157 107 158 108 
<< pdiffusion >>
rect 158 107 159 108 
<< pdiffusion >>
rect 159 107 160 108 
<< pdiffusion >>
rect 160 107 161 108 
<< pdiffusion >>
rect 161 107 162 108 
<< m1 >>
rect 163 107 164 108 
<< m1 >>
rect 165 107 166 108 
<< m1 >>
rect 167 107 168 108 
<< m2 >>
rect 171 107 172 108 
<< m1 >>
rect 172 107 173 108 
<< pdiffusion >>
rect 174 107 175 108 
<< pdiffusion >>
rect 175 107 176 108 
<< pdiffusion >>
rect 176 107 177 108 
<< pdiffusion >>
rect 177 107 178 108 
<< pdiffusion >>
rect 178 107 179 108 
<< pdiffusion >>
rect 179 107 180 108 
<< m1 >>
rect 181 107 182 108 
<< m2 >>
rect 182 107 183 108 
<< m2 >>
rect 189 107 190 108 
<< m1 >>
rect 190 107 191 108 
<< pdiffusion >>
rect 192 107 193 108 
<< pdiffusion >>
rect 193 107 194 108 
<< pdiffusion >>
rect 194 107 195 108 
<< pdiffusion >>
rect 195 107 196 108 
<< pdiffusion >>
rect 196 107 197 108 
<< pdiffusion >>
rect 197 107 198 108 
<< m1 >>
rect 199 107 200 108 
<< m1 >>
rect 201 107 202 108 
<< pdiffusion >>
rect 210 107 211 108 
<< pdiffusion >>
rect 211 107 212 108 
<< pdiffusion >>
rect 212 107 213 108 
<< pdiffusion >>
rect 213 107 214 108 
<< pdiffusion >>
rect 214 107 215 108 
<< pdiffusion >>
rect 215 107 216 108 
<< m1 >>
rect 218 107 219 108 
<< m1 >>
rect 220 107 221 108 
<< pdiffusion >>
rect 228 107 229 108 
<< pdiffusion >>
rect 229 107 230 108 
<< pdiffusion >>
rect 230 107 231 108 
<< pdiffusion >>
rect 231 107 232 108 
<< pdiffusion >>
rect 232 107 233 108 
<< pdiffusion >>
rect 233 107 234 108 
<< m1 >>
rect 244 107 245 108 
<< pdiffusion >>
rect 246 107 247 108 
<< m1 >>
rect 247 107 248 108 
<< pdiffusion >>
rect 247 107 248 108 
<< pdiffusion >>
rect 248 107 249 108 
<< pdiffusion >>
rect 249 107 250 108 
<< pdiffusion >>
rect 250 107 251 108 
<< pdiffusion >>
rect 251 107 252 108 
<< m1 >>
rect 253 107 254 108 
<< m2 >>
rect 254 107 255 108 
<< m1 >>
rect 256 107 257 108 
<< m1 >>
rect 19 108 20 109 
<< m1 >>
rect 28 108 29 109 
<< m1 >>
rect 31 108 32 109 
<< m1 >>
rect 37 108 38 109 
<< m2 >>
rect 37 108 38 109 
<< m2c >>
rect 37 108 38 109 
<< m1 >>
rect 37 108 38 109 
<< m2 >>
rect 37 108 38 109 
<< m1 >>
rect 40 108 41 109 
<< m2 >>
rect 40 108 41 109 
<< m2c >>
rect 40 108 41 109 
<< m1 >>
rect 40 108 41 109 
<< m2 >>
rect 40 108 41 109 
<< m1 >>
rect 44 108 45 109 
<< m1 >>
rect 46 108 47 109 
<< m1 >>
rect 49 108 50 109 
<< m1 >>
rect 55 108 56 109 
<< m2 >>
rect 56 108 57 109 
<< m1 >>
rect 59 108 60 109 
<< m1 >>
rect 64 108 65 109 
<< m1 >>
rect 67 108 68 109 
<< m1 >>
rect 73 108 74 109 
<< m1 >>
rect 77 108 78 109 
<< m1 >>
rect 82 108 83 109 
<< m1 >>
rect 91 108 92 109 
<< m1 >>
rect 100 108 101 109 
<< m1 >>
rect 103 108 104 109 
<< m1 >>
rect 109 108 110 109 
<< m1 >>
rect 118 108 119 109 
<< m1 >>
rect 124 108 125 109 
<< m1 >>
rect 129 108 130 109 
<< m1 >>
rect 154 108 155 109 
<< m1 >>
rect 163 108 164 109 
<< m1 >>
rect 165 108 166 109 
<< m1 >>
rect 167 108 168 109 
<< m2 >>
rect 171 108 172 109 
<< m1 >>
rect 172 108 173 109 
<< m1 >>
rect 181 108 182 109 
<< m2 >>
rect 182 108 183 109 
<< m2 >>
rect 189 108 190 109 
<< m1 >>
rect 190 108 191 109 
<< m1 >>
rect 199 108 200 109 
<< m1 >>
rect 201 108 202 109 
<< m1 >>
rect 218 108 219 109 
<< m1 >>
rect 220 108 221 109 
<< m1 >>
rect 244 108 245 109 
<< m1 >>
rect 247 108 248 109 
<< m1 >>
rect 253 108 254 109 
<< m2 >>
rect 254 108 255 109 
<< m1 >>
rect 256 108 257 109 
<< m1 >>
rect 19 109 20 110 
<< m1 >>
rect 28 109 29 110 
<< m1 >>
rect 31 109 32 110 
<< m2 >>
rect 37 109 38 110 
<< m2 >>
rect 40 109 41 110 
<< m1 >>
rect 44 109 45 110 
<< m1 >>
rect 46 109 47 110 
<< m1 >>
rect 49 109 50 110 
<< m1 >>
rect 55 109 56 110 
<< m2 >>
rect 56 109 57 110 
<< m1 >>
rect 59 109 60 110 
<< m2 >>
rect 59 109 60 110 
<< m2c >>
rect 59 109 60 110 
<< m1 >>
rect 59 109 60 110 
<< m2 >>
rect 59 109 60 110 
<< m1 >>
rect 64 109 65 110 
<< m2 >>
rect 64 109 65 110 
<< m2c >>
rect 64 109 65 110 
<< m1 >>
rect 64 109 65 110 
<< m2 >>
rect 64 109 65 110 
<< m1 >>
rect 67 109 68 110 
<< m1 >>
rect 73 109 74 110 
<< m1 >>
rect 77 109 78 110 
<< m1 >>
rect 82 109 83 110 
<< m1 >>
rect 91 109 92 110 
<< m1 >>
rect 100 109 101 110 
<< m1 >>
rect 103 109 104 110 
<< m1 >>
rect 109 109 110 110 
<< m1 >>
rect 118 109 119 110 
<< m1 >>
rect 124 109 125 110 
<< m1 >>
rect 126 109 127 110 
<< m1 >>
rect 127 109 128 110 
<< m2 >>
rect 127 109 128 110 
<< m2c >>
rect 127 109 128 110 
<< m1 >>
rect 127 109 128 110 
<< m2 >>
rect 127 109 128 110 
<< m2 >>
rect 128 109 129 110 
<< m1 >>
rect 129 109 130 110 
<< m2 >>
rect 129 109 130 110 
<< m2 >>
rect 130 109 131 110 
<< m1 >>
rect 131 109 132 110 
<< m2 >>
rect 131 109 132 110 
<< m2c >>
rect 131 109 132 110 
<< m1 >>
rect 131 109 132 110 
<< m2 >>
rect 131 109 132 110 
<< m1 >>
rect 154 109 155 110 
<< m1 >>
rect 163 109 164 110 
<< m1 >>
rect 165 109 166 110 
<< m1 >>
rect 167 109 168 110 
<< m2 >>
rect 171 109 172 110 
<< m1 >>
rect 172 109 173 110 
<< m1 >>
rect 181 109 182 110 
<< m2 >>
rect 182 109 183 110 
<< m1 >>
rect 185 109 186 110 
<< m2 >>
rect 185 109 186 110 
<< m2c >>
rect 185 109 186 110 
<< m1 >>
rect 185 109 186 110 
<< m2 >>
rect 185 109 186 110 
<< m1 >>
rect 186 109 187 110 
<< m1 >>
rect 187 109 188 110 
<< m1 >>
rect 188 109 189 110 
<< m2 >>
rect 188 109 189 110 
<< m2c >>
rect 188 109 189 110 
<< m1 >>
rect 188 109 189 110 
<< m2 >>
rect 188 109 189 110 
<< m2 >>
rect 189 109 190 110 
<< m1 >>
rect 190 109 191 110 
<< m1 >>
rect 199 109 200 110 
<< m1 >>
rect 201 109 202 110 
<< m1 >>
rect 218 109 219 110 
<< m1 >>
rect 220 109 221 110 
<< m1 >>
rect 244 109 245 110 
<< m1 >>
rect 247 109 248 110 
<< m1 >>
rect 253 109 254 110 
<< m2 >>
rect 254 109 255 110 
<< m1 >>
rect 256 109 257 110 
<< m1 >>
rect 19 110 20 111 
<< m1 >>
rect 28 110 29 111 
<< m1 >>
rect 31 110 32 111 
<< m1 >>
rect 32 110 33 111 
<< m1 >>
rect 33 110 34 111 
<< m1 >>
rect 34 110 35 111 
<< m1 >>
rect 35 110 36 111 
<< m1 >>
rect 36 110 37 111 
<< m1 >>
rect 37 110 38 111 
<< m2 >>
rect 37 110 38 111 
<< m1 >>
rect 38 110 39 111 
<< m1 >>
rect 39 110 40 111 
<< m1 >>
rect 40 110 41 111 
<< m2 >>
rect 40 110 41 111 
<< m1 >>
rect 41 110 42 111 
<< m1 >>
rect 42 110 43 111 
<< m2 >>
rect 42 110 43 111 
<< m2c >>
rect 42 110 43 111 
<< m1 >>
rect 42 110 43 111 
<< m2 >>
rect 42 110 43 111 
<< m2 >>
rect 43 110 44 111 
<< m1 >>
rect 44 110 45 111 
<< m2 >>
rect 44 110 45 111 
<< m2 >>
rect 45 110 46 111 
<< m1 >>
rect 46 110 47 111 
<< m2 >>
rect 46 110 47 111 
<< m2c >>
rect 46 110 47 111 
<< m1 >>
rect 46 110 47 111 
<< m2 >>
rect 46 110 47 111 
<< m1 >>
rect 49 110 50 111 
<< m1 >>
rect 50 110 51 111 
<< m1 >>
rect 51 110 52 111 
<< m1 >>
rect 52 110 53 111 
<< m1 >>
rect 53 110 54 111 
<< m1 >>
rect 54 110 55 111 
<< m1 >>
rect 55 110 56 111 
<< m2 >>
rect 56 110 57 111 
<< m2 >>
rect 59 110 60 111 
<< m2 >>
rect 64 110 65 111 
<< m1 >>
rect 67 110 68 111 
<< m1 >>
rect 68 110 69 111 
<< m1 >>
rect 69 110 70 111 
<< m1 >>
rect 70 110 71 111 
<< m1 >>
rect 71 110 72 111 
<< m2 >>
rect 71 110 72 111 
<< m2c >>
rect 71 110 72 111 
<< m1 >>
rect 71 110 72 111 
<< m2 >>
rect 71 110 72 111 
<< m2 >>
rect 72 110 73 111 
<< m1 >>
rect 73 110 74 111 
<< m2 >>
rect 73 110 74 111 
<< m2 >>
rect 74 110 75 111 
<< m1 >>
rect 75 110 76 111 
<< m2 >>
rect 75 110 76 111 
<< m2c >>
rect 75 110 76 111 
<< m1 >>
rect 75 110 76 111 
<< m2 >>
rect 75 110 76 111 
<< m1 >>
rect 77 110 78 111 
<< m2 >>
rect 77 110 78 111 
<< m2c >>
rect 77 110 78 111 
<< m1 >>
rect 77 110 78 111 
<< m2 >>
rect 77 110 78 111 
<< m1 >>
rect 82 110 83 111 
<< m1 >>
rect 83 110 84 111 
<< m1 >>
rect 84 110 85 111 
<< m2 >>
rect 84 110 85 111 
<< m2c >>
rect 84 110 85 111 
<< m1 >>
rect 84 110 85 111 
<< m2 >>
rect 84 110 85 111 
<< m1 >>
rect 91 110 92 111 
<< m2 >>
rect 91 110 92 111 
<< m2c >>
rect 91 110 92 111 
<< m1 >>
rect 91 110 92 111 
<< m2 >>
rect 91 110 92 111 
<< m1 >>
rect 100 110 101 111 
<< m2 >>
rect 100 110 101 111 
<< m2c >>
rect 100 110 101 111 
<< m1 >>
rect 100 110 101 111 
<< m2 >>
rect 100 110 101 111 
<< m1 >>
rect 103 110 104 111 
<< m2 >>
rect 103 110 104 111 
<< m2c >>
rect 103 110 104 111 
<< m1 >>
rect 103 110 104 111 
<< m2 >>
rect 103 110 104 111 
<< m1 >>
rect 109 110 110 111 
<< m1 >>
rect 118 110 119 111 
<< m2 >>
rect 118 110 119 111 
<< m2c >>
rect 118 110 119 111 
<< m1 >>
rect 118 110 119 111 
<< m2 >>
rect 118 110 119 111 
<< m1 >>
rect 124 110 125 111 
<< m1 >>
rect 126 110 127 111 
<< m1 >>
rect 129 110 130 111 
<< m1 >>
rect 131 110 132 111 
<< m1 >>
rect 154 110 155 111 
<< m1 >>
rect 163 110 164 111 
<< m1 >>
rect 165 110 166 111 
<< m1 >>
rect 167 110 168 111 
<< m2 >>
rect 171 110 172 111 
<< m1 >>
rect 172 110 173 111 
<< m1 >>
rect 181 110 182 111 
<< m2 >>
rect 182 110 183 111 
<< m2 >>
rect 185 110 186 111 
<< m1 >>
rect 190 110 191 111 
<< m1 >>
rect 199 110 200 111 
<< m1 >>
rect 201 110 202 111 
<< m1 >>
rect 218 110 219 111 
<< m1 >>
rect 220 110 221 111 
<< m1 >>
rect 244 110 245 111 
<< m1 >>
rect 247 110 248 111 
<< m1 >>
rect 253 110 254 111 
<< m2 >>
rect 254 110 255 111 
<< m1 >>
rect 256 110 257 111 
<< m1 >>
rect 19 111 20 112 
<< m1 >>
rect 28 111 29 112 
<< m2 >>
rect 37 111 38 112 
<< m2 >>
rect 40 111 41 112 
<< m1 >>
rect 44 111 45 112 
<< m2 >>
rect 56 111 57 112 
<< m1 >>
rect 57 111 58 112 
<< m2 >>
rect 57 111 58 112 
<< m2c >>
rect 57 111 58 112 
<< m1 >>
rect 57 111 58 112 
<< m2 >>
rect 57 111 58 112 
<< m1 >>
rect 58 111 59 112 
<< m1 >>
rect 59 111 60 112 
<< m2 >>
rect 59 111 60 112 
<< m1 >>
rect 60 111 61 112 
<< m1 >>
rect 61 111 62 112 
<< m1 >>
rect 62 111 63 112 
<< m1 >>
rect 63 111 64 112 
<< m1 >>
rect 64 111 65 112 
<< m2 >>
rect 64 111 65 112 
<< m1 >>
rect 73 111 74 112 
<< m1 >>
rect 75 111 76 112 
<< m2 >>
rect 77 111 78 112 
<< m2 >>
rect 84 111 85 112 
<< m2 >>
rect 91 111 92 112 
<< m2 >>
rect 100 111 101 112 
<< m2 >>
rect 103 111 104 112 
<< m1 >>
rect 109 111 110 112 
<< m2 >>
rect 118 111 119 112 
<< m2 >>
rect 122 111 123 112 
<< m2 >>
rect 123 111 124 112 
<< m1 >>
rect 124 111 125 112 
<< m2 >>
rect 124 111 125 112 
<< m2 >>
rect 125 111 126 112 
<< m1 >>
rect 126 111 127 112 
<< m2 >>
rect 126 111 127 112 
<< m2c >>
rect 126 111 127 112 
<< m1 >>
rect 126 111 127 112 
<< m2 >>
rect 126 111 127 112 
<< m1 >>
rect 129 111 130 112 
<< m2 >>
rect 129 111 130 112 
<< m2c >>
rect 129 111 130 112 
<< m1 >>
rect 129 111 130 112 
<< m2 >>
rect 129 111 130 112 
<< m1 >>
rect 131 111 132 112 
<< m2 >>
rect 131 111 132 112 
<< m2c >>
rect 131 111 132 112 
<< m1 >>
rect 131 111 132 112 
<< m2 >>
rect 131 111 132 112 
<< m1 >>
rect 154 111 155 112 
<< m1 >>
rect 163 111 164 112 
<< m2 >>
rect 163 111 164 112 
<< m2c >>
rect 163 111 164 112 
<< m1 >>
rect 163 111 164 112 
<< m2 >>
rect 163 111 164 112 
<< m1 >>
rect 165 111 166 112 
<< m2 >>
rect 165 111 166 112 
<< m2c >>
rect 165 111 166 112 
<< m1 >>
rect 165 111 166 112 
<< m2 >>
rect 165 111 166 112 
<< m1 >>
rect 167 111 168 112 
<< m2 >>
rect 167 111 168 112 
<< m2c >>
rect 167 111 168 112 
<< m1 >>
rect 167 111 168 112 
<< m2 >>
rect 167 111 168 112 
<< m2 >>
rect 171 111 172 112 
<< m1 >>
rect 172 111 173 112 
<< m1 >>
rect 181 111 182 112 
<< m2 >>
rect 182 111 183 112 
<< m1 >>
rect 183 111 184 112 
<< m2 >>
rect 183 111 184 112 
<< m2c >>
rect 183 111 184 112 
<< m1 >>
rect 183 111 184 112 
<< m2 >>
rect 183 111 184 112 
<< m1 >>
rect 184 111 185 112 
<< m1 >>
rect 185 111 186 112 
<< m2 >>
rect 185 111 186 112 
<< m1 >>
rect 186 111 187 112 
<< m1 >>
rect 187 111 188 112 
<< m1 >>
rect 188 111 189 112 
<< m2 >>
rect 188 111 189 112 
<< m2c >>
rect 188 111 189 112 
<< m1 >>
rect 188 111 189 112 
<< m2 >>
rect 188 111 189 112 
<< m2 >>
rect 189 111 190 112 
<< m1 >>
rect 190 111 191 112 
<< m2 >>
rect 190 111 191 112 
<< m2 >>
rect 191 111 192 112 
<< m1 >>
rect 192 111 193 112 
<< m2 >>
rect 192 111 193 112 
<< m2c >>
rect 192 111 193 112 
<< m1 >>
rect 192 111 193 112 
<< m2 >>
rect 192 111 193 112 
<< m1 >>
rect 197 111 198 112 
<< m2 >>
rect 197 111 198 112 
<< m2c >>
rect 197 111 198 112 
<< m1 >>
rect 197 111 198 112 
<< m2 >>
rect 197 111 198 112 
<< m2 >>
rect 198 111 199 112 
<< m1 >>
rect 199 111 200 112 
<< m2 >>
rect 199 111 200 112 
<< m2 >>
rect 200 111 201 112 
<< m1 >>
rect 201 111 202 112 
<< m2 >>
rect 201 111 202 112 
<< m2 >>
rect 202 111 203 112 
<< m1 >>
rect 203 111 204 112 
<< m2 >>
rect 203 111 204 112 
<< m2c >>
rect 203 111 204 112 
<< m1 >>
rect 203 111 204 112 
<< m2 >>
rect 203 111 204 112 
<< m1 >>
rect 204 111 205 112 
<< m1 >>
rect 205 111 206 112 
<< m1 >>
rect 206 111 207 112 
<< m1 >>
rect 207 111 208 112 
<< m1 >>
rect 208 111 209 112 
<< m1 >>
rect 209 111 210 112 
<< m1 >>
rect 210 111 211 112 
<< m1 >>
rect 218 111 219 112 
<< m1 >>
rect 220 111 221 112 
<< m1 >>
rect 244 111 245 112 
<< m1 >>
rect 247 111 248 112 
<< m1 >>
rect 253 111 254 112 
<< m2 >>
rect 254 111 255 112 
<< m1 >>
rect 256 111 257 112 
<< m1 >>
rect 19 112 20 113 
<< m1 >>
rect 28 112 29 113 
<< m1 >>
rect 37 112 38 113 
<< m2 >>
rect 37 112 38 113 
<< m2c >>
rect 37 112 38 113 
<< m1 >>
rect 37 112 38 113 
<< m2 >>
rect 37 112 38 113 
<< m1 >>
rect 40 112 41 113 
<< m2 >>
rect 40 112 41 113 
<< m2c >>
rect 40 112 41 113 
<< m1 >>
rect 40 112 41 113 
<< m2 >>
rect 40 112 41 113 
<< m1 >>
rect 41 112 42 113 
<< m1 >>
rect 42 112 43 113 
<< m2 >>
rect 42 112 43 113 
<< m2c >>
rect 42 112 43 113 
<< m1 >>
rect 42 112 43 113 
<< m2 >>
rect 42 112 43 113 
<< m2 >>
rect 43 112 44 113 
<< m1 >>
rect 44 112 45 113 
<< m2 >>
rect 44 112 45 113 
<< m2 >>
rect 45 112 46 113 
<< m1 >>
rect 46 112 47 113 
<< m2 >>
rect 46 112 47 113 
<< m2c >>
rect 46 112 47 113 
<< m1 >>
rect 46 112 47 113 
<< m2 >>
rect 46 112 47 113 
<< m1 >>
rect 47 112 48 113 
<< m1 >>
rect 48 112 49 113 
<< m2 >>
rect 59 112 60 113 
<< m1 >>
rect 64 112 65 113 
<< m2 >>
rect 64 112 65 113 
<< m1 >>
rect 73 112 74 113 
<< m1 >>
rect 75 112 76 113 
<< m1 >>
rect 76 112 77 113 
<< m1 >>
rect 77 112 78 113 
<< m2 >>
rect 77 112 78 113 
<< m1 >>
rect 78 112 79 113 
<< m1 >>
rect 79 112 80 113 
<< m1 >>
rect 80 112 81 113 
<< m1 >>
rect 81 112 82 113 
<< m1 >>
rect 82 112 83 113 
<< m1 >>
rect 83 112 84 113 
<< m1 >>
rect 84 112 85 113 
<< m2 >>
rect 84 112 85 113 
<< m1 >>
rect 85 112 86 113 
<< m1 >>
rect 86 112 87 113 
<< m1 >>
rect 87 112 88 113 
<< m1 >>
rect 88 112 89 113 
<< m1 >>
rect 89 112 90 113 
<< m1 >>
rect 90 112 91 113 
<< m1 >>
rect 91 112 92 113 
<< m2 >>
rect 91 112 92 113 
<< m1 >>
rect 92 112 93 113 
<< m1 >>
rect 93 112 94 113 
<< m1 >>
rect 94 112 95 113 
<< m1 >>
rect 95 112 96 113 
<< m1 >>
rect 96 112 97 113 
<< m1 >>
rect 97 112 98 113 
<< m1 >>
rect 98 112 99 113 
<< m1 >>
rect 99 112 100 113 
<< m1 >>
rect 100 112 101 113 
<< m2 >>
rect 100 112 101 113 
<< m1 >>
rect 101 112 102 113 
<< m1 >>
rect 102 112 103 113 
<< m1 >>
rect 103 112 104 113 
<< m2 >>
rect 103 112 104 113 
<< m1 >>
rect 104 112 105 113 
<< m1 >>
rect 109 112 110 113 
<< m1 >>
rect 110 112 111 113 
<< m1 >>
rect 111 112 112 113 
<< m1 >>
rect 112 112 113 113 
<< m1 >>
rect 113 112 114 113 
<< m1 >>
rect 114 112 115 113 
<< m1 >>
rect 115 112 116 113 
<< m1 >>
rect 116 112 117 113 
<< m1 >>
rect 117 112 118 113 
<< m1 >>
rect 118 112 119 113 
<< m2 >>
rect 118 112 119 113 
<< m1 >>
rect 119 112 120 113 
<< m1 >>
rect 120 112 121 113 
<< m1 >>
rect 121 112 122 113 
<< m1 >>
rect 122 112 123 113 
<< m2 >>
rect 122 112 123 113 
<< m1 >>
rect 123 112 124 113 
<< m1 >>
rect 124 112 125 113 
<< m2 >>
rect 129 112 130 113 
<< m2 >>
rect 131 112 132 113 
<< m2 >>
rect 132 112 133 113 
<< m2 >>
rect 133 112 134 113 
<< m2 >>
rect 134 112 135 113 
<< m2 >>
rect 135 112 136 113 
<< m2 >>
rect 136 112 137 113 
<< m2 >>
rect 137 112 138 113 
<< m2 >>
rect 138 112 139 113 
<< m2 >>
rect 139 112 140 113 
<< m2 >>
rect 140 112 141 113 
<< m1 >>
rect 154 112 155 113 
<< m2 >>
rect 163 112 164 113 
<< m2 >>
rect 165 112 166 113 
<< m2 >>
rect 167 112 168 113 
<< m2 >>
rect 171 112 172 113 
<< m1 >>
rect 172 112 173 113 
<< m1 >>
rect 181 112 182 113 
<< m2 >>
rect 185 112 186 113 
<< m1 >>
rect 190 112 191 113 
<< m1 >>
rect 192 112 193 113 
<< m1 >>
rect 193 112 194 113 
<< m1 >>
rect 194 112 195 113 
<< m1 >>
rect 195 112 196 113 
<< m1 >>
rect 196 112 197 113 
<< m1 >>
rect 197 112 198 113 
<< m1 >>
rect 199 112 200 113 
<< m1 >>
rect 201 112 202 113 
<< m1 >>
rect 210 112 211 113 
<< m1 >>
rect 218 112 219 113 
<< m1 >>
rect 220 112 221 113 
<< m1 >>
rect 221 112 222 113 
<< m1 >>
rect 222 112 223 113 
<< m1 >>
rect 223 112 224 113 
<< m1 >>
rect 224 112 225 113 
<< m1 >>
rect 225 112 226 113 
<< m1 >>
rect 226 112 227 113 
<< m1 >>
rect 227 112 228 113 
<< m1 >>
rect 228 112 229 113 
<< m1 >>
rect 229 112 230 113 
<< m1 >>
rect 230 112 231 113 
<< m1 >>
rect 231 112 232 113 
<< m1 >>
rect 244 112 245 113 
<< m1 >>
rect 247 112 248 113 
<< m1 >>
rect 253 112 254 113 
<< m2 >>
rect 254 112 255 113 
<< m1 >>
rect 256 112 257 113 
<< m1 >>
rect 19 113 20 114 
<< m2 >>
rect 19 113 20 114 
<< m2c >>
rect 19 113 20 114 
<< m1 >>
rect 19 113 20 114 
<< m2 >>
rect 19 113 20 114 
<< m1 >>
rect 28 113 29 114 
<< m2 >>
rect 28 113 29 114 
<< m2c >>
rect 28 113 29 114 
<< m1 >>
rect 28 113 29 114 
<< m2 >>
rect 28 113 29 114 
<< m1 >>
rect 37 113 38 114 
<< m2 >>
rect 37 113 38 114 
<< m1 >>
rect 44 113 45 114 
<< m1 >>
rect 48 113 49 114 
<< m2 >>
rect 48 113 49 114 
<< m2c >>
rect 48 113 49 114 
<< m1 >>
rect 48 113 49 114 
<< m2 >>
rect 48 113 49 114 
<< m1 >>
rect 59 113 60 114 
<< m2 >>
rect 59 113 60 114 
<< m2c >>
rect 59 113 60 114 
<< m1 >>
rect 59 113 60 114 
<< m2 >>
rect 59 113 60 114 
<< m1 >>
rect 64 113 65 114 
<< m2 >>
rect 64 113 65 114 
<< m1 >>
rect 73 113 74 114 
<< m2 >>
rect 77 113 78 114 
<< m2 >>
rect 84 113 85 114 
<< m2 >>
rect 85 113 86 114 
<< m2 >>
rect 91 113 92 114 
<< m2 >>
rect 100 113 101 114 
<< m2 >>
rect 103 113 104 114 
<< m1 >>
rect 104 113 105 114 
<< m2 >>
rect 118 113 119 114 
<< m2 >>
rect 122 113 123 114 
<< m1 >>
rect 127 113 128 114 
<< m2 >>
rect 127 113 128 114 
<< m2c >>
rect 127 113 128 114 
<< m1 >>
rect 127 113 128 114 
<< m2 >>
rect 127 113 128 114 
<< m1 >>
rect 128 113 129 114 
<< m1 >>
rect 129 113 130 114 
<< m2 >>
rect 129 113 130 114 
<< m1 >>
rect 130 113 131 114 
<< m1 >>
rect 131 113 132 114 
<< m1 >>
rect 132 113 133 114 
<< m1 >>
rect 133 113 134 114 
<< m1 >>
rect 134 113 135 114 
<< m1 >>
rect 135 113 136 114 
<< m1 >>
rect 136 113 137 114 
<< m1 >>
rect 137 113 138 114 
<< m1 >>
rect 138 113 139 114 
<< m1 >>
rect 139 113 140 114 
<< m1 >>
rect 140 113 141 114 
<< m2 >>
rect 140 113 141 114 
<< m1 >>
rect 141 113 142 114 
<< m1 >>
rect 142 113 143 114 
<< m1 >>
rect 143 113 144 114 
<< m1 >>
rect 144 113 145 114 
<< m1 >>
rect 145 113 146 114 
<< m1 >>
rect 146 113 147 114 
<< m1 >>
rect 147 113 148 114 
<< m1 >>
rect 148 113 149 114 
<< m1 >>
rect 149 113 150 114 
<< m1 >>
rect 150 113 151 114 
<< m1 >>
rect 151 113 152 114 
<< m1 >>
rect 152 113 153 114 
<< m2 >>
rect 152 113 153 114 
<< m2c >>
rect 152 113 153 114 
<< m1 >>
rect 152 113 153 114 
<< m2 >>
rect 152 113 153 114 
<< m2 >>
rect 153 113 154 114 
<< m1 >>
rect 154 113 155 114 
<< m2 >>
rect 154 113 155 114 
<< m2 >>
rect 155 113 156 114 
<< m1 >>
rect 156 113 157 114 
<< m2 >>
rect 156 113 157 114 
<< m2c >>
rect 156 113 157 114 
<< m1 >>
rect 156 113 157 114 
<< m2 >>
rect 156 113 157 114 
<< m1 >>
rect 157 113 158 114 
<< m1 >>
rect 158 113 159 114 
<< m1 >>
rect 159 113 160 114 
<< m1 >>
rect 160 113 161 114 
<< m1 >>
rect 161 113 162 114 
<< m1 >>
rect 162 113 163 114 
<< m1 >>
rect 163 113 164 114 
<< m2 >>
rect 163 113 164 114 
<< m1 >>
rect 164 113 165 114 
<< m1 >>
rect 165 113 166 114 
<< m2 >>
rect 165 113 166 114 
<< m1 >>
rect 166 113 167 114 
<< m1 >>
rect 167 113 168 114 
<< m2 >>
rect 167 113 168 114 
<< m1 >>
rect 168 113 169 114 
<< m1 >>
rect 169 113 170 114 
<< m1 >>
rect 170 113 171 114 
<< m2 >>
rect 170 113 171 114 
<< m2c >>
rect 170 113 171 114 
<< m1 >>
rect 170 113 171 114 
<< m2 >>
rect 170 113 171 114 
<< m2 >>
rect 171 113 172 114 
<< m1 >>
rect 172 113 173 114 
<< m1 >>
rect 181 113 182 114 
<< m2 >>
rect 181 113 182 114 
<< m2c >>
rect 181 113 182 114 
<< m1 >>
rect 181 113 182 114 
<< m2 >>
rect 181 113 182 114 
<< m1 >>
rect 183 113 184 114 
<< m2 >>
rect 183 113 184 114 
<< m2c >>
rect 183 113 184 114 
<< m1 >>
rect 183 113 184 114 
<< m2 >>
rect 183 113 184 114 
<< m1 >>
rect 184 113 185 114 
<< m1 >>
rect 185 113 186 114 
<< m2 >>
rect 185 113 186 114 
<< m2c >>
rect 185 113 186 114 
<< m1 >>
rect 185 113 186 114 
<< m2 >>
rect 185 113 186 114 
<< m1 >>
rect 190 113 191 114 
<< m2 >>
rect 190 113 191 114 
<< m2c >>
rect 190 113 191 114 
<< m1 >>
rect 190 113 191 114 
<< m2 >>
rect 190 113 191 114 
<< m1 >>
rect 199 113 200 114 
<< m2 >>
rect 199 113 200 114 
<< m2c >>
rect 199 113 200 114 
<< m1 >>
rect 199 113 200 114 
<< m2 >>
rect 199 113 200 114 
<< m1 >>
rect 201 113 202 114 
<< m2 >>
rect 201 113 202 114 
<< m2c >>
rect 201 113 202 114 
<< m1 >>
rect 201 113 202 114 
<< m2 >>
rect 201 113 202 114 
<< m1 >>
rect 210 113 211 114 
<< m1 >>
rect 211 113 212 114 
<< m1 >>
rect 212 113 213 114 
<< m1 >>
rect 213 113 214 114 
<< m1 >>
rect 214 113 215 114 
<< m1 >>
rect 215 113 216 114 
<< m1 >>
rect 216 113 217 114 
<< m2 >>
rect 216 113 217 114 
<< m2c >>
rect 216 113 217 114 
<< m1 >>
rect 216 113 217 114 
<< m2 >>
rect 216 113 217 114 
<< m2 >>
rect 217 113 218 114 
<< m1 >>
rect 218 113 219 114 
<< m2 >>
rect 218 113 219 114 
<< m2 >>
rect 219 113 220 114 
<< m1 >>
rect 231 113 232 114 
<< m2 >>
rect 231 113 232 114 
<< m2c >>
rect 231 113 232 114 
<< m1 >>
rect 231 113 232 114 
<< m2 >>
rect 231 113 232 114 
<< m1 >>
rect 244 113 245 114 
<< m2 >>
rect 244 113 245 114 
<< m2c >>
rect 244 113 245 114 
<< m1 >>
rect 244 113 245 114 
<< m2 >>
rect 244 113 245 114 
<< m1 >>
rect 247 113 248 114 
<< m1 >>
rect 253 113 254 114 
<< m2 >>
rect 254 113 255 114 
<< m1 >>
rect 256 113 257 114 
<< m2 >>
rect 19 114 20 115 
<< m2 >>
rect 28 114 29 115 
<< m2 >>
rect 37 114 38 115 
<< m1 >>
rect 44 114 45 115 
<< m2 >>
rect 48 114 49 115 
<< m2 >>
rect 49 114 50 115 
<< m2 >>
rect 50 114 51 115 
<< m1 >>
rect 59 114 60 115 
<< m1 >>
rect 64 114 65 115 
<< m2 >>
rect 64 114 65 115 
<< m1 >>
rect 73 114 74 115 
<< m1 >>
rect 77 114 78 115 
<< m2 >>
rect 77 114 78 115 
<< m2c >>
rect 77 114 78 115 
<< m1 >>
rect 77 114 78 115 
<< m2 >>
rect 77 114 78 115 
<< m1 >>
rect 85 114 86 115 
<< m2 >>
rect 85 114 86 115 
<< m2c >>
rect 85 114 86 115 
<< m1 >>
rect 85 114 86 115 
<< m2 >>
rect 85 114 86 115 
<< m1 >>
rect 91 114 92 115 
<< m2 >>
rect 91 114 92 115 
<< m2c >>
rect 91 114 92 115 
<< m1 >>
rect 91 114 92 115 
<< m2 >>
rect 91 114 92 115 
<< m1 >>
rect 100 114 101 115 
<< m2 >>
rect 100 114 101 115 
<< m1 >>
rect 101 114 102 115 
<< m1 >>
rect 102 114 103 115 
<< m2 >>
rect 102 114 103 115 
<< m2c >>
rect 102 114 103 115 
<< m1 >>
rect 102 114 103 115 
<< m2 >>
rect 102 114 103 115 
<< m2 >>
rect 103 114 104 115 
<< m1 >>
rect 104 114 105 115 
<< m1 >>
rect 118 114 119 115 
<< m2 >>
rect 118 114 119 115 
<< m2c >>
rect 118 114 119 115 
<< m1 >>
rect 118 114 119 115 
<< m2 >>
rect 118 114 119 115 
<< m2 >>
rect 122 114 123 115 
<< m2 >>
rect 127 114 128 115 
<< m2 >>
rect 129 114 130 115 
<< m2 >>
rect 140 114 141 115 
<< m1 >>
rect 154 114 155 115 
<< m2 >>
rect 163 114 164 115 
<< m2 >>
rect 165 114 166 115 
<< m2 >>
rect 167 114 168 115 
<< m1 >>
rect 172 114 173 115 
<< m2 >>
rect 181 114 182 115 
<< m2 >>
rect 183 114 184 115 
<< m2 >>
rect 190 114 191 115 
<< m2 >>
rect 199 114 200 115 
<< m2 >>
rect 201 114 202 115 
<< m1 >>
rect 218 114 219 115 
<< m2 >>
rect 219 114 220 115 
<< m2 >>
rect 231 114 232 115 
<< m2 >>
rect 244 114 245 115 
<< m1 >>
rect 247 114 248 115 
<< m1 >>
rect 253 114 254 115 
<< m2 >>
rect 254 114 255 115 
<< m1 >>
rect 256 114 257 115 
<< m1 >>
rect 19 115 20 116 
<< m2 >>
rect 19 115 20 116 
<< m1 >>
rect 20 115 21 116 
<< m1 >>
rect 21 115 22 116 
<< m1 >>
rect 22 115 23 116 
<< m1 >>
rect 23 115 24 116 
<< m1 >>
rect 24 115 25 116 
<< m1 >>
rect 25 115 26 116 
<< m1 >>
rect 26 115 27 116 
<< m1 >>
rect 27 115 28 116 
<< m1 >>
rect 28 115 29 116 
<< m2 >>
rect 28 115 29 116 
<< m1 >>
rect 29 115 30 116 
<< m1 >>
rect 30 115 31 116 
<< m1 >>
rect 31 115 32 116 
<< m1 >>
rect 32 115 33 116 
<< m1 >>
rect 33 115 34 116 
<< m1 >>
rect 34 115 35 116 
<< m1 >>
rect 35 115 36 116 
<< m1 >>
rect 36 115 37 116 
<< m1 >>
rect 37 115 38 116 
<< m2 >>
rect 37 115 38 116 
<< m1 >>
rect 38 115 39 116 
<< m1 >>
rect 39 115 40 116 
<< m1 >>
rect 40 115 41 116 
<< m1 >>
rect 41 115 42 116 
<< m1 >>
rect 42 115 43 116 
<< m2 >>
rect 42 115 43 116 
<< m2c >>
rect 42 115 43 116 
<< m1 >>
rect 42 115 43 116 
<< m2 >>
rect 42 115 43 116 
<< m2 >>
rect 43 115 44 116 
<< m1 >>
rect 44 115 45 116 
<< m2 >>
rect 44 115 45 116 
<< m2 >>
rect 45 115 46 116 
<< m1 >>
rect 46 115 47 116 
<< m2 >>
rect 46 115 47 116 
<< m2c >>
rect 46 115 47 116 
<< m1 >>
rect 46 115 47 116 
<< m2 >>
rect 46 115 47 116 
<< m1 >>
rect 47 115 48 116 
<< m1 >>
rect 48 115 49 116 
<< m1 >>
rect 49 115 50 116 
<< m1 >>
rect 50 115 51 116 
<< m2 >>
rect 50 115 51 116 
<< m1 >>
rect 51 115 52 116 
<< m1 >>
rect 52 115 53 116 
<< m1 >>
rect 53 115 54 116 
<< m1 >>
rect 54 115 55 116 
<< m1 >>
rect 55 115 56 116 
<< m1 >>
rect 56 115 57 116 
<< m1 >>
rect 57 115 58 116 
<< m1 >>
rect 58 115 59 116 
<< m1 >>
rect 59 115 60 116 
<< m1 >>
rect 64 115 65 116 
<< m2 >>
rect 64 115 65 116 
<< m1 >>
rect 73 115 74 116 
<< m1 >>
rect 77 115 78 116 
<< m1 >>
rect 85 115 86 116 
<< m1 >>
rect 91 115 92 116 
<< m1 >>
rect 100 115 101 116 
<< m2 >>
rect 100 115 101 116 
<< m1 >>
rect 104 115 105 116 
<< m1 >>
rect 118 115 119 116 
<< m1 >>
rect 120 115 121 116 
<< m1 >>
rect 121 115 122 116 
<< m1 >>
rect 122 115 123 116 
<< m2 >>
rect 122 115 123 116 
<< m1 >>
rect 123 115 124 116 
<< m1 >>
rect 124 115 125 116 
<< m1 >>
rect 125 115 126 116 
<< m1 >>
rect 126 115 127 116 
<< m1 >>
rect 127 115 128 116 
<< m2 >>
rect 127 115 128 116 
<< m1 >>
rect 128 115 129 116 
<< m1 >>
rect 129 115 130 116 
<< m2 >>
rect 129 115 130 116 
<< m1 >>
rect 130 115 131 116 
<< m1 >>
rect 131 115 132 116 
<< m1 >>
rect 132 115 133 116 
<< m1 >>
rect 133 115 134 116 
<< m1 >>
rect 134 115 135 116 
<< m1 >>
rect 135 115 136 116 
<< m1 >>
rect 136 115 137 116 
<< m1 >>
rect 137 115 138 116 
<< m1 >>
rect 138 115 139 116 
<< m1 >>
rect 139 115 140 116 
<< m1 >>
rect 140 115 141 116 
<< m2 >>
rect 140 115 141 116 
<< m1 >>
rect 141 115 142 116 
<< m1 >>
rect 142 115 143 116 
<< m1 >>
rect 143 115 144 116 
<< m1 >>
rect 144 115 145 116 
<< m1 >>
rect 145 115 146 116 
<< m1 >>
rect 146 115 147 116 
<< m1 >>
rect 147 115 148 116 
<< m1 >>
rect 148 115 149 116 
<< m1 >>
rect 149 115 150 116 
<< m1 >>
rect 150 115 151 116 
<< m1 >>
rect 151 115 152 116 
<< m1 >>
rect 152 115 153 116 
<< m2 >>
rect 152 115 153 116 
<< m2c >>
rect 152 115 153 116 
<< m1 >>
rect 152 115 153 116 
<< m2 >>
rect 152 115 153 116 
<< m2 >>
rect 153 115 154 116 
<< m1 >>
rect 154 115 155 116 
<< m2 >>
rect 154 115 155 116 
<< m2 >>
rect 155 115 156 116 
<< m1 >>
rect 156 115 157 116 
<< m2 >>
rect 156 115 157 116 
<< m2c >>
rect 156 115 157 116 
<< m1 >>
rect 156 115 157 116 
<< m2 >>
rect 156 115 157 116 
<< m1 >>
rect 157 115 158 116 
<< m1 >>
rect 158 115 159 116 
<< m1 >>
rect 159 115 160 116 
<< m1 >>
rect 160 115 161 116 
<< m1 >>
rect 161 115 162 116 
<< m1 >>
rect 162 115 163 116 
<< m1 >>
rect 163 115 164 116 
<< m2 >>
rect 163 115 164 116 
<< m1 >>
rect 164 115 165 116 
<< m1 >>
rect 165 115 166 116 
<< m2 >>
rect 165 115 166 116 
<< m1 >>
rect 166 115 167 116 
<< m1 >>
rect 167 115 168 116 
<< m2 >>
rect 167 115 168 116 
<< m1 >>
rect 168 115 169 116 
<< m1 >>
rect 169 115 170 116 
<< m1 >>
rect 170 115 171 116 
<< m2 >>
rect 170 115 171 116 
<< m2c >>
rect 170 115 171 116 
<< m1 >>
rect 170 115 171 116 
<< m2 >>
rect 170 115 171 116 
<< m2 >>
rect 171 115 172 116 
<< m1 >>
rect 172 115 173 116 
<< m2 >>
rect 172 115 173 116 
<< m2 >>
rect 173 115 174 116 
<< m1 >>
rect 174 115 175 116 
<< m2 >>
rect 174 115 175 116 
<< m2c >>
rect 174 115 175 116 
<< m1 >>
rect 174 115 175 116 
<< m2 >>
rect 174 115 175 116 
<< m1 >>
rect 175 115 176 116 
<< m1 >>
rect 176 115 177 116 
<< m1 >>
rect 177 115 178 116 
<< m1 >>
rect 178 115 179 116 
<< m1 >>
rect 179 115 180 116 
<< m1 >>
rect 180 115 181 116 
<< m1 >>
rect 181 115 182 116 
<< m2 >>
rect 181 115 182 116 
<< m1 >>
rect 182 115 183 116 
<< m1 >>
rect 183 115 184 116 
<< m2 >>
rect 183 115 184 116 
<< m1 >>
rect 184 115 185 116 
<< m1 >>
rect 185 115 186 116 
<< m1 >>
rect 186 115 187 116 
<< m1 >>
rect 187 115 188 116 
<< m1 >>
rect 188 115 189 116 
<< m1 >>
rect 189 115 190 116 
<< m1 >>
rect 190 115 191 116 
<< m2 >>
rect 190 115 191 116 
<< m1 >>
rect 191 115 192 116 
<< m1 >>
rect 192 115 193 116 
<< m2 >>
rect 192 115 193 116 
<< m1 >>
rect 193 115 194 116 
<< m2 >>
rect 193 115 194 116 
<< m1 >>
rect 194 115 195 116 
<< m2 >>
rect 194 115 195 116 
<< m1 >>
rect 195 115 196 116 
<< m2 >>
rect 195 115 196 116 
<< m1 >>
rect 196 115 197 116 
<< m2 >>
rect 196 115 197 116 
<< m1 >>
rect 197 115 198 116 
<< m1 >>
rect 198 115 199 116 
<< m1 >>
rect 199 115 200 116 
<< m2 >>
rect 199 115 200 116 
<< m1 >>
rect 200 115 201 116 
<< m1 >>
rect 201 115 202 116 
<< m2 >>
rect 201 115 202 116 
<< m1 >>
rect 202 115 203 116 
<< m1 >>
rect 203 115 204 116 
<< m2 >>
rect 203 115 204 116 
<< m1 >>
rect 204 115 205 116 
<< m2 >>
rect 204 115 205 116 
<< m1 >>
rect 205 115 206 116 
<< m2 >>
rect 205 115 206 116 
<< m1 >>
rect 206 115 207 116 
<< m2 >>
rect 206 115 207 116 
<< m1 >>
rect 207 115 208 116 
<< m2 >>
rect 207 115 208 116 
<< m1 >>
rect 208 115 209 116 
<< m2 >>
rect 208 115 209 116 
<< m1 >>
rect 209 115 210 116 
<< m2 >>
rect 209 115 210 116 
<< m1 >>
rect 210 115 211 116 
<< m2 >>
rect 210 115 211 116 
<< m1 >>
rect 211 115 212 116 
<< m2 >>
rect 211 115 212 116 
<< m2 >>
rect 212 115 213 116 
<< m1 >>
rect 213 115 214 116 
<< m2 >>
rect 213 115 214 116 
<< m2c >>
rect 213 115 214 116 
<< m1 >>
rect 213 115 214 116 
<< m2 >>
rect 213 115 214 116 
<< m1 >>
rect 214 115 215 116 
<< m1 >>
rect 215 115 216 116 
<< m1 >>
rect 216 115 217 116 
<< m1 >>
rect 217 115 218 116 
<< m1 >>
rect 218 115 219 116 
<< m2 >>
rect 219 115 220 116 
<< m2 >>
rect 231 115 232 116 
<< m1 >>
rect 232 115 233 116 
<< m1 >>
rect 233 115 234 116 
<< m1 >>
rect 234 115 235 116 
<< m1 >>
rect 235 115 236 116 
<< m1 >>
rect 236 115 237 116 
<< m1 >>
rect 237 115 238 116 
<< m1 >>
rect 238 115 239 116 
<< m1 >>
rect 239 115 240 116 
<< m1 >>
rect 240 115 241 116 
<< m1 >>
rect 241 115 242 116 
<< m1 >>
rect 242 115 243 116 
<< m1 >>
rect 243 115 244 116 
<< m1 >>
rect 244 115 245 116 
<< m2 >>
rect 244 115 245 116 
<< m1 >>
rect 245 115 246 116 
<< m1 >>
rect 246 115 247 116 
<< m1 >>
rect 247 115 248 116 
<< m1 >>
rect 253 115 254 116 
<< m2 >>
rect 254 115 255 116 
<< m1 >>
rect 256 115 257 116 
<< m1 >>
rect 19 116 20 117 
<< m2 >>
rect 19 116 20 117 
<< m2 >>
rect 28 116 29 117 
<< m2 >>
rect 37 116 38 117 
<< m1 >>
rect 44 116 45 117 
<< m2 >>
rect 50 116 51 117 
<< m1 >>
rect 64 116 65 117 
<< m2 >>
rect 64 116 65 117 
<< m1 >>
rect 73 116 74 117 
<< m1 >>
rect 77 116 78 117 
<< m1 >>
rect 85 116 86 117 
<< m1 >>
rect 91 116 92 117 
<< m2 >>
rect 91 116 92 117 
<< m2c >>
rect 91 116 92 117 
<< m1 >>
rect 91 116 92 117 
<< m2 >>
rect 91 116 92 117 
<< m1 >>
rect 100 116 101 117 
<< m2 >>
rect 100 116 101 117 
<< m1 >>
rect 104 116 105 117 
<< m1 >>
rect 105 116 106 117 
<< m1 >>
rect 106 116 107 117 
<< m1 >>
rect 107 116 108 117 
<< m1 >>
rect 108 116 109 117 
<< m1 >>
rect 109 116 110 117 
<< m1 >>
rect 110 116 111 117 
<< m1 >>
rect 111 116 112 117 
<< m1 >>
rect 112 116 113 117 
<< m1 >>
rect 113 116 114 117 
<< m1 >>
rect 114 116 115 117 
<< m1 >>
rect 115 116 116 117 
<< m1 >>
rect 116 116 117 117 
<< m2 >>
rect 116 116 117 117 
<< m2c >>
rect 116 116 117 117 
<< m1 >>
rect 116 116 117 117 
<< m2 >>
rect 116 116 117 117 
<< m2 >>
rect 117 116 118 117 
<< m1 >>
rect 118 116 119 117 
<< m2 >>
rect 118 116 119 117 
<< m2 >>
rect 119 116 120 117 
<< m1 >>
rect 120 116 121 117 
<< m2 >>
rect 120 116 121 117 
<< m2c >>
rect 120 116 121 117 
<< m1 >>
rect 120 116 121 117 
<< m2 >>
rect 120 116 121 117 
<< m2 >>
rect 122 116 123 117 
<< m2 >>
rect 127 116 128 117 
<< m2 >>
rect 129 116 130 117 
<< m2 >>
rect 140 116 141 117 
<< m1 >>
rect 154 116 155 117 
<< m2 >>
rect 163 116 164 117 
<< m2 >>
rect 165 116 166 117 
<< m2 >>
rect 167 116 168 117 
<< m1 >>
rect 172 116 173 117 
<< m2 >>
rect 181 116 182 117 
<< m2 >>
rect 183 116 184 117 
<< m2 >>
rect 190 116 191 117 
<< m2 >>
rect 192 116 193 117 
<< m2 >>
rect 196 116 197 117 
<< m2 >>
rect 199 116 200 117 
<< m2 >>
rect 201 116 202 117 
<< m2 >>
rect 203 116 204 117 
<< m1 >>
rect 211 116 212 117 
<< m2 >>
rect 219 116 220 117 
<< m2 >>
rect 231 116 232 117 
<< m1 >>
rect 232 116 233 117 
<< m2 >>
rect 244 116 245 117 
<< m1 >>
rect 253 116 254 117 
<< m2 >>
rect 254 116 255 117 
<< m1 >>
rect 256 116 257 117 
<< m1 >>
rect 19 117 20 118 
<< m2 >>
rect 19 117 20 118 
<< m2 >>
rect 28 117 29 118 
<< m1 >>
rect 37 117 38 118 
<< m2 >>
rect 37 117 38 118 
<< m2c >>
rect 37 117 38 118 
<< m1 >>
rect 37 117 38 118 
<< m2 >>
rect 37 117 38 118 
<< m1 >>
rect 38 117 39 118 
<< m1 >>
rect 39 117 40 118 
<< m1 >>
rect 40 117 41 118 
<< m1 >>
rect 41 117 42 118 
<< m1 >>
rect 42 117 43 118 
<< m2 >>
rect 42 117 43 118 
<< m2c >>
rect 42 117 43 118 
<< m1 >>
rect 42 117 43 118 
<< m2 >>
rect 42 117 43 118 
<< m2 >>
rect 43 117 44 118 
<< m1 >>
rect 44 117 45 118 
<< m2 >>
rect 44 117 45 118 
<< m2 >>
rect 45 117 46 118 
<< m1 >>
rect 46 117 47 118 
<< m2 >>
rect 46 117 47 118 
<< m2c >>
rect 46 117 47 118 
<< m1 >>
rect 46 117 47 118 
<< m2 >>
rect 46 117 47 118 
<< m1 >>
rect 50 117 51 118 
<< m2 >>
rect 50 117 51 118 
<< m2c >>
rect 50 117 51 118 
<< m1 >>
rect 50 117 51 118 
<< m2 >>
rect 50 117 51 118 
<< m1 >>
rect 51 117 52 118 
<< m1 >>
rect 52 117 53 118 
<< m1 >>
rect 53 117 54 118 
<< m1 >>
rect 54 117 55 118 
<< m1 >>
rect 55 117 56 118 
<< m1 >>
rect 56 117 57 118 
<< m1 >>
rect 57 117 58 118 
<< m1 >>
rect 64 117 65 118 
<< m2 >>
rect 64 117 65 118 
<< m1 >>
rect 73 117 74 118 
<< m1 >>
rect 77 117 78 118 
<< m1 >>
rect 85 117 86 118 
<< m2 >>
rect 91 117 92 118 
<< m1 >>
rect 100 117 101 118 
<< m2 >>
rect 100 117 101 118 
<< m1 >>
rect 118 117 119 118 
<< m1 >>
rect 122 117 123 118 
<< m2 >>
rect 122 117 123 118 
<< m2c >>
rect 122 117 123 118 
<< m1 >>
rect 122 117 123 118 
<< m2 >>
rect 122 117 123 118 
<< m1 >>
rect 127 117 128 118 
<< m2 >>
rect 127 117 128 118 
<< m2c >>
rect 127 117 128 118 
<< m1 >>
rect 127 117 128 118 
<< m2 >>
rect 127 117 128 118 
<< m1 >>
rect 129 117 130 118 
<< m2 >>
rect 129 117 130 118 
<< m2c >>
rect 129 117 130 118 
<< m1 >>
rect 129 117 130 118 
<< m2 >>
rect 129 117 130 118 
<< m1 >>
rect 140 117 141 118 
<< m2 >>
rect 140 117 141 118 
<< m2c >>
rect 140 117 141 118 
<< m1 >>
rect 140 117 141 118 
<< m2 >>
rect 140 117 141 118 
<< m1 >>
rect 141 117 142 118 
<< m1 >>
rect 142 117 143 118 
<< m1 >>
rect 143 117 144 118 
<< m1 >>
rect 144 117 145 118 
<< m1 >>
rect 145 117 146 118 
<< m1 >>
rect 146 117 147 118 
<< m1 >>
rect 147 117 148 118 
<< m1 >>
rect 154 117 155 118 
<< m1 >>
rect 163 117 164 118 
<< m2 >>
rect 163 117 164 118 
<< m2c >>
rect 163 117 164 118 
<< m1 >>
rect 163 117 164 118 
<< m2 >>
rect 163 117 164 118 
<< m1 >>
rect 165 117 166 118 
<< m2 >>
rect 165 117 166 118 
<< m2c >>
rect 165 117 166 118 
<< m1 >>
rect 165 117 166 118 
<< m2 >>
rect 165 117 166 118 
<< m1 >>
rect 167 117 168 118 
<< m2 >>
rect 167 117 168 118 
<< m2c >>
rect 167 117 168 118 
<< m1 >>
rect 167 117 168 118 
<< m2 >>
rect 167 117 168 118 
<< m1 >>
rect 168 117 169 118 
<< m1 >>
rect 169 117 170 118 
<< m1 >>
rect 172 117 173 118 
<< m1 >>
rect 181 117 182 118 
<< m2 >>
rect 181 117 182 118 
<< m2c >>
rect 181 117 182 118 
<< m1 >>
rect 181 117 182 118 
<< m2 >>
rect 181 117 182 118 
<< m1 >>
rect 182 117 183 118 
<< m1 >>
rect 183 117 184 118 
<< m2 >>
rect 183 117 184 118 
<< m1 >>
rect 184 117 185 118 
<< m1 >>
rect 185 117 186 118 
<< m1 >>
rect 188 117 189 118 
<< m2 >>
rect 188 117 189 118 
<< m2c >>
rect 188 117 189 118 
<< m1 >>
rect 188 117 189 118 
<< m2 >>
rect 188 117 189 118 
<< m2 >>
rect 189 117 190 118 
<< m1 >>
rect 190 117 191 118 
<< m2 >>
rect 190 117 191 118 
<< m1 >>
rect 191 117 192 118 
<< m1 >>
rect 192 117 193 118 
<< m2 >>
rect 192 117 193 118 
<< m2c >>
rect 192 117 193 118 
<< m1 >>
rect 192 117 193 118 
<< m2 >>
rect 192 117 193 118 
<< m1 >>
rect 196 117 197 118 
<< m2 >>
rect 196 117 197 118 
<< m2c >>
rect 196 117 197 118 
<< m1 >>
rect 196 117 197 118 
<< m2 >>
rect 196 117 197 118 
<< m1 >>
rect 199 117 200 118 
<< m2 >>
rect 199 117 200 118 
<< m2c >>
rect 199 117 200 118 
<< m1 >>
rect 199 117 200 118 
<< m2 >>
rect 199 117 200 118 
<< m1 >>
rect 201 117 202 118 
<< m2 >>
rect 201 117 202 118 
<< m2c >>
rect 201 117 202 118 
<< m1 >>
rect 201 117 202 118 
<< m2 >>
rect 201 117 202 118 
<< m1 >>
rect 203 117 204 118 
<< m2 >>
rect 203 117 204 118 
<< m2c >>
rect 203 117 204 118 
<< m1 >>
rect 203 117 204 118 
<< m2 >>
rect 203 117 204 118 
<< m1 >>
rect 211 117 212 118 
<< m2 >>
rect 219 117 220 118 
<< m2 >>
rect 231 117 232 118 
<< m1 >>
rect 232 117 233 118 
<< m2 >>
rect 232 117 233 118 
<< m2 >>
rect 233 117 234 118 
<< m1 >>
rect 234 117 235 118 
<< m2 >>
rect 234 117 235 118 
<< m2c >>
rect 234 117 235 118 
<< m1 >>
rect 234 117 235 118 
<< m2 >>
rect 234 117 235 118 
<< m1 >>
rect 235 117 236 118 
<< m1 >>
rect 244 117 245 118 
<< m2 >>
rect 244 117 245 118 
<< m2c >>
rect 244 117 245 118 
<< m1 >>
rect 244 117 245 118 
<< m2 >>
rect 244 117 245 118 
<< m1 >>
rect 253 117 254 118 
<< m2 >>
rect 254 117 255 118 
<< m1 >>
rect 256 117 257 118 
<< m1 >>
rect 19 118 20 119 
<< m2 >>
rect 19 118 20 119 
<< m1 >>
rect 28 118 29 119 
<< m2 >>
rect 28 118 29 119 
<< m1 >>
rect 29 118 30 119 
<< m1 >>
rect 30 118 31 119 
<< m1 >>
rect 31 118 32 119 
<< m1 >>
rect 44 118 45 119 
<< m1 >>
rect 46 118 47 119 
<< m1 >>
rect 57 118 58 119 
<< m1 >>
rect 64 118 65 119 
<< m2 >>
rect 64 118 65 119 
<< m1 >>
rect 73 118 74 119 
<< m1 >>
rect 77 118 78 119 
<< m1 >>
rect 85 118 86 119 
<< m1 >>
rect 88 118 89 119 
<< m1 >>
rect 89 118 90 119 
<< m1 >>
rect 90 118 91 119 
<< m1 >>
rect 91 118 92 119 
<< m2 >>
rect 91 118 92 119 
<< m1 >>
rect 100 118 101 119 
<< m2 >>
rect 100 118 101 119 
<< m2 >>
rect 101 118 102 119 
<< m1 >>
rect 102 118 103 119 
<< m2 >>
rect 102 118 103 119 
<< m2c >>
rect 102 118 103 119 
<< m1 >>
rect 102 118 103 119 
<< m2 >>
rect 102 118 103 119 
<< m1 >>
rect 103 118 104 119 
<< m1 >>
rect 118 118 119 119 
<< m1 >>
rect 121 118 122 119 
<< m1 >>
rect 122 118 123 119 
<< m1 >>
rect 127 118 128 119 
<< m1 >>
rect 129 118 130 119 
<< m2 >>
rect 142 118 143 119 
<< m2 >>
rect 143 118 144 119 
<< m2 >>
rect 144 118 145 119 
<< m2 >>
rect 145 118 146 119 
<< m2 >>
rect 146 118 147 119 
<< m1 >>
rect 147 118 148 119 
<< m2 >>
rect 147 118 148 119 
<< m2 >>
rect 148 118 149 119 
<< m1 >>
rect 154 118 155 119 
<< m1 >>
rect 163 118 164 119 
<< m1 >>
rect 165 118 166 119 
<< m1 >>
rect 169 118 170 119 
<< m1 >>
rect 172 118 173 119 
<< m2 >>
rect 183 118 184 119 
<< m1 >>
rect 185 118 186 119 
<< m1 >>
rect 188 118 189 119 
<< m1 >>
rect 190 118 191 119 
<< m1 >>
rect 196 118 197 119 
<< m1 >>
rect 199 118 200 119 
<< m1 >>
rect 201 118 202 119 
<< m1 >>
rect 203 118 204 119 
<< m1 >>
rect 211 118 212 119 
<< m1 >>
rect 214 118 215 119 
<< m1 >>
rect 215 118 216 119 
<< m1 >>
rect 216 118 217 119 
<< m1 >>
rect 217 118 218 119 
<< m1 >>
rect 218 118 219 119 
<< m1 >>
rect 219 118 220 119 
<< m2 >>
rect 219 118 220 119 
<< m1 >>
rect 220 118 221 119 
<< m1 >>
rect 221 118 222 119 
<< m1 >>
rect 222 118 223 119 
<< m1 >>
rect 223 118 224 119 
<< m1 >>
rect 224 118 225 119 
<< m1 >>
rect 225 118 226 119 
<< m1 >>
rect 226 118 227 119 
<< m1 >>
rect 232 118 233 119 
<< m1 >>
rect 235 118 236 119 
<< m1 >>
rect 244 118 245 119 
<< m1 >>
rect 253 118 254 119 
<< m2 >>
rect 254 118 255 119 
<< m1 >>
rect 256 118 257 119 
<< m1 >>
rect 19 119 20 120 
<< m2 >>
rect 19 119 20 120 
<< m1 >>
rect 28 119 29 120 
<< m2 >>
rect 28 119 29 120 
<< m1 >>
rect 31 119 32 120 
<< m1 >>
rect 44 119 45 120 
<< m1 >>
rect 46 119 47 120 
<< m1 >>
rect 57 119 58 120 
<< m1 >>
rect 64 119 65 120 
<< m2 >>
rect 64 119 65 120 
<< m1 >>
rect 73 119 74 120 
<< m1 >>
rect 77 119 78 120 
<< m1 >>
rect 85 119 86 120 
<< m1 >>
rect 88 119 89 120 
<< m1 >>
rect 91 119 92 120 
<< m2 >>
rect 91 119 92 120 
<< m1 >>
rect 100 119 101 120 
<< m1 >>
rect 103 119 104 120 
<< m1 >>
rect 118 119 119 120 
<< m1 >>
rect 121 119 122 120 
<< m1 >>
rect 127 119 128 120 
<< m1 >>
rect 129 119 130 120 
<< m1 >>
rect 142 119 143 120 
<< m2 >>
rect 142 119 143 120 
<< m2c >>
rect 142 119 143 120 
<< m1 >>
rect 142 119 143 120 
<< m2 >>
rect 142 119 143 120 
<< m1 >>
rect 147 119 148 120 
<< m2 >>
rect 148 119 149 120 
<< m1 >>
rect 154 119 155 120 
<< m1 >>
rect 163 119 164 120 
<< m1 >>
rect 165 119 166 120 
<< m1 >>
rect 169 119 170 120 
<< m1 >>
rect 172 119 173 120 
<< m1 >>
rect 183 119 184 120 
<< m2 >>
rect 183 119 184 120 
<< m2c >>
rect 183 119 184 120 
<< m1 >>
rect 183 119 184 120 
<< m2 >>
rect 183 119 184 120 
<< m1 >>
rect 185 119 186 120 
<< m1 >>
rect 188 119 189 120 
<< m1 >>
rect 190 119 191 120 
<< m1 >>
rect 196 119 197 120 
<< m1 >>
rect 199 119 200 120 
<< m2 >>
rect 200 119 201 120 
<< m1 >>
rect 201 119 202 120 
<< m2 >>
rect 201 119 202 120 
<< m2c >>
rect 201 119 202 120 
<< m1 >>
rect 201 119 202 120 
<< m2 >>
rect 201 119 202 120 
<< m1 >>
rect 203 119 204 120 
<< m1 >>
rect 211 119 212 120 
<< m1 >>
rect 214 119 215 120 
<< m2 >>
rect 219 119 220 120 
<< m2 >>
rect 220 119 221 120 
<< m2 >>
rect 221 119 222 120 
<< m2 >>
rect 222 119 223 120 
<< m2 >>
rect 223 119 224 120 
<< m2 >>
rect 224 119 225 120 
<< m2 >>
rect 225 119 226 120 
<< m1 >>
rect 226 119 227 120 
<< m2 >>
rect 226 119 227 120 
<< m1 >>
rect 232 119 233 120 
<< m1 >>
rect 235 119 236 120 
<< m1 >>
rect 236 119 237 120 
<< m1 >>
rect 237 119 238 120 
<< m1 >>
rect 238 119 239 120 
<< m1 >>
rect 239 119 240 120 
<< m1 >>
rect 240 119 241 120 
<< m1 >>
rect 241 119 242 120 
<< m1 >>
rect 242 119 243 120 
<< m2 >>
rect 242 119 243 120 
<< m2c >>
rect 242 119 243 120 
<< m1 >>
rect 242 119 243 120 
<< m2 >>
rect 242 119 243 120 
<< m2 >>
rect 243 119 244 120 
<< m1 >>
rect 244 119 245 120 
<< m1 >>
rect 253 119 254 120 
<< m2 >>
rect 254 119 255 120 
<< m1 >>
rect 256 119 257 120 
<< pdiffusion >>
rect 12 120 13 121 
<< pdiffusion >>
rect 13 120 14 121 
<< pdiffusion >>
rect 14 120 15 121 
<< pdiffusion >>
rect 15 120 16 121 
<< pdiffusion >>
rect 16 120 17 121 
<< pdiffusion >>
rect 17 120 18 121 
<< m1 >>
rect 19 120 20 121 
<< m2 >>
rect 19 120 20 121 
<< m1 >>
rect 28 120 29 121 
<< m2 >>
rect 28 120 29 121 
<< pdiffusion >>
rect 30 120 31 121 
<< m1 >>
rect 31 120 32 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< m1 >>
rect 44 120 45 121 
<< m1 >>
rect 46 120 47 121 
<< pdiffusion >>
rect 48 120 49 121 
<< pdiffusion >>
rect 49 120 50 121 
<< pdiffusion >>
rect 50 120 51 121 
<< pdiffusion >>
rect 51 120 52 121 
<< pdiffusion >>
rect 52 120 53 121 
<< pdiffusion >>
rect 53 120 54 121 
<< m1 >>
rect 57 120 58 121 
<< m1 >>
rect 64 120 65 121 
<< m2 >>
rect 64 120 65 121 
<< pdiffusion >>
rect 66 120 67 121 
<< pdiffusion >>
rect 67 120 68 121 
<< pdiffusion >>
rect 68 120 69 121 
<< pdiffusion >>
rect 69 120 70 121 
<< pdiffusion >>
rect 70 120 71 121 
<< pdiffusion >>
rect 71 120 72 121 
<< m1 >>
rect 73 120 74 121 
<< m1 >>
rect 77 120 78 121 
<< pdiffusion >>
rect 84 120 85 121 
<< m1 >>
rect 85 120 86 121 
<< pdiffusion >>
rect 85 120 86 121 
<< pdiffusion >>
rect 86 120 87 121 
<< pdiffusion >>
rect 87 120 88 121 
<< m1 >>
rect 88 120 89 121 
<< pdiffusion >>
rect 88 120 89 121 
<< pdiffusion >>
rect 89 120 90 121 
<< m1 >>
rect 91 120 92 121 
<< m2 >>
rect 91 120 92 121 
<< m1 >>
rect 100 120 101 121 
<< pdiffusion >>
rect 102 120 103 121 
<< m1 >>
rect 103 120 104 121 
<< pdiffusion >>
rect 103 120 104 121 
<< pdiffusion >>
rect 104 120 105 121 
<< pdiffusion >>
rect 105 120 106 121 
<< pdiffusion >>
rect 106 120 107 121 
<< pdiffusion >>
rect 107 120 108 121 
<< m1 >>
rect 118 120 119 121 
<< pdiffusion >>
rect 120 120 121 121 
<< m1 >>
rect 121 120 122 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< m1 >>
rect 127 120 128 121 
<< m1 >>
rect 129 120 130 121 
<< pdiffusion >>
rect 138 120 139 121 
<< pdiffusion >>
rect 139 120 140 121 
<< pdiffusion >>
rect 140 120 141 121 
<< pdiffusion >>
rect 141 120 142 121 
<< m1 >>
rect 142 120 143 121 
<< pdiffusion >>
rect 142 120 143 121 
<< pdiffusion >>
rect 143 120 144 121 
<< m1 >>
rect 147 120 148 121 
<< m2 >>
rect 148 120 149 121 
<< m1 >>
rect 154 120 155 121 
<< pdiffusion >>
rect 156 120 157 121 
<< pdiffusion >>
rect 157 120 158 121 
<< pdiffusion >>
rect 158 120 159 121 
<< pdiffusion >>
rect 159 120 160 121 
<< pdiffusion >>
rect 160 120 161 121 
<< pdiffusion >>
rect 161 120 162 121 
<< m1 >>
rect 163 120 164 121 
<< m1 >>
rect 165 120 166 121 
<< m1 >>
rect 169 120 170 121 
<< m1 >>
rect 172 120 173 121 
<< pdiffusion >>
rect 174 120 175 121 
<< pdiffusion >>
rect 175 120 176 121 
<< pdiffusion >>
rect 176 120 177 121 
<< pdiffusion >>
rect 177 120 178 121 
<< pdiffusion >>
rect 178 120 179 121 
<< pdiffusion >>
rect 179 120 180 121 
<< m1 >>
rect 183 120 184 121 
<< m1 >>
rect 185 120 186 121 
<< m1 >>
rect 188 120 189 121 
<< m1 >>
rect 190 120 191 121 
<< pdiffusion >>
rect 192 120 193 121 
<< pdiffusion >>
rect 193 120 194 121 
<< pdiffusion >>
rect 194 120 195 121 
<< pdiffusion >>
rect 195 120 196 121 
<< m1 >>
rect 196 120 197 121 
<< pdiffusion >>
rect 196 120 197 121 
<< pdiffusion >>
rect 197 120 198 121 
<< m1 >>
rect 199 120 200 121 
<< m2 >>
rect 200 120 201 121 
<< m1 >>
rect 203 120 204 121 
<< pdiffusion >>
rect 210 120 211 121 
<< m1 >>
rect 211 120 212 121 
<< pdiffusion >>
rect 211 120 212 121 
<< pdiffusion >>
rect 212 120 213 121 
<< pdiffusion >>
rect 213 120 214 121 
<< m1 >>
rect 214 120 215 121 
<< pdiffusion >>
rect 214 120 215 121 
<< pdiffusion >>
rect 215 120 216 121 
<< m1 >>
rect 226 120 227 121 
<< m2 >>
rect 226 120 227 121 
<< pdiffusion >>
rect 228 120 229 121 
<< pdiffusion >>
rect 229 120 230 121 
<< pdiffusion >>
rect 230 120 231 121 
<< pdiffusion >>
rect 231 120 232 121 
<< m1 >>
rect 232 120 233 121 
<< pdiffusion >>
rect 232 120 233 121 
<< pdiffusion >>
rect 233 120 234 121 
<< m2 >>
rect 243 120 244 121 
<< m1 >>
rect 244 120 245 121 
<< pdiffusion >>
rect 246 120 247 121 
<< pdiffusion >>
rect 247 120 248 121 
<< pdiffusion >>
rect 248 120 249 121 
<< pdiffusion >>
rect 249 120 250 121 
<< pdiffusion >>
rect 250 120 251 121 
<< pdiffusion >>
rect 251 120 252 121 
<< m1 >>
rect 253 120 254 121 
<< m2 >>
rect 254 120 255 121 
<< m1 >>
rect 256 120 257 121 
<< pdiffusion >>
rect 12 121 13 122 
<< pdiffusion >>
rect 13 121 14 122 
<< pdiffusion >>
rect 14 121 15 122 
<< pdiffusion >>
rect 15 121 16 122 
<< pdiffusion >>
rect 16 121 17 122 
<< pdiffusion >>
rect 17 121 18 122 
<< m1 >>
rect 19 121 20 122 
<< m2 >>
rect 19 121 20 122 
<< m1 >>
rect 28 121 29 122 
<< m2 >>
rect 28 121 29 122 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< m1 >>
rect 44 121 45 122 
<< m1 >>
rect 46 121 47 122 
<< pdiffusion >>
rect 48 121 49 122 
<< pdiffusion >>
rect 49 121 50 122 
<< pdiffusion >>
rect 50 121 51 122 
<< pdiffusion >>
rect 51 121 52 122 
<< pdiffusion >>
rect 52 121 53 122 
<< pdiffusion >>
rect 53 121 54 122 
<< m1 >>
rect 57 121 58 122 
<< m1 >>
rect 64 121 65 122 
<< m2 >>
rect 64 121 65 122 
<< pdiffusion >>
rect 66 121 67 122 
<< pdiffusion >>
rect 67 121 68 122 
<< pdiffusion >>
rect 68 121 69 122 
<< pdiffusion >>
rect 69 121 70 122 
<< pdiffusion >>
rect 70 121 71 122 
<< pdiffusion >>
rect 71 121 72 122 
<< m1 >>
rect 73 121 74 122 
<< m1 >>
rect 77 121 78 122 
<< pdiffusion >>
rect 84 121 85 122 
<< pdiffusion >>
rect 85 121 86 122 
<< pdiffusion >>
rect 86 121 87 122 
<< pdiffusion >>
rect 87 121 88 122 
<< pdiffusion >>
rect 88 121 89 122 
<< pdiffusion >>
rect 89 121 90 122 
<< m1 >>
rect 91 121 92 122 
<< m2 >>
rect 91 121 92 122 
<< m1 >>
rect 100 121 101 122 
<< pdiffusion >>
rect 102 121 103 122 
<< pdiffusion >>
rect 103 121 104 122 
<< pdiffusion >>
rect 104 121 105 122 
<< pdiffusion >>
rect 105 121 106 122 
<< pdiffusion >>
rect 106 121 107 122 
<< pdiffusion >>
rect 107 121 108 122 
<< m1 >>
rect 118 121 119 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< m1 >>
rect 127 121 128 122 
<< m1 >>
rect 129 121 130 122 
<< pdiffusion >>
rect 138 121 139 122 
<< pdiffusion >>
rect 139 121 140 122 
<< pdiffusion >>
rect 140 121 141 122 
<< pdiffusion >>
rect 141 121 142 122 
<< pdiffusion >>
rect 142 121 143 122 
<< pdiffusion >>
rect 143 121 144 122 
<< m1 >>
rect 147 121 148 122 
<< m2 >>
rect 148 121 149 122 
<< m1 >>
rect 154 121 155 122 
<< pdiffusion >>
rect 156 121 157 122 
<< pdiffusion >>
rect 157 121 158 122 
<< pdiffusion >>
rect 158 121 159 122 
<< pdiffusion >>
rect 159 121 160 122 
<< pdiffusion >>
rect 160 121 161 122 
<< pdiffusion >>
rect 161 121 162 122 
<< m1 >>
rect 163 121 164 122 
<< m1 >>
rect 165 121 166 122 
<< m1 >>
rect 169 121 170 122 
<< m1 >>
rect 172 121 173 122 
<< pdiffusion >>
rect 174 121 175 122 
<< pdiffusion >>
rect 175 121 176 122 
<< pdiffusion >>
rect 176 121 177 122 
<< pdiffusion >>
rect 177 121 178 122 
<< pdiffusion >>
rect 178 121 179 122 
<< pdiffusion >>
rect 179 121 180 122 
<< m1 >>
rect 183 121 184 122 
<< m1 >>
rect 185 121 186 122 
<< m1 >>
rect 188 121 189 122 
<< m1 >>
rect 190 121 191 122 
<< pdiffusion >>
rect 192 121 193 122 
<< pdiffusion >>
rect 193 121 194 122 
<< pdiffusion >>
rect 194 121 195 122 
<< pdiffusion >>
rect 195 121 196 122 
<< pdiffusion >>
rect 196 121 197 122 
<< pdiffusion >>
rect 197 121 198 122 
<< m1 >>
rect 199 121 200 122 
<< m2 >>
rect 200 121 201 122 
<< m1 >>
rect 203 121 204 122 
<< pdiffusion >>
rect 210 121 211 122 
<< pdiffusion >>
rect 211 121 212 122 
<< pdiffusion >>
rect 212 121 213 122 
<< pdiffusion >>
rect 213 121 214 122 
<< pdiffusion >>
rect 214 121 215 122 
<< pdiffusion >>
rect 215 121 216 122 
<< m1 >>
rect 226 121 227 122 
<< m2 >>
rect 226 121 227 122 
<< pdiffusion >>
rect 228 121 229 122 
<< pdiffusion >>
rect 229 121 230 122 
<< pdiffusion >>
rect 230 121 231 122 
<< pdiffusion >>
rect 231 121 232 122 
<< pdiffusion >>
rect 232 121 233 122 
<< pdiffusion >>
rect 233 121 234 122 
<< m2 >>
rect 243 121 244 122 
<< m1 >>
rect 244 121 245 122 
<< pdiffusion >>
rect 246 121 247 122 
<< pdiffusion >>
rect 247 121 248 122 
<< pdiffusion >>
rect 248 121 249 122 
<< pdiffusion >>
rect 249 121 250 122 
<< pdiffusion >>
rect 250 121 251 122 
<< pdiffusion >>
rect 251 121 252 122 
<< m1 >>
rect 253 121 254 122 
<< m2 >>
rect 254 121 255 122 
<< m1 >>
rect 256 121 257 122 
<< pdiffusion >>
rect 12 122 13 123 
<< pdiffusion >>
rect 13 122 14 123 
<< pdiffusion >>
rect 14 122 15 123 
<< pdiffusion >>
rect 15 122 16 123 
<< pdiffusion >>
rect 16 122 17 123 
<< pdiffusion >>
rect 17 122 18 123 
<< m1 >>
rect 19 122 20 123 
<< m2 >>
rect 19 122 20 123 
<< m1 >>
rect 28 122 29 123 
<< m2 >>
rect 28 122 29 123 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< m1 >>
rect 44 122 45 123 
<< m1 >>
rect 46 122 47 123 
<< pdiffusion >>
rect 48 122 49 123 
<< pdiffusion >>
rect 49 122 50 123 
<< pdiffusion >>
rect 50 122 51 123 
<< pdiffusion >>
rect 51 122 52 123 
<< pdiffusion >>
rect 52 122 53 123 
<< pdiffusion >>
rect 53 122 54 123 
<< m1 >>
rect 57 122 58 123 
<< m1 >>
rect 64 122 65 123 
<< m2 >>
rect 64 122 65 123 
<< pdiffusion >>
rect 66 122 67 123 
<< pdiffusion >>
rect 67 122 68 123 
<< pdiffusion >>
rect 68 122 69 123 
<< pdiffusion >>
rect 69 122 70 123 
<< pdiffusion >>
rect 70 122 71 123 
<< pdiffusion >>
rect 71 122 72 123 
<< m1 >>
rect 73 122 74 123 
<< m1 >>
rect 77 122 78 123 
<< pdiffusion >>
rect 84 122 85 123 
<< pdiffusion >>
rect 85 122 86 123 
<< pdiffusion >>
rect 86 122 87 123 
<< pdiffusion >>
rect 87 122 88 123 
<< pdiffusion >>
rect 88 122 89 123 
<< pdiffusion >>
rect 89 122 90 123 
<< m1 >>
rect 91 122 92 123 
<< m2 >>
rect 91 122 92 123 
<< m1 >>
rect 100 122 101 123 
<< pdiffusion >>
rect 102 122 103 123 
<< pdiffusion >>
rect 103 122 104 123 
<< pdiffusion >>
rect 104 122 105 123 
<< pdiffusion >>
rect 105 122 106 123 
<< pdiffusion >>
rect 106 122 107 123 
<< pdiffusion >>
rect 107 122 108 123 
<< m1 >>
rect 118 122 119 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< m1 >>
rect 127 122 128 123 
<< m1 >>
rect 129 122 130 123 
<< pdiffusion >>
rect 138 122 139 123 
<< pdiffusion >>
rect 139 122 140 123 
<< pdiffusion >>
rect 140 122 141 123 
<< pdiffusion >>
rect 141 122 142 123 
<< pdiffusion >>
rect 142 122 143 123 
<< pdiffusion >>
rect 143 122 144 123 
<< m1 >>
rect 147 122 148 123 
<< m2 >>
rect 148 122 149 123 
<< m1 >>
rect 154 122 155 123 
<< pdiffusion >>
rect 156 122 157 123 
<< pdiffusion >>
rect 157 122 158 123 
<< pdiffusion >>
rect 158 122 159 123 
<< pdiffusion >>
rect 159 122 160 123 
<< pdiffusion >>
rect 160 122 161 123 
<< pdiffusion >>
rect 161 122 162 123 
<< m1 >>
rect 163 122 164 123 
<< m1 >>
rect 165 122 166 123 
<< m1 >>
rect 169 122 170 123 
<< m1 >>
rect 172 122 173 123 
<< pdiffusion >>
rect 174 122 175 123 
<< pdiffusion >>
rect 175 122 176 123 
<< pdiffusion >>
rect 176 122 177 123 
<< pdiffusion >>
rect 177 122 178 123 
<< pdiffusion >>
rect 178 122 179 123 
<< pdiffusion >>
rect 179 122 180 123 
<< m1 >>
rect 183 122 184 123 
<< m1 >>
rect 185 122 186 123 
<< m1 >>
rect 188 122 189 123 
<< m1 >>
rect 190 122 191 123 
<< pdiffusion >>
rect 192 122 193 123 
<< pdiffusion >>
rect 193 122 194 123 
<< pdiffusion >>
rect 194 122 195 123 
<< pdiffusion >>
rect 195 122 196 123 
<< pdiffusion >>
rect 196 122 197 123 
<< pdiffusion >>
rect 197 122 198 123 
<< m1 >>
rect 199 122 200 123 
<< m2 >>
rect 200 122 201 123 
<< m1 >>
rect 203 122 204 123 
<< pdiffusion >>
rect 210 122 211 123 
<< pdiffusion >>
rect 211 122 212 123 
<< pdiffusion >>
rect 212 122 213 123 
<< pdiffusion >>
rect 213 122 214 123 
<< pdiffusion >>
rect 214 122 215 123 
<< pdiffusion >>
rect 215 122 216 123 
<< m1 >>
rect 226 122 227 123 
<< m2 >>
rect 226 122 227 123 
<< pdiffusion >>
rect 228 122 229 123 
<< pdiffusion >>
rect 229 122 230 123 
<< pdiffusion >>
rect 230 122 231 123 
<< pdiffusion >>
rect 231 122 232 123 
<< pdiffusion >>
rect 232 122 233 123 
<< pdiffusion >>
rect 233 122 234 123 
<< m2 >>
rect 243 122 244 123 
<< m1 >>
rect 244 122 245 123 
<< pdiffusion >>
rect 246 122 247 123 
<< pdiffusion >>
rect 247 122 248 123 
<< pdiffusion >>
rect 248 122 249 123 
<< pdiffusion >>
rect 249 122 250 123 
<< pdiffusion >>
rect 250 122 251 123 
<< pdiffusion >>
rect 251 122 252 123 
<< m1 >>
rect 253 122 254 123 
<< m2 >>
rect 254 122 255 123 
<< m1 >>
rect 256 122 257 123 
<< pdiffusion >>
rect 12 123 13 124 
<< pdiffusion >>
rect 13 123 14 124 
<< pdiffusion >>
rect 14 123 15 124 
<< pdiffusion >>
rect 15 123 16 124 
<< pdiffusion >>
rect 16 123 17 124 
<< pdiffusion >>
rect 17 123 18 124 
<< m1 >>
rect 19 123 20 124 
<< m2 >>
rect 19 123 20 124 
<< m1 >>
rect 28 123 29 124 
<< m2 >>
rect 28 123 29 124 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< m1 >>
rect 44 123 45 124 
<< m1 >>
rect 46 123 47 124 
<< pdiffusion >>
rect 48 123 49 124 
<< pdiffusion >>
rect 49 123 50 124 
<< pdiffusion >>
rect 50 123 51 124 
<< pdiffusion >>
rect 51 123 52 124 
<< pdiffusion >>
rect 52 123 53 124 
<< pdiffusion >>
rect 53 123 54 124 
<< m1 >>
rect 57 123 58 124 
<< m1 >>
rect 64 123 65 124 
<< m2 >>
rect 64 123 65 124 
<< pdiffusion >>
rect 66 123 67 124 
<< pdiffusion >>
rect 67 123 68 124 
<< pdiffusion >>
rect 68 123 69 124 
<< pdiffusion >>
rect 69 123 70 124 
<< pdiffusion >>
rect 70 123 71 124 
<< pdiffusion >>
rect 71 123 72 124 
<< m1 >>
rect 73 123 74 124 
<< m1 >>
rect 77 123 78 124 
<< pdiffusion >>
rect 84 123 85 124 
<< pdiffusion >>
rect 85 123 86 124 
<< pdiffusion >>
rect 86 123 87 124 
<< pdiffusion >>
rect 87 123 88 124 
<< pdiffusion >>
rect 88 123 89 124 
<< pdiffusion >>
rect 89 123 90 124 
<< m1 >>
rect 91 123 92 124 
<< m2 >>
rect 91 123 92 124 
<< m1 >>
rect 100 123 101 124 
<< pdiffusion >>
rect 102 123 103 124 
<< pdiffusion >>
rect 103 123 104 124 
<< pdiffusion >>
rect 104 123 105 124 
<< pdiffusion >>
rect 105 123 106 124 
<< pdiffusion >>
rect 106 123 107 124 
<< pdiffusion >>
rect 107 123 108 124 
<< m1 >>
rect 118 123 119 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< m1 >>
rect 127 123 128 124 
<< m1 >>
rect 129 123 130 124 
<< pdiffusion >>
rect 138 123 139 124 
<< pdiffusion >>
rect 139 123 140 124 
<< pdiffusion >>
rect 140 123 141 124 
<< pdiffusion >>
rect 141 123 142 124 
<< pdiffusion >>
rect 142 123 143 124 
<< pdiffusion >>
rect 143 123 144 124 
<< m1 >>
rect 147 123 148 124 
<< m2 >>
rect 148 123 149 124 
<< m1 >>
rect 154 123 155 124 
<< pdiffusion >>
rect 156 123 157 124 
<< pdiffusion >>
rect 157 123 158 124 
<< pdiffusion >>
rect 158 123 159 124 
<< pdiffusion >>
rect 159 123 160 124 
<< pdiffusion >>
rect 160 123 161 124 
<< pdiffusion >>
rect 161 123 162 124 
<< m1 >>
rect 163 123 164 124 
<< m1 >>
rect 165 123 166 124 
<< m1 >>
rect 169 123 170 124 
<< m1 >>
rect 172 123 173 124 
<< pdiffusion >>
rect 174 123 175 124 
<< pdiffusion >>
rect 175 123 176 124 
<< pdiffusion >>
rect 176 123 177 124 
<< pdiffusion >>
rect 177 123 178 124 
<< pdiffusion >>
rect 178 123 179 124 
<< pdiffusion >>
rect 179 123 180 124 
<< m1 >>
rect 183 123 184 124 
<< m1 >>
rect 185 123 186 124 
<< m1 >>
rect 188 123 189 124 
<< m1 >>
rect 190 123 191 124 
<< pdiffusion >>
rect 192 123 193 124 
<< pdiffusion >>
rect 193 123 194 124 
<< pdiffusion >>
rect 194 123 195 124 
<< pdiffusion >>
rect 195 123 196 124 
<< pdiffusion >>
rect 196 123 197 124 
<< pdiffusion >>
rect 197 123 198 124 
<< m1 >>
rect 199 123 200 124 
<< m2 >>
rect 200 123 201 124 
<< m1 >>
rect 203 123 204 124 
<< pdiffusion >>
rect 210 123 211 124 
<< pdiffusion >>
rect 211 123 212 124 
<< pdiffusion >>
rect 212 123 213 124 
<< pdiffusion >>
rect 213 123 214 124 
<< pdiffusion >>
rect 214 123 215 124 
<< pdiffusion >>
rect 215 123 216 124 
<< m1 >>
rect 226 123 227 124 
<< m2 >>
rect 226 123 227 124 
<< pdiffusion >>
rect 228 123 229 124 
<< pdiffusion >>
rect 229 123 230 124 
<< pdiffusion >>
rect 230 123 231 124 
<< pdiffusion >>
rect 231 123 232 124 
<< pdiffusion >>
rect 232 123 233 124 
<< pdiffusion >>
rect 233 123 234 124 
<< m2 >>
rect 243 123 244 124 
<< m1 >>
rect 244 123 245 124 
<< pdiffusion >>
rect 246 123 247 124 
<< pdiffusion >>
rect 247 123 248 124 
<< pdiffusion >>
rect 248 123 249 124 
<< pdiffusion >>
rect 249 123 250 124 
<< pdiffusion >>
rect 250 123 251 124 
<< pdiffusion >>
rect 251 123 252 124 
<< m1 >>
rect 253 123 254 124 
<< m2 >>
rect 254 123 255 124 
<< m1 >>
rect 256 123 257 124 
<< pdiffusion >>
rect 12 124 13 125 
<< pdiffusion >>
rect 13 124 14 125 
<< pdiffusion >>
rect 14 124 15 125 
<< pdiffusion >>
rect 15 124 16 125 
<< pdiffusion >>
rect 16 124 17 125 
<< pdiffusion >>
rect 17 124 18 125 
<< m1 >>
rect 19 124 20 125 
<< m2 >>
rect 19 124 20 125 
<< m1 >>
rect 28 124 29 125 
<< m2 >>
rect 28 124 29 125 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< m1 >>
rect 44 124 45 125 
<< m1 >>
rect 46 124 47 125 
<< pdiffusion >>
rect 48 124 49 125 
<< pdiffusion >>
rect 49 124 50 125 
<< pdiffusion >>
rect 50 124 51 125 
<< pdiffusion >>
rect 51 124 52 125 
<< pdiffusion >>
rect 52 124 53 125 
<< pdiffusion >>
rect 53 124 54 125 
<< m1 >>
rect 57 124 58 125 
<< m1 >>
rect 64 124 65 125 
<< m2 >>
rect 64 124 65 125 
<< pdiffusion >>
rect 66 124 67 125 
<< pdiffusion >>
rect 67 124 68 125 
<< pdiffusion >>
rect 68 124 69 125 
<< pdiffusion >>
rect 69 124 70 125 
<< pdiffusion >>
rect 70 124 71 125 
<< pdiffusion >>
rect 71 124 72 125 
<< m1 >>
rect 73 124 74 125 
<< m1 >>
rect 77 124 78 125 
<< pdiffusion >>
rect 84 124 85 125 
<< pdiffusion >>
rect 85 124 86 125 
<< pdiffusion >>
rect 86 124 87 125 
<< pdiffusion >>
rect 87 124 88 125 
<< pdiffusion >>
rect 88 124 89 125 
<< pdiffusion >>
rect 89 124 90 125 
<< m1 >>
rect 91 124 92 125 
<< m2 >>
rect 91 124 92 125 
<< m1 >>
rect 100 124 101 125 
<< pdiffusion >>
rect 102 124 103 125 
<< pdiffusion >>
rect 103 124 104 125 
<< pdiffusion >>
rect 104 124 105 125 
<< pdiffusion >>
rect 105 124 106 125 
<< pdiffusion >>
rect 106 124 107 125 
<< pdiffusion >>
rect 107 124 108 125 
<< m1 >>
rect 118 124 119 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< m1 >>
rect 127 124 128 125 
<< m1 >>
rect 129 124 130 125 
<< pdiffusion >>
rect 138 124 139 125 
<< pdiffusion >>
rect 139 124 140 125 
<< pdiffusion >>
rect 140 124 141 125 
<< pdiffusion >>
rect 141 124 142 125 
<< pdiffusion >>
rect 142 124 143 125 
<< pdiffusion >>
rect 143 124 144 125 
<< m1 >>
rect 147 124 148 125 
<< m2 >>
rect 148 124 149 125 
<< m1 >>
rect 154 124 155 125 
<< pdiffusion >>
rect 156 124 157 125 
<< pdiffusion >>
rect 157 124 158 125 
<< pdiffusion >>
rect 158 124 159 125 
<< pdiffusion >>
rect 159 124 160 125 
<< pdiffusion >>
rect 160 124 161 125 
<< pdiffusion >>
rect 161 124 162 125 
<< m1 >>
rect 163 124 164 125 
<< m1 >>
rect 165 124 166 125 
<< m1 >>
rect 169 124 170 125 
<< m1 >>
rect 172 124 173 125 
<< pdiffusion >>
rect 174 124 175 125 
<< pdiffusion >>
rect 175 124 176 125 
<< pdiffusion >>
rect 176 124 177 125 
<< pdiffusion >>
rect 177 124 178 125 
<< pdiffusion >>
rect 178 124 179 125 
<< pdiffusion >>
rect 179 124 180 125 
<< m1 >>
rect 183 124 184 125 
<< m1 >>
rect 185 124 186 125 
<< m1 >>
rect 188 124 189 125 
<< m1 >>
rect 190 124 191 125 
<< pdiffusion >>
rect 192 124 193 125 
<< pdiffusion >>
rect 193 124 194 125 
<< pdiffusion >>
rect 194 124 195 125 
<< pdiffusion >>
rect 195 124 196 125 
<< pdiffusion >>
rect 196 124 197 125 
<< pdiffusion >>
rect 197 124 198 125 
<< m1 >>
rect 199 124 200 125 
<< m2 >>
rect 200 124 201 125 
<< m1 >>
rect 203 124 204 125 
<< pdiffusion >>
rect 210 124 211 125 
<< pdiffusion >>
rect 211 124 212 125 
<< pdiffusion >>
rect 212 124 213 125 
<< pdiffusion >>
rect 213 124 214 125 
<< pdiffusion >>
rect 214 124 215 125 
<< pdiffusion >>
rect 215 124 216 125 
<< m1 >>
rect 226 124 227 125 
<< m2 >>
rect 226 124 227 125 
<< pdiffusion >>
rect 228 124 229 125 
<< pdiffusion >>
rect 229 124 230 125 
<< pdiffusion >>
rect 230 124 231 125 
<< pdiffusion >>
rect 231 124 232 125 
<< pdiffusion >>
rect 232 124 233 125 
<< pdiffusion >>
rect 233 124 234 125 
<< m2 >>
rect 243 124 244 125 
<< m1 >>
rect 244 124 245 125 
<< pdiffusion >>
rect 246 124 247 125 
<< pdiffusion >>
rect 247 124 248 125 
<< pdiffusion >>
rect 248 124 249 125 
<< pdiffusion >>
rect 249 124 250 125 
<< pdiffusion >>
rect 250 124 251 125 
<< pdiffusion >>
rect 251 124 252 125 
<< m1 >>
rect 253 124 254 125 
<< m2 >>
rect 254 124 255 125 
<< m1 >>
rect 256 124 257 125 
<< pdiffusion >>
rect 12 125 13 126 
<< pdiffusion >>
rect 13 125 14 126 
<< pdiffusion >>
rect 14 125 15 126 
<< pdiffusion >>
rect 15 125 16 126 
<< m1 >>
rect 16 125 17 126 
<< pdiffusion >>
rect 16 125 17 126 
<< pdiffusion >>
rect 17 125 18 126 
<< m1 >>
rect 19 125 20 126 
<< m2 >>
rect 19 125 20 126 
<< m1 >>
rect 28 125 29 126 
<< m2 >>
rect 28 125 29 126 
<< pdiffusion >>
rect 30 125 31 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< m1 >>
rect 44 125 45 126 
<< m1 >>
rect 46 125 47 126 
<< pdiffusion >>
rect 48 125 49 126 
<< pdiffusion >>
rect 49 125 50 126 
<< pdiffusion >>
rect 50 125 51 126 
<< pdiffusion >>
rect 51 125 52 126 
<< m1 >>
rect 52 125 53 126 
<< pdiffusion >>
rect 52 125 53 126 
<< pdiffusion >>
rect 53 125 54 126 
<< m1 >>
rect 57 125 58 126 
<< m1 >>
rect 64 125 65 126 
<< m2 >>
rect 64 125 65 126 
<< pdiffusion >>
rect 66 125 67 126 
<< m1 >>
rect 67 125 68 126 
<< pdiffusion >>
rect 67 125 68 126 
<< pdiffusion >>
rect 68 125 69 126 
<< pdiffusion >>
rect 69 125 70 126 
<< pdiffusion >>
rect 70 125 71 126 
<< pdiffusion >>
rect 71 125 72 126 
<< m1 >>
rect 73 125 74 126 
<< m1 >>
rect 77 125 78 126 
<< pdiffusion >>
rect 84 125 85 126 
<< pdiffusion >>
rect 85 125 86 126 
<< pdiffusion >>
rect 86 125 87 126 
<< pdiffusion >>
rect 87 125 88 126 
<< pdiffusion >>
rect 88 125 89 126 
<< pdiffusion >>
rect 89 125 90 126 
<< m1 >>
rect 91 125 92 126 
<< m2 >>
rect 91 125 92 126 
<< m1 >>
rect 100 125 101 126 
<< pdiffusion >>
rect 102 125 103 126 
<< pdiffusion >>
rect 103 125 104 126 
<< pdiffusion >>
rect 104 125 105 126 
<< pdiffusion >>
rect 105 125 106 126 
<< pdiffusion >>
rect 106 125 107 126 
<< pdiffusion >>
rect 107 125 108 126 
<< m1 >>
rect 118 125 119 126 
<< pdiffusion >>
rect 120 125 121 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< m1 >>
rect 127 125 128 126 
<< m1 >>
rect 129 125 130 126 
<< pdiffusion >>
rect 138 125 139 126 
<< m1 >>
rect 139 125 140 126 
<< pdiffusion >>
rect 139 125 140 126 
<< pdiffusion >>
rect 140 125 141 126 
<< pdiffusion >>
rect 141 125 142 126 
<< pdiffusion >>
rect 142 125 143 126 
<< pdiffusion >>
rect 143 125 144 126 
<< m1 >>
rect 147 125 148 126 
<< m2 >>
rect 148 125 149 126 
<< m1 >>
rect 154 125 155 126 
<< pdiffusion >>
rect 156 125 157 126 
<< m1 >>
rect 157 125 158 126 
<< pdiffusion >>
rect 157 125 158 126 
<< pdiffusion >>
rect 158 125 159 126 
<< pdiffusion >>
rect 159 125 160 126 
<< pdiffusion >>
rect 160 125 161 126 
<< pdiffusion >>
rect 161 125 162 126 
<< m1 >>
rect 163 125 164 126 
<< m1 >>
rect 165 125 166 126 
<< m1 >>
rect 169 125 170 126 
<< m1 >>
rect 172 125 173 126 
<< pdiffusion >>
rect 174 125 175 126 
<< m1 >>
rect 175 125 176 126 
<< pdiffusion >>
rect 175 125 176 126 
<< pdiffusion >>
rect 176 125 177 126 
<< pdiffusion >>
rect 177 125 178 126 
<< pdiffusion >>
rect 178 125 179 126 
<< pdiffusion >>
rect 179 125 180 126 
<< m1 >>
rect 183 125 184 126 
<< m1 >>
rect 185 125 186 126 
<< m1 >>
rect 188 125 189 126 
<< m1 >>
rect 190 125 191 126 
<< pdiffusion >>
rect 192 125 193 126 
<< m1 >>
rect 193 125 194 126 
<< pdiffusion >>
rect 193 125 194 126 
<< pdiffusion >>
rect 194 125 195 126 
<< pdiffusion >>
rect 195 125 196 126 
<< m1 >>
rect 196 125 197 126 
<< pdiffusion >>
rect 196 125 197 126 
<< pdiffusion >>
rect 197 125 198 126 
<< m1 >>
rect 199 125 200 126 
<< m2 >>
rect 200 125 201 126 
<< m1 >>
rect 203 125 204 126 
<< pdiffusion >>
rect 210 125 211 126 
<< pdiffusion >>
rect 211 125 212 126 
<< pdiffusion >>
rect 212 125 213 126 
<< pdiffusion >>
rect 213 125 214 126 
<< m1 >>
rect 214 125 215 126 
<< pdiffusion >>
rect 214 125 215 126 
<< pdiffusion >>
rect 215 125 216 126 
<< m1 >>
rect 226 125 227 126 
<< m2 >>
rect 226 125 227 126 
<< pdiffusion >>
rect 228 125 229 126 
<< pdiffusion >>
rect 229 125 230 126 
<< pdiffusion >>
rect 230 125 231 126 
<< pdiffusion >>
rect 231 125 232 126 
<< pdiffusion >>
rect 232 125 233 126 
<< pdiffusion >>
rect 233 125 234 126 
<< m2 >>
rect 243 125 244 126 
<< m1 >>
rect 244 125 245 126 
<< pdiffusion >>
rect 246 125 247 126 
<< pdiffusion >>
rect 247 125 248 126 
<< pdiffusion >>
rect 248 125 249 126 
<< pdiffusion >>
rect 249 125 250 126 
<< m1 >>
rect 250 125 251 126 
<< pdiffusion >>
rect 250 125 251 126 
<< pdiffusion >>
rect 251 125 252 126 
<< m1 >>
rect 253 125 254 126 
<< m2 >>
rect 254 125 255 126 
<< m1 >>
rect 256 125 257 126 
<< m1 >>
rect 16 126 17 127 
<< m1 >>
rect 19 126 20 127 
<< m2 >>
rect 19 126 20 127 
<< m1 >>
rect 28 126 29 127 
<< m2 >>
rect 28 126 29 127 
<< m1 >>
rect 44 126 45 127 
<< m1 >>
rect 46 126 47 127 
<< m1 >>
rect 52 126 53 127 
<< m1 >>
rect 57 126 58 127 
<< m1 >>
rect 64 126 65 127 
<< m2 >>
rect 64 126 65 127 
<< m1 >>
rect 67 126 68 127 
<< m1 >>
rect 73 126 74 127 
<< m1 >>
rect 77 126 78 127 
<< m1 >>
rect 91 126 92 127 
<< m2 >>
rect 91 126 92 127 
<< m1 >>
rect 100 126 101 127 
<< m1 >>
rect 118 126 119 127 
<< m1 >>
rect 127 126 128 127 
<< m1 >>
rect 129 126 130 127 
<< m1 >>
rect 139 126 140 127 
<< m1 >>
rect 147 126 148 127 
<< m2 >>
rect 148 126 149 127 
<< m1 >>
rect 154 126 155 127 
<< m1 >>
rect 157 126 158 127 
<< m1 >>
rect 163 126 164 127 
<< m1 >>
rect 165 126 166 127 
<< m1 >>
rect 169 126 170 127 
<< m1 >>
rect 172 126 173 127 
<< m1 >>
rect 175 126 176 127 
<< m1 >>
rect 183 126 184 127 
<< m1 >>
rect 185 126 186 127 
<< m1 >>
rect 188 126 189 127 
<< m1 >>
rect 190 126 191 127 
<< m1 >>
rect 193 126 194 127 
<< m1 >>
rect 196 126 197 127 
<< m2 >>
rect 196 126 197 127 
<< m2c >>
rect 196 126 197 127 
<< m1 >>
rect 196 126 197 127 
<< m2 >>
rect 196 126 197 127 
<< m1 >>
rect 199 126 200 127 
<< m2 >>
rect 200 126 201 127 
<< m1 >>
rect 203 126 204 127 
<< m1 >>
rect 214 126 215 127 
<< m1 >>
rect 226 126 227 127 
<< m2 >>
rect 226 126 227 127 
<< m2 >>
rect 243 126 244 127 
<< m1 >>
rect 244 126 245 127 
<< m1 >>
rect 250 126 251 127 
<< m1 >>
rect 253 126 254 127 
<< m2 >>
rect 254 126 255 127 
<< m1 >>
rect 256 126 257 127 
<< m1 >>
rect 16 127 17 128 
<< m1 >>
rect 17 127 18 128 
<< m1 >>
rect 18 127 19 128 
<< m1 >>
rect 19 127 20 128 
<< m2 >>
rect 19 127 20 128 
<< m1 >>
rect 28 127 29 128 
<< m2 >>
rect 28 127 29 128 
<< m1 >>
rect 44 127 45 128 
<< m1 >>
rect 46 127 47 128 
<< m1 >>
rect 52 127 53 128 
<< m1 >>
rect 57 127 58 128 
<< m1 >>
rect 64 127 65 128 
<< m2 >>
rect 64 127 65 128 
<< m1 >>
rect 67 127 68 128 
<< m1 >>
rect 73 127 74 128 
<< m1 >>
rect 77 127 78 128 
<< m1 >>
rect 91 127 92 128 
<< m2 >>
rect 91 127 92 128 
<< m1 >>
rect 100 127 101 128 
<< m1 >>
rect 118 127 119 128 
<< m1 >>
rect 127 127 128 128 
<< m1 >>
rect 129 127 130 128 
<< m1 >>
rect 139 127 140 128 
<< m1 >>
rect 147 127 148 128 
<< m2 >>
rect 148 127 149 128 
<< m1 >>
rect 154 127 155 128 
<< m1 >>
rect 155 127 156 128 
<< m1 >>
rect 156 127 157 128 
<< m1 >>
rect 157 127 158 128 
<< m1 >>
rect 163 127 164 128 
<< m1 >>
rect 165 127 166 128 
<< m1 >>
rect 169 127 170 128 
<< m1 >>
rect 172 127 173 128 
<< m1 >>
rect 173 127 174 128 
<< m1 >>
rect 174 127 175 128 
<< m1 >>
rect 175 127 176 128 
<< m1 >>
rect 179 127 180 128 
<< m1 >>
rect 180 127 181 128 
<< m1 >>
rect 181 127 182 128 
<< m1 >>
rect 182 127 183 128 
<< m1 >>
rect 183 127 184 128 
<< m1 >>
rect 185 127 186 128 
<< m2 >>
rect 185 127 186 128 
<< m2c >>
rect 185 127 186 128 
<< m1 >>
rect 185 127 186 128 
<< m2 >>
rect 185 127 186 128 
<< m1 >>
rect 188 127 189 128 
<< m1 >>
rect 190 127 191 128 
<< m1 >>
rect 193 127 194 128 
<< m2 >>
rect 196 127 197 128 
<< m2 >>
rect 197 127 198 128 
<< m2 >>
rect 198 127 199 128 
<< m1 >>
rect 199 127 200 128 
<< m2 >>
rect 199 127 200 128 
<< m2 >>
rect 200 127 201 128 
<< m1 >>
rect 203 127 204 128 
<< m1 >>
rect 214 127 215 128 
<< m1 >>
rect 226 127 227 128 
<< m2 >>
rect 226 127 227 128 
<< m2 >>
rect 243 127 244 128 
<< m1 >>
rect 244 127 245 128 
<< m2 >>
rect 244 127 245 128 
<< m2 >>
rect 245 127 246 128 
<< m1 >>
rect 246 127 247 128 
<< m2 >>
rect 246 127 247 128 
<< m2c >>
rect 246 127 247 128 
<< m1 >>
rect 246 127 247 128 
<< m2 >>
rect 246 127 247 128 
<< m1 >>
rect 250 127 251 128 
<< m1 >>
rect 253 127 254 128 
<< m2 >>
rect 254 127 255 128 
<< m1 >>
rect 256 127 257 128 
<< m2 >>
rect 19 128 20 129 
<< m1 >>
rect 28 128 29 129 
<< m2 >>
rect 28 128 29 129 
<< m1 >>
rect 44 128 45 129 
<< m1 >>
rect 46 128 47 129 
<< m1 >>
rect 52 128 53 129 
<< m1 >>
rect 57 128 58 129 
<< m1 >>
rect 64 128 65 129 
<< m2 >>
rect 64 128 65 129 
<< m1 >>
rect 67 128 68 129 
<< m1 >>
rect 68 128 69 129 
<< m1 >>
rect 69 128 70 129 
<< m1 >>
rect 70 128 71 129 
<< m1 >>
rect 71 128 72 129 
<< m2 >>
rect 71 128 72 129 
<< m2c >>
rect 71 128 72 129 
<< m1 >>
rect 71 128 72 129 
<< m2 >>
rect 71 128 72 129 
<< m2 >>
rect 72 128 73 129 
<< m1 >>
rect 73 128 74 129 
<< m2 >>
rect 73 128 74 129 
<< m2 >>
rect 74 128 75 129 
<< m1 >>
rect 75 128 76 129 
<< m2 >>
rect 75 128 76 129 
<< m2c >>
rect 75 128 76 129 
<< m1 >>
rect 75 128 76 129 
<< m2 >>
rect 75 128 76 129 
<< m2 >>
rect 76 128 77 129 
<< m1 >>
rect 77 128 78 129 
<< m2 >>
rect 77 128 78 129 
<< m2 >>
rect 78 128 79 129 
<< m1 >>
rect 79 128 80 129 
<< m2 >>
rect 79 128 80 129 
<< m2c >>
rect 79 128 80 129 
<< m1 >>
rect 79 128 80 129 
<< m2 >>
rect 79 128 80 129 
<< m1 >>
rect 91 128 92 129 
<< m2 >>
rect 91 128 92 129 
<< m1 >>
rect 100 128 101 129 
<< m2 >>
rect 100 128 101 129 
<< m2c >>
rect 100 128 101 129 
<< m1 >>
rect 100 128 101 129 
<< m2 >>
rect 100 128 101 129 
<< m1 >>
rect 118 128 119 129 
<< m1 >>
rect 122 128 123 129 
<< m2 >>
rect 122 128 123 129 
<< m2c >>
rect 122 128 123 129 
<< m1 >>
rect 122 128 123 129 
<< m2 >>
rect 122 128 123 129 
<< m1 >>
rect 123 128 124 129 
<< m1 >>
rect 124 128 125 129 
<< m1 >>
rect 125 128 126 129 
<< m1 >>
rect 126 128 127 129 
<< m1 >>
rect 127 128 128 129 
<< m1 >>
rect 129 128 130 129 
<< m2 >>
rect 129 128 130 129 
<< m2c >>
rect 129 128 130 129 
<< m1 >>
rect 129 128 130 129 
<< m2 >>
rect 129 128 130 129 
<< m1 >>
rect 131 128 132 129 
<< m2 >>
rect 131 128 132 129 
<< m2c >>
rect 131 128 132 129 
<< m1 >>
rect 131 128 132 129 
<< m2 >>
rect 131 128 132 129 
<< m1 >>
rect 132 128 133 129 
<< m1 >>
rect 133 128 134 129 
<< m1 >>
rect 134 128 135 129 
<< m1 >>
rect 135 128 136 129 
<< m1 >>
rect 136 128 137 129 
<< m1 >>
rect 137 128 138 129 
<< m1 >>
rect 138 128 139 129 
<< m1 >>
rect 139 128 140 129 
<< m1 >>
rect 147 128 148 129 
<< m2 >>
rect 148 128 149 129 
<< m1 >>
rect 163 128 164 129 
<< m1 >>
rect 165 128 166 129 
<< m1 >>
rect 169 128 170 129 
<< m2 >>
rect 169 128 170 129 
<< m2c >>
rect 169 128 170 129 
<< m1 >>
rect 169 128 170 129 
<< m2 >>
rect 169 128 170 129 
<< m1 >>
rect 177 128 178 129 
<< m2 >>
rect 177 128 178 129 
<< m2c >>
rect 177 128 178 129 
<< m1 >>
rect 177 128 178 129 
<< m2 >>
rect 177 128 178 129 
<< m1 >>
rect 178 128 179 129 
<< m1 >>
rect 179 128 180 129 
<< m2 >>
rect 185 128 186 129 
<< m1 >>
rect 188 128 189 129 
<< m1 >>
rect 190 128 191 129 
<< m1 >>
rect 193 128 194 129 
<< m1 >>
rect 194 128 195 129 
<< m1 >>
rect 195 128 196 129 
<< m1 >>
rect 196 128 197 129 
<< m1 >>
rect 197 128 198 129 
<< m1 >>
rect 198 128 199 129 
<< m1 >>
rect 199 128 200 129 
<< m1 >>
rect 203 128 204 129 
<< m1 >>
rect 214 128 215 129 
<< m1 >>
rect 226 128 227 129 
<< m2 >>
rect 226 128 227 129 
<< m1 >>
rect 244 128 245 129 
<< m1 >>
rect 246 128 247 129 
<< m1 >>
rect 250 128 251 129 
<< m1 >>
rect 253 128 254 129 
<< m2 >>
rect 254 128 255 129 
<< m1 >>
rect 256 128 257 129 
<< m1 >>
rect 19 129 20 130 
<< m2 >>
rect 19 129 20 130 
<< m2c >>
rect 19 129 20 130 
<< m1 >>
rect 19 129 20 130 
<< m2 >>
rect 19 129 20 130 
<< m1 >>
rect 28 129 29 130 
<< m2 >>
rect 28 129 29 130 
<< m1 >>
rect 44 129 45 130 
<< m1 >>
rect 46 129 47 130 
<< m1 >>
rect 52 129 53 130 
<< m1 >>
rect 57 129 58 130 
<< m1 >>
rect 64 129 65 130 
<< m2 >>
rect 64 129 65 130 
<< m1 >>
rect 73 129 74 130 
<< m1 >>
rect 77 129 78 130 
<< m1 >>
rect 79 129 80 130 
<< m1 >>
rect 91 129 92 130 
<< m2 >>
rect 91 129 92 130 
<< m2 >>
rect 100 129 101 130 
<< m1 >>
rect 118 129 119 130 
<< m2 >>
rect 122 129 123 130 
<< m2 >>
rect 129 129 130 130 
<< m2 >>
rect 131 129 132 130 
<< m1 >>
rect 147 129 148 130 
<< m2 >>
rect 148 129 149 130 
<< m1 >>
rect 163 129 164 130 
<< m1 >>
rect 165 129 166 130 
<< m2 >>
rect 169 129 170 130 
<< m2 >>
rect 177 129 178 130 
<< m2 >>
rect 182 129 183 130 
<< m1 >>
rect 183 129 184 130 
<< m2 >>
rect 183 129 184 130 
<< m2c >>
rect 183 129 184 130 
<< m1 >>
rect 183 129 184 130 
<< m2 >>
rect 183 129 184 130 
<< m1 >>
rect 184 129 185 130 
<< m1 >>
rect 185 129 186 130 
<< m2 >>
rect 185 129 186 130 
<< m1 >>
rect 186 129 187 130 
<< m1 >>
rect 187 129 188 130 
<< m1 >>
rect 188 129 189 130 
<< m1 >>
rect 190 129 191 130 
<< m2 >>
rect 196 129 197 130 
<< m2 >>
rect 197 129 198 130 
<< m2 >>
rect 198 129 199 130 
<< m2 >>
rect 199 129 200 130 
<< m2 >>
rect 200 129 201 130 
<< m1 >>
rect 201 129 202 130 
<< m2 >>
rect 201 129 202 130 
<< m2c >>
rect 201 129 202 130 
<< m1 >>
rect 201 129 202 130 
<< m2 >>
rect 201 129 202 130 
<< m1 >>
rect 202 129 203 130 
<< m1 >>
rect 203 129 204 130 
<< m1 >>
rect 214 129 215 130 
<< m1 >>
rect 226 129 227 130 
<< m2 >>
rect 226 129 227 130 
<< m1 >>
rect 244 129 245 130 
<< m1 >>
rect 246 129 247 130 
<< m1 >>
rect 250 129 251 130 
<< m1 >>
rect 253 129 254 130 
<< m2 >>
rect 254 129 255 130 
<< m1 >>
rect 256 129 257 130 
<< m1 >>
rect 19 130 20 131 
<< m1 >>
rect 28 130 29 131 
<< m2 >>
rect 28 130 29 131 
<< m1 >>
rect 34 130 35 131 
<< m1 >>
rect 35 130 36 131 
<< m1 >>
rect 36 130 37 131 
<< m1 >>
rect 37 130 38 131 
<< m1 >>
rect 38 130 39 131 
<< m1 >>
rect 39 130 40 131 
<< m1 >>
rect 40 130 41 131 
<< m1 >>
rect 41 130 42 131 
<< m1 >>
rect 42 130 43 131 
<< m2 >>
rect 42 130 43 131 
<< m2c >>
rect 42 130 43 131 
<< m1 >>
rect 42 130 43 131 
<< m2 >>
rect 42 130 43 131 
<< m2 >>
rect 43 130 44 131 
<< m1 >>
rect 44 130 45 131 
<< m2 >>
rect 44 130 45 131 
<< m2 >>
rect 45 130 46 131 
<< m1 >>
rect 46 130 47 131 
<< m2 >>
rect 46 130 47 131 
<< m2 >>
rect 47 130 48 131 
<< m1 >>
rect 48 130 49 131 
<< m2 >>
rect 48 130 49 131 
<< m2c >>
rect 48 130 49 131 
<< m1 >>
rect 48 130 49 131 
<< m2 >>
rect 48 130 49 131 
<< m1 >>
rect 49 130 50 131 
<< m1 >>
rect 50 130 51 131 
<< m1 >>
rect 51 130 52 131 
<< m1 >>
rect 52 130 53 131 
<< m1 >>
rect 57 130 58 131 
<< m1 >>
rect 64 130 65 131 
<< m2 >>
rect 64 130 65 131 
<< m1 >>
rect 73 130 74 131 
<< m1 >>
rect 77 130 78 131 
<< m1 >>
rect 79 130 80 131 
<< m1 >>
rect 91 130 92 131 
<< m2 >>
rect 91 130 92 131 
<< m1 >>
rect 92 130 93 131 
<< m1 >>
rect 93 130 94 131 
<< m1 >>
rect 94 130 95 131 
<< m1 >>
rect 95 130 96 131 
<< m1 >>
rect 96 130 97 131 
<< m1 >>
rect 97 130 98 131 
<< m1 >>
rect 98 130 99 131 
<< m1 >>
rect 99 130 100 131 
<< m1 >>
rect 100 130 101 131 
<< m2 >>
rect 100 130 101 131 
<< m1 >>
rect 101 130 102 131 
<< m1 >>
rect 102 130 103 131 
<< m1 >>
rect 103 130 104 131 
<< m1 >>
rect 104 130 105 131 
<< m1 >>
rect 105 130 106 131 
<< m1 >>
rect 106 130 107 131 
<< m1 >>
rect 107 130 108 131 
<< m1 >>
rect 108 130 109 131 
<< m1 >>
rect 109 130 110 131 
<< m1 >>
rect 110 130 111 131 
<< m1 >>
rect 111 130 112 131 
<< m1 >>
rect 112 130 113 131 
<< m1 >>
rect 113 130 114 131 
<< m1 >>
rect 114 130 115 131 
<< m1 >>
rect 115 130 116 131 
<< m1 >>
rect 116 130 117 131 
<< m2 >>
rect 116 130 117 131 
<< m2c >>
rect 116 130 117 131 
<< m1 >>
rect 116 130 117 131 
<< m2 >>
rect 116 130 117 131 
<< m2 >>
rect 117 130 118 131 
<< m1 >>
rect 118 130 119 131 
<< m2 >>
rect 118 130 119 131 
<< m2 >>
rect 119 130 120 131 
<< m1 >>
rect 120 130 121 131 
<< m2 >>
rect 120 130 121 131 
<< m2c >>
rect 120 130 121 131 
<< m1 >>
rect 120 130 121 131 
<< m2 >>
rect 120 130 121 131 
<< m1 >>
rect 121 130 122 131 
<< m1 >>
rect 122 130 123 131 
<< m2 >>
rect 122 130 123 131 
<< m1 >>
rect 123 130 124 131 
<< m1 >>
rect 124 130 125 131 
<< m1 >>
rect 125 130 126 131 
<< m1 >>
rect 126 130 127 131 
<< m1 >>
rect 127 130 128 131 
<< m1 >>
rect 128 130 129 131 
<< m1 >>
rect 129 130 130 131 
<< m2 >>
rect 129 130 130 131 
<< m1 >>
rect 130 130 131 131 
<< m1 >>
rect 131 130 132 131 
<< m2 >>
rect 131 130 132 131 
<< m1 >>
rect 132 130 133 131 
<< m1 >>
rect 133 130 134 131 
<< m1 >>
rect 134 130 135 131 
<< m1 >>
rect 135 130 136 131 
<< m1 >>
rect 136 130 137 131 
<< m1 >>
rect 137 130 138 131 
<< m1 >>
rect 138 130 139 131 
<< m1 >>
rect 139 130 140 131 
<< m1 >>
rect 140 130 141 131 
<< m1 >>
rect 141 130 142 131 
<< m1 >>
rect 142 130 143 131 
<< m1 >>
rect 143 130 144 131 
<< m1 >>
rect 144 130 145 131 
<< m1 >>
rect 145 130 146 131 
<< m1 >>
rect 147 130 148 131 
<< m1 >>
rect 148 130 149 131 
<< m2 >>
rect 148 130 149 131 
<< m1 >>
rect 149 130 150 131 
<< m1 >>
rect 150 130 151 131 
<< m1 >>
rect 151 130 152 131 
<< m1 >>
rect 152 130 153 131 
<< m1 >>
rect 153 130 154 131 
<< m1 >>
rect 154 130 155 131 
<< m1 >>
rect 155 130 156 131 
<< m1 >>
rect 156 130 157 131 
<< m1 >>
rect 157 130 158 131 
<< m1 >>
rect 158 130 159 131 
<< m1 >>
rect 159 130 160 131 
<< m1 >>
rect 160 130 161 131 
<< m1 >>
rect 161 130 162 131 
<< m2 >>
rect 161 130 162 131 
<< m2c >>
rect 161 130 162 131 
<< m1 >>
rect 161 130 162 131 
<< m2 >>
rect 161 130 162 131 
<< m2 >>
rect 162 130 163 131 
<< m1 >>
rect 163 130 164 131 
<< m2 >>
rect 163 130 164 131 
<< m2 >>
rect 164 130 165 131 
<< m1 >>
rect 165 130 166 131 
<< m2 >>
rect 165 130 166 131 
<< m2 >>
rect 166 130 167 131 
<< m1 >>
rect 167 130 168 131 
<< m2 >>
rect 167 130 168 131 
<< m2c >>
rect 167 130 168 131 
<< m1 >>
rect 167 130 168 131 
<< m2 >>
rect 167 130 168 131 
<< m1 >>
rect 168 130 169 131 
<< m1 >>
rect 169 130 170 131 
<< m2 >>
rect 169 130 170 131 
<< m1 >>
rect 170 130 171 131 
<< m1 >>
rect 171 130 172 131 
<< m1 >>
rect 172 130 173 131 
<< m1 >>
rect 173 130 174 131 
<< m1 >>
rect 174 130 175 131 
<< m1 >>
rect 175 130 176 131 
<< m1 >>
rect 176 130 177 131 
<< m1 >>
rect 177 130 178 131 
<< m2 >>
rect 177 130 178 131 
<< m1 >>
rect 178 130 179 131 
<< m1 >>
rect 179 130 180 131 
<< m1 >>
rect 180 130 181 131 
<< m1 >>
rect 181 130 182 131 
<< m2 >>
rect 182 130 183 131 
<< m2 >>
rect 185 130 186 131 
<< m2 >>
rect 186 130 187 131 
<< m2 >>
rect 187 130 188 131 
<< m2 >>
rect 188 130 189 131 
<< m2 >>
rect 189 130 190 131 
<< m1 >>
rect 190 130 191 131 
<< m2 >>
rect 190 130 191 131 
<< m2 >>
rect 191 130 192 131 
<< m1 >>
rect 192 130 193 131 
<< m2 >>
rect 192 130 193 131 
<< m2c >>
rect 192 130 193 131 
<< m1 >>
rect 192 130 193 131 
<< m2 >>
rect 192 130 193 131 
<< m1 >>
rect 193 130 194 131 
<< m1 >>
rect 194 130 195 131 
<< m1 >>
rect 195 130 196 131 
<< m1 >>
rect 196 130 197 131 
<< m2 >>
rect 196 130 197 131 
<< m1 >>
rect 197 130 198 131 
<< m1 >>
rect 198 130 199 131 
<< m1 >>
rect 214 130 215 131 
<< m1 >>
rect 226 130 227 131 
<< m2 >>
rect 226 130 227 131 
<< m1 >>
rect 229 130 230 131 
<< m1 >>
rect 230 130 231 131 
<< m1 >>
rect 231 130 232 131 
<< m1 >>
rect 232 130 233 131 
<< m1 >>
rect 233 130 234 131 
<< m1 >>
rect 234 130 235 131 
<< m1 >>
rect 235 130 236 131 
<< m1 >>
rect 236 130 237 131 
<< m1 >>
rect 237 130 238 131 
<< m1 >>
rect 238 130 239 131 
<< m1 >>
rect 239 130 240 131 
<< m1 >>
rect 240 130 241 131 
<< m1 >>
rect 241 130 242 131 
<< m1 >>
rect 242 130 243 131 
<< m1 >>
rect 243 130 244 131 
<< m1 >>
rect 244 130 245 131 
<< m1 >>
rect 246 130 247 131 
<< m1 >>
rect 247 130 248 131 
<< m1 >>
rect 248 130 249 131 
<< m1 >>
rect 249 130 250 131 
<< m1 >>
rect 250 130 251 131 
<< m1 >>
rect 253 130 254 131 
<< m2 >>
rect 254 130 255 131 
<< m1 >>
rect 256 130 257 131 
<< m1 >>
rect 19 131 20 132 
<< m1 >>
rect 28 131 29 132 
<< m2 >>
rect 28 131 29 132 
<< m1 >>
rect 34 131 35 132 
<< m1 >>
rect 44 131 45 132 
<< m1 >>
rect 46 131 47 132 
<< m1 >>
rect 57 131 58 132 
<< m1 >>
rect 64 131 65 132 
<< m2 >>
rect 64 131 65 132 
<< m1 >>
rect 73 131 74 132 
<< m1 >>
rect 77 131 78 132 
<< m2 >>
rect 77 131 78 132 
<< m2c >>
rect 77 131 78 132 
<< m1 >>
rect 77 131 78 132 
<< m2 >>
rect 77 131 78 132 
<< m1 >>
rect 79 131 80 132 
<< m2 >>
rect 79 131 80 132 
<< m2c >>
rect 79 131 80 132 
<< m1 >>
rect 79 131 80 132 
<< m2 >>
rect 79 131 80 132 
<< m2 >>
rect 91 131 92 132 
<< m2 >>
rect 100 131 101 132 
<< m1 >>
rect 118 131 119 132 
<< m2 >>
rect 122 131 123 132 
<< m2 >>
rect 129 131 130 132 
<< m2 >>
rect 131 131 132 132 
<< m1 >>
rect 145 131 146 132 
<< m2 >>
rect 148 131 149 132 
<< m2 >>
rect 149 131 150 132 
<< m2 >>
rect 150 131 151 132 
<< m2 >>
rect 151 131 152 132 
<< m2 >>
rect 152 131 153 132 
<< m2 >>
rect 153 131 154 132 
<< m2 >>
rect 154 131 155 132 
<< m2 >>
rect 155 131 156 132 
<< m2 >>
rect 156 131 157 132 
<< m2 >>
rect 157 131 158 132 
<< m2 >>
rect 158 131 159 132 
<< m2 >>
rect 159 131 160 132 
<< m1 >>
rect 163 131 164 132 
<< m1 >>
rect 165 131 166 132 
<< m2 >>
rect 169 131 170 132 
<< m2 >>
rect 177 131 178 132 
<< m1 >>
rect 181 131 182 132 
<< m2 >>
rect 182 131 183 132 
<< m1 >>
rect 190 131 191 132 
<< m2 >>
rect 196 131 197 132 
<< m1 >>
rect 198 131 199 132 
<< m2 >>
rect 198 131 199 132 
<< m2c >>
rect 198 131 199 132 
<< m1 >>
rect 198 131 199 132 
<< m2 >>
rect 198 131 199 132 
<< m1 >>
rect 203 131 204 132 
<< m2 >>
rect 203 131 204 132 
<< m2c >>
rect 203 131 204 132 
<< m1 >>
rect 203 131 204 132 
<< m2 >>
rect 203 131 204 132 
<< m1 >>
rect 204 131 205 132 
<< m1 >>
rect 205 131 206 132 
<< m1 >>
rect 206 131 207 132 
<< m1 >>
rect 207 131 208 132 
<< m1 >>
rect 208 131 209 132 
<< m1 >>
rect 209 131 210 132 
<< m1 >>
rect 210 131 211 132 
<< m1 >>
rect 211 131 212 132 
<< m1 >>
rect 212 131 213 132 
<< m1 >>
rect 213 131 214 132 
<< m1 >>
rect 214 131 215 132 
<< m1 >>
rect 226 131 227 132 
<< m2 >>
rect 226 131 227 132 
<< m1 >>
rect 229 131 230 132 
<< m1 >>
rect 253 131 254 132 
<< m2 >>
rect 254 131 255 132 
<< m1 >>
rect 256 131 257 132 
<< m1 >>
rect 19 132 20 133 
<< m1 >>
rect 28 132 29 133 
<< m2 >>
rect 28 132 29 133 
<< m1 >>
rect 34 132 35 133 
<< m1 >>
rect 44 132 45 133 
<< m1 >>
rect 46 132 47 133 
<< m1 >>
rect 57 132 58 133 
<< m1 >>
rect 64 132 65 133 
<< m2 >>
rect 64 132 65 133 
<< m1 >>
rect 73 132 74 133 
<< m2 >>
rect 77 132 78 133 
<< m2 >>
rect 79 132 80 133 
<< m1 >>
rect 91 132 92 133 
<< m2 >>
rect 91 132 92 133 
<< m2c >>
rect 91 132 92 133 
<< m1 >>
rect 91 132 92 133 
<< m2 >>
rect 91 132 92 133 
<< m1 >>
rect 100 132 101 133 
<< m2 >>
rect 100 132 101 133 
<< m2c >>
rect 100 132 101 133 
<< m1 >>
rect 100 132 101 133 
<< m2 >>
rect 100 132 101 133 
<< m1 >>
rect 118 132 119 133 
<< m1 >>
rect 122 132 123 133 
<< m2 >>
rect 122 132 123 133 
<< m2c >>
rect 122 132 123 133 
<< m1 >>
rect 122 132 123 133 
<< m2 >>
rect 122 132 123 133 
<< m1 >>
rect 129 132 130 133 
<< m2 >>
rect 129 132 130 133 
<< m2c >>
rect 129 132 130 133 
<< m1 >>
rect 129 132 130 133 
<< m2 >>
rect 129 132 130 133 
<< m1 >>
rect 131 132 132 133 
<< m2 >>
rect 131 132 132 133 
<< m2c >>
rect 131 132 132 133 
<< m1 >>
rect 131 132 132 133 
<< m2 >>
rect 131 132 132 133 
<< m1 >>
rect 145 132 146 133 
<< m1 >>
rect 159 132 160 133 
<< m2 >>
rect 159 132 160 133 
<< m2c >>
rect 159 132 160 133 
<< m1 >>
rect 159 132 160 133 
<< m2 >>
rect 159 132 160 133 
<< m1 >>
rect 163 132 164 133 
<< m1 >>
rect 165 132 166 133 
<< m1 >>
rect 169 132 170 133 
<< m2 >>
rect 169 132 170 133 
<< m2c >>
rect 169 132 170 133 
<< m1 >>
rect 169 132 170 133 
<< m2 >>
rect 169 132 170 133 
<< m2 >>
rect 177 132 178 133 
<< m1 >>
rect 178 132 179 133 
<< m1 >>
rect 179 132 180 133 
<< m2 >>
rect 179 132 180 133 
<< m2c >>
rect 179 132 180 133 
<< m1 >>
rect 179 132 180 133 
<< m2 >>
rect 179 132 180 133 
<< m2 >>
rect 180 132 181 133 
<< m1 >>
rect 181 132 182 133 
<< m2 >>
rect 181 132 182 133 
<< m2 >>
rect 182 132 183 133 
<< m1 >>
rect 190 132 191 133 
<< m1 >>
rect 196 132 197 133 
<< m2 >>
rect 196 132 197 133 
<< m2c >>
rect 196 132 197 133 
<< m1 >>
rect 196 132 197 133 
<< m2 >>
rect 196 132 197 133 
<< m2 >>
rect 198 132 199 133 
<< m2 >>
rect 203 132 204 133 
<< m1 >>
rect 226 132 227 133 
<< m2 >>
rect 226 132 227 133 
<< m1 >>
rect 229 132 230 133 
<< m1 >>
rect 253 132 254 133 
<< m2 >>
rect 254 132 255 133 
<< m1 >>
rect 256 132 257 133 
<< m1 >>
rect 19 133 20 134 
<< m1 >>
rect 28 133 29 134 
<< m2 >>
rect 28 133 29 134 
<< m1 >>
rect 34 133 35 134 
<< m1 >>
rect 44 133 45 134 
<< m1 >>
rect 46 133 47 134 
<< m1 >>
rect 57 133 58 134 
<< m1 >>
rect 64 133 65 134 
<< m2 >>
rect 64 133 65 134 
<< m1 >>
rect 73 133 74 134 
<< m2 >>
rect 74 133 75 134 
<< m1 >>
rect 75 133 76 134 
<< m2 >>
rect 75 133 76 134 
<< m2c >>
rect 75 133 76 134 
<< m1 >>
rect 75 133 76 134 
<< m2 >>
rect 75 133 76 134 
<< m1 >>
rect 76 133 77 134 
<< m1 >>
rect 77 133 78 134 
<< m2 >>
rect 77 133 78 134 
<< m1 >>
rect 78 133 79 134 
<< m1 >>
rect 79 133 80 134 
<< m2 >>
rect 79 133 80 134 
<< m1 >>
rect 80 133 81 134 
<< m1 >>
rect 81 133 82 134 
<< m1 >>
rect 82 133 83 134 
<< m1 >>
rect 83 133 84 134 
<< m1 >>
rect 84 133 85 134 
<< m2 >>
rect 84 133 85 134 
<< m1 >>
rect 85 133 86 134 
<< m2 >>
rect 85 133 86 134 
<< m1 >>
rect 86 133 87 134 
<< m2 >>
rect 86 133 87 134 
<< m1 >>
rect 87 133 88 134 
<< m2 >>
rect 87 133 88 134 
<< m1 >>
rect 88 133 89 134 
<< m1 >>
rect 89 133 90 134 
<< m1 >>
rect 91 133 92 134 
<< m1 >>
rect 100 133 101 134 
<< m1 >>
rect 118 133 119 134 
<< m1 >>
rect 120 133 121 134 
<< m1 >>
rect 121 133 122 134 
<< m1 >>
rect 122 133 123 134 
<< m1 >>
rect 129 133 130 134 
<< m1 >>
rect 131 133 132 134 
<< m1 >>
rect 145 133 146 134 
<< m1 >>
rect 159 133 160 134 
<< m1 >>
rect 163 133 164 134 
<< m1 >>
rect 165 133 166 134 
<< m1 >>
rect 169 133 170 134 
<< m2 >>
rect 177 133 178 134 
<< m1 >>
rect 178 133 179 134 
<< m1 >>
rect 181 133 182 134 
<< m1 >>
rect 190 133 191 134 
<< m1 >>
rect 196 133 197 134 
<< m2 >>
rect 198 133 199 134 
<< m1 >>
rect 199 133 200 134 
<< m1 >>
rect 200 133 201 134 
<< m1 >>
rect 201 133 202 134 
<< m1 >>
rect 202 133 203 134 
<< m1 >>
rect 203 133 204 134 
<< m2 >>
rect 203 133 204 134 
<< m1 >>
rect 204 133 205 134 
<< m1 >>
rect 205 133 206 134 
<< m1 >>
rect 206 133 207 134 
<< m1 >>
rect 207 133 208 134 
<< m1 >>
rect 208 133 209 134 
<< m1 >>
rect 209 133 210 134 
<< m1 >>
rect 210 133 211 134 
<< m1 >>
rect 211 133 212 134 
<< m1 >>
rect 212 133 213 134 
<< m1 >>
rect 213 133 214 134 
<< m1 >>
rect 214 133 215 134 
<< m1 >>
rect 226 133 227 134 
<< m2 >>
rect 226 133 227 134 
<< m1 >>
rect 229 133 230 134 
<< m1 >>
rect 253 133 254 134 
<< m2 >>
rect 254 133 255 134 
<< m1 >>
rect 256 133 257 134 
<< m1 >>
rect 19 134 20 135 
<< m1 >>
rect 28 134 29 135 
<< m2 >>
rect 28 134 29 135 
<< m1 >>
rect 34 134 35 135 
<< m1 >>
rect 44 134 45 135 
<< m1 >>
rect 46 134 47 135 
<< m1 >>
rect 57 134 58 135 
<< m2 >>
rect 57 134 58 135 
<< m2c >>
rect 57 134 58 135 
<< m1 >>
rect 57 134 58 135 
<< m2 >>
rect 57 134 58 135 
<< m1 >>
rect 64 134 65 135 
<< m2 >>
rect 64 134 65 135 
<< m1 >>
rect 73 134 74 135 
<< m2 >>
rect 74 134 75 135 
<< m2 >>
rect 77 134 78 135 
<< m2 >>
rect 79 134 80 135 
<< m2 >>
rect 84 134 85 135 
<< m2 >>
rect 87 134 88 135 
<< m1 >>
rect 89 134 90 135 
<< m2 >>
rect 89 134 90 135 
<< m2c >>
rect 89 134 90 135 
<< m1 >>
rect 89 134 90 135 
<< m2 >>
rect 89 134 90 135 
<< m2 >>
rect 90 134 91 135 
<< m1 >>
rect 91 134 92 135 
<< m2 >>
rect 91 134 92 135 
<< m2 >>
rect 92 134 93 135 
<< m1 >>
rect 93 134 94 135 
<< m2 >>
rect 93 134 94 135 
<< m2c >>
rect 93 134 94 135 
<< m1 >>
rect 93 134 94 135 
<< m2 >>
rect 93 134 94 135 
<< m1 >>
rect 94 134 95 135 
<< m1 >>
rect 95 134 96 135 
<< m1 >>
rect 96 134 97 135 
<< m1 >>
rect 97 134 98 135 
<< m1 >>
rect 98 134 99 135 
<< m1 >>
rect 99 134 100 135 
<< m1 >>
rect 100 134 101 135 
<< m1 >>
rect 118 134 119 135 
<< m1 >>
rect 120 134 121 135 
<< m1 >>
rect 129 134 130 135 
<< m1 >>
rect 131 134 132 135 
<< m1 >>
rect 145 134 146 135 
<< m1 >>
rect 159 134 160 135 
<< m1 >>
rect 163 134 164 135 
<< m1 >>
rect 165 134 166 135 
<< m1 >>
rect 169 134 170 135 
<< m2 >>
rect 177 134 178 135 
<< m1 >>
rect 178 134 179 135 
<< m1 >>
rect 181 134 182 135 
<< m1 >>
rect 190 134 191 135 
<< m1 >>
rect 196 134 197 135 
<< m2 >>
rect 198 134 199 135 
<< m1 >>
rect 199 134 200 135 
<< m2 >>
rect 203 134 204 135 
<< m1 >>
rect 214 134 215 135 
<< m1 >>
rect 226 134 227 135 
<< m2 >>
rect 226 134 227 135 
<< m1 >>
rect 229 134 230 135 
<< m1 >>
rect 253 134 254 135 
<< m2 >>
rect 254 134 255 135 
<< m1 >>
rect 256 134 257 135 
<< m1 >>
rect 19 135 20 136 
<< m1 >>
rect 28 135 29 136 
<< m2 >>
rect 28 135 29 136 
<< m1 >>
rect 34 135 35 136 
<< m1 >>
rect 44 135 45 136 
<< m1 >>
rect 46 135 47 136 
<< m2 >>
rect 51 135 52 136 
<< m2 >>
rect 52 135 53 136 
<< m2 >>
rect 53 135 54 136 
<< m2 >>
rect 54 135 55 136 
<< m2 >>
rect 55 135 56 136 
<< m2 >>
rect 57 135 58 136 
<< m1 >>
rect 64 135 65 136 
<< m2 >>
rect 64 135 65 136 
<< m1 >>
rect 73 135 74 136 
<< m2 >>
rect 74 135 75 136 
<< m1 >>
rect 77 135 78 136 
<< m2 >>
rect 77 135 78 136 
<< m2c >>
rect 77 135 78 136 
<< m1 >>
rect 77 135 78 136 
<< m2 >>
rect 77 135 78 136 
<< m1 >>
rect 79 135 80 136 
<< m2 >>
rect 79 135 80 136 
<< m2c >>
rect 79 135 80 136 
<< m1 >>
rect 79 135 80 136 
<< m2 >>
rect 79 135 80 136 
<< m1 >>
rect 82 135 83 136 
<< m1 >>
rect 83 135 84 136 
<< m1 >>
rect 84 135 85 136 
<< m2 >>
rect 84 135 85 136 
<< m2c >>
rect 84 135 85 136 
<< m1 >>
rect 84 135 85 136 
<< m2 >>
rect 84 135 85 136 
<< m1 >>
rect 87 135 88 136 
<< m2 >>
rect 87 135 88 136 
<< m2c >>
rect 87 135 88 136 
<< m1 >>
rect 87 135 88 136 
<< m2 >>
rect 87 135 88 136 
<< m1 >>
rect 91 135 92 136 
<< m1 >>
rect 118 135 119 136 
<< m1 >>
rect 120 135 121 136 
<< m1 >>
rect 129 135 130 136 
<< m1 >>
rect 131 135 132 136 
<< m1 >>
rect 145 135 146 136 
<< m1 >>
rect 159 135 160 136 
<< m1 >>
rect 160 135 161 136 
<< m1 >>
rect 161 135 162 136 
<< m1 >>
rect 163 135 164 136 
<< m1 >>
rect 165 135 166 136 
<< m1 >>
rect 169 135 170 136 
<< m2 >>
rect 177 135 178 136 
<< m1 >>
rect 178 135 179 136 
<< m2 >>
rect 178 135 179 136 
<< m2 >>
rect 179 135 180 136 
<< m2 >>
rect 180 135 181 136 
<< m1 >>
rect 181 135 182 136 
<< m2 >>
rect 181 135 182 136 
<< m2 >>
rect 182 135 183 136 
<< m1 >>
rect 190 135 191 136 
<< m1 >>
rect 196 135 197 136 
<< m2 >>
rect 198 135 199 136 
<< m1 >>
rect 199 135 200 136 
<< m2 >>
rect 199 135 200 136 
<< m2 >>
rect 200 135 201 136 
<< m1 >>
rect 201 135 202 136 
<< m2 >>
rect 201 135 202 136 
<< m2c >>
rect 201 135 202 136 
<< m1 >>
rect 201 135 202 136 
<< m2 >>
rect 201 135 202 136 
<< m1 >>
rect 203 135 204 136 
<< m2 >>
rect 203 135 204 136 
<< m2c >>
rect 203 135 204 136 
<< m1 >>
rect 203 135 204 136 
<< m2 >>
rect 203 135 204 136 
<< m1 >>
rect 214 135 215 136 
<< m1 >>
rect 226 135 227 136 
<< m2 >>
rect 226 135 227 136 
<< m1 >>
rect 229 135 230 136 
<< m1 >>
rect 253 135 254 136 
<< m2 >>
rect 254 135 255 136 
<< m1 >>
rect 256 135 257 136 
<< m1 >>
rect 19 136 20 137 
<< m1 >>
rect 28 136 29 137 
<< m2 >>
rect 28 136 29 137 
<< m1 >>
rect 34 136 35 137 
<< m1 >>
rect 44 136 45 137 
<< m1 >>
rect 46 136 47 137 
<< m1 >>
rect 49 136 50 137 
<< m1 >>
rect 50 136 51 137 
<< m2 >>
rect 50 136 51 137 
<< m2c >>
rect 50 136 51 137 
<< m1 >>
rect 50 136 51 137 
<< m2 >>
rect 50 136 51 137 
<< m2 >>
rect 51 136 52 137 
<< m1 >>
rect 52 136 53 137 
<< m1 >>
rect 53 136 54 137 
<< m1 >>
rect 54 136 55 137 
<< m1 >>
rect 55 136 56 137 
<< m2 >>
rect 55 136 56 137 
<< m1 >>
rect 56 136 57 137 
<< m1 >>
rect 57 136 58 137 
<< m2 >>
rect 57 136 58 137 
<< m1 >>
rect 58 136 59 137 
<< m1 >>
rect 59 136 60 137 
<< m1 >>
rect 60 136 61 137 
<< m1 >>
rect 61 136 62 137 
<< m1 >>
rect 62 136 63 137 
<< m1 >>
rect 64 136 65 137 
<< m2 >>
rect 64 136 65 137 
<< m1 >>
rect 65 136 66 137 
<< m1 >>
rect 66 136 67 137 
<< m1 >>
rect 67 136 68 137 
<< m1 >>
rect 73 136 74 137 
<< m2 >>
rect 74 136 75 137 
<< m1 >>
rect 77 136 78 137 
<< m1 >>
rect 79 136 80 137 
<< m1 >>
rect 82 136 83 137 
<< m1 >>
rect 87 136 88 137 
<< m1 >>
rect 88 136 89 137 
<< m1 >>
rect 91 136 92 137 
<< m2 >>
rect 117 136 118 137 
<< m1 >>
rect 118 136 119 137 
<< m2 >>
rect 118 136 119 137 
<< m2 >>
rect 119 136 120 137 
<< m1 >>
rect 120 136 121 137 
<< m2 >>
rect 120 136 121 137 
<< m2c >>
rect 120 136 121 137 
<< m1 >>
rect 120 136 121 137 
<< m2 >>
rect 120 136 121 137 
<< m1 >>
rect 129 136 130 137 
<< m1 >>
rect 131 136 132 137 
<< m1 >>
rect 145 136 146 137 
<< m1 >>
rect 161 136 162 137 
<< m2 >>
rect 161 136 162 137 
<< m2c >>
rect 161 136 162 137 
<< m1 >>
rect 161 136 162 137 
<< m2 >>
rect 161 136 162 137 
<< m2 >>
rect 162 136 163 137 
<< m1 >>
rect 163 136 164 137 
<< m2 >>
rect 163 136 164 137 
<< m2 >>
rect 164 136 165 137 
<< m1 >>
rect 165 136 166 137 
<< m2 >>
rect 165 136 166 137 
<< m2 >>
rect 166 136 167 137 
<< m1 >>
rect 169 136 170 137 
<< m1 >>
rect 178 136 179 137 
<< m1 >>
rect 181 136 182 137 
<< m2 >>
rect 182 136 183 137 
<< m1 >>
rect 190 136 191 137 
<< m1 >>
rect 196 136 197 137 
<< m1 >>
rect 199 136 200 137 
<< m1 >>
rect 201 136 202 137 
<< m1 >>
rect 203 136 204 137 
<< m1 >>
rect 214 136 215 137 
<< m1 >>
rect 226 136 227 137 
<< m2 >>
rect 226 136 227 137 
<< m1 >>
rect 229 136 230 137 
<< m1 >>
rect 253 136 254 137 
<< m2 >>
rect 254 136 255 137 
<< m1 >>
rect 256 136 257 137 
<< m1 >>
rect 19 137 20 138 
<< m1 >>
rect 28 137 29 138 
<< m2 >>
rect 28 137 29 138 
<< m1 >>
rect 34 137 35 138 
<< m1 >>
rect 44 137 45 138 
<< m1 >>
rect 46 137 47 138 
<< m1 >>
rect 49 137 50 138 
<< m1 >>
rect 52 137 53 138 
<< m2 >>
rect 55 137 56 138 
<< m2 >>
rect 57 137 58 138 
<< m1 >>
rect 62 137 63 138 
<< m2 >>
rect 64 137 65 138 
<< m1 >>
rect 67 137 68 138 
<< m1 >>
rect 73 137 74 138 
<< m2 >>
rect 74 137 75 138 
<< m1 >>
rect 75 137 76 138 
<< m2 >>
rect 75 137 76 138 
<< m2c >>
rect 75 137 76 138 
<< m1 >>
rect 75 137 76 138 
<< m2 >>
rect 75 137 76 138 
<< m2 >>
rect 76 137 77 138 
<< m1 >>
rect 77 137 78 138 
<< m2 >>
rect 77 137 78 138 
<< m2 >>
rect 78 137 79 138 
<< m1 >>
rect 79 137 80 138 
<< m2 >>
rect 79 137 80 138 
<< m2c >>
rect 79 137 80 138 
<< m1 >>
rect 79 137 80 138 
<< m2 >>
rect 79 137 80 138 
<< m1 >>
rect 82 137 83 138 
<< m1 >>
rect 88 137 89 138 
<< m1 >>
rect 91 137 92 138 
<< m2 >>
rect 117 137 118 138 
<< m1 >>
rect 118 137 119 138 
<< m1 >>
rect 129 137 130 138 
<< m1 >>
rect 131 137 132 138 
<< m1 >>
rect 145 137 146 138 
<< m1 >>
rect 163 137 164 138 
<< m1 >>
rect 165 137 166 138 
<< m2 >>
rect 166 137 167 138 
<< m1 >>
rect 169 137 170 138 
<< m1 >>
rect 178 137 179 138 
<< m1 >>
rect 181 137 182 138 
<< m2 >>
rect 182 137 183 138 
<< m1 >>
rect 190 137 191 138 
<< m1 >>
rect 196 137 197 138 
<< m1 >>
rect 199 137 200 138 
<< m1 >>
rect 201 137 202 138 
<< m1 >>
rect 203 137 204 138 
<< m1 >>
rect 214 137 215 138 
<< m1 >>
rect 226 137 227 138 
<< m2 >>
rect 226 137 227 138 
<< m1 >>
rect 229 137 230 138 
<< m1 >>
rect 253 137 254 138 
<< m2 >>
rect 254 137 255 138 
<< m1 >>
rect 256 137 257 138 
<< m1 >>
rect 19 138 20 139 
<< m1 >>
rect 28 138 29 139 
<< m2 >>
rect 28 138 29 139 
<< pdiffusion >>
rect 30 138 31 139 
<< pdiffusion >>
rect 31 138 32 139 
<< pdiffusion >>
rect 32 138 33 139 
<< pdiffusion >>
rect 33 138 34 139 
<< m1 >>
rect 34 138 35 139 
<< pdiffusion >>
rect 34 138 35 139 
<< pdiffusion >>
rect 35 138 36 139 
<< m1 >>
rect 44 138 45 139 
<< m1 >>
rect 46 138 47 139 
<< pdiffusion >>
rect 48 138 49 139 
<< m1 >>
rect 49 138 50 139 
<< pdiffusion >>
rect 49 138 50 139 
<< pdiffusion >>
rect 50 138 51 139 
<< pdiffusion >>
rect 51 138 52 139 
<< m1 >>
rect 52 138 53 139 
<< pdiffusion >>
rect 52 138 53 139 
<< pdiffusion >>
rect 53 138 54 139 
<< m1 >>
rect 55 138 56 139 
<< m2 >>
rect 55 138 56 139 
<< m2c >>
rect 55 138 56 139 
<< m1 >>
rect 55 138 56 139 
<< m2 >>
rect 55 138 56 139 
<< m1 >>
rect 57 138 58 139 
<< m2 >>
rect 57 138 58 139 
<< m2c >>
rect 57 138 58 139 
<< m1 >>
rect 57 138 58 139 
<< m2 >>
rect 57 138 58 139 
<< m1 >>
rect 62 138 63 139 
<< m1 >>
rect 64 138 65 139 
<< m2 >>
rect 64 138 65 139 
<< m2c >>
rect 64 138 65 139 
<< m1 >>
rect 64 138 65 139 
<< m2 >>
rect 64 138 65 139 
<< pdiffusion >>
rect 66 138 67 139 
<< m1 >>
rect 67 138 68 139 
<< pdiffusion >>
rect 67 138 68 139 
<< pdiffusion >>
rect 68 138 69 139 
<< pdiffusion >>
rect 69 138 70 139 
<< pdiffusion >>
rect 70 138 71 139 
<< pdiffusion >>
rect 71 138 72 139 
<< m1 >>
rect 73 138 74 139 
<< m2 >>
rect 74 138 75 139 
<< m1 >>
rect 75 138 76 139 
<< m1 >>
rect 77 138 78 139 
<< m1 >>
rect 82 138 83 139 
<< pdiffusion >>
rect 84 138 85 139 
<< pdiffusion >>
rect 85 138 86 139 
<< pdiffusion >>
rect 86 138 87 139 
<< pdiffusion >>
rect 87 138 88 139 
<< m1 >>
rect 88 138 89 139 
<< pdiffusion >>
rect 88 138 89 139 
<< pdiffusion >>
rect 89 138 90 139 
<< m1 >>
rect 91 138 92 139 
<< m2 >>
rect 117 138 118 139 
<< m1 >>
rect 118 138 119 139 
<< pdiffusion >>
rect 120 138 121 139 
<< pdiffusion >>
rect 121 138 122 139 
<< pdiffusion >>
rect 122 138 123 139 
<< pdiffusion >>
rect 123 138 124 139 
<< pdiffusion >>
rect 124 138 125 139 
<< pdiffusion >>
rect 125 138 126 139 
<< m1 >>
rect 129 138 130 139 
<< m1 >>
rect 131 138 132 139 
<< pdiffusion >>
rect 138 138 139 139 
<< pdiffusion >>
rect 139 138 140 139 
<< pdiffusion >>
rect 140 138 141 139 
<< pdiffusion >>
rect 141 138 142 139 
<< pdiffusion >>
rect 142 138 143 139 
<< pdiffusion >>
rect 143 138 144 139 
<< m1 >>
rect 145 138 146 139 
<< pdiffusion >>
rect 156 138 157 139 
<< pdiffusion >>
rect 157 138 158 139 
<< pdiffusion >>
rect 158 138 159 139 
<< pdiffusion >>
rect 159 138 160 139 
<< pdiffusion >>
rect 160 138 161 139 
<< pdiffusion >>
rect 161 138 162 139 
<< m1 >>
rect 163 138 164 139 
<< m1 >>
rect 165 138 166 139 
<< m2 >>
rect 166 138 167 139 
<< m1 >>
rect 169 138 170 139 
<< pdiffusion >>
rect 174 138 175 139 
<< pdiffusion >>
rect 175 138 176 139 
<< pdiffusion >>
rect 176 138 177 139 
<< pdiffusion >>
rect 177 138 178 139 
<< m1 >>
rect 178 138 179 139 
<< pdiffusion >>
rect 178 138 179 139 
<< pdiffusion >>
rect 179 138 180 139 
<< m1 >>
rect 181 138 182 139 
<< m2 >>
rect 182 138 183 139 
<< m1 >>
rect 190 138 191 139 
<< pdiffusion >>
rect 192 138 193 139 
<< pdiffusion >>
rect 193 138 194 139 
<< pdiffusion >>
rect 194 138 195 139 
<< pdiffusion >>
rect 195 138 196 139 
<< m1 >>
rect 196 138 197 139 
<< pdiffusion >>
rect 196 138 197 139 
<< pdiffusion >>
rect 197 138 198 139 
<< m1 >>
rect 199 138 200 139 
<< m1 >>
rect 201 138 202 139 
<< m1 >>
rect 203 138 204 139 
<< pdiffusion >>
rect 210 138 211 139 
<< pdiffusion >>
rect 211 138 212 139 
<< pdiffusion >>
rect 212 138 213 139 
<< pdiffusion >>
rect 213 138 214 139 
<< m1 >>
rect 214 138 215 139 
<< pdiffusion >>
rect 214 138 215 139 
<< pdiffusion >>
rect 215 138 216 139 
<< m1 >>
rect 226 138 227 139 
<< m2 >>
rect 226 138 227 139 
<< pdiffusion >>
rect 228 138 229 139 
<< m1 >>
rect 229 138 230 139 
<< pdiffusion >>
rect 229 138 230 139 
<< pdiffusion >>
rect 230 138 231 139 
<< pdiffusion >>
rect 231 138 232 139 
<< pdiffusion >>
rect 232 138 233 139 
<< pdiffusion >>
rect 233 138 234 139 
<< pdiffusion >>
rect 246 138 247 139 
<< pdiffusion >>
rect 247 138 248 139 
<< pdiffusion >>
rect 248 138 249 139 
<< pdiffusion >>
rect 249 138 250 139 
<< pdiffusion >>
rect 250 138 251 139 
<< pdiffusion >>
rect 251 138 252 139 
<< m1 >>
rect 253 138 254 139 
<< m2 >>
rect 254 138 255 139 
<< m1 >>
rect 256 138 257 139 
<< m1 >>
rect 19 139 20 140 
<< m1 >>
rect 28 139 29 140 
<< m2 >>
rect 28 139 29 140 
<< pdiffusion >>
rect 30 139 31 140 
<< pdiffusion >>
rect 31 139 32 140 
<< pdiffusion >>
rect 32 139 33 140 
<< pdiffusion >>
rect 33 139 34 140 
<< pdiffusion >>
rect 34 139 35 140 
<< pdiffusion >>
rect 35 139 36 140 
<< m1 >>
rect 44 139 45 140 
<< m1 >>
rect 46 139 47 140 
<< pdiffusion >>
rect 48 139 49 140 
<< pdiffusion >>
rect 49 139 50 140 
<< pdiffusion >>
rect 50 139 51 140 
<< pdiffusion >>
rect 51 139 52 140 
<< pdiffusion >>
rect 52 139 53 140 
<< pdiffusion >>
rect 53 139 54 140 
<< m1 >>
rect 55 139 56 140 
<< m1 >>
rect 57 139 58 140 
<< m1 >>
rect 62 139 63 140 
<< m1 >>
rect 64 139 65 140 
<< pdiffusion >>
rect 66 139 67 140 
<< pdiffusion >>
rect 67 139 68 140 
<< pdiffusion >>
rect 68 139 69 140 
<< pdiffusion >>
rect 69 139 70 140 
<< pdiffusion >>
rect 70 139 71 140 
<< pdiffusion >>
rect 71 139 72 140 
<< m1 >>
rect 73 139 74 140 
<< m2 >>
rect 74 139 75 140 
<< m1 >>
rect 75 139 76 140 
<< m1 >>
rect 77 139 78 140 
<< m1 >>
rect 82 139 83 140 
<< pdiffusion >>
rect 84 139 85 140 
<< pdiffusion >>
rect 85 139 86 140 
<< pdiffusion >>
rect 86 139 87 140 
<< pdiffusion >>
rect 87 139 88 140 
<< pdiffusion >>
rect 88 139 89 140 
<< pdiffusion >>
rect 89 139 90 140 
<< m1 >>
rect 91 139 92 140 
<< m2 >>
rect 117 139 118 140 
<< m1 >>
rect 118 139 119 140 
<< pdiffusion >>
rect 120 139 121 140 
<< pdiffusion >>
rect 121 139 122 140 
<< pdiffusion >>
rect 122 139 123 140 
<< pdiffusion >>
rect 123 139 124 140 
<< pdiffusion >>
rect 124 139 125 140 
<< pdiffusion >>
rect 125 139 126 140 
<< m1 >>
rect 129 139 130 140 
<< m1 >>
rect 131 139 132 140 
<< pdiffusion >>
rect 138 139 139 140 
<< pdiffusion >>
rect 139 139 140 140 
<< pdiffusion >>
rect 140 139 141 140 
<< pdiffusion >>
rect 141 139 142 140 
<< pdiffusion >>
rect 142 139 143 140 
<< pdiffusion >>
rect 143 139 144 140 
<< m1 >>
rect 145 139 146 140 
<< pdiffusion >>
rect 156 139 157 140 
<< pdiffusion >>
rect 157 139 158 140 
<< pdiffusion >>
rect 158 139 159 140 
<< pdiffusion >>
rect 159 139 160 140 
<< pdiffusion >>
rect 160 139 161 140 
<< pdiffusion >>
rect 161 139 162 140 
<< m1 >>
rect 163 139 164 140 
<< m1 >>
rect 165 139 166 140 
<< m2 >>
rect 166 139 167 140 
<< m1 >>
rect 169 139 170 140 
<< pdiffusion >>
rect 174 139 175 140 
<< pdiffusion >>
rect 175 139 176 140 
<< pdiffusion >>
rect 176 139 177 140 
<< pdiffusion >>
rect 177 139 178 140 
<< pdiffusion >>
rect 178 139 179 140 
<< pdiffusion >>
rect 179 139 180 140 
<< m1 >>
rect 181 139 182 140 
<< m2 >>
rect 182 139 183 140 
<< m1 >>
rect 190 139 191 140 
<< pdiffusion >>
rect 192 139 193 140 
<< pdiffusion >>
rect 193 139 194 140 
<< pdiffusion >>
rect 194 139 195 140 
<< pdiffusion >>
rect 195 139 196 140 
<< pdiffusion >>
rect 196 139 197 140 
<< pdiffusion >>
rect 197 139 198 140 
<< m1 >>
rect 199 139 200 140 
<< m1 >>
rect 201 139 202 140 
<< m1 >>
rect 203 139 204 140 
<< pdiffusion >>
rect 210 139 211 140 
<< pdiffusion >>
rect 211 139 212 140 
<< pdiffusion >>
rect 212 139 213 140 
<< pdiffusion >>
rect 213 139 214 140 
<< pdiffusion >>
rect 214 139 215 140 
<< pdiffusion >>
rect 215 139 216 140 
<< m1 >>
rect 226 139 227 140 
<< m2 >>
rect 226 139 227 140 
<< pdiffusion >>
rect 228 139 229 140 
<< pdiffusion >>
rect 229 139 230 140 
<< pdiffusion >>
rect 230 139 231 140 
<< pdiffusion >>
rect 231 139 232 140 
<< pdiffusion >>
rect 232 139 233 140 
<< pdiffusion >>
rect 233 139 234 140 
<< pdiffusion >>
rect 246 139 247 140 
<< pdiffusion >>
rect 247 139 248 140 
<< pdiffusion >>
rect 248 139 249 140 
<< pdiffusion >>
rect 249 139 250 140 
<< pdiffusion >>
rect 250 139 251 140 
<< pdiffusion >>
rect 251 139 252 140 
<< m1 >>
rect 253 139 254 140 
<< m2 >>
rect 254 139 255 140 
<< m1 >>
rect 256 139 257 140 
<< m1 >>
rect 19 140 20 141 
<< m1 >>
rect 28 140 29 141 
<< m2 >>
rect 28 140 29 141 
<< pdiffusion >>
rect 30 140 31 141 
<< pdiffusion >>
rect 31 140 32 141 
<< pdiffusion >>
rect 32 140 33 141 
<< pdiffusion >>
rect 33 140 34 141 
<< pdiffusion >>
rect 34 140 35 141 
<< pdiffusion >>
rect 35 140 36 141 
<< m1 >>
rect 44 140 45 141 
<< m1 >>
rect 46 140 47 141 
<< pdiffusion >>
rect 48 140 49 141 
<< pdiffusion >>
rect 49 140 50 141 
<< pdiffusion >>
rect 50 140 51 141 
<< pdiffusion >>
rect 51 140 52 141 
<< pdiffusion >>
rect 52 140 53 141 
<< pdiffusion >>
rect 53 140 54 141 
<< m1 >>
rect 55 140 56 141 
<< m1 >>
rect 57 140 58 141 
<< m1 >>
rect 62 140 63 141 
<< m1 >>
rect 64 140 65 141 
<< pdiffusion >>
rect 66 140 67 141 
<< pdiffusion >>
rect 67 140 68 141 
<< pdiffusion >>
rect 68 140 69 141 
<< pdiffusion >>
rect 69 140 70 141 
<< pdiffusion >>
rect 70 140 71 141 
<< pdiffusion >>
rect 71 140 72 141 
<< m1 >>
rect 73 140 74 141 
<< m2 >>
rect 74 140 75 141 
<< m1 >>
rect 75 140 76 141 
<< m1 >>
rect 77 140 78 141 
<< m1 >>
rect 82 140 83 141 
<< pdiffusion >>
rect 84 140 85 141 
<< pdiffusion >>
rect 85 140 86 141 
<< pdiffusion >>
rect 86 140 87 141 
<< pdiffusion >>
rect 87 140 88 141 
<< pdiffusion >>
rect 88 140 89 141 
<< pdiffusion >>
rect 89 140 90 141 
<< m1 >>
rect 91 140 92 141 
<< m2 >>
rect 117 140 118 141 
<< m1 >>
rect 118 140 119 141 
<< pdiffusion >>
rect 120 140 121 141 
<< pdiffusion >>
rect 121 140 122 141 
<< pdiffusion >>
rect 122 140 123 141 
<< pdiffusion >>
rect 123 140 124 141 
<< pdiffusion >>
rect 124 140 125 141 
<< pdiffusion >>
rect 125 140 126 141 
<< m1 >>
rect 129 140 130 141 
<< m1 >>
rect 131 140 132 141 
<< pdiffusion >>
rect 138 140 139 141 
<< pdiffusion >>
rect 139 140 140 141 
<< pdiffusion >>
rect 140 140 141 141 
<< pdiffusion >>
rect 141 140 142 141 
<< pdiffusion >>
rect 142 140 143 141 
<< pdiffusion >>
rect 143 140 144 141 
<< m1 >>
rect 145 140 146 141 
<< pdiffusion >>
rect 156 140 157 141 
<< pdiffusion >>
rect 157 140 158 141 
<< pdiffusion >>
rect 158 140 159 141 
<< pdiffusion >>
rect 159 140 160 141 
<< pdiffusion >>
rect 160 140 161 141 
<< pdiffusion >>
rect 161 140 162 141 
<< m1 >>
rect 163 140 164 141 
<< m1 >>
rect 165 140 166 141 
<< m2 >>
rect 166 140 167 141 
<< m1 >>
rect 169 140 170 141 
<< pdiffusion >>
rect 174 140 175 141 
<< pdiffusion >>
rect 175 140 176 141 
<< pdiffusion >>
rect 176 140 177 141 
<< pdiffusion >>
rect 177 140 178 141 
<< pdiffusion >>
rect 178 140 179 141 
<< pdiffusion >>
rect 179 140 180 141 
<< m1 >>
rect 181 140 182 141 
<< m2 >>
rect 182 140 183 141 
<< m1 >>
rect 190 140 191 141 
<< pdiffusion >>
rect 192 140 193 141 
<< pdiffusion >>
rect 193 140 194 141 
<< pdiffusion >>
rect 194 140 195 141 
<< pdiffusion >>
rect 195 140 196 141 
<< pdiffusion >>
rect 196 140 197 141 
<< pdiffusion >>
rect 197 140 198 141 
<< m1 >>
rect 199 140 200 141 
<< m1 >>
rect 201 140 202 141 
<< m1 >>
rect 203 140 204 141 
<< pdiffusion >>
rect 210 140 211 141 
<< pdiffusion >>
rect 211 140 212 141 
<< pdiffusion >>
rect 212 140 213 141 
<< pdiffusion >>
rect 213 140 214 141 
<< pdiffusion >>
rect 214 140 215 141 
<< pdiffusion >>
rect 215 140 216 141 
<< m1 >>
rect 226 140 227 141 
<< m2 >>
rect 226 140 227 141 
<< pdiffusion >>
rect 228 140 229 141 
<< pdiffusion >>
rect 229 140 230 141 
<< pdiffusion >>
rect 230 140 231 141 
<< pdiffusion >>
rect 231 140 232 141 
<< pdiffusion >>
rect 232 140 233 141 
<< pdiffusion >>
rect 233 140 234 141 
<< pdiffusion >>
rect 246 140 247 141 
<< pdiffusion >>
rect 247 140 248 141 
<< pdiffusion >>
rect 248 140 249 141 
<< pdiffusion >>
rect 249 140 250 141 
<< pdiffusion >>
rect 250 140 251 141 
<< pdiffusion >>
rect 251 140 252 141 
<< m1 >>
rect 253 140 254 141 
<< m2 >>
rect 254 140 255 141 
<< m1 >>
rect 256 140 257 141 
<< m1 >>
rect 19 141 20 142 
<< m1 >>
rect 28 141 29 142 
<< m2 >>
rect 28 141 29 142 
<< pdiffusion >>
rect 30 141 31 142 
<< pdiffusion >>
rect 31 141 32 142 
<< pdiffusion >>
rect 32 141 33 142 
<< pdiffusion >>
rect 33 141 34 142 
<< pdiffusion >>
rect 34 141 35 142 
<< pdiffusion >>
rect 35 141 36 142 
<< m1 >>
rect 44 141 45 142 
<< m1 >>
rect 46 141 47 142 
<< pdiffusion >>
rect 48 141 49 142 
<< pdiffusion >>
rect 49 141 50 142 
<< pdiffusion >>
rect 50 141 51 142 
<< pdiffusion >>
rect 51 141 52 142 
<< pdiffusion >>
rect 52 141 53 142 
<< pdiffusion >>
rect 53 141 54 142 
<< m1 >>
rect 55 141 56 142 
<< m1 >>
rect 57 141 58 142 
<< m1 >>
rect 62 141 63 142 
<< m1 >>
rect 64 141 65 142 
<< pdiffusion >>
rect 66 141 67 142 
<< pdiffusion >>
rect 67 141 68 142 
<< pdiffusion >>
rect 68 141 69 142 
<< pdiffusion >>
rect 69 141 70 142 
<< pdiffusion >>
rect 70 141 71 142 
<< pdiffusion >>
rect 71 141 72 142 
<< m1 >>
rect 73 141 74 142 
<< m2 >>
rect 74 141 75 142 
<< m1 >>
rect 75 141 76 142 
<< m1 >>
rect 77 141 78 142 
<< m1 >>
rect 82 141 83 142 
<< pdiffusion >>
rect 84 141 85 142 
<< pdiffusion >>
rect 85 141 86 142 
<< pdiffusion >>
rect 86 141 87 142 
<< pdiffusion >>
rect 87 141 88 142 
<< pdiffusion >>
rect 88 141 89 142 
<< pdiffusion >>
rect 89 141 90 142 
<< m1 >>
rect 91 141 92 142 
<< m2 >>
rect 117 141 118 142 
<< m1 >>
rect 118 141 119 142 
<< pdiffusion >>
rect 120 141 121 142 
<< pdiffusion >>
rect 121 141 122 142 
<< pdiffusion >>
rect 122 141 123 142 
<< pdiffusion >>
rect 123 141 124 142 
<< pdiffusion >>
rect 124 141 125 142 
<< pdiffusion >>
rect 125 141 126 142 
<< m1 >>
rect 129 141 130 142 
<< m1 >>
rect 131 141 132 142 
<< pdiffusion >>
rect 138 141 139 142 
<< pdiffusion >>
rect 139 141 140 142 
<< pdiffusion >>
rect 140 141 141 142 
<< pdiffusion >>
rect 141 141 142 142 
<< pdiffusion >>
rect 142 141 143 142 
<< pdiffusion >>
rect 143 141 144 142 
<< m1 >>
rect 145 141 146 142 
<< pdiffusion >>
rect 156 141 157 142 
<< pdiffusion >>
rect 157 141 158 142 
<< pdiffusion >>
rect 158 141 159 142 
<< pdiffusion >>
rect 159 141 160 142 
<< pdiffusion >>
rect 160 141 161 142 
<< pdiffusion >>
rect 161 141 162 142 
<< m1 >>
rect 163 141 164 142 
<< m1 >>
rect 165 141 166 142 
<< m2 >>
rect 166 141 167 142 
<< m1 >>
rect 169 141 170 142 
<< pdiffusion >>
rect 174 141 175 142 
<< pdiffusion >>
rect 175 141 176 142 
<< pdiffusion >>
rect 176 141 177 142 
<< pdiffusion >>
rect 177 141 178 142 
<< pdiffusion >>
rect 178 141 179 142 
<< pdiffusion >>
rect 179 141 180 142 
<< m1 >>
rect 181 141 182 142 
<< m2 >>
rect 182 141 183 142 
<< m1 >>
rect 190 141 191 142 
<< pdiffusion >>
rect 192 141 193 142 
<< pdiffusion >>
rect 193 141 194 142 
<< pdiffusion >>
rect 194 141 195 142 
<< pdiffusion >>
rect 195 141 196 142 
<< pdiffusion >>
rect 196 141 197 142 
<< pdiffusion >>
rect 197 141 198 142 
<< m1 >>
rect 199 141 200 142 
<< m1 >>
rect 201 141 202 142 
<< m1 >>
rect 203 141 204 142 
<< pdiffusion >>
rect 210 141 211 142 
<< pdiffusion >>
rect 211 141 212 142 
<< pdiffusion >>
rect 212 141 213 142 
<< pdiffusion >>
rect 213 141 214 142 
<< pdiffusion >>
rect 214 141 215 142 
<< pdiffusion >>
rect 215 141 216 142 
<< m1 >>
rect 226 141 227 142 
<< m2 >>
rect 226 141 227 142 
<< pdiffusion >>
rect 228 141 229 142 
<< pdiffusion >>
rect 229 141 230 142 
<< pdiffusion >>
rect 230 141 231 142 
<< pdiffusion >>
rect 231 141 232 142 
<< pdiffusion >>
rect 232 141 233 142 
<< pdiffusion >>
rect 233 141 234 142 
<< pdiffusion >>
rect 246 141 247 142 
<< pdiffusion >>
rect 247 141 248 142 
<< pdiffusion >>
rect 248 141 249 142 
<< pdiffusion >>
rect 249 141 250 142 
<< pdiffusion >>
rect 250 141 251 142 
<< pdiffusion >>
rect 251 141 252 142 
<< m1 >>
rect 253 141 254 142 
<< m2 >>
rect 254 141 255 142 
<< m1 >>
rect 256 141 257 142 
<< m1 >>
rect 19 142 20 143 
<< m1 >>
rect 28 142 29 143 
<< m2 >>
rect 28 142 29 143 
<< pdiffusion >>
rect 30 142 31 143 
<< pdiffusion >>
rect 31 142 32 143 
<< pdiffusion >>
rect 32 142 33 143 
<< pdiffusion >>
rect 33 142 34 143 
<< pdiffusion >>
rect 34 142 35 143 
<< pdiffusion >>
rect 35 142 36 143 
<< m1 >>
rect 44 142 45 143 
<< m1 >>
rect 46 142 47 143 
<< pdiffusion >>
rect 48 142 49 143 
<< pdiffusion >>
rect 49 142 50 143 
<< pdiffusion >>
rect 50 142 51 143 
<< pdiffusion >>
rect 51 142 52 143 
<< pdiffusion >>
rect 52 142 53 143 
<< pdiffusion >>
rect 53 142 54 143 
<< m1 >>
rect 55 142 56 143 
<< m1 >>
rect 57 142 58 143 
<< m1 >>
rect 62 142 63 143 
<< m1 >>
rect 64 142 65 143 
<< pdiffusion >>
rect 66 142 67 143 
<< pdiffusion >>
rect 67 142 68 143 
<< pdiffusion >>
rect 68 142 69 143 
<< pdiffusion >>
rect 69 142 70 143 
<< pdiffusion >>
rect 70 142 71 143 
<< pdiffusion >>
rect 71 142 72 143 
<< m1 >>
rect 73 142 74 143 
<< m2 >>
rect 74 142 75 143 
<< m1 >>
rect 75 142 76 143 
<< m1 >>
rect 77 142 78 143 
<< m1 >>
rect 82 142 83 143 
<< pdiffusion >>
rect 84 142 85 143 
<< pdiffusion >>
rect 85 142 86 143 
<< pdiffusion >>
rect 86 142 87 143 
<< pdiffusion >>
rect 87 142 88 143 
<< pdiffusion >>
rect 88 142 89 143 
<< pdiffusion >>
rect 89 142 90 143 
<< m1 >>
rect 91 142 92 143 
<< m2 >>
rect 117 142 118 143 
<< m1 >>
rect 118 142 119 143 
<< pdiffusion >>
rect 120 142 121 143 
<< pdiffusion >>
rect 121 142 122 143 
<< pdiffusion >>
rect 122 142 123 143 
<< pdiffusion >>
rect 123 142 124 143 
<< pdiffusion >>
rect 124 142 125 143 
<< pdiffusion >>
rect 125 142 126 143 
<< m1 >>
rect 129 142 130 143 
<< m1 >>
rect 131 142 132 143 
<< pdiffusion >>
rect 138 142 139 143 
<< pdiffusion >>
rect 139 142 140 143 
<< pdiffusion >>
rect 140 142 141 143 
<< pdiffusion >>
rect 141 142 142 143 
<< pdiffusion >>
rect 142 142 143 143 
<< pdiffusion >>
rect 143 142 144 143 
<< m1 >>
rect 145 142 146 143 
<< pdiffusion >>
rect 156 142 157 143 
<< pdiffusion >>
rect 157 142 158 143 
<< pdiffusion >>
rect 158 142 159 143 
<< pdiffusion >>
rect 159 142 160 143 
<< pdiffusion >>
rect 160 142 161 143 
<< pdiffusion >>
rect 161 142 162 143 
<< m1 >>
rect 163 142 164 143 
<< m1 >>
rect 165 142 166 143 
<< m2 >>
rect 166 142 167 143 
<< m1 >>
rect 169 142 170 143 
<< m2 >>
rect 169 142 170 143 
<< m2c >>
rect 169 142 170 143 
<< m1 >>
rect 169 142 170 143 
<< m2 >>
rect 169 142 170 143 
<< pdiffusion >>
rect 174 142 175 143 
<< pdiffusion >>
rect 175 142 176 143 
<< pdiffusion >>
rect 176 142 177 143 
<< pdiffusion >>
rect 177 142 178 143 
<< pdiffusion >>
rect 178 142 179 143 
<< pdiffusion >>
rect 179 142 180 143 
<< m1 >>
rect 181 142 182 143 
<< m2 >>
rect 182 142 183 143 
<< m1 >>
rect 190 142 191 143 
<< pdiffusion >>
rect 192 142 193 143 
<< pdiffusion >>
rect 193 142 194 143 
<< pdiffusion >>
rect 194 142 195 143 
<< pdiffusion >>
rect 195 142 196 143 
<< pdiffusion >>
rect 196 142 197 143 
<< pdiffusion >>
rect 197 142 198 143 
<< m1 >>
rect 199 142 200 143 
<< m1 >>
rect 201 142 202 143 
<< m1 >>
rect 203 142 204 143 
<< pdiffusion >>
rect 210 142 211 143 
<< pdiffusion >>
rect 211 142 212 143 
<< pdiffusion >>
rect 212 142 213 143 
<< pdiffusion >>
rect 213 142 214 143 
<< pdiffusion >>
rect 214 142 215 143 
<< pdiffusion >>
rect 215 142 216 143 
<< m1 >>
rect 226 142 227 143 
<< m2 >>
rect 226 142 227 143 
<< pdiffusion >>
rect 228 142 229 143 
<< pdiffusion >>
rect 229 142 230 143 
<< pdiffusion >>
rect 230 142 231 143 
<< pdiffusion >>
rect 231 142 232 143 
<< pdiffusion >>
rect 232 142 233 143 
<< pdiffusion >>
rect 233 142 234 143 
<< pdiffusion >>
rect 246 142 247 143 
<< pdiffusion >>
rect 247 142 248 143 
<< pdiffusion >>
rect 248 142 249 143 
<< pdiffusion >>
rect 249 142 250 143 
<< pdiffusion >>
rect 250 142 251 143 
<< pdiffusion >>
rect 251 142 252 143 
<< m1 >>
rect 253 142 254 143 
<< m2 >>
rect 254 142 255 143 
<< m1 >>
rect 256 142 257 143 
<< m1 >>
rect 19 143 20 144 
<< m1 >>
rect 28 143 29 144 
<< m2 >>
rect 28 143 29 144 
<< pdiffusion >>
rect 30 143 31 144 
<< pdiffusion >>
rect 31 143 32 144 
<< pdiffusion >>
rect 32 143 33 144 
<< pdiffusion >>
rect 33 143 34 144 
<< m1 >>
rect 34 143 35 144 
<< pdiffusion >>
rect 34 143 35 144 
<< pdiffusion >>
rect 35 143 36 144 
<< m1 >>
rect 44 143 45 144 
<< m1 >>
rect 46 143 47 144 
<< pdiffusion >>
rect 48 143 49 144 
<< pdiffusion >>
rect 49 143 50 144 
<< pdiffusion >>
rect 50 143 51 144 
<< pdiffusion >>
rect 51 143 52 144 
<< m1 >>
rect 52 143 53 144 
<< pdiffusion >>
rect 52 143 53 144 
<< pdiffusion >>
rect 53 143 54 144 
<< m1 >>
rect 55 143 56 144 
<< m1 >>
rect 57 143 58 144 
<< m1 >>
rect 62 143 63 144 
<< m1 >>
rect 64 143 65 144 
<< pdiffusion >>
rect 66 143 67 144 
<< m1 >>
rect 67 143 68 144 
<< pdiffusion >>
rect 67 143 68 144 
<< pdiffusion >>
rect 68 143 69 144 
<< pdiffusion >>
rect 69 143 70 144 
<< pdiffusion >>
rect 70 143 71 144 
<< pdiffusion >>
rect 71 143 72 144 
<< m1 >>
rect 73 143 74 144 
<< m2 >>
rect 74 143 75 144 
<< m1 >>
rect 75 143 76 144 
<< m1 >>
rect 77 143 78 144 
<< m1 >>
rect 82 143 83 144 
<< pdiffusion >>
rect 84 143 85 144 
<< pdiffusion >>
rect 85 143 86 144 
<< pdiffusion >>
rect 86 143 87 144 
<< pdiffusion >>
rect 87 143 88 144 
<< m1 >>
rect 88 143 89 144 
<< pdiffusion >>
rect 88 143 89 144 
<< pdiffusion >>
rect 89 143 90 144 
<< m1 >>
rect 91 143 92 144 
<< m2 >>
rect 117 143 118 144 
<< m1 >>
rect 118 143 119 144 
<< pdiffusion >>
rect 120 143 121 144 
<< pdiffusion >>
rect 121 143 122 144 
<< pdiffusion >>
rect 122 143 123 144 
<< pdiffusion >>
rect 123 143 124 144 
<< m1 >>
rect 124 143 125 144 
<< pdiffusion >>
rect 124 143 125 144 
<< pdiffusion >>
rect 125 143 126 144 
<< m1 >>
rect 129 143 130 144 
<< m1 >>
rect 131 143 132 144 
<< pdiffusion >>
rect 138 143 139 144 
<< pdiffusion >>
rect 139 143 140 144 
<< pdiffusion >>
rect 140 143 141 144 
<< pdiffusion >>
rect 141 143 142 144 
<< pdiffusion >>
rect 142 143 143 144 
<< pdiffusion >>
rect 143 143 144 144 
<< m1 >>
rect 145 143 146 144 
<< pdiffusion >>
rect 156 143 157 144 
<< m1 >>
rect 157 143 158 144 
<< pdiffusion >>
rect 157 143 158 144 
<< pdiffusion >>
rect 158 143 159 144 
<< pdiffusion >>
rect 159 143 160 144 
<< pdiffusion >>
rect 160 143 161 144 
<< pdiffusion >>
rect 161 143 162 144 
<< m1 >>
rect 163 143 164 144 
<< m1 >>
rect 165 143 166 144 
<< m2 >>
rect 166 143 167 144 
<< m2 >>
rect 169 143 170 144 
<< pdiffusion >>
rect 174 143 175 144 
<< pdiffusion >>
rect 175 143 176 144 
<< pdiffusion >>
rect 176 143 177 144 
<< pdiffusion >>
rect 177 143 178 144 
<< m1 >>
rect 178 143 179 144 
<< pdiffusion >>
rect 178 143 179 144 
<< pdiffusion >>
rect 179 143 180 144 
<< m1 >>
rect 181 143 182 144 
<< m2 >>
rect 182 143 183 144 
<< m1 >>
rect 190 143 191 144 
<< pdiffusion >>
rect 192 143 193 144 
<< pdiffusion >>
rect 193 143 194 144 
<< pdiffusion >>
rect 194 143 195 144 
<< pdiffusion >>
rect 195 143 196 144 
<< m1 >>
rect 196 143 197 144 
<< pdiffusion >>
rect 196 143 197 144 
<< pdiffusion >>
rect 197 143 198 144 
<< m1 >>
rect 199 143 200 144 
<< m1 >>
rect 201 143 202 144 
<< m1 >>
rect 203 143 204 144 
<< pdiffusion >>
rect 210 143 211 144 
<< pdiffusion >>
rect 211 143 212 144 
<< pdiffusion >>
rect 212 143 213 144 
<< pdiffusion >>
rect 213 143 214 144 
<< pdiffusion >>
rect 214 143 215 144 
<< pdiffusion >>
rect 215 143 216 144 
<< m1 >>
rect 226 143 227 144 
<< m2 >>
rect 226 143 227 144 
<< pdiffusion >>
rect 228 143 229 144 
<< pdiffusion >>
rect 229 143 230 144 
<< pdiffusion >>
rect 230 143 231 144 
<< pdiffusion >>
rect 231 143 232 144 
<< pdiffusion >>
rect 232 143 233 144 
<< pdiffusion >>
rect 233 143 234 144 
<< pdiffusion >>
rect 246 143 247 144 
<< pdiffusion >>
rect 247 143 248 144 
<< pdiffusion >>
rect 248 143 249 144 
<< pdiffusion >>
rect 249 143 250 144 
<< m1 >>
rect 250 143 251 144 
<< pdiffusion >>
rect 250 143 251 144 
<< pdiffusion >>
rect 251 143 252 144 
<< m1 >>
rect 253 143 254 144 
<< m2 >>
rect 254 143 255 144 
<< m1 >>
rect 256 143 257 144 
<< m1 >>
rect 19 144 20 145 
<< m1 >>
rect 28 144 29 145 
<< m2 >>
rect 28 144 29 145 
<< m1 >>
rect 34 144 35 145 
<< m1 >>
rect 44 144 45 145 
<< m1 >>
rect 46 144 47 145 
<< m1 >>
rect 52 144 53 145 
<< m1 >>
rect 55 144 56 145 
<< m1 >>
rect 57 144 58 145 
<< m1 >>
rect 62 144 63 145 
<< m1 >>
rect 64 144 65 145 
<< m1 >>
rect 67 144 68 145 
<< m1 >>
rect 73 144 74 145 
<< m2 >>
rect 74 144 75 145 
<< m1 >>
rect 75 144 76 145 
<< m1 >>
rect 77 144 78 145 
<< m1 >>
rect 82 144 83 145 
<< m1 >>
rect 88 144 89 145 
<< m1 >>
rect 91 144 92 145 
<< m2 >>
rect 91 144 92 145 
<< m2c >>
rect 91 144 92 145 
<< m1 >>
rect 91 144 92 145 
<< m2 >>
rect 91 144 92 145 
<< m2 >>
rect 117 144 118 145 
<< m1 >>
rect 118 144 119 145 
<< m1 >>
rect 124 144 125 145 
<< m1 >>
rect 129 144 130 145 
<< m1 >>
rect 131 144 132 145 
<< m1 >>
rect 145 144 146 145 
<< m1 >>
rect 157 144 158 145 
<< m1 >>
rect 163 144 164 145 
<< m1 >>
rect 165 144 166 145 
<< m2 >>
rect 166 144 167 145 
<< m1 >>
rect 167 144 168 145 
<< m2 >>
rect 167 144 168 145 
<< m2c >>
rect 167 144 168 145 
<< m1 >>
rect 167 144 168 145 
<< m2 >>
rect 167 144 168 145 
<< m1 >>
rect 168 144 169 145 
<< m1 >>
rect 169 144 170 145 
<< m2 >>
rect 169 144 170 145 
<< m1 >>
rect 170 144 171 145 
<< m1 >>
rect 171 144 172 145 
<< m1 >>
rect 172 144 173 145 
<< m1 >>
rect 178 144 179 145 
<< m1 >>
rect 181 144 182 145 
<< m2 >>
rect 182 144 183 145 
<< m1 >>
rect 190 144 191 145 
<< m1 >>
rect 196 144 197 145 
<< m1 >>
rect 199 144 200 145 
<< m1 >>
rect 201 144 202 145 
<< m1 >>
rect 203 144 204 145 
<< m1 >>
rect 226 144 227 145 
<< m2 >>
rect 226 144 227 145 
<< m1 >>
rect 250 144 251 145 
<< m1 >>
rect 253 144 254 145 
<< m2 >>
rect 254 144 255 145 
<< m1 >>
rect 256 144 257 145 
<< m1 >>
rect 19 145 20 146 
<< m1 >>
rect 28 145 29 146 
<< m2 >>
rect 28 145 29 146 
<< m1 >>
rect 34 145 35 146 
<< m1 >>
rect 44 145 45 146 
<< m1 >>
rect 46 145 47 146 
<< m1 >>
rect 52 145 53 146 
<< m1 >>
rect 55 145 56 146 
<< m1 >>
rect 57 145 58 146 
<< m1 >>
rect 62 145 63 146 
<< m1 >>
rect 64 145 65 146 
<< m1 >>
rect 67 145 68 146 
<< m1 >>
rect 71 145 72 146 
<< m2 >>
rect 71 145 72 146 
<< m2c >>
rect 71 145 72 146 
<< m1 >>
rect 71 145 72 146 
<< m2 >>
rect 71 145 72 146 
<< m2 >>
rect 72 145 73 146 
<< m1 >>
rect 73 145 74 146 
<< m2 >>
rect 73 145 74 146 
<< m2 >>
rect 74 145 75 146 
<< m1 >>
rect 75 145 76 146 
<< m1 >>
rect 77 145 78 146 
<< m1 >>
rect 82 145 83 146 
<< m1 >>
rect 88 145 89 146 
<< m2 >>
rect 88 145 89 146 
<< m2c >>
rect 88 145 89 146 
<< m1 >>
rect 88 145 89 146 
<< m2 >>
rect 88 145 89 146 
<< m2 >>
rect 91 145 92 146 
<< m2 >>
rect 117 145 118 146 
<< m1 >>
rect 118 145 119 146 
<< m1 >>
rect 124 145 125 146 
<< m1 >>
rect 125 145 126 146 
<< m1 >>
rect 126 145 127 146 
<< m1 >>
rect 127 145 128 146 
<< m1 >>
rect 128 145 129 146 
<< m1 >>
rect 129 145 130 146 
<< m1 >>
rect 131 145 132 146 
<< m1 >>
rect 145 145 146 146 
<< m1 >>
rect 157 145 158 146 
<< m1 >>
rect 163 145 164 146 
<< m1 >>
rect 165 145 166 146 
<< m2 >>
rect 169 145 170 146 
<< m1 >>
rect 172 145 173 146 
<< m1 >>
rect 178 145 179 146 
<< m1 >>
rect 181 145 182 146 
<< m2 >>
rect 182 145 183 146 
<< m1 >>
rect 190 145 191 146 
<< m1 >>
rect 196 145 197 146 
<< m1 >>
rect 199 145 200 146 
<< m1 >>
rect 201 145 202 146 
<< m1 >>
rect 203 145 204 146 
<< m1 >>
rect 226 145 227 146 
<< m2 >>
rect 226 145 227 146 
<< m1 >>
rect 250 145 251 146 
<< m1 >>
rect 253 145 254 146 
<< m2 >>
rect 254 145 255 146 
<< m1 >>
rect 256 145 257 146 
<< m1 >>
rect 19 146 20 147 
<< m1 >>
rect 28 146 29 147 
<< m2 >>
rect 28 146 29 147 
<< m1 >>
rect 34 146 35 147 
<< m1 >>
rect 44 146 45 147 
<< m1 >>
rect 46 146 47 147 
<< m1 >>
rect 52 146 53 147 
<< m1 >>
rect 55 146 56 147 
<< m1 >>
rect 57 146 58 147 
<< m1 >>
rect 62 146 63 147 
<< m1 >>
rect 64 146 65 147 
<< m1 >>
rect 67 146 68 147 
<< m1 >>
rect 68 146 69 147 
<< m1 >>
rect 69 146 70 147 
<< m2 >>
rect 69 146 70 147 
<< m2c >>
rect 69 146 70 147 
<< m1 >>
rect 69 146 70 147 
<< m2 >>
rect 69 146 70 147 
<< m1 >>
rect 71 146 72 147 
<< m1 >>
rect 73 146 74 147 
<< m1 >>
rect 75 146 76 147 
<< m1 >>
rect 77 146 78 147 
<< m1 >>
rect 82 146 83 147 
<< m1 >>
rect 88 146 89 147 
<< m1 >>
rect 89 146 90 147 
<< m2 >>
rect 89 146 90 147 
<< m1 >>
rect 90 146 91 147 
<< m2 >>
rect 90 146 91 147 
<< m1 >>
rect 91 146 92 147 
<< m2 >>
rect 91 146 92 147 
<< m1 >>
rect 92 146 93 147 
<< m1 >>
rect 93 146 94 147 
<< m1 >>
rect 94 146 95 147 
<< m1 >>
rect 95 146 96 147 
<< m1 >>
rect 96 146 97 147 
<< m1 >>
rect 97 146 98 147 
<< m1 >>
rect 98 146 99 147 
<< m1 >>
rect 99 146 100 147 
<< m1 >>
rect 100 146 101 147 
<< m1 >>
rect 101 146 102 147 
<< m1 >>
rect 102 146 103 147 
<< m1 >>
rect 103 146 104 147 
<< m1 >>
rect 104 146 105 147 
<< m1 >>
rect 105 146 106 147 
<< m1 >>
rect 106 146 107 147 
<< m1 >>
rect 107 146 108 147 
<< m1 >>
rect 108 146 109 147 
<< m1 >>
rect 109 146 110 147 
<< m1 >>
rect 110 146 111 147 
<< m1 >>
rect 111 146 112 147 
<< m1 >>
rect 112 146 113 147 
<< m1 >>
rect 113 146 114 147 
<< m1 >>
rect 114 146 115 147 
<< m1 >>
rect 115 146 116 147 
<< m1 >>
rect 116 146 117 147 
<< m1 >>
rect 117 146 118 147 
<< m2 >>
rect 117 146 118 147 
<< m1 >>
rect 118 146 119 147 
<< m2 >>
rect 123 146 124 147 
<< m2 >>
rect 124 146 125 147 
<< m2 >>
rect 125 146 126 147 
<< m2 >>
rect 126 146 127 147 
<< m2 >>
rect 127 146 128 147 
<< m2 >>
rect 128 146 129 147 
<< m2 >>
rect 129 146 130 147 
<< m2 >>
rect 130 146 131 147 
<< m1 >>
rect 131 146 132 147 
<< m2 >>
rect 131 146 132 147 
<< m2c >>
rect 131 146 132 147 
<< m1 >>
rect 131 146 132 147 
<< m2 >>
rect 131 146 132 147 
<< m1 >>
rect 145 146 146 147 
<< m1 >>
rect 157 146 158 147 
<< m1 >>
rect 158 146 159 147 
<< m1 >>
rect 159 146 160 147 
<< m1 >>
rect 160 146 161 147 
<< m1 >>
rect 161 146 162 147 
<< m2 >>
rect 161 146 162 147 
<< m2c >>
rect 161 146 162 147 
<< m1 >>
rect 161 146 162 147 
<< m2 >>
rect 161 146 162 147 
<< m1 >>
rect 163 146 164 147 
<< m2 >>
rect 163 146 164 147 
<< m2c >>
rect 163 146 164 147 
<< m1 >>
rect 163 146 164 147 
<< m2 >>
rect 163 146 164 147 
<< m1 >>
rect 165 146 166 147 
<< m2 >>
rect 165 146 166 147 
<< m2c >>
rect 165 146 166 147 
<< m1 >>
rect 165 146 166 147 
<< m2 >>
rect 165 146 166 147 
<< m1 >>
rect 169 146 170 147 
<< m2 >>
rect 169 146 170 147 
<< m2c >>
rect 169 146 170 147 
<< m1 >>
rect 169 146 170 147 
<< m2 >>
rect 169 146 170 147 
<< m1 >>
rect 172 146 173 147 
<< m1 >>
rect 173 146 174 147 
<< m1 >>
rect 174 146 175 147 
<< m2 >>
rect 174 146 175 147 
<< m2c >>
rect 174 146 175 147 
<< m1 >>
rect 174 146 175 147 
<< m2 >>
rect 174 146 175 147 
<< m1 >>
rect 178 146 179 147 
<< m1 >>
rect 181 146 182 147 
<< m2 >>
rect 182 146 183 147 
<< m1 >>
rect 190 146 191 147 
<< m1 >>
rect 196 146 197 147 
<< m2 >>
rect 198 146 199 147 
<< m1 >>
rect 199 146 200 147 
<< m2 >>
rect 199 146 200 147 
<< m2 >>
rect 200 146 201 147 
<< m1 >>
rect 201 146 202 147 
<< m2 >>
rect 201 146 202 147 
<< m2 >>
rect 202 146 203 147 
<< m1 >>
rect 203 146 204 147 
<< m2 >>
rect 203 146 204 147 
<< m2c >>
rect 203 146 204 147 
<< m1 >>
rect 203 146 204 147 
<< m2 >>
rect 203 146 204 147 
<< m1 >>
rect 226 146 227 147 
<< m2 >>
rect 226 146 227 147 
<< m1 >>
rect 227 146 228 147 
<< m1 >>
rect 228 146 229 147 
<< m2 >>
rect 228 146 229 147 
<< m2c >>
rect 228 146 229 147 
<< m1 >>
rect 228 146 229 147 
<< m2 >>
rect 228 146 229 147 
<< m1 >>
rect 250 146 251 147 
<< m1 >>
rect 253 146 254 147 
<< m2 >>
rect 254 146 255 147 
<< m1 >>
rect 256 146 257 147 
<< m1 >>
rect 19 147 20 148 
<< m1 >>
rect 28 147 29 148 
<< m2 >>
rect 28 147 29 148 
<< m1 >>
rect 34 147 35 148 
<< m1 >>
rect 44 147 45 148 
<< m1 >>
rect 46 147 47 148 
<< m1 >>
rect 52 147 53 148 
<< m1 >>
rect 55 147 56 148 
<< m1 >>
rect 57 147 58 148 
<< m1 >>
rect 62 147 63 148 
<< m1 >>
rect 64 147 65 148 
<< m2 >>
rect 69 147 70 148 
<< m2 >>
rect 70 147 71 148 
<< m1 >>
rect 71 147 72 148 
<< m2 >>
rect 71 147 72 148 
<< m2 >>
rect 72 147 73 148 
<< m1 >>
rect 73 147 74 148 
<< m2 >>
rect 73 147 74 148 
<< m2 >>
rect 74 147 75 148 
<< m1 >>
rect 75 147 76 148 
<< m2 >>
rect 75 147 76 148 
<< m2c >>
rect 75 147 76 148 
<< m1 >>
rect 75 147 76 148 
<< m2 >>
rect 75 147 76 148 
<< m1 >>
rect 77 147 78 148 
<< m1 >>
rect 82 147 83 148 
<< m1 >>
rect 88 147 89 148 
<< m2 >>
rect 89 147 90 148 
<< m2 >>
rect 91 147 92 148 
<< m2 >>
rect 92 147 93 148 
<< m2 >>
rect 93 147 94 148 
<< m2 >>
rect 94 147 95 148 
<< m2 >>
rect 95 147 96 148 
<< m2 >>
rect 96 147 97 148 
<< m2 >>
rect 97 147 98 148 
<< m2 >>
rect 98 147 99 148 
<< m2 >>
rect 99 147 100 148 
<< m2 >>
rect 100 147 101 148 
<< m2 >>
rect 101 147 102 148 
<< m2 >>
rect 102 147 103 148 
<< m2 >>
rect 103 147 104 148 
<< m2 >>
rect 104 147 105 148 
<< m2 >>
rect 105 147 106 148 
<< m2 >>
rect 106 147 107 148 
<< m2 >>
rect 107 147 108 148 
<< m2 >>
rect 108 147 109 148 
<< m2 >>
rect 109 147 110 148 
<< m2 >>
rect 110 147 111 148 
<< m2 >>
rect 111 147 112 148 
<< m2 >>
rect 112 147 113 148 
<< m2 >>
rect 113 147 114 148 
<< m2 >>
rect 114 147 115 148 
<< m2 >>
rect 115 147 116 148 
<< m2 >>
rect 116 147 117 148 
<< m2 >>
rect 117 147 118 148 
<< m2 >>
rect 123 147 124 148 
<< m1 >>
rect 145 147 146 148 
<< m2 >>
rect 161 147 162 148 
<< m2 >>
rect 163 147 164 148 
<< m2 >>
rect 165 147 166 148 
<< m2 >>
rect 169 147 170 148 
<< m2 >>
rect 174 147 175 148 
<< m1 >>
rect 178 147 179 148 
<< m1 >>
rect 181 147 182 148 
<< m2 >>
rect 182 147 183 148 
<< m1 >>
rect 183 147 184 148 
<< m2 >>
rect 183 147 184 148 
<< m2c >>
rect 183 147 184 148 
<< m1 >>
rect 183 147 184 148 
<< m2 >>
rect 183 147 184 148 
<< m1 >>
rect 184 147 185 148 
<< m1 >>
rect 185 147 186 148 
<< m1 >>
rect 186 147 187 148 
<< m1 >>
rect 187 147 188 148 
<< m1 >>
rect 188 147 189 148 
<< m1 >>
rect 190 147 191 148 
<< m1 >>
rect 196 147 197 148 
<< m2 >>
rect 198 147 199 148 
<< m1 >>
rect 199 147 200 148 
<< m1 >>
rect 201 147 202 148 
<< m2 >>
rect 226 147 227 148 
<< m2 >>
rect 228 147 229 148 
<< m1 >>
rect 250 147 251 148 
<< m1 >>
rect 253 147 254 148 
<< m2 >>
rect 254 147 255 148 
<< m1 >>
rect 256 147 257 148 
<< m1 >>
rect 19 148 20 149 
<< m1 >>
rect 28 148 29 149 
<< m2 >>
rect 28 148 29 149 
<< m1 >>
rect 34 148 35 149 
<< m1 >>
rect 44 148 45 149 
<< m1 >>
rect 46 148 47 149 
<< m1 >>
rect 47 148 48 149 
<< m1 >>
rect 48 148 49 149 
<< m1 >>
rect 49 148 50 149 
<< m1 >>
rect 50 148 51 149 
<< m1 >>
rect 51 148 52 149 
<< m1 >>
rect 52 148 53 149 
<< m1 >>
rect 55 148 56 149 
<< m1 >>
rect 57 148 58 149 
<< m1 >>
rect 62 148 63 149 
<< m2 >>
rect 62 148 63 149 
<< m2c >>
rect 62 148 63 149 
<< m1 >>
rect 62 148 63 149 
<< m2 >>
rect 62 148 63 149 
<< m2 >>
rect 63 148 64 149 
<< m1 >>
rect 64 148 65 149 
<< m2 >>
rect 64 148 65 149 
<< m2 >>
rect 65 148 66 149 
<< m1 >>
rect 66 148 67 149 
<< m2 >>
rect 66 148 67 149 
<< m2c >>
rect 66 148 67 149 
<< m1 >>
rect 66 148 67 149 
<< m2 >>
rect 66 148 67 149 
<< m1 >>
rect 67 148 68 149 
<< m1 >>
rect 68 148 69 149 
<< m1 >>
rect 69 148 70 149 
<< m1 >>
rect 70 148 71 149 
<< m1 >>
rect 71 148 72 149 
<< m1 >>
rect 73 148 74 149 
<< m1 >>
rect 77 148 78 149 
<< m1 >>
rect 82 148 83 149 
<< m1 >>
rect 88 148 89 149 
<< m2 >>
rect 89 148 90 149 
<< m1 >>
rect 91 148 92 149 
<< m2 >>
rect 91 148 92 149 
<< m2c >>
rect 91 148 92 149 
<< m1 >>
rect 91 148 92 149 
<< m2 >>
rect 91 148 92 149 
<< m1 >>
rect 121 148 122 149 
<< m1 >>
rect 122 148 123 149 
<< m1 >>
rect 123 148 124 149 
<< m2 >>
rect 123 148 124 149 
<< m1 >>
rect 124 148 125 149 
<< m1 >>
rect 125 148 126 149 
<< m1 >>
rect 126 148 127 149 
<< m1 >>
rect 127 148 128 149 
<< m1 >>
rect 128 148 129 149 
<< m1 >>
rect 129 148 130 149 
<< m1 >>
rect 130 148 131 149 
<< m1 >>
rect 131 148 132 149 
<< m1 >>
rect 132 148 133 149 
<< m1 >>
rect 133 148 134 149 
<< m1 >>
rect 134 148 135 149 
<< m1 >>
rect 135 148 136 149 
<< m1 >>
rect 136 148 137 149 
<< m1 >>
rect 137 148 138 149 
<< m1 >>
rect 138 148 139 149 
<< m1 >>
rect 139 148 140 149 
<< m1 >>
rect 140 148 141 149 
<< m1 >>
rect 141 148 142 149 
<< m1 >>
rect 142 148 143 149 
<< m1 >>
rect 143 148 144 149 
<< m2 >>
rect 143 148 144 149 
<< m2c >>
rect 143 148 144 149 
<< m1 >>
rect 143 148 144 149 
<< m2 >>
rect 143 148 144 149 
<< m2 >>
rect 144 148 145 149 
<< m1 >>
rect 145 148 146 149 
<< m2 >>
rect 145 148 146 149 
<< m2 >>
rect 146 148 147 149 
<< m1 >>
rect 147 148 148 149 
<< m2 >>
rect 147 148 148 149 
<< m2c >>
rect 147 148 148 149 
<< m1 >>
rect 147 148 148 149 
<< m2 >>
rect 147 148 148 149 
<< m1 >>
rect 148 148 149 149 
<< m1 >>
rect 149 148 150 149 
<< m1 >>
rect 150 148 151 149 
<< m1 >>
rect 151 148 152 149 
<< m1 >>
rect 152 148 153 149 
<< m1 >>
rect 153 148 154 149 
<< m1 >>
rect 154 148 155 149 
<< m1 >>
rect 155 148 156 149 
<< m1 >>
rect 156 148 157 149 
<< m1 >>
rect 157 148 158 149 
<< m1 >>
rect 158 148 159 149 
<< m1 >>
rect 159 148 160 149 
<< m1 >>
rect 160 148 161 149 
<< m1 >>
rect 161 148 162 149 
<< m2 >>
rect 161 148 162 149 
<< m1 >>
rect 162 148 163 149 
<< m1 >>
rect 163 148 164 149 
<< m2 >>
rect 163 148 164 149 
<< m1 >>
rect 164 148 165 149 
<< m1 >>
rect 165 148 166 149 
<< m2 >>
rect 165 148 166 149 
<< m1 >>
rect 166 148 167 149 
<< m1 >>
rect 167 148 168 149 
<< m1 >>
rect 168 148 169 149 
<< m1 >>
rect 169 148 170 149 
<< m2 >>
rect 169 148 170 149 
<< m1 >>
rect 170 148 171 149 
<< m1 >>
rect 171 148 172 149 
<< m1 >>
rect 172 148 173 149 
<< m1 >>
rect 173 148 174 149 
<< m1 >>
rect 174 148 175 149 
<< m2 >>
rect 174 148 175 149 
<< m1 >>
rect 175 148 176 149 
<< m1 >>
rect 176 148 177 149 
<< m1 >>
rect 177 148 178 149 
<< m1 >>
rect 178 148 179 149 
<< m1 >>
rect 181 148 182 149 
<< m1 >>
rect 188 148 189 149 
<< m2 >>
rect 188 148 189 149 
<< m2c >>
rect 188 148 189 149 
<< m1 >>
rect 188 148 189 149 
<< m2 >>
rect 188 148 189 149 
<< m2 >>
rect 189 148 190 149 
<< m1 >>
rect 190 148 191 149 
<< m2 >>
rect 190 148 191 149 
<< m2 >>
rect 191 148 192 149 
<< m1 >>
rect 192 148 193 149 
<< m2 >>
rect 192 148 193 149 
<< m2c >>
rect 192 148 193 149 
<< m1 >>
rect 192 148 193 149 
<< m2 >>
rect 192 148 193 149 
<< m1 >>
rect 193 148 194 149 
<< m1 >>
rect 194 148 195 149 
<< m1 >>
rect 195 148 196 149 
<< m1 >>
rect 196 148 197 149 
<< m2 >>
rect 198 148 199 149 
<< m1 >>
rect 199 148 200 149 
<< m1 >>
rect 201 148 202 149 
<< m1 >>
rect 202 148 203 149 
<< m1 >>
rect 203 148 204 149 
<< m1 >>
rect 204 148 205 149 
<< m1 >>
rect 205 148 206 149 
<< m1 >>
rect 206 148 207 149 
<< m1 >>
rect 207 148 208 149 
<< m1 >>
rect 208 148 209 149 
<< m1 >>
rect 209 148 210 149 
<< m1 >>
rect 210 148 211 149 
<< m1 >>
rect 211 148 212 149 
<< m1 >>
rect 212 148 213 149 
<< m1 >>
rect 213 148 214 149 
<< m1 >>
rect 214 148 215 149 
<< m1 >>
rect 215 148 216 149 
<< m1 >>
rect 216 148 217 149 
<< m1 >>
rect 217 148 218 149 
<< m1 >>
rect 218 148 219 149 
<< m1 >>
rect 219 148 220 149 
<< m1 >>
rect 220 148 221 149 
<< m1 >>
rect 221 148 222 149 
<< m1 >>
rect 222 148 223 149 
<< m1 >>
rect 223 148 224 149 
<< m1 >>
rect 224 148 225 149 
<< m1 >>
rect 225 148 226 149 
<< m1 >>
rect 226 148 227 149 
<< m2 >>
rect 226 148 227 149 
<< m1 >>
rect 227 148 228 149 
<< m1 >>
rect 228 148 229 149 
<< m2 >>
rect 228 148 229 149 
<< m1 >>
rect 229 148 230 149 
<< m1 >>
rect 230 148 231 149 
<< m1 >>
rect 231 148 232 149 
<< m1 >>
rect 232 148 233 149 
<< m1 >>
rect 233 148 234 149 
<< m1 >>
rect 234 148 235 149 
<< m1 >>
rect 235 148 236 149 
<< m1 >>
rect 236 148 237 149 
<< m1 >>
rect 237 148 238 149 
<< m1 >>
rect 238 148 239 149 
<< m1 >>
rect 239 148 240 149 
<< m1 >>
rect 240 148 241 149 
<< m1 >>
rect 241 148 242 149 
<< m1 >>
rect 242 148 243 149 
<< m1 >>
rect 243 148 244 149 
<< m1 >>
rect 244 148 245 149 
<< m1 >>
rect 245 148 246 149 
<< m1 >>
rect 246 148 247 149 
<< m1 >>
rect 247 148 248 149 
<< m1 >>
rect 248 148 249 149 
<< m1 >>
rect 249 148 250 149 
<< m1 >>
rect 250 148 251 149 
<< m1 >>
rect 253 148 254 149 
<< m2 >>
rect 254 148 255 149 
<< m1 >>
rect 256 148 257 149 
<< m1 >>
rect 19 149 20 150 
<< m1 >>
rect 28 149 29 150 
<< m2 >>
rect 28 149 29 150 
<< m1 >>
rect 34 149 35 150 
<< m1 >>
rect 44 149 45 150 
<< m1 >>
rect 55 149 56 150 
<< m1 >>
rect 57 149 58 150 
<< m1 >>
rect 64 149 65 150 
<< m1 >>
rect 73 149 74 150 
<< m1 >>
rect 77 149 78 150 
<< m1 >>
rect 82 149 83 150 
<< m1 >>
rect 88 149 89 150 
<< m2 >>
rect 89 149 90 150 
<< m1 >>
rect 91 149 92 150 
<< m2 >>
rect 120 149 121 150 
<< m1 >>
rect 121 149 122 150 
<< m2 >>
rect 121 149 122 150 
<< m2 >>
rect 122 149 123 150 
<< m2 >>
rect 123 149 124 150 
<< m1 >>
rect 145 149 146 150 
<< m2 >>
rect 161 149 162 150 
<< m2 >>
rect 163 149 164 150 
<< m2 >>
rect 165 149 166 150 
<< m2 >>
rect 169 149 170 150 
<< m2 >>
rect 174 149 175 150 
<< m2 >>
rect 175 149 176 150 
<< m2 >>
rect 176 149 177 150 
<< m2 >>
rect 177 149 178 150 
<< m2 >>
rect 178 149 179 150 
<< m2 >>
rect 179 149 180 150 
<< m2 >>
rect 180 149 181 150 
<< m1 >>
rect 181 149 182 150 
<< m2 >>
rect 181 149 182 150 
<< m2 >>
rect 182 149 183 150 
<< m1 >>
rect 190 149 191 150 
<< m2 >>
rect 198 149 199 150 
<< m1 >>
rect 199 149 200 150 
<< m2 >>
rect 226 149 227 150 
<< m2 >>
rect 228 149 229 150 
<< m2 >>
rect 229 149 230 150 
<< m2 >>
rect 230 149 231 150 
<< m2 >>
rect 231 149 232 150 
<< m2 >>
rect 232 149 233 150 
<< m2 >>
rect 233 149 234 150 
<< m2 >>
rect 234 149 235 150 
<< m2 >>
rect 235 149 236 150 
<< m2 >>
rect 236 149 237 150 
<< m2 >>
rect 237 149 238 150 
<< m2 >>
rect 238 149 239 150 
<< m2 >>
rect 239 149 240 150 
<< m2 >>
rect 240 149 241 150 
<< m2 >>
rect 241 149 242 150 
<< m2 >>
rect 242 149 243 150 
<< m2 >>
rect 243 149 244 150 
<< m2 >>
rect 244 149 245 150 
<< m2 >>
rect 245 149 246 150 
<< m2 >>
rect 246 149 247 150 
<< m2 >>
rect 247 149 248 150 
<< m2 >>
rect 248 149 249 150 
<< m2 >>
rect 249 149 250 150 
<< m2 >>
rect 250 149 251 150 
<< m1 >>
rect 253 149 254 150 
<< m2 >>
rect 254 149 255 150 
<< m1 >>
rect 256 149 257 150 
<< m1 >>
rect 19 150 20 151 
<< m1 >>
rect 28 150 29 151 
<< m2 >>
rect 28 150 29 151 
<< m1 >>
rect 34 150 35 151 
<< m1 >>
rect 44 150 45 151 
<< m1 >>
rect 55 150 56 151 
<< m1 >>
rect 57 150 58 151 
<< m1 >>
rect 64 150 65 151 
<< m1 >>
rect 73 150 74 151 
<< m1 >>
rect 77 150 78 151 
<< m1 >>
rect 82 150 83 151 
<< m1 >>
rect 88 150 89 151 
<< m2 >>
rect 89 150 90 151 
<< m1 >>
rect 91 150 92 151 
<< m2 >>
rect 120 150 121 151 
<< m1 >>
rect 121 150 122 151 
<< m1 >>
rect 145 150 146 151 
<< m1 >>
rect 161 150 162 151 
<< m2 >>
rect 161 150 162 151 
<< m2c >>
rect 161 150 162 151 
<< m1 >>
rect 161 150 162 151 
<< m2 >>
rect 161 150 162 151 
<< m1 >>
rect 163 150 164 151 
<< m2 >>
rect 163 150 164 151 
<< m2c >>
rect 163 150 164 151 
<< m1 >>
rect 163 150 164 151 
<< m2 >>
rect 163 150 164 151 
<< m1 >>
rect 165 150 166 151 
<< m2 >>
rect 165 150 166 151 
<< m2c >>
rect 165 150 166 151 
<< m1 >>
rect 165 150 166 151 
<< m2 >>
rect 165 150 166 151 
<< m1 >>
rect 169 150 170 151 
<< m2 >>
rect 169 150 170 151 
<< m2c >>
rect 169 150 170 151 
<< m1 >>
rect 169 150 170 151 
<< m2 >>
rect 169 150 170 151 
<< m1 >>
rect 181 150 182 151 
<< m2 >>
rect 182 150 183 151 
<< m1 >>
rect 190 150 191 151 
<< m2 >>
rect 198 150 199 151 
<< m1 >>
rect 199 150 200 151 
<< m1 >>
rect 226 150 227 151 
<< m2 >>
rect 226 150 227 151 
<< m2c >>
rect 226 150 227 151 
<< m1 >>
rect 226 150 227 151 
<< m2 >>
rect 226 150 227 151 
<< m1 >>
rect 250 150 251 151 
<< m2 >>
rect 250 150 251 151 
<< m2c >>
rect 250 150 251 151 
<< m1 >>
rect 250 150 251 151 
<< m2 >>
rect 250 150 251 151 
<< m1 >>
rect 253 150 254 151 
<< m2 >>
rect 254 150 255 151 
<< m1 >>
rect 256 150 257 151 
<< m1 >>
rect 19 151 20 152 
<< m2 >>
rect 19 151 20 152 
<< m2c >>
rect 19 151 20 152 
<< m1 >>
rect 19 151 20 152 
<< m2 >>
rect 19 151 20 152 
<< m1 >>
rect 28 151 29 152 
<< m2 >>
rect 28 151 29 152 
<< m2 >>
rect 29 151 30 152 
<< m1 >>
rect 30 151 31 152 
<< m2 >>
rect 30 151 31 152 
<< m2c >>
rect 30 151 31 152 
<< m1 >>
rect 30 151 31 152 
<< m2 >>
rect 30 151 31 152 
<< m1 >>
rect 31 151 32 152 
<< m1 >>
rect 32 151 33 152 
<< m1 >>
rect 34 151 35 152 
<< m1 >>
rect 44 151 45 152 
<< m1 >>
rect 46 151 47 152 
<< m1 >>
rect 47 151 48 152 
<< m1 >>
rect 48 151 49 152 
<< m1 >>
rect 49 151 50 152 
<< m1 >>
rect 50 151 51 152 
<< m1 >>
rect 51 151 52 152 
<< m1 >>
rect 52 151 53 152 
<< m1 >>
rect 55 151 56 152 
<< m1 >>
rect 57 151 58 152 
<< m1 >>
rect 64 151 65 152 
<< m2 >>
rect 64 151 65 152 
<< m2 >>
rect 65 151 66 152 
<< m1 >>
rect 66 151 67 152 
<< m2 >>
rect 66 151 67 152 
<< m2c >>
rect 66 151 67 152 
<< m1 >>
rect 66 151 67 152 
<< m2 >>
rect 66 151 67 152 
<< m1 >>
rect 67 151 68 152 
<< m1 >>
rect 68 151 69 152 
<< m1 >>
rect 69 151 70 152 
<< m1 >>
rect 70 151 71 152 
<< m1 >>
rect 71 151 72 152 
<< m2 >>
rect 71 151 72 152 
<< m2c >>
rect 71 151 72 152 
<< m1 >>
rect 71 151 72 152 
<< m2 >>
rect 71 151 72 152 
<< m2 >>
rect 72 151 73 152 
<< m1 >>
rect 73 151 74 152 
<< m2 >>
rect 73 151 74 152 
<< m2 >>
rect 74 151 75 152 
<< m1 >>
rect 75 151 76 152 
<< m2 >>
rect 75 151 76 152 
<< m2c >>
rect 75 151 76 152 
<< m1 >>
rect 75 151 76 152 
<< m2 >>
rect 75 151 76 152 
<< m1 >>
rect 76 151 77 152 
<< m1 >>
rect 77 151 78 152 
<< m1 >>
rect 82 151 83 152 
<< m1 >>
rect 88 151 89 152 
<< m2 >>
rect 89 151 90 152 
<< m1 >>
rect 91 151 92 152 
<< m1 >>
rect 95 151 96 152 
<< m1 >>
rect 96 151 97 152 
<< m1 >>
rect 97 151 98 152 
<< m1 >>
rect 98 151 99 152 
<< m1 >>
rect 99 151 100 152 
<< m1 >>
rect 100 151 101 152 
<< m1 >>
rect 101 151 102 152 
<< m1 >>
rect 102 151 103 152 
<< m1 >>
rect 103 151 104 152 
<< m1 >>
rect 104 151 105 152 
<< m1 >>
rect 105 151 106 152 
<< m1 >>
rect 106 151 107 152 
<< m1 >>
rect 107 151 108 152 
<< m1 >>
rect 108 151 109 152 
<< m1 >>
rect 109 151 110 152 
<< m1 >>
rect 110 151 111 152 
<< m1 >>
rect 111 151 112 152 
<< m1 >>
rect 112 151 113 152 
<< m1 >>
rect 113 151 114 152 
<< m1 >>
rect 114 151 115 152 
<< m1 >>
rect 115 151 116 152 
<< m1 >>
rect 116 151 117 152 
<< m1 >>
rect 117 151 118 152 
<< m1 >>
rect 118 151 119 152 
<< m1 >>
rect 119 151 120 152 
<< m2 >>
rect 119 151 120 152 
<< m2c >>
rect 119 151 120 152 
<< m1 >>
rect 119 151 120 152 
<< m2 >>
rect 119 151 120 152 
<< m2 >>
rect 120 151 121 152 
<< m1 >>
rect 121 151 122 152 
<< m1 >>
rect 145 151 146 152 
<< m1 >>
rect 161 151 162 152 
<< m1 >>
rect 163 151 164 152 
<< m1 >>
rect 165 151 166 152 
<< m1 >>
rect 169 151 170 152 
<< m1 >>
rect 181 151 182 152 
<< m2 >>
rect 182 151 183 152 
<< m1 >>
rect 190 151 191 152 
<< m2 >>
rect 198 151 199 152 
<< m1 >>
rect 199 151 200 152 
<< m1 >>
rect 226 151 227 152 
<< m1 >>
rect 250 151 251 152 
<< m1 >>
rect 253 151 254 152 
<< m2 >>
rect 254 151 255 152 
<< m1 >>
rect 256 151 257 152 
<< m2 >>
rect 19 152 20 153 
<< m1 >>
rect 28 152 29 153 
<< m1 >>
rect 32 152 33 153 
<< m1 >>
rect 34 152 35 153 
<< m1 >>
rect 44 152 45 153 
<< m1 >>
rect 46 152 47 153 
<< m1 >>
rect 52 152 53 153 
<< m1 >>
rect 55 152 56 153 
<< m1 >>
rect 57 152 58 153 
<< m1 >>
rect 64 152 65 153 
<< m2 >>
rect 64 152 65 153 
<< m1 >>
rect 73 152 74 153 
<< m1 >>
rect 82 152 83 153 
<< m1 >>
rect 88 152 89 153 
<< m2 >>
rect 89 152 90 153 
<< m1 >>
rect 91 152 92 153 
<< m1 >>
rect 95 152 96 153 
<< m1 >>
rect 121 152 122 153 
<< m1 >>
rect 145 152 146 153 
<< m1 >>
rect 161 152 162 153 
<< m2 >>
rect 161 152 162 153 
<< m2c >>
rect 161 152 162 153 
<< m1 >>
rect 161 152 162 153 
<< m2 >>
rect 161 152 162 153 
<< m2 >>
rect 162 152 163 153 
<< m1 >>
rect 163 152 164 153 
<< m2 >>
rect 163 152 164 153 
<< m2 >>
rect 164 152 165 153 
<< m1 >>
rect 165 152 166 153 
<< m2 >>
rect 165 152 166 153 
<< m2 >>
rect 166 152 167 153 
<< m1 >>
rect 167 152 168 153 
<< m2 >>
rect 167 152 168 153 
<< m2c >>
rect 167 152 168 153 
<< m1 >>
rect 167 152 168 153 
<< m2 >>
rect 167 152 168 153 
<< m1 >>
rect 168 152 169 153 
<< m1 >>
rect 169 152 170 153 
<< m1 >>
rect 181 152 182 153 
<< m2 >>
rect 182 152 183 153 
<< m1 >>
rect 190 152 191 153 
<< m2 >>
rect 198 152 199 153 
<< m1 >>
rect 199 152 200 153 
<< m1 >>
rect 226 152 227 153 
<< m2 >>
rect 226 152 227 153 
<< m2c >>
rect 226 152 227 153 
<< m1 >>
rect 226 152 227 153 
<< m2 >>
rect 226 152 227 153 
<< m1 >>
rect 247 152 248 153 
<< m1 >>
rect 248 152 249 153 
<< m2 >>
rect 248 152 249 153 
<< m2c >>
rect 248 152 249 153 
<< m1 >>
rect 248 152 249 153 
<< m2 >>
rect 248 152 249 153 
<< m2 >>
rect 249 152 250 153 
<< m1 >>
rect 250 152 251 153 
<< m2 >>
rect 250 152 251 153 
<< m2 >>
rect 251 152 252 153 
<< m1 >>
rect 252 152 253 153 
<< m2 >>
rect 252 152 253 153 
<< m2c >>
rect 252 152 253 153 
<< m1 >>
rect 252 152 253 153 
<< m2 >>
rect 252 152 253 153 
<< m1 >>
rect 253 152 254 153 
<< m2 >>
rect 254 152 255 153 
<< m1 >>
rect 256 152 257 153 
<< m1 >>
rect 13 153 14 154 
<< m1 >>
rect 14 153 15 154 
<< m1 >>
rect 15 153 16 154 
<< m1 >>
rect 16 153 17 154 
<< m1 >>
rect 17 153 18 154 
<< m1 >>
rect 18 153 19 154 
<< m1 >>
rect 19 153 20 154 
<< m2 >>
rect 19 153 20 154 
<< m1 >>
rect 20 153 21 154 
<< m1 >>
rect 21 153 22 154 
<< m1 >>
rect 22 153 23 154 
<< m1 >>
rect 23 153 24 154 
<< m1 >>
rect 24 153 25 154 
<< m1 >>
rect 25 153 26 154 
<< m1 >>
rect 26 153 27 154 
<< m1 >>
rect 28 153 29 154 
<< m1 >>
rect 32 153 33 154 
<< m1 >>
rect 34 153 35 154 
<< m1 >>
rect 35 153 36 154 
<< m1 >>
rect 36 153 37 154 
<< m1 >>
rect 37 153 38 154 
<< m1 >>
rect 44 153 45 154 
<< m1 >>
rect 46 153 47 154 
<< m1 >>
rect 52 153 53 154 
<< m1 >>
rect 55 153 56 154 
<< m1 >>
rect 57 153 58 154 
<< m1 >>
rect 64 153 65 154 
<< m2 >>
rect 64 153 65 154 
<< m1 >>
rect 67 153 68 154 
<< m1 >>
rect 68 153 69 154 
<< m1 >>
rect 69 153 70 154 
<< m1 >>
rect 70 153 71 154 
<< m1 >>
rect 71 153 72 154 
<< m2 >>
rect 71 153 72 154 
<< m2c >>
rect 71 153 72 154 
<< m1 >>
rect 71 153 72 154 
<< m2 >>
rect 71 153 72 154 
<< m2 >>
rect 72 153 73 154 
<< m1 >>
rect 73 153 74 154 
<< m2 >>
rect 73 153 74 154 
<< m1 >>
rect 82 153 83 154 
<< m1 >>
rect 88 153 89 154 
<< m2 >>
rect 89 153 90 154 
<< m1 >>
rect 91 153 92 154 
<< m1 >>
rect 95 153 96 154 
<< m1 >>
rect 121 153 122 154 
<< m1 >>
rect 145 153 146 154 
<< m1 >>
rect 163 153 164 154 
<< m1 >>
rect 165 153 166 154 
<< m1 >>
rect 181 153 182 154 
<< m2 >>
rect 182 153 183 154 
<< m1 >>
rect 190 153 191 154 
<< m2 >>
rect 198 153 199 154 
<< m1 >>
rect 199 153 200 154 
<< m2 >>
rect 226 153 227 154 
<< m1 >>
rect 247 153 248 154 
<< m1 >>
rect 250 153 251 154 
<< m2 >>
rect 254 153 255 154 
<< m1 >>
rect 256 153 257 154 
<< m1 >>
rect 13 154 14 155 
<< m2 >>
rect 19 154 20 155 
<< m1 >>
rect 26 154 27 155 
<< m1 >>
rect 28 154 29 155 
<< m1 >>
rect 32 154 33 155 
<< m2 >>
rect 32 154 33 155 
<< m2c >>
rect 32 154 33 155 
<< m1 >>
rect 32 154 33 155 
<< m2 >>
rect 32 154 33 155 
<< m2 >>
rect 33 154 34 155 
<< m2 >>
rect 34 154 35 155 
<< m1 >>
rect 37 154 38 155 
<< m1 >>
rect 44 154 45 155 
<< m1 >>
rect 46 154 47 155 
<< m1 >>
rect 52 154 53 155 
<< m1 >>
rect 55 154 56 155 
<< m1 >>
rect 57 154 58 155 
<< m1 >>
rect 64 154 65 155 
<< m2 >>
rect 64 154 65 155 
<< m1 >>
rect 67 154 68 155 
<< m1 >>
rect 73 154 74 155 
<< m2 >>
rect 73 154 74 155 
<< m1 >>
rect 82 154 83 155 
<< m1 >>
rect 88 154 89 155 
<< m2 >>
rect 89 154 90 155 
<< m2 >>
rect 90 154 91 155 
<< m1 >>
rect 91 154 92 155 
<< m2 >>
rect 91 154 92 155 
<< m2 >>
rect 92 154 93 155 
<< m1 >>
rect 95 154 96 155 
<< m1 >>
rect 106 154 107 155 
<< m1 >>
rect 107 154 108 155 
<< m1 >>
rect 108 154 109 155 
<< m1 >>
rect 109 154 110 155 
<< m1 >>
rect 121 154 122 155 
<< m1 >>
rect 145 154 146 155 
<< m1 >>
rect 160 154 161 155 
<< m1 >>
rect 161 154 162 155 
<< m2 >>
rect 161 154 162 155 
<< m2c >>
rect 161 154 162 155 
<< m1 >>
rect 161 154 162 155 
<< m2 >>
rect 161 154 162 155 
<< m2 >>
rect 162 154 163 155 
<< m1 >>
rect 163 154 164 155 
<< m2 >>
rect 163 154 164 155 
<< m2 >>
rect 164 154 165 155 
<< m1 >>
rect 165 154 166 155 
<< m2 >>
rect 165 154 166 155 
<< m2c >>
rect 165 154 166 155 
<< m1 >>
rect 165 154 166 155 
<< m2 >>
rect 165 154 166 155 
<< m1 >>
rect 181 154 182 155 
<< m2 >>
rect 182 154 183 155 
<< m1 >>
rect 190 154 191 155 
<< m1 >>
rect 196 154 197 155 
<< m1 >>
rect 197 154 198 155 
<< m2 >>
rect 197 154 198 155 
<< m2c >>
rect 197 154 198 155 
<< m1 >>
rect 197 154 198 155 
<< m2 >>
rect 197 154 198 155 
<< m2 >>
rect 198 154 199 155 
<< m1 >>
rect 199 154 200 155 
<< m1 >>
rect 226 154 227 155 
<< m2 >>
rect 226 154 227 155 
<< m1 >>
rect 227 154 228 155 
<< m1 >>
rect 228 154 229 155 
<< m1 >>
rect 229 154 230 155 
<< m1 >>
rect 247 154 248 155 
<< m1 >>
rect 250 154 251 155 
<< m1 >>
rect 254 154 255 155 
<< m2 >>
rect 254 154 255 155 
<< m2c >>
rect 254 154 255 155 
<< m1 >>
rect 254 154 255 155 
<< m2 >>
rect 254 154 255 155 
<< m1 >>
rect 256 154 257 155 
<< m1 >>
rect 13 155 14 156 
<< m1 >>
rect 19 155 20 156 
<< m2 >>
rect 19 155 20 156 
<< m2c >>
rect 19 155 20 156 
<< m1 >>
rect 19 155 20 156 
<< m2 >>
rect 19 155 20 156 
<< m1 >>
rect 26 155 27 156 
<< m1 >>
rect 28 155 29 156 
<< m1 >>
rect 34 155 35 156 
<< m2 >>
rect 34 155 35 156 
<< m1 >>
rect 37 155 38 156 
<< m1 >>
rect 44 155 45 156 
<< m1 >>
rect 46 155 47 156 
<< m1 >>
rect 52 155 53 156 
<< m1 >>
rect 55 155 56 156 
<< m1 >>
rect 57 155 58 156 
<< m1 >>
rect 64 155 65 156 
<< m2 >>
rect 64 155 65 156 
<< m1 >>
rect 67 155 68 156 
<< m1 >>
rect 73 155 74 156 
<< m2 >>
rect 73 155 74 156 
<< m1 >>
rect 82 155 83 156 
<< m1 >>
rect 88 155 89 156 
<< m1 >>
rect 91 155 92 156 
<< m2 >>
rect 92 155 93 156 
<< m1 >>
rect 95 155 96 156 
<< m1 >>
rect 106 155 107 156 
<< m1 >>
rect 109 155 110 156 
<< m1 >>
rect 121 155 122 156 
<< m1 >>
rect 145 155 146 156 
<< m1 >>
rect 160 155 161 156 
<< m1 >>
rect 163 155 164 156 
<< m1 >>
rect 181 155 182 156 
<< m2 >>
rect 182 155 183 156 
<< m1 >>
rect 190 155 191 156 
<< m1 >>
rect 196 155 197 156 
<< m1 >>
rect 199 155 200 156 
<< m1 >>
rect 226 155 227 156 
<< m2 >>
rect 226 155 227 156 
<< m1 >>
rect 229 155 230 156 
<< m1 >>
rect 247 155 248 156 
<< m1 >>
rect 250 155 251 156 
<< m1 >>
rect 254 155 255 156 
<< m1 >>
rect 256 155 257 156 
<< pdiffusion >>
rect 12 156 13 157 
<< m1 >>
rect 13 156 14 157 
<< pdiffusion >>
rect 13 156 14 157 
<< pdiffusion >>
rect 14 156 15 157 
<< pdiffusion >>
rect 15 156 16 157 
<< pdiffusion >>
rect 16 156 17 157 
<< pdiffusion >>
rect 17 156 18 157 
<< m1 >>
rect 19 156 20 157 
<< m1 >>
rect 26 156 27 157 
<< m1 >>
rect 28 156 29 157 
<< pdiffusion >>
rect 30 156 31 157 
<< pdiffusion >>
rect 31 156 32 157 
<< pdiffusion >>
rect 32 156 33 157 
<< m1 >>
rect 33 156 34 157 
<< m2 >>
rect 33 156 34 157 
<< m2c >>
rect 33 156 34 157 
<< m1 >>
rect 33 156 34 157 
<< m2 >>
rect 33 156 34 157 
<< pdiffusion >>
rect 33 156 34 157 
<< m1 >>
rect 34 156 35 157 
<< pdiffusion >>
rect 34 156 35 157 
<< pdiffusion >>
rect 35 156 36 157 
<< m1 >>
rect 37 156 38 157 
<< m1 >>
rect 44 156 45 157 
<< m1 >>
rect 46 156 47 157 
<< pdiffusion >>
rect 48 156 49 157 
<< pdiffusion >>
rect 49 156 50 157 
<< pdiffusion >>
rect 50 156 51 157 
<< pdiffusion >>
rect 51 156 52 157 
<< m1 >>
rect 52 156 53 157 
<< pdiffusion >>
rect 52 156 53 157 
<< pdiffusion >>
rect 53 156 54 157 
<< m1 >>
rect 55 156 56 157 
<< m1 >>
rect 57 156 58 157 
<< m1 >>
rect 64 156 65 157 
<< m2 >>
rect 64 156 65 157 
<< pdiffusion >>
rect 66 156 67 157 
<< m1 >>
rect 67 156 68 157 
<< pdiffusion >>
rect 67 156 68 157 
<< pdiffusion >>
rect 68 156 69 157 
<< pdiffusion >>
rect 69 156 70 157 
<< pdiffusion >>
rect 70 156 71 157 
<< pdiffusion >>
rect 71 156 72 157 
<< m1 >>
rect 73 156 74 157 
<< m2 >>
rect 73 156 74 157 
<< m1 >>
rect 82 156 83 157 
<< pdiffusion >>
rect 84 156 85 157 
<< pdiffusion >>
rect 85 156 86 157 
<< pdiffusion >>
rect 86 156 87 157 
<< pdiffusion >>
rect 87 156 88 157 
<< m1 >>
rect 88 156 89 157 
<< pdiffusion >>
rect 88 156 89 157 
<< pdiffusion >>
rect 89 156 90 157 
<< m1 >>
rect 91 156 92 157 
<< m2 >>
rect 92 156 93 157 
<< m1 >>
rect 95 156 96 157 
<< pdiffusion >>
rect 102 156 103 157 
<< m1 >>
rect 103 156 104 157 
<< pdiffusion >>
rect 103 156 104 157 
<< pdiffusion >>
rect 104 156 105 157 
<< pdiffusion >>
rect 105 156 106 157 
<< m1 >>
rect 106 156 107 157 
<< pdiffusion >>
rect 106 156 107 157 
<< pdiffusion >>
rect 107 156 108 157 
<< m1 >>
rect 109 156 110 157 
<< pdiffusion >>
rect 120 156 121 157 
<< m1 >>
rect 121 156 122 157 
<< pdiffusion >>
rect 121 156 122 157 
<< pdiffusion >>
rect 122 156 123 157 
<< pdiffusion >>
rect 123 156 124 157 
<< pdiffusion >>
rect 124 156 125 157 
<< pdiffusion >>
rect 125 156 126 157 
<< pdiffusion >>
rect 138 156 139 157 
<< pdiffusion >>
rect 139 156 140 157 
<< pdiffusion >>
rect 140 156 141 157 
<< pdiffusion >>
rect 141 156 142 157 
<< pdiffusion >>
rect 142 156 143 157 
<< pdiffusion >>
rect 143 156 144 157 
<< m1 >>
rect 145 156 146 157 
<< pdiffusion >>
rect 156 156 157 157 
<< pdiffusion >>
rect 157 156 158 157 
<< pdiffusion >>
rect 158 156 159 157 
<< pdiffusion >>
rect 159 156 160 157 
<< m1 >>
rect 160 156 161 157 
<< pdiffusion >>
rect 160 156 161 157 
<< pdiffusion >>
rect 161 156 162 157 
<< m1 >>
rect 163 156 164 157 
<< pdiffusion >>
rect 174 156 175 157 
<< pdiffusion >>
rect 175 156 176 157 
<< pdiffusion >>
rect 176 156 177 157 
<< pdiffusion >>
rect 177 156 178 157 
<< pdiffusion >>
rect 178 156 179 157 
<< pdiffusion >>
rect 179 156 180 157 
<< m1 >>
rect 181 156 182 157 
<< m2 >>
rect 182 156 183 157 
<< m1 >>
rect 190 156 191 157 
<< pdiffusion >>
rect 192 156 193 157 
<< pdiffusion >>
rect 193 156 194 157 
<< pdiffusion >>
rect 194 156 195 157 
<< pdiffusion >>
rect 195 156 196 157 
<< m1 >>
rect 196 156 197 157 
<< pdiffusion >>
rect 196 156 197 157 
<< pdiffusion >>
rect 197 156 198 157 
<< m1 >>
rect 199 156 200 157 
<< pdiffusion >>
rect 210 156 211 157 
<< pdiffusion >>
rect 211 156 212 157 
<< pdiffusion >>
rect 212 156 213 157 
<< pdiffusion >>
rect 213 156 214 157 
<< pdiffusion >>
rect 214 156 215 157 
<< pdiffusion >>
rect 215 156 216 157 
<< m1 >>
rect 226 156 227 157 
<< m2 >>
rect 226 156 227 157 
<< pdiffusion >>
rect 228 156 229 157 
<< m1 >>
rect 229 156 230 157 
<< pdiffusion >>
rect 229 156 230 157 
<< pdiffusion >>
rect 230 156 231 157 
<< pdiffusion >>
rect 231 156 232 157 
<< pdiffusion >>
rect 232 156 233 157 
<< pdiffusion >>
rect 233 156 234 157 
<< pdiffusion >>
rect 246 156 247 157 
<< m1 >>
rect 247 156 248 157 
<< pdiffusion >>
rect 247 156 248 157 
<< pdiffusion >>
rect 248 156 249 157 
<< pdiffusion >>
rect 249 156 250 157 
<< m1 >>
rect 250 156 251 157 
<< pdiffusion >>
rect 250 156 251 157 
<< pdiffusion >>
rect 251 156 252 157 
<< m1 >>
rect 254 156 255 157 
<< m1 >>
rect 256 156 257 157 
<< pdiffusion >>
rect 12 157 13 158 
<< pdiffusion >>
rect 13 157 14 158 
<< pdiffusion >>
rect 14 157 15 158 
<< pdiffusion >>
rect 15 157 16 158 
<< pdiffusion >>
rect 16 157 17 158 
<< pdiffusion >>
rect 17 157 18 158 
<< m1 >>
rect 19 157 20 158 
<< m1 >>
rect 26 157 27 158 
<< m1 >>
rect 28 157 29 158 
<< pdiffusion >>
rect 30 157 31 158 
<< pdiffusion >>
rect 31 157 32 158 
<< pdiffusion >>
rect 32 157 33 158 
<< pdiffusion >>
rect 33 157 34 158 
<< pdiffusion >>
rect 34 157 35 158 
<< pdiffusion >>
rect 35 157 36 158 
<< m1 >>
rect 37 157 38 158 
<< m1 >>
rect 44 157 45 158 
<< m1 >>
rect 46 157 47 158 
<< pdiffusion >>
rect 48 157 49 158 
<< pdiffusion >>
rect 49 157 50 158 
<< pdiffusion >>
rect 50 157 51 158 
<< pdiffusion >>
rect 51 157 52 158 
<< pdiffusion >>
rect 52 157 53 158 
<< pdiffusion >>
rect 53 157 54 158 
<< m1 >>
rect 55 157 56 158 
<< m1 >>
rect 57 157 58 158 
<< m1 >>
rect 64 157 65 158 
<< m2 >>
rect 64 157 65 158 
<< pdiffusion >>
rect 66 157 67 158 
<< pdiffusion >>
rect 67 157 68 158 
<< pdiffusion >>
rect 68 157 69 158 
<< pdiffusion >>
rect 69 157 70 158 
<< pdiffusion >>
rect 70 157 71 158 
<< pdiffusion >>
rect 71 157 72 158 
<< m1 >>
rect 73 157 74 158 
<< m2 >>
rect 73 157 74 158 
<< m1 >>
rect 82 157 83 158 
<< pdiffusion >>
rect 84 157 85 158 
<< pdiffusion >>
rect 85 157 86 158 
<< pdiffusion >>
rect 86 157 87 158 
<< pdiffusion >>
rect 87 157 88 158 
<< pdiffusion >>
rect 88 157 89 158 
<< pdiffusion >>
rect 89 157 90 158 
<< m1 >>
rect 91 157 92 158 
<< m2 >>
rect 92 157 93 158 
<< m1 >>
rect 95 157 96 158 
<< pdiffusion >>
rect 102 157 103 158 
<< pdiffusion >>
rect 103 157 104 158 
<< pdiffusion >>
rect 104 157 105 158 
<< pdiffusion >>
rect 105 157 106 158 
<< pdiffusion >>
rect 106 157 107 158 
<< pdiffusion >>
rect 107 157 108 158 
<< m1 >>
rect 109 157 110 158 
<< pdiffusion >>
rect 120 157 121 158 
<< pdiffusion >>
rect 121 157 122 158 
<< pdiffusion >>
rect 122 157 123 158 
<< pdiffusion >>
rect 123 157 124 158 
<< pdiffusion >>
rect 124 157 125 158 
<< pdiffusion >>
rect 125 157 126 158 
<< pdiffusion >>
rect 138 157 139 158 
<< pdiffusion >>
rect 139 157 140 158 
<< pdiffusion >>
rect 140 157 141 158 
<< pdiffusion >>
rect 141 157 142 158 
<< pdiffusion >>
rect 142 157 143 158 
<< pdiffusion >>
rect 143 157 144 158 
<< m1 >>
rect 145 157 146 158 
<< pdiffusion >>
rect 156 157 157 158 
<< pdiffusion >>
rect 157 157 158 158 
<< pdiffusion >>
rect 158 157 159 158 
<< pdiffusion >>
rect 159 157 160 158 
<< pdiffusion >>
rect 160 157 161 158 
<< pdiffusion >>
rect 161 157 162 158 
<< m1 >>
rect 163 157 164 158 
<< pdiffusion >>
rect 174 157 175 158 
<< pdiffusion >>
rect 175 157 176 158 
<< pdiffusion >>
rect 176 157 177 158 
<< pdiffusion >>
rect 177 157 178 158 
<< pdiffusion >>
rect 178 157 179 158 
<< pdiffusion >>
rect 179 157 180 158 
<< m1 >>
rect 181 157 182 158 
<< m2 >>
rect 182 157 183 158 
<< m1 >>
rect 190 157 191 158 
<< pdiffusion >>
rect 192 157 193 158 
<< pdiffusion >>
rect 193 157 194 158 
<< pdiffusion >>
rect 194 157 195 158 
<< pdiffusion >>
rect 195 157 196 158 
<< pdiffusion >>
rect 196 157 197 158 
<< pdiffusion >>
rect 197 157 198 158 
<< m1 >>
rect 199 157 200 158 
<< pdiffusion >>
rect 210 157 211 158 
<< pdiffusion >>
rect 211 157 212 158 
<< pdiffusion >>
rect 212 157 213 158 
<< pdiffusion >>
rect 213 157 214 158 
<< pdiffusion >>
rect 214 157 215 158 
<< pdiffusion >>
rect 215 157 216 158 
<< m1 >>
rect 226 157 227 158 
<< m2 >>
rect 226 157 227 158 
<< pdiffusion >>
rect 228 157 229 158 
<< pdiffusion >>
rect 229 157 230 158 
<< pdiffusion >>
rect 230 157 231 158 
<< pdiffusion >>
rect 231 157 232 158 
<< pdiffusion >>
rect 232 157 233 158 
<< pdiffusion >>
rect 233 157 234 158 
<< pdiffusion >>
rect 246 157 247 158 
<< pdiffusion >>
rect 247 157 248 158 
<< pdiffusion >>
rect 248 157 249 158 
<< pdiffusion >>
rect 249 157 250 158 
<< pdiffusion >>
rect 250 157 251 158 
<< pdiffusion >>
rect 251 157 252 158 
<< m1 >>
rect 254 157 255 158 
<< m1 >>
rect 256 157 257 158 
<< pdiffusion >>
rect 12 158 13 159 
<< pdiffusion >>
rect 13 158 14 159 
<< pdiffusion >>
rect 14 158 15 159 
<< pdiffusion >>
rect 15 158 16 159 
<< pdiffusion >>
rect 16 158 17 159 
<< pdiffusion >>
rect 17 158 18 159 
<< m1 >>
rect 19 158 20 159 
<< m1 >>
rect 26 158 27 159 
<< m1 >>
rect 28 158 29 159 
<< pdiffusion >>
rect 30 158 31 159 
<< pdiffusion >>
rect 31 158 32 159 
<< pdiffusion >>
rect 32 158 33 159 
<< pdiffusion >>
rect 33 158 34 159 
<< pdiffusion >>
rect 34 158 35 159 
<< pdiffusion >>
rect 35 158 36 159 
<< m1 >>
rect 37 158 38 159 
<< m1 >>
rect 44 158 45 159 
<< m1 >>
rect 46 158 47 159 
<< pdiffusion >>
rect 48 158 49 159 
<< pdiffusion >>
rect 49 158 50 159 
<< pdiffusion >>
rect 50 158 51 159 
<< pdiffusion >>
rect 51 158 52 159 
<< pdiffusion >>
rect 52 158 53 159 
<< pdiffusion >>
rect 53 158 54 159 
<< m1 >>
rect 55 158 56 159 
<< m1 >>
rect 57 158 58 159 
<< m1 >>
rect 64 158 65 159 
<< m2 >>
rect 64 158 65 159 
<< pdiffusion >>
rect 66 158 67 159 
<< pdiffusion >>
rect 67 158 68 159 
<< pdiffusion >>
rect 68 158 69 159 
<< pdiffusion >>
rect 69 158 70 159 
<< pdiffusion >>
rect 70 158 71 159 
<< pdiffusion >>
rect 71 158 72 159 
<< m1 >>
rect 73 158 74 159 
<< m2 >>
rect 73 158 74 159 
<< m1 >>
rect 82 158 83 159 
<< pdiffusion >>
rect 84 158 85 159 
<< pdiffusion >>
rect 85 158 86 159 
<< pdiffusion >>
rect 86 158 87 159 
<< pdiffusion >>
rect 87 158 88 159 
<< pdiffusion >>
rect 88 158 89 159 
<< pdiffusion >>
rect 89 158 90 159 
<< m1 >>
rect 91 158 92 159 
<< m2 >>
rect 92 158 93 159 
<< m1 >>
rect 95 158 96 159 
<< pdiffusion >>
rect 102 158 103 159 
<< pdiffusion >>
rect 103 158 104 159 
<< pdiffusion >>
rect 104 158 105 159 
<< pdiffusion >>
rect 105 158 106 159 
<< pdiffusion >>
rect 106 158 107 159 
<< pdiffusion >>
rect 107 158 108 159 
<< m1 >>
rect 109 158 110 159 
<< pdiffusion >>
rect 120 158 121 159 
<< pdiffusion >>
rect 121 158 122 159 
<< pdiffusion >>
rect 122 158 123 159 
<< pdiffusion >>
rect 123 158 124 159 
<< pdiffusion >>
rect 124 158 125 159 
<< pdiffusion >>
rect 125 158 126 159 
<< pdiffusion >>
rect 138 158 139 159 
<< pdiffusion >>
rect 139 158 140 159 
<< pdiffusion >>
rect 140 158 141 159 
<< pdiffusion >>
rect 141 158 142 159 
<< pdiffusion >>
rect 142 158 143 159 
<< pdiffusion >>
rect 143 158 144 159 
<< m1 >>
rect 145 158 146 159 
<< pdiffusion >>
rect 156 158 157 159 
<< pdiffusion >>
rect 157 158 158 159 
<< pdiffusion >>
rect 158 158 159 159 
<< pdiffusion >>
rect 159 158 160 159 
<< pdiffusion >>
rect 160 158 161 159 
<< pdiffusion >>
rect 161 158 162 159 
<< m1 >>
rect 163 158 164 159 
<< pdiffusion >>
rect 174 158 175 159 
<< pdiffusion >>
rect 175 158 176 159 
<< pdiffusion >>
rect 176 158 177 159 
<< pdiffusion >>
rect 177 158 178 159 
<< pdiffusion >>
rect 178 158 179 159 
<< pdiffusion >>
rect 179 158 180 159 
<< m1 >>
rect 181 158 182 159 
<< m2 >>
rect 182 158 183 159 
<< m1 >>
rect 190 158 191 159 
<< pdiffusion >>
rect 192 158 193 159 
<< pdiffusion >>
rect 193 158 194 159 
<< pdiffusion >>
rect 194 158 195 159 
<< pdiffusion >>
rect 195 158 196 159 
<< pdiffusion >>
rect 196 158 197 159 
<< pdiffusion >>
rect 197 158 198 159 
<< m1 >>
rect 199 158 200 159 
<< pdiffusion >>
rect 210 158 211 159 
<< pdiffusion >>
rect 211 158 212 159 
<< pdiffusion >>
rect 212 158 213 159 
<< pdiffusion >>
rect 213 158 214 159 
<< pdiffusion >>
rect 214 158 215 159 
<< pdiffusion >>
rect 215 158 216 159 
<< m1 >>
rect 226 158 227 159 
<< m2 >>
rect 226 158 227 159 
<< pdiffusion >>
rect 228 158 229 159 
<< pdiffusion >>
rect 229 158 230 159 
<< pdiffusion >>
rect 230 158 231 159 
<< pdiffusion >>
rect 231 158 232 159 
<< pdiffusion >>
rect 232 158 233 159 
<< pdiffusion >>
rect 233 158 234 159 
<< pdiffusion >>
rect 246 158 247 159 
<< pdiffusion >>
rect 247 158 248 159 
<< pdiffusion >>
rect 248 158 249 159 
<< pdiffusion >>
rect 249 158 250 159 
<< pdiffusion >>
rect 250 158 251 159 
<< pdiffusion >>
rect 251 158 252 159 
<< m1 >>
rect 254 158 255 159 
<< m1 >>
rect 256 158 257 159 
<< pdiffusion >>
rect 12 159 13 160 
<< pdiffusion >>
rect 13 159 14 160 
<< pdiffusion >>
rect 14 159 15 160 
<< pdiffusion >>
rect 15 159 16 160 
<< pdiffusion >>
rect 16 159 17 160 
<< pdiffusion >>
rect 17 159 18 160 
<< m1 >>
rect 19 159 20 160 
<< m1 >>
rect 26 159 27 160 
<< m1 >>
rect 28 159 29 160 
<< pdiffusion >>
rect 30 159 31 160 
<< pdiffusion >>
rect 31 159 32 160 
<< pdiffusion >>
rect 32 159 33 160 
<< pdiffusion >>
rect 33 159 34 160 
<< pdiffusion >>
rect 34 159 35 160 
<< pdiffusion >>
rect 35 159 36 160 
<< m1 >>
rect 37 159 38 160 
<< m1 >>
rect 44 159 45 160 
<< m1 >>
rect 46 159 47 160 
<< pdiffusion >>
rect 48 159 49 160 
<< pdiffusion >>
rect 49 159 50 160 
<< pdiffusion >>
rect 50 159 51 160 
<< pdiffusion >>
rect 51 159 52 160 
<< pdiffusion >>
rect 52 159 53 160 
<< pdiffusion >>
rect 53 159 54 160 
<< m1 >>
rect 55 159 56 160 
<< m1 >>
rect 57 159 58 160 
<< m1 >>
rect 64 159 65 160 
<< m2 >>
rect 64 159 65 160 
<< pdiffusion >>
rect 66 159 67 160 
<< pdiffusion >>
rect 67 159 68 160 
<< pdiffusion >>
rect 68 159 69 160 
<< pdiffusion >>
rect 69 159 70 160 
<< pdiffusion >>
rect 70 159 71 160 
<< pdiffusion >>
rect 71 159 72 160 
<< m1 >>
rect 73 159 74 160 
<< m2 >>
rect 73 159 74 160 
<< m1 >>
rect 82 159 83 160 
<< pdiffusion >>
rect 84 159 85 160 
<< pdiffusion >>
rect 85 159 86 160 
<< pdiffusion >>
rect 86 159 87 160 
<< pdiffusion >>
rect 87 159 88 160 
<< pdiffusion >>
rect 88 159 89 160 
<< pdiffusion >>
rect 89 159 90 160 
<< m1 >>
rect 91 159 92 160 
<< m2 >>
rect 92 159 93 160 
<< m1 >>
rect 95 159 96 160 
<< pdiffusion >>
rect 102 159 103 160 
<< pdiffusion >>
rect 103 159 104 160 
<< pdiffusion >>
rect 104 159 105 160 
<< pdiffusion >>
rect 105 159 106 160 
<< pdiffusion >>
rect 106 159 107 160 
<< pdiffusion >>
rect 107 159 108 160 
<< m1 >>
rect 109 159 110 160 
<< pdiffusion >>
rect 120 159 121 160 
<< pdiffusion >>
rect 121 159 122 160 
<< pdiffusion >>
rect 122 159 123 160 
<< pdiffusion >>
rect 123 159 124 160 
<< pdiffusion >>
rect 124 159 125 160 
<< pdiffusion >>
rect 125 159 126 160 
<< pdiffusion >>
rect 138 159 139 160 
<< pdiffusion >>
rect 139 159 140 160 
<< pdiffusion >>
rect 140 159 141 160 
<< pdiffusion >>
rect 141 159 142 160 
<< pdiffusion >>
rect 142 159 143 160 
<< pdiffusion >>
rect 143 159 144 160 
<< m1 >>
rect 145 159 146 160 
<< pdiffusion >>
rect 156 159 157 160 
<< pdiffusion >>
rect 157 159 158 160 
<< pdiffusion >>
rect 158 159 159 160 
<< pdiffusion >>
rect 159 159 160 160 
<< pdiffusion >>
rect 160 159 161 160 
<< pdiffusion >>
rect 161 159 162 160 
<< m1 >>
rect 163 159 164 160 
<< pdiffusion >>
rect 174 159 175 160 
<< pdiffusion >>
rect 175 159 176 160 
<< pdiffusion >>
rect 176 159 177 160 
<< pdiffusion >>
rect 177 159 178 160 
<< pdiffusion >>
rect 178 159 179 160 
<< pdiffusion >>
rect 179 159 180 160 
<< m1 >>
rect 181 159 182 160 
<< m2 >>
rect 182 159 183 160 
<< m1 >>
rect 190 159 191 160 
<< pdiffusion >>
rect 192 159 193 160 
<< pdiffusion >>
rect 193 159 194 160 
<< pdiffusion >>
rect 194 159 195 160 
<< pdiffusion >>
rect 195 159 196 160 
<< pdiffusion >>
rect 196 159 197 160 
<< pdiffusion >>
rect 197 159 198 160 
<< m1 >>
rect 199 159 200 160 
<< pdiffusion >>
rect 210 159 211 160 
<< pdiffusion >>
rect 211 159 212 160 
<< pdiffusion >>
rect 212 159 213 160 
<< pdiffusion >>
rect 213 159 214 160 
<< pdiffusion >>
rect 214 159 215 160 
<< pdiffusion >>
rect 215 159 216 160 
<< m1 >>
rect 226 159 227 160 
<< m2 >>
rect 226 159 227 160 
<< pdiffusion >>
rect 228 159 229 160 
<< pdiffusion >>
rect 229 159 230 160 
<< pdiffusion >>
rect 230 159 231 160 
<< pdiffusion >>
rect 231 159 232 160 
<< pdiffusion >>
rect 232 159 233 160 
<< pdiffusion >>
rect 233 159 234 160 
<< pdiffusion >>
rect 246 159 247 160 
<< pdiffusion >>
rect 247 159 248 160 
<< pdiffusion >>
rect 248 159 249 160 
<< pdiffusion >>
rect 249 159 250 160 
<< pdiffusion >>
rect 250 159 251 160 
<< pdiffusion >>
rect 251 159 252 160 
<< m1 >>
rect 254 159 255 160 
<< m1 >>
rect 256 159 257 160 
<< pdiffusion >>
rect 12 160 13 161 
<< pdiffusion >>
rect 13 160 14 161 
<< pdiffusion >>
rect 14 160 15 161 
<< pdiffusion >>
rect 15 160 16 161 
<< pdiffusion >>
rect 16 160 17 161 
<< pdiffusion >>
rect 17 160 18 161 
<< m1 >>
rect 19 160 20 161 
<< m1 >>
rect 26 160 27 161 
<< m1 >>
rect 28 160 29 161 
<< pdiffusion >>
rect 30 160 31 161 
<< pdiffusion >>
rect 31 160 32 161 
<< pdiffusion >>
rect 32 160 33 161 
<< pdiffusion >>
rect 33 160 34 161 
<< pdiffusion >>
rect 34 160 35 161 
<< pdiffusion >>
rect 35 160 36 161 
<< m1 >>
rect 37 160 38 161 
<< m1 >>
rect 44 160 45 161 
<< m1 >>
rect 46 160 47 161 
<< pdiffusion >>
rect 48 160 49 161 
<< pdiffusion >>
rect 49 160 50 161 
<< pdiffusion >>
rect 50 160 51 161 
<< pdiffusion >>
rect 51 160 52 161 
<< pdiffusion >>
rect 52 160 53 161 
<< pdiffusion >>
rect 53 160 54 161 
<< m1 >>
rect 55 160 56 161 
<< m1 >>
rect 57 160 58 161 
<< m1 >>
rect 64 160 65 161 
<< m2 >>
rect 64 160 65 161 
<< pdiffusion >>
rect 66 160 67 161 
<< pdiffusion >>
rect 67 160 68 161 
<< pdiffusion >>
rect 68 160 69 161 
<< pdiffusion >>
rect 69 160 70 161 
<< pdiffusion >>
rect 70 160 71 161 
<< pdiffusion >>
rect 71 160 72 161 
<< m1 >>
rect 73 160 74 161 
<< m2 >>
rect 73 160 74 161 
<< m1 >>
rect 82 160 83 161 
<< pdiffusion >>
rect 84 160 85 161 
<< pdiffusion >>
rect 85 160 86 161 
<< pdiffusion >>
rect 86 160 87 161 
<< pdiffusion >>
rect 87 160 88 161 
<< pdiffusion >>
rect 88 160 89 161 
<< pdiffusion >>
rect 89 160 90 161 
<< m1 >>
rect 91 160 92 161 
<< m2 >>
rect 92 160 93 161 
<< m1 >>
rect 95 160 96 161 
<< pdiffusion >>
rect 102 160 103 161 
<< pdiffusion >>
rect 103 160 104 161 
<< pdiffusion >>
rect 104 160 105 161 
<< pdiffusion >>
rect 105 160 106 161 
<< pdiffusion >>
rect 106 160 107 161 
<< pdiffusion >>
rect 107 160 108 161 
<< m1 >>
rect 109 160 110 161 
<< pdiffusion >>
rect 120 160 121 161 
<< pdiffusion >>
rect 121 160 122 161 
<< pdiffusion >>
rect 122 160 123 161 
<< pdiffusion >>
rect 123 160 124 161 
<< pdiffusion >>
rect 124 160 125 161 
<< pdiffusion >>
rect 125 160 126 161 
<< pdiffusion >>
rect 138 160 139 161 
<< pdiffusion >>
rect 139 160 140 161 
<< pdiffusion >>
rect 140 160 141 161 
<< pdiffusion >>
rect 141 160 142 161 
<< pdiffusion >>
rect 142 160 143 161 
<< pdiffusion >>
rect 143 160 144 161 
<< m1 >>
rect 145 160 146 161 
<< pdiffusion >>
rect 156 160 157 161 
<< pdiffusion >>
rect 157 160 158 161 
<< pdiffusion >>
rect 158 160 159 161 
<< pdiffusion >>
rect 159 160 160 161 
<< pdiffusion >>
rect 160 160 161 161 
<< pdiffusion >>
rect 161 160 162 161 
<< m1 >>
rect 163 160 164 161 
<< pdiffusion >>
rect 174 160 175 161 
<< pdiffusion >>
rect 175 160 176 161 
<< pdiffusion >>
rect 176 160 177 161 
<< pdiffusion >>
rect 177 160 178 161 
<< pdiffusion >>
rect 178 160 179 161 
<< pdiffusion >>
rect 179 160 180 161 
<< m1 >>
rect 181 160 182 161 
<< m2 >>
rect 182 160 183 161 
<< m1 >>
rect 183 160 184 161 
<< m2 >>
rect 183 160 184 161 
<< m2c >>
rect 183 160 184 161 
<< m1 >>
rect 183 160 184 161 
<< m2 >>
rect 183 160 184 161 
<< m1 >>
rect 184 160 185 161 
<< m1 >>
rect 185 160 186 161 
<< m1 >>
rect 186 160 187 161 
<< m1 >>
rect 187 160 188 161 
<< m1 >>
rect 188 160 189 161 
<< m1 >>
rect 190 160 191 161 
<< pdiffusion >>
rect 192 160 193 161 
<< pdiffusion >>
rect 193 160 194 161 
<< pdiffusion >>
rect 194 160 195 161 
<< pdiffusion >>
rect 195 160 196 161 
<< pdiffusion >>
rect 196 160 197 161 
<< pdiffusion >>
rect 197 160 198 161 
<< m1 >>
rect 199 160 200 161 
<< pdiffusion >>
rect 210 160 211 161 
<< pdiffusion >>
rect 211 160 212 161 
<< pdiffusion >>
rect 212 160 213 161 
<< pdiffusion >>
rect 213 160 214 161 
<< pdiffusion >>
rect 214 160 215 161 
<< pdiffusion >>
rect 215 160 216 161 
<< m1 >>
rect 226 160 227 161 
<< m2 >>
rect 226 160 227 161 
<< pdiffusion >>
rect 228 160 229 161 
<< pdiffusion >>
rect 229 160 230 161 
<< pdiffusion >>
rect 230 160 231 161 
<< pdiffusion >>
rect 231 160 232 161 
<< pdiffusion >>
rect 232 160 233 161 
<< pdiffusion >>
rect 233 160 234 161 
<< pdiffusion >>
rect 246 160 247 161 
<< pdiffusion >>
rect 247 160 248 161 
<< pdiffusion >>
rect 248 160 249 161 
<< pdiffusion >>
rect 249 160 250 161 
<< pdiffusion >>
rect 250 160 251 161 
<< pdiffusion >>
rect 251 160 252 161 
<< m1 >>
rect 254 160 255 161 
<< m1 >>
rect 256 160 257 161 
<< pdiffusion >>
rect 12 161 13 162 
<< pdiffusion >>
rect 13 161 14 162 
<< pdiffusion >>
rect 14 161 15 162 
<< pdiffusion >>
rect 15 161 16 162 
<< pdiffusion >>
rect 16 161 17 162 
<< pdiffusion >>
rect 17 161 18 162 
<< m1 >>
rect 19 161 20 162 
<< m1 >>
rect 26 161 27 162 
<< m1 >>
rect 28 161 29 162 
<< pdiffusion >>
rect 30 161 31 162 
<< pdiffusion >>
rect 31 161 32 162 
<< pdiffusion >>
rect 32 161 33 162 
<< pdiffusion >>
rect 33 161 34 162 
<< m1 >>
rect 34 161 35 162 
<< pdiffusion >>
rect 34 161 35 162 
<< pdiffusion >>
rect 35 161 36 162 
<< m1 >>
rect 37 161 38 162 
<< m1 >>
rect 44 161 45 162 
<< m1 >>
rect 46 161 47 162 
<< pdiffusion >>
rect 48 161 49 162 
<< m1 >>
rect 49 161 50 162 
<< pdiffusion >>
rect 49 161 50 162 
<< pdiffusion >>
rect 50 161 51 162 
<< m1 >>
rect 51 161 52 162 
<< m2 >>
rect 51 161 52 162 
<< m2c >>
rect 51 161 52 162 
<< m1 >>
rect 51 161 52 162 
<< m2 >>
rect 51 161 52 162 
<< pdiffusion >>
rect 51 161 52 162 
<< m1 >>
rect 52 161 53 162 
<< pdiffusion >>
rect 52 161 53 162 
<< pdiffusion >>
rect 53 161 54 162 
<< m1 >>
rect 55 161 56 162 
<< m1 >>
rect 57 161 58 162 
<< m1 >>
rect 64 161 65 162 
<< m2 >>
rect 64 161 65 162 
<< pdiffusion >>
rect 66 161 67 162 
<< pdiffusion >>
rect 67 161 68 162 
<< pdiffusion >>
rect 68 161 69 162 
<< pdiffusion >>
rect 69 161 70 162 
<< m1 >>
rect 70 161 71 162 
<< pdiffusion >>
rect 70 161 71 162 
<< pdiffusion >>
rect 71 161 72 162 
<< m1 >>
rect 73 161 74 162 
<< m2 >>
rect 73 161 74 162 
<< m1 >>
rect 82 161 83 162 
<< pdiffusion >>
rect 84 161 85 162 
<< pdiffusion >>
rect 85 161 86 162 
<< pdiffusion >>
rect 86 161 87 162 
<< pdiffusion >>
rect 87 161 88 162 
<< pdiffusion >>
rect 88 161 89 162 
<< pdiffusion >>
rect 89 161 90 162 
<< m1 >>
rect 91 161 92 162 
<< m2 >>
rect 92 161 93 162 
<< m1 >>
rect 95 161 96 162 
<< pdiffusion >>
rect 102 161 103 162 
<< m1 >>
rect 103 161 104 162 
<< pdiffusion >>
rect 103 161 104 162 
<< pdiffusion >>
rect 104 161 105 162 
<< pdiffusion >>
rect 105 161 106 162 
<< pdiffusion >>
rect 106 161 107 162 
<< pdiffusion >>
rect 107 161 108 162 
<< m1 >>
rect 109 161 110 162 
<< pdiffusion >>
rect 120 161 121 162 
<< pdiffusion >>
rect 121 161 122 162 
<< pdiffusion >>
rect 122 161 123 162 
<< pdiffusion >>
rect 123 161 124 162 
<< m1 >>
rect 124 161 125 162 
<< pdiffusion >>
rect 124 161 125 162 
<< pdiffusion >>
rect 125 161 126 162 
<< pdiffusion >>
rect 138 161 139 162 
<< m1 >>
rect 139 161 140 162 
<< pdiffusion >>
rect 139 161 140 162 
<< pdiffusion >>
rect 140 161 141 162 
<< pdiffusion >>
rect 141 161 142 162 
<< m1 >>
rect 142 161 143 162 
<< pdiffusion >>
rect 142 161 143 162 
<< pdiffusion >>
rect 143 161 144 162 
<< m1 >>
rect 145 161 146 162 
<< pdiffusion >>
rect 156 161 157 162 
<< m1 >>
rect 157 161 158 162 
<< pdiffusion >>
rect 157 161 158 162 
<< pdiffusion >>
rect 158 161 159 162 
<< pdiffusion >>
rect 159 161 160 162 
<< pdiffusion >>
rect 160 161 161 162 
<< pdiffusion >>
rect 161 161 162 162 
<< m1 >>
rect 163 161 164 162 
<< pdiffusion >>
rect 174 161 175 162 
<< m1 >>
rect 175 161 176 162 
<< pdiffusion >>
rect 175 161 176 162 
<< pdiffusion >>
rect 176 161 177 162 
<< pdiffusion >>
rect 177 161 178 162 
<< pdiffusion >>
rect 178 161 179 162 
<< pdiffusion >>
rect 179 161 180 162 
<< m1 >>
rect 181 161 182 162 
<< m1 >>
rect 188 161 189 162 
<< m1 >>
rect 190 161 191 162 
<< pdiffusion >>
rect 192 161 193 162 
<< m1 >>
rect 193 161 194 162 
<< pdiffusion >>
rect 193 161 194 162 
<< pdiffusion >>
rect 194 161 195 162 
<< pdiffusion >>
rect 195 161 196 162 
<< pdiffusion >>
rect 196 161 197 162 
<< pdiffusion >>
rect 197 161 198 162 
<< m1 >>
rect 199 161 200 162 
<< pdiffusion >>
rect 210 161 211 162 
<< pdiffusion >>
rect 211 161 212 162 
<< pdiffusion >>
rect 212 161 213 162 
<< pdiffusion >>
rect 213 161 214 162 
<< pdiffusion >>
rect 214 161 215 162 
<< pdiffusion >>
rect 215 161 216 162 
<< m1 >>
rect 226 161 227 162 
<< m2 >>
rect 226 161 227 162 
<< pdiffusion >>
rect 228 161 229 162 
<< m1 >>
rect 229 161 230 162 
<< pdiffusion >>
rect 229 161 230 162 
<< pdiffusion >>
rect 230 161 231 162 
<< pdiffusion >>
rect 231 161 232 162 
<< pdiffusion >>
rect 232 161 233 162 
<< pdiffusion >>
rect 233 161 234 162 
<< pdiffusion >>
rect 246 161 247 162 
<< pdiffusion >>
rect 247 161 248 162 
<< pdiffusion >>
rect 248 161 249 162 
<< pdiffusion >>
rect 249 161 250 162 
<< pdiffusion >>
rect 250 161 251 162 
<< pdiffusion >>
rect 251 161 252 162 
<< m1 >>
rect 254 161 255 162 
<< m1 >>
rect 256 161 257 162 
<< m1 >>
rect 19 162 20 163 
<< m1 >>
rect 26 162 27 163 
<< m1 >>
rect 28 162 29 163 
<< m1 >>
rect 34 162 35 163 
<< m1 >>
rect 37 162 38 163 
<< m1 >>
rect 44 162 45 163 
<< m1 >>
rect 46 162 47 163 
<< m1 >>
rect 49 162 50 163 
<< m1 >>
rect 52 162 53 163 
<< m2 >>
rect 52 162 53 163 
<< m1 >>
rect 55 162 56 163 
<< m2 >>
rect 55 162 56 163 
<< m2c >>
rect 55 162 56 163 
<< m1 >>
rect 55 162 56 163 
<< m2 >>
rect 55 162 56 163 
<< m1 >>
rect 57 162 58 163 
<< m2 >>
rect 57 162 58 163 
<< m2c >>
rect 57 162 58 163 
<< m1 >>
rect 57 162 58 163 
<< m2 >>
rect 57 162 58 163 
<< m1 >>
rect 64 162 65 163 
<< m2 >>
rect 64 162 65 163 
<< m1 >>
rect 70 162 71 163 
<< m1 >>
rect 73 162 74 163 
<< m2 >>
rect 73 162 74 163 
<< m1 >>
rect 82 162 83 163 
<< m1 >>
rect 91 162 92 163 
<< m2 >>
rect 92 162 93 163 
<< m1 >>
rect 95 162 96 163 
<< m1 >>
rect 103 162 104 163 
<< m1 >>
rect 109 162 110 163 
<< m1 >>
rect 124 162 125 163 
<< m1 >>
rect 139 162 140 163 
<< m1 >>
rect 142 162 143 163 
<< m1 >>
rect 145 162 146 163 
<< m1 >>
rect 157 162 158 163 
<< m1 >>
rect 163 162 164 163 
<< m1 >>
rect 175 162 176 163 
<< m1 >>
rect 181 162 182 163 
<< m2 >>
rect 181 162 182 163 
<< m2c >>
rect 181 162 182 163 
<< m1 >>
rect 181 162 182 163 
<< m2 >>
rect 181 162 182 163 
<< m1 >>
rect 188 162 189 163 
<< m2 >>
rect 188 162 189 163 
<< m2c >>
rect 188 162 189 163 
<< m1 >>
rect 188 162 189 163 
<< m2 >>
rect 188 162 189 163 
<< m2 >>
rect 189 162 190 163 
<< m1 >>
rect 190 162 191 163 
<< m2 >>
rect 190 162 191 163 
<< m1 >>
rect 193 162 194 163 
<< m1 >>
rect 199 162 200 163 
<< m1 >>
rect 226 162 227 163 
<< m2 >>
rect 226 162 227 163 
<< m1 >>
rect 229 162 230 163 
<< m1 >>
rect 254 162 255 163 
<< m1 >>
rect 256 162 257 163 
<< m1 >>
rect 19 163 20 164 
<< m1 >>
rect 26 163 27 164 
<< m1 >>
rect 28 163 29 164 
<< m1 >>
rect 34 163 35 164 
<< m1 >>
rect 35 163 36 164 
<< m1 >>
rect 36 163 37 164 
<< m1 >>
rect 37 163 38 164 
<< m1 >>
rect 44 163 45 164 
<< m1 >>
rect 46 163 47 164 
<< m1 >>
rect 49 163 50 164 
<< m2 >>
rect 52 163 53 164 
<< m2 >>
rect 55 163 56 164 
<< m2 >>
rect 57 163 58 164 
<< m1 >>
rect 64 163 65 164 
<< m2 >>
rect 64 163 65 164 
<< m1 >>
rect 70 163 71 164 
<< m1 >>
rect 73 163 74 164 
<< m2 >>
rect 73 163 74 164 
<< m1 >>
rect 82 163 83 164 
<< m1 >>
rect 91 163 92 164 
<< m2 >>
rect 92 163 93 164 
<< m1 >>
rect 95 163 96 164 
<< m2 >>
rect 95 163 96 164 
<< m2c >>
rect 95 163 96 164 
<< m1 >>
rect 95 163 96 164 
<< m2 >>
rect 95 163 96 164 
<< m1 >>
rect 103 163 104 164 
<< m1 >>
rect 104 163 105 164 
<< m1 >>
rect 107 163 108 164 
<< m2 >>
rect 107 163 108 164 
<< m2c >>
rect 107 163 108 164 
<< m1 >>
rect 107 163 108 164 
<< m2 >>
rect 107 163 108 164 
<< m2 >>
rect 108 163 109 164 
<< m1 >>
rect 109 163 110 164 
<< m2 >>
rect 109 163 110 164 
<< m2 >>
rect 110 163 111 164 
<< m1 >>
rect 111 163 112 164 
<< m2 >>
rect 111 163 112 164 
<< m2c >>
rect 111 163 112 164 
<< m1 >>
rect 111 163 112 164 
<< m2 >>
rect 111 163 112 164 
<< m1 >>
rect 124 163 125 164 
<< m1 >>
rect 139 163 140 164 
<< m1 >>
rect 142 163 143 164 
<< m1 >>
rect 145 163 146 164 
<< m1 >>
rect 157 163 158 164 
<< m1 >>
rect 163 163 164 164 
<< m1 >>
rect 175 163 176 164 
<< m2 >>
rect 181 163 182 164 
<< m2 >>
rect 182 163 183 164 
<< m2 >>
rect 183 163 184 164 
<< m2 >>
rect 184 163 185 164 
<< m2 >>
rect 185 163 186 164 
<< m1 >>
rect 190 163 191 164 
<< m2 >>
rect 190 163 191 164 
<< m1 >>
rect 193 163 194 164 
<< m1 >>
rect 199 163 200 164 
<< m1 >>
rect 226 163 227 164 
<< m2 >>
rect 226 163 227 164 
<< m2 >>
rect 227 163 228 164 
<< m1 >>
rect 228 163 229 164 
<< m2 >>
rect 228 163 229 164 
<< m2c >>
rect 228 163 229 164 
<< m1 >>
rect 228 163 229 164 
<< m2 >>
rect 228 163 229 164 
<< m1 >>
rect 229 163 230 164 
<< m1 >>
rect 254 163 255 164 
<< m1 >>
rect 256 163 257 164 
<< m1 >>
rect 19 164 20 165 
<< m1 >>
rect 26 164 27 165 
<< m1 >>
rect 28 164 29 165 
<< m1 >>
rect 44 164 45 165 
<< m1 >>
rect 46 164 47 165 
<< m1 >>
rect 49 164 50 165 
<< m1 >>
rect 50 164 51 165 
<< m1 >>
rect 51 164 52 165 
<< m1 >>
rect 52 164 53 165 
<< m2 >>
rect 52 164 53 165 
<< m1 >>
rect 53 164 54 165 
<< m1 >>
rect 54 164 55 165 
<< m1 >>
rect 55 164 56 165 
<< m2 >>
rect 55 164 56 165 
<< m1 >>
rect 56 164 57 165 
<< m1 >>
rect 57 164 58 165 
<< m2 >>
rect 57 164 58 165 
<< m1 >>
rect 58 164 59 165 
<< m1 >>
rect 59 164 60 165 
<< m1 >>
rect 60 164 61 165 
<< m1 >>
rect 61 164 62 165 
<< m1 >>
rect 62 164 63 165 
<< m1 >>
rect 63 164 64 165 
<< m1 >>
rect 64 164 65 165 
<< m2 >>
rect 64 164 65 165 
<< m1 >>
rect 70 164 71 165 
<< m1 >>
rect 73 164 74 165 
<< m2 >>
rect 73 164 74 165 
<< m1 >>
rect 82 164 83 165 
<< m1 >>
rect 91 164 92 165 
<< m2 >>
rect 92 164 93 165 
<< m2 >>
rect 95 164 96 165 
<< m1 >>
rect 104 164 105 165 
<< m1 >>
rect 105 164 106 165 
<< m1 >>
rect 106 164 107 165 
<< m1 >>
rect 107 164 108 165 
<< m1 >>
rect 109 164 110 165 
<< m1 >>
rect 111 164 112 165 
<< m1 >>
rect 124 164 125 165 
<< m1 >>
rect 139 164 140 165 
<< m1 >>
rect 142 164 143 165 
<< m1 >>
rect 145 164 146 165 
<< m1 >>
rect 157 164 158 165 
<< m1 >>
rect 163 164 164 165 
<< m2 >>
rect 163 164 164 165 
<< m2c >>
rect 163 164 164 165 
<< m1 >>
rect 163 164 164 165 
<< m2 >>
rect 163 164 164 165 
<< m1 >>
rect 175 164 176 165 
<< m1 >>
rect 176 164 177 165 
<< m1 >>
rect 177 164 178 165 
<< m1 >>
rect 178 164 179 165 
<< m1 >>
rect 179 164 180 165 
<< m1 >>
rect 180 164 181 165 
<< m1 >>
rect 181 164 182 165 
<< m1 >>
rect 182 164 183 165 
<< m1 >>
rect 183 164 184 165 
<< m1 >>
rect 184 164 185 165 
<< m1 >>
rect 185 164 186 165 
<< m2 >>
rect 185 164 186 165 
<< m1 >>
rect 186 164 187 165 
<< m1 >>
rect 187 164 188 165 
<< m1 >>
rect 188 164 189 165 
<< m1 >>
rect 189 164 190 165 
<< m1 >>
rect 190 164 191 165 
<< m2 >>
rect 190 164 191 165 
<< m1 >>
rect 192 164 193 165 
<< m2 >>
rect 192 164 193 165 
<< m2c >>
rect 192 164 193 165 
<< m1 >>
rect 192 164 193 165 
<< m2 >>
rect 192 164 193 165 
<< m1 >>
rect 193 164 194 165 
<< m1 >>
rect 199 164 200 165 
<< m2 >>
rect 199 164 200 165 
<< m2c >>
rect 199 164 200 165 
<< m1 >>
rect 199 164 200 165 
<< m2 >>
rect 199 164 200 165 
<< m1 >>
rect 226 164 227 165 
<< m1 >>
rect 254 164 255 165 
<< m1 >>
rect 256 164 257 165 
<< m1 >>
rect 19 165 20 166 
<< m1 >>
rect 26 165 27 166 
<< m1 >>
rect 28 165 29 166 
<< m1 >>
rect 44 165 45 166 
<< m1 >>
rect 46 165 47 166 
<< m2 >>
rect 52 165 53 166 
<< m2 >>
rect 55 165 56 166 
<< m2 >>
rect 57 165 58 166 
<< m2 >>
rect 64 165 65 166 
<< m1 >>
rect 70 165 71 166 
<< m1 >>
rect 73 165 74 166 
<< m2 >>
rect 73 165 74 166 
<< m1 >>
rect 82 165 83 166 
<< m1 >>
rect 91 165 92 166 
<< m2 >>
rect 92 165 93 166 
<< m1 >>
rect 93 165 94 166 
<< m2 >>
rect 93 165 94 166 
<< m2c >>
rect 93 165 94 166 
<< m1 >>
rect 93 165 94 166 
<< m2 >>
rect 93 165 94 166 
<< m1 >>
rect 94 165 95 166 
<< m1 >>
rect 95 165 96 166 
<< m2 >>
rect 95 165 96 166 
<< m1 >>
rect 96 165 97 166 
<< m1 >>
rect 97 165 98 166 
<< m1 >>
rect 98 165 99 166 
<< m1 >>
rect 99 165 100 166 
<< m1 >>
rect 100 165 101 166 
<< m1 >>
rect 101 165 102 166 
<< m1 >>
rect 102 165 103 166 
<< m1 >>
rect 109 165 110 166 
<< m2 >>
rect 109 165 110 166 
<< m2c >>
rect 109 165 110 166 
<< m1 >>
rect 109 165 110 166 
<< m2 >>
rect 109 165 110 166 
<< m1 >>
rect 111 165 112 166 
<< m2 >>
rect 111 165 112 166 
<< m2c >>
rect 111 165 112 166 
<< m1 >>
rect 111 165 112 166 
<< m2 >>
rect 111 165 112 166 
<< m1 >>
rect 124 165 125 166 
<< m1 >>
rect 139 165 140 166 
<< m1 >>
rect 142 165 143 166 
<< m1 >>
rect 145 165 146 166 
<< m1 >>
rect 157 165 158 166 
<< m2 >>
rect 163 165 164 166 
<< m2 >>
rect 185 165 186 166 
<< m2 >>
rect 190 165 191 166 
<< m2 >>
rect 192 165 193 166 
<< m2 >>
rect 199 165 200 166 
<< m1 >>
rect 226 165 227 166 
<< m1 >>
rect 254 165 255 166 
<< m1 >>
rect 256 165 257 166 
<< m1 >>
rect 19 166 20 167 
<< m1 >>
rect 26 166 27 167 
<< m1 >>
rect 28 166 29 167 
<< m1 >>
rect 44 166 45 167 
<< m1 >>
rect 46 166 47 167 
<< m1 >>
rect 52 166 53 167 
<< m2 >>
rect 52 166 53 167 
<< m2c >>
rect 52 166 53 167 
<< m1 >>
rect 52 166 53 167 
<< m2 >>
rect 52 166 53 167 
<< m1 >>
rect 55 166 56 167 
<< m2 >>
rect 55 166 56 167 
<< m2c >>
rect 55 166 56 167 
<< m1 >>
rect 55 166 56 167 
<< m2 >>
rect 55 166 56 167 
<< m1 >>
rect 57 166 58 167 
<< m2 >>
rect 57 166 58 167 
<< m2c >>
rect 57 166 58 167 
<< m1 >>
rect 57 166 58 167 
<< m2 >>
rect 57 166 58 167 
<< m1 >>
rect 58 166 59 167 
<< m1 >>
rect 59 166 60 167 
<< m1 >>
rect 64 166 65 167 
<< m2 >>
rect 64 166 65 167 
<< m2c >>
rect 64 166 65 167 
<< m1 >>
rect 64 166 65 167 
<< m2 >>
rect 64 166 65 167 
<< m1 >>
rect 70 166 71 167 
<< m1 >>
rect 73 166 74 167 
<< m2 >>
rect 73 166 74 167 
<< m1 >>
rect 82 166 83 167 
<< m1 >>
rect 91 166 92 167 
<< m2 >>
rect 95 166 96 167 
<< m1 >>
rect 102 166 103 167 
<< m2 >>
rect 109 166 110 167 
<< m2 >>
rect 111 166 112 167 
<< m1 >>
rect 124 166 125 167 
<< m1 >>
rect 139 166 140 167 
<< m1 >>
rect 142 166 143 167 
<< m1 >>
rect 145 166 146 167 
<< m1 >>
rect 157 166 158 167 
<< m1 >>
rect 158 166 159 167 
<< m1 >>
rect 159 166 160 167 
<< m1 >>
rect 160 166 161 167 
<< m1 >>
rect 161 166 162 167 
<< m1 >>
rect 162 166 163 167 
<< m1 >>
rect 163 166 164 167 
<< m2 >>
rect 163 166 164 167 
<< m1 >>
rect 164 166 165 167 
<< m2 >>
rect 164 166 165 167 
<< m1 >>
rect 165 166 166 167 
<< m2 >>
rect 165 166 166 167 
<< m1 >>
rect 166 166 167 167 
<< m2 >>
rect 166 166 167 167 
<< m1 >>
rect 167 166 168 167 
<< m2 >>
rect 167 166 168 167 
<< m1 >>
rect 168 166 169 167 
<< m2 >>
rect 168 166 169 167 
<< m1 >>
rect 169 166 170 167 
<< m2 >>
rect 169 166 170 167 
<< m1 >>
rect 170 166 171 167 
<< m2 >>
rect 170 166 171 167 
<< m1 >>
rect 171 166 172 167 
<< m2 >>
rect 171 166 172 167 
<< m1 >>
rect 172 166 173 167 
<< m2 >>
rect 172 166 173 167 
<< m1 >>
rect 173 166 174 167 
<< m2 >>
rect 173 166 174 167 
<< m1 >>
rect 174 166 175 167 
<< m2 >>
rect 174 166 175 167 
<< m1 >>
rect 175 166 176 167 
<< m2 >>
rect 175 166 176 167 
<< m1 >>
rect 176 166 177 167 
<< m2 >>
rect 176 166 177 167 
<< m1 >>
rect 177 166 178 167 
<< m1 >>
rect 178 166 179 167 
<< m1 >>
rect 179 166 180 167 
<< m1 >>
rect 180 166 181 167 
<< m1 >>
rect 181 166 182 167 
<< m2 >>
rect 182 166 183 167 
<< m1 >>
rect 183 166 184 167 
<< m2 >>
rect 183 166 184 167 
<< m2c >>
rect 183 166 184 167 
<< m1 >>
rect 183 166 184 167 
<< m2 >>
rect 183 166 184 167 
<< m1 >>
rect 184 166 185 167 
<< m1 >>
rect 185 166 186 167 
<< m2 >>
rect 185 166 186 167 
<< m1 >>
rect 186 166 187 167 
<< m1 >>
rect 187 166 188 167 
<< m1 >>
rect 188 166 189 167 
<< m1 >>
rect 189 166 190 167 
<< m1 >>
rect 190 166 191 167 
<< m2 >>
rect 190 166 191 167 
<< m1 >>
rect 191 166 192 167 
<< m1 >>
rect 192 166 193 167 
<< m2 >>
rect 192 166 193 167 
<< m1 >>
rect 193 166 194 167 
<< m1 >>
rect 194 166 195 167 
<< m1 >>
rect 195 166 196 167 
<< m1 >>
rect 196 166 197 167 
<< m1 >>
rect 197 166 198 167 
<< m1 >>
rect 198 166 199 167 
<< m1 >>
rect 199 166 200 167 
<< m2 >>
rect 199 166 200 167 
<< m1 >>
rect 200 166 201 167 
<< m1 >>
rect 201 166 202 167 
<< m1 >>
rect 202 166 203 167 
<< m1 >>
rect 203 166 204 167 
<< m1 >>
rect 204 166 205 167 
<< m1 >>
rect 205 166 206 167 
<< m1 >>
rect 206 166 207 167 
<< m1 >>
rect 207 166 208 167 
<< m1 >>
rect 208 166 209 167 
<< m1 >>
rect 209 166 210 167 
<< m1 >>
rect 210 166 211 167 
<< m1 >>
rect 211 166 212 167 
<< m1 >>
rect 212 166 213 167 
<< m1 >>
rect 213 166 214 167 
<< m1 >>
rect 214 166 215 167 
<< m1 >>
rect 215 166 216 167 
<< m1 >>
rect 216 166 217 167 
<< m1 >>
rect 217 166 218 167 
<< m1 >>
rect 218 166 219 167 
<< m1 >>
rect 219 166 220 167 
<< m1 >>
rect 220 166 221 167 
<< m1 >>
rect 221 166 222 167 
<< m1 >>
rect 222 166 223 167 
<< m1 >>
rect 223 166 224 167 
<< m1 >>
rect 224 166 225 167 
<< m1 >>
rect 225 166 226 167 
<< m1 >>
rect 226 166 227 167 
<< m1 >>
rect 254 166 255 167 
<< m1 >>
rect 256 166 257 167 
<< m1 >>
rect 19 167 20 168 
<< m1 >>
rect 26 167 27 168 
<< m1 >>
rect 28 167 29 168 
<< m1 >>
rect 44 167 45 168 
<< m1 >>
rect 46 167 47 168 
<< m1 >>
rect 52 167 53 168 
<< m1 >>
rect 55 167 56 168 
<< m1 >>
rect 59 167 60 168 
<< m1 >>
rect 64 167 65 168 
<< m1 >>
rect 70 167 71 168 
<< m1 >>
rect 73 167 74 168 
<< m2 >>
rect 73 167 74 168 
<< m1 >>
rect 82 167 83 168 
<< m2 >>
rect 82 167 83 168 
<< m2c >>
rect 82 167 83 168 
<< m1 >>
rect 82 167 83 168 
<< m2 >>
rect 82 167 83 168 
<< m1 >>
rect 91 167 92 168 
<< m2 >>
rect 91 167 92 168 
<< m2c >>
rect 91 167 92 168 
<< m1 >>
rect 91 167 92 168 
<< m2 >>
rect 91 167 92 168 
<< m1 >>
rect 93 167 94 168 
<< m2 >>
rect 93 167 94 168 
<< m2c >>
rect 93 167 94 168 
<< m1 >>
rect 93 167 94 168 
<< m2 >>
rect 93 167 94 168 
<< m1 >>
rect 94 167 95 168 
<< m1 >>
rect 95 167 96 168 
<< m2 >>
rect 95 167 96 168 
<< m2c >>
rect 95 167 96 168 
<< m1 >>
rect 95 167 96 168 
<< m2 >>
rect 95 167 96 168 
<< m1 >>
rect 102 167 103 168 
<< m1 >>
rect 103 167 104 168 
<< m1 >>
rect 104 167 105 168 
<< m1 >>
rect 105 167 106 168 
<< m1 >>
rect 106 167 107 168 
<< m1 >>
rect 107 167 108 168 
<< m1 >>
rect 108 167 109 168 
<< m1 >>
rect 109 167 110 168 
<< m2 >>
rect 109 167 110 168 
<< m1 >>
rect 110 167 111 168 
<< m1 >>
rect 111 167 112 168 
<< m2 >>
rect 111 167 112 168 
<< m1 >>
rect 112 167 113 168 
<< m1 >>
rect 113 167 114 168 
<< m1 >>
rect 114 167 115 168 
<< m1 >>
rect 115 167 116 168 
<< m1 >>
rect 116 167 117 168 
<< m1 >>
rect 117 167 118 168 
<< m1 >>
rect 118 167 119 168 
<< m1 >>
rect 119 167 120 168 
<< m1 >>
rect 120 167 121 168 
<< m1 >>
rect 121 167 122 168 
<< m1 >>
rect 122 167 123 168 
<< m2 >>
rect 122 167 123 168 
<< m2c >>
rect 122 167 123 168 
<< m1 >>
rect 122 167 123 168 
<< m2 >>
rect 122 167 123 168 
<< m2 >>
rect 123 167 124 168 
<< m1 >>
rect 124 167 125 168 
<< m2 >>
rect 124 167 125 168 
<< m2 >>
rect 125 167 126 168 
<< m1 >>
rect 139 167 140 168 
<< m1 >>
rect 142 167 143 168 
<< m1 >>
rect 145 167 146 168 
<< m2 >>
rect 176 167 177 168 
<< m1 >>
rect 181 167 182 168 
<< m2 >>
rect 182 167 183 168 
<< m2 >>
rect 185 167 186 168 
<< m2 >>
rect 190 167 191 168 
<< m2 >>
rect 192 167 193 168 
<< m2 >>
rect 199 167 200 168 
<< m1 >>
rect 254 167 255 168 
<< m1 >>
rect 256 167 257 168 
<< m1 >>
rect 19 168 20 169 
<< m1 >>
rect 26 168 27 169 
<< m1 >>
rect 28 168 29 169 
<< m1 >>
rect 44 168 45 169 
<< m1 >>
rect 46 168 47 169 
<< m1 >>
rect 52 168 53 169 
<< m1 >>
rect 55 168 56 169 
<< m1 >>
rect 59 168 60 169 
<< m1 >>
rect 64 168 65 169 
<< m1 >>
rect 70 168 71 169 
<< m1 >>
rect 73 168 74 169 
<< m2 >>
rect 73 168 74 169 
<< m2 >>
rect 82 168 83 169 
<< m2 >>
rect 91 168 92 169 
<< m2 >>
rect 93 168 94 169 
<< m2 >>
rect 109 168 110 169 
<< m2 >>
rect 111 168 112 169 
<< m1 >>
rect 124 168 125 169 
<< m2 >>
rect 125 168 126 169 
<< m1 >>
rect 139 168 140 169 
<< m1 >>
rect 142 168 143 169 
<< m1 >>
rect 145 168 146 169 
<< m1 >>
rect 175 168 176 169 
<< m1 >>
rect 176 168 177 169 
<< m2 >>
rect 176 168 177 169 
<< m1 >>
rect 177 168 178 169 
<< m1 >>
rect 178 168 179 169 
<< m1 >>
rect 179 168 180 169 
<< m2 >>
rect 179 168 180 169 
<< m2c >>
rect 179 168 180 169 
<< m1 >>
rect 179 168 180 169 
<< m2 >>
rect 179 168 180 169 
<< m2 >>
rect 180 168 181 169 
<< m1 >>
rect 181 168 182 169 
<< m2 >>
rect 181 168 182 169 
<< m2 >>
rect 182 168 183 169 
<< m1 >>
rect 185 168 186 169 
<< m2 >>
rect 185 168 186 169 
<< m2c >>
rect 185 168 186 169 
<< m1 >>
rect 185 168 186 169 
<< m2 >>
rect 185 168 186 169 
<< m1 >>
rect 190 168 191 169 
<< m2 >>
rect 190 168 191 169 
<< m2c >>
rect 190 168 191 169 
<< m1 >>
rect 190 168 191 169 
<< m2 >>
rect 190 168 191 169 
<< m1 >>
rect 192 168 193 169 
<< m2 >>
rect 192 168 193 169 
<< m2c >>
rect 192 168 193 169 
<< m1 >>
rect 192 168 193 169 
<< m2 >>
rect 192 168 193 169 
<< m2 >>
rect 199 168 200 169 
<< m1 >>
rect 254 168 255 169 
<< m1 >>
rect 256 168 257 169 
<< m1 >>
rect 19 169 20 170 
<< m1 >>
rect 26 169 27 170 
<< m2 >>
rect 26 169 27 170 
<< m2c >>
rect 26 169 27 170 
<< m1 >>
rect 26 169 27 170 
<< m2 >>
rect 26 169 27 170 
<< m2 >>
rect 27 169 28 170 
<< m1 >>
rect 28 169 29 170 
<< m2 >>
rect 28 169 29 170 
<< m2 >>
rect 29 169 30 170 
<< m1 >>
rect 30 169 31 170 
<< m2 >>
rect 30 169 31 170 
<< m2c >>
rect 30 169 31 170 
<< m1 >>
rect 30 169 31 170 
<< m2 >>
rect 30 169 31 170 
<< m1 >>
rect 31 169 32 170 
<< m1 >>
rect 32 169 33 170 
<< m1 >>
rect 33 169 34 170 
<< m1 >>
rect 34 169 35 170 
<< m1 >>
rect 35 169 36 170 
<< m1 >>
rect 36 169 37 170 
<< m1 >>
rect 37 169 38 170 
<< m1 >>
rect 38 169 39 170 
<< m1 >>
rect 39 169 40 170 
<< m1 >>
rect 40 169 41 170 
<< m1 >>
rect 41 169 42 170 
<< m1 >>
rect 42 169 43 170 
<< m2 >>
rect 42 169 43 170 
<< m2c >>
rect 42 169 43 170 
<< m1 >>
rect 42 169 43 170 
<< m2 >>
rect 42 169 43 170 
<< m2 >>
rect 43 169 44 170 
<< m1 >>
rect 44 169 45 170 
<< m2 >>
rect 44 169 45 170 
<< m2 >>
rect 45 169 46 170 
<< m1 >>
rect 46 169 47 170 
<< m2 >>
rect 46 169 47 170 
<< m2 >>
rect 47 169 48 170 
<< m1 >>
rect 48 169 49 170 
<< m2 >>
rect 48 169 49 170 
<< m2c >>
rect 48 169 49 170 
<< m1 >>
rect 48 169 49 170 
<< m2 >>
rect 48 169 49 170 
<< m1 >>
rect 49 169 50 170 
<< m1 >>
rect 50 169 51 170 
<< m1 >>
rect 52 169 53 170 
<< m1 >>
rect 55 169 56 170 
<< m1 >>
rect 59 169 60 170 
<< m1 >>
rect 64 169 65 170 
<< m1 >>
rect 70 169 71 170 
<< m1 >>
rect 73 169 74 170 
<< m2 >>
rect 73 169 74 170 
<< m1 >>
rect 75 169 76 170 
<< m1 >>
rect 76 169 77 170 
<< m1 >>
rect 77 169 78 170 
<< m1 >>
rect 78 169 79 170 
<< m1 >>
rect 79 169 80 170 
<< m1 >>
rect 80 169 81 170 
<< m1 >>
rect 81 169 82 170 
<< m1 >>
rect 82 169 83 170 
<< m2 >>
rect 82 169 83 170 
<< m1 >>
rect 83 169 84 170 
<< m1 >>
rect 84 169 85 170 
<< m1 >>
rect 85 169 86 170 
<< m1 >>
rect 86 169 87 170 
<< m1 >>
rect 87 169 88 170 
<< m1 >>
rect 88 169 89 170 
<< m1 >>
rect 89 169 90 170 
<< m1 >>
rect 90 169 91 170 
<< m1 >>
rect 91 169 92 170 
<< m2 >>
rect 91 169 92 170 
<< m1 >>
rect 92 169 93 170 
<< m1 >>
rect 93 169 94 170 
<< m2 >>
rect 93 169 94 170 
<< m1 >>
rect 94 169 95 170 
<< m1 >>
rect 95 169 96 170 
<< m1 >>
rect 96 169 97 170 
<< m1 >>
rect 97 169 98 170 
<< m1 >>
rect 98 169 99 170 
<< m1 >>
rect 99 169 100 170 
<< m1 >>
rect 100 169 101 170 
<< m1 >>
rect 101 169 102 170 
<< m1 >>
rect 102 169 103 170 
<< m1 >>
rect 103 169 104 170 
<< m1 >>
rect 104 169 105 170 
<< m1 >>
rect 105 169 106 170 
<< m1 >>
rect 106 169 107 170 
<< m1 >>
rect 107 169 108 170 
<< m1 >>
rect 108 169 109 170 
<< m1 >>
rect 109 169 110 170 
<< m2 >>
rect 109 169 110 170 
<< m1 >>
rect 110 169 111 170 
<< m1 >>
rect 111 169 112 170 
<< m2 >>
rect 111 169 112 170 
<< m1 >>
rect 112 169 113 170 
<< m2 >>
rect 112 169 113 170 
<< m1 >>
rect 113 169 114 170 
<< m2 >>
rect 113 169 114 170 
<< m1 >>
rect 114 169 115 170 
<< m2 >>
rect 114 169 115 170 
<< m1 >>
rect 115 169 116 170 
<< m2 >>
rect 115 169 116 170 
<< m1 >>
rect 116 169 117 170 
<< m2 >>
rect 116 169 117 170 
<< m1 >>
rect 117 169 118 170 
<< m2 >>
rect 117 169 118 170 
<< m1 >>
rect 118 169 119 170 
<< m2 >>
rect 118 169 119 170 
<< m1 >>
rect 119 169 120 170 
<< m2 >>
rect 119 169 120 170 
<< m1 >>
rect 120 169 121 170 
<< m2 >>
rect 120 169 121 170 
<< m1 >>
rect 121 169 122 170 
<< m2 >>
rect 121 169 122 170 
<< m1 >>
rect 122 169 123 170 
<< m2 >>
rect 122 169 123 170 
<< m1 >>
rect 123 169 124 170 
<< m1 >>
rect 124 169 125 170 
<< m2 >>
rect 125 169 126 170 
<< m1 >>
rect 127 169 128 170 
<< m1 >>
rect 128 169 129 170 
<< m1 >>
rect 129 169 130 170 
<< m1 >>
rect 130 169 131 170 
<< m1 >>
rect 131 169 132 170 
<< m1 >>
rect 132 169 133 170 
<< m1 >>
rect 133 169 134 170 
<< m1 >>
rect 134 169 135 170 
<< m1 >>
rect 135 169 136 170 
<< m1 >>
rect 136 169 137 170 
<< m1 >>
rect 137 169 138 170 
<< m1 >>
rect 138 169 139 170 
<< m1 >>
rect 139 169 140 170 
<< m1 >>
rect 142 169 143 170 
<< m1 >>
rect 145 169 146 170 
<< m1 >>
rect 175 169 176 170 
<< m2 >>
rect 176 169 177 170 
<< m1 >>
rect 181 169 182 170 
<< m1 >>
rect 185 169 186 170 
<< m1 >>
rect 190 169 191 170 
<< m1 >>
rect 192 169 193 170 
<< m1 >>
rect 199 169 200 170 
<< m2 >>
rect 199 169 200 170 
<< m1 >>
rect 200 169 201 170 
<< m1 >>
rect 201 169 202 170 
<< m1 >>
rect 202 169 203 170 
<< m1 >>
rect 203 169 204 170 
<< m1 >>
rect 204 169 205 170 
<< m1 >>
rect 205 169 206 170 
<< m1 >>
rect 206 169 207 170 
<< m1 >>
rect 207 169 208 170 
<< m1 >>
rect 208 169 209 170 
<< m1 >>
rect 209 169 210 170 
<< m1 >>
rect 210 169 211 170 
<< m1 >>
rect 211 169 212 170 
<< m1 >>
rect 212 169 213 170 
<< m1 >>
rect 213 169 214 170 
<< m1 >>
rect 214 169 215 170 
<< m1 >>
rect 254 169 255 170 
<< m1 >>
rect 256 169 257 170 
<< m1 >>
rect 19 170 20 171 
<< m1 >>
rect 28 170 29 171 
<< m1 >>
rect 44 170 45 171 
<< m1 >>
rect 46 170 47 171 
<< m1 >>
rect 50 170 51 171 
<< m1 >>
rect 52 170 53 171 
<< m1 >>
rect 55 170 56 171 
<< m1 >>
rect 59 170 60 171 
<< m1 >>
rect 64 170 65 171 
<< m1 >>
rect 70 170 71 171 
<< m1 >>
rect 73 170 74 171 
<< m2 >>
rect 73 170 74 171 
<< m1 >>
rect 75 170 76 171 
<< m2 >>
rect 82 170 83 171 
<< m2 >>
rect 91 170 92 171 
<< m2 >>
rect 93 170 94 171 
<< m2 >>
rect 109 170 110 171 
<< m2 >>
rect 122 170 123 171 
<< m2 >>
rect 125 170 126 171 
<< m2 >>
rect 126 170 127 171 
<< m1 >>
rect 127 170 128 171 
<< m2 >>
rect 127 170 128 171 
<< m2 >>
rect 128 170 129 171 
<< m2 >>
rect 129 170 130 171 
<< m2 >>
rect 130 170 131 171 
<< m2 >>
rect 131 170 132 171 
<< m2 >>
rect 132 170 133 171 
<< m2 >>
rect 133 170 134 171 
<< m2 >>
rect 134 170 135 171 
<< m2 >>
rect 135 170 136 171 
<< m2 >>
rect 136 170 137 171 
<< m1 >>
rect 142 170 143 171 
<< m1 >>
rect 145 170 146 171 
<< m1 >>
rect 175 170 176 171 
<< m2 >>
rect 176 170 177 171 
<< m1 >>
rect 177 170 178 171 
<< m2 >>
rect 177 170 178 171 
<< m2c >>
rect 177 170 178 171 
<< m1 >>
rect 177 170 178 171 
<< m2 >>
rect 177 170 178 171 
<< m1 >>
rect 178 170 179 171 
<< m1 >>
rect 179 170 180 171 
<< m2 >>
rect 179 170 180 171 
<< m2c >>
rect 179 170 180 171 
<< m1 >>
rect 179 170 180 171 
<< m2 >>
rect 179 170 180 171 
<< m2 >>
rect 180 170 181 171 
<< m1 >>
rect 181 170 182 171 
<< m2 >>
rect 181 170 182 171 
<< m2 >>
rect 182 170 183 171 
<< m1 >>
rect 183 170 184 171 
<< m2 >>
rect 183 170 184 171 
<< m2c >>
rect 183 170 184 171 
<< m1 >>
rect 183 170 184 171 
<< m2 >>
rect 183 170 184 171 
<< m1 >>
rect 185 170 186 171 
<< m1 >>
rect 190 170 191 171 
<< m1 >>
rect 192 170 193 171 
<< m1 >>
rect 199 170 200 171 
<< m2 >>
rect 199 170 200 171 
<< m1 >>
rect 214 170 215 171 
<< m1 >>
rect 254 170 255 171 
<< m1 >>
rect 256 170 257 171 
<< m1 >>
rect 19 171 20 172 
<< m1 >>
rect 28 171 29 172 
<< m1 >>
rect 44 171 45 172 
<< m1 >>
rect 46 171 47 172 
<< m1 >>
rect 50 171 51 172 
<< m2 >>
rect 50 171 51 172 
<< m2c >>
rect 50 171 51 172 
<< m1 >>
rect 50 171 51 172 
<< m2 >>
rect 50 171 51 172 
<< m2 >>
rect 51 171 52 172 
<< m1 >>
rect 52 171 53 172 
<< m2 >>
rect 52 171 53 172 
<< m2 >>
rect 53 171 54 172 
<< m2 >>
rect 54 171 55 172 
<< m1 >>
rect 55 171 56 172 
<< m2 >>
rect 55 171 56 172 
<< m2 >>
rect 56 171 57 172 
<< m1 >>
rect 59 171 60 172 
<< m1 >>
rect 64 171 65 172 
<< m1 >>
rect 70 171 71 172 
<< m1 >>
rect 73 171 74 172 
<< m2 >>
rect 73 171 74 172 
<< m2 >>
rect 74 171 75 172 
<< m1 >>
rect 75 171 76 172 
<< m2 >>
rect 75 171 76 172 
<< m2 >>
rect 76 171 77 172 
<< m1 >>
rect 77 171 78 172 
<< m2 >>
rect 77 171 78 172 
<< m2c >>
rect 77 171 78 172 
<< m1 >>
rect 77 171 78 172 
<< m2 >>
rect 77 171 78 172 
<< m1 >>
rect 78 171 79 172 
<< m1 >>
rect 79 171 80 172 
<< m1 >>
rect 80 171 81 172 
<< m1 >>
rect 81 171 82 172 
<< m1 >>
rect 82 171 83 172 
<< m2 >>
rect 82 171 83 172 
<< m1 >>
rect 83 171 84 172 
<< m1 >>
rect 84 171 85 172 
<< m1 >>
rect 85 171 86 172 
<< m1 >>
rect 91 171 92 172 
<< m2 >>
rect 91 171 92 172 
<< m2c >>
rect 91 171 92 172 
<< m1 >>
rect 91 171 92 172 
<< m2 >>
rect 91 171 92 172 
<< m1 >>
rect 93 171 94 172 
<< m2 >>
rect 93 171 94 172 
<< m2c >>
rect 93 171 94 172 
<< m1 >>
rect 93 171 94 172 
<< m2 >>
rect 93 171 94 172 
<< m2 >>
rect 109 171 110 172 
<< m2 >>
rect 122 171 123 172 
<< m1 >>
rect 123 171 124 172 
<< m2 >>
rect 123 171 124 172 
<< m2c >>
rect 123 171 124 172 
<< m1 >>
rect 123 171 124 172 
<< m2 >>
rect 123 171 124 172 
<< m1 >>
rect 124 171 125 172 
<< m1 >>
rect 125 171 126 172 
<< m1 >>
rect 127 171 128 172 
<< m1 >>
rect 136 171 137 172 
<< m2 >>
rect 136 171 137 172 
<< m2c >>
rect 136 171 137 172 
<< m1 >>
rect 136 171 137 172 
<< m2 >>
rect 136 171 137 172 
<< m1 >>
rect 142 171 143 172 
<< m1 >>
rect 143 171 144 172 
<< m1 >>
rect 145 171 146 172 
<< m1 >>
rect 175 171 176 172 
<< m1 >>
rect 181 171 182 172 
<< m1 >>
rect 183 171 184 172 
<< m1 >>
rect 185 171 186 172 
<< m1 >>
rect 190 171 191 172 
<< m1 >>
rect 192 171 193 172 
<< m1 >>
rect 199 171 200 172 
<< m2 >>
rect 199 171 200 172 
<< m1 >>
rect 214 171 215 172 
<< m1 >>
rect 254 171 255 172 
<< m1 >>
rect 256 171 257 172 
<< m1 >>
rect 19 172 20 173 
<< m1 >>
rect 28 172 29 173 
<< m1 >>
rect 44 172 45 173 
<< m1 >>
rect 46 172 47 173 
<< m1 >>
rect 52 172 53 173 
<< m1 >>
rect 55 172 56 173 
<< m2 >>
rect 56 172 57 173 
<< m1 >>
rect 59 172 60 173 
<< m1 >>
rect 64 172 65 173 
<< m1 >>
rect 70 172 71 173 
<< m1 >>
rect 73 172 74 173 
<< m1 >>
rect 75 172 76 173 
<< m2 >>
rect 82 172 83 173 
<< m1 >>
rect 85 172 86 173 
<< m1 >>
rect 91 172 92 173 
<< m1 >>
rect 93 172 94 173 
<< m1 >>
rect 106 172 107 173 
<< m1 >>
rect 107 172 108 173 
<< m1 >>
rect 108 172 109 173 
<< m1 >>
rect 109 172 110 173 
<< m2 >>
rect 109 172 110 173 
<< m1 >>
rect 111 172 112 173 
<< m1 >>
rect 112 172 113 173 
<< m1 >>
rect 113 172 114 173 
<< m1 >>
rect 114 172 115 173 
<< m1 >>
rect 115 172 116 173 
<< m1 >>
rect 116 172 117 173 
<< m1 >>
rect 117 172 118 173 
<< m1 >>
rect 118 172 119 173 
<< m1 >>
rect 119 172 120 173 
<< m1 >>
rect 120 172 121 173 
<< m1 >>
rect 121 172 122 173 
<< m1 >>
rect 125 172 126 173 
<< m2 >>
rect 125 172 126 173 
<< m2c >>
rect 125 172 126 173 
<< m1 >>
rect 125 172 126 173 
<< m2 >>
rect 125 172 126 173 
<< m2 >>
rect 126 172 127 173 
<< m1 >>
rect 127 172 128 173 
<< m2 >>
rect 127 172 128 173 
<< m2 >>
rect 128 172 129 173 
<< m1 >>
rect 129 172 130 173 
<< m2 >>
rect 129 172 130 173 
<< m2c >>
rect 129 172 130 173 
<< m1 >>
rect 129 172 130 173 
<< m2 >>
rect 129 172 130 173 
<< m1 >>
rect 136 172 137 173 
<< m1 >>
rect 143 172 144 173 
<< m2 >>
rect 143 172 144 173 
<< m2c >>
rect 143 172 144 173 
<< m1 >>
rect 143 172 144 173 
<< m2 >>
rect 143 172 144 173 
<< m2 >>
rect 144 172 145 173 
<< m1 >>
rect 145 172 146 173 
<< m2 >>
rect 145 172 146 173 
<< m2 >>
rect 146 172 147 173 
<< m1 >>
rect 147 172 148 173 
<< m2 >>
rect 147 172 148 173 
<< m2c >>
rect 147 172 148 173 
<< m1 >>
rect 147 172 148 173 
<< m2 >>
rect 147 172 148 173 
<< m1 >>
rect 148 172 149 173 
<< m1 >>
rect 149 172 150 173 
<< m1 >>
rect 150 172 151 173 
<< m1 >>
rect 151 172 152 173 
<< m1 >>
rect 152 172 153 173 
<< m1 >>
rect 153 172 154 173 
<< m1 >>
rect 154 172 155 173 
<< m1 >>
rect 155 172 156 173 
<< m1 >>
rect 156 172 157 173 
<< m1 >>
rect 157 172 158 173 
<< m1 >>
rect 175 172 176 173 
<< m1 >>
rect 181 172 182 173 
<< m1 >>
rect 183 172 184 173 
<< m1 >>
rect 185 172 186 173 
<< m2 >>
rect 189 172 190 173 
<< m1 >>
rect 190 172 191 173 
<< m2 >>
rect 190 172 191 173 
<< m2 >>
rect 191 172 192 173 
<< m1 >>
rect 192 172 193 173 
<< m2 >>
rect 192 172 193 173 
<< m2c >>
rect 192 172 193 173 
<< m1 >>
rect 192 172 193 173 
<< m2 >>
rect 192 172 193 173 
<< m1 >>
rect 199 172 200 173 
<< m2 >>
rect 199 172 200 173 
<< m1 >>
rect 214 172 215 173 
<< m1 >>
rect 254 172 255 173 
<< m1 >>
rect 256 172 257 173 
<< m1 >>
rect 19 173 20 174 
<< m1 >>
rect 28 173 29 174 
<< m1 >>
rect 44 173 45 174 
<< m1 >>
rect 46 173 47 174 
<< m1 >>
rect 52 173 53 174 
<< m1 >>
rect 55 173 56 174 
<< m2 >>
rect 56 173 57 174 
<< m1 >>
rect 59 173 60 174 
<< m1 >>
rect 64 173 65 174 
<< m1 >>
rect 70 173 71 174 
<< m1 >>
rect 73 173 74 174 
<< m1 >>
rect 75 173 76 174 
<< m1 >>
rect 82 173 83 174 
<< m2 >>
rect 82 173 83 174 
<< m2c >>
rect 82 173 83 174 
<< m1 >>
rect 82 173 83 174 
<< m2 >>
rect 82 173 83 174 
<< m1 >>
rect 85 173 86 174 
<< m1 >>
rect 91 173 92 174 
<< m1 >>
rect 93 173 94 174 
<< m1 >>
rect 106 173 107 174 
<< m1 >>
rect 109 173 110 174 
<< m2 >>
rect 109 173 110 174 
<< m1 >>
rect 111 173 112 174 
<< m1 >>
rect 121 173 122 174 
<< m1 >>
rect 127 173 128 174 
<< m1 >>
rect 129 173 130 174 
<< m1 >>
rect 136 173 137 174 
<< m1 >>
rect 145 173 146 174 
<< m1 >>
rect 157 173 158 174 
<< m1 >>
rect 175 173 176 174 
<< m1 >>
rect 181 173 182 174 
<< m1 >>
rect 183 173 184 174 
<< m1 >>
rect 185 173 186 174 
<< m2 >>
rect 189 173 190 174 
<< m1 >>
rect 190 173 191 174 
<< m1 >>
rect 199 173 200 174 
<< m2 >>
rect 199 173 200 174 
<< m1 >>
rect 214 173 215 174 
<< m1 >>
rect 254 173 255 174 
<< m1 >>
rect 256 173 257 174 
<< pdiffusion >>
rect 12 174 13 175 
<< pdiffusion >>
rect 13 174 14 175 
<< pdiffusion >>
rect 14 174 15 175 
<< pdiffusion >>
rect 15 174 16 175 
<< pdiffusion >>
rect 16 174 17 175 
<< pdiffusion >>
rect 17 174 18 175 
<< m1 >>
rect 19 174 20 175 
<< m1 >>
rect 28 174 29 175 
<< pdiffusion >>
rect 30 174 31 175 
<< pdiffusion >>
rect 31 174 32 175 
<< pdiffusion >>
rect 32 174 33 175 
<< pdiffusion >>
rect 33 174 34 175 
<< pdiffusion >>
rect 34 174 35 175 
<< pdiffusion >>
rect 35 174 36 175 
<< m1 >>
rect 44 174 45 175 
<< m1 >>
rect 46 174 47 175 
<< pdiffusion >>
rect 48 174 49 175 
<< pdiffusion >>
rect 49 174 50 175 
<< pdiffusion >>
rect 50 174 51 175 
<< pdiffusion >>
rect 51 174 52 175 
<< m1 >>
rect 52 174 53 175 
<< pdiffusion >>
rect 52 174 53 175 
<< pdiffusion >>
rect 53 174 54 175 
<< m1 >>
rect 55 174 56 175 
<< m2 >>
rect 56 174 57 175 
<< m1 >>
rect 59 174 60 175 
<< m1 >>
rect 64 174 65 175 
<< pdiffusion >>
rect 66 174 67 175 
<< pdiffusion >>
rect 67 174 68 175 
<< pdiffusion >>
rect 68 174 69 175 
<< pdiffusion >>
rect 69 174 70 175 
<< m1 >>
rect 70 174 71 175 
<< pdiffusion >>
rect 70 174 71 175 
<< pdiffusion >>
rect 71 174 72 175 
<< m1 >>
rect 73 174 74 175 
<< m1 >>
rect 75 174 76 175 
<< m1 >>
rect 82 174 83 175 
<< pdiffusion >>
rect 84 174 85 175 
<< m1 >>
rect 85 174 86 175 
<< pdiffusion >>
rect 85 174 86 175 
<< pdiffusion >>
rect 86 174 87 175 
<< pdiffusion >>
rect 87 174 88 175 
<< pdiffusion >>
rect 88 174 89 175 
<< pdiffusion >>
rect 89 174 90 175 
<< m1 >>
rect 91 174 92 175 
<< m1 >>
rect 93 174 94 175 
<< pdiffusion >>
rect 102 174 103 175 
<< pdiffusion >>
rect 103 174 104 175 
<< pdiffusion >>
rect 104 174 105 175 
<< pdiffusion >>
rect 105 174 106 175 
<< m1 >>
rect 106 174 107 175 
<< pdiffusion >>
rect 106 174 107 175 
<< pdiffusion >>
rect 107 174 108 175 
<< m1 >>
rect 109 174 110 175 
<< m2 >>
rect 109 174 110 175 
<< m2 >>
rect 110 174 111 175 
<< m1 >>
rect 111 174 112 175 
<< m2 >>
rect 111 174 112 175 
<< m2 >>
rect 112 174 113 175 
<< m1 >>
rect 113 174 114 175 
<< m2 >>
rect 113 174 114 175 
<< m2c >>
rect 113 174 114 175 
<< m1 >>
rect 113 174 114 175 
<< m2 >>
rect 113 174 114 175 
<< pdiffusion >>
rect 120 174 121 175 
<< m1 >>
rect 121 174 122 175 
<< pdiffusion >>
rect 121 174 122 175 
<< pdiffusion >>
rect 122 174 123 175 
<< pdiffusion >>
rect 123 174 124 175 
<< pdiffusion >>
rect 124 174 125 175 
<< pdiffusion >>
rect 125 174 126 175 
<< m1 >>
rect 127 174 128 175 
<< m1 >>
rect 129 174 130 175 
<< m1 >>
rect 136 174 137 175 
<< pdiffusion >>
rect 138 174 139 175 
<< pdiffusion >>
rect 139 174 140 175 
<< pdiffusion >>
rect 140 174 141 175 
<< pdiffusion >>
rect 141 174 142 175 
<< pdiffusion >>
rect 142 174 143 175 
<< pdiffusion >>
rect 143 174 144 175 
<< m1 >>
rect 145 174 146 175 
<< pdiffusion >>
rect 156 174 157 175 
<< m1 >>
rect 157 174 158 175 
<< pdiffusion >>
rect 157 174 158 175 
<< pdiffusion >>
rect 158 174 159 175 
<< pdiffusion >>
rect 159 174 160 175 
<< pdiffusion >>
rect 160 174 161 175 
<< pdiffusion >>
rect 161 174 162 175 
<< pdiffusion >>
rect 174 174 175 175 
<< m1 >>
rect 175 174 176 175 
<< pdiffusion >>
rect 175 174 176 175 
<< pdiffusion >>
rect 176 174 177 175 
<< pdiffusion >>
rect 177 174 178 175 
<< pdiffusion >>
rect 178 174 179 175 
<< pdiffusion >>
rect 179 174 180 175 
<< m1 >>
rect 181 174 182 175 
<< m1 >>
rect 183 174 184 175 
<< m1 >>
rect 185 174 186 175 
<< m2 >>
rect 189 174 190 175 
<< m1 >>
rect 190 174 191 175 
<< pdiffusion >>
rect 192 174 193 175 
<< pdiffusion >>
rect 193 174 194 175 
<< pdiffusion >>
rect 194 174 195 175 
<< pdiffusion >>
rect 195 174 196 175 
<< pdiffusion >>
rect 196 174 197 175 
<< pdiffusion >>
rect 197 174 198 175 
<< m1 >>
rect 199 174 200 175 
<< m2 >>
rect 199 174 200 175 
<< pdiffusion >>
rect 210 174 211 175 
<< pdiffusion >>
rect 211 174 212 175 
<< pdiffusion >>
rect 212 174 213 175 
<< pdiffusion >>
rect 213 174 214 175 
<< m1 >>
rect 214 174 215 175 
<< pdiffusion >>
rect 214 174 215 175 
<< pdiffusion >>
rect 215 174 216 175 
<< pdiffusion >>
rect 228 174 229 175 
<< pdiffusion >>
rect 229 174 230 175 
<< pdiffusion >>
rect 230 174 231 175 
<< pdiffusion >>
rect 231 174 232 175 
<< pdiffusion >>
rect 232 174 233 175 
<< pdiffusion >>
rect 233 174 234 175 
<< m1 >>
rect 254 174 255 175 
<< m1 >>
rect 256 174 257 175 
<< pdiffusion >>
rect 12 175 13 176 
<< pdiffusion >>
rect 13 175 14 176 
<< pdiffusion >>
rect 14 175 15 176 
<< pdiffusion >>
rect 15 175 16 176 
<< pdiffusion >>
rect 16 175 17 176 
<< pdiffusion >>
rect 17 175 18 176 
<< m1 >>
rect 19 175 20 176 
<< m1 >>
rect 28 175 29 176 
<< pdiffusion >>
rect 30 175 31 176 
<< pdiffusion >>
rect 31 175 32 176 
<< pdiffusion >>
rect 32 175 33 176 
<< pdiffusion >>
rect 33 175 34 176 
<< pdiffusion >>
rect 34 175 35 176 
<< pdiffusion >>
rect 35 175 36 176 
<< m1 >>
rect 44 175 45 176 
<< m1 >>
rect 46 175 47 176 
<< pdiffusion >>
rect 48 175 49 176 
<< pdiffusion >>
rect 49 175 50 176 
<< pdiffusion >>
rect 50 175 51 176 
<< pdiffusion >>
rect 51 175 52 176 
<< pdiffusion >>
rect 52 175 53 176 
<< pdiffusion >>
rect 53 175 54 176 
<< m1 >>
rect 55 175 56 176 
<< m2 >>
rect 56 175 57 176 
<< m1 >>
rect 59 175 60 176 
<< m1 >>
rect 64 175 65 176 
<< pdiffusion >>
rect 66 175 67 176 
<< pdiffusion >>
rect 67 175 68 176 
<< pdiffusion >>
rect 68 175 69 176 
<< pdiffusion >>
rect 69 175 70 176 
<< pdiffusion >>
rect 70 175 71 176 
<< pdiffusion >>
rect 71 175 72 176 
<< m1 >>
rect 73 175 74 176 
<< m1 >>
rect 75 175 76 176 
<< m1 >>
rect 82 175 83 176 
<< pdiffusion >>
rect 84 175 85 176 
<< pdiffusion >>
rect 85 175 86 176 
<< pdiffusion >>
rect 86 175 87 176 
<< pdiffusion >>
rect 87 175 88 176 
<< pdiffusion >>
rect 88 175 89 176 
<< pdiffusion >>
rect 89 175 90 176 
<< m1 >>
rect 91 175 92 176 
<< m1 >>
rect 93 175 94 176 
<< pdiffusion >>
rect 102 175 103 176 
<< pdiffusion >>
rect 103 175 104 176 
<< pdiffusion >>
rect 104 175 105 176 
<< pdiffusion >>
rect 105 175 106 176 
<< pdiffusion >>
rect 106 175 107 176 
<< pdiffusion >>
rect 107 175 108 176 
<< m1 >>
rect 109 175 110 176 
<< m1 >>
rect 111 175 112 176 
<< m1 >>
rect 113 175 114 176 
<< pdiffusion >>
rect 120 175 121 176 
<< pdiffusion >>
rect 121 175 122 176 
<< pdiffusion >>
rect 122 175 123 176 
<< pdiffusion >>
rect 123 175 124 176 
<< pdiffusion >>
rect 124 175 125 176 
<< pdiffusion >>
rect 125 175 126 176 
<< m1 >>
rect 127 175 128 176 
<< m1 >>
rect 129 175 130 176 
<< m1 >>
rect 136 175 137 176 
<< pdiffusion >>
rect 138 175 139 176 
<< pdiffusion >>
rect 139 175 140 176 
<< pdiffusion >>
rect 140 175 141 176 
<< pdiffusion >>
rect 141 175 142 176 
<< pdiffusion >>
rect 142 175 143 176 
<< pdiffusion >>
rect 143 175 144 176 
<< m1 >>
rect 145 175 146 176 
<< pdiffusion >>
rect 156 175 157 176 
<< pdiffusion >>
rect 157 175 158 176 
<< pdiffusion >>
rect 158 175 159 176 
<< pdiffusion >>
rect 159 175 160 176 
<< pdiffusion >>
rect 160 175 161 176 
<< pdiffusion >>
rect 161 175 162 176 
<< pdiffusion >>
rect 174 175 175 176 
<< pdiffusion >>
rect 175 175 176 176 
<< pdiffusion >>
rect 176 175 177 176 
<< pdiffusion >>
rect 177 175 178 176 
<< pdiffusion >>
rect 178 175 179 176 
<< pdiffusion >>
rect 179 175 180 176 
<< m1 >>
rect 181 175 182 176 
<< m1 >>
rect 183 175 184 176 
<< m1 >>
rect 185 175 186 176 
<< m2 >>
rect 189 175 190 176 
<< m1 >>
rect 190 175 191 176 
<< pdiffusion >>
rect 192 175 193 176 
<< pdiffusion >>
rect 193 175 194 176 
<< pdiffusion >>
rect 194 175 195 176 
<< pdiffusion >>
rect 195 175 196 176 
<< pdiffusion >>
rect 196 175 197 176 
<< pdiffusion >>
rect 197 175 198 176 
<< m1 >>
rect 199 175 200 176 
<< m2 >>
rect 199 175 200 176 
<< pdiffusion >>
rect 210 175 211 176 
<< pdiffusion >>
rect 211 175 212 176 
<< pdiffusion >>
rect 212 175 213 176 
<< pdiffusion >>
rect 213 175 214 176 
<< pdiffusion >>
rect 214 175 215 176 
<< pdiffusion >>
rect 215 175 216 176 
<< pdiffusion >>
rect 228 175 229 176 
<< pdiffusion >>
rect 229 175 230 176 
<< pdiffusion >>
rect 230 175 231 176 
<< pdiffusion >>
rect 231 175 232 176 
<< pdiffusion >>
rect 232 175 233 176 
<< pdiffusion >>
rect 233 175 234 176 
<< m1 >>
rect 254 175 255 176 
<< m1 >>
rect 256 175 257 176 
<< pdiffusion >>
rect 12 176 13 177 
<< pdiffusion >>
rect 13 176 14 177 
<< pdiffusion >>
rect 14 176 15 177 
<< pdiffusion >>
rect 15 176 16 177 
<< pdiffusion >>
rect 16 176 17 177 
<< pdiffusion >>
rect 17 176 18 177 
<< m1 >>
rect 19 176 20 177 
<< m1 >>
rect 28 176 29 177 
<< pdiffusion >>
rect 30 176 31 177 
<< pdiffusion >>
rect 31 176 32 177 
<< pdiffusion >>
rect 32 176 33 177 
<< pdiffusion >>
rect 33 176 34 177 
<< pdiffusion >>
rect 34 176 35 177 
<< pdiffusion >>
rect 35 176 36 177 
<< m1 >>
rect 44 176 45 177 
<< m1 >>
rect 46 176 47 177 
<< pdiffusion >>
rect 48 176 49 177 
<< pdiffusion >>
rect 49 176 50 177 
<< pdiffusion >>
rect 50 176 51 177 
<< pdiffusion >>
rect 51 176 52 177 
<< pdiffusion >>
rect 52 176 53 177 
<< pdiffusion >>
rect 53 176 54 177 
<< m1 >>
rect 55 176 56 177 
<< m2 >>
rect 56 176 57 177 
<< m1 >>
rect 59 176 60 177 
<< m1 >>
rect 64 176 65 177 
<< pdiffusion >>
rect 66 176 67 177 
<< pdiffusion >>
rect 67 176 68 177 
<< pdiffusion >>
rect 68 176 69 177 
<< pdiffusion >>
rect 69 176 70 177 
<< pdiffusion >>
rect 70 176 71 177 
<< pdiffusion >>
rect 71 176 72 177 
<< m1 >>
rect 73 176 74 177 
<< m1 >>
rect 75 176 76 177 
<< m1 >>
rect 82 176 83 177 
<< pdiffusion >>
rect 84 176 85 177 
<< pdiffusion >>
rect 85 176 86 177 
<< pdiffusion >>
rect 86 176 87 177 
<< pdiffusion >>
rect 87 176 88 177 
<< pdiffusion >>
rect 88 176 89 177 
<< pdiffusion >>
rect 89 176 90 177 
<< m1 >>
rect 91 176 92 177 
<< m1 >>
rect 93 176 94 177 
<< pdiffusion >>
rect 102 176 103 177 
<< pdiffusion >>
rect 103 176 104 177 
<< pdiffusion >>
rect 104 176 105 177 
<< pdiffusion >>
rect 105 176 106 177 
<< pdiffusion >>
rect 106 176 107 177 
<< pdiffusion >>
rect 107 176 108 177 
<< m1 >>
rect 109 176 110 177 
<< m1 >>
rect 111 176 112 177 
<< m1 >>
rect 113 176 114 177 
<< pdiffusion >>
rect 120 176 121 177 
<< pdiffusion >>
rect 121 176 122 177 
<< pdiffusion >>
rect 122 176 123 177 
<< pdiffusion >>
rect 123 176 124 177 
<< pdiffusion >>
rect 124 176 125 177 
<< pdiffusion >>
rect 125 176 126 177 
<< m1 >>
rect 127 176 128 177 
<< m1 >>
rect 129 176 130 177 
<< m1 >>
rect 136 176 137 177 
<< pdiffusion >>
rect 138 176 139 177 
<< pdiffusion >>
rect 139 176 140 177 
<< pdiffusion >>
rect 140 176 141 177 
<< pdiffusion >>
rect 141 176 142 177 
<< pdiffusion >>
rect 142 176 143 177 
<< pdiffusion >>
rect 143 176 144 177 
<< m1 >>
rect 145 176 146 177 
<< pdiffusion >>
rect 156 176 157 177 
<< pdiffusion >>
rect 157 176 158 177 
<< pdiffusion >>
rect 158 176 159 177 
<< pdiffusion >>
rect 159 176 160 177 
<< pdiffusion >>
rect 160 176 161 177 
<< pdiffusion >>
rect 161 176 162 177 
<< pdiffusion >>
rect 174 176 175 177 
<< pdiffusion >>
rect 175 176 176 177 
<< pdiffusion >>
rect 176 176 177 177 
<< pdiffusion >>
rect 177 176 178 177 
<< pdiffusion >>
rect 178 176 179 177 
<< pdiffusion >>
rect 179 176 180 177 
<< m1 >>
rect 181 176 182 177 
<< m1 >>
rect 183 176 184 177 
<< m1 >>
rect 185 176 186 177 
<< m2 >>
rect 189 176 190 177 
<< m1 >>
rect 190 176 191 177 
<< pdiffusion >>
rect 192 176 193 177 
<< pdiffusion >>
rect 193 176 194 177 
<< pdiffusion >>
rect 194 176 195 177 
<< pdiffusion >>
rect 195 176 196 177 
<< pdiffusion >>
rect 196 176 197 177 
<< pdiffusion >>
rect 197 176 198 177 
<< m1 >>
rect 199 176 200 177 
<< m2 >>
rect 199 176 200 177 
<< pdiffusion >>
rect 210 176 211 177 
<< pdiffusion >>
rect 211 176 212 177 
<< pdiffusion >>
rect 212 176 213 177 
<< pdiffusion >>
rect 213 176 214 177 
<< pdiffusion >>
rect 214 176 215 177 
<< pdiffusion >>
rect 215 176 216 177 
<< pdiffusion >>
rect 228 176 229 177 
<< pdiffusion >>
rect 229 176 230 177 
<< pdiffusion >>
rect 230 176 231 177 
<< pdiffusion >>
rect 231 176 232 177 
<< pdiffusion >>
rect 232 176 233 177 
<< pdiffusion >>
rect 233 176 234 177 
<< m1 >>
rect 254 176 255 177 
<< m1 >>
rect 256 176 257 177 
<< pdiffusion >>
rect 12 177 13 178 
<< pdiffusion >>
rect 13 177 14 178 
<< pdiffusion >>
rect 14 177 15 178 
<< pdiffusion >>
rect 15 177 16 178 
<< pdiffusion >>
rect 16 177 17 178 
<< pdiffusion >>
rect 17 177 18 178 
<< m1 >>
rect 19 177 20 178 
<< m1 >>
rect 28 177 29 178 
<< pdiffusion >>
rect 30 177 31 178 
<< pdiffusion >>
rect 31 177 32 178 
<< pdiffusion >>
rect 32 177 33 178 
<< pdiffusion >>
rect 33 177 34 178 
<< pdiffusion >>
rect 34 177 35 178 
<< pdiffusion >>
rect 35 177 36 178 
<< m1 >>
rect 44 177 45 178 
<< m1 >>
rect 46 177 47 178 
<< pdiffusion >>
rect 48 177 49 178 
<< pdiffusion >>
rect 49 177 50 178 
<< pdiffusion >>
rect 50 177 51 178 
<< pdiffusion >>
rect 51 177 52 178 
<< pdiffusion >>
rect 52 177 53 178 
<< pdiffusion >>
rect 53 177 54 178 
<< m1 >>
rect 55 177 56 178 
<< m2 >>
rect 56 177 57 178 
<< m1 >>
rect 59 177 60 178 
<< m1 >>
rect 64 177 65 178 
<< pdiffusion >>
rect 66 177 67 178 
<< pdiffusion >>
rect 67 177 68 178 
<< pdiffusion >>
rect 68 177 69 178 
<< pdiffusion >>
rect 69 177 70 178 
<< pdiffusion >>
rect 70 177 71 178 
<< pdiffusion >>
rect 71 177 72 178 
<< m1 >>
rect 73 177 74 178 
<< m1 >>
rect 75 177 76 178 
<< m1 >>
rect 82 177 83 178 
<< pdiffusion >>
rect 84 177 85 178 
<< pdiffusion >>
rect 85 177 86 178 
<< pdiffusion >>
rect 86 177 87 178 
<< pdiffusion >>
rect 87 177 88 178 
<< pdiffusion >>
rect 88 177 89 178 
<< pdiffusion >>
rect 89 177 90 178 
<< m1 >>
rect 91 177 92 178 
<< m1 >>
rect 93 177 94 178 
<< pdiffusion >>
rect 102 177 103 178 
<< pdiffusion >>
rect 103 177 104 178 
<< pdiffusion >>
rect 104 177 105 178 
<< pdiffusion >>
rect 105 177 106 178 
<< pdiffusion >>
rect 106 177 107 178 
<< pdiffusion >>
rect 107 177 108 178 
<< m1 >>
rect 109 177 110 178 
<< m1 >>
rect 111 177 112 178 
<< m1 >>
rect 113 177 114 178 
<< pdiffusion >>
rect 120 177 121 178 
<< pdiffusion >>
rect 121 177 122 178 
<< pdiffusion >>
rect 122 177 123 178 
<< pdiffusion >>
rect 123 177 124 178 
<< pdiffusion >>
rect 124 177 125 178 
<< pdiffusion >>
rect 125 177 126 178 
<< m1 >>
rect 127 177 128 178 
<< m1 >>
rect 129 177 130 178 
<< m1 >>
rect 136 177 137 178 
<< pdiffusion >>
rect 138 177 139 178 
<< pdiffusion >>
rect 139 177 140 178 
<< pdiffusion >>
rect 140 177 141 178 
<< pdiffusion >>
rect 141 177 142 178 
<< pdiffusion >>
rect 142 177 143 178 
<< pdiffusion >>
rect 143 177 144 178 
<< m1 >>
rect 145 177 146 178 
<< pdiffusion >>
rect 156 177 157 178 
<< pdiffusion >>
rect 157 177 158 178 
<< pdiffusion >>
rect 158 177 159 178 
<< pdiffusion >>
rect 159 177 160 178 
<< pdiffusion >>
rect 160 177 161 178 
<< pdiffusion >>
rect 161 177 162 178 
<< pdiffusion >>
rect 174 177 175 178 
<< pdiffusion >>
rect 175 177 176 178 
<< pdiffusion >>
rect 176 177 177 178 
<< pdiffusion >>
rect 177 177 178 178 
<< pdiffusion >>
rect 178 177 179 178 
<< pdiffusion >>
rect 179 177 180 178 
<< m1 >>
rect 181 177 182 178 
<< m1 >>
rect 183 177 184 178 
<< m1 >>
rect 185 177 186 178 
<< m2 >>
rect 189 177 190 178 
<< m1 >>
rect 190 177 191 178 
<< pdiffusion >>
rect 192 177 193 178 
<< pdiffusion >>
rect 193 177 194 178 
<< pdiffusion >>
rect 194 177 195 178 
<< pdiffusion >>
rect 195 177 196 178 
<< pdiffusion >>
rect 196 177 197 178 
<< pdiffusion >>
rect 197 177 198 178 
<< m1 >>
rect 199 177 200 178 
<< m2 >>
rect 199 177 200 178 
<< pdiffusion >>
rect 210 177 211 178 
<< pdiffusion >>
rect 211 177 212 178 
<< pdiffusion >>
rect 212 177 213 178 
<< pdiffusion >>
rect 213 177 214 178 
<< pdiffusion >>
rect 214 177 215 178 
<< pdiffusion >>
rect 215 177 216 178 
<< pdiffusion >>
rect 228 177 229 178 
<< pdiffusion >>
rect 229 177 230 178 
<< pdiffusion >>
rect 230 177 231 178 
<< pdiffusion >>
rect 231 177 232 178 
<< pdiffusion >>
rect 232 177 233 178 
<< pdiffusion >>
rect 233 177 234 178 
<< m1 >>
rect 254 177 255 178 
<< m1 >>
rect 256 177 257 178 
<< pdiffusion >>
rect 12 178 13 179 
<< pdiffusion >>
rect 13 178 14 179 
<< pdiffusion >>
rect 14 178 15 179 
<< pdiffusion >>
rect 15 178 16 179 
<< pdiffusion >>
rect 16 178 17 179 
<< pdiffusion >>
rect 17 178 18 179 
<< m1 >>
rect 19 178 20 179 
<< m1 >>
rect 28 178 29 179 
<< pdiffusion >>
rect 30 178 31 179 
<< pdiffusion >>
rect 31 178 32 179 
<< pdiffusion >>
rect 32 178 33 179 
<< pdiffusion >>
rect 33 178 34 179 
<< pdiffusion >>
rect 34 178 35 179 
<< pdiffusion >>
rect 35 178 36 179 
<< m1 >>
rect 44 178 45 179 
<< m1 >>
rect 46 178 47 179 
<< pdiffusion >>
rect 48 178 49 179 
<< pdiffusion >>
rect 49 178 50 179 
<< pdiffusion >>
rect 50 178 51 179 
<< pdiffusion >>
rect 51 178 52 179 
<< pdiffusion >>
rect 52 178 53 179 
<< pdiffusion >>
rect 53 178 54 179 
<< m1 >>
rect 55 178 56 179 
<< m2 >>
rect 56 178 57 179 
<< m1 >>
rect 59 178 60 179 
<< m2 >>
rect 59 178 60 179 
<< m2c >>
rect 59 178 60 179 
<< m1 >>
rect 59 178 60 179 
<< m2 >>
rect 59 178 60 179 
<< m1 >>
rect 64 178 65 179 
<< pdiffusion >>
rect 66 178 67 179 
<< pdiffusion >>
rect 67 178 68 179 
<< pdiffusion >>
rect 68 178 69 179 
<< pdiffusion >>
rect 69 178 70 179 
<< pdiffusion >>
rect 70 178 71 179 
<< pdiffusion >>
rect 71 178 72 179 
<< m1 >>
rect 73 178 74 179 
<< m1 >>
rect 75 178 76 179 
<< m1 >>
rect 82 178 83 179 
<< pdiffusion >>
rect 84 178 85 179 
<< pdiffusion >>
rect 85 178 86 179 
<< pdiffusion >>
rect 86 178 87 179 
<< pdiffusion >>
rect 87 178 88 179 
<< pdiffusion >>
rect 88 178 89 179 
<< pdiffusion >>
rect 89 178 90 179 
<< m1 >>
rect 91 178 92 179 
<< m1 >>
rect 93 178 94 179 
<< pdiffusion >>
rect 102 178 103 179 
<< pdiffusion >>
rect 103 178 104 179 
<< pdiffusion >>
rect 104 178 105 179 
<< pdiffusion >>
rect 105 178 106 179 
<< pdiffusion >>
rect 106 178 107 179 
<< pdiffusion >>
rect 107 178 108 179 
<< m1 >>
rect 109 178 110 179 
<< m1 >>
rect 111 178 112 179 
<< m1 >>
rect 113 178 114 179 
<< pdiffusion >>
rect 120 178 121 179 
<< pdiffusion >>
rect 121 178 122 179 
<< pdiffusion >>
rect 122 178 123 179 
<< pdiffusion >>
rect 123 178 124 179 
<< pdiffusion >>
rect 124 178 125 179 
<< pdiffusion >>
rect 125 178 126 179 
<< m1 >>
rect 127 178 128 179 
<< m1 >>
rect 129 178 130 179 
<< m1 >>
rect 136 178 137 179 
<< pdiffusion >>
rect 138 178 139 179 
<< pdiffusion >>
rect 139 178 140 179 
<< pdiffusion >>
rect 140 178 141 179 
<< pdiffusion >>
rect 141 178 142 179 
<< pdiffusion >>
rect 142 178 143 179 
<< pdiffusion >>
rect 143 178 144 179 
<< m1 >>
rect 145 178 146 179 
<< pdiffusion >>
rect 156 178 157 179 
<< pdiffusion >>
rect 157 178 158 179 
<< pdiffusion >>
rect 158 178 159 179 
<< pdiffusion >>
rect 159 178 160 179 
<< pdiffusion >>
rect 160 178 161 179 
<< pdiffusion >>
rect 161 178 162 179 
<< pdiffusion >>
rect 174 178 175 179 
<< pdiffusion >>
rect 175 178 176 179 
<< pdiffusion >>
rect 176 178 177 179 
<< pdiffusion >>
rect 177 178 178 179 
<< pdiffusion >>
rect 178 178 179 179 
<< pdiffusion >>
rect 179 178 180 179 
<< m1 >>
rect 181 178 182 179 
<< m1 >>
rect 183 178 184 179 
<< m1 >>
rect 185 178 186 179 
<< m2 >>
rect 189 178 190 179 
<< m1 >>
rect 190 178 191 179 
<< pdiffusion >>
rect 192 178 193 179 
<< pdiffusion >>
rect 193 178 194 179 
<< pdiffusion >>
rect 194 178 195 179 
<< pdiffusion >>
rect 195 178 196 179 
<< pdiffusion >>
rect 196 178 197 179 
<< pdiffusion >>
rect 197 178 198 179 
<< m1 >>
rect 199 178 200 179 
<< m2 >>
rect 199 178 200 179 
<< pdiffusion >>
rect 210 178 211 179 
<< pdiffusion >>
rect 211 178 212 179 
<< pdiffusion >>
rect 212 178 213 179 
<< pdiffusion >>
rect 213 178 214 179 
<< pdiffusion >>
rect 214 178 215 179 
<< pdiffusion >>
rect 215 178 216 179 
<< pdiffusion >>
rect 228 178 229 179 
<< pdiffusion >>
rect 229 178 230 179 
<< pdiffusion >>
rect 230 178 231 179 
<< pdiffusion >>
rect 231 178 232 179 
<< pdiffusion >>
rect 232 178 233 179 
<< pdiffusion >>
rect 233 178 234 179 
<< m1 >>
rect 254 178 255 179 
<< m1 >>
rect 256 178 257 179 
<< pdiffusion >>
rect 12 179 13 180 
<< pdiffusion >>
rect 13 179 14 180 
<< pdiffusion >>
rect 14 179 15 180 
<< pdiffusion >>
rect 15 179 16 180 
<< pdiffusion >>
rect 16 179 17 180 
<< pdiffusion >>
rect 17 179 18 180 
<< m1 >>
rect 19 179 20 180 
<< m1 >>
rect 28 179 29 180 
<< pdiffusion >>
rect 30 179 31 180 
<< m1 >>
rect 31 179 32 180 
<< pdiffusion >>
rect 31 179 32 180 
<< pdiffusion >>
rect 32 179 33 180 
<< pdiffusion >>
rect 33 179 34 180 
<< pdiffusion >>
rect 34 179 35 180 
<< pdiffusion >>
rect 35 179 36 180 
<< m1 >>
rect 44 179 45 180 
<< m1 >>
rect 46 179 47 180 
<< pdiffusion >>
rect 48 179 49 180 
<< pdiffusion >>
rect 49 179 50 180 
<< pdiffusion >>
rect 50 179 51 180 
<< pdiffusion >>
rect 51 179 52 180 
<< m1 >>
rect 52 179 53 180 
<< pdiffusion >>
rect 52 179 53 180 
<< pdiffusion >>
rect 53 179 54 180 
<< m1 >>
rect 55 179 56 180 
<< m2 >>
rect 56 179 57 180 
<< m2 >>
rect 59 179 60 180 
<< m1 >>
rect 64 179 65 180 
<< pdiffusion >>
rect 66 179 67 180 
<< m1 >>
rect 67 179 68 180 
<< pdiffusion >>
rect 67 179 68 180 
<< pdiffusion >>
rect 68 179 69 180 
<< pdiffusion >>
rect 69 179 70 180 
<< m1 >>
rect 70 179 71 180 
<< pdiffusion >>
rect 70 179 71 180 
<< pdiffusion >>
rect 71 179 72 180 
<< m1 >>
rect 73 179 74 180 
<< m1 >>
rect 75 179 76 180 
<< m1 >>
rect 82 179 83 180 
<< pdiffusion >>
rect 84 179 85 180 
<< pdiffusion >>
rect 85 179 86 180 
<< pdiffusion >>
rect 86 179 87 180 
<< pdiffusion >>
rect 87 179 88 180 
<< pdiffusion >>
rect 88 179 89 180 
<< pdiffusion >>
rect 89 179 90 180 
<< m1 >>
rect 91 179 92 180 
<< m1 >>
rect 93 179 94 180 
<< pdiffusion >>
rect 102 179 103 180 
<< pdiffusion >>
rect 103 179 104 180 
<< pdiffusion >>
rect 104 179 105 180 
<< pdiffusion >>
rect 105 179 106 180 
<< pdiffusion >>
rect 106 179 107 180 
<< pdiffusion >>
rect 107 179 108 180 
<< m1 >>
rect 109 179 110 180 
<< m1 >>
rect 111 179 112 180 
<< m1 >>
rect 113 179 114 180 
<< pdiffusion >>
rect 120 179 121 180 
<< pdiffusion >>
rect 121 179 122 180 
<< pdiffusion >>
rect 122 179 123 180 
<< pdiffusion >>
rect 123 179 124 180 
<< pdiffusion >>
rect 124 179 125 180 
<< pdiffusion >>
rect 125 179 126 180 
<< m1 >>
rect 127 179 128 180 
<< m1 >>
rect 129 179 130 180 
<< m1 >>
rect 136 179 137 180 
<< pdiffusion >>
rect 138 179 139 180 
<< pdiffusion >>
rect 139 179 140 180 
<< pdiffusion >>
rect 140 179 141 180 
<< pdiffusion >>
rect 141 179 142 180 
<< m1 >>
rect 142 179 143 180 
<< pdiffusion >>
rect 142 179 143 180 
<< pdiffusion >>
rect 143 179 144 180 
<< m1 >>
rect 145 179 146 180 
<< pdiffusion >>
rect 156 179 157 180 
<< pdiffusion >>
rect 157 179 158 180 
<< pdiffusion >>
rect 158 179 159 180 
<< pdiffusion >>
rect 159 179 160 180 
<< pdiffusion >>
rect 160 179 161 180 
<< pdiffusion >>
rect 161 179 162 180 
<< pdiffusion >>
rect 174 179 175 180 
<< pdiffusion >>
rect 175 179 176 180 
<< pdiffusion >>
rect 176 179 177 180 
<< pdiffusion >>
rect 177 179 178 180 
<< pdiffusion >>
rect 178 179 179 180 
<< pdiffusion >>
rect 179 179 180 180 
<< m1 >>
rect 181 179 182 180 
<< m1 >>
rect 183 179 184 180 
<< m1 >>
rect 185 179 186 180 
<< m2 >>
rect 189 179 190 180 
<< m1 >>
rect 190 179 191 180 
<< pdiffusion >>
rect 192 179 193 180 
<< m1 >>
rect 193 179 194 180 
<< pdiffusion >>
rect 193 179 194 180 
<< pdiffusion >>
rect 194 179 195 180 
<< pdiffusion >>
rect 195 179 196 180 
<< m1 >>
rect 196 179 197 180 
<< pdiffusion >>
rect 196 179 197 180 
<< pdiffusion >>
rect 197 179 198 180 
<< m1 >>
rect 199 179 200 180 
<< m2 >>
rect 199 179 200 180 
<< pdiffusion >>
rect 210 179 211 180 
<< pdiffusion >>
rect 211 179 212 180 
<< pdiffusion >>
rect 212 179 213 180 
<< pdiffusion >>
rect 213 179 214 180 
<< pdiffusion >>
rect 214 179 215 180 
<< pdiffusion >>
rect 215 179 216 180 
<< pdiffusion >>
rect 228 179 229 180 
<< m1 >>
rect 229 179 230 180 
<< pdiffusion >>
rect 229 179 230 180 
<< pdiffusion >>
rect 230 179 231 180 
<< pdiffusion >>
rect 231 179 232 180 
<< pdiffusion >>
rect 232 179 233 180 
<< pdiffusion >>
rect 233 179 234 180 
<< m1 >>
rect 254 179 255 180 
<< m1 >>
rect 256 179 257 180 
<< m1 >>
rect 19 180 20 181 
<< m1 >>
rect 28 180 29 181 
<< m1 >>
rect 31 180 32 181 
<< m1 >>
rect 44 180 45 181 
<< m1 >>
rect 46 180 47 181 
<< m1 >>
rect 52 180 53 181 
<< m1 >>
rect 55 180 56 181 
<< m2 >>
rect 56 180 57 181 
<< m1 >>
rect 57 180 58 181 
<< m2 >>
rect 57 180 58 181 
<< m2c >>
rect 57 180 58 181 
<< m1 >>
rect 57 180 58 181 
<< m2 >>
rect 57 180 58 181 
<< m1 >>
rect 58 180 59 181 
<< m1 >>
rect 59 180 60 181 
<< m2 >>
rect 59 180 60 181 
<< m1 >>
rect 60 180 61 181 
<< m1 >>
rect 61 180 62 181 
<< m1 >>
rect 62 180 63 181 
<< m1 >>
rect 64 180 65 181 
<< m1 >>
rect 67 180 68 181 
<< m1 >>
rect 70 180 71 181 
<< m1 >>
rect 73 180 74 181 
<< m1 >>
rect 75 180 76 181 
<< m1 >>
rect 82 180 83 181 
<< m1 >>
rect 91 180 92 181 
<< m1 >>
rect 93 180 94 181 
<< m1 >>
rect 109 180 110 181 
<< m1 >>
rect 111 180 112 181 
<< m1 >>
rect 113 180 114 181 
<< m1 >>
rect 127 180 128 181 
<< m1 >>
rect 129 180 130 181 
<< m1 >>
rect 136 180 137 181 
<< m1 >>
rect 142 180 143 181 
<< m1 >>
rect 145 180 146 181 
<< m1 >>
rect 181 180 182 181 
<< m1 >>
rect 183 180 184 181 
<< m1 >>
rect 185 180 186 181 
<< m2 >>
rect 189 180 190 181 
<< m1 >>
rect 190 180 191 181 
<< m1 >>
rect 193 180 194 181 
<< m1 >>
rect 196 180 197 181 
<< m1 >>
rect 199 180 200 181 
<< m2 >>
rect 199 180 200 181 
<< m1 >>
rect 229 180 230 181 
<< m1 >>
rect 254 180 255 181 
<< m1 >>
rect 256 180 257 181 
<< m1 >>
rect 19 181 20 182 
<< m1 >>
rect 28 181 29 182 
<< m1 >>
rect 31 181 32 182 
<< m1 >>
rect 44 181 45 182 
<< m1 >>
rect 46 181 47 182 
<< m1 >>
rect 52 181 53 182 
<< m1 >>
rect 55 181 56 182 
<< m2 >>
rect 59 181 60 182 
<< m1 >>
rect 62 181 63 182 
<< m1 >>
rect 64 181 65 182 
<< m1 >>
rect 67 181 68 182 
<< m1 >>
rect 68 181 69 182 
<< m2 >>
rect 68 181 69 182 
<< m2c >>
rect 68 181 69 182 
<< m1 >>
rect 68 181 69 182 
<< m2 >>
rect 68 181 69 182 
<< m2 >>
rect 69 181 70 182 
<< m1 >>
rect 70 181 71 182 
<< m1 >>
rect 73 181 74 182 
<< m1 >>
rect 75 181 76 182 
<< m1 >>
rect 82 181 83 182 
<< m1 >>
rect 91 181 92 182 
<< m1 >>
rect 93 181 94 182 
<< m1 >>
rect 109 181 110 182 
<< m1 >>
rect 111 181 112 182 
<< m1 >>
rect 113 181 114 182 
<< m1 >>
rect 127 181 128 182 
<< m1 >>
rect 129 181 130 182 
<< m1 >>
rect 136 181 137 182 
<< m1 >>
rect 142 181 143 182 
<< m1 >>
rect 145 181 146 182 
<< m1 >>
rect 181 181 182 182 
<< m1 >>
rect 183 181 184 182 
<< m1 >>
rect 185 181 186 182 
<< m2 >>
rect 189 181 190 182 
<< m1 >>
rect 190 181 191 182 
<< m1 >>
rect 193 181 194 182 
<< m1 >>
rect 194 181 195 182 
<< m2 >>
rect 194 181 195 182 
<< m2c >>
rect 194 181 195 182 
<< m1 >>
rect 194 181 195 182 
<< m2 >>
rect 194 181 195 182 
<< m2 >>
rect 195 181 196 182 
<< m1 >>
rect 196 181 197 182 
<< m1 >>
rect 197 181 198 182 
<< m1 >>
rect 198 181 199 182 
<< m1 >>
rect 199 181 200 182 
<< m2 >>
rect 199 181 200 182 
<< m1 >>
rect 229 181 230 182 
<< m1 >>
rect 254 181 255 182 
<< m1 >>
rect 256 181 257 182 
<< m1 >>
rect 19 182 20 183 
<< m1 >>
rect 28 182 29 183 
<< m2 >>
rect 28 182 29 183 
<< m2c >>
rect 28 182 29 183 
<< m1 >>
rect 28 182 29 183 
<< m2 >>
rect 28 182 29 183 
<< m1 >>
rect 31 182 32 183 
<< m1 >>
rect 32 182 33 183 
<< m1 >>
rect 33 182 34 183 
<< m1 >>
rect 34 182 35 183 
<< m1 >>
rect 35 182 36 183 
<< m1 >>
rect 36 182 37 183 
<< m1 >>
rect 37 182 38 183 
<< m1 >>
rect 38 182 39 183 
<< m1 >>
rect 39 182 40 183 
<< m1 >>
rect 40 182 41 183 
<< m1 >>
rect 41 182 42 183 
<< m1 >>
rect 42 182 43 183 
<< m1 >>
rect 43 182 44 183 
<< m1 >>
rect 44 182 45 183 
<< m1 >>
rect 46 182 47 183 
<< m2 >>
rect 46 182 47 183 
<< m2c >>
rect 46 182 47 183 
<< m1 >>
rect 46 182 47 183 
<< m2 >>
rect 46 182 47 183 
<< m1 >>
rect 52 182 53 183 
<< m2 >>
rect 52 182 53 183 
<< m2c >>
rect 52 182 53 183 
<< m1 >>
rect 52 182 53 183 
<< m2 >>
rect 52 182 53 183 
<< m1 >>
rect 55 182 56 183 
<< m2 >>
rect 55 182 56 183 
<< m2c >>
rect 55 182 56 183 
<< m1 >>
rect 55 182 56 183 
<< m2 >>
rect 55 182 56 183 
<< m1 >>
rect 59 182 60 183 
<< m2 >>
rect 59 182 60 183 
<< m2c >>
rect 59 182 60 183 
<< m1 >>
rect 59 182 60 183 
<< m2 >>
rect 59 182 60 183 
<< m1 >>
rect 62 182 63 183 
<< m2 >>
rect 62 182 63 183 
<< m2c >>
rect 62 182 63 183 
<< m1 >>
rect 62 182 63 183 
<< m2 >>
rect 62 182 63 183 
<< m1 >>
rect 64 182 65 183 
<< m2 >>
rect 64 182 65 183 
<< m2c >>
rect 64 182 65 183 
<< m1 >>
rect 64 182 65 183 
<< m2 >>
rect 64 182 65 183 
<< m2 >>
rect 69 182 70 183 
<< m1 >>
rect 70 182 71 183 
<< m2 >>
rect 70 182 71 183 
<< m2 >>
rect 71 182 72 183 
<< m2 >>
rect 72 182 73 183 
<< m1 >>
rect 73 182 74 183 
<< m2 >>
rect 73 182 74 183 
<< m2 >>
rect 74 182 75 183 
<< m1 >>
rect 75 182 76 183 
<< m2 >>
rect 75 182 76 183 
<< m2c >>
rect 75 182 76 183 
<< m1 >>
rect 75 182 76 183 
<< m2 >>
rect 75 182 76 183 
<< m1 >>
rect 82 182 83 183 
<< m1 >>
rect 86 182 87 183 
<< m1 >>
rect 87 182 88 183 
<< m1 >>
rect 88 182 89 183 
<< m1 >>
rect 89 182 90 183 
<< m2 >>
rect 89 182 90 183 
<< m2c >>
rect 89 182 90 183 
<< m1 >>
rect 89 182 90 183 
<< m2 >>
rect 89 182 90 183 
<< m2 >>
rect 90 182 91 183 
<< m1 >>
rect 91 182 92 183 
<< m2 >>
rect 91 182 92 183 
<< m2 >>
rect 92 182 93 183 
<< m1 >>
rect 93 182 94 183 
<< m2 >>
rect 93 182 94 183 
<< m2c >>
rect 93 182 94 183 
<< m1 >>
rect 93 182 94 183 
<< m2 >>
rect 93 182 94 183 
<< m2 >>
rect 108 182 109 183 
<< m1 >>
rect 109 182 110 183 
<< m2 >>
rect 109 182 110 183 
<< m2 >>
rect 110 182 111 183 
<< m1 >>
rect 111 182 112 183 
<< m2 >>
rect 111 182 112 183 
<< m2c >>
rect 111 182 112 183 
<< m1 >>
rect 111 182 112 183 
<< m2 >>
rect 111 182 112 183 
<< m1 >>
rect 113 182 114 183 
<< m2 >>
rect 113 182 114 183 
<< m2c >>
rect 113 182 114 183 
<< m1 >>
rect 113 182 114 183 
<< m2 >>
rect 113 182 114 183 
<< m1 >>
rect 127 182 128 183 
<< m2 >>
rect 127 182 128 183 
<< m2c >>
rect 127 182 128 183 
<< m1 >>
rect 127 182 128 183 
<< m2 >>
rect 127 182 128 183 
<< m1 >>
rect 129 182 130 183 
<< m2 >>
rect 129 182 130 183 
<< m2c >>
rect 129 182 130 183 
<< m1 >>
rect 129 182 130 183 
<< m2 >>
rect 129 182 130 183 
<< m1 >>
rect 136 182 137 183 
<< m1 >>
rect 137 182 138 183 
<< m1 >>
rect 138 182 139 183 
<< m2 >>
rect 138 182 139 183 
<< m2c >>
rect 138 182 139 183 
<< m1 >>
rect 138 182 139 183 
<< m2 >>
rect 138 182 139 183 
<< m1 >>
rect 142 182 143 183 
<< m2 >>
rect 142 182 143 183 
<< m2c >>
rect 142 182 143 183 
<< m1 >>
rect 142 182 143 183 
<< m2 >>
rect 142 182 143 183 
<< m1 >>
rect 145 182 146 183 
<< m2 >>
rect 145 182 146 183 
<< m2c >>
rect 145 182 146 183 
<< m1 >>
rect 145 182 146 183 
<< m2 >>
rect 145 182 146 183 
<< m1 >>
rect 181 182 182 183 
<< m2 >>
rect 181 182 182 183 
<< m2c >>
rect 181 182 182 183 
<< m1 >>
rect 181 182 182 183 
<< m2 >>
rect 181 182 182 183 
<< m1 >>
rect 183 182 184 183 
<< m2 >>
rect 183 182 184 183 
<< m2c >>
rect 183 182 184 183 
<< m1 >>
rect 183 182 184 183 
<< m2 >>
rect 183 182 184 183 
<< m1 >>
rect 185 182 186 183 
<< m2 >>
rect 185 182 186 183 
<< m2c >>
rect 185 182 186 183 
<< m1 >>
rect 185 182 186 183 
<< m2 >>
rect 185 182 186 183 
<< m2 >>
rect 189 182 190 183 
<< m1 >>
rect 190 182 191 183 
<< m1 >>
rect 191 182 192 183 
<< m2 >>
rect 191 182 192 183 
<< m2c >>
rect 191 182 192 183 
<< m1 >>
rect 191 182 192 183 
<< m2 >>
rect 191 182 192 183 
<< m2 >>
rect 192 182 193 183 
<< m2 >>
rect 195 182 196 183 
<< m2 >>
rect 196 182 197 183 
<< m2 >>
rect 197 182 198 183 
<< m2 >>
rect 198 182 199 183 
<< m2 >>
rect 199 182 200 183 
<< m1 >>
rect 229 182 230 183 
<< m1 >>
rect 254 182 255 183 
<< m1 >>
rect 256 182 257 183 
<< m1 >>
rect 19 183 20 184 
<< m2 >>
rect 28 183 29 184 
<< m2 >>
rect 46 183 47 184 
<< m2 >>
rect 52 183 53 184 
<< m2 >>
rect 55 183 56 184 
<< m2 >>
rect 59 183 60 184 
<< m2 >>
rect 62 183 63 184 
<< m2 >>
rect 64 183 65 184 
<< m1 >>
rect 70 183 71 184 
<< m1 >>
rect 73 183 74 184 
<< m1 >>
rect 82 183 83 184 
<< m1 >>
rect 86 183 87 184 
<< m1 >>
rect 91 183 92 184 
<< m2 >>
rect 108 183 109 184 
<< m1 >>
rect 109 183 110 184 
<< m2 >>
rect 113 183 114 184 
<< m2 >>
rect 127 183 128 184 
<< m2 >>
rect 129 183 130 184 
<< m2 >>
rect 138 183 139 184 
<< m2 >>
rect 142 183 143 184 
<< m2 >>
rect 145 183 146 184 
<< m2 >>
rect 181 183 182 184 
<< m2 >>
rect 183 183 184 184 
<< m2 >>
rect 185 183 186 184 
<< m2 >>
rect 189 183 190 184 
<< m2 >>
rect 192 183 193 184 
<< m1 >>
rect 229 183 230 184 
<< m1 >>
rect 254 183 255 184 
<< m1 >>
rect 256 183 257 184 
<< m1 >>
rect 19 184 20 185 
<< m1 >>
rect 28 184 29 185 
<< m2 >>
rect 28 184 29 185 
<< m1 >>
rect 29 184 30 185 
<< m1 >>
rect 30 184 31 185 
<< m1 >>
rect 31 184 32 185 
<< m1 >>
rect 32 184 33 185 
<< m1 >>
rect 33 184 34 185 
<< m1 >>
rect 34 184 35 185 
<< m1 >>
rect 35 184 36 185 
<< m1 >>
rect 36 184 37 185 
<< m1 >>
rect 37 184 38 185 
<< m1 >>
rect 38 184 39 185 
<< m1 >>
rect 39 184 40 185 
<< m1 >>
rect 40 184 41 185 
<< m1 >>
rect 41 184 42 185 
<< m1 >>
rect 42 184 43 185 
<< m1 >>
rect 43 184 44 185 
<< m1 >>
rect 44 184 45 185 
<< m1 >>
rect 45 184 46 185 
<< m1 >>
rect 46 184 47 185 
<< m2 >>
rect 46 184 47 185 
<< m1 >>
rect 47 184 48 185 
<< m1 >>
rect 48 184 49 185 
<< m1 >>
rect 49 184 50 185 
<< m1 >>
rect 50 184 51 185 
<< m1 >>
rect 51 184 52 185 
<< m1 >>
rect 52 184 53 185 
<< m2 >>
rect 52 184 53 185 
<< m1 >>
rect 53 184 54 185 
<< m1 >>
rect 54 184 55 185 
<< m1 >>
rect 55 184 56 185 
<< m2 >>
rect 55 184 56 185 
<< m1 >>
rect 56 184 57 185 
<< m1 >>
rect 57 184 58 185 
<< m1 >>
rect 58 184 59 185 
<< m1 >>
rect 59 184 60 185 
<< m2 >>
rect 59 184 60 185 
<< m1 >>
rect 60 184 61 185 
<< m1 >>
rect 61 184 62 185 
<< m1 >>
rect 62 184 63 185 
<< m2 >>
rect 62 184 63 185 
<< m1 >>
rect 63 184 64 185 
<< m1 >>
rect 64 184 65 185 
<< m2 >>
rect 64 184 65 185 
<< m1 >>
rect 65 184 66 185 
<< m1 >>
rect 66 184 67 185 
<< m1 >>
rect 67 184 68 185 
<< m1 >>
rect 68 184 69 185 
<< m1 >>
rect 69 184 70 185 
<< m1 >>
rect 70 184 71 185 
<< m1 >>
rect 73 184 74 185 
<< m2 >>
rect 73 184 74 185 
<< m2c >>
rect 73 184 74 185 
<< m1 >>
rect 73 184 74 185 
<< m2 >>
rect 73 184 74 185 
<< m1 >>
rect 82 184 83 185 
<< m1 >>
rect 83 184 84 185 
<< m1 >>
rect 84 184 85 185 
<< m1 >>
rect 85 184 86 185 
<< m1 >>
rect 86 184 87 185 
<< m1 >>
rect 91 184 92 185 
<< m2 >>
rect 91 184 92 185 
<< m2c >>
rect 91 184 92 185 
<< m1 >>
rect 91 184 92 185 
<< m2 >>
rect 91 184 92 185 
<< m2 >>
rect 108 184 109 185 
<< m1 >>
rect 109 184 110 185 
<< m1 >>
rect 110 184 111 185 
<< m1 >>
rect 111 184 112 185 
<< m1 >>
rect 112 184 113 185 
<< m1 >>
rect 113 184 114 185 
<< m2 >>
rect 113 184 114 185 
<< m1 >>
rect 114 184 115 185 
<< m1 >>
rect 115 184 116 185 
<< m1 >>
rect 116 184 117 185 
<< m1 >>
rect 117 184 118 185 
<< m1 >>
rect 118 184 119 185 
<< m1 >>
rect 119 184 120 185 
<< m1 >>
rect 120 184 121 185 
<< m1 >>
rect 121 184 122 185 
<< m1 >>
rect 122 184 123 185 
<< m1 >>
rect 123 184 124 185 
<< m1 >>
rect 124 184 125 185 
<< m1 >>
rect 125 184 126 185 
<< m1 >>
rect 126 184 127 185 
<< m1 >>
rect 127 184 128 185 
<< m2 >>
rect 127 184 128 185 
<< m1 >>
rect 128 184 129 185 
<< m1 >>
rect 129 184 130 185 
<< m2 >>
rect 129 184 130 185 
<< m1 >>
rect 130 184 131 185 
<< m1 >>
rect 131 184 132 185 
<< m1 >>
rect 132 184 133 185 
<< m1 >>
rect 133 184 134 185 
<< m1 >>
rect 134 184 135 185 
<< m1 >>
rect 135 184 136 185 
<< m1 >>
rect 136 184 137 185 
<< m1 >>
rect 137 184 138 185 
<< m1 >>
rect 138 184 139 185 
<< m2 >>
rect 138 184 139 185 
<< m1 >>
rect 139 184 140 185 
<< m1 >>
rect 140 184 141 185 
<< m1 >>
rect 141 184 142 185 
<< m1 >>
rect 142 184 143 185 
<< m2 >>
rect 142 184 143 185 
<< m1 >>
rect 143 184 144 185 
<< m1 >>
rect 144 184 145 185 
<< m1 >>
rect 145 184 146 185 
<< m2 >>
rect 145 184 146 185 
<< m1 >>
rect 146 184 147 185 
<< m2 >>
rect 146 184 147 185 
<< m1 >>
rect 147 184 148 185 
<< m2 >>
rect 147 184 148 185 
<< m1 >>
rect 148 184 149 185 
<< m2 >>
rect 148 184 149 185 
<< m1 >>
rect 149 184 150 185 
<< m2 >>
rect 149 184 150 185 
<< m1 >>
rect 150 184 151 185 
<< m2 >>
rect 150 184 151 185 
<< m1 >>
rect 151 184 152 185 
<< m2 >>
rect 151 184 152 185 
<< m1 >>
rect 152 184 153 185 
<< m2 >>
rect 152 184 153 185 
<< m1 >>
rect 153 184 154 185 
<< m2 >>
rect 153 184 154 185 
<< m1 >>
rect 154 184 155 185 
<< m2 >>
rect 154 184 155 185 
<< m1 >>
rect 155 184 156 185 
<< m2 >>
rect 155 184 156 185 
<< m1 >>
rect 156 184 157 185 
<< m2 >>
rect 156 184 157 185 
<< m1 >>
rect 157 184 158 185 
<< m2 >>
rect 157 184 158 185 
<< m1 >>
rect 158 184 159 185 
<< m2 >>
rect 158 184 159 185 
<< m1 >>
rect 159 184 160 185 
<< m2 >>
rect 159 184 160 185 
<< m1 >>
rect 160 184 161 185 
<< m2 >>
rect 160 184 161 185 
<< m1 >>
rect 161 184 162 185 
<< m2 >>
rect 161 184 162 185 
<< m1 >>
rect 162 184 163 185 
<< m2 >>
rect 162 184 163 185 
<< m1 >>
rect 163 184 164 185 
<< m2 >>
rect 163 184 164 185 
<< m1 >>
rect 164 184 165 185 
<< m2 >>
rect 164 184 165 185 
<< m1 >>
rect 165 184 166 185 
<< m2 >>
rect 165 184 166 185 
<< m1 >>
rect 166 184 167 185 
<< m2 >>
rect 166 184 167 185 
<< m1 >>
rect 167 184 168 185 
<< m2 >>
rect 167 184 168 185 
<< m1 >>
rect 168 184 169 185 
<< m2 >>
rect 168 184 169 185 
<< m1 >>
rect 169 184 170 185 
<< m2 >>
rect 169 184 170 185 
<< m1 >>
rect 170 184 171 185 
<< m2 >>
rect 170 184 171 185 
<< m1 >>
rect 171 184 172 185 
<< m2 >>
rect 171 184 172 185 
<< m1 >>
rect 172 184 173 185 
<< m2 >>
rect 172 184 173 185 
<< m1 >>
rect 173 184 174 185 
<< m2 >>
rect 173 184 174 185 
<< m1 >>
rect 174 184 175 185 
<< m2 >>
rect 174 184 175 185 
<< m1 >>
rect 175 184 176 185 
<< m2 >>
rect 175 184 176 185 
<< m2 >>
rect 176 184 177 185 
<< m1 >>
rect 177 184 178 185 
<< m2 >>
rect 177 184 178 185 
<< m2c >>
rect 177 184 178 185 
<< m1 >>
rect 177 184 178 185 
<< m2 >>
rect 177 184 178 185 
<< m1 >>
rect 178 184 179 185 
<< m1 >>
rect 179 184 180 185 
<< m1 >>
rect 180 184 181 185 
<< m1 >>
rect 181 184 182 185 
<< m2 >>
rect 181 184 182 185 
<< m1 >>
rect 182 184 183 185 
<< m1 >>
rect 183 184 184 185 
<< m2 >>
rect 183 184 184 185 
<< m1 >>
rect 184 184 185 185 
<< m1 >>
rect 185 184 186 185 
<< m2 >>
rect 185 184 186 185 
<< m1 >>
rect 186 184 187 185 
<< m1 >>
rect 187 184 188 185 
<< m1 >>
rect 188 184 189 185 
<< m1 >>
rect 189 184 190 185 
<< m2 >>
rect 189 184 190 185 
<< m1 >>
rect 190 184 191 185 
<< m1 >>
rect 191 184 192 185 
<< m1 >>
rect 192 184 193 185 
<< m2 >>
rect 192 184 193 185 
<< m1 >>
rect 193 184 194 185 
<< m1 >>
rect 194 184 195 185 
<< m1 >>
rect 195 184 196 185 
<< m1 >>
rect 196 184 197 185 
<< m1 >>
rect 197 184 198 185 
<< m1 >>
rect 198 184 199 185 
<< m1 >>
rect 199 184 200 185 
<< m1 >>
rect 200 184 201 185 
<< m1 >>
rect 201 184 202 185 
<< m1 >>
rect 202 184 203 185 
<< m1 >>
rect 203 184 204 185 
<< m1 >>
rect 204 184 205 185 
<< m1 >>
rect 205 184 206 185 
<< m1 >>
rect 206 184 207 185 
<< m1 >>
rect 207 184 208 185 
<< m1 >>
rect 208 184 209 185 
<< m1 >>
rect 209 184 210 185 
<< m1 >>
rect 210 184 211 185 
<< m1 >>
rect 211 184 212 185 
<< m1 >>
rect 212 184 213 185 
<< m1 >>
rect 213 184 214 185 
<< m1 >>
rect 214 184 215 185 
<< m1 >>
rect 229 184 230 185 
<< m1 >>
rect 254 184 255 185 
<< m1 >>
rect 256 184 257 185 
<< m1 >>
rect 19 185 20 186 
<< m1 >>
rect 28 185 29 186 
<< m2 >>
rect 28 185 29 186 
<< m2 >>
rect 46 185 47 186 
<< m2 >>
rect 52 185 53 186 
<< m2 >>
rect 55 185 56 186 
<< m2 >>
rect 59 185 60 186 
<< m2 >>
rect 62 185 63 186 
<< m2 >>
rect 64 185 65 186 
<< m2 >>
rect 73 185 74 186 
<< m2 >>
rect 74 185 75 186 
<< m2 >>
rect 75 185 76 186 
<< m2 >>
rect 76 185 77 186 
<< m2 >>
rect 77 185 78 186 
<< m2 >>
rect 78 185 79 186 
<< m2 >>
rect 79 185 80 186 
<< m2 >>
rect 80 185 81 186 
<< m2 >>
rect 81 185 82 186 
<< m2 >>
rect 82 185 83 186 
<< m2 >>
rect 83 185 84 186 
<< m2 >>
rect 84 185 85 186 
<< m2 >>
rect 85 185 86 186 
<< m2 >>
rect 86 185 87 186 
<< m2 >>
rect 91 185 92 186 
<< m2 >>
rect 108 185 109 186 
<< m2 >>
rect 113 185 114 186 
<< m2 >>
rect 127 185 128 186 
<< m2 >>
rect 129 185 130 186 
<< m2 >>
rect 138 185 139 186 
<< m2 >>
rect 142 185 143 186 
<< m1 >>
rect 175 185 176 186 
<< m2 >>
rect 181 185 182 186 
<< m2 >>
rect 183 185 184 186 
<< m2 >>
rect 185 185 186 186 
<< m2 >>
rect 189 185 190 186 
<< m2 >>
rect 192 185 193 186 
<< m1 >>
rect 214 185 215 186 
<< m1 >>
rect 229 185 230 186 
<< m1 >>
rect 254 185 255 186 
<< m1 >>
rect 256 185 257 186 
<< m1 >>
rect 19 186 20 187 
<< m1 >>
rect 28 186 29 187 
<< m2 >>
rect 28 186 29 187 
<< m1 >>
rect 46 186 47 187 
<< m2 >>
rect 46 186 47 187 
<< m1 >>
rect 47 186 48 187 
<< m1 >>
rect 48 186 49 187 
<< m1 >>
rect 49 186 50 187 
<< m1 >>
rect 50 186 51 187 
<< m1 >>
rect 51 186 52 187 
<< m1 >>
rect 52 186 53 187 
<< m2 >>
rect 52 186 53 187 
<< m1 >>
rect 53 186 54 187 
<< m1 >>
rect 54 186 55 187 
<< m1 >>
rect 55 186 56 187 
<< m2 >>
rect 55 186 56 187 
<< m1 >>
rect 56 186 57 187 
<< m1 >>
rect 57 186 58 187 
<< m1 >>
rect 58 186 59 187 
<< m1 >>
rect 59 186 60 187 
<< m2 >>
rect 59 186 60 187 
<< m1 >>
rect 60 186 61 187 
<< m1 >>
rect 61 186 62 187 
<< m1 >>
rect 62 186 63 187 
<< m2 >>
rect 62 186 63 187 
<< m1 >>
rect 63 186 64 187 
<< m1 >>
rect 64 186 65 187 
<< m2 >>
rect 64 186 65 187 
<< m1 >>
rect 65 186 66 187 
<< m1 >>
rect 66 186 67 187 
<< m1 >>
rect 67 186 68 187 
<< m1 >>
rect 68 186 69 187 
<< m1 >>
rect 69 186 70 187 
<< m1 >>
rect 70 186 71 187 
<< m1 >>
rect 71 186 72 187 
<< m1 >>
rect 72 186 73 187 
<< m1 >>
rect 73 186 74 187 
<< m1 >>
rect 74 186 75 187 
<< m1 >>
rect 75 186 76 187 
<< m1 >>
rect 76 186 77 187 
<< m1 >>
rect 77 186 78 187 
<< m1 >>
rect 78 186 79 187 
<< m1 >>
rect 79 186 80 187 
<< m1 >>
rect 80 186 81 187 
<< m1 >>
rect 81 186 82 187 
<< m1 >>
rect 82 186 83 187 
<< m1 >>
rect 83 186 84 187 
<< m1 >>
rect 84 186 85 187 
<< m1 >>
rect 85 186 86 187 
<< m1 >>
rect 86 186 87 187 
<< m2 >>
rect 86 186 87 187 
<< m1 >>
rect 87 186 88 187 
<< m1 >>
rect 88 186 89 187 
<< m1 >>
rect 89 186 90 187 
<< m1 >>
rect 90 186 91 187 
<< m1 >>
rect 91 186 92 187 
<< m2 >>
rect 91 186 92 187 
<< m1 >>
rect 92 186 93 187 
<< m1 >>
rect 93 186 94 187 
<< m1 >>
rect 94 186 95 187 
<< m1 >>
rect 95 186 96 187 
<< m1 >>
rect 96 186 97 187 
<< m1 >>
rect 97 186 98 187 
<< m1 >>
rect 98 186 99 187 
<< m1 >>
rect 99 186 100 187 
<< m1 >>
rect 100 186 101 187 
<< m1 >>
rect 101 186 102 187 
<< m1 >>
rect 102 186 103 187 
<< m1 >>
rect 103 186 104 187 
<< m1 >>
rect 104 186 105 187 
<< m1 >>
rect 105 186 106 187 
<< m1 >>
rect 106 186 107 187 
<< m1 >>
rect 107 186 108 187 
<< m1 >>
rect 108 186 109 187 
<< m2 >>
rect 108 186 109 187 
<< m1 >>
rect 109 186 110 187 
<< m1 >>
rect 110 186 111 187 
<< m1 >>
rect 111 186 112 187 
<< m1 >>
rect 112 186 113 187 
<< m1 >>
rect 113 186 114 187 
<< m2 >>
rect 113 186 114 187 
<< m1 >>
rect 114 186 115 187 
<< m1 >>
rect 115 186 116 187 
<< m1 >>
rect 116 186 117 187 
<< m1 >>
rect 117 186 118 187 
<< m1 >>
rect 118 186 119 187 
<< m1 >>
rect 119 186 120 187 
<< m1 >>
rect 120 186 121 187 
<< m1 >>
rect 121 186 122 187 
<< m1 >>
rect 122 186 123 187 
<< m1 >>
rect 123 186 124 187 
<< m1 >>
rect 124 186 125 187 
<< m1 >>
rect 125 186 126 187 
<< m1 >>
rect 126 186 127 187 
<< m1 >>
rect 127 186 128 187 
<< m2 >>
rect 127 186 128 187 
<< m1 >>
rect 128 186 129 187 
<< m1 >>
rect 129 186 130 187 
<< m2 >>
rect 129 186 130 187 
<< m1 >>
rect 130 186 131 187 
<< m1 >>
rect 131 186 132 187 
<< m1 >>
rect 132 186 133 187 
<< m1 >>
rect 133 186 134 187 
<< m1 >>
rect 134 186 135 187 
<< m1 >>
rect 135 186 136 187 
<< m1 >>
rect 136 186 137 187 
<< m1 >>
rect 137 186 138 187 
<< m1 >>
rect 138 186 139 187 
<< m2 >>
rect 138 186 139 187 
<< m1 >>
rect 139 186 140 187 
<< m1 >>
rect 140 186 141 187 
<< m1 >>
rect 141 186 142 187 
<< m1 >>
rect 142 186 143 187 
<< m2 >>
rect 142 186 143 187 
<< m2c >>
rect 142 186 143 187 
<< m1 >>
rect 142 186 143 187 
<< m2 >>
rect 142 186 143 187 
<< m1 >>
rect 175 186 176 187 
<< m1 >>
rect 181 186 182 187 
<< m2 >>
rect 181 186 182 187 
<< m2c >>
rect 181 186 182 187 
<< m1 >>
rect 181 186 182 187 
<< m2 >>
rect 181 186 182 187 
<< m1 >>
rect 183 186 184 187 
<< m2 >>
rect 183 186 184 187 
<< m2c >>
rect 183 186 184 187 
<< m1 >>
rect 183 186 184 187 
<< m2 >>
rect 183 186 184 187 
<< m1 >>
rect 184 186 185 187 
<< m1 >>
rect 185 186 186 187 
<< m2 >>
rect 185 186 186 187 
<< m1 >>
rect 186 186 187 187 
<< m1 >>
rect 187 186 188 187 
<< m1 >>
rect 188 186 189 187 
<< m1 >>
rect 189 186 190 187 
<< m2 >>
rect 189 186 190 187 
<< m1 >>
rect 190 186 191 187 
<< m1 >>
rect 191 186 192 187 
<< m1 >>
rect 192 186 193 187 
<< m2 >>
rect 192 186 193 187 
<< m1 >>
rect 193 186 194 187 
<< m1 >>
rect 214 186 215 187 
<< m1 >>
rect 229 186 230 187 
<< m1 >>
rect 254 186 255 187 
<< m1 >>
rect 256 186 257 187 
<< m1 >>
rect 19 187 20 188 
<< m1 >>
rect 28 187 29 188 
<< m2 >>
rect 28 187 29 188 
<< m1 >>
rect 46 187 47 188 
<< m2 >>
rect 46 187 47 188 
<< m2 >>
rect 52 187 53 188 
<< m2 >>
rect 55 187 56 188 
<< m2 >>
rect 59 187 60 188 
<< m2 >>
rect 62 187 63 188 
<< m2 >>
rect 64 187 65 188 
<< m2 >>
rect 86 187 87 188 
<< m2 >>
rect 91 187 92 188 
<< m2 >>
rect 93 187 94 188 
<< m2 >>
rect 94 187 95 188 
<< m2 >>
rect 95 187 96 188 
<< m2 >>
rect 96 187 97 188 
<< m2 >>
rect 97 187 98 188 
<< m2 >>
rect 98 187 99 188 
<< m2 >>
rect 99 187 100 188 
<< m2 >>
rect 100 187 101 188 
<< m2 >>
rect 101 187 102 188 
<< m2 >>
rect 102 187 103 188 
<< m2 >>
rect 103 187 104 188 
<< m2 >>
rect 104 187 105 188 
<< m2 >>
rect 105 187 106 188 
<< m2 >>
rect 106 187 107 188 
<< m2 >>
rect 107 187 108 188 
<< m2 >>
rect 108 187 109 188 
<< m2 >>
rect 113 187 114 188 
<< m2 >>
rect 115 187 116 188 
<< m2 >>
rect 116 187 117 188 
<< m2 >>
rect 117 187 118 188 
<< m2 >>
rect 118 187 119 188 
<< m2 >>
rect 119 187 120 188 
<< m2 >>
rect 120 187 121 188 
<< m2 >>
rect 121 187 122 188 
<< m2 >>
rect 122 187 123 188 
<< m2 >>
rect 127 187 128 188 
<< m2 >>
rect 129 187 130 188 
<< m2 >>
rect 138 187 139 188 
<< m2 >>
rect 139 187 140 188 
<< m2 >>
rect 140 187 141 188 
<< m1 >>
rect 156 187 157 188 
<< m1 >>
rect 157 187 158 188 
<< m1 >>
rect 158 187 159 188 
<< m1 >>
rect 159 187 160 188 
<< m1 >>
rect 160 187 161 188 
<< m1 >>
rect 161 187 162 188 
<< m1 >>
rect 162 187 163 188 
<< m1 >>
rect 163 187 164 188 
<< m1 >>
rect 164 187 165 188 
<< m1 >>
rect 165 187 166 188 
<< m1 >>
rect 166 187 167 188 
<< m1 >>
rect 167 187 168 188 
<< m2 >>
rect 174 187 175 188 
<< m1 >>
rect 175 187 176 188 
<< m2 >>
rect 175 187 176 188 
<< m2 >>
rect 176 187 177 188 
<< m1 >>
rect 177 187 178 188 
<< m2 >>
rect 177 187 178 188 
<< m2c >>
rect 177 187 178 188 
<< m1 >>
rect 177 187 178 188 
<< m2 >>
rect 177 187 178 188 
<< m1 >>
rect 178 187 179 188 
<< m1 >>
rect 181 187 182 188 
<< m2 >>
rect 185 187 186 188 
<< m2 >>
rect 187 187 188 188 
<< m2 >>
rect 188 187 189 188 
<< m2 >>
rect 189 187 190 188 
<< m2 >>
rect 192 187 193 188 
<< m1 >>
rect 193 187 194 188 
<< m2 >>
rect 193 187 194 188 
<< m2 >>
rect 194 187 195 188 
<< m1 >>
rect 199 187 200 188 
<< m2 >>
rect 199 187 200 188 
<< m2c >>
rect 199 187 200 188 
<< m1 >>
rect 199 187 200 188 
<< m2 >>
rect 199 187 200 188 
<< m1 >>
rect 200 187 201 188 
<< m1 >>
rect 201 187 202 188 
<< m1 >>
rect 202 187 203 188 
<< m1 >>
rect 203 187 204 188 
<< m1 >>
rect 204 187 205 188 
<< m1 >>
rect 205 187 206 188 
<< m1 >>
rect 206 187 207 188 
<< m1 >>
rect 207 187 208 188 
<< m1 >>
rect 208 187 209 188 
<< m1 >>
rect 209 187 210 188 
<< m1 >>
rect 210 187 211 188 
<< m1 >>
rect 211 187 212 188 
<< m1 >>
rect 212 187 213 188 
<< m2 >>
rect 212 187 213 188 
<< m2c >>
rect 212 187 213 188 
<< m1 >>
rect 212 187 213 188 
<< m2 >>
rect 212 187 213 188 
<< m2 >>
rect 213 187 214 188 
<< m1 >>
rect 214 187 215 188 
<< m2 >>
rect 214 187 215 188 
<< m2 >>
rect 215 187 216 188 
<< m1 >>
rect 216 187 217 188 
<< m2 >>
rect 216 187 217 188 
<< m2c >>
rect 216 187 217 188 
<< m1 >>
rect 216 187 217 188 
<< m2 >>
rect 216 187 217 188 
<< m1 >>
rect 217 187 218 188 
<< m1 >>
rect 218 187 219 188 
<< m1 >>
rect 219 187 220 188 
<< m1 >>
rect 220 187 221 188 
<< m1 >>
rect 221 187 222 188 
<< m1 >>
rect 222 187 223 188 
<< m1 >>
rect 223 187 224 188 
<< m1 >>
rect 224 187 225 188 
<< m1 >>
rect 225 187 226 188 
<< m1 >>
rect 226 187 227 188 
<< m1 >>
rect 227 187 228 188 
<< m1 >>
rect 228 187 229 188 
<< m1 >>
rect 229 187 230 188 
<< m1 >>
rect 254 187 255 188 
<< m1 >>
rect 256 187 257 188 
<< m1 >>
rect 19 188 20 189 
<< m1 >>
rect 28 188 29 189 
<< m2 >>
rect 28 188 29 189 
<< m1 >>
rect 46 188 47 189 
<< m2 >>
rect 46 188 47 189 
<< m1 >>
rect 52 188 53 189 
<< m2 >>
rect 52 188 53 189 
<< m2c >>
rect 52 188 53 189 
<< m1 >>
rect 52 188 53 189 
<< m2 >>
rect 52 188 53 189 
<< m1 >>
rect 53 188 54 189 
<< m1 >>
rect 54 188 55 189 
<< m1 >>
rect 55 188 56 189 
<< m2 >>
rect 55 188 56 189 
<< m1 >>
rect 59 188 60 189 
<< m2 >>
rect 59 188 60 189 
<< m2c >>
rect 59 188 60 189 
<< m1 >>
rect 59 188 60 189 
<< m2 >>
rect 59 188 60 189 
<< m1 >>
rect 62 188 63 189 
<< m2 >>
rect 62 188 63 189 
<< m2c >>
rect 62 188 63 189 
<< m1 >>
rect 62 188 63 189 
<< m2 >>
rect 62 188 63 189 
<< m1 >>
rect 64 188 65 189 
<< m2 >>
rect 64 188 65 189 
<< m2c >>
rect 64 188 65 189 
<< m1 >>
rect 64 188 65 189 
<< m2 >>
rect 64 188 65 189 
<< m1 >>
rect 86 188 87 189 
<< m2 >>
rect 86 188 87 189 
<< m2c >>
rect 86 188 87 189 
<< m1 >>
rect 86 188 87 189 
<< m2 >>
rect 86 188 87 189 
<< m1 >>
rect 87 188 88 189 
<< m1 >>
rect 88 188 89 189 
<< m1 >>
rect 89 188 90 189 
<< m1 >>
rect 90 188 91 189 
<< m1 >>
rect 91 188 92 189 
<< m2 >>
rect 91 188 92 189 
<< m1 >>
rect 92 188 93 189 
<< m1 >>
rect 93 188 94 189 
<< m2 >>
rect 93 188 94 189 
<< m1 >>
rect 113 188 114 189 
<< m2 >>
rect 113 188 114 189 
<< m2c >>
rect 113 188 114 189 
<< m1 >>
rect 113 188 114 189 
<< m2 >>
rect 113 188 114 189 
<< m1 >>
rect 115 188 116 189 
<< m2 >>
rect 115 188 116 189 
<< m2c >>
rect 115 188 116 189 
<< m1 >>
rect 115 188 116 189 
<< m2 >>
rect 115 188 116 189 
<< m1 >>
rect 122 188 123 189 
<< m2 >>
rect 122 188 123 189 
<< m2c >>
rect 122 188 123 189 
<< m1 >>
rect 122 188 123 189 
<< m2 >>
rect 122 188 123 189 
<< m1 >>
rect 123 188 124 189 
<< m1 >>
rect 124 188 125 189 
<< m1 >>
rect 127 188 128 189 
<< m2 >>
rect 127 188 128 189 
<< m2c >>
rect 127 188 128 189 
<< m1 >>
rect 127 188 128 189 
<< m2 >>
rect 127 188 128 189 
<< m1 >>
rect 129 188 130 189 
<< m2 >>
rect 129 188 130 189 
<< m2c >>
rect 129 188 130 189 
<< m1 >>
rect 129 188 130 189 
<< m2 >>
rect 129 188 130 189 
<< m1 >>
rect 140 188 141 189 
<< m2 >>
rect 140 188 141 189 
<< m2c >>
rect 140 188 141 189 
<< m1 >>
rect 140 188 141 189 
<< m2 >>
rect 140 188 141 189 
<< m2 >>
rect 154 188 155 189 
<< m2 >>
rect 155 188 156 189 
<< m1 >>
rect 156 188 157 189 
<< m2 >>
rect 156 188 157 189 
<< m2c >>
rect 156 188 157 189 
<< m1 >>
rect 156 188 157 189 
<< m2 >>
rect 156 188 157 189 
<< m1 >>
rect 167 188 168 189 
<< m2 >>
rect 167 188 168 189 
<< m2c >>
rect 167 188 168 189 
<< m1 >>
rect 167 188 168 189 
<< m2 >>
rect 167 188 168 189 
<< m2 >>
rect 174 188 175 189 
<< m1 >>
rect 175 188 176 189 
<< m1 >>
rect 178 188 179 189 
<< m1 >>
rect 181 188 182 189 
<< m2 >>
rect 182 188 183 189 
<< m1 >>
rect 183 188 184 189 
<< m2 >>
rect 183 188 184 189 
<< m2c >>
rect 183 188 184 189 
<< m1 >>
rect 183 188 184 189 
<< m2 >>
rect 183 188 184 189 
<< m1 >>
rect 184 188 185 189 
<< m1 >>
rect 185 188 186 189 
<< m2 >>
rect 185 188 186 189 
<< m2c >>
rect 185 188 186 189 
<< m1 >>
rect 185 188 186 189 
<< m2 >>
rect 185 188 186 189 
<< m1 >>
rect 187 188 188 189 
<< m2 >>
rect 187 188 188 189 
<< m2c >>
rect 187 188 188 189 
<< m1 >>
rect 187 188 188 189 
<< m2 >>
rect 187 188 188 189 
<< m1 >>
rect 193 188 194 189 
<< m2 >>
rect 194 188 195 189 
<< m2 >>
rect 199 188 200 189 
<< m1 >>
rect 214 188 215 189 
<< m1 >>
rect 254 188 255 189 
<< m1 >>
rect 256 188 257 189 
<< m1 >>
rect 19 189 20 190 
<< m1 >>
rect 28 189 29 190 
<< m2 >>
rect 28 189 29 190 
<< m1 >>
rect 46 189 47 190 
<< m2 >>
rect 46 189 47 190 
<< m1 >>
rect 55 189 56 190 
<< m2 >>
rect 55 189 56 190 
<< m1 >>
rect 59 189 60 190 
<< m1 >>
rect 62 189 63 190 
<< m1 >>
rect 64 189 65 190 
<< m2 >>
rect 91 189 92 190 
<< m1 >>
rect 93 189 94 190 
<< m2 >>
rect 93 189 94 190 
<< m1 >>
rect 113 189 114 190 
<< m1 >>
rect 115 189 116 190 
<< m1 >>
rect 124 189 125 190 
<< m1 >>
rect 127 189 128 190 
<< m1 >>
rect 129 189 130 190 
<< m1 >>
rect 140 189 141 190 
<< m1 >>
rect 141 189 142 190 
<< m1 >>
rect 142 189 143 190 
<< m1 >>
rect 143 189 144 190 
<< m1 >>
rect 144 189 145 190 
<< m1 >>
rect 145 189 146 190 
<< m1 >>
rect 146 189 147 190 
<< m1 >>
rect 147 189 148 190 
<< m1 >>
rect 148 189 149 190 
<< m1 >>
rect 149 189 150 190 
<< m1 >>
rect 150 189 151 190 
<< m1 >>
rect 151 189 152 190 
<< m1 >>
rect 152 189 153 190 
<< m1 >>
rect 153 189 154 190 
<< m1 >>
rect 154 189 155 190 
<< m2 >>
rect 154 189 155 190 
<< m2 >>
rect 167 189 168 190 
<< m2 >>
rect 174 189 175 190 
<< m1 >>
rect 175 189 176 190 
<< m1 >>
rect 178 189 179 190 
<< m1 >>
rect 181 189 182 190 
<< m2 >>
rect 182 189 183 190 
<< m1 >>
rect 187 189 188 190 
<< m1 >>
rect 193 189 194 190 
<< m2 >>
rect 194 189 195 190 
<< m1 >>
rect 195 189 196 190 
<< m2 >>
rect 195 189 196 190 
<< m2c >>
rect 195 189 196 190 
<< m1 >>
rect 195 189 196 190 
<< m2 >>
rect 195 189 196 190 
<< m1 >>
rect 196 189 197 190 
<< m1 >>
rect 197 189 198 190 
<< m1 >>
rect 198 189 199 190 
<< m1 >>
rect 199 189 200 190 
<< m2 >>
rect 199 189 200 190 
<< m1 >>
rect 200 189 201 190 
<< m1 >>
rect 201 189 202 190 
<< m1 >>
rect 202 189 203 190 
<< m1 >>
rect 203 189 204 190 
<< m1 >>
rect 204 189 205 190 
<< m1 >>
rect 205 189 206 190 
<< m1 >>
rect 206 189 207 190 
<< m1 >>
rect 207 189 208 190 
<< m1 >>
rect 208 189 209 190 
<< m1 >>
rect 209 189 210 190 
<< m1 >>
rect 210 189 211 190 
<< m1 >>
rect 211 189 212 190 
<< m1 >>
rect 214 189 215 190 
<< m1 >>
rect 254 189 255 190 
<< m1 >>
rect 256 189 257 190 
<< m1 >>
rect 19 190 20 191 
<< m1 >>
rect 28 190 29 191 
<< m2 >>
rect 28 190 29 191 
<< m1 >>
rect 46 190 47 191 
<< m2 >>
rect 46 190 47 191 
<< m1 >>
rect 55 190 56 191 
<< m2 >>
rect 55 190 56 191 
<< m1 >>
rect 59 190 60 191 
<< m1 >>
rect 62 190 63 191 
<< m2 >>
rect 62 190 63 191 
<< m2c >>
rect 62 190 63 191 
<< m1 >>
rect 62 190 63 191 
<< m2 >>
rect 62 190 63 191 
<< m2 >>
rect 63 190 64 191 
<< m1 >>
rect 64 190 65 191 
<< m2 >>
rect 64 190 65 191 
<< m2 >>
rect 65 190 66 191 
<< m1 >>
rect 66 190 67 191 
<< m2 >>
rect 66 190 67 191 
<< m2c >>
rect 66 190 67 191 
<< m1 >>
rect 66 190 67 191 
<< m2 >>
rect 66 190 67 191 
<< m1 >>
rect 67 190 68 191 
<< m1 >>
rect 82 190 83 191 
<< m1 >>
rect 83 190 84 191 
<< m1 >>
rect 84 190 85 191 
<< m1 >>
rect 85 190 86 191 
<< m1 >>
rect 88 190 89 191 
<< m1 >>
rect 89 190 90 191 
<< m1 >>
rect 90 190 91 191 
<< m1 >>
rect 91 190 92 191 
<< m2 >>
rect 91 190 92 191 
<< m1 >>
rect 93 190 94 191 
<< m2 >>
rect 93 190 94 191 
<< m1 >>
rect 113 190 114 191 
<< m1 >>
rect 115 190 116 191 
<< m1 >>
rect 124 190 125 191 
<< m1 >>
rect 127 190 128 191 
<< m1 >>
rect 129 190 130 191 
<< m1 >>
rect 136 190 137 191 
<< m1 >>
rect 137 190 138 191 
<< m1 >>
rect 138 190 139 191 
<< m2 >>
rect 138 190 139 191 
<< m2 >>
rect 139 190 140 191 
<< m1 >>
rect 154 190 155 191 
<< m2 >>
rect 154 190 155 191 
<< m1 >>
rect 160 190 161 191 
<< m1 >>
rect 161 190 162 191 
<< m2 >>
rect 161 190 162 191 
<< m2c >>
rect 161 190 162 191 
<< m1 >>
rect 161 190 162 191 
<< m2 >>
rect 161 190 162 191 
<< m2 >>
rect 162 190 163 191 
<< m1 >>
rect 163 190 164 191 
<< m2 >>
rect 163 190 164 191 
<< m1 >>
rect 164 190 165 191 
<< m1 >>
rect 165 190 166 191 
<< m1 >>
rect 166 190 167 191 
<< m1 >>
rect 167 190 168 191 
<< m2 >>
rect 167 190 168 191 
<< m1 >>
rect 168 190 169 191 
<< m1 >>
rect 169 190 170 191 
<< m1 >>
rect 170 190 171 191 
<< m1 >>
rect 171 190 172 191 
<< m1 >>
rect 172 190 173 191 
<< m1 >>
rect 173 190 174 191 
<< m2 >>
rect 173 190 174 191 
<< m2c >>
rect 173 190 174 191 
<< m1 >>
rect 173 190 174 191 
<< m2 >>
rect 173 190 174 191 
<< m2 >>
rect 174 190 175 191 
<< m1 >>
rect 175 190 176 191 
<< m1 >>
rect 178 190 179 191 
<< m1 >>
rect 181 190 182 191 
<< m2 >>
rect 182 190 183 191 
<< m1 >>
rect 187 190 188 191 
<< m1 >>
rect 193 190 194 191 
<< m2 >>
rect 199 190 200 191 
<< m1 >>
rect 211 190 212 191 
<< m1 >>
rect 214 190 215 191 
<< m1 >>
rect 250 190 251 191 
<< m1 >>
rect 251 190 252 191 
<< m1 >>
rect 252 190 253 191 
<< m1 >>
rect 253 190 254 191 
<< m1 >>
rect 254 190 255 191 
<< m1 >>
rect 256 190 257 191 
<< m1 >>
rect 19 191 20 192 
<< m1 >>
rect 28 191 29 192 
<< m2 >>
rect 28 191 29 192 
<< m1 >>
rect 46 191 47 192 
<< m2 >>
rect 46 191 47 192 
<< m1 >>
rect 55 191 56 192 
<< m2 >>
rect 55 191 56 192 
<< m1 >>
rect 59 191 60 192 
<< m1 >>
rect 64 191 65 192 
<< m1 >>
rect 67 191 68 192 
<< m1 >>
rect 82 191 83 192 
<< m1 >>
rect 85 191 86 192 
<< m1 >>
rect 88 191 89 192 
<< m1 >>
rect 91 191 92 192 
<< m2 >>
rect 91 191 92 192 
<< m1 >>
rect 93 191 94 192 
<< m2 >>
rect 93 191 94 192 
<< m1 >>
rect 113 191 114 192 
<< m1 >>
rect 115 191 116 192 
<< m1 >>
rect 124 191 125 192 
<< m1 >>
rect 127 191 128 192 
<< m1 >>
rect 129 191 130 192 
<< m1 >>
rect 136 191 137 192 
<< m1 >>
rect 139 191 140 192 
<< m2 >>
rect 139 191 140 192 
<< m1 >>
rect 150 191 151 192 
<< m1 >>
rect 151 191 152 192 
<< m1 >>
rect 152 191 153 192 
<< m2 >>
rect 152 191 153 192 
<< m2c >>
rect 152 191 153 192 
<< m1 >>
rect 152 191 153 192 
<< m2 >>
rect 152 191 153 192 
<< m2 >>
rect 153 191 154 192 
<< m1 >>
rect 154 191 155 192 
<< m2 >>
rect 154 191 155 192 
<< m1 >>
rect 160 191 161 192 
<< m1 >>
rect 163 191 164 192 
<< m2 >>
rect 163 191 164 192 
<< m2 >>
rect 167 191 168 192 
<< m1 >>
rect 175 191 176 192 
<< m1 >>
rect 178 191 179 192 
<< m1 >>
rect 181 191 182 192 
<< m2 >>
rect 182 191 183 192 
<< m1 >>
rect 187 191 188 192 
<< m1 >>
rect 193 191 194 192 
<< m1 >>
rect 199 191 200 192 
<< m2 >>
rect 199 191 200 192 
<< m2c >>
rect 199 191 200 192 
<< m1 >>
rect 199 191 200 192 
<< m2 >>
rect 199 191 200 192 
<< m1 >>
rect 211 191 212 192 
<< m1 >>
rect 214 191 215 192 
<< m1 >>
rect 250 191 251 192 
<< m1 >>
rect 256 191 257 192 
<< pdiffusion >>
rect 12 192 13 193 
<< pdiffusion >>
rect 13 192 14 193 
<< pdiffusion >>
rect 14 192 15 193 
<< pdiffusion >>
rect 15 192 16 193 
<< pdiffusion >>
rect 16 192 17 193 
<< pdiffusion >>
rect 17 192 18 193 
<< m1 >>
rect 19 192 20 193 
<< m1 >>
rect 28 192 29 193 
<< m2 >>
rect 28 192 29 193 
<< pdiffusion >>
rect 30 192 31 193 
<< pdiffusion >>
rect 31 192 32 193 
<< pdiffusion >>
rect 32 192 33 193 
<< pdiffusion >>
rect 33 192 34 193 
<< pdiffusion >>
rect 34 192 35 193 
<< pdiffusion >>
rect 35 192 36 193 
<< m1 >>
rect 46 192 47 193 
<< m2 >>
rect 46 192 47 193 
<< pdiffusion >>
rect 48 192 49 193 
<< pdiffusion >>
rect 49 192 50 193 
<< pdiffusion >>
rect 50 192 51 193 
<< pdiffusion >>
rect 51 192 52 193 
<< pdiffusion >>
rect 52 192 53 193 
<< pdiffusion >>
rect 53 192 54 193 
<< m1 >>
rect 55 192 56 193 
<< m2 >>
rect 55 192 56 193 
<< m1 >>
rect 59 192 60 193 
<< m1 >>
rect 64 192 65 193 
<< pdiffusion >>
rect 66 192 67 193 
<< m1 >>
rect 67 192 68 193 
<< pdiffusion >>
rect 67 192 68 193 
<< pdiffusion >>
rect 68 192 69 193 
<< pdiffusion >>
rect 69 192 70 193 
<< pdiffusion >>
rect 70 192 71 193 
<< pdiffusion >>
rect 71 192 72 193 
<< m1 >>
rect 82 192 83 193 
<< pdiffusion >>
rect 84 192 85 193 
<< m1 >>
rect 85 192 86 193 
<< pdiffusion >>
rect 85 192 86 193 
<< pdiffusion >>
rect 86 192 87 193 
<< pdiffusion >>
rect 87 192 88 193 
<< m1 >>
rect 88 192 89 193 
<< pdiffusion >>
rect 88 192 89 193 
<< pdiffusion >>
rect 89 192 90 193 
<< m1 >>
rect 91 192 92 193 
<< m2 >>
rect 91 192 92 193 
<< m1 >>
rect 93 192 94 193 
<< m2 >>
rect 93 192 94 193 
<< pdiffusion >>
rect 102 192 103 193 
<< pdiffusion >>
rect 103 192 104 193 
<< pdiffusion >>
rect 104 192 105 193 
<< pdiffusion >>
rect 105 192 106 193 
<< pdiffusion >>
rect 106 192 107 193 
<< pdiffusion >>
rect 107 192 108 193 
<< m1 >>
rect 113 192 114 193 
<< m1 >>
rect 115 192 116 193 
<< pdiffusion >>
rect 120 192 121 193 
<< pdiffusion >>
rect 121 192 122 193 
<< pdiffusion >>
rect 122 192 123 193 
<< pdiffusion >>
rect 123 192 124 193 
<< m1 >>
rect 124 192 125 193 
<< pdiffusion >>
rect 124 192 125 193 
<< pdiffusion >>
rect 125 192 126 193 
<< m1 >>
rect 127 192 128 193 
<< m1 >>
rect 129 192 130 193 
<< m1 >>
rect 136 192 137 193 
<< m1 >>
rect 138 192 139 193 
<< m2 >>
rect 138 192 139 193 
<< m2c >>
rect 138 192 139 193 
<< m1 >>
rect 138 192 139 193 
<< m2 >>
rect 138 192 139 193 
<< pdiffusion >>
rect 138 192 139 193 
<< m1 >>
rect 139 192 140 193 
<< pdiffusion >>
rect 139 192 140 193 
<< pdiffusion >>
rect 140 192 141 193 
<< pdiffusion >>
rect 141 192 142 193 
<< pdiffusion >>
rect 142 192 143 193 
<< pdiffusion >>
rect 143 192 144 193 
<< m1 >>
rect 150 192 151 193 
<< m1 >>
rect 154 192 155 193 
<< pdiffusion >>
rect 156 192 157 193 
<< pdiffusion >>
rect 157 192 158 193 
<< pdiffusion >>
rect 158 192 159 193 
<< pdiffusion >>
rect 159 192 160 193 
<< m1 >>
rect 160 192 161 193 
<< pdiffusion >>
rect 160 192 161 193 
<< pdiffusion >>
rect 161 192 162 193 
<< m1 >>
rect 163 192 164 193 
<< m2 >>
rect 163 192 164 193 
<< m2 >>
rect 164 192 165 193 
<< m1 >>
rect 165 192 166 193 
<< m2 >>
rect 165 192 166 193 
<< m2c >>
rect 165 192 166 193 
<< m1 >>
rect 165 192 166 193 
<< m2 >>
rect 165 192 166 193 
<< m1 >>
rect 166 192 167 193 
<< m1 >>
rect 167 192 168 193 
<< m2 >>
rect 167 192 168 193 
<< pdiffusion >>
rect 174 192 175 193 
<< m1 >>
rect 175 192 176 193 
<< pdiffusion >>
rect 175 192 176 193 
<< pdiffusion >>
rect 176 192 177 193 
<< pdiffusion >>
rect 177 192 178 193 
<< m1 >>
rect 178 192 179 193 
<< pdiffusion >>
rect 178 192 179 193 
<< pdiffusion >>
rect 179 192 180 193 
<< m1 >>
rect 181 192 182 193 
<< m2 >>
rect 182 192 183 193 
<< m1 >>
rect 187 192 188 193 
<< pdiffusion >>
rect 192 192 193 193 
<< m1 >>
rect 193 192 194 193 
<< pdiffusion >>
rect 193 192 194 193 
<< pdiffusion >>
rect 194 192 195 193 
<< pdiffusion >>
rect 195 192 196 193 
<< pdiffusion >>
rect 196 192 197 193 
<< pdiffusion >>
rect 197 192 198 193 
<< m1 >>
rect 199 192 200 193 
<< pdiffusion >>
rect 210 192 211 193 
<< m1 >>
rect 211 192 212 193 
<< pdiffusion >>
rect 211 192 212 193 
<< pdiffusion >>
rect 212 192 213 193 
<< pdiffusion >>
rect 213 192 214 193 
<< m1 >>
rect 214 192 215 193 
<< pdiffusion >>
rect 214 192 215 193 
<< pdiffusion >>
rect 215 192 216 193 
<< pdiffusion >>
rect 228 192 229 193 
<< pdiffusion >>
rect 229 192 230 193 
<< pdiffusion >>
rect 230 192 231 193 
<< pdiffusion >>
rect 231 192 232 193 
<< pdiffusion >>
rect 232 192 233 193 
<< pdiffusion >>
rect 233 192 234 193 
<< pdiffusion >>
rect 246 192 247 193 
<< pdiffusion >>
rect 247 192 248 193 
<< pdiffusion >>
rect 248 192 249 193 
<< pdiffusion >>
rect 249 192 250 193 
<< m1 >>
rect 250 192 251 193 
<< pdiffusion >>
rect 250 192 251 193 
<< pdiffusion >>
rect 251 192 252 193 
<< m1 >>
rect 256 192 257 193 
<< pdiffusion >>
rect 12 193 13 194 
<< pdiffusion >>
rect 13 193 14 194 
<< pdiffusion >>
rect 14 193 15 194 
<< pdiffusion >>
rect 15 193 16 194 
<< pdiffusion >>
rect 16 193 17 194 
<< pdiffusion >>
rect 17 193 18 194 
<< m1 >>
rect 19 193 20 194 
<< m1 >>
rect 28 193 29 194 
<< m2 >>
rect 28 193 29 194 
<< pdiffusion >>
rect 30 193 31 194 
<< pdiffusion >>
rect 31 193 32 194 
<< pdiffusion >>
rect 32 193 33 194 
<< pdiffusion >>
rect 33 193 34 194 
<< pdiffusion >>
rect 34 193 35 194 
<< pdiffusion >>
rect 35 193 36 194 
<< m1 >>
rect 46 193 47 194 
<< m2 >>
rect 46 193 47 194 
<< pdiffusion >>
rect 48 193 49 194 
<< pdiffusion >>
rect 49 193 50 194 
<< pdiffusion >>
rect 50 193 51 194 
<< pdiffusion >>
rect 51 193 52 194 
<< pdiffusion >>
rect 52 193 53 194 
<< pdiffusion >>
rect 53 193 54 194 
<< m1 >>
rect 55 193 56 194 
<< m2 >>
rect 55 193 56 194 
<< m1 >>
rect 59 193 60 194 
<< m1 >>
rect 64 193 65 194 
<< pdiffusion >>
rect 66 193 67 194 
<< pdiffusion >>
rect 67 193 68 194 
<< pdiffusion >>
rect 68 193 69 194 
<< pdiffusion >>
rect 69 193 70 194 
<< pdiffusion >>
rect 70 193 71 194 
<< pdiffusion >>
rect 71 193 72 194 
<< m1 >>
rect 82 193 83 194 
<< pdiffusion >>
rect 84 193 85 194 
<< pdiffusion >>
rect 85 193 86 194 
<< pdiffusion >>
rect 86 193 87 194 
<< pdiffusion >>
rect 87 193 88 194 
<< pdiffusion >>
rect 88 193 89 194 
<< pdiffusion >>
rect 89 193 90 194 
<< m1 >>
rect 91 193 92 194 
<< m2 >>
rect 91 193 92 194 
<< m1 >>
rect 93 193 94 194 
<< m2 >>
rect 93 193 94 194 
<< pdiffusion >>
rect 102 193 103 194 
<< pdiffusion >>
rect 103 193 104 194 
<< pdiffusion >>
rect 104 193 105 194 
<< pdiffusion >>
rect 105 193 106 194 
<< pdiffusion >>
rect 106 193 107 194 
<< pdiffusion >>
rect 107 193 108 194 
<< m1 >>
rect 113 193 114 194 
<< m1 >>
rect 115 193 116 194 
<< pdiffusion >>
rect 120 193 121 194 
<< pdiffusion >>
rect 121 193 122 194 
<< pdiffusion >>
rect 122 193 123 194 
<< pdiffusion >>
rect 123 193 124 194 
<< pdiffusion >>
rect 124 193 125 194 
<< pdiffusion >>
rect 125 193 126 194 
<< m1 >>
rect 127 193 128 194 
<< m1 >>
rect 129 193 130 194 
<< m1 >>
rect 136 193 137 194 
<< pdiffusion >>
rect 138 193 139 194 
<< pdiffusion >>
rect 139 193 140 194 
<< pdiffusion >>
rect 140 193 141 194 
<< pdiffusion >>
rect 141 193 142 194 
<< pdiffusion >>
rect 142 193 143 194 
<< pdiffusion >>
rect 143 193 144 194 
<< m1 >>
rect 150 193 151 194 
<< m1 >>
rect 154 193 155 194 
<< pdiffusion >>
rect 156 193 157 194 
<< pdiffusion >>
rect 157 193 158 194 
<< pdiffusion >>
rect 158 193 159 194 
<< pdiffusion >>
rect 159 193 160 194 
<< pdiffusion >>
rect 160 193 161 194 
<< pdiffusion >>
rect 161 193 162 194 
<< m1 >>
rect 163 193 164 194 
<< m1 >>
rect 167 193 168 194 
<< m2 >>
rect 167 193 168 194 
<< pdiffusion >>
rect 174 193 175 194 
<< pdiffusion >>
rect 175 193 176 194 
<< pdiffusion >>
rect 176 193 177 194 
<< pdiffusion >>
rect 177 193 178 194 
<< pdiffusion >>
rect 178 193 179 194 
<< pdiffusion >>
rect 179 193 180 194 
<< m1 >>
rect 181 193 182 194 
<< m2 >>
rect 182 193 183 194 
<< m1 >>
rect 187 193 188 194 
<< pdiffusion >>
rect 192 193 193 194 
<< pdiffusion >>
rect 193 193 194 194 
<< pdiffusion >>
rect 194 193 195 194 
<< pdiffusion >>
rect 195 193 196 194 
<< pdiffusion >>
rect 196 193 197 194 
<< pdiffusion >>
rect 197 193 198 194 
<< m1 >>
rect 199 193 200 194 
<< pdiffusion >>
rect 210 193 211 194 
<< pdiffusion >>
rect 211 193 212 194 
<< pdiffusion >>
rect 212 193 213 194 
<< pdiffusion >>
rect 213 193 214 194 
<< pdiffusion >>
rect 214 193 215 194 
<< pdiffusion >>
rect 215 193 216 194 
<< pdiffusion >>
rect 228 193 229 194 
<< pdiffusion >>
rect 229 193 230 194 
<< pdiffusion >>
rect 230 193 231 194 
<< pdiffusion >>
rect 231 193 232 194 
<< pdiffusion >>
rect 232 193 233 194 
<< pdiffusion >>
rect 233 193 234 194 
<< pdiffusion >>
rect 246 193 247 194 
<< pdiffusion >>
rect 247 193 248 194 
<< pdiffusion >>
rect 248 193 249 194 
<< pdiffusion >>
rect 249 193 250 194 
<< pdiffusion >>
rect 250 193 251 194 
<< pdiffusion >>
rect 251 193 252 194 
<< m1 >>
rect 256 193 257 194 
<< pdiffusion >>
rect 12 194 13 195 
<< pdiffusion >>
rect 13 194 14 195 
<< pdiffusion >>
rect 14 194 15 195 
<< pdiffusion >>
rect 15 194 16 195 
<< pdiffusion >>
rect 16 194 17 195 
<< pdiffusion >>
rect 17 194 18 195 
<< m1 >>
rect 19 194 20 195 
<< m1 >>
rect 28 194 29 195 
<< m2 >>
rect 28 194 29 195 
<< pdiffusion >>
rect 30 194 31 195 
<< pdiffusion >>
rect 31 194 32 195 
<< pdiffusion >>
rect 32 194 33 195 
<< pdiffusion >>
rect 33 194 34 195 
<< pdiffusion >>
rect 34 194 35 195 
<< pdiffusion >>
rect 35 194 36 195 
<< m1 >>
rect 46 194 47 195 
<< m2 >>
rect 46 194 47 195 
<< pdiffusion >>
rect 48 194 49 195 
<< pdiffusion >>
rect 49 194 50 195 
<< pdiffusion >>
rect 50 194 51 195 
<< pdiffusion >>
rect 51 194 52 195 
<< pdiffusion >>
rect 52 194 53 195 
<< pdiffusion >>
rect 53 194 54 195 
<< m1 >>
rect 55 194 56 195 
<< m2 >>
rect 55 194 56 195 
<< m1 >>
rect 59 194 60 195 
<< m1 >>
rect 64 194 65 195 
<< pdiffusion >>
rect 66 194 67 195 
<< pdiffusion >>
rect 67 194 68 195 
<< pdiffusion >>
rect 68 194 69 195 
<< pdiffusion >>
rect 69 194 70 195 
<< pdiffusion >>
rect 70 194 71 195 
<< pdiffusion >>
rect 71 194 72 195 
<< m1 >>
rect 82 194 83 195 
<< pdiffusion >>
rect 84 194 85 195 
<< pdiffusion >>
rect 85 194 86 195 
<< pdiffusion >>
rect 86 194 87 195 
<< pdiffusion >>
rect 87 194 88 195 
<< pdiffusion >>
rect 88 194 89 195 
<< pdiffusion >>
rect 89 194 90 195 
<< m1 >>
rect 91 194 92 195 
<< m2 >>
rect 91 194 92 195 
<< m1 >>
rect 93 194 94 195 
<< m2 >>
rect 93 194 94 195 
<< pdiffusion >>
rect 102 194 103 195 
<< pdiffusion >>
rect 103 194 104 195 
<< pdiffusion >>
rect 104 194 105 195 
<< pdiffusion >>
rect 105 194 106 195 
<< pdiffusion >>
rect 106 194 107 195 
<< pdiffusion >>
rect 107 194 108 195 
<< m1 >>
rect 113 194 114 195 
<< m1 >>
rect 115 194 116 195 
<< pdiffusion >>
rect 120 194 121 195 
<< pdiffusion >>
rect 121 194 122 195 
<< pdiffusion >>
rect 122 194 123 195 
<< pdiffusion >>
rect 123 194 124 195 
<< pdiffusion >>
rect 124 194 125 195 
<< pdiffusion >>
rect 125 194 126 195 
<< m1 >>
rect 127 194 128 195 
<< m1 >>
rect 129 194 130 195 
<< m1 >>
rect 136 194 137 195 
<< pdiffusion >>
rect 138 194 139 195 
<< pdiffusion >>
rect 139 194 140 195 
<< pdiffusion >>
rect 140 194 141 195 
<< pdiffusion >>
rect 141 194 142 195 
<< pdiffusion >>
rect 142 194 143 195 
<< pdiffusion >>
rect 143 194 144 195 
<< m1 >>
rect 150 194 151 195 
<< m1 >>
rect 154 194 155 195 
<< pdiffusion >>
rect 156 194 157 195 
<< pdiffusion >>
rect 157 194 158 195 
<< pdiffusion >>
rect 158 194 159 195 
<< pdiffusion >>
rect 159 194 160 195 
<< pdiffusion >>
rect 160 194 161 195 
<< pdiffusion >>
rect 161 194 162 195 
<< m1 >>
rect 163 194 164 195 
<< m1 >>
rect 167 194 168 195 
<< m2 >>
rect 167 194 168 195 
<< pdiffusion >>
rect 174 194 175 195 
<< pdiffusion >>
rect 175 194 176 195 
<< pdiffusion >>
rect 176 194 177 195 
<< pdiffusion >>
rect 177 194 178 195 
<< pdiffusion >>
rect 178 194 179 195 
<< pdiffusion >>
rect 179 194 180 195 
<< m1 >>
rect 181 194 182 195 
<< m2 >>
rect 182 194 183 195 
<< m1 >>
rect 187 194 188 195 
<< pdiffusion >>
rect 192 194 193 195 
<< pdiffusion >>
rect 193 194 194 195 
<< pdiffusion >>
rect 194 194 195 195 
<< pdiffusion >>
rect 195 194 196 195 
<< pdiffusion >>
rect 196 194 197 195 
<< pdiffusion >>
rect 197 194 198 195 
<< m1 >>
rect 199 194 200 195 
<< pdiffusion >>
rect 210 194 211 195 
<< pdiffusion >>
rect 211 194 212 195 
<< pdiffusion >>
rect 212 194 213 195 
<< pdiffusion >>
rect 213 194 214 195 
<< pdiffusion >>
rect 214 194 215 195 
<< pdiffusion >>
rect 215 194 216 195 
<< pdiffusion >>
rect 228 194 229 195 
<< pdiffusion >>
rect 229 194 230 195 
<< pdiffusion >>
rect 230 194 231 195 
<< pdiffusion >>
rect 231 194 232 195 
<< pdiffusion >>
rect 232 194 233 195 
<< pdiffusion >>
rect 233 194 234 195 
<< pdiffusion >>
rect 246 194 247 195 
<< pdiffusion >>
rect 247 194 248 195 
<< pdiffusion >>
rect 248 194 249 195 
<< pdiffusion >>
rect 249 194 250 195 
<< pdiffusion >>
rect 250 194 251 195 
<< pdiffusion >>
rect 251 194 252 195 
<< m1 >>
rect 256 194 257 195 
<< pdiffusion >>
rect 12 195 13 196 
<< pdiffusion >>
rect 13 195 14 196 
<< pdiffusion >>
rect 14 195 15 196 
<< pdiffusion >>
rect 15 195 16 196 
<< pdiffusion >>
rect 16 195 17 196 
<< pdiffusion >>
rect 17 195 18 196 
<< m1 >>
rect 19 195 20 196 
<< m1 >>
rect 28 195 29 196 
<< m2 >>
rect 28 195 29 196 
<< pdiffusion >>
rect 30 195 31 196 
<< pdiffusion >>
rect 31 195 32 196 
<< pdiffusion >>
rect 32 195 33 196 
<< pdiffusion >>
rect 33 195 34 196 
<< pdiffusion >>
rect 34 195 35 196 
<< pdiffusion >>
rect 35 195 36 196 
<< m1 >>
rect 46 195 47 196 
<< m2 >>
rect 46 195 47 196 
<< pdiffusion >>
rect 48 195 49 196 
<< pdiffusion >>
rect 49 195 50 196 
<< pdiffusion >>
rect 50 195 51 196 
<< pdiffusion >>
rect 51 195 52 196 
<< pdiffusion >>
rect 52 195 53 196 
<< pdiffusion >>
rect 53 195 54 196 
<< m1 >>
rect 55 195 56 196 
<< m2 >>
rect 55 195 56 196 
<< m1 >>
rect 59 195 60 196 
<< m1 >>
rect 64 195 65 196 
<< pdiffusion >>
rect 66 195 67 196 
<< pdiffusion >>
rect 67 195 68 196 
<< pdiffusion >>
rect 68 195 69 196 
<< pdiffusion >>
rect 69 195 70 196 
<< pdiffusion >>
rect 70 195 71 196 
<< pdiffusion >>
rect 71 195 72 196 
<< m1 >>
rect 82 195 83 196 
<< pdiffusion >>
rect 84 195 85 196 
<< pdiffusion >>
rect 85 195 86 196 
<< pdiffusion >>
rect 86 195 87 196 
<< pdiffusion >>
rect 87 195 88 196 
<< pdiffusion >>
rect 88 195 89 196 
<< pdiffusion >>
rect 89 195 90 196 
<< m1 >>
rect 91 195 92 196 
<< m2 >>
rect 91 195 92 196 
<< m1 >>
rect 93 195 94 196 
<< m2 >>
rect 93 195 94 196 
<< pdiffusion >>
rect 102 195 103 196 
<< pdiffusion >>
rect 103 195 104 196 
<< pdiffusion >>
rect 104 195 105 196 
<< pdiffusion >>
rect 105 195 106 196 
<< pdiffusion >>
rect 106 195 107 196 
<< pdiffusion >>
rect 107 195 108 196 
<< m1 >>
rect 113 195 114 196 
<< m1 >>
rect 115 195 116 196 
<< pdiffusion >>
rect 120 195 121 196 
<< pdiffusion >>
rect 121 195 122 196 
<< pdiffusion >>
rect 122 195 123 196 
<< pdiffusion >>
rect 123 195 124 196 
<< pdiffusion >>
rect 124 195 125 196 
<< pdiffusion >>
rect 125 195 126 196 
<< m1 >>
rect 127 195 128 196 
<< m1 >>
rect 129 195 130 196 
<< m1 >>
rect 136 195 137 196 
<< pdiffusion >>
rect 138 195 139 196 
<< pdiffusion >>
rect 139 195 140 196 
<< pdiffusion >>
rect 140 195 141 196 
<< pdiffusion >>
rect 141 195 142 196 
<< pdiffusion >>
rect 142 195 143 196 
<< pdiffusion >>
rect 143 195 144 196 
<< m1 >>
rect 150 195 151 196 
<< m1 >>
rect 154 195 155 196 
<< pdiffusion >>
rect 156 195 157 196 
<< pdiffusion >>
rect 157 195 158 196 
<< pdiffusion >>
rect 158 195 159 196 
<< pdiffusion >>
rect 159 195 160 196 
<< pdiffusion >>
rect 160 195 161 196 
<< pdiffusion >>
rect 161 195 162 196 
<< m1 >>
rect 163 195 164 196 
<< m1 >>
rect 167 195 168 196 
<< m2 >>
rect 167 195 168 196 
<< pdiffusion >>
rect 174 195 175 196 
<< pdiffusion >>
rect 175 195 176 196 
<< pdiffusion >>
rect 176 195 177 196 
<< pdiffusion >>
rect 177 195 178 196 
<< pdiffusion >>
rect 178 195 179 196 
<< pdiffusion >>
rect 179 195 180 196 
<< m1 >>
rect 181 195 182 196 
<< m2 >>
rect 182 195 183 196 
<< m1 >>
rect 187 195 188 196 
<< pdiffusion >>
rect 192 195 193 196 
<< pdiffusion >>
rect 193 195 194 196 
<< pdiffusion >>
rect 194 195 195 196 
<< pdiffusion >>
rect 195 195 196 196 
<< pdiffusion >>
rect 196 195 197 196 
<< pdiffusion >>
rect 197 195 198 196 
<< m1 >>
rect 199 195 200 196 
<< pdiffusion >>
rect 210 195 211 196 
<< pdiffusion >>
rect 211 195 212 196 
<< pdiffusion >>
rect 212 195 213 196 
<< pdiffusion >>
rect 213 195 214 196 
<< pdiffusion >>
rect 214 195 215 196 
<< pdiffusion >>
rect 215 195 216 196 
<< pdiffusion >>
rect 228 195 229 196 
<< pdiffusion >>
rect 229 195 230 196 
<< pdiffusion >>
rect 230 195 231 196 
<< pdiffusion >>
rect 231 195 232 196 
<< pdiffusion >>
rect 232 195 233 196 
<< pdiffusion >>
rect 233 195 234 196 
<< pdiffusion >>
rect 246 195 247 196 
<< pdiffusion >>
rect 247 195 248 196 
<< pdiffusion >>
rect 248 195 249 196 
<< pdiffusion >>
rect 249 195 250 196 
<< pdiffusion >>
rect 250 195 251 196 
<< pdiffusion >>
rect 251 195 252 196 
<< m1 >>
rect 256 195 257 196 
<< pdiffusion >>
rect 12 196 13 197 
<< pdiffusion >>
rect 13 196 14 197 
<< pdiffusion >>
rect 14 196 15 197 
<< pdiffusion >>
rect 15 196 16 197 
<< pdiffusion >>
rect 16 196 17 197 
<< pdiffusion >>
rect 17 196 18 197 
<< m1 >>
rect 19 196 20 197 
<< m1 >>
rect 28 196 29 197 
<< m2 >>
rect 28 196 29 197 
<< pdiffusion >>
rect 30 196 31 197 
<< pdiffusion >>
rect 31 196 32 197 
<< pdiffusion >>
rect 32 196 33 197 
<< pdiffusion >>
rect 33 196 34 197 
<< pdiffusion >>
rect 34 196 35 197 
<< pdiffusion >>
rect 35 196 36 197 
<< m1 >>
rect 46 196 47 197 
<< m2 >>
rect 46 196 47 197 
<< pdiffusion >>
rect 48 196 49 197 
<< pdiffusion >>
rect 49 196 50 197 
<< pdiffusion >>
rect 50 196 51 197 
<< pdiffusion >>
rect 51 196 52 197 
<< pdiffusion >>
rect 52 196 53 197 
<< pdiffusion >>
rect 53 196 54 197 
<< m1 >>
rect 55 196 56 197 
<< m2 >>
rect 55 196 56 197 
<< m1 >>
rect 59 196 60 197 
<< m1 >>
rect 64 196 65 197 
<< pdiffusion >>
rect 66 196 67 197 
<< pdiffusion >>
rect 67 196 68 197 
<< pdiffusion >>
rect 68 196 69 197 
<< pdiffusion >>
rect 69 196 70 197 
<< pdiffusion >>
rect 70 196 71 197 
<< pdiffusion >>
rect 71 196 72 197 
<< m1 >>
rect 82 196 83 197 
<< pdiffusion >>
rect 84 196 85 197 
<< pdiffusion >>
rect 85 196 86 197 
<< pdiffusion >>
rect 86 196 87 197 
<< pdiffusion >>
rect 87 196 88 197 
<< pdiffusion >>
rect 88 196 89 197 
<< pdiffusion >>
rect 89 196 90 197 
<< m1 >>
rect 91 196 92 197 
<< m2 >>
rect 91 196 92 197 
<< m1 >>
rect 93 196 94 197 
<< m2 >>
rect 93 196 94 197 
<< pdiffusion >>
rect 102 196 103 197 
<< pdiffusion >>
rect 103 196 104 197 
<< pdiffusion >>
rect 104 196 105 197 
<< pdiffusion >>
rect 105 196 106 197 
<< pdiffusion >>
rect 106 196 107 197 
<< pdiffusion >>
rect 107 196 108 197 
<< m1 >>
rect 113 196 114 197 
<< m1 >>
rect 115 196 116 197 
<< pdiffusion >>
rect 120 196 121 197 
<< pdiffusion >>
rect 121 196 122 197 
<< pdiffusion >>
rect 122 196 123 197 
<< pdiffusion >>
rect 123 196 124 197 
<< pdiffusion >>
rect 124 196 125 197 
<< pdiffusion >>
rect 125 196 126 197 
<< m1 >>
rect 127 196 128 197 
<< m1 >>
rect 129 196 130 197 
<< m1 >>
rect 136 196 137 197 
<< pdiffusion >>
rect 138 196 139 197 
<< pdiffusion >>
rect 139 196 140 197 
<< pdiffusion >>
rect 140 196 141 197 
<< pdiffusion >>
rect 141 196 142 197 
<< pdiffusion >>
rect 142 196 143 197 
<< pdiffusion >>
rect 143 196 144 197 
<< m1 >>
rect 150 196 151 197 
<< m1 >>
rect 154 196 155 197 
<< pdiffusion >>
rect 156 196 157 197 
<< pdiffusion >>
rect 157 196 158 197 
<< pdiffusion >>
rect 158 196 159 197 
<< pdiffusion >>
rect 159 196 160 197 
<< pdiffusion >>
rect 160 196 161 197 
<< pdiffusion >>
rect 161 196 162 197 
<< m1 >>
rect 163 196 164 197 
<< m1 >>
rect 167 196 168 197 
<< m2 >>
rect 167 196 168 197 
<< pdiffusion >>
rect 174 196 175 197 
<< pdiffusion >>
rect 175 196 176 197 
<< pdiffusion >>
rect 176 196 177 197 
<< pdiffusion >>
rect 177 196 178 197 
<< pdiffusion >>
rect 178 196 179 197 
<< pdiffusion >>
rect 179 196 180 197 
<< m1 >>
rect 181 196 182 197 
<< m2 >>
rect 182 196 183 197 
<< m1 >>
rect 187 196 188 197 
<< pdiffusion >>
rect 192 196 193 197 
<< pdiffusion >>
rect 193 196 194 197 
<< pdiffusion >>
rect 194 196 195 197 
<< pdiffusion >>
rect 195 196 196 197 
<< pdiffusion >>
rect 196 196 197 197 
<< pdiffusion >>
rect 197 196 198 197 
<< m1 >>
rect 199 196 200 197 
<< pdiffusion >>
rect 210 196 211 197 
<< pdiffusion >>
rect 211 196 212 197 
<< pdiffusion >>
rect 212 196 213 197 
<< pdiffusion >>
rect 213 196 214 197 
<< pdiffusion >>
rect 214 196 215 197 
<< pdiffusion >>
rect 215 196 216 197 
<< pdiffusion >>
rect 228 196 229 197 
<< pdiffusion >>
rect 229 196 230 197 
<< pdiffusion >>
rect 230 196 231 197 
<< pdiffusion >>
rect 231 196 232 197 
<< pdiffusion >>
rect 232 196 233 197 
<< pdiffusion >>
rect 233 196 234 197 
<< pdiffusion >>
rect 246 196 247 197 
<< pdiffusion >>
rect 247 196 248 197 
<< pdiffusion >>
rect 248 196 249 197 
<< pdiffusion >>
rect 249 196 250 197 
<< pdiffusion >>
rect 250 196 251 197 
<< pdiffusion >>
rect 251 196 252 197 
<< m1 >>
rect 256 196 257 197 
<< pdiffusion >>
rect 12 197 13 198 
<< m1 >>
rect 13 197 14 198 
<< pdiffusion >>
rect 13 197 14 198 
<< pdiffusion >>
rect 14 197 15 198 
<< pdiffusion >>
rect 15 197 16 198 
<< pdiffusion >>
rect 16 197 17 198 
<< pdiffusion >>
rect 17 197 18 198 
<< m1 >>
rect 19 197 20 198 
<< m1 >>
rect 28 197 29 198 
<< m2 >>
rect 28 197 29 198 
<< pdiffusion >>
rect 30 197 31 198 
<< pdiffusion >>
rect 31 197 32 198 
<< pdiffusion >>
rect 32 197 33 198 
<< pdiffusion >>
rect 33 197 34 198 
<< m1 >>
rect 34 197 35 198 
<< pdiffusion >>
rect 34 197 35 198 
<< pdiffusion >>
rect 35 197 36 198 
<< m1 >>
rect 46 197 47 198 
<< m2 >>
rect 46 197 47 198 
<< pdiffusion >>
rect 48 197 49 198 
<< pdiffusion >>
rect 49 197 50 198 
<< pdiffusion >>
rect 50 197 51 198 
<< pdiffusion >>
rect 51 197 52 198 
<< pdiffusion >>
rect 52 197 53 198 
<< pdiffusion >>
rect 53 197 54 198 
<< m1 >>
rect 55 197 56 198 
<< m2 >>
rect 55 197 56 198 
<< m1 >>
rect 59 197 60 198 
<< m1 >>
rect 64 197 65 198 
<< pdiffusion >>
rect 66 197 67 198 
<< m1 >>
rect 67 197 68 198 
<< pdiffusion >>
rect 67 197 68 198 
<< pdiffusion >>
rect 68 197 69 198 
<< pdiffusion >>
rect 69 197 70 198 
<< pdiffusion >>
rect 70 197 71 198 
<< pdiffusion >>
rect 71 197 72 198 
<< m1 >>
rect 82 197 83 198 
<< pdiffusion >>
rect 84 197 85 198 
<< pdiffusion >>
rect 85 197 86 198 
<< pdiffusion >>
rect 86 197 87 198 
<< pdiffusion >>
rect 87 197 88 198 
<< m1 >>
rect 88 197 89 198 
<< pdiffusion >>
rect 88 197 89 198 
<< pdiffusion >>
rect 89 197 90 198 
<< m1 >>
rect 91 197 92 198 
<< m2 >>
rect 91 197 92 198 
<< m1 >>
rect 93 197 94 198 
<< m2 >>
rect 93 197 94 198 
<< pdiffusion >>
rect 102 197 103 198 
<< m1 >>
rect 103 197 104 198 
<< pdiffusion >>
rect 103 197 104 198 
<< pdiffusion >>
rect 104 197 105 198 
<< pdiffusion >>
rect 105 197 106 198 
<< pdiffusion >>
rect 106 197 107 198 
<< pdiffusion >>
rect 107 197 108 198 
<< m1 >>
rect 113 197 114 198 
<< m1 >>
rect 115 197 116 198 
<< pdiffusion >>
rect 120 197 121 198 
<< pdiffusion >>
rect 121 197 122 198 
<< pdiffusion >>
rect 122 197 123 198 
<< pdiffusion >>
rect 123 197 124 198 
<< pdiffusion >>
rect 124 197 125 198 
<< pdiffusion >>
rect 125 197 126 198 
<< m1 >>
rect 127 197 128 198 
<< m1 >>
rect 129 197 130 198 
<< m1 >>
rect 136 197 137 198 
<< pdiffusion >>
rect 138 197 139 198 
<< pdiffusion >>
rect 139 197 140 198 
<< pdiffusion >>
rect 140 197 141 198 
<< pdiffusion >>
rect 141 197 142 198 
<< pdiffusion >>
rect 142 197 143 198 
<< pdiffusion >>
rect 143 197 144 198 
<< m1 >>
rect 150 197 151 198 
<< m1 >>
rect 154 197 155 198 
<< pdiffusion >>
rect 156 197 157 198 
<< pdiffusion >>
rect 157 197 158 198 
<< pdiffusion >>
rect 158 197 159 198 
<< pdiffusion >>
rect 159 197 160 198 
<< m1 >>
rect 160 197 161 198 
<< pdiffusion >>
rect 160 197 161 198 
<< pdiffusion >>
rect 161 197 162 198 
<< m1 >>
rect 163 197 164 198 
<< m1 >>
rect 167 197 168 198 
<< m2 >>
rect 167 197 168 198 
<< pdiffusion >>
rect 174 197 175 198 
<< pdiffusion >>
rect 175 197 176 198 
<< pdiffusion >>
rect 176 197 177 198 
<< pdiffusion >>
rect 177 197 178 198 
<< pdiffusion >>
rect 178 197 179 198 
<< pdiffusion >>
rect 179 197 180 198 
<< m1 >>
rect 181 197 182 198 
<< m2 >>
rect 182 197 183 198 
<< m1 >>
rect 187 197 188 198 
<< pdiffusion >>
rect 192 197 193 198 
<< pdiffusion >>
rect 193 197 194 198 
<< pdiffusion >>
rect 194 197 195 198 
<< pdiffusion >>
rect 195 197 196 198 
<< pdiffusion >>
rect 196 197 197 198 
<< pdiffusion >>
rect 197 197 198 198 
<< m1 >>
rect 199 197 200 198 
<< pdiffusion >>
rect 210 197 211 198 
<< pdiffusion >>
rect 211 197 212 198 
<< pdiffusion >>
rect 212 197 213 198 
<< pdiffusion >>
rect 213 197 214 198 
<< pdiffusion >>
rect 214 197 215 198 
<< pdiffusion >>
rect 215 197 216 198 
<< pdiffusion >>
rect 228 197 229 198 
<< pdiffusion >>
rect 229 197 230 198 
<< pdiffusion >>
rect 230 197 231 198 
<< pdiffusion >>
rect 231 197 232 198 
<< m1 >>
rect 232 197 233 198 
<< pdiffusion >>
rect 232 197 233 198 
<< pdiffusion >>
rect 233 197 234 198 
<< pdiffusion >>
rect 246 197 247 198 
<< pdiffusion >>
rect 247 197 248 198 
<< pdiffusion >>
rect 248 197 249 198 
<< pdiffusion >>
rect 249 197 250 198 
<< pdiffusion >>
rect 250 197 251 198 
<< pdiffusion >>
rect 251 197 252 198 
<< m1 >>
rect 256 197 257 198 
<< m1 >>
rect 13 198 14 199 
<< m1 >>
rect 19 198 20 199 
<< m1 >>
rect 28 198 29 199 
<< m2 >>
rect 28 198 29 199 
<< m1 >>
rect 34 198 35 199 
<< m1 >>
rect 46 198 47 199 
<< m2 >>
rect 46 198 47 199 
<< m1 >>
rect 55 198 56 199 
<< m2 >>
rect 55 198 56 199 
<< m1 >>
rect 59 198 60 199 
<< m1 >>
rect 64 198 65 199 
<< m1 >>
rect 67 198 68 199 
<< m1 >>
rect 82 198 83 199 
<< m1 >>
rect 88 198 89 199 
<< m1 >>
rect 91 198 92 199 
<< m2 >>
rect 91 198 92 199 
<< m1 >>
rect 93 198 94 199 
<< m2 >>
rect 93 198 94 199 
<< m1 >>
rect 103 198 104 199 
<< m1 >>
rect 109 198 110 199 
<< m1 >>
rect 110 198 111 199 
<< m1 >>
rect 111 198 112 199 
<< m2 >>
rect 111 198 112 199 
<< m2c >>
rect 111 198 112 199 
<< m1 >>
rect 111 198 112 199 
<< m2 >>
rect 111 198 112 199 
<< m2 >>
rect 112 198 113 199 
<< m1 >>
rect 113 198 114 199 
<< m2 >>
rect 113 198 114 199 
<< m2 >>
rect 114 198 115 199 
<< m1 >>
rect 115 198 116 199 
<< m2 >>
rect 115 198 116 199 
<< m2c >>
rect 115 198 116 199 
<< m1 >>
rect 115 198 116 199 
<< m2 >>
rect 115 198 116 199 
<< m1 >>
rect 127 198 128 199 
<< m1 >>
rect 129 198 130 199 
<< m1 >>
rect 136 198 137 199 
<< m1 >>
rect 150 198 151 199 
<< m1 >>
rect 154 198 155 199 
<< m1 >>
rect 160 198 161 199 
<< m1 >>
rect 163 198 164 199 
<< m1 >>
rect 165 198 166 199 
<< m2 >>
rect 165 198 166 199 
<< m2 >>
rect 166 198 167 199 
<< m1 >>
rect 167 198 168 199 
<< m2 >>
rect 167 198 168 199 
<< m1 >>
rect 181 198 182 199 
<< m2 >>
rect 182 198 183 199 
<< m1 >>
rect 187 198 188 199 
<< m1 >>
rect 199 198 200 199 
<< m1 >>
rect 232 198 233 199 
<< m1 >>
rect 256 198 257 199 
<< m1 >>
rect 13 199 14 200 
<< m1 >>
rect 19 199 20 200 
<< m1 >>
rect 28 199 29 200 
<< m2 >>
rect 28 199 29 200 
<< m2 >>
rect 29 199 30 200 
<< m1 >>
rect 30 199 31 200 
<< m2 >>
rect 30 199 31 200 
<< m2c >>
rect 30 199 31 200 
<< m1 >>
rect 30 199 31 200 
<< m2 >>
rect 30 199 31 200 
<< m1 >>
rect 34 199 35 200 
<< m1 >>
rect 46 199 47 200 
<< m2 >>
rect 46 199 47 200 
<< m1 >>
rect 55 199 56 200 
<< m2 >>
rect 55 199 56 200 
<< m1 >>
rect 59 199 60 200 
<< m1 >>
rect 64 199 65 200 
<< m1 >>
rect 65 199 66 200 
<< m1 >>
rect 66 199 67 200 
<< m1 >>
rect 67 199 68 200 
<< m1 >>
rect 82 199 83 200 
<< m1 >>
rect 88 199 89 200 
<< m1 >>
rect 91 199 92 200 
<< m2 >>
rect 91 199 92 200 
<< m1 >>
rect 93 199 94 200 
<< m2 >>
rect 93 199 94 200 
<< m1 >>
rect 94 199 95 200 
<< m1 >>
rect 95 199 96 200 
<< m1 >>
rect 96 199 97 200 
<< m1 >>
rect 97 199 98 200 
<< m1 >>
rect 98 199 99 200 
<< m1 >>
rect 99 199 100 200 
<< m1 >>
rect 100 199 101 200 
<< m1 >>
rect 101 199 102 200 
<< m1 >>
rect 102 199 103 200 
<< m1 >>
rect 103 199 104 200 
<< m1 >>
rect 109 199 110 200 
<< m1 >>
rect 113 199 114 200 
<< m1 >>
rect 127 199 128 200 
<< m1 >>
rect 129 199 130 200 
<< m1 >>
rect 136 199 137 200 
<< m1 >>
rect 150 199 151 200 
<< m1 >>
rect 154 199 155 200 
<< m1 >>
rect 160 199 161 200 
<< m1 >>
rect 161 199 162 200 
<< m2 >>
rect 161 199 162 200 
<< m2c >>
rect 161 199 162 200 
<< m1 >>
rect 161 199 162 200 
<< m2 >>
rect 161 199 162 200 
<< m2 >>
rect 162 199 163 200 
<< m1 >>
rect 163 199 164 200 
<< m2 >>
rect 163 199 164 200 
<< m2 >>
rect 164 199 165 200 
<< m1 >>
rect 165 199 166 200 
<< m2 >>
rect 165 199 166 200 
<< m2c >>
rect 165 199 166 200 
<< m1 >>
rect 165 199 166 200 
<< m2 >>
rect 165 199 166 200 
<< m1 >>
rect 167 199 168 200 
<< m1 >>
rect 179 199 180 200 
<< m2 >>
rect 179 199 180 200 
<< m2c >>
rect 179 199 180 200 
<< m1 >>
rect 179 199 180 200 
<< m2 >>
rect 179 199 180 200 
<< m2 >>
rect 180 199 181 200 
<< m1 >>
rect 181 199 182 200 
<< m2 >>
rect 181 199 182 200 
<< m2 >>
rect 182 199 183 200 
<< m1 >>
rect 187 199 188 200 
<< m1 >>
rect 199 199 200 200 
<< m1 >>
rect 232 199 233 200 
<< m1 >>
rect 256 199 257 200 
<< m1 >>
rect 13 200 14 201 
<< m1 >>
rect 19 200 20 201 
<< m1 >>
rect 28 200 29 201 
<< m1 >>
rect 30 200 31 201 
<< m1 >>
rect 34 200 35 201 
<< m1 >>
rect 46 200 47 201 
<< m2 >>
rect 46 200 47 201 
<< m1 >>
rect 55 200 56 201 
<< m2 >>
rect 55 200 56 201 
<< m1 >>
rect 59 200 60 201 
<< m1 >>
rect 82 200 83 201 
<< m1 >>
rect 88 200 89 201 
<< m1 >>
rect 91 200 92 201 
<< m2 >>
rect 91 200 92 201 
<< m2 >>
rect 93 200 94 201 
<< m2 >>
rect 104 200 105 201 
<< m1 >>
rect 105 200 106 201 
<< m2 >>
rect 105 200 106 201 
<< m2c >>
rect 105 200 106 201 
<< m1 >>
rect 105 200 106 201 
<< m2 >>
rect 105 200 106 201 
<< m1 >>
rect 106 200 107 201 
<< m1 >>
rect 107 200 108 201 
<< m1 >>
rect 108 200 109 201 
<< m1 >>
rect 109 200 110 201 
<< m1 >>
rect 113 200 114 201 
<< m2 >>
rect 113 200 114 201 
<< m2c >>
rect 113 200 114 201 
<< m1 >>
rect 113 200 114 201 
<< m2 >>
rect 113 200 114 201 
<< m1 >>
rect 127 200 128 201 
<< m1 >>
rect 129 200 130 201 
<< m1 >>
rect 136 200 137 201 
<< m2 >>
rect 136 200 137 201 
<< m2c >>
rect 136 200 137 201 
<< m1 >>
rect 136 200 137 201 
<< m2 >>
rect 136 200 137 201 
<< m1 >>
rect 150 200 151 201 
<< m2 >>
rect 150 200 151 201 
<< m2c >>
rect 150 200 151 201 
<< m1 >>
rect 150 200 151 201 
<< m2 >>
rect 150 200 151 201 
<< m1 >>
rect 154 200 155 201 
<< m1 >>
rect 163 200 164 201 
<< m1 >>
rect 167 200 168 201 
<< m2 >>
rect 167 200 168 201 
<< m2c >>
rect 167 200 168 201 
<< m1 >>
rect 167 200 168 201 
<< m2 >>
rect 167 200 168 201 
<< m1 >>
rect 179 200 180 201 
<< m1 >>
rect 181 200 182 201 
<< m1 >>
rect 183 200 184 201 
<< m2 >>
rect 183 200 184 201 
<< m2c >>
rect 183 200 184 201 
<< m1 >>
rect 183 200 184 201 
<< m2 >>
rect 183 200 184 201 
<< m1 >>
rect 184 200 185 201 
<< m1 >>
rect 185 200 186 201 
<< m1 >>
rect 186 200 187 201 
<< m1 >>
rect 187 200 188 201 
<< m1 >>
rect 194 200 195 201 
<< m2 >>
rect 194 200 195 201 
<< m2c >>
rect 194 200 195 201 
<< m1 >>
rect 194 200 195 201 
<< m2 >>
rect 194 200 195 201 
<< m1 >>
rect 195 200 196 201 
<< m1 >>
rect 196 200 197 201 
<< m1 >>
rect 197 200 198 201 
<< m1 >>
rect 198 200 199 201 
<< m1 >>
rect 199 200 200 201 
<< m1 >>
rect 232 200 233 201 
<< m1 >>
rect 256 200 257 201 
<< m1 >>
rect 13 201 14 202 
<< m1 >>
rect 19 201 20 202 
<< m1 >>
rect 28 201 29 202 
<< m1 >>
rect 30 201 31 202 
<< m1 >>
rect 34 201 35 202 
<< m1 >>
rect 46 201 47 202 
<< m2 >>
rect 46 201 47 202 
<< m1 >>
rect 55 201 56 202 
<< m2 >>
rect 55 201 56 202 
<< m1 >>
rect 59 201 60 202 
<< m1 >>
rect 82 201 83 202 
<< m2 >>
rect 87 201 88 202 
<< m1 >>
rect 88 201 89 202 
<< m2 >>
rect 88 201 89 202 
<< m2c >>
rect 88 201 89 202 
<< m1 >>
rect 88 201 89 202 
<< m2 >>
rect 88 201 89 202 
<< m1 >>
rect 91 201 92 202 
<< m2 >>
rect 91 201 92 202 
<< m2 >>
rect 93 201 94 202 
<< m2 >>
rect 104 201 105 202 
<< m2 >>
rect 113 201 114 202 
<< m1 >>
rect 127 201 128 202 
<< m1 >>
rect 129 201 130 202 
<< m2 >>
rect 136 201 137 202 
<< m2 >>
rect 150 201 151 202 
<< m1 >>
rect 154 201 155 202 
<< m1 >>
rect 163 201 164 202 
<< m2 >>
rect 167 201 168 202 
<< m1 >>
rect 179 201 180 202 
<< m1 >>
rect 181 201 182 202 
<< m2 >>
rect 183 201 184 202 
<< m2 >>
rect 194 201 195 202 
<< m1 >>
rect 232 201 233 202 
<< m1 >>
rect 256 201 257 202 
<< m1 >>
rect 13 202 14 203 
<< m1 >>
rect 19 202 20 203 
<< m1 >>
rect 28 202 29 203 
<< m1 >>
rect 30 202 31 203 
<< m1 >>
rect 31 202 32 203 
<< m1 >>
rect 32 202 33 203 
<< m1 >>
rect 33 202 34 203 
<< m1 >>
rect 34 202 35 203 
<< m1 >>
rect 46 202 47 203 
<< m2 >>
rect 46 202 47 203 
<< m1 >>
rect 55 202 56 203 
<< m2 >>
rect 55 202 56 203 
<< m1 >>
rect 59 202 60 203 
<< m1 >>
rect 60 202 61 203 
<< m1 >>
rect 61 202 62 203 
<< m1 >>
rect 62 202 63 203 
<< m1 >>
rect 63 202 64 203 
<< m1 >>
rect 64 202 65 203 
<< m1 >>
rect 65 202 66 203 
<< m1 >>
rect 66 202 67 203 
<< m1 >>
rect 67 202 68 203 
<< m1 >>
rect 68 202 69 203 
<< m1 >>
rect 69 202 70 203 
<< m1 >>
rect 70 202 71 203 
<< m1 >>
rect 71 202 72 203 
<< m1 >>
rect 72 202 73 203 
<< m1 >>
rect 73 202 74 203 
<< m1 >>
rect 74 202 75 203 
<< m1 >>
rect 75 202 76 203 
<< m1 >>
rect 76 202 77 203 
<< m1 >>
rect 77 202 78 203 
<< m1 >>
rect 78 202 79 203 
<< m1 >>
rect 79 202 80 203 
<< m1 >>
rect 80 202 81 203 
<< m2 >>
rect 80 202 81 203 
<< m2c >>
rect 80 202 81 203 
<< m1 >>
rect 80 202 81 203 
<< m2 >>
rect 80 202 81 203 
<< m2 >>
rect 81 202 82 203 
<< m1 >>
rect 82 202 83 203 
<< m2 >>
rect 82 202 83 203 
<< m2 >>
rect 83 202 84 203 
<< m1 >>
rect 84 202 85 203 
<< m2 >>
rect 84 202 85 203 
<< m2c >>
rect 84 202 85 203 
<< m1 >>
rect 84 202 85 203 
<< m2 >>
rect 84 202 85 203 
<< m1 >>
rect 85 202 86 203 
<< m1 >>
rect 86 202 87 203 
<< m2 >>
rect 87 202 88 203 
<< m1 >>
rect 91 202 92 203 
<< m2 >>
rect 91 202 92 203 
<< m1 >>
rect 92 202 93 203 
<< m1 >>
rect 93 202 94 203 
<< m2 >>
rect 93 202 94 203 
<< m1 >>
rect 94 202 95 203 
<< m1 >>
rect 95 202 96 203 
<< m1 >>
rect 96 202 97 203 
<< m1 >>
rect 97 202 98 203 
<< m1 >>
rect 98 202 99 203 
<< m1 >>
rect 99 202 100 203 
<< m1 >>
rect 100 202 101 203 
<< m1 >>
rect 101 202 102 203 
<< m1 >>
rect 102 202 103 203 
<< m1 >>
rect 103 202 104 203 
<< m1 >>
rect 104 202 105 203 
<< m2 >>
rect 104 202 105 203 
<< m1 >>
rect 105 202 106 203 
<< m1 >>
rect 106 202 107 203 
<< m1 >>
rect 107 202 108 203 
<< m1 >>
rect 108 202 109 203 
<< m1 >>
rect 109 202 110 203 
<< m1 >>
rect 110 202 111 203 
<< m1 >>
rect 111 202 112 203 
<< m1 >>
rect 112 202 113 203 
<< m1 >>
rect 113 202 114 203 
<< m2 >>
rect 113 202 114 203 
<< m1 >>
rect 114 202 115 203 
<< m1 >>
rect 115 202 116 203 
<< m1 >>
rect 116 202 117 203 
<< m1 >>
rect 117 202 118 203 
<< m1 >>
rect 118 202 119 203 
<< m1 >>
rect 119 202 120 203 
<< m1 >>
rect 120 202 121 203 
<< m1 >>
rect 121 202 122 203 
<< m1 >>
rect 127 202 128 203 
<< m1 >>
rect 129 202 130 203 
<< m1 >>
rect 130 202 131 203 
<< m1 >>
rect 131 202 132 203 
<< m1 >>
rect 132 202 133 203 
<< m1 >>
rect 133 202 134 203 
<< m1 >>
rect 134 202 135 203 
<< m1 >>
rect 135 202 136 203 
<< m1 >>
rect 136 202 137 203 
<< m2 >>
rect 136 202 137 203 
<< m1 >>
rect 137 202 138 203 
<< m1 >>
rect 138 202 139 203 
<< m1 >>
rect 139 202 140 203 
<< m1 >>
rect 140 202 141 203 
<< m1 >>
rect 141 202 142 203 
<< m1 >>
rect 142 202 143 203 
<< m1 >>
rect 143 202 144 203 
<< m1 >>
rect 144 202 145 203 
<< m1 >>
rect 145 202 146 203 
<< m1 >>
rect 146 202 147 203 
<< m1 >>
rect 147 202 148 203 
<< m1 >>
rect 148 202 149 203 
<< m1 >>
rect 149 202 150 203 
<< m1 >>
rect 150 202 151 203 
<< m2 >>
rect 150 202 151 203 
<< m1 >>
rect 151 202 152 203 
<< m1 >>
rect 152 202 153 203 
<< m2 >>
rect 152 202 153 203 
<< m2c >>
rect 152 202 153 203 
<< m1 >>
rect 152 202 153 203 
<< m2 >>
rect 152 202 153 203 
<< m2 >>
rect 153 202 154 203 
<< m1 >>
rect 154 202 155 203 
<< m2 >>
rect 154 202 155 203 
<< m2 >>
rect 155 202 156 203 
<< m1 >>
rect 156 202 157 203 
<< m2 >>
rect 156 202 157 203 
<< m2c >>
rect 156 202 157 203 
<< m1 >>
rect 156 202 157 203 
<< m2 >>
rect 156 202 157 203 
<< m1 >>
rect 157 202 158 203 
<< m1 >>
rect 158 202 159 203 
<< m1 >>
rect 159 202 160 203 
<< m1 >>
rect 160 202 161 203 
<< m1 >>
rect 161 202 162 203 
<< m2 >>
rect 161 202 162 203 
<< m1 >>
rect 162 202 163 203 
<< m2 >>
rect 162 202 163 203 
<< m1 >>
rect 163 202 164 203 
<< m2 >>
rect 163 202 164 203 
<< m2 >>
rect 164 202 165 203 
<< m1 >>
rect 165 202 166 203 
<< m2 >>
rect 165 202 166 203 
<< m2c >>
rect 165 202 166 203 
<< m1 >>
rect 165 202 166 203 
<< m2 >>
rect 165 202 166 203 
<< m1 >>
rect 166 202 167 203 
<< m1 >>
rect 167 202 168 203 
<< m2 >>
rect 167 202 168 203 
<< m1 >>
rect 168 202 169 203 
<< m2 >>
rect 168 202 169 203 
<< m1 >>
rect 169 202 170 203 
<< m2 >>
rect 169 202 170 203 
<< m1 >>
rect 170 202 171 203 
<< m2 >>
rect 170 202 171 203 
<< m1 >>
rect 171 202 172 203 
<< m2 >>
rect 171 202 172 203 
<< m1 >>
rect 172 202 173 203 
<< m2 >>
rect 172 202 173 203 
<< m1 >>
rect 173 202 174 203 
<< m2 >>
rect 173 202 174 203 
<< m1 >>
rect 174 202 175 203 
<< m2 >>
rect 174 202 175 203 
<< m1 >>
rect 175 202 176 203 
<< m2 >>
rect 175 202 176 203 
<< m1 >>
rect 176 202 177 203 
<< m2 >>
rect 176 202 177 203 
<< m1 >>
rect 177 202 178 203 
<< m2 >>
rect 177 202 178 203 
<< m1 >>
rect 178 202 179 203 
<< m2 >>
rect 178 202 179 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m2 >>
rect 180 202 181 203 
<< m1 >>
rect 181 202 182 203 
<< m2 >>
rect 181 202 182 203 
<< m1 >>
rect 182 202 183 203 
<< m2 >>
rect 182 202 183 203 
<< m1 >>
rect 183 202 184 203 
<< m2 >>
rect 183 202 184 203 
<< m1 >>
rect 184 202 185 203 
<< m1 >>
rect 185 202 186 203 
<< m1 >>
rect 186 202 187 203 
<< m1 >>
rect 187 202 188 203 
<< m1 >>
rect 188 202 189 203 
<< m1 >>
rect 189 202 190 203 
<< m1 >>
rect 190 202 191 203 
<< m1 >>
rect 191 202 192 203 
<< m1 >>
rect 192 202 193 203 
<< m1 >>
rect 193 202 194 203 
<< m1 >>
rect 194 202 195 203 
<< m2 >>
rect 194 202 195 203 
<< m1 >>
rect 195 202 196 203 
<< m1 >>
rect 196 202 197 203 
<< m1 >>
rect 197 202 198 203 
<< m1 >>
rect 198 202 199 203 
<< m1 >>
rect 199 202 200 203 
<< m1 >>
rect 200 202 201 203 
<< m1 >>
rect 201 202 202 203 
<< m1 >>
rect 202 202 203 203 
<< m1 >>
rect 203 202 204 203 
<< m1 >>
rect 204 202 205 203 
<< m1 >>
rect 205 202 206 203 
<< m1 >>
rect 206 202 207 203 
<< m1 >>
rect 207 202 208 203 
<< m1 >>
rect 208 202 209 203 
<< m1 >>
rect 209 202 210 203 
<< m1 >>
rect 210 202 211 203 
<< m1 >>
rect 211 202 212 203 
<< m1 >>
rect 212 202 213 203 
<< m1 >>
rect 213 202 214 203 
<< m1 >>
rect 214 202 215 203 
<< m1 >>
rect 215 202 216 203 
<< m1 >>
rect 216 202 217 203 
<< m1 >>
rect 217 202 218 203 
<< m1 >>
rect 218 202 219 203 
<< m1 >>
rect 219 202 220 203 
<< m1 >>
rect 220 202 221 203 
<< m1 >>
rect 221 202 222 203 
<< m1 >>
rect 222 202 223 203 
<< m1 >>
rect 223 202 224 203 
<< m1 >>
rect 224 202 225 203 
<< m1 >>
rect 225 202 226 203 
<< m1 >>
rect 226 202 227 203 
<< m1 >>
rect 227 202 228 203 
<< m1 >>
rect 228 202 229 203 
<< m1 >>
rect 229 202 230 203 
<< m1 >>
rect 230 202 231 203 
<< m1 >>
rect 231 202 232 203 
<< m1 >>
rect 232 202 233 203 
<< m1 >>
rect 256 202 257 203 
<< m1 >>
rect 13 203 14 204 
<< m1 >>
rect 19 203 20 204 
<< m1 >>
rect 28 203 29 204 
<< m1 >>
rect 46 203 47 204 
<< m2 >>
rect 46 203 47 204 
<< m1 >>
rect 55 203 56 204 
<< m2 >>
rect 55 203 56 204 
<< m1 >>
rect 82 203 83 204 
<< m1 >>
rect 86 203 87 204 
<< m2 >>
rect 87 203 88 204 
<< m2 >>
rect 90 203 91 204 
<< m2 >>
rect 91 203 92 204 
<< m2 >>
rect 93 203 94 204 
<< m2 >>
rect 104 203 105 204 
<< m2 >>
rect 113 203 114 204 
<< m1 >>
rect 121 203 122 204 
<< m1 >>
rect 127 203 128 204 
<< m2 >>
rect 136 203 137 204 
<< m2 >>
rect 150 203 151 204 
<< m1 >>
rect 154 203 155 204 
<< m2 >>
rect 161 203 162 204 
<< m2 >>
rect 194 203 195 204 
<< m1 >>
rect 256 203 257 204 
<< m1 >>
rect 13 204 14 205 
<< m1 >>
rect 19 204 20 205 
<< m1 >>
rect 28 204 29 205 
<< m1 >>
rect 46 204 47 205 
<< m2 >>
rect 46 204 47 205 
<< m1 >>
rect 55 204 56 205 
<< m2 >>
rect 55 204 56 205 
<< m1 >>
rect 80 204 81 205 
<< m2 >>
rect 80 204 81 205 
<< m2c >>
rect 80 204 81 205 
<< m1 >>
rect 80 204 81 205 
<< m2 >>
rect 80 204 81 205 
<< m2 >>
rect 81 204 82 205 
<< m1 >>
rect 82 204 83 205 
<< m2 >>
rect 82 204 83 205 
<< m2 >>
rect 83 204 84 205 
<< m1 >>
rect 84 204 85 205 
<< m2 >>
rect 84 204 85 205 
<< m2c >>
rect 84 204 85 205 
<< m1 >>
rect 84 204 85 205 
<< m2 >>
rect 84 204 85 205 
<< m2 >>
rect 85 204 86 205 
<< m1 >>
rect 86 204 87 205 
<< m2 >>
rect 86 204 87 205 
<< m2 >>
rect 87 204 88 205 
<< m1 >>
rect 90 204 91 205 
<< m2 >>
rect 90 204 91 205 
<< m2c >>
rect 90 204 91 205 
<< m1 >>
rect 90 204 91 205 
<< m2 >>
rect 90 204 91 205 
<< m1 >>
rect 93 204 94 205 
<< m2 >>
rect 93 204 94 205 
<< m2c >>
rect 93 204 94 205 
<< m1 >>
rect 93 204 94 205 
<< m2 >>
rect 93 204 94 205 
<< m2 >>
rect 104 204 105 205 
<< m1 >>
rect 113 204 114 205 
<< m2 >>
rect 113 204 114 205 
<< m2c >>
rect 113 204 114 205 
<< m1 >>
rect 113 204 114 205 
<< m2 >>
rect 113 204 114 205 
<< m1 >>
rect 121 204 122 205 
<< m1 >>
rect 127 204 128 205 
<< m1 >>
rect 136 204 137 205 
<< m2 >>
rect 136 204 137 205 
<< m2c >>
rect 136 204 137 205 
<< m1 >>
rect 136 204 137 205 
<< m2 >>
rect 136 204 137 205 
<< m1 >>
rect 137 204 138 205 
<< m1 >>
rect 138 204 139 205 
<< m1 >>
rect 139 204 140 205 
<< m1 >>
rect 140 204 141 205 
<< m1 >>
rect 150 204 151 205 
<< m2 >>
rect 150 204 151 205 
<< m2c >>
rect 150 204 151 205 
<< m1 >>
rect 150 204 151 205 
<< m2 >>
rect 150 204 151 205 
<< m1 >>
rect 154 204 155 205 
<< m2 >>
rect 156 204 157 205 
<< m2 >>
rect 157 204 158 205 
<< m2 >>
rect 158 204 159 205 
<< m2 >>
rect 159 204 160 205 
<< m2 >>
rect 160 204 161 205 
<< m2 >>
rect 161 204 162 205 
<< m1 >>
rect 163 204 164 205 
<< m1 >>
rect 164 204 165 205 
<< m1 >>
rect 165 204 166 205 
<< m1 >>
rect 166 204 167 205 
<< m1 >>
rect 167 204 168 205 
<< m1 >>
rect 168 204 169 205 
<< m1 >>
rect 169 204 170 205 
<< m1 >>
rect 170 204 171 205 
<< m1 >>
rect 171 204 172 205 
<< m1 >>
rect 172 204 173 205 
<< m1 >>
rect 173 204 174 205 
<< m1 >>
rect 174 204 175 205 
<< m1 >>
rect 175 204 176 205 
<< m1 >>
rect 176 204 177 205 
<< m1 >>
rect 177 204 178 205 
<< m1 >>
rect 178 204 179 205 
<< m1 >>
rect 179 204 180 205 
<< m1 >>
rect 180 204 181 205 
<< m1 >>
rect 181 204 182 205 
<< m1 >>
rect 182 204 183 205 
<< m1 >>
rect 183 204 184 205 
<< m1 >>
rect 184 204 185 205 
<< m1 >>
rect 185 204 186 205 
<< m1 >>
rect 186 204 187 205 
<< m1 >>
rect 187 204 188 205 
<< m1 >>
rect 188 204 189 205 
<< m1 >>
rect 189 204 190 205 
<< m1 >>
rect 190 204 191 205 
<< m2 >>
rect 190 204 191 205 
<< m2c >>
rect 190 204 191 205 
<< m1 >>
rect 190 204 191 205 
<< m2 >>
rect 190 204 191 205 
<< m2 >>
rect 191 204 192 205 
<< m1 >>
rect 192 204 193 205 
<< m2 >>
rect 192 204 193 205 
<< m1 >>
rect 193 204 194 205 
<< m2 >>
rect 193 204 194 205 
<< m1 >>
rect 194 204 195 205 
<< m2 >>
rect 194 204 195 205 
<< m1 >>
rect 195 204 196 205 
<< m1 >>
rect 196 204 197 205 
<< m1 >>
rect 197 204 198 205 
<< m1 >>
rect 198 204 199 205 
<< m1 >>
rect 199 204 200 205 
<< m1 >>
rect 200 204 201 205 
<< m1 >>
rect 201 204 202 205 
<< m1 >>
rect 202 204 203 205 
<< m1 >>
rect 203 204 204 205 
<< m1 >>
rect 204 204 205 205 
<< m1 >>
rect 205 204 206 205 
<< m1 >>
rect 206 204 207 205 
<< m1 >>
rect 207 204 208 205 
<< m1 >>
rect 208 204 209 205 
<< m1 >>
rect 209 204 210 205 
<< m1 >>
rect 210 204 211 205 
<< m1 >>
rect 211 204 212 205 
<< m1 >>
rect 212 204 213 205 
<< m1 >>
rect 213 204 214 205 
<< m1 >>
rect 214 204 215 205 
<< m1 >>
rect 215 204 216 205 
<< m1 >>
rect 216 204 217 205 
<< m1 >>
rect 217 204 218 205 
<< m1 >>
rect 218 204 219 205 
<< m1 >>
rect 219 204 220 205 
<< m1 >>
rect 220 204 221 205 
<< m1 >>
rect 221 204 222 205 
<< m1 >>
rect 222 204 223 205 
<< m1 >>
rect 223 204 224 205 
<< m1 >>
rect 224 204 225 205 
<< m1 >>
rect 225 204 226 205 
<< m1 >>
rect 226 204 227 205 
<< m1 >>
rect 227 204 228 205 
<< m1 >>
rect 228 204 229 205 
<< m1 >>
rect 229 204 230 205 
<< m1 >>
rect 230 204 231 205 
<< m1 >>
rect 231 204 232 205 
<< m1 >>
rect 232 204 233 205 
<< m1 >>
rect 233 204 234 205 
<< m1 >>
rect 234 204 235 205 
<< m1 >>
rect 235 204 236 205 
<< m1 >>
rect 236 204 237 205 
<< m1 >>
rect 237 204 238 205 
<< m1 >>
rect 238 204 239 205 
<< m1 >>
rect 239 204 240 205 
<< m1 >>
rect 240 204 241 205 
<< m1 >>
rect 241 204 242 205 
<< m1 >>
rect 242 204 243 205 
<< m1 >>
rect 243 204 244 205 
<< m1 >>
rect 244 204 245 205 
<< m1 >>
rect 245 204 246 205 
<< m1 >>
rect 246 204 247 205 
<< m1 >>
rect 247 204 248 205 
<< m1 >>
rect 248 204 249 205 
<< m1 >>
rect 249 204 250 205 
<< m1 >>
rect 250 204 251 205 
<< m1 >>
rect 251 204 252 205 
<< m1 >>
rect 252 204 253 205 
<< m1 >>
rect 253 204 254 205 
<< m1 >>
rect 254 204 255 205 
<< m1 >>
rect 255 204 256 205 
<< m1 >>
rect 256 204 257 205 
<< m1 >>
rect 13 205 14 206 
<< m1 >>
rect 14 205 15 206 
<< m1 >>
rect 15 205 16 206 
<< m1 >>
rect 16 205 17 206 
<< m1 >>
rect 17 205 18 206 
<< m1 >>
rect 19 205 20 206 
<< m1 >>
rect 28 205 29 206 
<< m1 >>
rect 46 205 47 206 
<< m2 >>
rect 46 205 47 206 
<< m1 >>
rect 55 205 56 206 
<< m2 >>
rect 55 205 56 206 
<< m1 >>
rect 80 205 81 206 
<< m1 >>
rect 82 205 83 206 
<< m1 >>
rect 86 205 87 206 
<< m1 >>
rect 90 205 91 206 
<< m1 >>
rect 93 205 94 206 
<< m1 >>
rect 95 205 96 206 
<< m2 >>
rect 95 205 96 206 
<< m1 >>
rect 96 205 97 206 
<< m2 >>
rect 96 205 97 206 
<< m1 >>
rect 97 205 98 206 
<< m2 >>
rect 97 205 98 206 
<< m1 >>
rect 98 205 99 206 
<< m2 >>
rect 98 205 99 206 
<< m1 >>
rect 99 205 100 206 
<< m2 >>
rect 99 205 100 206 
<< m1 >>
rect 100 205 101 206 
<< m2 >>
rect 100 205 101 206 
<< m1 >>
rect 101 205 102 206 
<< m2 >>
rect 101 205 102 206 
<< m1 >>
rect 102 205 103 206 
<< m2 >>
rect 102 205 103 206 
<< m1 >>
rect 103 205 104 206 
<< m2 >>
rect 103 205 104 206 
<< m1 >>
rect 104 205 105 206 
<< m2 >>
rect 104 205 105 206 
<< m1 >>
rect 105 205 106 206 
<< m1 >>
rect 106 205 107 206 
<< m1 >>
rect 113 205 114 206 
<< m1 >>
rect 121 205 122 206 
<< m1 >>
rect 127 205 128 206 
<< m1 >>
rect 140 205 141 206 
<< m1 >>
rect 150 205 151 206 
<< m1 >>
rect 154 205 155 206 
<< m1 >>
rect 155 205 156 206 
<< m1 >>
rect 156 205 157 206 
<< m2 >>
rect 156 205 157 206 
<< m1 >>
rect 157 205 158 206 
<< m1 >>
rect 158 205 159 206 
<< m1 >>
rect 159 205 160 206 
<< m1 >>
rect 160 205 161 206 
<< m1 >>
rect 163 205 164 206 
<< m1 >>
rect 192 205 193 206 
<< m1 >>
rect 17 206 18 207 
<< m1 >>
rect 19 206 20 207 
<< m1 >>
rect 28 206 29 207 
<< m1 >>
rect 46 206 47 207 
<< m2 >>
rect 46 206 47 207 
<< m1 >>
rect 55 206 56 207 
<< m2 >>
rect 55 206 56 207 
<< m1 >>
rect 80 206 81 207 
<< m1 >>
rect 82 206 83 207 
<< m1 >>
rect 86 206 87 207 
<< m1 >>
rect 87 206 88 207 
<< m1 >>
rect 88 206 89 207 
<< m2 >>
rect 88 206 89 207 
<< m2c >>
rect 88 206 89 207 
<< m1 >>
rect 88 206 89 207 
<< m2 >>
rect 88 206 89 207 
<< m2 >>
rect 89 206 90 207 
<< m1 >>
rect 90 206 91 207 
<< m2 >>
rect 90 206 91 207 
<< m2 >>
rect 91 206 92 207 
<< m2 >>
rect 92 206 93 207 
<< m1 >>
rect 93 206 94 207 
<< m2 >>
rect 93 206 94 207 
<< m2 >>
rect 94 206 95 207 
<< m1 >>
rect 95 206 96 207 
<< m2 >>
rect 95 206 96 207 
<< m1 >>
rect 106 206 107 207 
<< m1 >>
rect 113 206 114 207 
<< m1 >>
rect 121 206 122 207 
<< m1 >>
rect 127 206 128 207 
<< m1 >>
rect 140 206 141 207 
<< m1 >>
rect 141 206 142 207 
<< m1 >>
rect 142 206 143 207 
<< m1 >>
rect 143 206 144 207 
<< m1 >>
rect 144 206 145 207 
<< m1 >>
rect 145 206 146 207 
<< m1 >>
rect 146 206 147 207 
<< m1 >>
rect 147 206 148 207 
<< m1 >>
rect 148 206 149 207 
<< m2 >>
rect 148 206 149 207 
<< m2c >>
rect 148 206 149 207 
<< m1 >>
rect 148 206 149 207 
<< m2 >>
rect 148 206 149 207 
<< m2 >>
rect 149 206 150 207 
<< m1 >>
rect 150 206 151 207 
<< m2 >>
rect 150 206 151 207 
<< m2 >>
rect 151 206 152 207 
<< m1 >>
rect 152 206 153 207 
<< m2 >>
rect 152 206 153 207 
<< m2c >>
rect 152 206 153 207 
<< m1 >>
rect 152 206 153 207 
<< m2 >>
rect 152 206 153 207 
<< m2 >>
rect 156 206 157 207 
<< m1 >>
rect 160 206 161 207 
<< m1 >>
rect 163 206 164 207 
<< m2 >>
rect 190 206 191 207 
<< m2 >>
rect 191 206 192 207 
<< m1 >>
rect 192 206 193 207 
<< m2 >>
rect 192 206 193 207 
<< m2c >>
rect 192 206 193 207 
<< m1 >>
rect 192 206 193 207 
<< m2 >>
rect 192 206 193 207 
<< m1 >>
rect 17 207 18 208 
<< m1 >>
rect 19 207 20 208 
<< m1 >>
rect 28 207 29 208 
<< m1 >>
rect 46 207 47 208 
<< m2 >>
rect 46 207 47 208 
<< m1 >>
rect 55 207 56 208 
<< m2 >>
rect 55 207 56 208 
<< m2 >>
rect 74 207 75 208 
<< m1 >>
rect 75 207 76 208 
<< m2 >>
rect 75 207 76 208 
<< m2c >>
rect 75 207 76 208 
<< m1 >>
rect 75 207 76 208 
<< m2 >>
rect 75 207 76 208 
<< m1 >>
rect 76 207 77 208 
<< m1 >>
rect 77 207 78 208 
<< m1 >>
rect 78 207 79 208 
<< m1 >>
rect 79 207 80 208 
<< m1 >>
rect 80 207 81 208 
<< m1 >>
rect 82 207 83 208 
<< m1 >>
rect 90 207 91 208 
<< m1 >>
rect 93 207 94 208 
<< m1 >>
rect 95 207 96 208 
<< m1 >>
rect 106 207 107 208 
<< m1 >>
rect 113 207 114 208 
<< m1 >>
rect 121 207 122 208 
<< m1 >>
rect 127 207 128 208 
<< m1 >>
rect 150 207 151 208 
<< m1 >>
rect 152 207 153 208 
<< m1 >>
rect 154 207 155 208 
<< m1 >>
rect 155 207 156 208 
<< m1 >>
rect 156 207 157 208 
<< m2 >>
rect 156 207 157 208 
<< m2c >>
rect 156 207 157 208 
<< m1 >>
rect 156 207 157 208 
<< m2 >>
rect 156 207 157 208 
<< m1 >>
rect 160 207 161 208 
<< m1 >>
rect 163 207 164 208 
<< m1 >>
rect 175 207 176 208 
<< m1 >>
rect 176 207 177 208 
<< m1 >>
rect 177 207 178 208 
<< m1 >>
rect 178 207 179 208 
<< m1 >>
rect 179 207 180 208 
<< m1 >>
rect 180 207 181 208 
<< m1 >>
rect 181 207 182 208 
<< m1 >>
rect 182 207 183 208 
<< m1 >>
rect 183 207 184 208 
<< m1 >>
rect 184 207 185 208 
<< m1 >>
rect 185 207 186 208 
<< m1 >>
rect 186 207 187 208 
<< m1 >>
rect 187 207 188 208 
<< m1 >>
rect 188 207 189 208 
<< m1 >>
rect 189 207 190 208 
<< m1 >>
rect 190 207 191 208 
<< m2 >>
rect 190 207 191 208 
<< m1 >>
rect 17 208 18 209 
<< m2 >>
rect 17 208 18 209 
<< m2c >>
rect 17 208 18 209 
<< m1 >>
rect 17 208 18 209 
<< m2 >>
rect 17 208 18 209 
<< m2 >>
rect 18 208 19 209 
<< m1 >>
rect 19 208 20 209 
<< m2 >>
rect 19 208 20 209 
<< m2 >>
rect 20 208 21 209 
<< m1 >>
rect 28 208 29 209 
<< m1 >>
rect 46 208 47 209 
<< m2 >>
rect 46 208 47 209 
<< m1 >>
rect 55 208 56 209 
<< m2 >>
rect 55 208 56 209 
<< m1 >>
rect 70 208 71 209 
<< m1 >>
rect 71 208 72 209 
<< m1 >>
rect 72 208 73 209 
<< m1 >>
rect 73 208 74 209 
<< m2 >>
rect 74 208 75 209 
<< m1 >>
rect 82 208 83 209 
<< m1 >>
rect 88 208 89 209 
<< m1 >>
rect 89 208 90 209 
<< m1 >>
rect 90 208 91 209 
<< m1 >>
rect 93 208 94 209 
<< m1 >>
rect 95 208 96 209 
<< m1 >>
rect 106 208 107 209 
<< m1 >>
rect 113 208 114 209 
<< m1 >>
rect 121 208 122 209 
<< m1 >>
rect 124 208 125 209 
<< m1 >>
rect 125 208 126 209 
<< m1 >>
rect 126 208 127 209 
<< m1 >>
rect 127 208 128 209 
<< m1 >>
rect 150 208 151 209 
<< m1 >>
rect 152 208 153 209 
<< m1 >>
rect 154 208 155 209 
<< m1 >>
rect 160 208 161 209 
<< m1 >>
rect 163 208 164 209 
<< m1 >>
rect 175 208 176 209 
<< m1 >>
rect 190 208 191 209 
<< m2 >>
rect 190 208 191 209 
<< m1 >>
rect 208 208 209 209 
<< m1 >>
rect 209 208 210 209 
<< m1 >>
rect 210 208 211 209 
<< m1 >>
rect 211 208 212 209 
<< m1 >>
rect 19 209 20 210 
<< m2 >>
rect 20 209 21 210 
<< m1 >>
rect 28 209 29 210 
<< m1 >>
rect 46 209 47 210 
<< m2 >>
rect 46 209 47 210 
<< m1 >>
rect 55 209 56 210 
<< m2 >>
rect 55 209 56 210 
<< m1 >>
rect 70 209 71 210 
<< m1 >>
rect 73 209 74 210 
<< m2 >>
rect 74 209 75 210 
<< m1 >>
rect 82 209 83 210 
<< m1 >>
rect 88 209 89 210 
<< m1 >>
rect 93 209 94 210 
<< m1 >>
rect 95 209 96 210 
<< m1 >>
rect 106 209 107 210 
<< m1 >>
rect 113 209 114 210 
<< m1 >>
rect 121 209 122 210 
<< m1 >>
rect 124 209 125 210 
<< m1 >>
rect 150 209 151 210 
<< m1 >>
rect 152 209 153 210 
<< m1 >>
rect 154 209 155 210 
<< m1 >>
rect 160 209 161 210 
<< m1 >>
rect 163 209 164 210 
<< m1 >>
rect 175 209 176 210 
<< m1 >>
rect 188 209 189 210 
<< m2 >>
rect 188 209 189 210 
<< m2c >>
rect 188 209 189 210 
<< m1 >>
rect 188 209 189 210 
<< m2 >>
rect 188 209 189 210 
<< m2 >>
rect 189 209 190 210 
<< m1 >>
rect 190 209 191 210 
<< m2 >>
rect 190 209 191 210 
<< m1 >>
rect 208 209 209 210 
<< m1 >>
rect 211 209 212 210 
<< pdiffusion >>
rect 12 210 13 211 
<< pdiffusion >>
rect 13 210 14 211 
<< pdiffusion >>
rect 14 210 15 211 
<< pdiffusion >>
rect 15 210 16 211 
<< pdiffusion >>
rect 16 210 17 211 
<< pdiffusion >>
rect 17 210 18 211 
<< m1 >>
rect 19 210 20 211 
<< m2 >>
rect 20 210 21 211 
<< m1 >>
rect 28 210 29 211 
<< pdiffusion >>
rect 30 210 31 211 
<< pdiffusion >>
rect 31 210 32 211 
<< pdiffusion >>
rect 32 210 33 211 
<< pdiffusion >>
rect 33 210 34 211 
<< pdiffusion >>
rect 34 210 35 211 
<< pdiffusion >>
rect 35 210 36 211 
<< m1 >>
rect 46 210 47 211 
<< m2 >>
rect 46 210 47 211 
<< pdiffusion >>
rect 48 210 49 211 
<< pdiffusion >>
rect 49 210 50 211 
<< pdiffusion >>
rect 50 210 51 211 
<< pdiffusion >>
rect 51 210 52 211 
<< pdiffusion >>
rect 52 210 53 211 
<< pdiffusion >>
rect 53 210 54 211 
<< m1 >>
rect 55 210 56 211 
<< m2 >>
rect 55 210 56 211 
<< pdiffusion >>
rect 66 210 67 211 
<< pdiffusion >>
rect 67 210 68 211 
<< pdiffusion >>
rect 68 210 69 211 
<< pdiffusion >>
rect 69 210 70 211 
<< m1 >>
rect 70 210 71 211 
<< pdiffusion >>
rect 70 210 71 211 
<< pdiffusion >>
rect 71 210 72 211 
<< m1 >>
rect 73 210 74 211 
<< m2 >>
rect 74 210 75 211 
<< m1 >>
rect 82 210 83 211 
<< pdiffusion >>
rect 84 210 85 211 
<< pdiffusion >>
rect 85 210 86 211 
<< pdiffusion >>
rect 86 210 87 211 
<< pdiffusion >>
rect 87 210 88 211 
<< m1 >>
rect 88 210 89 211 
<< pdiffusion >>
rect 88 210 89 211 
<< pdiffusion >>
rect 89 210 90 211 
<< m1 >>
rect 93 210 94 211 
<< m1 >>
rect 95 210 96 211 
<< pdiffusion >>
rect 102 210 103 211 
<< pdiffusion >>
rect 103 210 104 211 
<< pdiffusion >>
rect 104 210 105 211 
<< pdiffusion >>
rect 105 210 106 211 
<< m1 >>
rect 106 210 107 211 
<< pdiffusion >>
rect 106 210 107 211 
<< pdiffusion >>
rect 107 210 108 211 
<< m1 >>
rect 113 210 114 211 
<< pdiffusion >>
rect 120 210 121 211 
<< m1 >>
rect 121 210 122 211 
<< pdiffusion >>
rect 121 210 122 211 
<< pdiffusion >>
rect 122 210 123 211 
<< pdiffusion >>
rect 123 210 124 211 
<< m1 >>
rect 124 210 125 211 
<< pdiffusion >>
rect 124 210 125 211 
<< pdiffusion >>
rect 125 210 126 211 
<< pdiffusion >>
rect 138 210 139 211 
<< pdiffusion >>
rect 139 210 140 211 
<< pdiffusion >>
rect 140 210 141 211 
<< pdiffusion >>
rect 141 210 142 211 
<< pdiffusion >>
rect 142 210 143 211 
<< pdiffusion >>
rect 143 210 144 211 
<< m1 >>
rect 150 210 151 211 
<< m1 >>
rect 152 210 153 211 
<< m1 >>
rect 154 210 155 211 
<< pdiffusion >>
rect 156 210 157 211 
<< pdiffusion >>
rect 157 210 158 211 
<< pdiffusion >>
rect 158 210 159 211 
<< pdiffusion >>
rect 159 210 160 211 
<< m1 >>
rect 160 210 161 211 
<< pdiffusion >>
rect 160 210 161 211 
<< pdiffusion >>
rect 161 210 162 211 
<< m1 >>
rect 163 210 164 211 
<< pdiffusion >>
rect 174 210 175 211 
<< m1 >>
rect 175 210 176 211 
<< pdiffusion >>
rect 175 210 176 211 
<< pdiffusion >>
rect 176 210 177 211 
<< pdiffusion >>
rect 177 210 178 211 
<< pdiffusion >>
rect 178 210 179 211 
<< pdiffusion >>
rect 179 210 180 211 
<< m1 >>
rect 188 210 189 211 
<< m1 >>
rect 190 210 191 211 
<< pdiffusion >>
rect 192 210 193 211 
<< pdiffusion >>
rect 193 210 194 211 
<< pdiffusion >>
rect 194 210 195 211 
<< pdiffusion >>
rect 195 210 196 211 
<< pdiffusion >>
rect 196 210 197 211 
<< pdiffusion >>
rect 197 210 198 211 
<< m1 >>
rect 208 210 209 211 
<< pdiffusion >>
rect 210 210 211 211 
<< m1 >>
rect 211 210 212 211 
<< pdiffusion >>
rect 211 210 212 211 
<< pdiffusion >>
rect 212 210 213 211 
<< pdiffusion >>
rect 213 210 214 211 
<< pdiffusion >>
rect 214 210 215 211 
<< pdiffusion >>
rect 215 210 216 211 
<< pdiffusion >>
rect 228 210 229 211 
<< pdiffusion >>
rect 229 210 230 211 
<< pdiffusion >>
rect 230 210 231 211 
<< pdiffusion >>
rect 231 210 232 211 
<< pdiffusion >>
rect 232 210 233 211 
<< pdiffusion >>
rect 233 210 234 211 
<< pdiffusion >>
rect 246 210 247 211 
<< pdiffusion >>
rect 247 210 248 211 
<< pdiffusion >>
rect 248 210 249 211 
<< pdiffusion >>
rect 249 210 250 211 
<< pdiffusion >>
rect 250 210 251 211 
<< pdiffusion >>
rect 251 210 252 211 
<< pdiffusion >>
rect 12 211 13 212 
<< pdiffusion >>
rect 13 211 14 212 
<< pdiffusion >>
rect 14 211 15 212 
<< pdiffusion >>
rect 15 211 16 212 
<< pdiffusion >>
rect 16 211 17 212 
<< pdiffusion >>
rect 17 211 18 212 
<< m1 >>
rect 19 211 20 212 
<< m2 >>
rect 20 211 21 212 
<< m1 >>
rect 28 211 29 212 
<< pdiffusion >>
rect 30 211 31 212 
<< pdiffusion >>
rect 31 211 32 212 
<< pdiffusion >>
rect 32 211 33 212 
<< pdiffusion >>
rect 33 211 34 212 
<< pdiffusion >>
rect 34 211 35 212 
<< pdiffusion >>
rect 35 211 36 212 
<< m1 >>
rect 46 211 47 212 
<< m2 >>
rect 46 211 47 212 
<< pdiffusion >>
rect 48 211 49 212 
<< pdiffusion >>
rect 49 211 50 212 
<< pdiffusion >>
rect 50 211 51 212 
<< pdiffusion >>
rect 51 211 52 212 
<< pdiffusion >>
rect 52 211 53 212 
<< pdiffusion >>
rect 53 211 54 212 
<< m1 >>
rect 55 211 56 212 
<< m2 >>
rect 55 211 56 212 
<< pdiffusion >>
rect 66 211 67 212 
<< pdiffusion >>
rect 67 211 68 212 
<< pdiffusion >>
rect 68 211 69 212 
<< pdiffusion >>
rect 69 211 70 212 
<< pdiffusion >>
rect 70 211 71 212 
<< pdiffusion >>
rect 71 211 72 212 
<< m1 >>
rect 73 211 74 212 
<< m2 >>
rect 74 211 75 212 
<< m1 >>
rect 82 211 83 212 
<< pdiffusion >>
rect 84 211 85 212 
<< pdiffusion >>
rect 85 211 86 212 
<< pdiffusion >>
rect 86 211 87 212 
<< pdiffusion >>
rect 87 211 88 212 
<< pdiffusion >>
rect 88 211 89 212 
<< pdiffusion >>
rect 89 211 90 212 
<< m1 >>
rect 93 211 94 212 
<< m1 >>
rect 95 211 96 212 
<< pdiffusion >>
rect 102 211 103 212 
<< pdiffusion >>
rect 103 211 104 212 
<< pdiffusion >>
rect 104 211 105 212 
<< pdiffusion >>
rect 105 211 106 212 
<< pdiffusion >>
rect 106 211 107 212 
<< pdiffusion >>
rect 107 211 108 212 
<< m1 >>
rect 113 211 114 212 
<< pdiffusion >>
rect 120 211 121 212 
<< pdiffusion >>
rect 121 211 122 212 
<< pdiffusion >>
rect 122 211 123 212 
<< pdiffusion >>
rect 123 211 124 212 
<< pdiffusion >>
rect 124 211 125 212 
<< pdiffusion >>
rect 125 211 126 212 
<< pdiffusion >>
rect 138 211 139 212 
<< pdiffusion >>
rect 139 211 140 212 
<< pdiffusion >>
rect 140 211 141 212 
<< pdiffusion >>
rect 141 211 142 212 
<< pdiffusion >>
rect 142 211 143 212 
<< pdiffusion >>
rect 143 211 144 212 
<< m1 >>
rect 150 211 151 212 
<< m1 >>
rect 152 211 153 212 
<< m1 >>
rect 154 211 155 212 
<< pdiffusion >>
rect 156 211 157 212 
<< pdiffusion >>
rect 157 211 158 212 
<< pdiffusion >>
rect 158 211 159 212 
<< pdiffusion >>
rect 159 211 160 212 
<< pdiffusion >>
rect 160 211 161 212 
<< pdiffusion >>
rect 161 211 162 212 
<< m1 >>
rect 163 211 164 212 
<< pdiffusion >>
rect 174 211 175 212 
<< pdiffusion >>
rect 175 211 176 212 
<< pdiffusion >>
rect 176 211 177 212 
<< pdiffusion >>
rect 177 211 178 212 
<< pdiffusion >>
rect 178 211 179 212 
<< pdiffusion >>
rect 179 211 180 212 
<< m1 >>
rect 188 211 189 212 
<< m1 >>
rect 190 211 191 212 
<< pdiffusion >>
rect 192 211 193 212 
<< pdiffusion >>
rect 193 211 194 212 
<< pdiffusion >>
rect 194 211 195 212 
<< pdiffusion >>
rect 195 211 196 212 
<< pdiffusion >>
rect 196 211 197 212 
<< pdiffusion >>
rect 197 211 198 212 
<< m1 >>
rect 208 211 209 212 
<< pdiffusion >>
rect 210 211 211 212 
<< pdiffusion >>
rect 211 211 212 212 
<< pdiffusion >>
rect 212 211 213 212 
<< pdiffusion >>
rect 213 211 214 212 
<< pdiffusion >>
rect 214 211 215 212 
<< pdiffusion >>
rect 215 211 216 212 
<< pdiffusion >>
rect 228 211 229 212 
<< pdiffusion >>
rect 229 211 230 212 
<< pdiffusion >>
rect 230 211 231 212 
<< pdiffusion >>
rect 231 211 232 212 
<< pdiffusion >>
rect 232 211 233 212 
<< pdiffusion >>
rect 233 211 234 212 
<< pdiffusion >>
rect 246 211 247 212 
<< pdiffusion >>
rect 247 211 248 212 
<< pdiffusion >>
rect 248 211 249 212 
<< pdiffusion >>
rect 249 211 250 212 
<< pdiffusion >>
rect 250 211 251 212 
<< pdiffusion >>
rect 251 211 252 212 
<< pdiffusion >>
rect 12 212 13 213 
<< pdiffusion >>
rect 13 212 14 213 
<< pdiffusion >>
rect 14 212 15 213 
<< pdiffusion >>
rect 15 212 16 213 
<< pdiffusion >>
rect 16 212 17 213 
<< pdiffusion >>
rect 17 212 18 213 
<< m1 >>
rect 19 212 20 213 
<< m2 >>
rect 20 212 21 213 
<< m1 >>
rect 28 212 29 213 
<< pdiffusion >>
rect 30 212 31 213 
<< pdiffusion >>
rect 31 212 32 213 
<< pdiffusion >>
rect 32 212 33 213 
<< pdiffusion >>
rect 33 212 34 213 
<< pdiffusion >>
rect 34 212 35 213 
<< pdiffusion >>
rect 35 212 36 213 
<< m1 >>
rect 46 212 47 213 
<< m2 >>
rect 46 212 47 213 
<< pdiffusion >>
rect 48 212 49 213 
<< pdiffusion >>
rect 49 212 50 213 
<< pdiffusion >>
rect 50 212 51 213 
<< pdiffusion >>
rect 51 212 52 213 
<< pdiffusion >>
rect 52 212 53 213 
<< pdiffusion >>
rect 53 212 54 213 
<< m1 >>
rect 55 212 56 213 
<< m2 >>
rect 55 212 56 213 
<< pdiffusion >>
rect 66 212 67 213 
<< pdiffusion >>
rect 67 212 68 213 
<< pdiffusion >>
rect 68 212 69 213 
<< pdiffusion >>
rect 69 212 70 213 
<< pdiffusion >>
rect 70 212 71 213 
<< pdiffusion >>
rect 71 212 72 213 
<< m1 >>
rect 73 212 74 213 
<< m2 >>
rect 74 212 75 213 
<< m1 >>
rect 82 212 83 213 
<< pdiffusion >>
rect 84 212 85 213 
<< pdiffusion >>
rect 85 212 86 213 
<< pdiffusion >>
rect 86 212 87 213 
<< pdiffusion >>
rect 87 212 88 213 
<< pdiffusion >>
rect 88 212 89 213 
<< pdiffusion >>
rect 89 212 90 213 
<< m1 >>
rect 93 212 94 213 
<< m1 >>
rect 95 212 96 213 
<< pdiffusion >>
rect 102 212 103 213 
<< pdiffusion >>
rect 103 212 104 213 
<< pdiffusion >>
rect 104 212 105 213 
<< pdiffusion >>
rect 105 212 106 213 
<< pdiffusion >>
rect 106 212 107 213 
<< pdiffusion >>
rect 107 212 108 213 
<< m1 >>
rect 113 212 114 213 
<< pdiffusion >>
rect 120 212 121 213 
<< pdiffusion >>
rect 121 212 122 213 
<< pdiffusion >>
rect 122 212 123 213 
<< pdiffusion >>
rect 123 212 124 213 
<< pdiffusion >>
rect 124 212 125 213 
<< pdiffusion >>
rect 125 212 126 213 
<< pdiffusion >>
rect 138 212 139 213 
<< pdiffusion >>
rect 139 212 140 213 
<< pdiffusion >>
rect 140 212 141 213 
<< pdiffusion >>
rect 141 212 142 213 
<< pdiffusion >>
rect 142 212 143 213 
<< pdiffusion >>
rect 143 212 144 213 
<< m1 >>
rect 150 212 151 213 
<< m1 >>
rect 152 212 153 213 
<< m1 >>
rect 154 212 155 213 
<< pdiffusion >>
rect 156 212 157 213 
<< pdiffusion >>
rect 157 212 158 213 
<< pdiffusion >>
rect 158 212 159 213 
<< pdiffusion >>
rect 159 212 160 213 
<< pdiffusion >>
rect 160 212 161 213 
<< pdiffusion >>
rect 161 212 162 213 
<< m1 >>
rect 163 212 164 213 
<< pdiffusion >>
rect 174 212 175 213 
<< pdiffusion >>
rect 175 212 176 213 
<< pdiffusion >>
rect 176 212 177 213 
<< pdiffusion >>
rect 177 212 178 213 
<< pdiffusion >>
rect 178 212 179 213 
<< pdiffusion >>
rect 179 212 180 213 
<< m1 >>
rect 188 212 189 213 
<< m1 >>
rect 190 212 191 213 
<< pdiffusion >>
rect 192 212 193 213 
<< pdiffusion >>
rect 193 212 194 213 
<< pdiffusion >>
rect 194 212 195 213 
<< pdiffusion >>
rect 195 212 196 213 
<< pdiffusion >>
rect 196 212 197 213 
<< pdiffusion >>
rect 197 212 198 213 
<< m1 >>
rect 208 212 209 213 
<< pdiffusion >>
rect 210 212 211 213 
<< pdiffusion >>
rect 211 212 212 213 
<< pdiffusion >>
rect 212 212 213 213 
<< pdiffusion >>
rect 213 212 214 213 
<< pdiffusion >>
rect 214 212 215 213 
<< pdiffusion >>
rect 215 212 216 213 
<< pdiffusion >>
rect 228 212 229 213 
<< pdiffusion >>
rect 229 212 230 213 
<< pdiffusion >>
rect 230 212 231 213 
<< pdiffusion >>
rect 231 212 232 213 
<< pdiffusion >>
rect 232 212 233 213 
<< pdiffusion >>
rect 233 212 234 213 
<< pdiffusion >>
rect 246 212 247 213 
<< pdiffusion >>
rect 247 212 248 213 
<< pdiffusion >>
rect 248 212 249 213 
<< pdiffusion >>
rect 249 212 250 213 
<< pdiffusion >>
rect 250 212 251 213 
<< pdiffusion >>
rect 251 212 252 213 
<< pdiffusion >>
rect 12 213 13 214 
<< pdiffusion >>
rect 13 213 14 214 
<< pdiffusion >>
rect 14 213 15 214 
<< pdiffusion >>
rect 15 213 16 214 
<< pdiffusion >>
rect 16 213 17 214 
<< pdiffusion >>
rect 17 213 18 214 
<< m1 >>
rect 19 213 20 214 
<< m2 >>
rect 20 213 21 214 
<< m1 >>
rect 28 213 29 214 
<< pdiffusion >>
rect 30 213 31 214 
<< pdiffusion >>
rect 31 213 32 214 
<< pdiffusion >>
rect 32 213 33 214 
<< pdiffusion >>
rect 33 213 34 214 
<< pdiffusion >>
rect 34 213 35 214 
<< pdiffusion >>
rect 35 213 36 214 
<< m1 >>
rect 46 213 47 214 
<< m2 >>
rect 46 213 47 214 
<< pdiffusion >>
rect 48 213 49 214 
<< pdiffusion >>
rect 49 213 50 214 
<< pdiffusion >>
rect 50 213 51 214 
<< pdiffusion >>
rect 51 213 52 214 
<< pdiffusion >>
rect 52 213 53 214 
<< pdiffusion >>
rect 53 213 54 214 
<< m1 >>
rect 55 213 56 214 
<< m2 >>
rect 55 213 56 214 
<< pdiffusion >>
rect 66 213 67 214 
<< pdiffusion >>
rect 67 213 68 214 
<< pdiffusion >>
rect 68 213 69 214 
<< pdiffusion >>
rect 69 213 70 214 
<< pdiffusion >>
rect 70 213 71 214 
<< pdiffusion >>
rect 71 213 72 214 
<< m1 >>
rect 73 213 74 214 
<< m2 >>
rect 74 213 75 214 
<< m1 >>
rect 82 213 83 214 
<< pdiffusion >>
rect 84 213 85 214 
<< pdiffusion >>
rect 85 213 86 214 
<< pdiffusion >>
rect 86 213 87 214 
<< pdiffusion >>
rect 87 213 88 214 
<< pdiffusion >>
rect 88 213 89 214 
<< pdiffusion >>
rect 89 213 90 214 
<< m1 >>
rect 93 213 94 214 
<< m1 >>
rect 95 213 96 214 
<< pdiffusion >>
rect 102 213 103 214 
<< pdiffusion >>
rect 103 213 104 214 
<< pdiffusion >>
rect 104 213 105 214 
<< pdiffusion >>
rect 105 213 106 214 
<< pdiffusion >>
rect 106 213 107 214 
<< pdiffusion >>
rect 107 213 108 214 
<< m1 >>
rect 113 213 114 214 
<< pdiffusion >>
rect 120 213 121 214 
<< pdiffusion >>
rect 121 213 122 214 
<< pdiffusion >>
rect 122 213 123 214 
<< pdiffusion >>
rect 123 213 124 214 
<< pdiffusion >>
rect 124 213 125 214 
<< pdiffusion >>
rect 125 213 126 214 
<< pdiffusion >>
rect 138 213 139 214 
<< pdiffusion >>
rect 139 213 140 214 
<< pdiffusion >>
rect 140 213 141 214 
<< pdiffusion >>
rect 141 213 142 214 
<< pdiffusion >>
rect 142 213 143 214 
<< pdiffusion >>
rect 143 213 144 214 
<< m1 >>
rect 150 213 151 214 
<< m1 >>
rect 152 213 153 214 
<< m1 >>
rect 154 213 155 214 
<< pdiffusion >>
rect 156 213 157 214 
<< pdiffusion >>
rect 157 213 158 214 
<< pdiffusion >>
rect 158 213 159 214 
<< pdiffusion >>
rect 159 213 160 214 
<< pdiffusion >>
rect 160 213 161 214 
<< pdiffusion >>
rect 161 213 162 214 
<< m1 >>
rect 163 213 164 214 
<< pdiffusion >>
rect 174 213 175 214 
<< pdiffusion >>
rect 175 213 176 214 
<< pdiffusion >>
rect 176 213 177 214 
<< pdiffusion >>
rect 177 213 178 214 
<< pdiffusion >>
rect 178 213 179 214 
<< pdiffusion >>
rect 179 213 180 214 
<< m1 >>
rect 188 213 189 214 
<< m1 >>
rect 190 213 191 214 
<< pdiffusion >>
rect 192 213 193 214 
<< pdiffusion >>
rect 193 213 194 214 
<< pdiffusion >>
rect 194 213 195 214 
<< pdiffusion >>
rect 195 213 196 214 
<< pdiffusion >>
rect 196 213 197 214 
<< pdiffusion >>
rect 197 213 198 214 
<< m1 >>
rect 208 213 209 214 
<< pdiffusion >>
rect 210 213 211 214 
<< pdiffusion >>
rect 211 213 212 214 
<< pdiffusion >>
rect 212 213 213 214 
<< pdiffusion >>
rect 213 213 214 214 
<< pdiffusion >>
rect 214 213 215 214 
<< pdiffusion >>
rect 215 213 216 214 
<< pdiffusion >>
rect 228 213 229 214 
<< pdiffusion >>
rect 229 213 230 214 
<< pdiffusion >>
rect 230 213 231 214 
<< pdiffusion >>
rect 231 213 232 214 
<< pdiffusion >>
rect 232 213 233 214 
<< pdiffusion >>
rect 233 213 234 214 
<< pdiffusion >>
rect 246 213 247 214 
<< pdiffusion >>
rect 247 213 248 214 
<< pdiffusion >>
rect 248 213 249 214 
<< pdiffusion >>
rect 249 213 250 214 
<< pdiffusion >>
rect 250 213 251 214 
<< pdiffusion >>
rect 251 213 252 214 
<< pdiffusion >>
rect 12 214 13 215 
<< pdiffusion >>
rect 13 214 14 215 
<< pdiffusion >>
rect 14 214 15 215 
<< pdiffusion >>
rect 15 214 16 215 
<< pdiffusion >>
rect 16 214 17 215 
<< pdiffusion >>
rect 17 214 18 215 
<< m1 >>
rect 19 214 20 215 
<< m2 >>
rect 20 214 21 215 
<< m1 >>
rect 28 214 29 215 
<< pdiffusion >>
rect 30 214 31 215 
<< pdiffusion >>
rect 31 214 32 215 
<< pdiffusion >>
rect 32 214 33 215 
<< pdiffusion >>
rect 33 214 34 215 
<< pdiffusion >>
rect 34 214 35 215 
<< pdiffusion >>
rect 35 214 36 215 
<< m1 >>
rect 46 214 47 215 
<< m2 >>
rect 46 214 47 215 
<< pdiffusion >>
rect 48 214 49 215 
<< pdiffusion >>
rect 49 214 50 215 
<< pdiffusion >>
rect 50 214 51 215 
<< pdiffusion >>
rect 51 214 52 215 
<< pdiffusion >>
rect 52 214 53 215 
<< pdiffusion >>
rect 53 214 54 215 
<< m1 >>
rect 55 214 56 215 
<< m2 >>
rect 55 214 56 215 
<< pdiffusion >>
rect 66 214 67 215 
<< pdiffusion >>
rect 67 214 68 215 
<< pdiffusion >>
rect 68 214 69 215 
<< pdiffusion >>
rect 69 214 70 215 
<< pdiffusion >>
rect 70 214 71 215 
<< pdiffusion >>
rect 71 214 72 215 
<< m1 >>
rect 73 214 74 215 
<< m2 >>
rect 74 214 75 215 
<< m1 >>
rect 82 214 83 215 
<< pdiffusion >>
rect 84 214 85 215 
<< pdiffusion >>
rect 85 214 86 215 
<< pdiffusion >>
rect 86 214 87 215 
<< pdiffusion >>
rect 87 214 88 215 
<< pdiffusion >>
rect 88 214 89 215 
<< pdiffusion >>
rect 89 214 90 215 
<< m1 >>
rect 93 214 94 215 
<< m1 >>
rect 95 214 96 215 
<< pdiffusion >>
rect 102 214 103 215 
<< pdiffusion >>
rect 103 214 104 215 
<< pdiffusion >>
rect 104 214 105 215 
<< pdiffusion >>
rect 105 214 106 215 
<< pdiffusion >>
rect 106 214 107 215 
<< pdiffusion >>
rect 107 214 108 215 
<< m1 >>
rect 113 214 114 215 
<< pdiffusion >>
rect 120 214 121 215 
<< pdiffusion >>
rect 121 214 122 215 
<< pdiffusion >>
rect 122 214 123 215 
<< pdiffusion >>
rect 123 214 124 215 
<< pdiffusion >>
rect 124 214 125 215 
<< pdiffusion >>
rect 125 214 126 215 
<< pdiffusion >>
rect 138 214 139 215 
<< pdiffusion >>
rect 139 214 140 215 
<< pdiffusion >>
rect 140 214 141 215 
<< pdiffusion >>
rect 141 214 142 215 
<< pdiffusion >>
rect 142 214 143 215 
<< pdiffusion >>
rect 143 214 144 215 
<< m1 >>
rect 150 214 151 215 
<< m1 >>
rect 152 214 153 215 
<< m1 >>
rect 154 214 155 215 
<< pdiffusion >>
rect 156 214 157 215 
<< pdiffusion >>
rect 157 214 158 215 
<< pdiffusion >>
rect 158 214 159 215 
<< pdiffusion >>
rect 159 214 160 215 
<< pdiffusion >>
rect 160 214 161 215 
<< pdiffusion >>
rect 161 214 162 215 
<< m1 >>
rect 163 214 164 215 
<< pdiffusion >>
rect 174 214 175 215 
<< pdiffusion >>
rect 175 214 176 215 
<< pdiffusion >>
rect 176 214 177 215 
<< pdiffusion >>
rect 177 214 178 215 
<< pdiffusion >>
rect 178 214 179 215 
<< pdiffusion >>
rect 179 214 180 215 
<< m1 >>
rect 188 214 189 215 
<< m1 >>
rect 190 214 191 215 
<< pdiffusion >>
rect 192 214 193 215 
<< pdiffusion >>
rect 193 214 194 215 
<< pdiffusion >>
rect 194 214 195 215 
<< pdiffusion >>
rect 195 214 196 215 
<< pdiffusion >>
rect 196 214 197 215 
<< pdiffusion >>
rect 197 214 198 215 
<< m1 >>
rect 208 214 209 215 
<< pdiffusion >>
rect 210 214 211 215 
<< pdiffusion >>
rect 211 214 212 215 
<< pdiffusion >>
rect 212 214 213 215 
<< pdiffusion >>
rect 213 214 214 215 
<< pdiffusion >>
rect 214 214 215 215 
<< pdiffusion >>
rect 215 214 216 215 
<< pdiffusion >>
rect 228 214 229 215 
<< pdiffusion >>
rect 229 214 230 215 
<< pdiffusion >>
rect 230 214 231 215 
<< pdiffusion >>
rect 231 214 232 215 
<< pdiffusion >>
rect 232 214 233 215 
<< pdiffusion >>
rect 233 214 234 215 
<< pdiffusion >>
rect 246 214 247 215 
<< pdiffusion >>
rect 247 214 248 215 
<< pdiffusion >>
rect 248 214 249 215 
<< pdiffusion >>
rect 249 214 250 215 
<< pdiffusion >>
rect 250 214 251 215 
<< pdiffusion >>
rect 251 214 252 215 
<< pdiffusion >>
rect 12 215 13 216 
<< pdiffusion >>
rect 13 215 14 216 
<< pdiffusion >>
rect 14 215 15 216 
<< pdiffusion >>
rect 15 215 16 216 
<< m1 >>
rect 16 215 17 216 
<< pdiffusion >>
rect 16 215 17 216 
<< pdiffusion >>
rect 17 215 18 216 
<< m1 >>
rect 19 215 20 216 
<< m2 >>
rect 20 215 21 216 
<< m1 >>
rect 28 215 29 216 
<< pdiffusion >>
rect 30 215 31 216 
<< pdiffusion >>
rect 31 215 32 216 
<< pdiffusion >>
rect 32 215 33 216 
<< pdiffusion >>
rect 33 215 34 216 
<< pdiffusion >>
rect 34 215 35 216 
<< pdiffusion >>
rect 35 215 36 216 
<< m1 >>
rect 46 215 47 216 
<< m2 >>
rect 46 215 47 216 
<< pdiffusion >>
rect 48 215 49 216 
<< pdiffusion >>
rect 49 215 50 216 
<< pdiffusion >>
rect 50 215 51 216 
<< pdiffusion >>
rect 51 215 52 216 
<< pdiffusion >>
rect 52 215 53 216 
<< pdiffusion >>
rect 53 215 54 216 
<< m1 >>
rect 55 215 56 216 
<< m2 >>
rect 55 215 56 216 
<< pdiffusion >>
rect 66 215 67 216 
<< pdiffusion >>
rect 67 215 68 216 
<< pdiffusion >>
rect 68 215 69 216 
<< pdiffusion >>
rect 69 215 70 216 
<< m1 >>
rect 70 215 71 216 
<< pdiffusion >>
rect 70 215 71 216 
<< pdiffusion >>
rect 71 215 72 216 
<< m1 >>
rect 73 215 74 216 
<< m2 >>
rect 74 215 75 216 
<< m1 >>
rect 82 215 83 216 
<< pdiffusion >>
rect 84 215 85 216 
<< pdiffusion >>
rect 85 215 86 216 
<< pdiffusion >>
rect 86 215 87 216 
<< pdiffusion >>
rect 87 215 88 216 
<< m1 >>
rect 88 215 89 216 
<< pdiffusion >>
rect 88 215 89 216 
<< pdiffusion >>
rect 89 215 90 216 
<< m1 >>
rect 93 215 94 216 
<< m1 >>
rect 95 215 96 216 
<< pdiffusion >>
rect 102 215 103 216 
<< m1 >>
rect 103 215 104 216 
<< pdiffusion >>
rect 103 215 104 216 
<< pdiffusion >>
rect 104 215 105 216 
<< pdiffusion >>
rect 105 215 106 216 
<< pdiffusion >>
rect 106 215 107 216 
<< pdiffusion >>
rect 107 215 108 216 
<< m1 >>
rect 113 215 114 216 
<< pdiffusion >>
rect 120 215 121 216 
<< pdiffusion >>
rect 121 215 122 216 
<< pdiffusion >>
rect 122 215 123 216 
<< pdiffusion >>
rect 123 215 124 216 
<< m1 >>
rect 124 215 125 216 
<< pdiffusion >>
rect 124 215 125 216 
<< pdiffusion >>
rect 125 215 126 216 
<< pdiffusion >>
rect 138 215 139 216 
<< m1 >>
rect 139 215 140 216 
<< pdiffusion >>
rect 139 215 140 216 
<< pdiffusion >>
rect 140 215 141 216 
<< pdiffusion >>
rect 141 215 142 216 
<< pdiffusion >>
rect 142 215 143 216 
<< pdiffusion >>
rect 143 215 144 216 
<< m1 >>
rect 150 215 151 216 
<< m1 >>
rect 152 215 153 216 
<< m1 >>
rect 154 215 155 216 
<< pdiffusion >>
rect 156 215 157 216 
<< pdiffusion >>
rect 157 215 158 216 
<< pdiffusion >>
rect 158 215 159 216 
<< pdiffusion >>
rect 159 215 160 216 
<< pdiffusion >>
rect 160 215 161 216 
<< pdiffusion >>
rect 161 215 162 216 
<< m1 >>
rect 163 215 164 216 
<< pdiffusion >>
rect 174 215 175 216 
<< pdiffusion >>
rect 175 215 176 216 
<< pdiffusion >>
rect 176 215 177 216 
<< pdiffusion >>
rect 177 215 178 216 
<< pdiffusion >>
rect 178 215 179 216 
<< pdiffusion >>
rect 179 215 180 216 
<< m1 >>
rect 188 215 189 216 
<< m1 >>
rect 190 215 191 216 
<< pdiffusion >>
rect 192 215 193 216 
<< pdiffusion >>
rect 193 215 194 216 
<< pdiffusion >>
rect 194 215 195 216 
<< pdiffusion >>
rect 195 215 196 216 
<< pdiffusion >>
rect 196 215 197 216 
<< pdiffusion >>
rect 197 215 198 216 
<< m1 >>
rect 208 215 209 216 
<< pdiffusion >>
rect 210 215 211 216 
<< pdiffusion >>
rect 211 215 212 216 
<< pdiffusion >>
rect 212 215 213 216 
<< pdiffusion >>
rect 213 215 214 216 
<< pdiffusion >>
rect 214 215 215 216 
<< pdiffusion >>
rect 215 215 216 216 
<< pdiffusion >>
rect 228 215 229 216 
<< pdiffusion >>
rect 229 215 230 216 
<< pdiffusion >>
rect 230 215 231 216 
<< pdiffusion >>
rect 231 215 232 216 
<< pdiffusion >>
rect 232 215 233 216 
<< pdiffusion >>
rect 233 215 234 216 
<< pdiffusion >>
rect 246 215 247 216 
<< pdiffusion >>
rect 247 215 248 216 
<< pdiffusion >>
rect 248 215 249 216 
<< pdiffusion >>
rect 249 215 250 216 
<< pdiffusion >>
rect 250 215 251 216 
<< pdiffusion >>
rect 251 215 252 216 
<< m1 >>
rect 16 216 17 217 
<< m1 >>
rect 19 216 20 217 
<< m2 >>
rect 20 216 21 217 
<< m1 >>
rect 28 216 29 217 
<< m1 >>
rect 46 216 47 217 
<< m2 >>
rect 46 216 47 217 
<< m1 >>
rect 55 216 56 217 
<< m2 >>
rect 55 216 56 217 
<< m1 >>
rect 70 216 71 217 
<< m1 >>
rect 73 216 74 217 
<< m2 >>
rect 74 216 75 217 
<< m1 >>
rect 82 216 83 217 
<< m1 >>
rect 88 216 89 217 
<< m1 >>
rect 93 216 94 217 
<< m1 >>
rect 95 216 96 217 
<< m1 >>
rect 103 216 104 217 
<< m1 >>
rect 113 216 114 217 
<< m1 >>
rect 124 216 125 217 
<< m1 >>
rect 139 216 140 217 
<< m1 >>
rect 150 216 151 217 
<< m2 >>
rect 150 216 151 217 
<< m2c >>
rect 150 216 151 217 
<< m1 >>
rect 150 216 151 217 
<< m2 >>
rect 150 216 151 217 
<< m1 >>
rect 152 216 153 217 
<< m2 >>
rect 152 216 153 217 
<< m2c >>
rect 152 216 153 217 
<< m1 >>
rect 152 216 153 217 
<< m2 >>
rect 152 216 153 217 
<< m1 >>
rect 154 216 155 217 
<< m1 >>
rect 163 216 164 217 
<< m1 >>
rect 188 216 189 217 
<< m1 >>
rect 190 216 191 217 
<< m1 >>
rect 208 216 209 217 
<< m1 >>
rect 16 217 17 218 
<< m1 >>
rect 19 217 20 218 
<< m2 >>
rect 20 217 21 218 
<< m1 >>
rect 28 217 29 218 
<< m1 >>
rect 46 217 47 218 
<< m2 >>
rect 46 217 47 218 
<< m1 >>
rect 53 217 54 218 
<< m2 >>
rect 53 217 54 218 
<< m2c >>
rect 53 217 54 218 
<< m1 >>
rect 53 217 54 218 
<< m2 >>
rect 53 217 54 218 
<< m2 >>
rect 54 217 55 218 
<< m1 >>
rect 55 217 56 218 
<< m2 >>
rect 55 217 56 218 
<< m1 >>
rect 70 217 71 218 
<< m1 >>
rect 73 217 74 218 
<< m2 >>
rect 74 217 75 218 
<< m1 >>
rect 82 217 83 218 
<< m1 >>
rect 88 217 89 218 
<< m1 >>
rect 93 217 94 218 
<< m1 >>
rect 95 217 96 218 
<< m1 >>
rect 103 217 104 218 
<< m1 >>
rect 113 217 114 218 
<< m1 >>
rect 124 217 125 218 
<< m1 >>
rect 139 217 140 218 
<< m2 >>
rect 150 217 151 218 
<< m2 >>
rect 152 217 153 218 
<< m1 >>
rect 154 217 155 218 
<< m1 >>
rect 163 217 164 218 
<< m1 >>
rect 188 217 189 218 
<< m1 >>
rect 190 217 191 218 
<< m1 >>
rect 208 217 209 218 
<< m1 >>
rect 16 218 17 219 
<< m1 >>
rect 19 218 20 219 
<< m2 >>
rect 20 218 21 219 
<< m1 >>
rect 28 218 29 219 
<< m1 >>
rect 46 218 47 219 
<< m2 >>
rect 46 218 47 219 
<< m1 >>
rect 52 218 53 219 
<< m1 >>
rect 53 218 54 219 
<< m1 >>
rect 55 218 56 219 
<< m1 >>
rect 70 218 71 219 
<< m1 >>
rect 73 218 74 219 
<< m2 >>
rect 74 218 75 219 
<< m1 >>
rect 82 218 83 219 
<< m1 >>
rect 88 218 89 219 
<< m1 >>
rect 89 218 90 219 
<< m2 >>
rect 89 218 90 219 
<< m2c >>
rect 89 218 90 219 
<< m1 >>
rect 89 218 90 219 
<< m2 >>
rect 89 218 90 219 
<< m1 >>
rect 91 218 92 219 
<< m2 >>
rect 91 218 92 219 
<< m2c >>
rect 91 218 92 219 
<< m1 >>
rect 91 218 92 219 
<< m2 >>
rect 91 218 92 219 
<< m1 >>
rect 92 218 93 219 
<< m1 >>
rect 93 218 94 219 
<< m1 >>
rect 95 218 96 219 
<< m2 >>
rect 95 218 96 219 
<< m2c >>
rect 95 218 96 219 
<< m1 >>
rect 95 218 96 219 
<< m2 >>
rect 95 218 96 219 
<< m1 >>
rect 103 218 104 219 
<< m1 >>
rect 104 218 105 219 
<< m1 >>
rect 105 218 106 219 
<< m1 >>
rect 106 218 107 219 
<< m1 >>
rect 107 218 108 219 
<< m1 >>
rect 108 218 109 219 
<< m1 >>
rect 109 218 110 219 
<< m1 >>
rect 110 218 111 219 
<< m1 >>
rect 111 218 112 219 
<< m2 >>
rect 111 218 112 219 
<< m2c >>
rect 111 218 112 219 
<< m1 >>
rect 111 218 112 219 
<< m2 >>
rect 111 218 112 219 
<< m1 >>
rect 113 218 114 219 
<< m2 >>
rect 113 218 114 219 
<< m2c >>
rect 113 218 114 219 
<< m1 >>
rect 113 218 114 219 
<< m2 >>
rect 113 218 114 219 
<< m1 >>
rect 124 218 125 219 
<< m1 >>
rect 125 218 126 219 
<< m1 >>
rect 126 218 127 219 
<< m1 >>
rect 127 218 128 219 
<< m1 >>
rect 128 218 129 219 
<< m1 >>
rect 129 218 130 219 
<< m1 >>
rect 130 218 131 219 
<< m1 >>
rect 131 218 132 219 
<< m1 >>
rect 132 218 133 219 
<< m1 >>
rect 133 218 134 219 
<< m1 >>
rect 134 218 135 219 
<< m1 >>
rect 135 218 136 219 
<< m1 >>
rect 136 218 137 219 
<< m1 >>
rect 137 218 138 219 
<< m2 >>
rect 137 218 138 219 
<< m2c >>
rect 137 218 138 219 
<< m1 >>
rect 137 218 138 219 
<< m2 >>
rect 137 218 138 219 
<< m2 >>
rect 138 218 139 219 
<< m1 >>
rect 139 218 140 219 
<< m1 >>
rect 140 218 141 219 
<< m1 >>
rect 141 218 142 219 
<< m1 >>
rect 142 218 143 219 
<< m1 >>
rect 143 218 144 219 
<< m1 >>
rect 144 218 145 219 
<< m1 >>
rect 145 218 146 219 
<< m1 >>
rect 146 218 147 219 
<< m1 >>
rect 147 218 148 219 
<< m1 >>
rect 148 218 149 219 
<< m1 >>
rect 149 218 150 219 
<< m1 >>
rect 150 218 151 219 
<< m2 >>
rect 150 218 151 219 
<< m1 >>
rect 151 218 152 219 
<< m1 >>
rect 152 218 153 219 
<< m2 >>
rect 152 218 153 219 
<< m1 >>
rect 153 218 154 219 
<< m1 >>
rect 154 218 155 219 
<< m1 >>
rect 158 218 159 219 
<< m2 >>
rect 158 218 159 219 
<< m2c >>
rect 158 218 159 219 
<< m1 >>
rect 158 218 159 219 
<< m2 >>
rect 158 218 159 219 
<< m1 >>
rect 159 218 160 219 
<< m1 >>
rect 160 218 161 219 
<< m1 >>
rect 161 218 162 219 
<< m1 >>
rect 162 218 163 219 
<< m1 >>
rect 163 218 164 219 
<< m1 >>
rect 188 218 189 219 
<< m1 >>
rect 190 218 191 219 
<< m1 >>
rect 208 218 209 219 
<< m1 >>
rect 16 219 17 220 
<< m1 >>
rect 19 219 20 220 
<< m2 >>
rect 20 219 21 220 
<< m1 >>
rect 28 219 29 220 
<< m1 >>
rect 46 219 47 220 
<< m2 >>
rect 46 219 47 220 
<< m1 >>
rect 52 219 53 220 
<< m1 >>
rect 55 219 56 220 
<< m1 >>
rect 70 219 71 220 
<< m1 >>
rect 73 219 74 220 
<< m2 >>
rect 74 219 75 220 
<< m1 >>
rect 82 219 83 220 
<< m2 >>
rect 89 219 90 220 
<< m2 >>
rect 91 219 92 220 
<< m2 >>
rect 95 219 96 220 
<< m2 >>
rect 111 219 112 220 
<< m2 >>
rect 113 219 114 220 
<< m2 >>
rect 138 219 139 220 
<< m2 >>
rect 150 219 151 220 
<< m2 >>
rect 152 219 153 220 
<< m2 >>
rect 158 219 159 220 
<< m1 >>
rect 188 219 189 220 
<< m1 >>
rect 190 219 191 220 
<< m1 >>
rect 208 219 209 220 
<< m1 >>
rect 16 220 17 221 
<< m1 >>
rect 19 220 20 221 
<< m2 >>
rect 20 220 21 221 
<< m1 >>
rect 28 220 29 221 
<< m1 >>
rect 46 220 47 221 
<< m2 >>
rect 46 220 47 221 
<< m1 >>
rect 52 220 53 221 
<< m1 >>
rect 55 220 56 221 
<< m1 >>
rect 56 220 57 221 
<< m1 >>
rect 57 220 58 221 
<< m1 >>
rect 58 220 59 221 
<< m1 >>
rect 59 220 60 221 
<< m1 >>
rect 60 220 61 221 
<< m1 >>
rect 61 220 62 221 
<< m1 >>
rect 62 220 63 221 
<< m1 >>
rect 63 220 64 221 
<< m1 >>
rect 64 220 65 221 
<< m1 >>
rect 65 220 66 221 
<< m1 >>
rect 66 220 67 221 
<< m1 >>
rect 67 220 68 221 
<< m1 >>
rect 68 220 69 221 
<< m1 >>
rect 69 220 70 221 
<< m1 >>
rect 70 220 71 221 
<< m1 >>
rect 73 220 74 221 
<< m2 >>
rect 74 220 75 221 
<< m1 >>
rect 82 220 83 221 
<< m1 >>
rect 83 220 84 221 
<< m1 >>
rect 84 220 85 221 
<< m1 >>
rect 85 220 86 221 
<< m1 >>
rect 86 220 87 221 
<< m1 >>
rect 87 220 88 221 
<< m1 >>
rect 88 220 89 221 
<< m1 >>
rect 89 220 90 221 
<< m2 >>
rect 89 220 90 221 
<< m1 >>
rect 90 220 91 221 
<< m1 >>
rect 91 220 92 221 
<< m2 >>
rect 91 220 92 221 
<< m1 >>
rect 92 220 93 221 
<< m1 >>
rect 93 220 94 221 
<< m1 >>
rect 94 220 95 221 
<< m1 >>
rect 95 220 96 221 
<< m2 >>
rect 95 220 96 221 
<< m1 >>
rect 96 220 97 221 
<< m1 >>
rect 97 220 98 221 
<< m1 >>
rect 98 220 99 221 
<< m1 >>
rect 99 220 100 221 
<< m1 >>
rect 100 220 101 221 
<< m1 >>
rect 101 220 102 221 
<< m1 >>
rect 102 220 103 221 
<< m1 >>
rect 103 220 104 221 
<< m1 >>
rect 104 220 105 221 
<< m1 >>
rect 105 220 106 221 
<< m1 >>
rect 106 220 107 221 
<< m1 >>
rect 107 220 108 221 
<< m1 >>
rect 108 220 109 221 
<< m1 >>
rect 109 220 110 221 
<< m1 >>
rect 110 220 111 221 
<< m1 >>
rect 111 220 112 221 
<< m2 >>
rect 111 220 112 221 
<< m1 >>
rect 112 220 113 221 
<< m1 >>
rect 113 220 114 221 
<< m2 >>
rect 113 220 114 221 
<< m1 >>
rect 114 220 115 221 
<< m1 >>
rect 115 220 116 221 
<< m1 >>
rect 116 220 117 221 
<< m1 >>
rect 117 220 118 221 
<< m1 >>
rect 118 220 119 221 
<< m1 >>
rect 119 220 120 221 
<< m1 >>
rect 120 220 121 221 
<< m1 >>
rect 121 220 122 221 
<< m1 >>
rect 122 220 123 221 
<< m1 >>
rect 123 220 124 221 
<< m1 >>
rect 124 220 125 221 
<< m1 >>
rect 125 220 126 221 
<< m1 >>
rect 126 220 127 221 
<< m1 >>
rect 127 220 128 221 
<< m1 >>
rect 128 220 129 221 
<< m1 >>
rect 129 220 130 221 
<< m1 >>
rect 130 220 131 221 
<< m1 >>
rect 131 220 132 221 
<< m1 >>
rect 132 220 133 221 
<< m1 >>
rect 133 220 134 221 
<< m1 >>
rect 134 220 135 221 
<< m1 >>
rect 135 220 136 221 
<< m1 >>
rect 136 220 137 221 
<< m1 >>
rect 137 220 138 221 
<< m1 >>
rect 138 220 139 221 
<< m2 >>
rect 138 220 139 221 
<< m1 >>
rect 139 220 140 221 
<< m2 >>
rect 139 220 140 221 
<< m2 >>
rect 140 220 141 221 
<< m1 >>
rect 141 220 142 221 
<< m2 >>
rect 141 220 142 221 
<< m2c >>
rect 141 220 142 221 
<< m1 >>
rect 141 220 142 221 
<< m2 >>
rect 141 220 142 221 
<< m1 >>
rect 142 220 143 221 
<< m1 >>
rect 143 220 144 221 
<< m1 >>
rect 144 220 145 221 
<< m1 >>
rect 145 220 146 221 
<< m1 >>
rect 146 220 147 221 
<< m1 >>
rect 147 220 148 221 
<< m1 >>
rect 148 220 149 221 
<< m1 >>
rect 149 220 150 221 
<< m1 >>
rect 150 220 151 221 
<< m2 >>
rect 150 220 151 221 
<< m1 >>
rect 151 220 152 221 
<< m1 >>
rect 152 220 153 221 
<< m2 >>
rect 152 220 153 221 
<< m1 >>
rect 153 220 154 221 
<< m2 >>
rect 153 220 154 221 
<< m1 >>
rect 154 220 155 221 
<< m2 >>
rect 154 220 155 221 
<< m1 >>
rect 155 220 156 221 
<< m2 >>
rect 155 220 156 221 
<< m1 >>
rect 156 220 157 221 
<< m2 >>
rect 156 220 157 221 
<< m1 >>
rect 157 220 158 221 
<< m2 >>
rect 157 220 158 221 
<< m1 >>
rect 158 220 159 221 
<< m2 >>
rect 158 220 159 221 
<< m1 >>
rect 159 220 160 221 
<< m1 >>
rect 160 220 161 221 
<< m1 >>
rect 161 220 162 221 
<< m1 >>
rect 162 220 163 221 
<< m1 >>
rect 163 220 164 221 
<< m1 >>
rect 164 220 165 221 
<< m1 >>
rect 165 220 166 221 
<< m1 >>
rect 166 220 167 221 
<< m1 >>
rect 167 220 168 221 
<< m1 >>
rect 168 220 169 221 
<< m1 >>
rect 169 220 170 221 
<< m1 >>
rect 170 220 171 221 
<< m1 >>
rect 171 220 172 221 
<< m1 >>
rect 172 220 173 221 
<< m1 >>
rect 173 220 174 221 
<< m1 >>
rect 174 220 175 221 
<< m1 >>
rect 175 220 176 221 
<< m1 >>
rect 176 220 177 221 
<< m1 >>
rect 177 220 178 221 
<< m1 >>
rect 178 220 179 221 
<< m1 >>
rect 179 220 180 221 
<< m1 >>
rect 180 220 181 221 
<< m1 >>
rect 181 220 182 221 
<< m1 >>
rect 182 220 183 221 
<< m1 >>
rect 183 220 184 221 
<< m1 >>
rect 184 220 185 221 
<< m1 >>
rect 185 220 186 221 
<< m1 >>
rect 186 220 187 221 
<< m1 >>
rect 187 220 188 221 
<< m1 >>
rect 188 220 189 221 
<< m1 >>
rect 190 220 191 221 
<< m2 >>
rect 191 220 192 221 
<< m1 >>
rect 192 220 193 221 
<< m2 >>
rect 192 220 193 221 
<< m2c >>
rect 192 220 193 221 
<< m1 >>
rect 192 220 193 221 
<< m2 >>
rect 192 220 193 221 
<< m1 >>
rect 193 220 194 221 
<< m1 >>
rect 194 220 195 221 
<< m1 >>
rect 195 220 196 221 
<< m1 >>
rect 196 220 197 221 
<< m1 >>
rect 197 220 198 221 
<< m1 >>
rect 198 220 199 221 
<< m1 >>
rect 199 220 200 221 
<< m1 >>
rect 200 220 201 221 
<< m1 >>
rect 201 220 202 221 
<< m1 >>
rect 202 220 203 221 
<< m1 >>
rect 203 220 204 221 
<< m1 >>
rect 204 220 205 221 
<< m1 >>
rect 205 220 206 221 
<< m1 >>
rect 206 220 207 221 
<< m1 >>
rect 207 220 208 221 
<< m1 >>
rect 208 220 209 221 
<< m1 >>
rect 16 221 17 222 
<< m1 >>
rect 19 221 20 222 
<< m2 >>
rect 20 221 21 222 
<< m1 >>
rect 21 221 22 222 
<< m2 >>
rect 21 221 22 222 
<< m2c >>
rect 21 221 22 222 
<< m1 >>
rect 21 221 22 222 
<< m2 >>
rect 21 221 22 222 
<< m1 >>
rect 22 221 23 222 
<< m1 >>
rect 23 221 24 222 
<< m1 >>
rect 24 221 25 222 
<< m1 >>
rect 28 221 29 222 
<< m1 >>
rect 46 221 47 222 
<< m2 >>
rect 46 221 47 222 
<< m1 >>
rect 52 221 53 222 
<< m1 >>
rect 73 221 74 222 
<< m2 >>
rect 74 221 75 222 
<< m2 >>
rect 89 221 90 222 
<< m2 >>
rect 91 221 92 222 
<< m2 >>
rect 95 221 96 222 
<< m2 >>
rect 111 221 112 222 
<< m2 >>
rect 113 221 114 222 
<< m1 >>
rect 139 221 140 222 
<< m2 >>
rect 150 221 151 222 
<< m1 >>
rect 190 221 191 222 
<< m2 >>
rect 191 221 192 222 
<< m1 >>
rect 16 222 17 223 
<< m1 >>
rect 19 222 20 223 
<< m1 >>
rect 24 222 25 223 
<< m1 >>
rect 28 222 29 223 
<< m1 >>
rect 46 222 47 223 
<< m2 >>
rect 46 222 47 223 
<< m1 >>
rect 52 222 53 223 
<< m1 >>
rect 71 222 72 223 
<< m2 >>
rect 71 222 72 223 
<< m2c >>
rect 71 222 72 223 
<< m1 >>
rect 71 222 72 223 
<< m2 >>
rect 71 222 72 223 
<< m2 >>
rect 72 222 73 223 
<< m1 >>
rect 73 222 74 223 
<< m2 >>
rect 73 222 74 223 
<< m2 >>
rect 74 222 75 223 
<< m1 >>
rect 89 222 90 223 
<< m2 >>
rect 89 222 90 223 
<< m2c >>
rect 89 222 90 223 
<< m1 >>
rect 89 222 90 223 
<< m2 >>
rect 89 222 90 223 
<< m1 >>
rect 91 222 92 223 
<< m2 >>
rect 91 222 92 223 
<< m2c >>
rect 91 222 92 223 
<< m1 >>
rect 91 222 92 223 
<< m2 >>
rect 91 222 92 223 
<< m1 >>
rect 95 222 96 223 
<< m2 >>
rect 95 222 96 223 
<< m2c >>
rect 95 222 96 223 
<< m1 >>
rect 95 222 96 223 
<< m2 >>
rect 95 222 96 223 
<< m1 >>
rect 102 222 103 223 
<< m1 >>
rect 103 222 104 223 
<< m1 >>
rect 104 222 105 223 
<< m1 >>
rect 105 222 106 223 
<< m1 >>
rect 106 222 107 223 
<< m1 >>
rect 107 222 108 223 
<< m1 >>
rect 108 222 109 223 
<< m1 >>
rect 109 222 110 223 
<< m1 >>
rect 110 222 111 223 
<< m1 >>
rect 111 222 112 223 
<< m2 >>
rect 111 222 112 223 
<< m1 >>
rect 112 222 113 223 
<< m1 >>
rect 113 222 114 223 
<< m2 >>
rect 113 222 114 223 
<< m2c >>
rect 113 222 114 223 
<< m1 >>
rect 113 222 114 223 
<< m2 >>
rect 113 222 114 223 
<< m1 >>
rect 139 222 140 223 
<< m1 >>
rect 150 222 151 223 
<< m2 >>
rect 150 222 151 223 
<< m2c >>
rect 150 222 151 223 
<< m1 >>
rect 150 222 151 223 
<< m2 >>
rect 150 222 151 223 
<< m1 >>
rect 156 222 157 223 
<< m1 >>
rect 157 222 158 223 
<< m1 >>
rect 158 222 159 223 
<< m1 >>
rect 159 222 160 223 
<< m1 >>
rect 160 222 161 223 
<< m1 >>
rect 161 222 162 223 
<< m1 >>
rect 162 222 163 223 
<< m1 >>
rect 163 222 164 223 
<< m1 >>
rect 164 222 165 223 
<< m1 >>
rect 165 222 166 223 
<< m1 >>
rect 166 222 167 223 
<< m1 >>
rect 167 222 168 223 
<< m1 >>
rect 168 222 169 223 
<< m1 >>
rect 169 222 170 223 
<< m1 >>
rect 170 222 171 223 
<< m1 >>
rect 171 222 172 223 
<< m1 >>
rect 172 222 173 223 
<< m1 >>
rect 173 222 174 223 
<< m1 >>
rect 174 222 175 223 
<< m1 >>
rect 175 222 176 223 
<< m1 >>
rect 176 222 177 223 
<< m1 >>
rect 177 222 178 223 
<< m1 >>
rect 178 222 179 223 
<< m1 >>
rect 179 222 180 223 
<< m1 >>
rect 180 222 181 223 
<< m1 >>
rect 181 222 182 223 
<< m1 >>
rect 182 222 183 223 
<< m1 >>
rect 183 222 184 223 
<< m1 >>
rect 184 222 185 223 
<< m1 >>
rect 185 222 186 223 
<< m1 >>
rect 186 222 187 223 
<< m1 >>
rect 187 222 188 223 
<< m1 >>
rect 188 222 189 223 
<< m2 >>
rect 188 222 189 223 
<< m2c >>
rect 188 222 189 223 
<< m1 >>
rect 188 222 189 223 
<< m2 >>
rect 188 222 189 223 
<< m2 >>
rect 189 222 190 223 
<< m1 >>
rect 190 222 191 223 
<< m2 >>
rect 190 222 191 223 
<< m2 >>
rect 191 222 192 223 
<< m1 >>
rect 16 223 17 224 
<< m1 >>
rect 19 223 20 224 
<< m2 >>
rect 19 223 20 224 
<< m2c >>
rect 19 223 20 224 
<< m1 >>
rect 19 223 20 224 
<< m2 >>
rect 19 223 20 224 
<< m1 >>
rect 24 223 25 224 
<< m2 >>
rect 24 223 25 224 
<< m2c >>
rect 24 223 25 224 
<< m1 >>
rect 24 223 25 224 
<< m2 >>
rect 24 223 25 224 
<< m1 >>
rect 28 223 29 224 
<< m1 >>
rect 46 223 47 224 
<< m2 >>
rect 46 223 47 224 
<< m1 >>
rect 52 223 53 224 
<< m1 >>
rect 71 223 72 224 
<< m1 >>
rect 73 223 74 224 
<< m1 >>
rect 89 223 90 224 
<< m1 >>
rect 91 223 92 224 
<< m2 >>
rect 95 223 96 224 
<< m1 >>
rect 102 223 103 224 
<< m2 >>
rect 111 223 112 224 
<< m1 >>
rect 137 223 138 224 
<< m2 >>
rect 137 223 138 224 
<< m2c >>
rect 137 223 138 224 
<< m1 >>
rect 137 223 138 224 
<< m2 >>
rect 137 223 138 224 
<< m2 >>
rect 138 223 139 224 
<< m1 >>
rect 139 223 140 224 
<< m2 >>
rect 139 223 140 224 
<< m2 >>
rect 140 223 141 224 
<< m1 >>
rect 150 223 151 224 
<< m1 >>
rect 156 223 157 224 
<< m1 >>
rect 190 223 191 224 
<< m1 >>
rect 16 224 17 225 
<< m2 >>
rect 19 224 20 225 
<< m2 >>
rect 24 224 25 225 
<< m1 >>
rect 28 224 29 225 
<< m1 >>
rect 46 224 47 225 
<< m2 >>
rect 46 224 47 225 
<< m1 >>
rect 52 224 53 225 
<< m1 >>
rect 71 224 72 225 
<< m1 >>
rect 73 224 74 225 
<< m1 >>
rect 89 224 90 225 
<< m2 >>
rect 89 224 90 225 
<< m2c >>
rect 89 224 90 225 
<< m1 >>
rect 89 224 90 225 
<< m2 >>
rect 89 224 90 225 
<< m2 >>
rect 90 224 91 225 
<< m1 >>
rect 91 224 92 225 
<< m2 >>
rect 91 224 92 225 
<< m2 >>
rect 92 224 93 225 
<< m1 >>
rect 93 224 94 225 
<< m2 >>
rect 93 224 94 225 
<< m2c >>
rect 93 224 94 225 
<< m1 >>
rect 93 224 94 225 
<< m2 >>
rect 93 224 94 225 
<< m1 >>
rect 94 224 95 225 
<< m1 >>
rect 95 224 96 225 
<< m2 >>
rect 95 224 96 225 
<< m1 >>
rect 96 224 97 225 
<< m1 >>
rect 97 224 98 225 
<< m1 >>
rect 98 224 99 225 
<< m1 >>
rect 99 224 100 225 
<< m1 >>
rect 100 224 101 225 
<< m1 >>
rect 101 224 102 225 
<< m1 >>
rect 102 224 103 225 
<< m1 >>
rect 111 224 112 225 
<< m2 >>
rect 111 224 112 225 
<< m2c >>
rect 111 224 112 225 
<< m1 >>
rect 111 224 112 225 
<< m2 >>
rect 111 224 112 225 
<< m1 >>
rect 112 224 113 225 
<< m1 >>
rect 113 224 114 225 
<< m1 >>
rect 114 224 115 225 
<< m1 >>
rect 115 224 116 225 
<< m1 >>
rect 116 224 117 225 
<< m1 >>
rect 117 224 118 225 
<< m1 >>
rect 118 224 119 225 
<< m1 >>
rect 119 224 120 225 
<< m1 >>
rect 120 224 121 225 
<< m1 >>
rect 121 224 122 225 
<< m1 >>
rect 122 224 123 225 
<< m1 >>
rect 123 224 124 225 
<< m1 >>
rect 124 224 125 225 
<< m1 >>
rect 125 224 126 225 
<< m1 >>
rect 126 224 127 225 
<< m1 >>
rect 127 224 128 225 
<< m1 >>
rect 128 224 129 225 
<< m1 >>
rect 129 224 130 225 
<< m1 >>
rect 130 224 131 225 
<< m1 >>
rect 131 224 132 225 
<< m1 >>
rect 132 224 133 225 
<< m1 >>
rect 133 224 134 225 
<< m1 >>
rect 134 224 135 225 
<< m1 >>
rect 135 224 136 225 
<< m1 >>
rect 136 224 137 225 
<< m1 >>
rect 137 224 138 225 
<< m1 >>
rect 139 224 140 225 
<< m2 >>
rect 140 224 141 225 
<< m1 >>
rect 141 224 142 225 
<< m2 >>
rect 141 224 142 225 
<< m2c >>
rect 141 224 142 225 
<< m1 >>
rect 141 224 142 225 
<< m2 >>
rect 141 224 142 225 
<< m1 >>
rect 142 224 143 225 
<< m1 >>
rect 143 224 144 225 
<< m1 >>
rect 144 224 145 225 
<< m1 >>
rect 145 224 146 225 
<< m1 >>
rect 146 224 147 225 
<< m1 >>
rect 147 224 148 225 
<< m1 >>
rect 148 224 149 225 
<< m2 >>
rect 148 224 149 225 
<< m2c >>
rect 148 224 149 225 
<< m1 >>
rect 148 224 149 225 
<< m2 >>
rect 148 224 149 225 
<< m2 >>
rect 149 224 150 225 
<< m1 >>
rect 150 224 151 225 
<< m2 >>
rect 150 224 151 225 
<< m2 >>
rect 151 224 152 225 
<< m1 >>
rect 152 224 153 225 
<< m2 >>
rect 152 224 153 225 
<< m2c >>
rect 152 224 153 225 
<< m1 >>
rect 152 224 153 225 
<< m2 >>
rect 152 224 153 225 
<< m1 >>
rect 153 224 154 225 
<< m1 >>
rect 154 224 155 225 
<< m1 >>
rect 155 224 156 225 
<< m1 >>
rect 156 224 157 225 
<< m1 >>
rect 190 224 191 225 
<< m1 >>
rect 16 225 17 226 
<< m1 >>
rect 17 225 18 226 
<< m1 >>
rect 18 225 19 226 
<< m1 >>
rect 19 225 20 226 
<< m2 >>
rect 19 225 20 226 
<< m1 >>
rect 20 225 21 226 
<< m1 >>
rect 21 225 22 226 
<< m1 >>
rect 22 225 23 226 
<< m1 >>
rect 23 225 24 226 
<< m1 >>
rect 24 225 25 226 
<< m2 >>
rect 24 225 25 226 
<< m1 >>
rect 25 225 26 226 
<< m1 >>
rect 26 225 27 226 
<< m1 >>
rect 28 225 29 226 
<< m1 >>
rect 46 225 47 226 
<< m2 >>
rect 46 225 47 226 
<< m1 >>
rect 52 225 53 226 
<< m1 >>
rect 71 225 72 226 
<< m1 >>
rect 73 225 74 226 
<< m1 >>
rect 91 225 92 226 
<< m2 >>
rect 95 225 96 226 
<< m1 >>
rect 139 225 140 226 
<< m1 >>
rect 150 225 151 226 
<< m1 >>
rect 190 225 191 226 
<< m2 >>
rect 19 226 20 227 
<< m2 >>
rect 24 226 25 227 
<< m1 >>
rect 26 226 27 227 
<< m1 >>
rect 28 226 29 227 
<< m1 >>
rect 46 226 47 227 
<< m2 >>
rect 46 226 47 227 
<< m1 >>
rect 52 226 53 227 
<< m1 >>
rect 71 226 72 227 
<< m1 >>
rect 73 226 74 227 
<< m1 >>
rect 91 226 92 227 
<< m1 >>
rect 95 226 96 227 
<< m2 >>
rect 95 226 96 227 
<< m2c >>
rect 95 226 96 227 
<< m1 >>
rect 95 226 96 227 
<< m2 >>
rect 95 226 96 227 
<< m1 >>
rect 139 226 140 227 
<< m1 >>
rect 150 226 151 227 
<< m1 >>
rect 190 226 191 227 
<< m1 >>
rect 191 226 192 227 
<< m1 >>
rect 192 226 193 227 
<< m1 >>
rect 193 226 194 227 
<< m1 >>
rect 194 226 195 227 
<< m1 >>
rect 195 226 196 227 
<< m1 >>
rect 196 226 197 227 
<< m1 >>
rect 197 226 198 227 
<< m1 >>
rect 198 226 199 227 
<< m1 >>
rect 199 226 200 227 
<< m1 >>
rect 200 226 201 227 
<< m1 >>
rect 201 226 202 227 
<< m1 >>
rect 202 226 203 227 
<< m1 >>
rect 203 226 204 227 
<< m1 >>
rect 204 226 205 227 
<< m1 >>
rect 205 226 206 227 
<< m1 >>
rect 206 226 207 227 
<< m1 >>
rect 207 226 208 227 
<< m1 >>
rect 208 226 209 227 
<< m1 >>
rect 209 226 210 227 
<< m1 >>
rect 210 226 211 227 
<< m1 >>
rect 211 226 212 227 
<< m1 >>
rect 19 227 20 228 
<< m2 >>
rect 19 227 20 228 
<< m2c >>
rect 19 227 20 228 
<< m1 >>
rect 19 227 20 228 
<< m2 >>
rect 19 227 20 228 
<< m1 >>
rect 24 227 25 228 
<< m2 >>
rect 24 227 25 228 
<< m2c >>
rect 24 227 25 228 
<< m1 >>
rect 24 227 25 228 
<< m2 >>
rect 24 227 25 228 
<< m1 >>
rect 26 227 27 228 
<< m1 >>
rect 28 227 29 228 
<< m1 >>
rect 46 227 47 228 
<< m2 >>
rect 46 227 47 228 
<< m1 >>
rect 52 227 53 228 
<< m1 >>
rect 71 227 72 228 
<< m1 >>
rect 73 227 74 228 
<< m1 >>
rect 91 227 92 228 
<< m1 >>
rect 95 227 96 228 
<< m1 >>
rect 139 227 140 228 
<< m1 >>
rect 150 227 151 228 
<< m1 >>
rect 211 227 212 228 
<< pdiffusion >>
rect 12 228 13 229 
<< pdiffusion >>
rect 13 228 14 229 
<< pdiffusion >>
rect 14 228 15 229 
<< pdiffusion >>
rect 15 228 16 229 
<< pdiffusion >>
rect 16 228 17 229 
<< pdiffusion >>
rect 17 228 18 229 
<< m1 >>
rect 19 228 20 229 
<< m1 >>
rect 24 228 25 229 
<< m1 >>
rect 26 228 27 229 
<< m1 >>
rect 28 228 29 229 
<< pdiffusion >>
rect 30 228 31 229 
<< pdiffusion >>
rect 31 228 32 229 
<< pdiffusion >>
rect 32 228 33 229 
<< pdiffusion >>
rect 33 228 34 229 
<< pdiffusion >>
rect 34 228 35 229 
<< pdiffusion >>
rect 35 228 36 229 
<< m1 >>
rect 46 228 47 229 
<< m2 >>
rect 46 228 47 229 
<< pdiffusion >>
rect 48 228 49 229 
<< pdiffusion >>
rect 49 228 50 229 
<< pdiffusion >>
rect 50 228 51 229 
<< pdiffusion >>
rect 51 228 52 229 
<< m1 >>
rect 52 228 53 229 
<< pdiffusion >>
rect 52 228 53 229 
<< pdiffusion >>
rect 53 228 54 229 
<< m1 >>
rect 71 228 72 229 
<< m1 >>
rect 73 228 74 229 
<< pdiffusion >>
rect 84 228 85 229 
<< pdiffusion >>
rect 85 228 86 229 
<< pdiffusion >>
rect 86 228 87 229 
<< pdiffusion >>
rect 87 228 88 229 
<< pdiffusion >>
rect 88 228 89 229 
<< pdiffusion >>
rect 89 228 90 229 
<< m1 >>
rect 91 228 92 229 
<< m1 >>
rect 95 228 96 229 
<< pdiffusion >>
rect 102 228 103 229 
<< pdiffusion >>
rect 103 228 104 229 
<< pdiffusion >>
rect 104 228 105 229 
<< pdiffusion >>
rect 105 228 106 229 
<< pdiffusion >>
rect 106 228 107 229 
<< pdiffusion >>
rect 107 228 108 229 
<< pdiffusion >>
rect 138 228 139 229 
<< m1 >>
rect 139 228 140 229 
<< pdiffusion >>
rect 139 228 140 229 
<< pdiffusion >>
rect 140 228 141 229 
<< pdiffusion >>
rect 141 228 142 229 
<< pdiffusion >>
rect 142 228 143 229 
<< pdiffusion >>
rect 143 228 144 229 
<< m1 >>
rect 150 228 151 229 
<< pdiffusion >>
rect 156 228 157 229 
<< pdiffusion >>
rect 157 228 158 229 
<< pdiffusion >>
rect 158 228 159 229 
<< pdiffusion >>
rect 159 228 160 229 
<< pdiffusion >>
rect 160 228 161 229 
<< pdiffusion >>
rect 161 228 162 229 
<< pdiffusion >>
rect 210 228 211 229 
<< m1 >>
rect 211 228 212 229 
<< pdiffusion >>
rect 211 228 212 229 
<< pdiffusion >>
rect 212 228 213 229 
<< pdiffusion >>
rect 213 228 214 229 
<< pdiffusion >>
rect 214 228 215 229 
<< pdiffusion >>
rect 215 228 216 229 
<< pdiffusion >>
rect 228 228 229 229 
<< pdiffusion >>
rect 229 228 230 229 
<< pdiffusion >>
rect 230 228 231 229 
<< pdiffusion >>
rect 231 228 232 229 
<< pdiffusion >>
rect 232 228 233 229 
<< pdiffusion >>
rect 233 228 234 229 
<< pdiffusion >>
rect 12 229 13 230 
<< pdiffusion >>
rect 13 229 14 230 
<< pdiffusion >>
rect 14 229 15 230 
<< pdiffusion >>
rect 15 229 16 230 
<< pdiffusion >>
rect 16 229 17 230 
<< pdiffusion >>
rect 17 229 18 230 
<< m1 >>
rect 19 229 20 230 
<< m1 >>
rect 24 229 25 230 
<< m1 >>
rect 26 229 27 230 
<< m1 >>
rect 28 229 29 230 
<< pdiffusion >>
rect 30 229 31 230 
<< pdiffusion >>
rect 31 229 32 230 
<< pdiffusion >>
rect 32 229 33 230 
<< pdiffusion >>
rect 33 229 34 230 
<< pdiffusion >>
rect 34 229 35 230 
<< pdiffusion >>
rect 35 229 36 230 
<< m1 >>
rect 46 229 47 230 
<< m2 >>
rect 46 229 47 230 
<< pdiffusion >>
rect 48 229 49 230 
<< pdiffusion >>
rect 49 229 50 230 
<< pdiffusion >>
rect 50 229 51 230 
<< pdiffusion >>
rect 51 229 52 230 
<< pdiffusion >>
rect 52 229 53 230 
<< pdiffusion >>
rect 53 229 54 230 
<< m1 >>
rect 71 229 72 230 
<< m1 >>
rect 73 229 74 230 
<< pdiffusion >>
rect 84 229 85 230 
<< pdiffusion >>
rect 85 229 86 230 
<< pdiffusion >>
rect 86 229 87 230 
<< pdiffusion >>
rect 87 229 88 230 
<< pdiffusion >>
rect 88 229 89 230 
<< pdiffusion >>
rect 89 229 90 230 
<< m1 >>
rect 91 229 92 230 
<< m1 >>
rect 95 229 96 230 
<< pdiffusion >>
rect 102 229 103 230 
<< pdiffusion >>
rect 103 229 104 230 
<< pdiffusion >>
rect 104 229 105 230 
<< pdiffusion >>
rect 105 229 106 230 
<< pdiffusion >>
rect 106 229 107 230 
<< pdiffusion >>
rect 107 229 108 230 
<< pdiffusion >>
rect 138 229 139 230 
<< pdiffusion >>
rect 139 229 140 230 
<< pdiffusion >>
rect 140 229 141 230 
<< pdiffusion >>
rect 141 229 142 230 
<< pdiffusion >>
rect 142 229 143 230 
<< pdiffusion >>
rect 143 229 144 230 
<< m1 >>
rect 150 229 151 230 
<< pdiffusion >>
rect 156 229 157 230 
<< pdiffusion >>
rect 157 229 158 230 
<< pdiffusion >>
rect 158 229 159 230 
<< pdiffusion >>
rect 159 229 160 230 
<< pdiffusion >>
rect 160 229 161 230 
<< pdiffusion >>
rect 161 229 162 230 
<< pdiffusion >>
rect 210 229 211 230 
<< pdiffusion >>
rect 211 229 212 230 
<< pdiffusion >>
rect 212 229 213 230 
<< pdiffusion >>
rect 213 229 214 230 
<< pdiffusion >>
rect 214 229 215 230 
<< pdiffusion >>
rect 215 229 216 230 
<< pdiffusion >>
rect 228 229 229 230 
<< pdiffusion >>
rect 229 229 230 230 
<< pdiffusion >>
rect 230 229 231 230 
<< pdiffusion >>
rect 231 229 232 230 
<< pdiffusion >>
rect 232 229 233 230 
<< pdiffusion >>
rect 233 229 234 230 
<< pdiffusion >>
rect 12 230 13 231 
<< pdiffusion >>
rect 13 230 14 231 
<< pdiffusion >>
rect 14 230 15 231 
<< pdiffusion >>
rect 15 230 16 231 
<< pdiffusion >>
rect 16 230 17 231 
<< pdiffusion >>
rect 17 230 18 231 
<< m1 >>
rect 19 230 20 231 
<< m1 >>
rect 24 230 25 231 
<< m1 >>
rect 26 230 27 231 
<< m1 >>
rect 28 230 29 231 
<< pdiffusion >>
rect 30 230 31 231 
<< pdiffusion >>
rect 31 230 32 231 
<< pdiffusion >>
rect 32 230 33 231 
<< pdiffusion >>
rect 33 230 34 231 
<< pdiffusion >>
rect 34 230 35 231 
<< pdiffusion >>
rect 35 230 36 231 
<< m1 >>
rect 46 230 47 231 
<< m2 >>
rect 46 230 47 231 
<< pdiffusion >>
rect 48 230 49 231 
<< pdiffusion >>
rect 49 230 50 231 
<< pdiffusion >>
rect 50 230 51 231 
<< pdiffusion >>
rect 51 230 52 231 
<< pdiffusion >>
rect 52 230 53 231 
<< pdiffusion >>
rect 53 230 54 231 
<< m1 >>
rect 71 230 72 231 
<< m1 >>
rect 73 230 74 231 
<< pdiffusion >>
rect 84 230 85 231 
<< pdiffusion >>
rect 85 230 86 231 
<< pdiffusion >>
rect 86 230 87 231 
<< pdiffusion >>
rect 87 230 88 231 
<< pdiffusion >>
rect 88 230 89 231 
<< pdiffusion >>
rect 89 230 90 231 
<< m1 >>
rect 91 230 92 231 
<< m1 >>
rect 95 230 96 231 
<< pdiffusion >>
rect 102 230 103 231 
<< pdiffusion >>
rect 103 230 104 231 
<< pdiffusion >>
rect 104 230 105 231 
<< pdiffusion >>
rect 105 230 106 231 
<< pdiffusion >>
rect 106 230 107 231 
<< pdiffusion >>
rect 107 230 108 231 
<< pdiffusion >>
rect 138 230 139 231 
<< pdiffusion >>
rect 139 230 140 231 
<< pdiffusion >>
rect 140 230 141 231 
<< pdiffusion >>
rect 141 230 142 231 
<< pdiffusion >>
rect 142 230 143 231 
<< pdiffusion >>
rect 143 230 144 231 
<< m1 >>
rect 150 230 151 231 
<< pdiffusion >>
rect 156 230 157 231 
<< pdiffusion >>
rect 157 230 158 231 
<< pdiffusion >>
rect 158 230 159 231 
<< pdiffusion >>
rect 159 230 160 231 
<< pdiffusion >>
rect 160 230 161 231 
<< pdiffusion >>
rect 161 230 162 231 
<< pdiffusion >>
rect 210 230 211 231 
<< pdiffusion >>
rect 211 230 212 231 
<< pdiffusion >>
rect 212 230 213 231 
<< pdiffusion >>
rect 213 230 214 231 
<< pdiffusion >>
rect 214 230 215 231 
<< pdiffusion >>
rect 215 230 216 231 
<< pdiffusion >>
rect 228 230 229 231 
<< pdiffusion >>
rect 229 230 230 231 
<< pdiffusion >>
rect 230 230 231 231 
<< pdiffusion >>
rect 231 230 232 231 
<< pdiffusion >>
rect 232 230 233 231 
<< pdiffusion >>
rect 233 230 234 231 
<< pdiffusion >>
rect 12 231 13 232 
<< pdiffusion >>
rect 13 231 14 232 
<< pdiffusion >>
rect 14 231 15 232 
<< pdiffusion >>
rect 15 231 16 232 
<< pdiffusion >>
rect 16 231 17 232 
<< pdiffusion >>
rect 17 231 18 232 
<< m1 >>
rect 19 231 20 232 
<< m1 >>
rect 24 231 25 232 
<< m1 >>
rect 26 231 27 232 
<< m1 >>
rect 28 231 29 232 
<< pdiffusion >>
rect 30 231 31 232 
<< pdiffusion >>
rect 31 231 32 232 
<< pdiffusion >>
rect 32 231 33 232 
<< pdiffusion >>
rect 33 231 34 232 
<< pdiffusion >>
rect 34 231 35 232 
<< pdiffusion >>
rect 35 231 36 232 
<< m1 >>
rect 46 231 47 232 
<< m2 >>
rect 46 231 47 232 
<< pdiffusion >>
rect 48 231 49 232 
<< pdiffusion >>
rect 49 231 50 232 
<< pdiffusion >>
rect 50 231 51 232 
<< pdiffusion >>
rect 51 231 52 232 
<< pdiffusion >>
rect 52 231 53 232 
<< pdiffusion >>
rect 53 231 54 232 
<< m1 >>
rect 71 231 72 232 
<< m1 >>
rect 73 231 74 232 
<< pdiffusion >>
rect 84 231 85 232 
<< pdiffusion >>
rect 85 231 86 232 
<< pdiffusion >>
rect 86 231 87 232 
<< pdiffusion >>
rect 87 231 88 232 
<< pdiffusion >>
rect 88 231 89 232 
<< pdiffusion >>
rect 89 231 90 232 
<< m1 >>
rect 91 231 92 232 
<< m1 >>
rect 95 231 96 232 
<< pdiffusion >>
rect 102 231 103 232 
<< pdiffusion >>
rect 103 231 104 232 
<< pdiffusion >>
rect 104 231 105 232 
<< pdiffusion >>
rect 105 231 106 232 
<< pdiffusion >>
rect 106 231 107 232 
<< pdiffusion >>
rect 107 231 108 232 
<< pdiffusion >>
rect 138 231 139 232 
<< pdiffusion >>
rect 139 231 140 232 
<< pdiffusion >>
rect 140 231 141 232 
<< pdiffusion >>
rect 141 231 142 232 
<< pdiffusion >>
rect 142 231 143 232 
<< pdiffusion >>
rect 143 231 144 232 
<< m1 >>
rect 150 231 151 232 
<< pdiffusion >>
rect 156 231 157 232 
<< pdiffusion >>
rect 157 231 158 232 
<< pdiffusion >>
rect 158 231 159 232 
<< pdiffusion >>
rect 159 231 160 232 
<< pdiffusion >>
rect 160 231 161 232 
<< pdiffusion >>
rect 161 231 162 232 
<< pdiffusion >>
rect 210 231 211 232 
<< pdiffusion >>
rect 211 231 212 232 
<< pdiffusion >>
rect 212 231 213 232 
<< pdiffusion >>
rect 213 231 214 232 
<< pdiffusion >>
rect 214 231 215 232 
<< pdiffusion >>
rect 215 231 216 232 
<< pdiffusion >>
rect 228 231 229 232 
<< pdiffusion >>
rect 229 231 230 232 
<< pdiffusion >>
rect 230 231 231 232 
<< pdiffusion >>
rect 231 231 232 232 
<< pdiffusion >>
rect 232 231 233 232 
<< pdiffusion >>
rect 233 231 234 232 
<< pdiffusion >>
rect 12 232 13 233 
<< pdiffusion >>
rect 13 232 14 233 
<< pdiffusion >>
rect 14 232 15 233 
<< pdiffusion >>
rect 15 232 16 233 
<< pdiffusion >>
rect 16 232 17 233 
<< pdiffusion >>
rect 17 232 18 233 
<< m1 >>
rect 19 232 20 233 
<< m1 >>
rect 24 232 25 233 
<< m1 >>
rect 26 232 27 233 
<< m1 >>
rect 28 232 29 233 
<< pdiffusion >>
rect 30 232 31 233 
<< pdiffusion >>
rect 31 232 32 233 
<< pdiffusion >>
rect 32 232 33 233 
<< pdiffusion >>
rect 33 232 34 233 
<< pdiffusion >>
rect 34 232 35 233 
<< pdiffusion >>
rect 35 232 36 233 
<< m1 >>
rect 46 232 47 233 
<< m2 >>
rect 46 232 47 233 
<< pdiffusion >>
rect 48 232 49 233 
<< pdiffusion >>
rect 49 232 50 233 
<< pdiffusion >>
rect 50 232 51 233 
<< pdiffusion >>
rect 51 232 52 233 
<< pdiffusion >>
rect 52 232 53 233 
<< pdiffusion >>
rect 53 232 54 233 
<< m1 >>
rect 71 232 72 233 
<< m1 >>
rect 73 232 74 233 
<< pdiffusion >>
rect 84 232 85 233 
<< pdiffusion >>
rect 85 232 86 233 
<< pdiffusion >>
rect 86 232 87 233 
<< pdiffusion >>
rect 87 232 88 233 
<< pdiffusion >>
rect 88 232 89 233 
<< pdiffusion >>
rect 89 232 90 233 
<< m1 >>
rect 91 232 92 233 
<< m1 >>
rect 95 232 96 233 
<< pdiffusion >>
rect 102 232 103 233 
<< pdiffusion >>
rect 103 232 104 233 
<< pdiffusion >>
rect 104 232 105 233 
<< pdiffusion >>
rect 105 232 106 233 
<< pdiffusion >>
rect 106 232 107 233 
<< pdiffusion >>
rect 107 232 108 233 
<< pdiffusion >>
rect 138 232 139 233 
<< pdiffusion >>
rect 139 232 140 233 
<< pdiffusion >>
rect 140 232 141 233 
<< pdiffusion >>
rect 141 232 142 233 
<< pdiffusion >>
rect 142 232 143 233 
<< pdiffusion >>
rect 143 232 144 233 
<< m1 >>
rect 150 232 151 233 
<< pdiffusion >>
rect 156 232 157 233 
<< pdiffusion >>
rect 157 232 158 233 
<< pdiffusion >>
rect 158 232 159 233 
<< pdiffusion >>
rect 159 232 160 233 
<< pdiffusion >>
rect 160 232 161 233 
<< pdiffusion >>
rect 161 232 162 233 
<< pdiffusion >>
rect 210 232 211 233 
<< pdiffusion >>
rect 211 232 212 233 
<< pdiffusion >>
rect 212 232 213 233 
<< pdiffusion >>
rect 213 232 214 233 
<< pdiffusion >>
rect 214 232 215 233 
<< pdiffusion >>
rect 215 232 216 233 
<< pdiffusion >>
rect 228 232 229 233 
<< pdiffusion >>
rect 229 232 230 233 
<< pdiffusion >>
rect 230 232 231 233 
<< pdiffusion >>
rect 231 232 232 233 
<< pdiffusion >>
rect 232 232 233 233 
<< pdiffusion >>
rect 233 232 234 233 
<< pdiffusion >>
rect 12 233 13 234 
<< m1 >>
rect 13 233 14 234 
<< pdiffusion >>
rect 13 233 14 234 
<< pdiffusion >>
rect 14 233 15 234 
<< pdiffusion >>
rect 15 233 16 234 
<< pdiffusion >>
rect 16 233 17 234 
<< pdiffusion >>
rect 17 233 18 234 
<< m1 >>
rect 19 233 20 234 
<< m1 >>
rect 24 233 25 234 
<< m1 >>
rect 26 233 27 234 
<< m1 >>
rect 28 233 29 234 
<< pdiffusion >>
rect 30 233 31 234 
<< pdiffusion >>
rect 31 233 32 234 
<< pdiffusion >>
rect 32 233 33 234 
<< pdiffusion >>
rect 33 233 34 234 
<< m1 >>
rect 34 233 35 234 
<< pdiffusion >>
rect 34 233 35 234 
<< pdiffusion >>
rect 35 233 36 234 
<< m1 >>
rect 46 233 47 234 
<< m2 >>
rect 46 233 47 234 
<< pdiffusion >>
rect 48 233 49 234 
<< pdiffusion >>
rect 49 233 50 234 
<< pdiffusion >>
rect 50 233 51 234 
<< pdiffusion >>
rect 51 233 52 234 
<< pdiffusion >>
rect 52 233 53 234 
<< pdiffusion >>
rect 53 233 54 234 
<< m1 >>
rect 71 233 72 234 
<< m1 >>
rect 73 233 74 234 
<< pdiffusion >>
rect 84 233 85 234 
<< pdiffusion >>
rect 85 233 86 234 
<< pdiffusion >>
rect 86 233 87 234 
<< pdiffusion >>
rect 87 233 88 234 
<< m1 >>
rect 88 233 89 234 
<< pdiffusion >>
rect 88 233 89 234 
<< pdiffusion >>
rect 89 233 90 234 
<< m1 >>
rect 91 233 92 234 
<< m1 >>
rect 95 233 96 234 
<< pdiffusion >>
rect 102 233 103 234 
<< pdiffusion >>
rect 103 233 104 234 
<< pdiffusion >>
rect 104 233 105 234 
<< pdiffusion >>
rect 105 233 106 234 
<< pdiffusion >>
rect 106 233 107 234 
<< pdiffusion >>
rect 107 233 108 234 
<< pdiffusion >>
rect 138 233 139 234 
<< pdiffusion >>
rect 139 233 140 234 
<< pdiffusion >>
rect 140 233 141 234 
<< pdiffusion >>
rect 141 233 142 234 
<< m1 >>
rect 142 233 143 234 
<< pdiffusion >>
rect 142 233 143 234 
<< pdiffusion >>
rect 143 233 144 234 
<< m1 >>
rect 150 233 151 234 
<< pdiffusion >>
rect 156 233 157 234 
<< pdiffusion >>
rect 157 233 158 234 
<< pdiffusion >>
rect 158 233 159 234 
<< pdiffusion >>
rect 159 233 160 234 
<< pdiffusion >>
rect 160 233 161 234 
<< pdiffusion >>
rect 161 233 162 234 
<< pdiffusion >>
rect 210 233 211 234 
<< pdiffusion >>
rect 211 233 212 234 
<< pdiffusion >>
rect 212 233 213 234 
<< pdiffusion >>
rect 213 233 214 234 
<< pdiffusion >>
rect 214 233 215 234 
<< pdiffusion >>
rect 215 233 216 234 
<< pdiffusion >>
rect 228 233 229 234 
<< pdiffusion >>
rect 229 233 230 234 
<< pdiffusion >>
rect 230 233 231 234 
<< pdiffusion >>
rect 231 233 232 234 
<< pdiffusion >>
rect 232 233 233 234 
<< pdiffusion >>
rect 233 233 234 234 
<< m1 >>
rect 13 234 14 235 
<< m1 >>
rect 19 234 20 235 
<< m2 >>
rect 19 234 20 235 
<< m2c >>
rect 19 234 20 235 
<< m1 >>
rect 19 234 20 235 
<< m2 >>
rect 19 234 20 235 
<< m1 >>
rect 24 234 25 235 
<< m2 >>
rect 24 234 25 235 
<< m2c >>
rect 24 234 25 235 
<< m1 >>
rect 24 234 25 235 
<< m2 >>
rect 24 234 25 235 
<< m1 >>
rect 26 234 27 235 
<< m2 >>
rect 26 234 27 235 
<< m2c >>
rect 26 234 27 235 
<< m1 >>
rect 26 234 27 235 
<< m2 >>
rect 26 234 27 235 
<< m2 >>
rect 27 234 28 235 
<< m1 >>
rect 28 234 29 235 
<< m2 >>
rect 28 234 29 235 
<< m1 >>
rect 34 234 35 235 
<< m2 >>
rect 34 234 35 235 
<< m2c >>
rect 34 234 35 235 
<< m1 >>
rect 34 234 35 235 
<< m2 >>
rect 34 234 35 235 
<< m1 >>
rect 46 234 47 235 
<< m2 >>
rect 46 234 47 235 
<< m1 >>
rect 71 234 72 235 
<< m1 >>
rect 73 234 74 235 
<< m1 >>
rect 88 234 89 235 
<< m1 >>
rect 91 234 92 235 
<< m1 >>
rect 95 234 96 235 
<< m1 >>
rect 142 234 143 235 
<< m1 >>
rect 150 234 151 235 
<< m1 >>
rect 13 235 14 236 
<< m1 >>
rect 14 235 15 236 
<< m2 >>
rect 14 235 15 236 
<< m2c >>
rect 14 235 15 236 
<< m1 >>
rect 14 235 15 236 
<< m2 >>
rect 14 235 15 236 
<< m2 >>
rect 15 235 16 236 
<< m2 >>
rect 19 235 20 236 
<< m2 >>
rect 20 235 21 236 
<< m2 >>
rect 24 235 25 236 
<< m1 >>
rect 28 235 29 236 
<< m2 >>
rect 28 235 29 236 
<< m2 >>
rect 34 235 35 236 
<< m2 >>
rect 35 235 36 236 
<< m2 >>
rect 36 235 37 236 
<< m2 >>
rect 37 235 38 236 
<< m2 >>
rect 38 235 39 236 
<< m2 >>
rect 39 235 40 236 
<< m2 >>
rect 40 235 41 236 
<< m2 >>
rect 41 235 42 236 
<< m2 >>
rect 42 235 43 236 
<< m2 >>
rect 43 235 44 236 
<< m2 >>
rect 44 235 45 236 
<< m2 >>
rect 45 235 46 236 
<< m1 >>
rect 46 235 47 236 
<< m2 >>
rect 46 235 47 236 
<< m1 >>
rect 71 235 72 236 
<< m1 >>
rect 73 235 74 236 
<< m1 >>
rect 88 235 89 236 
<< m1 >>
rect 89 235 90 236 
<< m2 >>
rect 89 235 90 236 
<< m2c >>
rect 89 235 90 236 
<< m1 >>
rect 89 235 90 236 
<< m2 >>
rect 89 235 90 236 
<< m2 >>
rect 90 235 91 236 
<< m1 >>
rect 91 235 92 236 
<< m2 >>
rect 91 235 92 236 
<< m2 >>
rect 92 235 93 236 
<< m1 >>
rect 93 235 94 236 
<< m2 >>
rect 93 235 94 236 
<< m2c >>
rect 93 235 94 236 
<< m1 >>
rect 93 235 94 236 
<< m2 >>
rect 93 235 94 236 
<< m1 >>
rect 94 235 95 236 
<< m1 >>
rect 95 235 96 236 
<< m1 >>
rect 142 235 143 236 
<< m1 >>
rect 143 235 144 236 
<< m1 >>
rect 144 235 145 236 
<< m1 >>
rect 145 235 146 236 
<< m1 >>
rect 146 235 147 236 
<< m1 >>
rect 147 235 148 236 
<< m1 >>
rect 148 235 149 236 
<< m1 >>
rect 149 235 150 236 
<< m1 >>
rect 150 235 151 236 
<< m2 >>
rect 15 236 16 237 
<< m1 >>
rect 16 236 17 237 
<< m1 >>
rect 17 236 18 237 
<< m1 >>
rect 18 236 19 237 
<< m1 >>
rect 19 236 20 237 
<< m1 >>
rect 20 236 21 237 
<< m2 >>
rect 20 236 21 237 
<< m1 >>
rect 21 236 22 237 
<< m1 >>
rect 22 236 23 237 
<< m1 >>
rect 23 236 24 237 
<< m1 >>
rect 24 236 25 237 
<< m2 >>
rect 24 236 25 237 
<< m1 >>
rect 25 236 26 237 
<< m1 >>
rect 26 236 27 237 
<< m1 >>
rect 27 236 28 237 
<< m1 >>
rect 28 236 29 237 
<< m2 >>
rect 28 236 29 237 
<< m1 >>
rect 34 236 35 237 
<< m1 >>
rect 35 236 36 237 
<< m1 >>
rect 36 236 37 237 
<< m1 >>
rect 37 236 38 237 
<< m1 >>
rect 38 236 39 237 
<< m1 >>
rect 39 236 40 237 
<< m1 >>
rect 40 236 41 237 
<< m1 >>
rect 41 236 42 237 
<< m1 >>
rect 42 236 43 237 
<< m1 >>
rect 43 236 44 237 
<< m1 >>
rect 44 236 45 237 
<< m1 >>
rect 45 236 46 237 
<< m1 >>
rect 46 236 47 237 
<< m1 >>
rect 71 236 72 237 
<< m1 >>
rect 73 236 74 237 
<< m1 >>
rect 91 236 92 237 
<< m2 >>
rect 15 237 16 238 
<< m1 >>
rect 16 237 17 238 
<< m2 >>
rect 20 237 21 238 
<< m2 >>
rect 24 237 25 238 
<< m2 >>
rect 28 237 29 238 
<< m2 >>
rect 29 237 30 238 
<< m1 >>
rect 30 237 31 238 
<< m2 >>
rect 30 237 31 238 
<< m2c >>
rect 30 237 31 238 
<< m1 >>
rect 30 237 31 238 
<< m2 >>
rect 30 237 31 238 
<< m1 >>
rect 34 237 35 238 
<< m1 >>
rect 71 237 72 238 
<< m1 >>
rect 73 237 74 238 
<< m1 >>
rect 91 237 92 238 
<< m2 >>
rect 15 238 16 239 
<< m1 >>
rect 16 238 17 239 
<< m2 >>
rect 16 238 17 239 
<< m2 >>
rect 17 238 18 239 
<< m1 >>
rect 18 238 19 239 
<< m2 >>
rect 18 238 19 239 
<< m2c >>
rect 18 238 19 239 
<< m1 >>
rect 18 238 19 239 
<< m2 >>
rect 18 238 19 239 
<< m2 >>
rect 20 238 21 239 
<< m2 >>
rect 24 238 25 239 
<< m1 >>
rect 30 238 31 239 
<< m1 >>
rect 34 238 35 239 
<< m2 >>
rect 46 238 47 239 
<< m2 >>
rect 47 238 48 239 
<< m2 >>
rect 48 238 49 239 
<< m2 >>
rect 49 238 50 239 
<< m2 >>
rect 50 238 51 239 
<< m2 >>
rect 51 238 52 239 
<< m2 >>
rect 52 238 53 239 
<< m2 >>
rect 53 238 54 239 
<< m2 >>
rect 54 238 55 239 
<< m2 >>
rect 55 238 56 239 
<< m2 >>
rect 56 238 57 239 
<< m1 >>
rect 57 238 58 239 
<< m2 >>
rect 57 238 58 239 
<< m2c >>
rect 57 238 58 239 
<< m1 >>
rect 57 238 58 239 
<< m2 >>
rect 57 238 58 239 
<< m1 >>
rect 58 238 59 239 
<< m1 >>
rect 59 238 60 239 
<< m1 >>
rect 60 238 61 239 
<< m1 >>
rect 61 238 62 239 
<< m1 >>
rect 62 238 63 239 
<< m1 >>
rect 63 238 64 239 
<< m1 >>
rect 64 238 65 239 
<< m1 >>
rect 65 238 66 239 
<< m1 >>
rect 66 238 67 239 
<< m1 >>
rect 67 238 68 239 
<< m1 >>
rect 68 238 69 239 
<< m1 >>
rect 69 238 70 239 
<< m1 >>
rect 70 238 71 239 
<< m1 >>
rect 71 238 72 239 
<< m1 >>
rect 73 238 74 239 
<< m1 >>
rect 91 238 92 239 
<< m1 >>
rect 16 239 17 240 
<< m1 >>
rect 18 239 19 240 
<< m1 >>
rect 19 239 20 240 
<< m1 >>
rect 20 239 21 240 
<< m2 >>
rect 20 239 21 240 
<< m1 >>
rect 21 239 22 240 
<< m1 >>
rect 22 239 23 240 
<< m1 >>
rect 23 239 24 240 
<< m1 >>
rect 24 239 25 240 
<< m2 >>
rect 24 239 25 240 
<< m1 >>
rect 25 239 26 240 
<< m1 >>
rect 26 239 27 240 
<< m1 >>
rect 27 239 28 240 
<< m1 >>
rect 28 239 29 240 
<< m2 >>
rect 28 239 29 240 
<< m2c >>
rect 28 239 29 240 
<< m1 >>
rect 28 239 29 240 
<< m2 >>
rect 28 239 29 240 
<< m2 >>
rect 29 239 30 240 
<< m1 >>
rect 30 239 31 240 
<< m2 >>
rect 30 239 31 240 
<< m2 >>
rect 31 239 32 240 
<< m1 >>
rect 32 239 33 240 
<< m2 >>
rect 32 239 33 240 
<< m2c >>
rect 32 239 33 240 
<< m1 >>
rect 32 239 33 240 
<< m2 >>
rect 32 239 33 240 
<< m2 >>
rect 33 239 34 240 
<< m1 >>
rect 34 239 35 240 
<< m2 >>
rect 34 239 35 240 
<< m2 >>
rect 35 239 36 240 
<< m1 >>
rect 36 239 37 240 
<< m2 >>
rect 36 239 37 240 
<< m2c >>
rect 36 239 37 240 
<< m1 >>
rect 36 239 37 240 
<< m2 >>
rect 36 239 37 240 
<< m1 >>
rect 37 239 38 240 
<< m1 >>
rect 38 239 39 240 
<< m1 >>
rect 39 239 40 240 
<< m1 >>
rect 40 239 41 240 
<< m1 >>
rect 41 239 42 240 
<< m1 >>
rect 42 239 43 240 
<< m1 >>
rect 43 239 44 240 
<< m1 >>
rect 44 239 45 240 
<< m1 >>
rect 45 239 46 240 
<< m1 >>
rect 46 239 47 240 
<< m2 >>
rect 46 239 47 240 
<< m1 >>
rect 47 239 48 240 
<< m1 >>
rect 48 239 49 240 
<< m1 >>
rect 49 239 50 240 
<< m1 >>
rect 50 239 51 240 
<< m1 >>
rect 51 239 52 240 
<< m1 >>
rect 52 239 53 240 
<< m1 >>
rect 53 239 54 240 
<< m1 >>
rect 54 239 55 240 
<< m1 >>
rect 55 239 56 240 
<< m1 >>
rect 73 239 74 240 
<< m1 >>
rect 91 239 92 240 
<< m1 >>
rect 16 240 17 241 
<< m2 >>
rect 20 240 21 241 
<< m2 >>
rect 24 240 25 241 
<< m1 >>
rect 30 240 31 241 
<< m1 >>
rect 34 240 35 241 
<< m2 >>
rect 46 240 47 241 
<< m1 >>
rect 55 240 56 241 
<< m1 >>
rect 73 240 74 241 
<< m1 >>
rect 91 240 92 241 
<< m1 >>
rect 16 241 17 242 
<< m1 >>
rect 20 241 21 242 
<< m2 >>
rect 20 241 21 242 
<< m2c >>
rect 20 241 21 242 
<< m1 >>
rect 20 241 21 242 
<< m2 >>
rect 20 241 21 242 
<< m1 >>
rect 21 241 22 242 
<< m1 >>
rect 22 241 23 242 
<< m1 >>
rect 23 241 24 242 
<< m1 >>
rect 24 241 25 242 
<< m2 >>
rect 24 241 25 242 
<< m1 >>
rect 25 241 26 242 
<< m1 >>
rect 26 241 27 242 
<< m1 >>
rect 27 241 28 242 
<< m1 >>
rect 28 241 29 242 
<< m2 >>
rect 28 241 29 242 
<< m2c >>
rect 28 241 29 242 
<< m1 >>
rect 28 241 29 242 
<< m2 >>
rect 28 241 29 242 
<< m2 >>
rect 29 241 30 242 
<< m1 >>
rect 30 241 31 242 
<< m2 >>
rect 30 241 31 242 
<< m1 >>
rect 31 241 32 242 
<< m2 >>
rect 31 241 32 242 
<< m1 >>
rect 32 241 33 242 
<< m2 >>
rect 32 241 33 242 
<< m2 >>
rect 33 241 34 242 
<< m1 >>
rect 34 241 35 242 
<< m2 >>
rect 34 241 35 242 
<< m2 >>
rect 35 241 36 242 
<< m1 >>
rect 36 241 37 242 
<< m2 >>
rect 36 241 37 242 
<< m2c >>
rect 36 241 37 242 
<< m1 >>
rect 36 241 37 242 
<< m2 >>
rect 36 241 37 242 
<< m1 >>
rect 37 241 38 242 
<< m1 >>
rect 38 241 39 242 
<< m1 >>
rect 39 241 40 242 
<< m1 >>
rect 40 241 41 242 
<< m1 >>
rect 41 241 42 242 
<< m1 >>
rect 42 241 43 242 
<< m1 >>
rect 43 241 44 242 
<< m1 >>
rect 44 241 45 242 
<< m1 >>
rect 45 241 46 242 
<< m1 >>
rect 46 241 47 242 
<< m2 >>
rect 46 241 47 242 
<< m1 >>
rect 47 241 48 242 
<< m1 >>
rect 48 241 49 242 
<< m1 >>
rect 49 241 50 242 
<< m1 >>
rect 50 241 51 242 
<< m1 >>
rect 51 241 52 242 
<< m1 >>
rect 52 241 53 242 
<< m1 >>
rect 55 241 56 242 
<< m1 >>
rect 73 241 74 242 
<< m1 >>
rect 91 241 92 242 
<< m1 >>
rect 16 242 17 243 
<< m2 >>
rect 24 242 25 243 
<< m2 >>
rect 25 242 26 243 
<< m2 >>
rect 26 242 27 243 
<< m1 >>
rect 32 242 33 243 
<< m1 >>
rect 34 242 35 243 
<< m2 >>
rect 46 242 47 243 
<< m1 >>
rect 52 242 53 243 
<< m1 >>
rect 55 242 56 243 
<< m1 >>
rect 73 242 74 243 
<< m1 >>
rect 91 242 92 243 
<< m1 >>
rect 16 243 17 244 
<< m1 >>
rect 26 243 27 244 
<< m2 >>
rect 26 243 27 244 
<< m2c >>
rect 26 243 27 244 
<< m1 >>
rect 26 243 27 244 
<< m2 >>
rect 26 243 27 244 
<< m1 >>
rect 32 243 33 244 
<< m2 >>
rect 32 243 33 244 
<< m2c >>
rect 32 243 33 244 
<< m1 >>
rect 32 243 33 244 
<< m2 >>
rect 32 243 33 244 
<< m2 >>
rect 33 243 34 244 
<< m1 >>
rect 34 243 35 244 
<< m2 >>
rect 34 243 35 244 
<< m2 >>
rect 35 243 36 244 
<< m2 >>
rect 46 243 47 244 
<< m1 >>
rect 52 243 53 244 
<< m1 >>
rect 55 243 56 244 
<< m1 >>
rect 73 243 74 244 
<< m1 >>
rect 91 243 92 244 
<< m1 >>
rect 139 243 140 244 
<< m1 >>
rect 140 243 141 244 
<< m1 >>
rect 141 243 142 244 
<< m1 >>
rect 142 243 143 244 
<< m1 >>
rect 143 243 144 244 
<< m1 >>
rect 144 243 145 244 
<< m1 >>
rect 145 243 146 244 
<< m1 >>
rect 146 243 147 244 
<< m1 >>
rect 147 243 148 244 
<< m1 >>
rect 148 243 149 244 
<< m1 >>
rect 149 243 150 244 
<< m1 >>
rect 150 243 151 244 
<< m1 >>
rect 151 243 152 244 
<< m1 >>
rect 152 243 153 244 
<< m1 >>
rect 153 243 154 244 
<< m1 >>
rect 154 243 155 244 
<< m1 >>
rect 16 244 17 245 
<< m1 >>
rect 26 244 27 245 
<< m1 >>
rect 34 244 35 245 
<< m2 >>
rect 35 244 36 245 
<< m1 >>
rect 36 244 37 245 
<< m2 >>
rect 36 244 37 245 
<< m2c >>
rect 36 244 37 245 
<< m1 >>
rect 36 244 37 245 
<< m2 >>
rect 36 244 37 245 
<< m1 >>
rect 37 244 38 245 
<< m1 >>
rect 38 244 39 245 
<< m1 >>
rect 39 244 40 245 
<< m1 >>
rect 40 244 41 245 
<< m1 >>
rect 41 244 42 245 
<< m1 >>
rect 42 244 43 245 
<< m1 >>
rect 43 244 44 245 
<< m1 >>
rect 44 244 45 245 
<< m1 >>
rect 45 244 46 245 
<< m1 >>
rect 46 244 47 245 
<< m2 >>
rect 46 244 47 245 
<< m1 >>
rect 52 244 53 245 
<< m1 >>
rect 55 244 56 245 
<< m1 >>
rect 73 244 74 245 
<< m1 >>
rect 91 244 92 245 
<< m1 >>
rect 139 244 140 245 
<< m1 >>
rect 154 244 155 245 
<< m1 >>
rect 16 245 17 246 
<< m1 >>
rect 26 245 27 246 
<< m1 >>
rect 34 245 35 246 
<< m1 >>
rect 46 245 47 246 
<< m2 >>
rect 46 245 47 246 
<< m1 >>
rect 52 245 53 246 
<< m1 >>
rect 55 245 56 246 
<< m1 >>
rect 73 245 74 246 
<< m1 >>
rect 91 245 92 246 
<< m1 >>
rect 139 245 140 246 
<< m1 >>
rect 154 245 155 246 
<< pdiffusion >>
rect 12 246 13 247 
<< pdiffusion >>
rect 13 246 14 247 
<< pdiffusion >>
rect 14 246 15 247 
<< pdiffusion >>
rect 15 246 16 247 
<< m1 >>
rect 16 246 17 247 
<< pdiffusion >>
rect 16 246 17 247 
<< pdiffusion >>
rect 17 246 18 247 
<< m1 >>
rect 26 246 27 247 
<< pdiffusion >>
rect 30 246 31 247 
<< pdiffusion >>
rect 31 246 32 247 
<< pdiffusion >>
rect 32 246 33 247 
<< pdiffusion >>
rect 33 246 34 247 
<< m1 >>
rect 34 246 35 247 
<< pdiffusion >>
rect 34 246 35 247 
<< pdiffusion >>
rect 35 246 36 247 
<< m1 >>
rect 44 246 45 247 
<< m2 >>
rect 44 246 45 247 
<< m2c >>
rect 44 246 45 247 
<< m1 >>
rect 44 246 45 247 
<< m2 >>
rect 44 246 45 247 
<< m2 >>
rect 45 246 46 247 
<< m1 >>
rect 46 246 47 247 
<< m2 >>
rect 46 246 47 247 
<< pdiffusion >>
rect 48 246 49 247 
<< pdiffusion >>
rect 49 246 50 247 
<< pdiffusion >>
rect 50 246 51 247 
<< pdiffusion >>
rect 51 246 52 247 
<< m1 >>
rect 52 246 53 247 
<< pdiffusion >>
rect 52 246 53 247 
<< pdiffusion >>
rect 53 246 54 247 
<< m1 >>
rect 55 246 56 247 
<< pdiffusion >>
rect 66 246 67 247 
<< pdiffusion >>
rect 67 246 68 247 
<< pdiffusion >>
rect 68 246 69 247 
<< pdiffusion >>
rect 69 246 70 247 
<< pdiffusion >>
rect 70 246 71 247 
<< pdiffusion >>
rect 71 246 72 247 
<< m1 >>
rect 73 246 74 247 
<< pdiffusion >>
rect 84 246 85 247 
<< pdiffusion >>
rect 85 246 86 247 
<< pdiffusion >>
rect 86 246 87 247 
<< pdiffusion >>
rect 87 246 88 247 
<< pdiffusion >>
rect 88 246 89 247 
<< pdiffusion >>
rect 89 246 90 247 
<< m1 >>
rect 91 246 92 247 
<< pdiffusion >>
rect 102 246 103 247 
<< pdiffusion >>
rect 103 246 104 247 
<< pdiffusion >>
rect 104 246 105 247 
<< pdiffusion >>
rect 105 246 106 247 
<< pdiffusion >>
rect 106 246 107 247 
<< pdiffusion >>
rect 107 246 108 247 
<< pdiffusion >>
rect 120 246 121 247 
<< pdiffusion >>
rect 121 246 122 247 
<< pdiffusion >>
rect 122 246 123 247 
<< pdiffusion >>
rect 123 246 124 247 
<< pdiffusion >>
rect 124 246 125 247 
<< pdiffusion >>
rect 125 246 126 247 
<< pdiffusion >>
rect 138 246 139 247 
<< m1 >>
rect 139 246 140 247 
<< pdiffusion >>
rect 139 246 140 247 
<< pdiffusion >>
rect 140 246 141 247 
<< pdiffusion >>
rect 141 246 142 247 
<< pdiffusion >>
rect 142 246 143 247 
<< pdiffusion >>
rect 143 246 144 247 
<< m1 >>
rect 154 246 155 247 
<< pdiffusion >>
rect 156 246 157 247 
<< pdiffusion >>
rect 157 246 158 247 
<< pdiffusion >>
rect 158 246 159 247 
<< pdiffusion >>
rect 159 246 160 247 
<< pdiffusion >>
rect 160 246 161 247 
<< pdiffusion >>
rect 161 246 162 247 
<< pdiffusion >>
rect 12 247 13 248 
<< pdiffusion >>
rect 13 247 14 248 
<< pdiffusion >>
rect 14 247 15 248 
<< pdiffusion >>
rect 15 247 16 248 
<< pdiffusion >>
rect 16 247 17 248 
<< pdiffusion >>
rect 17 247 18 248 
<< m1 >>
rect 26 247 27 248 
<< pdiffusion >>
rect 30 247 31 248 
<< pdiffusion >>
rect 31 247 32 248 
<< pdiffusion >>
rect 32 247 33 248 
<< pdiffusion >>
rect 33 247 34 248 
<< pdiffusion >>
rect 34 247 35 248 
<< pdiffusion >>
rect 35 247 36 248 
<< m1 >>
rect 44 247 45 248 
<< m1 >>
rect 46 247 47 248 
<< pdiffusion >>
rect 48 247 49 248 
<< pdiffusion >>
rect 49 247 50 248 
<< pdiffusion >>
rect 50 247 51 248 
<< pdiffusion >>
rect 51 247 52 248 
<< pdiffusion >>
rect 52 247 53 248 
<< pdiffusion >>
rect 53 247 54 248 
<< m1 >>
rect 55 247 56 248 
<< pdiffusion >>
rect 66 247 67 248 
<< pdiffusion >>
rect 67 247 68 248 
<< pdiffusion >>
rect 68 247 69 248 
<< pdiffusion >>
rect 69 247 70 248 
<< pdiffusion >>
rect 70 247 71 248 
<< pdiffusion >>
rect 71 247 72 248 
<< m1 >>
rect 73 247 74 248 
<< pdiffusion >>
rect 84 247 85 248 
<< pdiffusion >>
rect 85 247 86 248 
<< pdiffusion >>
rect 86 247 87 248 
<< pdiffusion >>
rect 87 247 88 248 
<< pdiffusion >>
rect 88 247 89 248 
<< pdiffusion >>
rect 89 247 90 248 
<< m1 >>
rect 91 247 92 248 
<< pdiffusion >>
rect 102 247 103 248 
<< pdiffusion >>
rect 103 247 104 248 
<< pdiffusion >>
rect 104 247 105 248 
<< pdiffusion >>
rect 105 247 106 248 
<< pdiffusion >>
rect 106 247 107 248 
<< pdiffusion >>
rect 107 247 108 248 
<< pdiffusion >>
rect 120 247 121 248 
<< pdiffusion >>
rect 121 247 122 248 
<< pdiffusion >>
rect 122 247 123 248 
<< pdiffusion >>
rect 123 247 124 248 
<< pdiffusion >>
rect 124 247 125 248 
<< pdiffusion >>
rect 125 247 126 248 
<< pdiffusion >>
rect 138 247 139 248 
<< pdiffusion >>
rect 139 247 140 248 
<< pdiffusion >>
rect 140 247 141 248 
<< pdiffusion >>
rect 141 247 142 248 
<< pdiffusion >>
rect 142 247 143 248 
<< pdiffusion >>
rect 143 247 144 248 
<< m1 >>
rect 154 247 155 248 
<< pdiffusion >>
rect 156 247 157 248 
<< pdiffusion >>
rect 157 247 158 248 
<< pdiffusion >>
rect 158 247 159 248 
<< pdiffusion >>
rect 159 247 160 248 
<< pdiffusion >>
rect 160 247 161 248 
<< pdiffusion >>
rect 161 247 162 248 
<< pdiffusion >>
rect 12 248 13 249 
<< pdiffusion >>
rect 13 248 14 249 
<< pdiffusion >>
rect 14 248 15 249 
<< pdiffusion >>
rect 15 248 16 249 
<< pdiffusion >>
rect 16 248 17 249 
<< pdiffusion >>
rect 17 248 18 249 
<< m1 >>
rect 26 248 27 249 
<< pdiffusion >>
rect 30 248 31 249 
<< pdiffusion >>
rect 31 248 32 249 
<< pdiffusion >>
rect 32 248 33 249 
<< pdiffusion >>
rect 33 248 34 249 
<< pdiffusion >>
rect 34 248 35 249 
<< pdiffusion >>
rect 35 248 36 249 
<< m1 >>
rect 44 248 45 249 
<< m1 >>
rect 46 248 47 249 
<< pdiffusion >>
rect 48 248 49 249 
<< pdiffusion >>
rect 49 248 50 249 
<< pdiffusion >>
rect 50 248 51 249 
<< pdiffusion >>
rect 51 248 52 249 
<< pdiffusion >>
rect 52 248 53 249 
<< pdiffusion >>
rect 53 248 54 249 
<< m1 >>
rect 55 248 56 249 
<< pdiffusion >>
rect 66 248 67 249 
<< pdiffusion >>
rect 67 248 68 249 
<< pdiffusion >>
rect 68 248 69 249 
<< pdiffusion >>
rect 69 248 70 249 
<< pdiffusion >>
rect 70 248 71 249 
<< pdiffusion >>
rect 71 248 72 249 
<< m1 >>
rect 73 248 74 249 
<< pdiffusion >>
rect 84 248 85 249 
<< pdiffusion >>
rect 85 248 86 249 
<< pdiffusion >>
rect 86 248 87 249 
<< pdiffusion >>
rect 87 248 88 249 
<< pdiffusion >>
rect 88 248 89 249 
<< pdiffusion >>
rect 89 248 90 249 
<< m1 >>
rect 91 248 92 249 
<< pdiffusion >>
rect 102 248 103 249 
<< pdiffusion >>
rect 103 248 104 249 
<< pdiffusion >>
rect 104 248 105 249 
<< pdiffusion >>
rect 105 248 106 249 
<< pdiffusion >>
rect 106 248 107 249 
<< pdiffusion >>
rect 107 248 108 249 
<< pdiffusion >>
rect 120 248 121 249 
<< pdiffusion >>
rect 121 248 122 249 
<< pdiffusion >>
rect 122 248 123 249 
<< pdiffusion >>
rect 123 248 124 249 
<< pdiffusion >>
rect 124 248 125 249 
<< pdiffusion >>
rect 125 248 126 249 
<< pdiffusion >>
rect 138 248 139 249 
<< pdiffusion >>
rect 139 248 140 249 
<< pdiffusion >>
rect 140 248 141 249 
<< pdiffusion >>
rect 141 248 142 249 
<< pdiffusion >>
rect 142 248 143 249 
<< pdiffusion >>
rect 143 248 144 249 
<< m1 >>
rect 154 248 155 249 
<< pdiffusion >>
rect 156 248 157 249 
<< pdiffusion >>
rect 157 248 158 249 
<< pdiffusion >>
rect 158 248 159 249 
<< pdiffusion >>
rect 159 248 160 249 
<< pdiffusion >>
rect 160 248 161 249 
<< pdiffusion >>
rect 161 248 162 249 
<< pdiffusion >>
rect 12 249 13 250 
<< pdiffusion >>
rect 13 249 14 250 
<< pdiffusion >>
rect 14 249 15 250 
<< pdiffusion >>
rect 15 249 16 250 
<< pdiffusion >>
rect 16 249 17 250 
<< pdiffusion >>
rect 17 249 18 250 
<< m1 >>
rect 26 249 27 250 
<< pdiffusion >>
rect 30 249 31 250 
<< pdiffusion >>
rect 31 249 32 250 
<< pdiffusion >>
rect 32 249 33 250 
<< pdiffusion >>
rect 33 249 34 250 
<< pdiffusion >>
rect 34 249 35 250 
<< pdiffusion >>
rect 35 249 36 250 
<< m1 >>
rect 44 249 45 250 
<< m1 >>
rect 46 249 47 250 
<< pdiffusion >>
rect 48 249 49 250 
<< pdiffusion >>
rect 49 249 50 250 
<< pdiffusion >>
rect 50 249 51 250 
<< pdiffusion >>
rect 51 249 52 250 
<< pdiffusion >>
rect 52 249 53 250 
<< pdiffusion >>
rect 53 249 54 250 
<< m1 >>
rect 55 249 56 250 
<< pdiffusion >>
rect 66 249 67 250 
<< pdiffusion >>
rect 67 249 68 250 
<< pdiffusion >>
rect 68 249 69 250 
<< pdiffusion >>
rect 69 249 70 250 
<< pdiffusion >>
rect 70 249 71 250 
<< pdiffusion >>
rect 71 249 72 250 
<< m1 >>
rect 73 249 74 250 
<< pdiffusion >>
rect 84 249 85 250 
<< pdiffusion >>
rect 85 249 86 250 
<< pdiffusion >>
rect 86 249 87 250 
<< pdiffusion >>
rect 87 249 88 250 
<< pdiffusion >>
rect 88 249 89 250 
<< pdiffusion >>
rect 89 249 90 250 
<< m1 >>
rect 91 249 92 250 
<< pdiffusion >>
rect 102 249 103 250 
<< pdiffusion >>
rect 103 249 104 250 
<< pdiffusion >>
rect 104 249 105 250 
<< pdiffusion >>
rect 105 249 106 250 
<< pdiffusion >>
rect 106 249 107 250 
<< pdiffusion >>
rect 107 249 108 250 
<< pdiffusion >>
rect 120 249 121 250 
<< pdiffusion >>
rect 121 249 122 250 
<< pdiffusion >>
rect 122 249 123 250 
<< pdiffusion >>
rect 123 249 124 250 
<< pdiffusion >>
rect 124 249 125 250 
<< pdiffusion >>
rect 125 249 126 250 
<< pdiffusion >>
rect 138 249 139 250 
<< pdiffusion >>
rect 139 249 140 250 
<< pdiffusion >>
rect 140 249 141 250 
<< pdiffusion >>
rect 141 249 142 250 
<< pdiffusion >>
rect 142 249 143 250 
<< pdiffusion >>
rect 143 249 144 250 
<< m1 >>
rect 154 249 155 250 
<< pdiffusion >>
rect 156 249 157 250 
<< pdiffusion >>
rect 157 249 158 250 
<< pdiffusion >>
rect 158 249 159 250 
<< pdiffusion >>
rect 159 249 160 250 
<< pdiffusion >>
rect 160 249 161 250 
<< pdiffusion >>
rect 161 249 162 250 
<< pdiffusion >>
rect 12 250 13 251 
<< pdiffusion >>
rect 13 250 14 251 
<< pdiffusion >>
rect 14 250 15 251 
<< pdiffusion >>
rect 15 250 16 251 
<< pdiffusion >>
rect 16 250 17 251 
<< pdiffusion >>
rect 17 250 18 251 
<< m1 >>
rect 26 250 27 251 
<< pdiffusion >>
rect 30 250 31 251 
<< pdiffusion >>
rect 31 250 32 251 
<< pdiffusion >>
rect 32 250 33 251 
<< pdiffusion >>
rect 33 250 34 251 
<< pdiffusion >>
rect 34 250 35 251 
<< pdiffusion >>
rect 35 250 36 251 
<< m1 >>
rect 44 250 45 251 
<< m1 >>
rect 46 250 47 251 
<< pdiffusion >>
rect 48 250 49 251 
<< pdiffusion >>
rect 49 250 50 251 
<< pdiffusion >>
rect 50 250 51 251 
<< pdiffusion >>
rect 51 250 52 251 
<< pdiffusion >>
rect 52 250 53 251 
<< pdiffusion >>
rect 53 250 54 251 
<< m1 >>
rect 55 250 56 251 
<< pdiffusion >>
rect 66 250 67 251 
<< pdiffusion >>
rect 67 250 68 251 
<< pdiffusion >>
rect 68 250 69 251 
<< pdiffusion >>
rect 69 250 70 251 
<< pdiffusion >>
rect 70 250 71 251 
<< pdiffusion >>
rect 71 250 72 251 
<< m1 >>
rect 73 250 74 251 
<< pdiffusion >>
rect 84 250 85 251 
<< pdiffusion >>
rect 85 250 86 251 
<< pdiffusion >>
rect 86 250 87 251 
<< pdiffusion >>
rect 87 250 88 251 
<< pdiffusion >>
rect 88 250 89 251 
<< pdiffusion >>
rect 89 250 90 251 
<< m1 >>
rect 91 250 92 251 
<< pdiffusion >>
rect 102 250 103 251 
<< pdiffusion >>
rect 103 250 104 251 
<< pdiffusion >>
rect 104 250 105 251 
<< pdiffusion >>
rect 105 250 106 251 
<< pdiffusion >>
rect 106 250 107 251 
<< pdiffusion >>
rect 107 250 108 251 
<< pdiffusion >>
rect 120 250 121 251 
<< pdiffusion >>
rect 121 250 122 251 
<< pdiffusion >>
rect 122 250 123 251 
<< pdiffusion >>
rect 123 250 124 251 
<< pdiffusion >>
rect 124 250 125 251 
<< pdiffusion >>
rect 125 250 126 251 
<< pdiffusion >>
rect 138 250 139 251 
<< pdiffusion >>
rect 139 250 140 251 
<< pdiffusion >>
rect 140 250 141 251 
<< pdiffusion >>
rect 141 250 142 251 
<< pdiffusion >>
rect 142 250 143 251 
<< pdiffusion >>
rect 143 250 144 251 
<< m1 >>
rect 154 250 155 251 
<< pdiffusion >>
rect 156 250 157 251 
<< pdiffusion >>
rect 157 250 158 251 
<< pdiffusion >>
rect 158 250 159 251 
<< pdiffusion >>
rect 159 250 160 251 
<< pdiffusion >>
rect 160 250 161 251 
<< pdiffusion >>
rect 161 250 162 251 
<< pdiffusion >>
rect 12 251 13 252 
<< pdiffusion >>
rect 13 251 14 252 
<< pdiffusion >>
rect 14 251 15 252 
<< pdiffusion >>
rect 15 251 16 252 
<< pdiffusion >>
rect 16 251 17 252 
<< pdiffusion >>
rect 17 251 18 252 
<< m1 >>
rect 26 251 27 252 
<< pdiffusion >>
rect 30 251 31 252 
<< pdiffusion >>
rect 31 251 32 252 
<< pdiffusion >>
rect 32 251 33 252 
<< pdiffusion >>
rect 33 251 34 252 
<< pdiffusion >>
rect 34 251 35 252 
<< pdiffusion >>
rect 35 251 36 252 
<< m1 >>
rect 44 251 45 252 
<< m1 >>
rect 46 251 47 252 
<< pdiffusion >>
rect 48 251 49 252 
<< pdiffusion >>
rect 49 251 50 252 
<< pdiffusion >>
rect 50 251 51 252 
<< pdiffusion >>
rect 51 251 52 252 
<< m1 >>
rect 52 251 53 252 
<< pdiffusion >>
rect 52 251 53 252 
<< pdiffusion >>
rect 53 251 54 252 
<< m1 >>
rect 55 251 56 252 
<< pdiffusion >>
rect 66 251 67 252 
<< m1 >>
rect 67 251 68 252 
<< pdiffusion >>
rect 67 251 68 252 
<< pdiffusion >>
rect 68 251 69 252 
<< pdiffusion >>
rect 69 251 70 252 
<< pdiffusion >>
rect 70 251 71 252 
<< pdiffusion >>
rect 71 251 72 252 
<< m1 >>
rect 73 251 74 252 
<< pdiffusion >>
rect 84 251 85 252 
<< m1 >>
rect 85 251 86 252 
<< pdiffusion >>
rect 85 251 86 252 
<< pdiffusion >>
rect 86 251 87 252 
<< pdiffusion >>
rect 87 251 88 252 
<< pdiffusion >>
rect 88 251 89 252 
<< pdiffusion >>
rect 89 251 90 252 
<< m1 >>
rect 91 251 92 252 
<< pdiffusion >>
rect 102 251 103 252 
<< pdiffusion >>
rect 103 251 104 252 
<< pdiffusion >>
rect 104 251 105 252 
<< pdiffusion >>
rect 105 251 106 252 
<< pdiffusion >>
rect 106 251 107 252 
<< pdiffusion >>
rect 107 251 108 252 
<< pdiffusion >>
rect 120 251 121 252 
<< pdiffusion >>
rect 121 251 122 252 
<< pdiffusion >>
rect 122 251 123 252 
<< pdiffusion >>
rect 123 251 124 252 
<< m1 >>
rect 124 251 125 252 
<< pdiffusion >>
rect 124 251 125 252 
<< pdiffusion >>
rect 125 251 126 252 
<< pdiffusion >>
rect 138 251 139 252 
<< pdiffusion >>
rect 139 251 140 252 
<< pdiffusion >>
rect 140 251 141 252 
<< pdiffusion >>
rect 141 251 142 252 
<< pdiffusion >>
rect 142 251 143 252 
<< pdiffusion >>
rect 143 251 144 252 
<< m1 >>
rect 154 251 155 252 
<< pdiffusion >>
rect 156 251 157 252 
<< pdiffusion >>
rect 157 251 158 252 
<< pdiffusion >>
rect 158 251 159 252 
<< pdiffusion >>
rect 159 251 160 252 
<< m1 >>
rect 160 251 161 252 
<< pdiffusion >>
rect 160 251 161 252 
<< pdiffusion >>
rect 161 251 162 252 
<< m1 >>
rect 26 252 27 253 
<< m1 >>
rect 44 252 45 253 
<< m1 >>
rect 46 252 47 253 
<< m1 >>
rect 52 252 53 253 
<< m1 >>
rect 55 252 56 253 
<< m1 >>
rect 67 252 68 253 
<< m1 >>
rect 73 252 74 253 
<< m1 >>
rect 85 252 86 253 
<< m1 >>
rect 91 252 92 253 
<< m1 >>
rect 124 252 125 253 
<< m1 >>
rect 154 252 155 253 
<< m1 >>
rect 160 252 161 253 
<< m1 >>
rect 26 253 27 254 
<< m1 >>
rect 44 253 45 254 
<< m1 >>
rect 46 253 47 254 
<< m1 >>
rect 52 253 53 254 
<< m1 >>
rect 55 253 56 254 
<< m1 >>
rect 56 253 57 254 
<< m1 >>
rect 57 253 58 254 
<< m1 >>
rect 58 253 59 254 
<< m1 >>
rect 59 253 60 254 
<< m1 >>
rect 60 253 61 254 
<< m1 >>
rect 61 253 62 254 
<< m1 >>
rect 62 253 63 254 
<< m1 >>
rect 63 253 64 254 
<< m1 >>
rect 64 253 65 254 
<< m1 >>
rect 65 253 66 254 
<< m1 >>
rect 66 253 67 254 
<< m1 >>
rect 67 253 68 254 
<< m1 >>
rect 73 253 74 254 
<< m1 >>
rect 85 253 86 254 
<< m1 >>
rect 91 253 92 254 
<< m1 >>
rect 124 253 125 254 
<< m1 >>
rect 154 253 155 254 
<< m1 >>
rect 160 253 161 254 
<< m1 >>
rect 26 254 27 255 
<< m1 >>
rect 44 254 45 255 
<< m1 >>
rect 46 254 47 255 
<< m1 >>
rect 52 254 53 255 
<< m1 >>
rect 73 254 74 255 
<< m1 >>
rect 85 254 86 255 
<< m1 >>
rect 86 254 87 255 
<< m1 >>
rect 87 254 88 255 
<< m1 >>
rect 88 254 89 255 
<< m1 >>
rect 89 254 90 255 
<< m1 >>
rect 90 254 91 255 
<< m1 >>
rect 91 254 92 255 
<< m1 >>
rect 124 254 125 255 
<< m1 >>
rect 154 254 155 255 
<< m1 >>
rect 160 254 161 255 
<< m1 >>
rect 26 255 27 256 
<< m1 >>
rect 44 255 45 256 
<< m1 >>
rect 46 255 47 256 
<< m1 >>
rect 52 255 53 256 
<< m1 >>
rect 73 255 74 256 
<< m1 >>
rect 124 255 125 256 
<< m1 >>
rect 154 255 155 256 
<< m1 >>
rect 160 255 161 256 
<< m1 >>
rect 26 256 27 257 
<< m1 >>
rect 27 256 28 257 
<< m1 >>
rect 28 256 29 257 
<< m1 >>
rect 29 256 30 257 
<< m1 >>
rect 30 256 31 257 
<< m1 >>
rect 31 256 32 257 
<< m1 >>
rect 32 256 33 257 
<< m1 >>
rect 33 256 34 257 
<< m1 >>
rect 34 256 35 257 
<< m1 >>
rect 35 256 36 257 
<< m1 >>
rect 36 256 37 257 
<< m1 >>
rect 37 256 38 257 
<< m1 >>
rect 38 256 39 257 
<< m1 >>
rect 39 256 40 257 
<< m1 >>
rect 40 256 41 257 
<< m1 >>
rect 41 256 42 257 
<< m1 >>
rect 42 256 43 257 
<< m1 >>
rect 43 256 44 257 
<< m1 >>
rect 44 256 45 257 
<< m1 >>
rect 46 256 47 257 
<< m1 >>
rect 47 256 48 257 
<< m1 >>
rect 48 256 49 257 
<< m1 >>
rect 49 256 50 257 
<< m1 >>
rect 50 256 51 257 
<< m1 >>
rect 51 256 52 257 
<< m1 >>
rect 52 256 53 257 
<< m1 >>
rect 73 256 74 257 
<< m1 >>
rect 74 256 75 257 
<< m1 >>
rect 75 256 76 257 
<< m1 >>
rect 76 256 77 257 
<< m1 >>
rect 77 256 78 257 
<< m1 >>
rect 78 256 79 257 
<< m1 >>
rect 79 256 80 257 
<< m1 >>
rect 80 256 81 257 
<< m1 >>
rect 81 256 82 257 
<< m1 >>
rect 82 256 83 257 
<< m1 >>
rect 83 256 84 257 
<< m1 >>
rect 84 256 85 257 
<< m1 >>
rect 85 256 86 257 
<< m1 >>
rect 86 256 87 257 
<< m1 >>
rect 87 256 88 257 
<< m1 >>
rect 88 256 89 257 
<< m1 >>
rect 89 256 90 257 
<< m1 >>
rect 90 256 91 257 
<< m1 >>
rect 91 256 92 257 
<< m1 >>
rect 92 256 93 257 
<< m1 >>
rect 93 256 94 257 
<< m1 >>
rect 94 256 95 257 
<< m1 >>
rect 95 256 96 257 
<< m1 >>
rect 96 256 97 257 
<< m1 >>
rect 97 256 98 257 
<< m1 >>
rect 98 256 99 257 
<< m1 >>
rect 99 256 100 257 
<< m1 >>
rect 100 256 101 257 
<< m1 >>
rect 101 256 102 257 
<< m1 >>
rect 102 256 103 257 
<< m1 >>
rect 103 256 104 257 
<< m1 >>
rect 104 256 105 257 
<< m1 >>
rect 105 256 106 257 
<< m1 >>
rect 106 256 107 257 
<< m1 >>
rect 107 256 108 257 
<< m1 >>
rect 108 256 109 257 
<< m1 >>
rect 109 256 110 257 
<< m1 >>
rect 110 256 111 257 
<< m1 >>
rect 111 256 112 257 
<< m1 >>
rect 112 256 113 257 
<< m1 >>
rect 113 256 114 257 
<< m1 >>
rect 114 256 115 257 
<< m1 >>
rect 115 256 116 257 
<< m1 >>
rect 116 256 117 257 
<< m1 >>
rect 117 256 118 257 
<< m1 >>
rect 118 256 119 257 
<< m1 >>
rect 119 256 120 257 
<< m1 >>
rect 120 256 121 257 
<< m1 >>
rect 121 256 122 257 
<< m1 >>
rect 122 256 123 257 
<< m1 >>
rect 123 256 124 257 
<< m1 >>
rect 124 256 125 257 
<< m1 >>
rect 154 256 155 257 
<< m1 >>
rect 155 256 156 257 
<< m1 >>
rect 156 256 157 257 
<< m1 >>
rect 157 256 158 257 
<< m1 >>
rect 158 256 159 257 
<< m1 >>
rect 159 256 160 257 
<< m1 >>
rect 160 256 161 257 
<< labels >>
rlabel pdiffusion 157 66 158 67  0 t = 1
rlabel pdiffusion 160 66 161 67  0 t = 2
rlabel pdiffusion 157 71 158 72  0 t = 3
rlabel pdiffusion 160 71 161 72  0 t = 4
rlabel pdiffusion 156 66 162 72 0 cell no = 1
<< m1 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2c >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< labels >>
rlabel pdiffusion 103 174 104 175  0 t = 1
rlabel pdiffusion 106 174 107 175  0 t = 2
rlabel pdiffusion 103 179 104 180  0 t = 3
rlabel pdiffusion 106 179 107 180  0 t = 4
rlabel pdiffusion 102 174 108 180 0 cell no = 2
<< m1 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2c >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< labels >>
rlabel pdiffusion 211 66 212 67  0 t = 1
rlabel pdiffusion 214 66 215 67  0 t = 2
rlabel pdiffusion 211 71 212 72  0 t = 3
rlabel pdiffusion 214 71 215 72  0 t = 4
rlabel pdiffusion 210 66 216 72 0 cell no = 3
<< m1 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2c >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< labels >>
rlabel pdiffusion 193 138 194 139  0 t = 1
rlabel pdiffusion 196 138 197 139  0 t = 2
rlabel pdiffusion 193 143 194 144  0 t = 3
rlabel pdiffusion 196 143 197 144  0 t = 4
rlabel pdiffusion 192 138 198 144 0 cell no = 4
<< m1 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2c >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< labels >>
rlabel pdiffusion 85 12 86 13  0 t = 1
rlabel pdiffusion 88 12 89 13  0 t = 2
rlabel pdiffusion 85 17 86 18  0 t = 3
rlabel pdiffusion 88 17 89 18  0 t = 4
rlabel pdiffusion 84 12 90 18 0 cell no = 5
<< m1 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2c >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< labels >>
rlabel pdiffusion 193 174 194 175  0 t = 1
rlabel pdiffusion 196 174 197 175  0 t = 2
rlabel pdiffusion 193 179 194 180  0 t = 3
rlabel pdiffusion 196 179 197 180  0 t = 4
rlabel pdiffusion 192 174 198 180 0 cell no = 6
<< m1 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2c >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 7
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 8
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 67 174 68 175  0 t = 1
rlabel pdiffusion 70 174 71 175  0 t = 2
rlabel pdiffusion 67 179 68 180  0 t = 3
rlabel pdiffusion 70 179 71 180  0 t = 4
rlabel pdiffusion 66 174 72 180 0 cell no = 9
<< m1 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2c >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 10
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 193 30 194 31  0 t = 1
rlabel pdiffusion 196 30 197 31  0 t = 2
rlabel pdiffusion 193 35 194 36  0 t = 3
rlabel pdiffusion 196 35 197 36  0 t = 4
rlabel pdiffusion 192 30 198 36 0 cell no = 11
<< m1 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2c >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< labels >>
rlabel pdiffusion 211 102 212 103  0 t = 1
rlabel pdiffusion 214 102 215 103  0 t = 2
rlabel pdiffusion 211 107 212 108  0 t = 3
rlabel pdiffusion 214 107 215 108  0 t = 4
rlabel pdiffusion 210 102 216 108 0 cell no = 12
<< m1 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2c >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< labels >>
rlabel pdiffusion 229 48 230 49  0 t = 1
rlabel pdiffusion 232 48 233 49  0 t = 2
rlabel pdiffusion 229 53 230 54  0 t = 3
rlabel pdiffusion 232 53 233 54  0 t = 4
rlabel pdiffusion 228 48 234 54 0 cell no = 13
<< m1 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2c >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< labels >>
rlabel pdiffusion 247 30 248 31  0 t = 1
rlabel pdiffusion 250 30 251 31  0 t = 2
rlabel pdiffusion 247 35 248 36  0 t = 3
rlabel pdiffusion 250 35 251 36  0 t = 4
rlabel pdiffusion 246 30 252 36 0 cell no = 14
<< m1 >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< m2 >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< m2c >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< labels >>
rlabel pdiffusion 31 30 32 31  0 t = 1
rlabel pdiffusion 34 30 35 31  0 t = 2
rlabel pdiffusion 31 35 32 36  0 t = 3
rlabel pdiffusion 34 35 35 36  0 t = 4
rlabel pdiffusion 30 30 36 36 0 cell no = 15
<< m1 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2c >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< labels >>
rlabel pdiffusion 49 120 50 121  0 t = 1
rlabel pdiffusion 52 120 53 121  0 t = 2
rlabel pdiffusion 49 125 50 126  0 t = 3
rlabel pdiffusion 52 125 53 126  0 t = 4
rlabel pdiffusion 48 120 54 126 0 cell no = 16
<< m1 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2c >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< labels >>
rlabel pdiffusion 175 66 176 67  0 t = 1
rlabel pdiffusion 178 66 179 67  0 t = 2
rlabel pdiffusion 175 71 176 72  0 t = 3
rlabel pdiffusion 178 71 179 72  0 t = 4
rlabel pdiffusion 174 66 180 72 0 cell no = 17
<< m1 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2c >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< labels >>
rlabel pdiffusion 175 12 176 13  0 t = 1
rlabel pdiffusion 178 12 179 13  0 t = 2
rlabel pdiffusion 175 17 176 18  0 t = 3
rlabel pdiffusion 178 17 179 18  0 t = 4
rlabel pdiffusion 174 12 180 18 0 cell no = 18
<< m1 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2c >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< labels >>
rlabel pdiffusion 121 84 122 85  0 t = 1
rlabel pdiffusion 124 84 125 85  0 t = 2
rlabel pdiffusion 121 89 122 90  0 t = 3
rlabel pdiffusion 124 89 125 90  0 t = 4
rlabel pdiffusion 120 84 126 90 0 cell no = 19
<< m1 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2c >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< labels >>
rlabel pdiffusion 139 102 140 103  0 t = 1
rlabel pdiffusion 142 102 143 103  0 t = 2
rlabel pdiffusion 139 107 140 108  0 t = 3
rlabel pdiffusion 142 107 143 108  0 t = 4
rlabel pdiffusion 138 102 144 108 0 cell no = 20
<< m1 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2c >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< labels >>
rlabel pdiffusion 49 210 50 211  0 t = 1
rlabel pdiffusion 52 210 53 211  0 t = 2
rlabel pdiffusion 49 215 50 216  0 t = 3
rlabel pdiffusion 52 215 53 216  0 t = 4
rlabel pdiffusion 48 210 54 216 0 cell no = 21
<< m1 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2c >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< labels >>
rlabel pdiffusion 139 66 140 67  0 t = 1
rlabel pdiffusion 142 66 143 67  0 t = 2
rlabel pdiffusion 139 71 140 72  0 t = 3
rlabel pdiffusion 142 71 143 72  0 t = 4
rlabel pdiffusion 138 66 144 72 0 cell no = 22
<< m1 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2c >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< labels >>
rlabel pdiffusion 85 192 86 193  0 t = 1
rlabel pdiffusion 88 192 89 193  0 t = 2
rlabel pdiffusion 85 197 86 198  0 t = 3
rlabel pdiffusion 88 197 89 198  0 t = 4
rlabel pdiffusion 84 192 90 198 0 cell no = 23
<< m1 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2c >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< labels >>
rlabel pdiffusion 193 84 194 85  0 t = 1
rlabel pdiffusion 196 84 197 85  0 t = 2
rlabel pdiffusion 193 89 194 90  0 t = 3
rlabel pdiffusion 196 89 197 90  0 t = 4
rlabel pdiffusion 192 84 198 90 0 cell no = 24
<< m1 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2c >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< labels >>
rlabel pdiffusion 139 84 140 85  0 t = 1
rlabel pdiffusion 142 84 143 85  0 t = 2
rlabel pdiffusion 139 89 140 90  0 t = 3
rlabel pdiffusion 142 89 143 90  0 t = 4
rlabel pdiffusion 138 84 144 90 0 cell no = 25
<< m1 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2c >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< labels >>
rlabel pdiffusion 193 102 194 103  0 t = 1
rlabel pdiffusion 196 102 197 103  0 t = 2
rlabel pdiffusion 193 107 194 108  0 t = 3
rlabel pdiffusion 196 107 197 108  0 t = 4
rlabel pdiffusion 192 102 198 108 0 cell no = 26
<< m1 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2c >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< labels >>
rlabel pdiffusion 157 102 158 103  0 t = 1
rlabel pdiffusion 160 102 161 103  0 t = 2
rlabel pdiffusion 157 107 158 108  0 t = 3
rlabel pdiffusion 160 107 161 108  0 t = 4
rlabel pdiffusion 156 102 162 108 0 cell no = 27
<< m1 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2c >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< labels >>
rlabel pdiffusion 247 66 248 67  0 t = 1
rlabel pdiffusion 250 66 251 67  0 t = 2
rlabel pdiffusion 247 71 248 72  0 t = 3
rlabel pdiffusion 250 71 251 72  0 t = 4
rlabel pdiffusion 246 66 252 72 0 cell no = 28
<< m1 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2c >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< labels >>
rlabel pdiffusion 103 156 104 157  0 t = 1
rlabel pdiffusion 106 156 107 157  0 t = 2
rlabel pdiffusion 103 161 104 162  0 t = 3
rlabel pdiffusion 106 161 107 162  0 t = 4
rlabel pdiffusion 102 156 108 162 0 cell no = 29
<< m1 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2c >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 30
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 31
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 229 156 230 157  0 t = 1
rlabel pdiffusion 232 156 233 157  0 t = 2
rlabel pdiffusion 229 161 230 162  0 t = 3
rlabel pdiffusion 232 161 233 162  0 t = 4
rlabel pdiffusion 228 156 234 162 0 cell no = 32
<< m1 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2c >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 33
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 175 120 176 121  0 t = 1
rlabel pdiffusion 178 120 179 121  0 t = 2
rlabel pdiffusion 175 125 176 126  0 t = 3
rlabel pdiffusion 178 125 179 126  0 t = 4
rlabel pdiffusion 174 120 180 126 0 cell no = 34
<< m1 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2c >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< labels >>
rlabel pdiffusion 67 192 68 193  0 t = 1
rlabel pdiffusion 70 192 71 193  0 t = 2
rlabel pdiffusion 67 197 68 198  0 t = 3
rlabel pdiffusion 70 197 71 198  0 t = 4
rlabel pdiffusion 66 192 72 198 0 cell no = 35
<< m1 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2c >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 36
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< labels >>
rlabel pdiffusion 229 120 230 121  0 t = 1
rlabel pdiffusion 232 120 233 121  0 t = 2
rlabel pdiffusion 229 125 230 126  0 t = 3
rlabel pdiffusion 232 125 233 126  0 t = 4
rlabel pdiffusion 228 120 234 126 0 cell no = 37
<< m1 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2c >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< labels >>
rlabel pdiffusion 247 48 248 49  0 t = 1
rlabel pdiffusion 250 48 251 49  0 t = 2
rlabel pdiffusion 247 53 248 54  0 t = 3
rlabel pdiffusion 250 53 251 54  0 t = 4
rlabel pdiffusion 246 48 252 54 0 cell no = 38
<< m1 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2c >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< labels >>
rlabel pdiffusion 103 30 104 31  0 t = 1
rlabel pdiffusion 106 30 107 31  0 t = 2
rlabel pdiffusion 103 35 104 36  0 t = 3
rlabel pdiffusion 106 35 107 36  0 t = 4
rlabel pdiffusion 102 30 108 36 0 cell no = 39
<< m1 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2c >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< labels >>
rlabel pdiffusion 157 120 158 121  0 t = 1
rlabel pdiffusion 160 120 161 121  0 t = 2
rlabel pdiffusion 157 125 158 126  0 t = 3
rlabel pdiffusion 160 125 161 126  0 t = 4
rlabel pdiffusion 156 120 162 126 0 cell no = 40
<< m1 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2c >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< labels >>
rlabel pdiffusion 193 48 194 49  0 t = 1
rlabel pdiffusion 196 48 197 49  0 t = 2
rlabel pdiffusion 193 53 194 54  0 t = 3
rlabel pdiffusion 196 53 197 54  0 t = 4
rlabel pdiffusion 192 48 198 54 0 cell no = 41
<< m1 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2c >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< labels >>
rlabel pdiffusion 193 66 194 67  0 t = 1
rlabel pdiffusion 196 66 197 67  0 t = 2
rlabel pdiffusion 193 71 194 72  0 t = 3
rlabel pdiffusion 196 71 197 72  0 t = 4
rlabel pdiffusion 192 66 198 72 0 cell no = 42
<< m1 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2c >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< labels >>
rlabel pdiffusion 13 192 14 193  0 t = 1
rlabel pdiffusion 16 192 17 193  0 t = 2
rlabel pdiffusion 13 197 14 198  0 t = 3
rlabel pdiffusion 16 197 17 198  0 t = 4
rlabel pdiffusion 12 192 18 198 0 cell no = 43
<< m1 >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< m2 >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< m2c >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< labels >>
rlabel pdiffusion 139 174 140 175  0 t = 1
rlabel pdiffusion 142 174 143 175  0 t = 2
rlabel pdiffusion 139 179 140 180  0 t = 3
rlabel pdiffusion 142 179 143 180  0 t = 4
rlabel pdiffusion 138 174 144 180 0 cell no = 44
<< m1 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2c >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< labels >>
rlabel pdiffusion 139 192 140 193  0 t = 1
rlabel pdiffusion 142 192 143 193  0 t = 2
rlabel pdiffusion 139 197 140 198  0 t = 3
rlabel pdiffusion 142 197 143 198  0 t = 4
rlabel pdiffusion 138 192 144 198 0 cell no = 45
<< m1 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2c >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 46
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 157 192 158 193  0 t = 1
rlabel pdiffusion 160 192 161 193  0 t = 2
rlabel pdiffusion 157 197 158 198  0 t = 3
rlabel pdiffusion 160 197 161 198  0 t = 4
rlabel pdiffusion 156 192 162 198 0 cell no = 47
<< m1 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2c >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< labels >>
rlabel pdiffusion 175 48 176 49  0 t = 1
rlabel pdiffusion 178 48 179 49  0 t = 2
rlabel pdiffusion 175 53 176 54  0 t = 3
rlabel pdiffusion 178 53 179 54  0 t = 4
rlabel pdiffusion 174 48 180 54 0 cell no = 48
<< m1 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2c >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< labels >>
rlabel pdiffusion 229 102 230 103  0 t = 1
rlabel pdiffusion 232 102 233 103  0 t = 2
rlabel pdiffusion 229 107 230 108  0 t = 3
rlabel pdiffusion 232 107 233 108  0 t = 4
rlabel pdiffusion 228 102 234 108 0 cell no = 49
<< m1 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2c >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< labels >>
rlabel pdiffusion 85 138 86 139  0 t = 1
rlabel pdiffusion 88 138 89 139  0 t = 2
rlabel pdiffusion 85 143 86 144  0 t = 3
rlabel pdiffusion 88 143 89 144  0 t = 4
rlabel pdiffusion 84 138 90 144 0 cell no = 50
<< m1 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2c >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< labels >>
rlabel pdiffusion 247 156 248 157  0 t = 1
rlabel pdiffusion 250 156 251 157  0 t = 2
rlabel pdiffusion 247 161 248 162  0 t = 3
rlabel pdiffusion 250 161 251 162  0 t = 4
rlabel pdiffusion 246 156 252 162 0 cell no = 51
<< m1 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2c >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 52
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 229 30 230 31  0 t = 1
rlabel pdiffusion 232 30 233 31  0 t = 2
rlabel pdiffusion 229 35 230 36  0 t = 3
rlabel pdiffusion 232 35 233 36  0 t = 4
rlabel pdiffusion 228 30 234 36 0 cell no = 53
<< m1 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2c >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< labels >>
rlabel pdiffusion 211 84 212 85  0 t = 1
rlabel pdiffusion 214 84 215 85  0 t = 2
rlabel pdiffusion 211 89 212 90  0 t = 3
rlabel pdiffusion 214 89 215 90  0 t = 4
rlabel pdiffusion 210 84 216 90 0 cell no = 54
<< m1 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2c >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< labels >>
rlabel pdiffusion 229 66 230 67  0 t = 1
rlabel pdiffusion 232 66 233 67  0 t = 2
rlabel pdiffusion 229 71 230 72  0 t = 3
rlabel pdiffusion 232 71 233 72  0 t = 4
rlabel pdiffusion 228 66 234 72 0 cell no = 55
<< m1 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2c >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< labels >>
rlabel pdiffusion 193 156 194 157  0 t = 1
rlabel pdiffusion 196 156 197 157  0 t = 2
rlabel pdiffusion 193 161 194 162  0 t = 3
rlabel pdiffusion 196 161 197 162  0 t = 4
rlabel pdiffusion 192 156 198 162 0 cell no = 56
<< m1 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2c >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 57
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 157 48 158 49  0 t = 1
rlabel pdiffusion 160 48 161 49  0 t = 2
rlabel pdiffusion 157 53 158 54  0 t = 3
rlabel pdiffusion 160 53 161 54  0 t = 4
rlabel pdiffusion 156 48 162 54 0 cell no = 58
<< m1 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2c >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 59
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 60
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 49 138 50 139  0 t = 1
rlabel pdiffusion 52 138 53 139  0 t = 2
rlabel pdiffusion 49 143 50 144  0 t = 3
rlabel pdiffusion 52 143 53 144  0 t = 4
rlabel pdiffusion 48 138 54 144 0 cell no = 61
<< m1 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2c >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< labels >>
rlabel pdiffusion 211 228 212 229  0 t = 1
rlabel pdiffusion 214 228 215 229  0 t = 2
rlabel pdiffusion 211 233 212 234  0 t = 3
rlabel pdiffusion 214 233 215 234  0 t = 4
rlabel pdiffusion 210 228 216 234 0 cell no = 62
<< m1 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2c >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< labels >>
rlabel pdiffusion 103 120 104 121  0 t = 1
rlabel pdiffusion 106 120 107 121  0 t = 2
rlabel pdiffusion 103 125 104 126  0 t = 3
rlabel pdiffusion 106 125 107 126  0 t = 4
rlabel pdiffusion 102 120 108 126 0 cell no = 63
<< m1 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2c >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< labels >>
rlabel pdiffusion 247 102 248 103  0 t = 1
rlabel pdiffusion 250 102 251 103  0 t = 2
rlabel pdiffusion 247 107 248 108  0 t = 3
rlabel pdiffusion 250 107 251 108  0 t = 4
rlabel pdiffusion 246 102 252 108 0 cell no = 64
<< m1 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2c >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 65
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 229 174 230 175  0 t = 1
rlabel pdiffusion 232 174 233 175  0 t = 2
rlabel pdiffusion 229 179 230 180  0 t = 3
rlabel pdiffusion 232 179 233 180  0 t = 4
rlabel pdiffusion 228 174 234 180 0 cell no = 66
<< m1 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2c >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< labels >>
rlabel pdiffusion 13 120 14 121  0 t = 1
rlabel pdiffusion 16 120 17 121  0 t = 2
rlabel pdiffusion 13 125 14 126  0 t = 3
rlabel pdiffusion 16 125 17 126  0 t = 4
rlabel pdiffusion 12 120 18 126 0 cell no = 67
<< m1 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2c >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 68
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 69
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 211 48 212 49  0 t = 1
rlabel pdiffusion 214 48 215 49  0 t = 2
rlabel pdiffusion 211 53 212 54  0 t = 3
rlabel pdiffusion 214 53 215 54  0 t = 4
rlabel pdiffusion 210 48 216 54 0 cell no = 70
<< m1 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2c >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< labels >>
rlabel pdiffusion 229 138 230 139  0 t = 1
rlabel pdiffusion 232 138 233 139  0 t = 2
rlabel pdiffusion 229 143 230 144  0 t = 3
rlabel pdiffusion 232 143 233 144  0 t = 4
rlabel pdiffusion 228 138 234 144 0 cell no = 71
<< m1 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2c >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 72
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 49 192 50 193  0 t = 1
rlabel pdiffusion 52 192 53 193  0 t = 2
rlabel pdiffusion 49 197 50 198  0 t = 3
rlabel pdiffusion 52 197 53 198  0 t = 4
rlabel pdiffusion 48 192 54 198 0 cell no = 73
<< m1 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2c >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 74
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 157 210 158 211  0 t = 1
rlabel pdiffusion 160 210 161 211  0 t = 2
rlabel pdiffusion 157 215 158 216  0 t = 3
rlabel pdiffusion 160 215 161 216  0 t = 4
rlabel pdiffusion 156 210 162 216 0 cell no = 75
<< m1 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2c >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< labels >>
rlabel pdiffusion 103 228 104 229  0 t = 1
rlabel pdiffusion 106 228 107 229  0 t = 2
rlabel pdiffusion 103 233 104 234  0 t = 3
rlabel pdiffusion 106 233 107 234  0 t = 4
rlabel pdiffusion 102 228 108 234 0 cell no = 76
<< m1 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2c >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< labels >>
rlabel pdiffusion 31 156 32 157  0 t = 1
rlabel pdiffusion 34 156 35 157  0 t = 2
rlabel pdiffusion 31 161 32 162  0 t = 3
rlabel pdiffusion 34 161 35 162  0 t = 4
rlabel pdiffusion 30 156 36 162 0 cell no = 77
<< m1 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2c >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 78
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 31 84 32 85  0 t = 1
rlabel pdiffusion 34 84 35 85  0 t = 2
rlabel pdiffusion 31 89 32 90  0 t = 3
rlabel pdiffusion 34 89 35 90  0 t = 4
rlabel pdiffusion 30 84 36 90 0 cell no = 79
<< m1 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2c >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< labels >>
rlabel pdiffusion 49 156 50 157  0 t = 1
rlabel pdiffusion 52 156 53 157  0 t = 2
rlabel pdiffusion 49 161 50 162  0 t = 3
rlabel pdiffusion 52 161 53 162  0 t = 4
rlabel pdiffusion 48 156 54 162 0 cell no = 80
<< m1 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2c >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< labels >>
rlabel pdiffusion 229 84 230 85  0 t = 1
rlabel pdiffusion 232 84 233 85  0 t = 2
rlabel pdiffusion 229 89 230 90  0 t = 3
rlabel pdiffusion 232 89 233 90  0 t = 4
rlabel pdiffusion 228 84 234 90 0 cell no = 81
<< m1 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2c >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< labels >>
rlabel pdiffusion 211 210 212 211  0 t = 1
rlabel pdiffusion 214 210 215 211  0 t = 2
rlabel pdiffusion 211 215 212 216  0 t = 3
rlabel pdiffusion 214 215 215 216  0 t = 4
rlabel pdiffusion 210 210 216 216 0 cell no = 82
<< m1 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2c >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< labels >>
rlabel pdiffusion 157 30 158 31  0 t = 1
rlabel pdiffusion 160 30 161 31  0 t = 2
rlabel pdiffusion 157 35 158 36  0 t = 3
rlabel pdiffusion 160 35 161 36  0 t = 4
rlabel pdiffusion 156 30 162 36 0 cell no = 83
<< m1 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2c >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< labels >>
rlabel pdiffusion 157 156 158 157  0 t = 1
rlabel pdiffusion 160 156 161 157  0 t = 2
rlabel pdiffusion 157 161 158 162  0 t = 3
rlabel pdiffusion 160 161 161 162  0 t = 4
rlabel pdiffusion 156 156 162 162 0 cell no = 84
<< m1 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2c >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< labels >>
rlabel pdiffusion 31 12 32 13  0 t = 1
rlabel pdiffusion 34 12 35 13  0 t = 2
rlabel pdiffusion 31 17 32 18  0 t = 3
rlabel pdiffusion 34 17 35 18  0 t = 4
rlabel pdiffusion 30 12 36 18 0 cell no = 85
<< m1 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2c >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< labels >>
rlabel pdiffusion 13 246 14 247  0 t = 1
rlabel pdiffusion 16 246 17 247  0 t = 2
rlabel pdiffusion 13 251 14 252  0 t = 3
rlabel pdiffusion 16 251 17 252  0 t = 4
rlabel pdiffusion 12 246 18 252 0 cell no = 86
<< m1 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2c >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< labels >>
rlabel pdiffusion 49 174 50 175  0 t = 1
rlabel pdiffusion 52 174 53 175  0 t = 2
rlabel pdiffusion 49 179 50 180  0 t = 3
rlabel pdiffusion 52 179 53 180  0 t = 4
rlabel pdiffusion 48 174 54 180 0 cell no = 87
<< m1 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2c >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< labels >>
rlabel pdiffusion 211 12 212 13  0 t = 1
rlabel pdiffusion 214 12 215 13  0 t = 2
rlabel pdiffusion 211 17 212 18  0 t = 3
rlabel pdiffusion 214 17 215 18  0 t = 4
rlabel pdiffusion 210 12 216 18 0 cell no = 88
<< m1 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2c >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 89
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 90
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 229 192 230 193  0 t = 1
rlabel pdiffusion 232 192 233 193  0 t = 2
rlabel pdiffusion 229 197 230 198  0 t = 3
rlabel pdiffusion 232 197 233 198  0 t = 4
rlabel pdiffusion 228 192 234 198 0 cell no = 91
<< m1 >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< m2 >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< m2c >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< labels >>
rlabel pdiffusion 211 30 212 31  0 t = 1
rlabel pdiffusion 214 30 215 31  0 t = 2
rlabel pdiffusion 211 35 212 36  0 t = 3
rlabel pdiffusion 214 35 215 36  0 t = 4
rlabel pdiffusion 210 30 216 36 0 cell no = 92
<< m1 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2c >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< labels >>
rlabel pdiffusion 157 246 158 247  0 t = 1
rlabel pdiffusion 160 246 161 247  0 t = 2
rlabel pdiffusion 157 251 158 252  0 t = 3
rlabel pdiffusion 160 251 161 252  0 t = 4
rlabel pdiffusion 156 246 162 252 0 cell no = 93
<< m1 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2c >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< labels >>
rlabel pdiffusion 247 84 248 85  0 t = 1
rlabel pdiffusion 250 84 251 85  0 t = 2
rlabel pdiffusion 247 89 248 90  0 t = 3
rlabel pdiffusion 250 89 251 90  0 t = 4
rlabel pdiffusion 246 84 252 90 0 cell no = 94
<< m1 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2c >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< labels >>
rlabel pdiffusion 139 30 140 31  0 t = 1
rlabel pdiffusion 142 30 143 31  0 t = 2
rlabel pdiffusion 139 35 140 36  0 t = 3
rlabel pdiffusion 142 35 143 36  0 t = 4
rlabel pdiffusion 138 30 144 36 0 cell no = 95
<< m1 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2c >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< labels >>
rlabel pdiffusion 85 210 86 211  0 t = 1
rlabel pdiffusion 88 210 89 211  0 t = 2
rlabel pdiffusion 85 215 86 216  0 t = 3
rlabel pdiffusion 88 215 89 216  0 t = 4
rlabel pdiffusion 84 210 90 216 0 cell no = 96
<< m1 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2c >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< labels >>
rlabel pdiffusion 247 138 248 139  0 t = 1
rlabel pdiffusion 250 138 251 139  0 t = 2
rlabel pdiffusion 247 143 248 144  0 t = 3
rlabel pdiffusion 250 143 251 144  0 t = 4
rlabel pdiffusion 246 138 252 144 0 cell no = 97
<< m1 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2c >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 98
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 247 120 248 121  0 t = 1
rlabel pdiffusion 250 120 251 121  0 t = 2
rlabel pdiffusion 247 125 248 126  0 t = 3
rlabel pdiffusion 250 125 251 126  0 t = 4
rlabel pdiffusion 246 120 252 126 0 cell no = 99
<< m1 >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< m2 >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< m2c >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< labels >>
rlabel pdiffusion 13 156 14 157  0 t = 1
rlabel pdiffusion 16 156 17 157  0 t = 2
rlabel pdiffusion 13 161 14 162  0 t = 3
rlabel pdiffusion 16 161 17 162  0 t = 4
rlabel pdiffusion 12 156 18 162 0 cell no = 100
<< m1 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2c >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< labels >>
rlabel pdiffusion 175 192 176 193  0 t = 1
rlabel pdiffusion 178 192 179 193  0 t = 2
rlabel pdiffusion 175 197 176 198  0 t = 3
rlabel pdiffusion 178 197 179 198  0 t = 4
rlabel pdiffusion 174 192 180 198 0 cell no = 101
<< m1 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2c >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< labels >>
rlabel pdiffusion 85 228 86 229  0 t = 1
rlabel pdiffusion 88 228 89 229  0 t = 2
rlabel pdiffusion 85 233 86 234  0 t = 3
rlabel pdiffusion 88 233 89 234  0 t = 4
rlabel pdiffusion 84 228 90 234 0 cell no = 102
<< m1 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2c >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< labels >>
rlabel pdiffusion 175 30 176 31  0 t = 1
rlabel pdiffusion 178 30 179 31  0 t = 2
rlabel pdiffusion 175 35 176 36  0 t = 3
rlabel pdiffusion 178 35 179 36  0 t = 4
rlabel pdiffusion 174 30 180 36 0 cell no = 103
<< m1 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2c >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< labels >>
rlabel pdiffusion 13 228 14 229  0 t = 1
rlabel pdiffusion 16 228 17 229  0 t = 2
rlabel pdiffusion 13 233 14 234  0 t = 3
rlabel pdiffusion 16 233 17 234  0 t = 4
rlabel pdiffusion 12 228 18 234 0 cell no = 104
<< m1 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2c >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< labels >>
rlabel pdiffusion 31 192 32 193  0 t = 1
rlabel pdiffusion 34 192 35 193  0 t = 2
rlabel pdiffusion 31 197 32 198  0 t = 3
rlabel pdiffusion 34 197 35 198  0 t = 4
rlabel pdiffusion 30 192 36 198 0 cell no = 105
<< m1 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2c >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< labels >>
rlabel pdiffusion 67 120 68 121  0 t = 1
rlabel pdiffusion 70 120 71 121  0 t = 2
rlabel pdiffusion 67 125 68 126  0 t = 3
rlabel pdiffusion 70 125 71 126  0 t = 4
rlabel pdiffusion 66 120 72 126 0 cell no = 106
<< m1 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2c >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< labels >>
rlabel pdiffusion 229 210 230 211  0 t = 1
rlabel pdiffusion 232 210 233 211  0 t = 2
rlabel pdiffusion 229 215 230 216  0 t = 3
rlabel pdiffusion 232 215 233 216  0 t = 4
rlabel pdiffusion 228 210 234 216 0 cell no = 107
<< m1 >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< m2 >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< m2c >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 108
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 109
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 193 192 194 193  0 t = 1
rlabel pdiffusion 196 192 197 193  0 t = 2
rlabel pdiffusion 193 197 194 198  0 t = 3
rlabel pdiffusion 196 197 197 198  0 t = 4
rlabel pdiffusion 192 192 198 198 0 cell no = 110
<< m1 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2c >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< labels >>
rlabel pdiffusion 85 120 86 121  0 t = 1
rlabel pdiffusion 88 120 89 121  0 t = 2
rlabel pdiffusion 85 125 86 126  0 t = 3
rlabel pdiffusion 88 125 89 126  0 t = 4
rlabel pdiffusion 84 120 90 126 0 cell no = 111
<< m1 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2c >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< labels >>
rlabel pdiffusion 157 228 158 229  0 t = 1
rlabel pdiffusion 160 228 161 229  0 t = 2
rlabel pdiffusion 157 233 158 234  0 t = 3
rlabel pdiffusion 160 233 161 234  0 t = 4
rlabel pdiffusion 156 228 162 234 0 cell no = 112
<< m1 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2c >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< labels >>
rlabel pdiffusion 211 192 212 193  0 t = 1
rlabel pdiffusion 214 192 215 193  0 t = 2
rlabel pdiffusion 211 197 212 198  0 t = 3
rlabel pdiffusion 214 197 215 198  0 t = 4
rlabel pdiffusion 210 192 216 198 0 cell no = 113
<< m1 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2c >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< labels >>
rlabel pdiffusion 49 228 50 229  0 t = 1
rlabel pdiffusion 52 228 53 229  0 t = 2
rlabel pdiffusion 49 233 50 234  0 t = 3
rlabel pdiffusion 52 233 53 234  0 t = 4
rlabel pdiffusion 48 228 54 234 0 cell no = 114
<< m1 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2c >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 115
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 116
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 157 174 158 175  0 t = 1
rlabel pdiffusion 160 174 161 175  0 t = 2
rlabel pdiffusion 157 179 158 180  0 t = 3
rlabel pdiffusion 160 179 161 180  0 t = 4
rlabel pdiffusion 156 174 162 180 0 cell no = 117
<< m1 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2c >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< labels >>
rlabel pdiffusion 85 246 86 247  0 t = 1
rlabel pdiffusion 88 246 89 247  0 t = 2
rlabel pdiffusion 85 251 86 252  0 t = 3
rlabel pdiffusion 88 251 89 252  0 t = 4
rlabel pdiffusion 84 246 90 252 0 cell no = 118
<< m1 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2c >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< labels >>
rlabel pdiffusion 67 138 68 139  0 t = 1
rlabel pdiffusion 70 138 71 139  0 t = 2
rlabel pdiffusion 67 143 68 144  0 t = 3
rlabel pdiffusion 70 143 71 144  0 t = 4
rlabel pdiffusion 66 138 72 144 0 cell no = 119
<< m1 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2c >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< labels >>
rlabel pdiffusion 103 246 104 247  0 t = 1
rlabel pdiffusion 106 246 107 247  0 t = 2
rlabel pdiffusion 103 251 104 252  0 t = 3
rlabel pdiffusion 106 251 107 252  0 t = 4
rlabel pdiffusion 102 246 108 252 0 cell no = 120
<< m1 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2c >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< labels >>
rlabel pdiffusion 121 210 122 211  0 t = 1
rlabel pdiffusion 124 210 125 211  0 t = 2
rlabel pdiffusion 121 215 122 216  0 t = 3
rlabel pdiffusion 124 215 125 216  0 t = 4
rlabel pdiffusion 120 210 126 216 0 cell no = 121
<< m1 >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< m2 >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< m2c >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< labels >>
rlabel pdiffusion 175 174 176 175  0 t = 1
rlabel pdiffusion 178 174 179 175  0 t = 2
rlabel pdiffusion 175 179 176 180  0 t = 3
rlabel pdiffusion 178 179 179 180  0 t = 4
rlabel pdiffusion 174 174 180 180 0 cell no = 122
<< m1 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2c >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< labels >>
rlabel pdiffusion 175 138 176 139  0 t = 1
rlabel pdiffusion 178 138 179 139  0 t = 2
rlabel pdiffusion 175 143 176 144  0 t = 3
rlabel pdiffusion 178 143 179 144  0 t = 4
rlabel pdiffusion 174 138 180 144 0 cell no = 123
<< m1 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2c >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 124
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 247 192 248 193  0 t = 1
rlabel pdiffusion 250 192 251 193  0 t = 2
rlabel pdiffusion 247 197 248 198  0 t = 3
rlabel pdiffusion 250 197 251 198  0 t = 4
rlabel pdiffusion 246 192 252 198 0 cell no = 125
<< m1 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2c >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 126
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 49 246 50 247  0 t = 1
rlabel pdiffusion 52 246 53 247  0 t = 2
rlabel pdiffusion 49 251 50 252  0 t = 3
rlabel pdiffusion 52 251 53 252  0 t = 4
rlabel pdiffusion 48 246 54 252 0 cell no = 127
<< m1 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2c >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< labels >>
rlabel pdiffusion 103 192 104 193  0 t = 1
rlabel pdiffusion 106 192 107 193  0 t = 2
rlabel pdiffusion 103 197 104 198  0 t = 3
rlabel pdiffusion 106 197 107 198  0 t = 4
rlabel pdiffusion 102 192 108 198 0 cell no = 128
<< m1 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2c >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 129
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 13 210 14 211  0 t = 1
rlabel pdiffusion 16 210 17 211  0 t = 2
rlabel pdiffusion 13 215 14 216  0 t = 3
rlabel pdiffusion 16 215 17 216  0 t = 4
rlabel pdiffusion 12 210 18 216 0 cell no = 130
<< m1 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2c >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 131
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 193 12 194 13  0 t = 1
rlabel pdiffusion 196 12 197 13  0 t = 2
rlabel pdiffusion 193 17 194 18  0 t = 3
rlabel pdiffusion 196 17 197 18  0 t = 4
rlabel pdiffusion 192 12 198 18 0 cell no = 132
<< m1 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2c >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< labels >>
rlabel pdiffusion 121 192 122 193  0 t = 1
rlabel pdiffusion 124 192 125 193  0 t = 2
rlabel pdiffusion 121 197 122 198  0 t = 3
rlabel pdiffusion 124 197 125 198  0 t = 4
rlabel pdiffusion 120 192 126 198 0 cell no = 133
<< m1 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2c >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< labels >>
rlabel pdiffusion 139 120 140 121  0 t = 1
rlabel pdiffusion 142 120 143 121  0 t = 2
rlabel pdiffusion 139 125 140 126  0 t = 3
rlabel pdiffusion 142 125 143 126  0 t = 4
rlabel pdiffusion 138 120 144 126 0 cell no = 134
<< m1 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2c >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 135
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 121 102 122 103  0 t = 1
rlabel pdiffusion 124 102 125 103  0 t = 2
rlabel pdiffusion 121 107 122 108  0 t = 3
rlabel pdiffusion 124 107 125 108  0 t = 4
rlabel pdiffusion 120 102 126 108 0 cell no = 136
<< m1 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2c >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< labels >>
rlabel pdiffusion 211 138 212 139  0 t = 1
rlabel pdiffusion 214 138 215 139  0 t = 2
rlabel pdiffusion 211 143 212 144  0 t = 3
rlabel pdiffusion 214 143 215 144  0 t = 4
rlabel pdiffusion 210 138 216 144 0 cell no = 137
<< m1 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2c >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< labels >>
rlabel pdiffusion 175 102 176 103  0 t = 1
rlabel pdiffusion 178 102 179 103  0 t = 2
rlabel pdiffusion 175 107 176 108  0 t = 3
rlabel pdiffusion 178 107 179 108  0 t = 4
rlabel pdiffusion 174 102 180 108 0 cell no = 138
<< m1 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2c >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< labels >>
rlabel pdiffusion 175 84 176 85  0 t = 1
rlabel pdiffusion 178 84 179 85  0 t = 2
rlabel pdiffusion 175 89 176 90  0 t = 3
rlabel pdiffusion 178 89 179 90  0 t = 4
rlabel pdiffusion 174 84 180 90 0 cell no = 139
<< m1 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2c >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< labels >>
rlabel pdiffusion 157 12 158 13  0 t = 1
rlabel pdiffusion 160 12 161 13  0 t = 2
rlabel pdiffusion 157 17 158 18  0 t = 3
rlabel pdiffusion 160 17 161 18  0 t = 4
rlabel pdiffusion 156 12 162 18 0 cell no = 140
<< m1 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2c >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 141
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 67 246 68 247  0 t = 1
rlabel pdiffusion 70 246 71 247  0 t = 2
rlabel pdiffusion 67 251 68 252  0 t = 3
rlabel pdiffusion 70 251 71 252  0 t = 4
rlabel pdiffusion 66 246 72 252 0 cell no = 142
<< m1 >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< m2 >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< m2c >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< labels >>
rlabel pdiffusion 229 12 230 13  0 t = 1
rlabel pdiffusion 232 12 233 13  0 t = 2
rlabel pdiffusion 229 17 230 18  0 t = 3
rlabel pdiffusion 232 17 233 18  0 t = 4
rlabel pdiffusion 228 12 234 18 0 cell no = 143
<< m1 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2c >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< labels >>
rlabel pdiffusion 121 138 122 139  0 t = 1
rlabel pdiffusion 124 138 125 139  0 t = 2
rlabel pdiffusion 121 143 122 144  0 t = 3
rlabel pdiffusion 124 143 125 144  0 t = 4
rlabel pdiffusion 120 138 126 144 0 cell no = 144
<< m1 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2c >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< labels >>
rlabel pdiffusion 31 210 32 211  0 t = 1
rlabel pdiffusion 34 210 35 211  0 t = 2
rlabel pdiffusion 31 215 32 216  0 t = 3
rlabel pdiffusion 34 215 35 216  0 t = 4
rlabel pdiffusion 30 210 36 216 0 cell no = 145
<< m1 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2c >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 146
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 139 48 140 49  0 t = 1
rlabel pdiffusion 142 48 143 49  0 t = 2
rlabel pdiffusion 139 53 140 54  0 t = 3
rlabel pdiffusion 142 53 143 54  0 t = 4
rlabel pdiffusion 138 48 144 54 0 cell no = 147
<< m1 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2c >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< labels >>
rlabel pdiffusion 67 210 68 211  0 t = 1
rlabel pdiffusion 70 210 71 211  0 t = 2
rlabel pdiffusion 67 215 68 216  0 t = 3
rlabel pdiffusion 70 215 71 216  0 t = 4
rlabel pdiffusion 66 210 72 216 0 cell no = 148
<< m1 >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< m2 >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< m2c >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 149
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 193 210 194 211  0 t = 1
rlabel pdiffusion 196 210 197 211  0 t = 2
rlabel pdiffusion 193 215 194 216  0 t = 3
rlabel pdiffusion 196 215 197 216  0 t = 4
rlabel pdiffusion 192 210 198 216 0 cell no = 150
<< m1 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2c >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< labels >>
rlabel pdiffusion 175 210 176 211  0 t = 1
rlabel pdiffusion 178 210 179 211  0 t = 2
rlabel pdiffusion 175 215 176 216  0 t = 3
rlabel pdiffusion 178 215 179 216  0 t = 4
rlabel pdiffusion 174 210 180 216 0 cell no = 151
<< m1 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2c >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< labels >>
rlabel pdiffusion 31 246 32 247  0 t = 1
rlabel pdiffusion 34 246 35 247  0 t = 2
rlabel pdiffusion 31 251 32 252  0 t = 3
rlabel pdiffusion 34 251 35 252  0 t = 4
rlabel pdiffusion 30 246 36 252 0 cell no = 152
<< m1 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2c >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< labels >>
rlabel pdiffusion 247 210 248 211  0 t = 1
rlabel pdiffusion 250 210 251 211  0 t = 2
rlabel pdiffusion 247 215 248 216  0 t = 3
rlabel pdiffusion 250 215 251 216  0 t = 4
rlabel pdiffusion 246 210 252 216 0 cell no = 153
<< m1 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2c >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< labels >>
rlabel pdiffusion 139 228 140 229  0 t = 1
rlabel pdiffusion 142 228 143 229  0 t = 2
rlabel pdiffusion 139 233 140 234  0 t = 3
rlabel pdiffusion 142 233 143 234  0 t = 4
rlabel pdiffusion 138 228 144 234 0 cell no = 154
<< m1 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2c >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< labels >>
rlabel pdiffusion 13 174 14 175  0 t = 1
rlabel pdiffusion 16 174 17 175  0 t = 2
rlabel pdiffusion 13 179 14 180  0 t = 3
rlabel pdiffusion 16 179 17 180  0 t = 4
rlabel pdiffusion 12 174 18 180 0 cell no = 155
<< m1 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2c >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< labels >>
rlabel pdiffusion 139 12 140 13  0 t = 1
rlabel pdiffusion 142 12 143 13  0 t = 2
rlabel pdiffusion 139 17 140 18  0 t = 3
rlabel pdiffusion 142 17 143 18  0 t = 4
rlabel pdiffusion 138 12 144 18 0 cell no = 156
<< m1 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2c >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< labels >>
rlabel pdiffusion 211 156 212 157  0 t = 1
rlabel pdiffusion 214 156 215 157  0 t = 2
rlabel pdiffusion 211 161 212 162  0 t = 3
rlabel pdiffusion 214 161 215 162  0 t = 4
rlabel pdiffusion 210 156 216 162 0 cell no = 157
<< m1 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2c >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< labels >>
rlabel pdiffusion 157 138 158 139  0 t = 1
rlabel pdiffusion 160 138 161 139  0 t = 2
rlabel pdiffusion 157 143 158 144  0 t = 3
rlabel pdiffusion 160 143 161 144  0 t = 4
rlabel pdiffusion 156 138 162 144 0 cell no = 158
<< m1 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2c >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< labels >>
rlabel pdiffusion 85 156 86 157  0 t = 1
rlabel pdiffusion 88 156 89 157  0 t = 2
rlabel pdiffusion 85 161 86 162  0 t = 3
rlabel pdiffusion 88 161 89 162  0 t = 4
rlabel pdiffusion 84 156 90 162 0 cell no = 159
<< m1 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2c >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< labels >>
rlabel pdiffusion 139 210 140 211  0 t = 1
rlabel pdiffusion 142 210 143 211  0 t = 2
rlabel pdiffusion 139 215 140 216  0 t = 3
rlabel pdiffusion 142 215 143 216  0 t = 4
rlabel pdiffusion 138 210 144 216 0 cell no = 160
<< m1 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2c >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< labels >>
rlabel pdiffusion 193 120 194 121  0 t = 1
rlabel pdiffusion 196 120 197 121  0 t = 2
rlabel pdiffusion 193 125 194 126  0 t = 3
rlabel pdiffusion 196 125 197 126  0 t = 4
rlabel pdiffusion 192 120 198 126 0 cell no = 161
<< m1 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2c >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< labels >>
rlabel pdiffusion 121 246 122 247  0 t = 1
rlabel pdiffusion 124 246 125 247  0 t = 2
rlabel pdiffusion 121 251 122 252  0 t = 3
rlabel pdiffusion 124 251 125 252  0 t = 4
rlabel pdiffusion 120 246 126 252 0 cell no = 162
<< m1 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2c >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< labels >>
rlabel pdiffusion 121 156 122 157  0 t = 1
rlabel pdiffusion 124 156 125 157  0 t = 2
rlabel pdiffusion 121 161 122 162  0 t = 3
rlabel pdiffusion 124 161 125 162  0 t = 4
rlabel pdiffusion 120 156 126 162 0 cell no = 163
<< m1 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2c >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< labels >>
rlabel pdiffusion 175 156 176 157  0 t = 1
rlabel pdiffusion 178 156 179 157  0 t = 2
rlabel pdiffusion 175 161 176 162  0 t = 3
rlabel pdiffusion 178 161 179 162  0 t = 4
rlabel pdiffusion 174 156 180 162 0 cell no = 164
<< m1 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2c >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< labels >>
rlabel pdiffusion 31 228 32 229  0 t = 1
rlabel pdiffusion 34 228 35 229  0 t = 2
rlabel pdiffusion 31 233 32 234  0 t = 3
rlabel pdiffusion 34 233 35 234  0 t = 4
rlabel pdiffusion 30 228 36 234 0 cell no = 165
<< m1 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2c >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< labels >>
rlabel pdiffusion 139 138 140 139  0 t = 1
rlabel pdiffusion 142 138 143 139  0 t = 2
rlabel pdiffusion 139 143 140 144  0 t = 3
rlabel pdiffusion 142 143 143 144  0 t = 4
rlabel pdiffusion 138 138 144 144 0 cell no = 166
<< m1 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2c >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< labels >>
rlabel pdiffusion 229 228 230 229  0 t = 1
rlabel pdiffusion 232 228 233 229  0 t = 2
rlabel pdiffusion 229 233 230 234  0 t = 3
rlabel pdiffusion 232 233 233 234  0 t = 4
rlabel pdiffusion 228 228 234 234 0 cell no = 167
<< m1 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2c >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< labels >>
rlabel pdiffusion 211 174 212 175  0 t = 1
rlabel pdiffusion 214 174 215 175  0 t = 2
rlabel pdiffusion 211 179 212 180  0 t = 3
rlabel pdiffusion 214 179 215 180  0 t = 4
rlabel pdiffusion 210 174 216 180 0 cell no = 168
<< m1 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2c >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< labels >>
rlabel pdiffusion 157 84 158 85  0 t = 1
rlabel pdiffusion 160 84 161 85  0 t = 2
rlabel pdiffusion 157 89 158 90  0 t = 3
rlabel pdiffusion 160 89 161 90  0 t = 4
rlabel pdiffusion 156 84 162 90 0 cell no = 169
<< m1 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2c >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< labels >>
rlabel pdiffusion 103 210 104 211  0 t = 1
rlabel pdiffusion 106 210 107 211  0 t = 2
rlabel pdiffusion 103 215 104 216  0 t = 3
rlabel pdiffusion 106 215 107 216  0 t = 4
rlabel pdiffusion 102 210 108 216 0 cell no = 170
<< m1 >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< m2 >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< m2c >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< labels >>
rlabel pdiffusion 67 156 68 157  0 t = 1
rlabel pdiffusion 70 156 71 157  0 t = 2
rlabel pdiffusion 67 161 68 162  0 t = 3
rlabel pdiffusion 70 161 71 162  0 t = 4
rlabel pdiffusion 66 156 72 162 0 cell no = 171
<< m1 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2c >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< labels >>
rlabel pdiffusion 31 174 32 175  0 t = 1
rlabel pdiffusion 34 174 35 175  0 t = 2
rlabel pdiffusion 31 179 32 180  0 t = 3
rlabel pdiffusion 34 179 35 180  0 t = 4
rlabel pdiffusion 30 174 36 180 0 cell no = 172
<< m1 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2c >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< labels >>
rlabel pdiffusion 211 120 212 121  0 t = 1
rlabel pdiffusion 214 120 215 121  0 t = 2
rlabel pdiffusion 211 125 212 126  0 t = 3
rlabel pdiffusion 214 125 215 126  0 t = 4
rlabel pdiffusion 210 120 216 126 0 cell no = 173
<< m1 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2c >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 174
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 121 174 122 175  0 t = 1
rlabel pdiffusion 124 174 125 175  0 t = 2
rlabel pdiffusion 121 179 122 180  0 t = 3
rlabel pdiffusion 124 179 125 180  0 t = 4
rlabel pdiffusion 120 174 126 180 0 cell no = 175
<< m1 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2c >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< labels >>
rlabel pdiffusion 139 246 140 247  0 t = 1
rlabel pdiffusion 142 246 143 247  0 t = 2
rlabel pdiffusion 139 251 140 252  0 t = 3
rlabel pdiffusion 142 251 143 252  0 t = 4
rlabel pdiffusion 138 246 144 252 0 cell no = 176
<< m1 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2c >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< labels >>
rlabel pdiffusion 31 138 32 139  0 t = 1
rlabel pdiffusion 34 138 35 139  0 t = 2
rlabel pdiffusion 31 143 32 144  0 t = 3
rlabel pdiffusion 34 143 35 144  0 t = 4
rlabel pdiffusion 30 138 36 144 0 cell no = 177
<< m1 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2c >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< labels >>
rlabel pdiffusion 85 174 86 175  0 t = 1
rlabel pdiffusion 88 174 89 175  0 t = 2
rlabel pdiffusion 85 179 86 180  0 t = 3
rlabel pdiffusion 88 179 89 180  0 t = 4
rlabel pdiffusion 84 174 90 180 0 cell no = 178
<< m1 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2c >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 179
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 139 156 140 157  0 t = 1
rlabel pdiffusion 142 156 143 157  0 t = 2
rlabel pdiffusion 139 161 140 162  0 t = 3
rlabel pdiffusion 142 161 143 162  0 t = 4
rlabel pdiffusion 138 156 144 162 0 cell no = 180
<< m1 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2c >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< end >> 
