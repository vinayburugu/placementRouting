magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 40 3 41 4 
<< m2 >>
rect 40 3 41 4 
<< m2c >>
rect 40 3 41 4 
<< m1 >>
rect 40 3 41 4 
<< m2 >>
rect 40 3 41 4 
<< m2 >>
rect 41 3 42 4 
<< m1 >>
rect 42 3 43 4 
<< m2 >>
rect 42 3 43 4 
<< m1 >>
rect 43 3 44 4 
<< m2 >>
rect 43 3 44 4 
<< m1 >>
rect 44 3 45 4 
<< m2 >>
rect 44 3 45 4 
<< m1 >>
rect 45 3 46 4 
<< m2 >>
rect 45 3 46 4 
<< m1 >>
rect 46 3 47 4 
<< m2 >>
rect 46 3 47 4 
<< m1 >>
rect 47 3 48 4 
<< m2 >>
rect 47 3 48 4 
<< m1 >>
rect 48 3 49 4 
<< m2 >>
rect 48 3 49 4 
<< m1 >>
rect 49 3 50 4 
<< m2 >>
rect 49 3 50 4 
<< m1 >>
rect 50 3 51 4 
<< m2 >>
rect 50 3 51 4 
<< m1 >>
rect 51 3 52 4 
<< m2 >>
rect 51 3 52 4 
<< m1 >>
rect 52 3 53 4 
<< m2 >>
rect 52 3 53 4 
<< m1 >>
rect 53 3 54 4 
<< m2 >>
rect 53 3 54 4 
<< m1 >>
rect 54 3 55 4 
<< m2 >>
rect 54 3 55 4 
<< m1 >>
rect 55 3 56 4 
<< m2 >>
rect 55 3 56 4 
<< m1 >>
rect 56 3 57 4 
<< m2 >>
rect 56 3 57 4 
<< m1 >>
rect 57 3 58 4 
<< m2 >>
rect 57 3 58 4 
<< m1 >>
rect 58 3 59 4 
<< m2 >>
rect 58 3 59 4 
<< m1 >>
rect 59 3 60 4 
<< m2 >>
rect 59 3 60 4 
<< m1 >>
rect 60 3 61 4 
<< m2 >>
rect 60 3 61 4 
<< m1 >>
rect 61 3 62 4 
<< m2 >>
rect 61 3 62 4 
<< m1 >>
rect 62 3 63 4 
<< m2 >>
rect 62 3 63 4 
<< m1 >>
rect 63 3 64 4 
<< m2 >>
rect 63 3 64 4 
<< m1 >>
rect 64 3 65 4 
<< m2 >>
rect 64 3 65 4 
<< m1 >>
rect 65 3 66 4 
<< m2 >>
rect 65 3 66 4 
<< m1 >>
rect 66 3 67 4 
<< m2 >>
rect 66 3 67 4 
<< m1 >>
rect 67 3 68 4 
<< m2 >>
rect 67 3 68 4 
<< m1 >>
rect 68 3 69 4 
<< m2 >>
rect 68 3 69 4 
<< m1 >>
rect 69 3 70 4 
<< m2 >>
rect 69 3 70 4 
<< m1 >>
rect 70 3 71 4 
<< m2 >>
rect 70 3 71 4 
<< m1 >>
rect 71 3 72 4 
<< m2 >>
rect 71 3 72 4 
<< m1 >>
rect 72 3 73 4 
<< m2 >>
rect 72 3 73 4 
<< m1 >>
rect 73 3 74 4 
<< m2 >>
rect 73 3 74 4 
<< m1 >>
rect 74 3 75 4 
<< m2 >>
rect 74 3 75 4 
<< m1 >>
rect 75 3 76 4 
<< m2 >>
rect 75 3 76 4 
<< m1 >>
rect 76 3 77 4 
<< m2 >>
rect 76 3 77 4 
<< m1 >>
rect 77 3 78 4 
<< m2 >>
rect 77 3 78 4 
<< m1 >>
rect 78 3 79 4 
<< m2 >>
rect 78 3 79 4 
<< m1 >>
rect 79 3 80 4 
<< m2 >>
rect 79 3 80 4 
<< m1 >>
rect 80 3 81 4 
<< m2 >>
rect 80 3 81 4 
<< m1 >>
rect 81 3 82 4 
<< m2 >>
rect 81 3 82 4 
<< m1 >>
rect 82 3 83 4 
<< m2 >>
rect 82 3 83 4 
<< m1 >>
rect 83 3 84 4 
<< m2 >>
rect 83 3 84 4 
<< m1 >>
rect 84 3 85 4 
<< m2 >>
rect 84 3 85 4 
<< m1 >>
rect 85 3 86 4 
<< m2 >>
rect 85 3 86 4 
<< m1 >>
rect 86 3 87 4 
<< m2 >>
rect 86 3 87 4 
<< m1 >>
rect 87 3 88 4 
<< m2 >>
rect 87 3 88 4 
<< m1 >>
rect 88 3 89 4 
<< m2 >>
rect 88 3 89 4 
<< m1 >>
rect 89 3 90 4 
<< m2 >>
rect 89 3 90 4 
<< m1 >>
rect 90 3 91 4 
<< m2 >>
rect 90 3 91 4 
<< m1 >>
rect 91 3 92 4 
<< m2 >>
rect 91 3 92 4 
<< m1 >>
rect 92 3 93 4 
<< m2 >>
rect 92 3 93 4 
<< m1 >>
rect 93 3 94 4 
<< m2 >>
rect 93 3 94 4 
<< m1 >>
rect 94 3 95 4 
<< m2 >>
rect 94 3 95 4 
<< m1 >>
rect 95 3 96 4 
<< m2 >>
rect 95 3 96 4 
<< m1 >>
rect 96 3 97 4 
<< m2 >>
rect 96 3 97 4 
<< m1 >>
rect 97 3 98 4 
<< m2 >>
rect 97 3 98 4 
<< m1 >>
rect 98 3 99 4 
<< m2 >>
rect 98 3 99 4 
<< m1 >>
rect 99 3 100 4 
<< m2 >>
rect 99 3 100 4 
<< m1 >>
rect 100 3 101 4 
<< m2 >>
rect 100 3 101 4 
<< m1 >>
rect 101 3 102 4 
<< m2 >>
rect 101 3 102 4 
<< m1 >>
rect 102 3 103 4 
<< m2 >>
rect 102 3 103 4 
<< m1 >>
rect 103 3 104 4 
<< m2 >>
rect 103 3 104 4 
<< m1 >>
rect 104 3 105 4 
<< m2 >>
rect 104 3 105 4 
<< m1 >>
rect 105 3 106 4 
<< m2 >>
rect 105 3 106 4 
<< m1 >>
rect 106 3 107 4 
<< m2 >>
rect 106 3 107 4 
<< m1 >>
rect 107 3 108 4 
<< m2 >>
rect 107 3 108 4 
<< m1 >>
rect 108 3 109 4 
<< m2 >>
rect 108 3 109 4 
<< m1 >>
rect 109 3 110 4 
<< m2 >>
rect 109 3 110 4 
<< m1 >>
rect 110 3 111 4 
<< m2 >>
rect 110 3 111 4 
<< m1 >>
rect 111 3 112 4 
<< m2 >>
rect 111 3 112 4 
<< m1 >>
rect 112 3 113 4 
<< m2 >>
rect 112 3 113 4 
<< m1 >>
rect 113 3 114 4 
<< m2 >>
rect 113 3 114 4 
<< m1 >>
rect 114 3 115 4 
<< m2 >>
rect 114 3 115 4 
<< m1 >>
rect 115 3 116 4 
<< m2 >>
rect 115 3 116 4 
<< m1 >>
rect 116 3 117 4 
<< m2 >>
rect 116 3 117 4 
<< m1 >>
rect 117 3 118 4 
<< m2 >>
rect 117 3 118 4 
<< m1 >>
rect 118 3 119 4 
<< m2 >>
rect 118 3 119 4 
<< m1 >>
rect 119 3 120 4 
<< m2 >>
rect 119 3 120 4 
<< m1 >>
rect 120 3 121 4 
<< m2 >>
rect 120 3 121 4 
<< m1 >>
rect 121 3 122 4 
<< m2 >>
rect 121 3 122 4 
<< m1 >>
rect 122 3 123 4 
<< m2 >>
rect 122 3 123 4 
<< m1 >>
rect 123 3 124 4 
<< m2 >>
rect 123 3 124 4 
<< m1 >>
rect 124 3 125 4 
<< m2 >>
rect 124 3 125 4 
<< m1 >>
rect 125 3 126 4 
<< m2 >>
rect 125 3 126 4 
<< m1 >>
rect 126 3 127 4 
<< m2 >>
rect 126 3 127 4 
<< m1 >>
rect 127 3 128 4 
<< m2 >>
rect 127 3 128 4 
<< m1 >>
rect 128 3 129 4 
<< m2 >>
rect 128 3 129 4 
<< m1 >>
rect 129 3 130 4 
<< m2 >>
rect 129 3 130 4 
<< m1 >>
rect 130 3 131 4 
<< m2 >>
rect 130 3 131 4 
<< m1 >>
rect 131 3 132 4 
<< m2 >>
rect 131 3 132 4 
<< m1 >>
rect 132 3 133 4 
<< m2 >>
rect 132 3 133 4 
<< m1 >>
rect 133 3 134 4 
<< m2 >>
rect 133 3 134 4 
<< m1 >>
rect 134 3 135 4 
<< m2 >>
rect 134 3 135 4 
<< m1 >>
rect 135 3 136 4 
<< m2 >>
rect 135 3 136 4 
<< m1 >>
rect 136 3 137 4 
<< m2 >>
rect 136 3 137 4 
<< m1 >>
rect 137 3 138 4 
<< m2 >>
rect 137 3 138 4 
<< m1 >>
rect 138 3 139 4 
<< m2 >>
rect 138 3 139 4 
<< m1 >>
rect 139 3 140 4 
<< m2 >>
rect 139 3 140 4 
<< m1 >>
rect 140 3 141 4 
<< m2 >>
rect 140 3 141 4 
<< m1 >>
rect 141 3 142 4 
<< m2 >>
rect 141 3 142 4 
<< m1 >>
rect 142 3 143 4 
<< m2 >>
rect 142 3 143 4 
<< m1 >>
rect 143 3 144 4 
<< m2 >>
rect 143 3 144 4 
<< m1 >>
rect 144 3 145 4 
<< m2 >>
rect 144 3 145 4 
<< m1 >>
rect 145 3 146 4 
<< m2 >>
rect 145 3 146 4 
<< m1 >>
rect 146 3 147 4 
<< m2 >>
rect 146 3 147 4 
<< m1 >>
rect 147 3 148 4 
<< m2 >>
rect 147 3 148 4 
<< m1 >>
rect 148 3 149 4 
<< m2 >>
rect 148 3 149 4 
<< m1 >>
rect 149 3 150 4 
<< m2 >>
rect 149 3 150 4 
<< m1 >>
rect 150 3 151 4 
<< m2 >>
rect 150 3 151 4 
<< m1 >>
rect 151 3 152 4 
<< m2 >>
rect 151 3 152 4 
<< m1 >>
rect 152 3 153 4 
<< m2 >>
rect 152 3 153 4 
<< m1 >>
rect 153 3 154 4 
<< m2 >>
rect 153 3 154 4 
<< m1 >>
rect 154 3 155 4 
<< m2 >>
rect 154 3 155 4 
<< m1 >>
rect 155 3 156 4 
<< m2 >>
rect 155 3 156 4 
<< m1 >>
rect 156 3 157 4 
<< m2 >>
rect 156 3 157 4 
<< m1 >>
rect 157 3 158 4 
<< m2 >>
rect 157 3 158 4 
<< m1 >>
rect 158 3 159 4 
<< m2 >>
rect 158 3 159 4 
<< m1 >>
rect 159 3 160 4 
<< m2 >>
rect 159 3 160 4 
<< m1 >>
rect 160 3 161 4 
<< m2 >>
rect 160 3 161 4 
<< m1 >>
rect 161 3 162 4 
<< m2 >>
rect 161 3 162 4 
<< m1 >>
rect 162 3 163 4 
<< m2 >>
rect 162 3 163 4 
<< m1 >>
rect 163 3 164 4 
<< m2 >>
rect 163 3 164 4 
<< m1 >>
rect 164 3 165 4 
<< m2 >>
rect 164 3 165 4 
<< m1 >>
rect 165 3 166 4 
<< m2 >>
rect 165 3 166 4 
<< m2 >>
rect 166 3 167 4 
<< m1 >>
rect 167 3 168 4 
<< m2 >>
rect 167 3 168 4 
<< m2c >>
rect 167 3 168 4 
<< m1 >>
rect 167 3 168 4 
<< m2 >>
rect 167 3 168 4 
<< m1 >>
rect 40 4 41 5 
<< m1 >>
rect 42 4 43 5 
<< m1 >>
rect 165 4 166 5 
<< m1 >>
rect 167 4 168 5 
<< m1 >>
rect 40 5 41 6 
<< m2 >>
rect 40 5 41 6 
<< m2c >>
rect 40 5 41 6 
<< m1 >>
rect 40 5 41 6 
<< m2 >>
rect 40 5 41 6 
<< m1 >>
rect 42 5 43 6 
<< m2 >>
rect 42 5 43 6 
<< m2c >>
rect 42 5 43 6 
<< m1 >>
rect 42 5 43 6 
<< m2 >>
rect 42 5 43 6 
<< m1 >>
rect 93 5 94 6 
<< m2 >>
rect 93 5 94 6 
<< m2c >>
rect 93 5 94 6 
<< m1 >>
rect 93 5 94 6 
<< m2 >>
rect 93 5 94 6 
<< m1 >>
rect 94 5 95 6 
<< m1 >>
rect 95 5 96 6 
<< m1 >>
rect 96 5 97 6 
<< m1 >>
rect 97 5 98 6 
<< m1 >>
rect 98 5 99 6 
<< m1 >>
rect 99 5 100 6 
<< m1 >>
rect 100 5 101 6 
<< m1 >>
rect 101 5 102 6 
<< m1 >>
rect 102 5 103 6 
<< m1 >>
rect 103 5 104 6 
<< m1 >>
rect 104 5 105 6 
<< m1 >>
rect 105 5 106 6 
<< m1 >>
rect 106 5 107 6 
<< m1 >>
rect 107 5 108 6 
<< m1 >>
rect 108 5 109 6 
<< m1 >>
rect 109 5 110 6 
<< m1 >>
rect 110 5 111 6 
<< m1 >>
rect 111 5 112 6 
<< m1 >>
rect 112 5 113 6 
<< m1 >>
rect 113 5 114 6 
<< m1 >>
rect 114 5 115 6 
<< m1 >>
rect 115 5 116 6 
<< m1 >>
rect 116 5 117 6 
<< m1 >>
rect 117 5 118 6 
<< m1 >>
rect 118 5 119 6 
<< m1 >>
rect 119 5 120 6 
<< m1 >>
rect 120 5 121 6 
<< m1 >>
rect 121 5 122 6 
<< m1 >>
rect 122 5 123 6 
<< m1 >>
rect 123 5 124 6 
<< m1 >>
rect 124 5 125 6 
<< m1 >>
rect 125 5 126 6 
<< m1 >>
rect 126 5 127 6 
<< m1 >>
rect 127 5 128 6 
<< m1 >>
rect 128 5 129 6 
<< m1 >>
rect 129 5 130 6 
<< m1 >>
rect 130 5 131 6 
<< m1 >>
rect 131 5 132 6 
<< m1 >>
rect 132 5 133 6 
<< m1 >>
rect 133 5 134 6 
<< m1 >>
rect 134 5 135 6 
<< m1 >>
rect 135 5 136 6 
<< m1 >>
rect 136 5 137 6 
<< m1 >>
rect 137 5 138 6 
<< m1 >>
rect 138 5 139 6 
<< m1 >>
rect 139 5 140 6 
<< m1 >>
rect 140 5 141 6 
<< m1 >>
rect 141 5 142 6 
<< m1 >>
rect 142 5 143 6 
<< m1 >>
rect 143 5 144 6 
<< m1 >>
rect 144 5 145 6 
<< m1 >>
rect 145 5 146 6 
<< m1 >>
rect 146 5 147 6 
<< m1 >>
rect 147 5 148 6 
<< m1 >>
rect 148 5 149 6 
<< m1 >>
rect 149 5 150 6 
<< m1 >>
rect 150 5 151 6 
<< m1 >>
rect 151 5 152 6 
<< m1 >>
rect 152 5 153 6 
<< m1 >>
rect 153 5 154 6 
<< m1 >>
rect 154 5 155 6 
<< m1 >>
rect 155 5 156 6 
<< m1 >>
rect 156 5 157 6 
<< m1 >>
rect 157 5 158 6 
<< m1 >>
rect 158 5 159 6 
<< m1 >>
rect 159 5 160 6 
<< m1 >>
rect 160 5 161 6 
<< m1 >>
rect 161 5 162 6 
<< m1 >>
rect 162 5 163 6 
<< m1 >>
rect 163 5 164 6 
<< m1 >>
rect 165 5 166 6 
<< m1 >>
rect 167 5 168 6 
<< m2 >>
rect 40 6 41 7 
<< m2 >>
rect 42 6 43 7 
<< m2 >>
rect 93 6 94 7 
<< m1 >>
rect 163 6 164 7 
<< m1 >>
rect 165 6 166 7 
<< m1 >>
rect 167 6 168 7 
<< m1 >>
rect 19 7 20 8 
<< m1 >>
rect 20 7 21 8 
<< m1 >>
rect 21 7 22 8 
<< m1 >>
rect 22 7 23 8 
<< m1 >>
rect 23 7 24 8 
<< m1 >>
rect 24 7 25 8 
<< m1 >>
rect 25 7 26 8 
<< m1 >>
rect 26 7 27 8 
<< m1 >>
rect 27 7 28 8 
<< m1 >>
rect 28 7 29 8 
<< m1 >>
rect 29 7 30 8 
<< m1 >>
rect 30 7 31 8 
<< m1 >>
rect 31 7 32 8 
<< m1 >>
rect 32 7 33 8 
<< m1 >>
rect 33 7 34 8 
<< m1 >>
rect 34 7 35 8 
<< m1 >>
rect 35 7 36 8 
<< m1 >>
rect 36 7 37 8 
<< m1 >>
rect 37 7 38 8 
<< m1 >>
rect 38 7 39 8 
<< m1 >>
rect 39 7 40 8 
<< m1 >>
rect 40 7 41 8 
<< m2 >>
rect 40 7 41 8 
<< m1 >>
rect 41 7 42 8 
<< m1 >>
rect 42 7 43 8 
<< m2 >>
rect 42 7 43 8 
<< m1 >>
rect 43 7 44 8 
<< m1 >>
rect 44 7 45 8 
<< m2 >>
rect 44 7 45 8 
<< m1 >>
rect 45 7 46 8 
<< m2 >>
rect 45 7 46 8 
<< m1 >>
rect 46 7 47 8 
<< m2 >>
rect 46 7 47 8 
<< m1 >>
rect 47 7 48 8 
<< m2 >>
rect 47 7 48 8 
<< m1 >>
rect 48 7 49 8 
<< m2 >>
rect 48 7 49 8 
<< m1 >>
rect 49 7 50 8 
<< m2 >>
rect 49 7 50 8 
<< m1 >>
rect 50 7 51 8 
<< m2 >>
rect 50 7 51 8 
<< m1 >>
rect 51 7 52 8 
<< m2 >>
rect 51 7 52 8 
<< m1 >>
rect 52 7 53 8 
<< m2 >>
rect 52 7 53 8 
<< m1 >>
rect 53 7 54 8 
<< m2 >>
rect 53 7 54 8 
<< m1 >>
rect 54 7 55 8 
<< m2 >>
rect 54 7 55 8 
<< m1 >>
rect 55 7 56 8 
<< m2 >>
rect 55 7 56 8 
<< m1 >>
rect 56 7 57 8 
<< m2 >>
rect 56 7 57 8 
<< m1 >>
rect 57 7 58 8 
<< m2 >>
rect 57 7 58 8 
<< m1 >>
rect 58 7 59 8 
<< m2 >>
rect 58 7 59 8 
<< m1 >>
rect 59 7 60 8 
<< m2 >>
rect 59 7 60 8 
<< m1 >>
rect 60 7 61 8 
<< m2 >>
rect 60 7 61 8 
<< m1 >>
rect 61 7 62 8 
<< m2 >>
rect 61 7 62 8 
<< m1 >>
rect 62 7 63 8 
<< m2 >>
rect 62 7 63 8 
<< m1 >>
rect 63 7 64 8 
<< m2 >>
rect 63 7 64 8 
<< m1 >>
rect 64 7 65 8 
<< m2 >>
rect 64 7 65 8 
<< m1 >>
rect 65 7 66 8 
<< m2 >>
rect 65 7 66 8 
<< m1 >>
rect 66 7 67 8 
<< m2 >>
rect 66 7 67 8 
<< m1 >>
rect 67 7 68 8 
<< m2 >>
rect 67 7 68 8 
<< m1 >>
rect 68 7 69 8 
<< m2 >>
rect 68 7 69 8 
<< m1 >>
rect 69 7 70 8 
<< m1 >>
rect 70 7 71 8 
<< m1 >>
rect 71 7 72 8 
<< m1 >>
rect 72 7 73 8 
<< m1 >>
rect 73 7 74 8 
<< m1 >>
rect 74 7 75 8 
<< m1 >>
rect 75 7 76 8 
<< m1 >>
rect 76 7 77 8 
<< m1 >>
rect 77 7 78 8 
<< m1 >>
rect 78 7 79 8 
<< m1 >>
rect 79 7 80 8 
<< m1 >>
rect 80 7 81 8 
<< m1 >>
rect 81 7 82 8 
<< m1 >>
rect 82 7 83 8 
<< m1 >>
rect 83 7 84 8 
<< m1 >>
rect 84 7 85 8 
<< m1 >>
rect 85 7 86 8 
<< m1 >>
rect 86 7 87 8 
<< m1 >>
rect 87 7 88 8 
<< m1 >>
rect 88 7 89 8 
<< m1 >>
rect 89 7 90 8 
<< m1 >>
rect 90 7 91 8 
<< m1 >>
rect 91 7 92 8 
<< m1 >>
rect 92 7 93 8 
<< m1 >>
rect 93 7 94 8 
<< m2 >>
rect 93 7 94 8 
<< m1 >>
rect 94 7 95 8 
<< m1 >>
rect 95 7 96 8 
<< m2 >>
rect 95 7 96 8 
<< m1 >>
rect 96 7 97 8 
<< m2 >>
rect 96 7 97 8 
<< m1 >>
rect 97 7 98 8 
<< m2 >>
rect 97 7 98 8 
<< m1 >>
rect 98 7 99 8 
<< m2 >>
rect 98 7 99 8 
<< m1 >>
rect 99 7 100 8 
<< m2 >>
rect 99 7 100 8 
<< m1 >>
rect 100 7 101 8 
<< m2 >>
rect 100 7 101 8 
<< m1 >>
rect 101 7 102 8 
<< m2 >>
rect 101 7 102 8 
<< m1 >>
rect 102 7 103 8 
<< m2 >>
rect 102 7 103 8 
<< m1 >>
rect 103 7 104 8 
<< m2 >>
rect 103 7 104 8 
<< m1 >>
rect 104 7 105 8 
<< m2 >>
rect 104 7 105 8 
<< m1 >>
rect 105 7 106 8 
<< m2 >>
rect 105 7 106 8 
<< m1 >>
rect 106 7 107 8 
<< m2 >>
rect 106 7 107 8 
<< m1 >>
rect 107 7 108 8 
<< m2 >>
rect 107 7 108 8 
<< m1 >>
rect 108 7 109 8 
<< m2 >>
rect 108 7 109 8 
<< m1 >>
rect 109 7 110 8 
<< m2 >>
rect 109 7 110 8 
<< m1 >>
rect 110 7 111 8 
<< m2 >>
rect 110 7 111 8 
<< m1 >>
rect 111 7 112 8 
<< m2 >>
rect 111 7 112 8 
<< m1 >>
rect 112 7 113 8 
<< m2 >>
rect 112 7 113 8 
<< m1 >>
rect 113 7 114 8 
<< m2 >>
rect 113 7 114 8 
<< m1 >>
rect 114 7 115 8 
<< m2 >>
rect 114 7 115 8 
<< m1 >>
rect 115 7 116 8 
<< m2 >>
rect 115 7 116 8 
<< m1 >>
rect 116 7 117 8 
<< m2 >>
rect 116 7 117 8 
<< m1 >>
rect 117 7 118 8 
<< m2 >>
rect 117 7 118 8 
<< m1 >>
rect 118 7 119 8 
<< m2 >>
rect 118 7 119 8 
<< m1 >>
rect 119 7 120 8 
<< m2 >>
rect 119 7 120 8 
<< m1 >>
rect 120 7 121 8 
<< m2 >>
rect 120 7 121 8 
<< m1 >>
rect 121 7 122 8 
<< m2 >>
rect 121 7 122 8 
<< m1 >>
rect 122 7 123 8 
<< m2 >>
rect 122 7 123 8 
<< m1 >>
rect 123 7 124 8 
<< m2 >>
rect 123 7 124 8 
<< m1 >>
rect 124 7 125 8 
<< m2 >>
rect 124 7 125 8 
<< m2 >>
rect 125 7 126 8 
<< m1 >>
rect 126 7 127 8 
<< m2 >>
rect 126 7 127 8 
<< m2c >>
rect 126 7 127 8 
<< m1 >>
rect 126 7 127 8 
<< m2 >>
rect 126 7 127 8 
<< m1 >>
rect 127 7 128 8 
<< m1 >>
rect 128 7 129 8 
<< m1 >>
rect 129 7 130 8 
<< m1 >>
rect 130 7 131 8 
<< m1 >>
rect 131 7 132 8 
<< m1 >>
rect 132 7 133 8 
<< m1 >>
rect 133 7 134 8 
<< m1 >>
rect 134 7 135 8 
<< m1 >>
rect 135 7 136 8 
<< m1 >>
rect 136 7 137 8 
<< m1 >>
rect 137 7 138 8 
<< m1 >>
rect 138 7 139 8 
<< m1 >>
rect 139 7 140 8 
<< m1 >>
rect 163 7 164 8 
<< m1 >>
rect 165 7 166 8 
<< m1 >>
rect 167 7 168 8 
<< m1 >>
rect 19 8 20 9 
<< m2 >>
rect 40 8 41 9 
<< m2 >>
rect 42 8 43 9 
<< m2 >>
rect 44 8 45 9 
<< m2 >>
rect 68 8 69 9 
<< m2 >>
rect 93 8 94 9 
<< m2 >>
rect 95 8 96 9 
<< m1 >>
rect 124 8 125 9 
<< m1 >>
rect 139 8 140 9 
<< m1 >>
rect 163 8 164 9 
<< m2 >>
rect 163 8 164 9 
<< m2c >>
rect 163 8 164 9 
<< m1 >>
rect 163 8 164 9 
<< m2 >>
rect 163 8 164 9 
<< m1 >>
rect 165 8 166 9 
<< m2 >>
rect 165 8 166 9 
<< m2c >>
rect 165 8 166 9 
<< m1 >>
rect 165 8 166 9 
<< m2 >>
rect 165 8 166 9 
<< m1 >>
rect 167 8 168 9 
<< m2 >>
rect 167 8 168 9 
<< m2c >>
rect 167 8 168 9 
<< m1 >>
rect 167 8 168 9 
<< m2 >>
rect 167 8 168 9 
<< m1 >>
rect 19 9 20 10 
<< m1 >>
rect 40 9 41 10 
<< m2 >>
rect 40 9 41 10 
<< m2c >>
rect 40 9 41 10 
<< m1 >>
rect 40 9 41 10 
<< m2 >>
rect 40 9 41 10 
<< m1 >>
rect 42 9 43 10 
<< m2 >>
rect 42 9 43 10 
<< m2c >>
rect 42 9 43 10 
<< m1 >>
rect 42 9 43 10 
<< m2 >>
rect 42 9 43 10 
<< m1 >>
rect 44 9 45 10 
<< m2 >>
rect 44 9 45 10 
<< m2c >>
rect 44 9 45 10 
<< m1 >>
rect 44 9 45 10 
<< m2 >>
rect 44 9 45 10 
<< m1 >>
rect 68 9 69 10 
<< m2 >>
rect 68 9 69 10 
<< m2c >>
rect 68 9 69 10 
<< m1 >>
rect 68 9 69 10 
<< m2 >>
rect 68 9 69 10 
<< m1 >>
rect 69 9 70 10 
<< m1 >>
rect 70 9 71 10 
<< m1 >>
rect 93 9 94 10 
<< m2 >>
rect 93 9 94 10 
<< m2c >>
rect 93 9 94 10 
<< m1 >>
rect 93 9 94 10 
<< m2 >>
rect 93 9 94 10 
<< m1 >>
rect 95 9 96 10 
<< m2 >>
rect 95 9 96 10 
<< m2c >>
rect 95 9 96 10 
<< m1 >>
rect 95 9 96 10 
<< m2 >>
rect 95 9 96 10 
<< m1 >>
rect 124 9 125 10 
<< m1 >>
rect 139 9 140 10 
<< m2 >>
rect 163 9 164 10 
<< m2 >>
rect 165 9 166 10 
<< m2 >>
rect 167 9 168 10 
<< m1 >>
rect 19 10 20 11 
<< m2 >>
rect 20 10 21 11 
<< m1 >>
rect 21 10 22 11 
<< m2 >>
rect 21 10 22 11 
<< m2c >>
rect 21 10 22 11 
<< m1 >>
rect 21 10 22 11 
<< m2 >>
rect 21 10 22 11 
<< m1 >>
rect 22 10 23 11 
<< m1 >>
rect 23 10 24 11 
<< m1 >>
rect 24 10 25 11 
<< m1 >>
rect 25 10 26 11 
<< m1 >>
rect 26 10 27 11 
<< m1 >>
rect 27 10 28 11 
<< m1 >>
rect 28 10 29 11 
<< m1 >>
rect 29 10 30 11 
<< m1 >>
rect 30 10 31 11 
<< m1 >>
rect 31 10 32 11 
<< m1 >>
rect 40 10 41 11 
<< m1 >>
rect 42 10 43 11 
<< m1 >>
rect 44 10 45 11 
<< m1 >>
rect 46 10 47 11 
<< m1 >>
rect 47 10 48 11 
<< m1 >>
rect 48 10 49 11 
<< m1 >>
rect 49 10 50 11 
<< m1 >>
rect 70 10 71 11 
<< m1 >>
rect 93 10 94 11 
<< m1 >>
rect 95 10 96 11 
<< m1 >>
rect 124 10 125 11 
<< m1 >>
rect 139 10 140 11 
<< m1 >>
rect 163 10 164 11 
<< m2 >>
rect 163 10 164 11 
<< m1 >>
rect 164 10 165 11 
<< m1 >>
rect 165 10 166 11 
<< m2 >>
rect 165 10 166 11 
<< m1 >>
rect 166 10 167 11 
<< m1 >>
rect 167 10 168 11 
<< m2 >>
rect 167 10 168 11 
<< m1 >>
rect 168 10 169 11 
<< m1 >>
rect 169 10 170 11 
<< m1 >>
rect 170 10 171 11 
<< m1 >>
rect 171 10 172 11 
<< m1 >>
rect 172 10 173 11 
<< m1 >>
rect 173 10 174 11 
<< m1 >>
rect 174 10 175 11 
<< m1 >>
rect 175 10 176 11 
<< m1 >>
rect 19 11 20 12 
<< m2 >>
rect 20 11 21 12 
<< m1 >>
rect 31 11 32 12 
<< m1 >>
rect 40 11 41 12 
<< m2 >>
rect 40 11 41 12 
<< m2c >>
rect 40 11 41 12 
<< m1 >>
rect 40 11 41 12 
<< m2 >>
rect 40 11 41 12 
<< m2 >>
rect 41 11 42 12 
<< m1 >>
rect 42 11 43 12 
<< m2 >>
rect 42 11 43 12 
<< m2 >>
rect 43 11 44 12 
<< m1 >>
rect 44 11 45 12 
<< m2 >>
rect 44 11 45 12 
<< m2 >>
rect 45 11 46 12 
<< m1 >>
rect 46 11 47 12 
<< m2 >>
rect 46 11 47 12 
<< m2c >>
rect 46 11 47 12 
<< m1 >>
rect 46 11 47 12 
<< m2 >>
rect 46 11 47 12 
<< m1 >>
rect 49 11 50 12 
<< m1 >>
rect 70 11 71 12 
<< m1 >>
rect 93 11 94 12 
<< m2 >>
rect 93 11 94 12 
<< m2c >>
rect 93 11 94 12 
<< m1 >>
rect 93 11 94 12 
<< m2 >>
rect 93 11 94 12 
<< m2 >>
rect 94 11 95 12 
<< m1 >>
rect 95 11 96 12 
<< m2 >>
rect 95 11 96 12 
<< m2 >>
rect 96 11 97 12 
<< m1 >>
rect 97 11 98 12 
<< m2 >>
rect 97 11 98 12 
<< m2c >>
rect 97 11 98 12 
<< m1 >>
rect 97 11 98 12 
<< m2 >>
rect 97 11 98 12 
<< m1 >>
rect 124 11 125 12 
<< m1 >>
rect 139 11 140 12 
<< m1 >>
rect 163 11 164 12 
<< m2 >>
rect 163 11 164 12 
<< m2 >>
rect 165 11 166 12 
<< m2 >>
rect 167 11 168 12 
<< m1 >>
rect 175 11 176 12 
<< pdiffusion >>
rect 12 12 13 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< m1 >>
rect 19 12 20 13 
<< m2 >>
rect 20 12 21 13 
<< pdiffusion >>
rect 30 12 31 13 
<< m1 >>
rect 31 12 32 13 
<< pdiffusion >>
rect 31 12 32 13 
<< pdiffusion >>
rect 32 12 33 13 
<< pdiffusion >>
rect 33 12 34 13 
<< pdiffusion >>
rect 34 12 35 13 
<< pdiffusion >>
rect 35 12 36 13 
<< m1 >>
rect 42 12 43 13 
<< m1 >>
rect 44 12 45 13 
<< pdiffusion >>
rect 48 12 49 13 
<< m1 >>
rect 49 12 50 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< pdiffusion >>
rect 51 12 52 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< pdiffusion >>
rect 66 12 67 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< m1 >>
rect 70 12 71 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< pdiffusion >>
rect 84 12 85 13 
<< pdiffusion >>
rect 85 12 86 13 
<< pdiffusion >>
rect 86 12 87 13 
<< pdiffusion >>
rect 87 12 88 13 
<< pdiffusion >>
rect 88 12 89 13 
<< pdiffusion >>
rect 89 12 90 13 
<< m1 >>
rect 95 12 96 13 
<< m1 >>
rect 97 12 98 13 
<< pdiffusion >>
rect 102 12 103 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< pdiffusion >>
rect 120 12 121 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< m1 >>
rect 124 12 125 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< pdiffusion >>
rect 138 12 139 13 
<< m1 >>
rect 139 12 140 13 
<< pdiffusion >>
rect 139 12 140 13 
<< pdiffusion >>
rect 140 12 141 13 
<< pdiffusion >>
rect 141 12 142 13 
<< pdiffusion >>
rect 142 12 143 13 
<< pdiffusion >>
rect 143 12 144 13 
<< pdiffusion >>
rect 156 12 157 13 
<< pdiffusion >>
rect 157 12 158 13 
<< pdiffusion >>
rect 158 12 159 13 
<< pdiffusion >>
rect 159 12 160 13 
<< pdiffusion >>
rect 160 12 161 13 
<< pdiffusion >>
rect 161 12 162 13 
<< m1 >>
rect 163 12 164 13 
<< m2 >>
rect 163 12 164 13 
<< m1 >>
rect 165 12 166 13 
<< m2 >>
rect 165 12 166 13 
<< m2c >>
rect 165 12 166 13 
<< m1 >>
rect 165 12 166 13 
<< m2 >>
rect 165 12 166 13 
<< m1 >>
rect 167 12 168 13 
<< m2 >>
rect 167 12 168 13 
<< m2c >>
rect 167 12 168 13 
<< m1 >>
rect 167 12 168 13 
<< m2 >>
rect 167 12 168 13 
<< m1 >>
rect 168 12 169 13 
<< m1 >>
rect 169 12 170 13 
<< m1 >>
rect 170 12 171 13 
<< m1 >>
rect 171 12 172 13 
<< pdiffusion >>
rect 174 12 175 13 
<< m1 >>
rect 175 12 176 13 
<< pdiffusion >>
rect 175 12 176 13 
<< pdiffusion >>
rect 176 12 177 13 
<< pdiffusion >>
rect 177 12 178 13 
<< pdiffusion >>
rect 178 12 179 13 
<< pdiffusion >>
rect 179 12 180 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< m1 >>
rect 19 13 20 14 
<< m2 >>
rect 20 13 21 14 
<< pdiffusion >>
rect 30 13 31 14 
<< pdiffusion >>
rect 31 13 32 14 
<< pdiffusion >>
rect 32 13 33 14 
<< pdiffusion >>
rect 33 13 34 14 
<< pdiffusion >>
rect 34 13 35 14 
<< pdiffusion >>
rect 35 13 36 14 
<< m1 >>
rect 42 13 43 14 
<< m1 >>
rect 44 13 45 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< pdiffusion >>
rect 84 13 85 14 
<< pdiffusion >>
rect 85 13 86 14 
<< pdiffusion >>
rect 86 13 87 14 
<< pdiffusion >>
rect 87 13 88 14 
<< pdiffusion >>
rect 88 13 89 14 
<< pdiffusion >>
rect 89 13 90 14 
<< m1 >>
rect 95 13 96 14 
<< m1 >>
rect 97 13 98 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< pdiffusion >>
rect 138 13 139 14 
<< pdiffusion >>
rect 139 13 140 14 
<< pdiffusion >>
rect 140 13 141 14 
<< pdiffusion >>
rect 141 13 142 14 
<< pdiffusion >>
rect 142 13 143 14 
<< pdiffusion >>
rect 143 13 144 14 
<< pdiffusion >>
rect 156 13 157 14 
<< pdiffusion >>
rect 157 13 158 14 
<< pdiffusion >>
rect 158 13 159 14 
<< pdiffusion >>
rect 159 13 160 14 
<< pdiffusion >>
rect 160 13 161 14 
<< pdiffusion >>
rect 161 13 162 14 
<< m1 >>
rect 163 13 164 14 
<< m2 >>
rect 163 13 164 14 
<< m1 >>
rect 165 13 166 14 
<< m1 >>
rect 171 13 172 14 
<< pdiffusion >>
rect 174 13 175 14 
<< pdiffusion >>
rect 175 13 176 14 
<< pdiffusion >>
rect 176 13 177 14 
<< pdiffusion >>
rect 177 13 178 14 
<< pdiffusion >>
rect 178 13 179 14 
<< pdiffusion >>
rect 179 13 180 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< m1 >>
rect 19 14 20 15 
<< m2 >>
rect 20 14 21 15 
<< pdiffusion >>
rect 30 14 31 15 
<< pdiffusion >>
rect 31 14 32 15 
<< pdiffusion >>
rect 32 14 33 15 
<< pdiffusion >>
rect 33 14 34 15 
<< pdiffusion >>
rect 34 14 35 15 
<< pdiffusion >>
rect 35 14 36 15 
<< m1 >>
rect 42 14 43 15 
<< m1 >>
rect 44 14 45 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< pdiffusion >>
rect 84 14 85 15 
<< pdiffusion >>
rect 85 14 86 15 
<< pdiffusion >>
rect 86 14 87 15 
<< pdiffusion >>
rect 87 14 88 15 
<< pdiffusion >>
rect 88 14 89 15 
<< pdiffusion >>
rect 89 14 90 15 
<< m1 >>
rect 95 14 96 15 
<< m1 >>
rect 97 14 98 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< pdiffusion >>
rect 138 14 139 15 
<< pdiffusion >>
rect 139 14 140 15 
<< pdiffusion >>
rect 140 14 141 15 
<< pdiffusion >>
rect 141 14 142 15 
<< pdiffusion >>
rect 142 14 143 15 
<< pdiffusion >>
rect 143 14 144 15 
<< pdiffusion >>
rect 156 14 157 15 
<< pdiffusion >>
rect 157 14 158 15 
<< pdiffusion >>
rect 158 14 159 15 
<< pdiffusion >>
rect 159 14 160 15 
<< pdiffusion >>
rect 160 14 161 15 
<< pdiffusion >>
rect 161 14 162 15 
<< m1 >>
rect 163 14 164 15 
<< m2 >>
rect 163 14 164 15 
<< m1 >>
rect 165 14 166 15 
<< m1 >>
rect 171 14 172 15 
<< pdiffusion >>
rect 174 14 175 15 
<< pdiffusion >>
rect 175 14 176 15 
<< pdiffusion >>
rect 176 14 177 15 
<< pdiffusion >>
rect 177 14 178 15 
<< pdiffusion >>
rect 178 14 179 15 
<< pdiffusion >>
rect 179 14 180 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< m1 >>
rect 19 15 20 16 
<< m2 >>
rect 20 15 21 16 
<< pdiffusion >>
rect 30 15 31 16 
<< pdiffusion >>
rect 31 15 32 16 
<< pdiffusion >>
rect 32 15 33 16 
<< pdiffusion >>
rect 33 15 34 16 
<< pdiffusion >>
rect 34 15 35 16 
<< pdiffusion >>
rect 35 15 36 16 
<< m1 >>
rect 42 15 43 16 
<< m1 >>
rect 44 15 45 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< pdiffusion >>
rect 84 15 85 16 
<< pdiffusion >>
rect 85 15 86 16 
<< pdiffusion >>
rect 86 15 87 16 
<< pdiffusion >>
rect 87 15 88 16 
<< pdiffusion >>
rect 88 15 89 16 
<< pdiffusion >>
rect 89 15 90 16 
<< m1 >>
rect 95 15 96 16 
<< m1 >>
rect 97 15 98 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< pdiffusion >>
rect 138 15 139 16 
<< pdiffusion >>
rect 139 15 140 16 
<< pdiffusion >>
rect 140 15 141 16 
<< pdiffusion >>
rect 141 15 142 16 
<< pdiffusion >>
rect 142 15 143 16 
<< pdiffusion >>
rect 143 15 144 16 
<< pdiffusion >>
rect 156 15 157 16 
<< pdiffusion >>
rect 157 15 158 16 
<< pdiffusion >>
rect 158 15 159 16 
<< pdiffusion >>
rect 159 15 160 16 
<< pdiffusion >>
rect 160 15 161 16 
<< pdiffusion >>
rect 161 15 162 16 
<< m1 >>
rect 163 15 164 16 
<< m2 >>
rect 163 15 164 16 
<< m1 >>
rect 165 15 166 16 
<< m1 >>
rect 171 15 172 16 
<< pdiffusion >>
rect 174 15 175 16 
<< pdiffusion >>
rect 175 15 176 16 
<< pdiffusion >>
rect 176 15 177 16 
<< pdiffusion >>
rect 177 15 178 16 
<< pdiffusion >>
rect 178 15 179 16 
<< pdiffusion >>
rect 179 15 180 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< m1 >>
rect 19 16 20 17 
<< m2 >>
rect 20 16 21 17 
<< pdiffusion >>
rect 30 16 31 17 
<< pdiffusion >>
rect 31 16 32 17 
<< pdiffusion >>
rect 32 16 33 17 
<< pdiffusion >>
rect 33 16 34 17 
<< pdiffusion >>
rect 34 16 35 17 
<< pdiffusion >>
rect 35 16 36 17 
<< m1 >>
rect 42 16 43 17 
<< m1 >>
rect 44 16 45 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< pdiffusion >>
rect 84 16 85 17 
<< pdiffusion >>
rect 85 16 86 17 
<< pdiffusion >>
rect 86 16 87 17 
<< pdiffusion >>
rect 87 16 88 17 
<< pdiffusion >>
rect 88 16 89 17 
<< pdiffusion >>
rect 89 16 90 17 
<< m1 >>
rect 95 16 96 17 
<< m1 >>
rect 97 16 98 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< pdiffusion >>
rect 138 16 139 17 
<< pdiffusion >>
rect 139 16 140 17 
<< pdiffusion >>
rect 140 16 141 17 
<< pdiffusion >>
rect 141 16 142 17 
<< pdiffusion >>
rect 142 16 143 17 
<< pdiffusion >>
rect 143 16 144 17 
<< pdiffusion >>
rect 156 16 157 17 
<< pdiffusion >>
rect 157 16 158 17 
<< pdiffusion >>
rect 158 16 159 17 
<< pdiffusion >>
rect 159 16 160 17 
<< pdiffusion >>
rect 160 16 161 17 
<< pdiffusion >>
rect 161 16 162 17 
<< m1 >>
rect 163 16 164 17 
<< m2 >>
rect 163 16 164 17 
<< m1 >>
rect 165 16 166 17 
<< m1 >>
rect 171 16 172 17 
<< pdiffusion >>
rect 174 16 175 17 
<< pdiffusion >>
rect 175 16 176 17 
<< pdiffusion >>
rect 176 16 177 17 
<< pdiffusion >>
rect 177 16 178 17 
<< pdiffusion >>
rect 178 16 179 17 
<< pdiffusion >>
rect 179 16 180 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< m1 >>
rect 19 17 20 18 
<< m2 >>
rect 20 17 21 18 
<< pdiffusion >>
rect 30 17 31 18 
<< pdiffusion >>
rect 31 17 32 18 
<< pdiffusion >>
rect 32 17 33 18 
<< pdiffusion >>
rect 33 17 34 18 
<< pdiffusion >>
rect 34 17 35 18 
<< pdiffusion >>
rect 35 17 36 18 
<< m1 >>
rect 42 17 43 18 
<< m1 >>
rect 44 17 45 18 
<< pdiffusion >>
rect 48 17 49 18 
<< m1 >>
rect 49 17 50 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< pdiffusion >>
rect 66 17 67 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< m1 >>
rect 70 17 71 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< pdiffusion >>
rect 84 17 85 18 
<< pdiffusion >>
rect 85 17 86 18 
<< pdiffusion >>
rect 86 17 87 18 
<< pdiffusion >>
rect 87 17 88 18 
<< pdiffusion >>
rect 88 17 89 18 
<< pdiffusion >>
rect 89 17 90 18 
<< m1 >>
rect 95 17 96 18 
<< m1 >>
rect 97 17 98 18 
<< pdiffusion >>
rect 102 17 103 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< m1 >>
rect 106 17 107 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< pdiffusion >>
rect 120 17 121 18 
<< m1 >>
rect 121 17 122 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< m1 >>
rect 124 17 125 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< pdiffusion >>
rect 138 17 139 18 
<< pdiffusion >>
rect 139 17 140 18 
<< pdiffusion >>
rect 140 17 141 18 
<< pdiffusion >>
rect 141 17 142 18 
<< pdiffusion >>
rect 142 17 143 18 
<< pdiffusion >>
rect 143 17 144 18 
<< pdiffusion >>
rect 156 17 157 18 
<< pdiffusion >>
rect 157 17 158 18 
<< pdiffusion >>
rect 158 17 159 18 
<< pdiffusion >>
rect 159 17 160 18 
<< pdiffusion >>
rect 160 17 161 18 
<< pdiffusion >>
rect 161 17 162 18 
<< m1 >>
rect 163 17 164 18 
<< m2 >>
rect 163 17 164 18 
<< m1 >>
rect 165 17 166 18 
<< m1 >>
rect 171 17 172 18 
<< pdiffusion >>
rect 174 17 175 18 
<< pdiffusion >>
rect 175 17 176 18 
<< pdiffusion >>
rect 176 17 177 18 
<< pdiffusion >>
rect 177 17 178 18 
<< pdiffusion >>
rect 178 17 179 18 
<< pdiffusion >>
rect 179 17 180 18 
<< m1 >>
rect 19 18 20 19 
<< m2 >>
rect 20 18 21 19 
<< m1 >>
rect 42 18 43 19 
<< m1 >>
rect 44 18 45 19 
<< m1 >>
rect 49 18 50 19 
<< m1 >>
rect 70 18 71 19 
<< m1 >>
rect 95 18 96 19 
<< m1 >>
rect 97 18 98 19 
<< m1 >>
rect 106 18 107 19 
<< m1 >>
rect 121 18 122 19 
<< m1 >>
rect 124 18 125 19 
<< m1 >>
rect 163 18 164 19 
<< m2 >>
rect 163 18 164 19 
<< m1 >>
rect 165 18 166 19 
<< m1 >>
rect 171 18 172 19 
<< m1 >>
rect 17 19 18 20 
<< m2 >>
rect 17 19 18 20 
<< m2c >>
rect 17 19 18 20 
<< m1 >>
rect 17 19 18 20 
<< m2 >>
rect 17 19 18 20 
<< m2 >>
rect 18 19 19 20 
<< m1 >>
rect 19 19 20 20 
<< m2 >>
rect 19 19 20 20 
<< m2 >>
rect 20 19 21 20 
<< m2 >>
rect 41 19 42 20 
<< m1 >>
rect 42 19 43 20 
<< m2 >>
rect 42 19 43 20 
<< m2 >>
rect 43 19 44 20 
<< m1 >>
rect 44 19 45 20 
<< m2 >>
rect 44 19 45 20 
<< m2c >>
rect 44 19 45 20 
<< m1 >>
rect 44 19 45 20 
<< m2 >>
rect 44 19 45 20 
<< m1 >>
rect 49 19 50 20 
<< m1 >>
rect 70 19 71 20 
<< m1 >>
rect 95 19 96 20 
<< m1 >>
rect 97 19 98 20 
<< m1 >>
rect 106 19 107 20 
<< m1 >>
rect 107 19 108 20 
<< m1 >>
rect 108 19 109 20 
<< m1 >>
rect 109 19 110 20 
<< m1 >>
rect 121 19 122 20 
<< m1 >>
rect 124 19 125 20 
<< m1 >>
rect 163 19 164 20 
<< m2 >>
rect 163 19 164 20 
<< m1 >>
rect 165 19 166 20 
<< m1 >>
rect 171 19 172 20 
<< m1 >>
rect 17 20 18 21 
<< m1 >>
rect 19 20 20 21 
<< m2 >>
rect 41 20 42 21 
<< m1 >>
rect 42 20 43 21 
<< m1 >>
rect 49 20 50 21 
<< m1 >>
rect 50 20 51 21 
<< m1 >>
rect 51 20 52 21 
<< m1 >>
rect 52 20 53 21 
<< m1 >>
rect 53 20 54 21 
<< m1 >>
rect 54 20 55 21 
<< m1 >>
rect 55 20 56 21 
<< m1 >>
rect 70 20 71 21 
<< m1 >>
rect 95 20 96 21 
<< m1 >>
rect 97 20 98 21 
<< m1 >>
rect 109 20 110 21 
<< m1 >>
rect 121 20 122 21 
<< m1 >>
rect 124 20 125 21 
<< m1 >>
rect 158 20 159 21 
<< m2 >>
rect 158 20 159 21 
<< m2c >>
rect 158 20 159 21 
<< m1 >>
rect 158 20 159 21 
<< m2 >>
rect 158 20 159 21 
<< m1 >>
rect 159 20 160 21 
<< m1 >>
rect 160 20 161 21 
<< m1 >>
rect 161 20 162 21 
<< m1 >>
rect 162 20 163 21 
<< m1 >>
rect 163 20 164 21 
<< m2 >>
rect 163 20 164 21 
<< m1 >>
rect 165 20 166 21 
<< m2 >>
rect 165 20 166 21 
<< m2c >>
rect 165 20 166 21 
<< m1 >>
rect 165 20 166 21 
<< m2 >>
rect 165 20 166 21 
<< m1 >>
rect 171 20 172 21 
<< m1 >>
rect 17 21 18 22 
<< m1 >>
rect 19 21 20 22 
<< m1 >>
rect 37 21 38 22 
<< m1 >>
rect 38 21 39 22 
<< m1 >>
rect 39 21 40 22 
<< m1 >>
rect 40 21 41 22 
<< m2 >>
rect 40 21 41 22 
<< m2c >>
rect 40 21 41 22 
<< m1 >>
rect 40 21 41 22 
<< m2 >>
rect 40 21 41 22 
<< m2 >>
rect 41 21 42 22 
<< m1 >>
rect 42 21 43 22 
<< m1 >>
rect 44 21 45 22 
<< m1 >>
rect 45 21 46 22 
<< m1 >>
rect 46 21 47 22 
<< m1 >>
rect 47 21 48 22 
<< m2 >>
rect 47 21 48 22 
<< m2c >>
rect 47 21 48 22 
<< m1 >>
rect 47 21 48 22 
<< m2 >>
rect 47 21 48 22 
<< m2 >>
rect 48 21 49 22 
<< m1 >>
rect 55 21 56 22 
<< m1 >>
rect 70 21 71 22 
<< m1 >>
rect 95 21 96 22 
<< m1 >>
rect 97 21 98 22 
<< m1 >>
rect 109 21 110 22 
<< m1 >>
rect 121 21 122 22 
<< m1 >>
rect 124 21 125 22 
<< m2 >>
rect 158 21 159 22 
<< m2 >>
rect 163 21 164 22 
<< m2 >>
rect 165 21 166 22 
<< m2 >>
rect 166 21 167 22 
<< m2 >>
rect 167 21 168 22 
<< m2 >>
rect 168 21 169 22 
<< m2 >>
rect 169 21 170 22 
<< m1 >>
rect 171 21 172 22 
<< m1 >>
rect 13 22 14 23 
<< m1 >>
rect 14 22 15 23 
<< m1 >>
rect 15 22 16 23 
<< m1 >>
rect 16 22 17 23 
<< m1 >>
rect 17 22 18 23 
<< m1 >>
rect 19 22 20 23 
<< m1 >>
rect 37 22 38 23 
<< m1 >>
rect 42 22 43 23 
<< m1 >>
rect 44 22 45 23 
<< m2 >>
rect 48 22 49 23 
<< m1 >>
rect 55 22 56 23 
<< m1 >>
rect 70 22 71 23 
<< m1 >>
rect 95 22 96 23 
<< m1 >>
rect 97 22 98 23 
<< m1 >>
rect 109 22 110 23 
<< m1 >>
rect 121 22 122 23 
<< m1 >>
rect 124 22 125 23 
<< m1 >>
rect 125 22 126 23 
<< m1 >>
rect 126 22 127 23 
<< m1 >>
rect 127 22 128 23 
<< m1 >>
rect 128 22 129 23 
<< m1 >>
rect 129 22 130 23 
<< m1 >>
rect 130 22 131 23 
<< m1 >>
rect 131 22 132 23 
<< m1 >>
rect 132 22 133 23 
<< m1 >>
rect 133 22 134 23 
<< m1 >>
rect 134 22 135 23 
<< m1 >>
rect 135 22 136 23 
<< m1 >>
rect 136 22 137 23 
<< m1 >>
rect 137 22 138 23 
<< m1 >>
rect 138 22 139 23 
<< m1 >>
rect 139 22 140 23 
<< m1 >>
rect 140 22 141 23 
<< m1 >>
rect 141 22 142 23 
<< m1 >>
rect 142 22 143 23 
<< m1 >>
rect 143 22 144 23 
<< m1 >>
rect 144 22 145 23 
<< m1 >>
rect 145 22 146 23 
<< m1 >>
rect 146 22 147 23 
<< m1 >>
rect 147 22 148 23 
<< m1 >>
rect 148 22 149 23 
<< m1 >>
rect 149 22 150 23 
<< m1 >>
rect 150 22 151 23 
<< m1 >>
rect 151 22 152 23 
<< m1 >>
rect 152 22 153 23 
<< m1 >>
rect 153 22 154 23 
<< m1 >>
rect 154 22 155 23 
<< m1 >>
rect 155 22 156 23 
<< m1 >>
rect 156 22 157 23 
<< m1 >>
rect 157 22 158 23 
<< m1 >>
rect 158 22 159 23 
<< m2 >>
rect 158 22 159 23 
<< m1 >>
rect 159 22 160 23 
<< m1 >>
rect 160 22 161 23 
<< m1 >>
rect 161 22 162 23 
<< m1 >>
rect 162 22 163 23 
<< m1 >>
rect 163 22 164 23 
<< m2 >>
rect 163 22 164 23 
<< m1 >>
rect 164 22 165 23 
<< m1 >>
rect 165 22 166 23 
<< m1 >>
rect 166 22 167 23 
<< m1 >>
rect 167 22 168 23 
<< m1 >>
rect 168 22 169 23 
<< m1 >>
rect 169 22 170 23 
<< m2 >>
rect 169 22 170 23 
<< m1 >>
rect 171 22 172 23 
<< m1 >>
rect 13 23 14 24 
<< m1 >>
rect 19 23 20 24 
<< m1 >>
rect 37 23 38 24 
<< m2 >>
rect 37 23 38 24 
<< m2c >>
rect 37 23 38 24 
<< m1 >>
rect 37 23 38 24 
<< m2 >>
rect 37 23 38 24 
<< m1 >>
rect 42 23 43 24 
<< m2 >>
rect 42 23 43 24 
<< m2c >>
rect 42 23 43 24 
<< m1 >>
rect 42 23 43 24 
<< m2 >>
rect 42 23 43 24 
<< m1 >>
rect 44 23 45 24 
<< m2 >>
rect 44 23 45 24 
<< m2c >>
rect 44 23 45 24 
<< m1 >>
rect 44 23 45 24 
<< m2 >>
rect 44 23 45 24 
<< m1 >>
rect 46 23 47 24 
<< m2 >>
rect 46 23 47 24 
<< m2c >>
rect 46 23 47 24 
<< m1 >>
rect 46 23 47 24 
<< m2 >>
rect 46 23 47 24 
<< m1 >>
rect 47 23 48 24 
<< m1 >>
rect 48 23 49 24 
<< m2 >>
rect 48 23 49 24 
<< m1 >>
rect 49 23 50 24 
<< m1 >>
rect 50 23 51 24 
<< m1 >>
rect 51 23 52 24 
<< m1 >>
rect 52 23 53 24 
<< m1 >>
rect 53 23 54 24 
<< m2 >>
rect 53 23 54 24 
<< m2c >>
rect 53 23 54 24 
<< m1 >>
rect 53 23 54 24 
<< m2 >>
rect 53 23 54 24 
<< m2 >>
rect 54 23 55 24 
<< m1 >>
rect 55 23 56 24 
<< m2 >>
rect 55 23 56 24 
<< m2 >>
rect 56 23 57 24 
<< m1 >>
rect 57 23 58 24 
<< m2 >>
rect 57 23 58 24 
<< m2c >>
rect 57 23 58 24 
<< m1 >>
rect 57 23 58 24 
<< m2 >>
rect 57 23 58 24 
<< m1 >>
rect 58 23 59 24 
<< m1 >>
rect 59 23 60 24 
<< m1 >>
rect 60 23 61 24 
<< m1 >>
rect 61 23 62 24 
<< m1 >>
rect 62 23 63 24 
<< m1 >>
rect 63 23 64 24 
<< m1 >>
rect 64 23 65 24 
<< m1 >>
rect 65 23 66 24 
<< m1 >>
rect 66 23 67 24 
<< m1 >>
rect 67 23 68 24 
<< m1 >>
rect 68 23 69 24 
<< m2 >>
rect 68 23 69 24 
<< m2c >>
rect 68 23 69 24 
<< m1 >>
rect 68 23 69 24 
<< m2 >>
rect 68 23 69 24 
<< m2 >>
rect 69 23 70 24 
<< m1 >>
rect 70 23 71 24 
<< m2 >>
rect 70 23 71 24 
<< m2 >>
rect 71 23 72 24 
<< m1 >>
rect 72 23 73 24 
<< m2 >>
rect 72 23 73 24 
<< m2c >>
rect 72 23 73 24 
<< m1 >>
rect 72 23 73 24 
<< m2 >>
rect 72 23 73 24 
<< m1 >>
rect 73 23 74 24 
<< m1 >>
rect 74 23 75 24 
<< m1 >>
rect 75 23 76 24 
<< m1 >>
rect 76 23 77 24 
<< m1 >>
rect 77 23 78 24 
<< m1 >>
rect 78 23 79 24 
<< m1 >>
rect 79 23 80 24 
<< m1 >>
rect 80 23 81 24 
<< m1 >>
rect 81 23 82 24 
<< m1 >>
rect 82 23 83 24 
<< m1 >>
rect 83 23 84 24 
<< m1 >>
rect 84 23 85 24 
<< m1 >>
rect 85 23 86 24 
<< m1 >>
rect 86 23 87 24 
<< m1 >>
rect 87 23 88 24 
<< m1 >>
rect 88 23 89 24 
<< m1 >>
rect 89 23 90 24 
<< m1 >>
rect 90 23 91 24 
<< m1 >>
rect 91 23 92 24 
<< m1 >>
rect 95 23 96 24 
<< m1 >>
rect 97 23 98 24 
<< m1 >>
rect 109 23 110 24 
<< m2 >>
rect 120 23 121 24 
<< m1 >>
rect 121 23 122 24 
<< m2 >>
rect 121 23 122 24 
<< m2 >>
rect 122 23 123 24 
<< m2 >>
rect 123 23 124 24 
<< m2 >>
rect 124 23 125 24 
<< m2 >>
rect 125 23 126 24 
<< m2 >>
rect 126 23 127 24 
<< m2 >>
rect 127 23 128 24 
<< m2 >>
rect 128 23 129 24 
<< m2 >>
rect 129 23 130 24 
<< m2 >>
rect 130 23 131 24 
<< m2 >>
rect 131 23 132 24 
<< m2 >>
rect 132 23 133 24 
<< m2 >>
rect 133 23 134 24 
<< m2 >>
rect 134 23 135 24 
<< m2 >>
rect 135 23 136 24 
<< m2 >>
rect 136 23 137 24 
<< m2 >>
rect 137 23 138 24 
<< m2 >>
rect 138 23 139 24 
<< m2 >>
rect 139 23 140 24 
<< m2 >>
rect 140 23 141 24 
<< m2 >>
rect 141 23 142 24 
<< m2 >>
rect 142 23 143 24 
<< m2 >>
rect 143 23 144 24 
<< m2 >>
rect 144 23 145 24 
<< m2 >>
rect 145 23 146 24 
<< m2 >>
rect 146 23 147 24 
<< m2 >>
rect 147 23 148 24 
<< m2 >>
rect 148 23 149 24 
<< m2 >>
rect 149 23 150 24 
<< m2 >>
rect 150 23 151 24 
<< m2 >>
rect 151 23 152 24 
<< m2 >>
rect 152 23 153 24 
<< m2 >>
rect 153 23 154 24 
<< m2 >>
rect 154 23 155 24 
<< m2 >>
rect 155 23 156 24 
<< m2 >>
rect 156 23 157 24 
<< m2 >>
rect 157 23 158 24 
<< m2 >>
rect 158 23 159 24 
<< m2 >>
rect 163 23 164 24 
<< m1 >>
rect 169 23 170 24 
<< m2 >>
rect 169 23 170 24 
<< m1 >>
rect 171 23 172 24 
<< m1 >>
rect 13 24 14 25 
<< m1 >>
rect 19 24 20 25 
<< m2 >>
rect 37 24 38 25 
<< m2 >>
rect 42 24 43 25 
<< m2 >>
rect 44 24 45 25 
<< m2 >>
rect 46 24 47 25 
<< m2 >>
rect 48 24 49 25 
<< m1 >>
rect 55 24 56 25 
<< m1 >>
rect 70 24 71 25 
<< m1 >>
rect 91 24 92 25 
<< m1 >>
rect 95 24 96 25 
<< m1 >>
rect 97 24 98 25 
<< m1 >>
rect 109 24 110 25 
<< m2 >>
rect 120 24 121 25 
<< m1 >>
rect 121 24 122 25 
<< m1 >>
rect 163 24 164 25 
<< m2 >>
rect 163 24 164 25 
<< m2c >>
rect 163 24 164 25 
<< m1 >>
rect 163 24 164 25 
<< m2 >>
rect 163 24 164 25 
<< m1 >>
rect 169 24 170 25 
<< m2 >>
rect 169 24 170 25 
<< m1 >>
rect 171 24 172 25 
<< m1 >>
rect 13 25 14 26 
<< m1 >>
rect 19 25 20 26 
<< m1 >>
rect 37 25 38 26 
<< m2 >>
rect 37 25 38 26 
<< m1 >>
rect 38 25 39 26 
<< m1 >>
rect 39 25 40 26 
<< m1 >>
rect 40 25 41 26 
<< m1 >>
rect 41 25 42 26 
<< m1 >>
rect 42 25 43 26 
<< m2 >>
rect 42 25 43 26 
<< m1 >>
rect 43 25 44 26 
<< m1 >>
rect 44 25 45 26 
<< m2 >>
rect 44 25 45 26 
<< m1 >>
rect 45 25 46 26 
<< m1 >>
rect 46 25 47 26 
<< m2 >>
rect 46 25 47 26 
<< m1 >>
rect 47 25 48 26 
<< m1 >>
rect 48 25 49 26 
<< m2 >>
rect 48 25 49 26 
<< m1 >>
rect 49 25 50 26 
<< m1 >>
rect 50 25 51 26 
<< m1 >>
rect 51 25 52 26 
<< m1 >>
rect 52 25 53 26 
<< m1 >>
rect 53 25 54 26 
<< m2 >>
rect 53 25 54 26 
<< m2c >>
rect 53 25 54 26 
<< m1 >>
rect 53 25 54 26 
<< m2 >>
rect 53 25 54 26 
<< m2 >>
rect 54 25 55 26 
<< m1 >>
rect 55 25 56 26 
<< m2 >>
rect 55 25 56 26 
<< m2 >>
rect 56 25 57 26 
<< m1 >>
rect 57 25 58 26 
<< m2 >>
rect 57 25 58 26 
<< m2c >>
rect 57 25 58 26 
<< m1 >>
rect 57 25 58 26 
<< m2 >>
rect 57 25 58 26 
<< m1 >>
rect 58 25 59 26 
<< m1 >>
rect 59 25 60 26 
<< m1 >>
rect 60 25 61 26 
<< m1 >>
rect 61 25 62 26 
<< m1 >>
rect 62 25 63 26 
<< m1 >>
rect 63 25 64 26 
<< m1 >>
rect 64 25 65 26 
<< m1 >>
rect 65 25 66 26 
<< m1 >>
rect 66 25 67 26 
<< m1 >>
rect 67 25 68 26 
<< m1 >>
rect 68 25 69 26 
<< m2 >>
rect 68 25 69 26 
<< m2c >>
rect 68 25 69 26 
<< m1 >>
rect 68 25 69 26 
<< m2 >>
rect 68 25 69 26 
<< m2 >>
rect 69 25 70 26 
<< m1 >>
rect 70 25 71 26 
<< m1 >>
rect 91 25 92 26 
<< m1 >>
rect 95 25 96 26 
<< m1 >>
rect 97 25 98 26 
<< m1 >>
rect 109 25 110 26 
<< m2 >>
rect 120 25 121 26 
<< m1 >>
rect 121 25 122 26 
<< m1 >>
rect 122 25 123 26 
<< m1 >>
rect 123 25 124 26 
<< m1 >>
rect 124 25 125 26 
<< m1 >>
rect 125 25 126 26 
<< m1 >>
rect 126 25 127 26 
<< m1 >>
rect 127 25 128 26 
<< m1 >>
rect 128 25 129 26 
<< m1 >>
rect 129 25 130 26 
<< m1 >>
rect 130 25 131 26 
<< m1 >>
rect 131 25 132 26 
<< m1 >>
rect 132 25 133 26 
<< m1 >>
rect 133 25 134 26 
<< m1 >>
rect 134 25 135 26 
<< m1 >>
rect 135 25 136 26 
<< m1 >>
rect 136 25 137 26 
<< m1 >>
rect 137 25 138 26 
<< m1 >>
rect 138 25 139 26 
<< m1 >>
rect 139 25 140 26 
<< m1 >>
rect 140 25 141 26 
<< m1 >>
rect 141 25 142 26 
<< m1 >>
rect 142 25 143 26 
<< m1 >>
rect 143 25 144 26 
<< m1 >>
rect 144 25 145 26 
<< m1 >>
rect 145 25 146 26 
<< m1 >>
rect 146 25 147 26 
<< m1 >>
rect 147 25 148 26 
<< m1 >>
rect 148 25 149 26 
<< m1 >>
rect 149 25 150 26 
<< m1 >>
rect 150 25 151 26 
<< m1 >>
rect 151 25 152 26 
<< m1 >>
rect 152 25 153 26 
<< m1 >>
rect 153 25 154 26 
<< m1 >>
rect 154 25 155 26 
<< m1 >>
rect 163 25 164 26 
<< m1 >>
rect 169 25 170 26 
<< m2 >>
rect 169 25 170 26 
<< m1 >>
rect 171 25 172 26 
<< m1 >>
rect 13 26 14 27 
<< m1 >>
rect 19 26 20 27 
<< m1 >>
rect 37 26 38 27 
<< m2 >>
rect 37 26 38 27 
<< m2 >>
rect 42 26 43 27 
<< m2 >>
rect 44 26 45 27 
<< m2 >>
rect 46 26 47 27 
<< m2 >>
rect 48 26 49 27 
<< m1 >>
rect 55 26 56 27 
<< m2 >>
rect 69 26 70 27 
<< m1 >>
rect 70 26 71 27 
<< m2 >>
rect 70 26 71 27 
<< m2 >>
rect 71 26 72 27 
<< m2 >>
rect 72 26 73 27 
<< m2 >>
rect 73 26 74 27 
<< m1 >>
rect 91 26 92 27 
<< m1 >>
rect 95 26 96 27 
<< m1 >>
rect 97 26 98 27 
<< m1 >>
rect 109 26 110 27 
<< m2 >>
rect 120 26 121 27 
<< m1 >>
rect 154 26 155 27 
<< m1 >>
rect 163 26 164 27 
<< m1 >>
rect 169 26 170 27 
<< m2 >>
rect 169 26 170 27 
<< m1 >>
rect 171 26 172 27 
<< m1 >>
rect 13 27 14 28 
<< m1 >>
rect 19 27 20 28 
<< m1 >>
rect 37 27 38 28 
<< m2 >>
rect 37 27 38 28 
<< m1 >>
rect 42 27 43 28 
<< m2 >>
rect 42 27 43 28 
<< m2c >>
rect 42 27 43 28 
<< m1 >>
rect 42 27 43 28 
<< m2 >>
rect 42 27 43 28 
<< m1 >>
rect 44 27 45 28 
<< m2 >>
rect 44 27 45 28 
<< m2c >>
rect 44 27 45 28 
<< m1 >>
rect 44 27 45 28 
<< m2 >>
rect 44 27 45 28 
<< m1 >>
rect 46 27 47 28 
<< m2 >>
rect 46 27 47 28 
<< m2c >>
rect 46 27 47 28 
<< m1 >>
rect 46 27 47 28 
<< m2 >>
rect 46 27 47 28 
<< m1 >>
rect 48 27 49 28 
<< m2 >>
rect 48 27 49 28 
<< m2c >>
rect 48 27 49 28 
<< m1 >>
rect 48 27 49 28 
<< m2 >>
rect 48 27 49 28 
<< m1 >>
rect 49 27 50 28 
<< m1 >>
rect 55 27 56 28 
<< m1 >>
rect 70 27 71 28 
<< m1 >>
rect 71 27 72 28 
<< m1 >>
rect 72 27 73 28 
<< m1 >>
rect 73 27 74 28 
<< m2 >>
rect 73 27 74 28 
<< m1 >>
rect 74 27 75 28 
<< m1 >>
rect 75 27 76 28 
<< m1 >>
rect 76 27 77 28 
<< m1 >>
rect 77 27 78 28 
<< m1 >>
rect 78 27 79 28 
<< m1 >>
rect 79 27 80 28 
<< m1 >>
rect 80 27 81 28 
<< m1 >>
rect 81 27 82 28 
<< m1 >>
rect 82 27 83 28 
<< m1 >>
rect 85 27 86 28 
<< m1 >>
rect 86 27 87 28 
<< m1 >>
rect 87 27 88 28 
<< m1 >>
rect 88 27 89 28 
<< m1 >>
rect 89 27 90 28 
<< m1 >>
rect 91 27 92 28 
<< m1 >>
rect 95 27 96 28 
<< m1 >>
rect 97 27 98 28 
<< m1 >>
rect 109 27 110 28 
<< m1 >>
rect 120 27 121 28 
<< m2 >>
rect 120 27 121 28 
<< m2c >>
rect 120 27 121 28 
<< m1 >>
rect 120 27 121 28 
<< m2 >>
rect 120 27 121 28 
<< m1 >>
rect 154 27 155 28 
<< m1 >>
rect 163 27 164 28 
<< m1 >>
rect 169 27 170 28 
<< m2 >>
rect 169 27 170 28 
<< m1 >>
rect 171 27 172 28 
<< m1 >>
rect 13 28 14 29 
<< m1 >>
rect 19 28 20 29 
<< m1 >>
rect 37 28 38 29 
<< m2 >>
rect 37 28 38 29 
<< m1 >>
rect 42 28 43 29 
<< m1 >>
rect 44 28 45 29 
<< m1 >>
rect 46 28 47 29 
<< m1 >>
rect 49 28 50 29 
<< m1 >>
rect 52 28 53 29 
<< m1 >>
rect 53 28 54 29 
<< m2 >>
rect 53 28 54 29 
<< m2c >>
rect 53 28 54 29 
<< m1 >>
rect 53 28 54 29 
<< m2 >>
rect 53 28 54 29 
<< m2 >>
rect 54 28 55 29 
<< m1 >>
rect 55 28 56 29 
<< m2 >>
rect 55 28 56 29 
<< m2 >>
rect 56 28 57 29 
<< m1 >>
rect 64 28 65 29 
<< m1 >>
rect 65 28 66 29 
<< m1 >>
rect 66 28 67 29 
<< m1 >>
rect 67 28 68 29 
<< m2 >>
rect 73 28 74 29 
<< m1 >>
rect 82 28 83 29 
<< m1 >>
rect 85 28 86 29 
<< m1 >>
rect 89 28 90 29 
<< m2 >>
rect 89 28 90 29 
<< m2c >>
rect 89 28 90 29 
<< m1 >>
rect 89 28 90 29 
<< m2 >>
rect 89 28 90 29 
<< m2 >>
rect 90 28 91 29 
<< m1 >>
rect 91 28 92 29 
<< m2 >>
rect 91 28 92 29 
<< m2 >>
rect 92 28 93 29 
<< m1 >>
rect 95 28 96 29 
<< m1 >>
rect 97 28 98 29 
<< m1 >>
rect 109 28 110 29 
<< m1 >>
rect 111 28 112 29 
<< m1 >>
rect 112 28 113 29 
<< m1 >>
rect 113 28 114 29 
<< m1 >>
rect 114 28 115 29 
<< m1 >>
rect 115 28 116 29 
<< m1 >>
rect 116 28 117 29 
<< m1 >>
rect 117 28 118 29 
<< m1 >>
rect 118 28 119 29 
<< m1 >>
rect 119 28 120 29 
<< m1 >>
rect 120 28 121 29 
<< m1 >>
rect 124 28 125 29 
<< m1 >>
rect 125 28 126 29 
<< m1 >>
rect 126 28 127 29 
<< m1 >>
rect 127 28 128 29 
<< m1 >>
rect 154 28 155 29 
<< m1 >>
rect 163 28 164 29 
<< m1 >>
rect 169 28 170 29 
<< m2 >>
rect 169 28 170 29 
<< m1 >>
rect 171 28 172 29 
<< m1 >>
rect 13 29 14 30 
<< m1 >>
rect 19 29 20 30 
<< m1 >>
rect 37 29 38 30 
<< m2 >>
rect 37 29 38 30 
<< m1 >>
rect 42 29 43 30 
<< m1 >>
rect 44 29 45 30 
<< m1 >>
rect 46 29 47 30 
<< m1 >>
rect 49 29 50 30 
<< m1 >>
rect 52 29 53 30 
<< m1 >>
rect 55 29 56 30 
<< m2 >>
rect 56 29 57 30 
<< m1 >>
rect 64 29 65 30 
<< m1 >>
rect 67 29 68 30 
<< m1 >>
rect 73 29 74 30 
<< m2 >>
rect 73 29 74 30 
<< m2c >>
rect 73 29 74 30 
<< m1 >>
rect 73 29 74 30 
<< m2 >>
rect 73 29 74 30 
<< m1 >>
rect 82 29 83 30 
<< m1 >>
rect 85 29 86 30 
<< m1 >>
rect 91 29 92 30 
<< m2 >>
rect 92 29 93 30 
<< m1 >>
rect 95 29 96 30 
<< m1 >>
rect 97 29 98 30 
<< m1 >>
rect 109 29 110 30 
<< m1 >>
rect 111 29 112 30 
<< m1 >>
rect 124 29 125 30 
<< m1 >>
rect 127 29 128 30 
<< m1 >>
rect 154 29 155 30 
<< m1 >>
rect 163 29 164 30 
<< m1 >>
rect 169 29 170 30 
<< m2 >>
rect 169 29 170 30 
<< m1 >>
rect 171 29 172 30 
<< pdiffusion >>
rect 12 30 13 31 
<< m1 >>
rect 13 30 14 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< pdiffusion >>
rect 15 30 16 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< m1 >>
rect 19 30 20 31 
<< m1 >>
rect 37 30 38 31 
<< m2 >>
rect 37 30 38 31 
<< m1 >>
rect 42 30 43 31 
<< m1 >>
rect 44 30 45 31 
<< m1 >>
rect 46 30 47 31 
<< pdiffusion >>
rect 48 30 49 31 
<< m1 >>
rect 49 30 50 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< m1 >>
rect 52 30 53 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 55 30 56 31 
<< m2 >>
rect 56 30 57 31 
<< m1 >>
rect 64 30 65 31 
<< pdiffusion >>
rect 66 30 67 31 
<< m1 >>
rect 67 30 68 31 
<< pdiffusion >>
rect 67 30 68 31 
<< pdiffusion >>
rect 68 30 69 31 
<< pdiffusion >>
rect 69 30 70 31 
<< pdiffusion >>
rect 70 30 71 31 
<< pdiffusion >>
rect 71 30 72 31 
<< m1 >>
rect 73 30 74 31 
<< m1 >>
rect 82 30 83 31 
<< pdiffusion >>
rect 84 30 85 31 
<< m1 >>
rect 85 30 86 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< m1 >>
rect 91 30 92 31 
<< m2 >>
rect 92 30 93 31 
<< m1 >>
rect 95 30 96 31 
<< m1 >>
rect 97 30 98 31 
<< pdiffusion >>
rect 102 30 103 31 
<< pdiffusion >>
rect 103 30 104 31 
<< pdiffusion >>
rect 104 30 105 31 
<< pdiffusion >>
rect 105 30 106 31 
<< pdiffusion >>
rect 106 30 107 31 
<< pdiffusion >>
rect 107 30 108 31 
<< m1 >>
rect 109 30 110 31 
<< m1 >>
rect 111 30 112 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< m1 >>
rect 124 30 125 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< m1 >>
rect 127 30 128 31 
<< pdiffusion >>
rect 138 30 139 31 
<< pdiffusion >>
rect 139 30 140 31 
<< pdiffusion >>
rect 140 30 141 31 
<< pdiffusion >>
rect 141 30 142 31 
<< pdiffusion >>
rect 142 30 143 31 
<< pdiffusion >>
rect 143 30 144 31 
<< m1 >>
rect 154 30 155 31 
<< pdiffusion >>
rect 156 30 157 31 
<< pdiffusion >>
rect 157 30 158 31 
<< pdiffusion >>
rect 158 30 159 31 
<< pdiffusion >>
rect 159 30 160 31 
<< pdiffusion >>
rect 160 30 161 31 
<< pdiffusion >>
rect 161 30 162 31 
<< m1 >>
rect 163 30 164 31 
<< m1 >>
rect 169 30 170 31 
<< m2 >>
rect 169 30 170 31 
<< m1 >>
rect 171 30 172 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< m1 >>
rect 19 31 20 32 
<< m1 >>
rect 37 31 38 32 
<< m2 >>
rect 37 31 38 32 
<< m1 >>
rect 42 31 43 32 
<< m1 >>
rect 44 31 45 32 
<< m1 >>
rect 46 31 47 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 55 31 56 32 
<< m2 >>
rect 56 31 57 32 
<< m1 >>
rect 64 31 65 32 
<< pdiffusion >>
rect 66 31 67 32 
<< pdiffusion >>
rect 67 31 68 32 
<< pdiffusion >>
rect 68 31 69 32 
<< pdiffusion >>
rect 69 31 70 32 
<< pdiffusion >>
rect 70 31 71 32 
<< pdiffusion >>
rect 71 31 72 32 
<< m1 >>
rect 73 31 74 32 
<< m1 >>
rect 82 31 83 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< m1 >>
rect 91 31 92 32 
<< m2 >>
rect 92 31 93 32 
<< m1 >>
rect 95 31 96 32 
<< m1 >>
rect 97 31 98 32 
<< pdiffusion >>
rect 102 31 103 32 
<< pdiffusion >>
rect 103 31 104 32 
<< pdiffusion >>
rect 104 31 105 32 
<< pdiffusion >>
rect 105 31 106 32 
<< pdiffusion >>
rect 106 31 107 32 
<< pdiffusion >>
rect 107 31 108 32 
<< m1 >>
rect 109 31 110 32 
<< m1 >>
rect 111 31 112 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< m1 >>
rect 127 31 128 32 
<< pdiffusion >>
rect 138 31 139 32 
<< pdiffusion >>
rect 139 31 140 32 
<< pdiffusion >>
rect 140 31 141 32 
<< pdiffusion >>
rect 141 31 142 32 
<< pdiffusion >>
rect 142 31 143 32 
<< pdiffusion >>
rect 143 31 144 32 
<< m1 >>
rect 154 31 155 32 
<< pdiffusion >>
rect 156 31 157 32 
<< pdiffusion >>
rect 157 31 158 32 
<< pdiffusion >>
rect 158 31 159 32 
<< pdiffusion >>
rect 159 31 160 32 
<< pdiffusion >>
rect 160 31 161 32 
<< pdiffusion >>
rect 161 31 162 32 
<< m1 >>
rect 163 31 164 32 
<< m1 >>
rect 169 31 170 32 
<< m2 >>
rect 169 31 170 32 
<< m1 >>
rect 171 31 172 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< m1 >>
rect 19 32 20 33 
<< m1 >>
rect 37 32 38 33 
<< m2 >>
rect 37 32 38 33 
<< m1 >>
rect 42 32 43 33 
<< m1 >>
rect 44 32 45 33 
<< m1 >>
rect 46 32 47 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 55 32 56 33 
<< m2 >>
rect 56 32 57 33 
<< m1 >>
rect 64 32 65 33 
<< pdiffusion >>
rect 66 32 67 33 
<< pdiffusion >>
rect 67 32 68 33 
<< pdiffusion >>
rect 68 32 69 33 
<< pdiffusion >>
rect 69 32 70 33 
<< pdiffusion >>
rect 70 32 71 33 
<< pdiffusion >>
rect 71 32 72 33 
<< m1 >>
rect 73 32 74 33 
<< m1 >>
rect 82 32 83 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< m1 >>
rect 91 32 92 33 
<< m2 >>
rect 92 32 93 33 
<< m1 >>
rect 95 32 96 33 
<< m1 >>
rect 97 32 98 33 
<< pdiffusion >>
rect 102 32 103 33 
<< pdiffusion >>
rect 103 32 104 33 
<< pdiffusion >>
rect 104 32 105 33 
<< pdiffusion >>
rect 105 32 106 33 
<< pdiffusion >>
rect 106 32 107 33 
<< pdiffusion >>
rect 107 32 108 33 
<< m1 >>
rect 109 32 110 33 
<< m1 >>
rect 111 32 112 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< m1 >>
rect 127 32 128 33 
<< pdiffusion >>
rect 138 32 139 33 
<< pdiffusion >>
rect 139 32 140 33 
<< pdiffusion >>
rect 140 32 141 33 
<< pdiffusion >>
rect 141 32 142 33 
<< pdiffusion >>
rect 142 32 143 33 
<< pdiffusion >>
rect 143 32 144 33 
<< m1 >>
rect 154 32 155 33 
<< pdiffusion >>
rect 156 32 157 33 
<< pdiffusion >>
rect 157 32 158 33 
<< pdiffusion >>
rect 158 32 159 33 
<< pdiffusion >>
rect 159 32 160 33 
<< pdiffusion >>
rect 160 32 161 33 
<< pdiffusion >>
rect 161 32 162 33 
<< m1 >>
rect 163 32 164 33 
<< m1 >>
rect 169 32 170 33 
<< m2 >>
rect 169 32 170 33 
<< m1 >>
rect 171 32 172 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< m1 >>
rect 19 33 20 34 
<< m1 >>
rect 37 33 38 34 
<< m2 >>
rect 37 33 38 34 
<< m1 >>
rect 42 33 43 34 
<< m1 >>
rect 44 33 45 34 
<< m1 >>
rect 46 33 47 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 55 33 56 34 
<< m2 >>
rect 56 33 57 34 
<< m1 >>
rect 64 33 65 34 
<< pdiffusion >>
rect 66 33 67 34 
<< pdiffusion >>
rect 67 33 68 34 
<< pdiffusion >>
rect 68 33 69 34 
<< pdiffusion >>
rect 69 33 70 34 
<< pdiffusion >>
rect 70 33 71 34 
<< pdiffusion >>
rect 71 33 72 34 
<< m1 >>
rect 73 33 74 34 
<< m1 >>
rect 82 33 83 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< m1 >>
rect 91 33 92 34 
<< m2 >>
rect 92 33 93 34 
<< m1 >>
rect 95 33 96 34 
<< m1 >>
rect 97 33 98 34 
<< pdiffusion >>
rect 102 33 103 34 
<< pdiffusion >>
rect 103 33 104 34 
<< pdiffusion >>
rect 104 33 105 34 
<< pdiffusion >>
rect 105 33 106 34 
<< pdiffusion >>
rect 106 33 107 34 
<< pdiffusion >>
rect 107 33 108 34 
<< m1 >>
rect 109 33 110 34 
<< m1 >>
rect 111 33 112 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< m1 >>
rect 127 33 128 34 
<< pdiffusion >>
rect 138 33 139 34 
<< pdiffusion >>
rect 139 33 140 34 
<< pdiffusion >>
rect 140 33 141 34 
<< pdiffusion >>
rect 141 33 142 34 
<< pdiffusion >>
rect 142 33 143 34 
<< pdiffusion >>
rect 143 33 144 34 
<< m1 >>
rect 154 33 155 34 
<< pdiffusion >>
rect 156 33 157 34 
<< pdiffusion >>
rect 157 33 158 34 
<< pdiffusion >>
rect 158 33 159 34 
<< pdiffusion >>
rect 159 33 160 34 
<< pdiffusion >>
rect 160 33 161 34 
<< pdiffusion >>
rect 161 33 162 34 
<< m1 >>
rect 163 33 164 34 
<< m1 >>
rect 169 33 170 34 
<< m2 >>
rect 169 33 170 34 
<< m1 >>
rect 171 33 172 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< m1 >>
rect 19 34 20 35 
<< m1 >>
rect 37 34 38 35 
<< m2 >>
rect 37 34 38 35 
<< m1 >>
rect 42 34 43 35 
<< m1 >>
rect 44 34 45 35 
<< m1 >>
rect 46 34 47 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 55 34 56 35 
<< m2 >>
rect 56 34 57 35 
<< m1 >>
rect 64 34 65 35 
<< pdiffusion >>
rect 66 34 67 35 
<< pdiffusion >>
rect 67 34 68 35 
<< pdiffusion >>
rect 68 34 69 35 
<< pdiffusion >>
rect 69 34 70 35 
<< pdiffusion >>
rect 70 34 71 35 
<< pdiffusion >>
rect 71 34 72 35 
<< m1 >>
rect 73 34 74 35 
<< m1 >>
rect 82 34 83 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< m1 >>
rect 91 34 92 35 
<< m2 >>
rect 92 34 93 35 
<< m1 >>
rect 95 34 96 35 
<< m2 >>
rect 95 34 96 35 
<< m2c >>
rect 95 34 96 35 
<< m1 >>
rect 95 34 96 35 
<< m2 >>
rect 95 34 96 35 
<< m1 >>
rect 97 34 98 35 
<< m2 >>
rect 97 34 98 35 
<< m2c >>
rect 97 34 98 35 
<< m1 >>
rect 97 34 98 35 
<< m2 >>
rect 97 34 98 35 
<< pdiffusion >>
rect 102 34 103 35 
<< pdiffusion >>
rect 103 34 104 35 
<< pdiffusion >>
rect 104 34 105 35 
<< pdiffusion >>
rect 105 34 106 35 
<< pdiffusion >>
rect 106 34 107 35 
<< pdiffusion >>
rect 107 34 108 35 
<< m1 >>
rect 109 34 110 35 
<< m1 >>
rect 111 34 112 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< m1 >>
rect 127 34 128 35 
<< pdiffusion >>
rect 138 34 139 35 
<< pdiffusion >>
rect 139 34 140 35 
<< pdiffusion >>
rect 140 34 141 35 
<< pdiffusion >>
rect 141 34 142 35 
<< pdiffusion >>
rect 142 34 143 35 
<< pdiffusion >>
rect 143 34 144 35 
<< m1 >>
rect 154 34 155 35 
<< pdiffusion >>
rect 156 34 157 35 
<< pdiffusion >>
rect 157 34 158 35 
<< pdiffusion >>
rect 158 34 159 35 
<< pdiffusion >>
rect 159 34 160 35 
<< pdiffusion >>
rect 160 34 161 35 
<< pdiffusion >>
rect 161 34 162 35 
<< m1 >>
rect 163 34 164 35 
<< m1 >>
rect 169 34 170 35 
<< m2 >>
rect 169 34 170 35 
<< m1 >>
rect 171 34 172 35 
<< pdiffusion >>
rect 12 35 13 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< m1 >>
rect 19 35 20 36 
<< m1 >>
rect 37 35 38 36 
<< m2 >>
rect 37 35 38 36 
<< m1 >>
rect 42 35 43 36 
<< m1 >>
rect 44 35 45 36 
<< m1 >>
rect 46 35 47 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 55 35 56 36 
<< m2 >>
rect 56 35 57 36 
<< m1 >>
rect 64 35 65 36 
<< pdiffusion >>
rect 66 35 67 36 
<< pdiffusion >>
rect 67 35 68 36 
<< pdiffusion >>
rect 68 35 69 36 
<< pdiffusion >>
rect 69 35 70 36 
<< pdiffusion >>
rect 70 35 71 36 
<< pdiffusion >>
rect 71 35 72 36 
<< m1 >>
rect 73 35 74 36 
<< m1 >>
rect 82 35 83 36 
<< pdiffusion >>
rect 84 35 85 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< m1 >>
rect 91 35 92 36 
<< m2 >>
rect 92 35 93 36 
<< m2 >>
rect 95 35 96 36 
<< m2 >>
rect 97 35 98 36 
<< pdiffusion >>
rect 102 35 103 36 
<< pdiffusion >>
rect 103 35 104 36 
<< pdiffusion >>
rect 104 35 105 36 
<< pdiffusion >>
rect 105 35 106 36 
<< m1 >>
rect 106 35 107 36 
<< pdiffusion >>
rect 106 35 107 36 
<< pdiffusion >>
rect 107 35 108 36 
<< m1 >>
rect 109 35 110 36 
<< m1 >>
rect 111 35 112 36 
<< pdiffusion >>
rect 120 35 121 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< m1 >>
rect 124 35 125 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< m1 >>
rect 127 35 128 36 
<< pdiffusion >>
rect 138 35 139 36 
<< m1 >>
rect 139 35 140 36 
<< pdiffusion >>
rect 139 35 140 36 
<< pdiffusion >>
rect 140 35 141 36 
<< pdiffusion >>
rect 141 35 142 36 
<< pdiffusion >>
rect 142 35 143 36 
<< pdiffusion >>
rect 143 35 144 36 
<< m1 >>
rect 154 35 155 36 
<< pdiffusion >>
rect 156 35 157 36 
<< pdiffusion >>
rect 157 35 158 36 
<< pdiffusion >>
rect 158 35 159 36 
<< pdiffusion >>
rect 159 35 160 36 
<< m1 >>
rect 160 35 161 36 
<< pdiffusion >>
rect 160 35 161 36 
<< pdiffusion >>
rect 161 35 162 36 
<< m1 >>
rect 163 35 164 36 
<< m1 >>
rect 169 35 170 36 
<< m2 >>
rect 169 35 170 36 
<< m1 >>
rect 171 35 172 36 
<< m1 >>
rect 19 36 20 37 
<< m1 >>
rect 37 36 38 37 
<< m2 >>
rect 37 36 38 37 
<< m1 >>
rect 42 36 43 37 
<< m1 >>
rect 44 36 45 37 
<< m1 >>
rect 46 36 47 37 
<< m1 >>
rect 55 36 56 37 
<< m2 >>
rect 56 36 57 37 
<< m1 >>
rect 64 36 65 37 
<< m1 >>
rect 73 36 74 37 
<< m1 >>
rect 82 36 83 37 
<< m1 >>
rect 91 36 92 37 
<< m2 >>
rect 92 36 93 37 
<< m1 >>
rect 93 36 94 37 
<< m2 >>
rect 93 36 94 37 
<< m2c >>
rect 93 36 94 37 
<< m1 >>
rect 93 36 94 37 
<< m2 >>
rect 93 36 94 37 
<< m1 >>
rect 94 36 95 37 
<< m1 >>
rect 95 36 96 37 
<< m2 >>
rect 95 36 96 37 
<< m1 >>
rect 96 36 97 37 
<< m1 >>
rect 97 36 98 37 
<< m2 >>
rect 97 36 98 37 
<< m1 >>
rect 98 36 99 37 
<< m1 >>
rect 99 36 100 37 
<< m1 >>
rect 100 36 101 37 
<< m1 >>
rect 106 36 107 37 
<< m1 >>
rect 109 36 110 37 
<< m1 >>
rect 111 36 112 37 
<< m1 >>
rect 124 36 125 37 
<< m1 >>
rect 127 36 128 37 
<< m1 >>
rect 139 36 140 37 
<< m1 >>
rect 154 36 155 37 
<< m1 >>
rect 160 36 161 37 
<< m1 >>
rect 163 36 164 37 
<< m1 >>
rect 169 36 170 37 
<< m2 >>
rect 169 36 170 37 
<< m1 >>
rect 171 36 172 37 
<< m1 >>
rect 19 37 20 38 
<< m1 >>
rect 37 37 38 38 
<< m2 >>
rect 37 37 38 38 
<< m1 >>
rect 42 37 43 38 
<< m1 >>
rect 44 37 45 38 
<< m1 >>
rect 46 37 47 38 
<< m1 >>
rect 55 37 56 38 
<< m2 >>
rect 56 37 57 38 
<< m1 >>
rect 64 37 65 38 
<< m1 >>
rect 73 37 74 38 
<< m1 >>
rect 82 37 83 38 
<< m1 >>
rect 91 37 92 38 
<< m2 >>
rect 95 37 96 38 
<< m2 >>
rect 97 37 98 38 
<< m1 >>
rect 100 37 101 38 
<< m1 >>
rect 106 37 107 38 
<< m1 >>
rect 109 37 110 38 
<< m1 >>
rect 111 37 112 38 
<< m1 >>
rect 124 37 125 38 
<< m1 >>
rect 125 37 126 38 
<< m2 >>
rect 125 37 126 38 
<< m2c >>
rect 125 37 126 38 
<< m1 >>
rect 125 37 126 38 
<< m2 >>
rect 125 37 126 38 
<< m2 >>
rect 126 37 127 38 
<< m1 >>
rect 127 37 128 38 
<< m2 >>
rect 127 37 128 38 
<< m1 >>
rect 139 37 140 38 
<< m1 >>
rect 154 37 155 38 
<< m1 >>
rect 160 37 161 38 
<< m1 >>
rect 163 37 164 38 
<< m1 >>
rect 169 37 170 38 
<< m2 >>
rect 169 37 170 38 
<< m1 >>
rect 171 37 172 38 
<< m1 >>
rect 19 38 20 39 
<< m1 >>
rect 37 38 38 39 
<< m2 >>
rect 37 38 38 39 
<< m1 >>
rect 42 38 43 39 
<< m1 >>
rect 44 38 45 39 
<< m1 >>
rect 46 38 47 39 
<< m1 >>
rect 55 38 56 39 
<< m2 >>
rect 56 38 57 39 
<< m1 >>
rect 64 38 65 39 
<< m1 >>
rect 65 38 66 39 
<< m1 >>
rect 66 38 67 39 
<< m2 >>
rect 66 38 67 39 
<< m2c >>
rect 66 38 67 39 
<< m1 >>
rect 66 38 67 39 
<< m2 >>
rect 66 38 67 39 
<< m1 >>
rect 73 38 74 39 
<< m2 >>
rect 73 38 74 39 
<< m2c >>
rect 73 38 74 39 
<< m1 >>
rect 73 38 74 39 
<< m2 >>
rect 73 38 74 39 
<< m1 >>
rect 82 38 83 39 
<< m1 >>
rect 83 38 84 39 
<< m1 >>
rect 84 38 85 39 
<< m2 >>
rect 84 38 85 39 
<< m2c >>
rect 84 38 85 39 
<< m1 >>
rect 84 38 85 39 
<< m2 >>
rect 84 38 85 39 
<< m1 >>
rect 91 38 92 39 
<< m2 >>
rect 91 38 92 39 
<< m2c >>
rect 91 38 92 39 
<< m1 >>
rect 91 38 92 39 
<< m2 >>
rect 91 38 92 39 
<< m1 >>
rect 95 38 96 39 
<< m2 >>
rect 95 38 96 39 
<< m2c >>
rect 95 38 96 39 
<< m1 >>
rect 95 38 96 39 
<< m2 >>
rect 95 38 96 39 
<< m1 >>
rect 97 38 98 39 
<< m2 >>
rect 97 38 98 39 
<< m2c >>
rect 97 38 98 39 
<< m1 >>
rect 97 38 98 39 
<< m2 >>
rect 97 38 98 39 
<< m1 >>
rect 100 38 101 39 
<< m1 >>
rect 101 38 102 39 
<< m1 >>
rect 102 38 103 39 
<< m2 >>
rect 102 38 103 39 
<< m2c >>
rect 102 38 103 39 
<< m1 >>
rect 102 38 103 39 
<< m2 >>
rect 102 38 103 39 
<< m1 >>
rect 106 38 107 39 
<< m1 >>
rect 109 38 110 39 
<< m1 >>
rect 111 38 112 39 
<< m1 >>
rect 127 38 128 39 
<< m2 >>
rect 127 38 128 39 
<< m1 >>
rect 139 38 140 39 
<< m1 >>
rect 140 38 141 39 
<< m1 >>
rect 141 38 142 39 
<< m1 >>
rect 142 38 143 39 
<< m1 >>
rect 143 38 144 39 
<< m1 >>
rect 144 38 145 39 
<< m1 >>
rect 145 38 146 39 
<< m1 >>
rect 146 38 147 39 
<< m1 >>
rect 154 38 155 39 
<< m1 >>
rect 160 38 161 39 
<< m1 >>
rect 163 38 164 39 
<< m1 >>
rect 169 38 170 39 
<< m2 >>
rect 169 38 170 39 
<< m1 >>
rect 171 38 172 39 
<< m1 >>
rect 19 39 20 40 
<< m1 >>
rect 37 39 38 40 
<< m2 >>
rect 37 39 38 40 
<< m1 >>
rect 42 39 43 40 
<< m1 >>
rect 44 39 45 40 
<< m1 >>
rect 46 39 47 40 
<< m1 >>
rect 55 39 56 40 
<< m2 >>
rect 56 39 57 40 
<< m2 >>
rect 66 39 67 40 
<< m2 >>
rect 73 39 74 40 
<< m2 >>
rect 84 39 85 40 
<< m2 >>
rect 91 39 92 40 
<< m2 >>
rect 92 39 93 40 
<< m2 >>
rect 93 39 94 40 
<< m2 >>
rect 95 39 96 40 
<< m2 >>
rect 97 39 98 40 
<< m2 >>
rect 102 39 103 40 
<< m2 >>
rect 104 39 105 40 
<< m1 >>
rect 105 39 106 40 
<< m2 >>
rect 105 39 106 40 
<< m2c >>
rect 105 39 106 40 
<< m1 >>
rect 105 39 106 40 
<< m2 >>
rect 105 39 106 40 
<< m1 >>
rect 106 39 107 40 
<< m1 >>
rect 109 39 110 40 
<< m1 >>
rect 111 39 112 40 
<< m1 >>
rect 127 39 128 40 
<< m2 >>
rect 127 39 128 40 
<< m1 >>
rect 146 39 147 40 
<< m1 >>
rect 154 39 155 40 
<< m1 >>
rect 160 39 161 40 
<< m1 >>
rect 163 39 164 40 
<< m1 >>
rect 169 39 170 40 
<< m2 >>
rect 169 39 170 40 
<< m1 >>
rect 171 39 172 40 
<< m1 >>
rect 19 40 20 41 
<< m1 >>
rect 37 40 38 41 
<< m2 >>
rect 37 40 38 41 
<< m1 >>
rect 42 40 43 41 
<< m1 >>
rect 44 40 45 41 
<< m1 >>
rect 46 40 47 41 
<< m1 >>
rect 55 40 56 41 
<< m1 >>
rect 56 40 57 41 
<< m2 >>
rect 56 40 57 41 
<< m1 >>
rect 57 40 58 41 
<< m1 >>
rect 58 40 59 41 
<< m1 >>
rect 59 40 60 41 
<< m1 >>
rect 60 40 61 41 
<< m1 >>
rect 61 40 62 41 
<< m1 >>
rect 62 40 63 41 
<< m1 >>
rect 63 40 64 41 
<< m1 >>
rect 64 40 65 41 
<< m1 >>
rect 65 40 66 41 
<< m1 >>
rect 66 40 67 41 
<< m2 >>
rect 66 40 67 41 
<< m1 >>
rect 67 40 68 41 
<< m1 >>
rect 68 40 69 41 
<< m1 >>
rect 69 40 70 41 
<< m1 >>
rect 70 40 71 41 
<< m1 >>
rect 71 40 72 41 
<< m1 >>
rect 72 40 73 41 
<< m1 >>
rect 73 40 74 41 
<< m2 >>
rect 73 40 74 41 
<< m1 >>
rect 74 40 75 41 
<< m1 >>
rect 75 40 76 41 
<< m1 >>
rect 76 40 77 41 
<< m1 >>
rect 77 40 78 41 
<< m1 >>
rect 78 40 79 41 
<< m1 >>
rect 79 40 80 41 
<< m1 >>
rect 80 40 81 41 
<< m1 >>
rect 81 40 82 41 
<< m1 >>
rect 82 40 83 41 
<< m1 >>
rect 83 40 84 41 
<< m1 >>
rect 84 40 85 41 
<< m2 >>
rect 84 40 85 41 
<< m1 >>
rect 85 40 86 41 
<< m1 >>
rect 86 40 87 41 
<< m1 >>
rect 87 40 88 41 
<< m1 >>
rect 88 40 89 41 
<< m1 >>
rect 89 40 90 41 
<< m1 >>
rect 90 40 91 41 
<< m1 >>
rect 91 40 92 41 
<< m1 >>
rect 92 40 93 41 
<< m1 >>
rect 93 40 94 41 
<< m2 >>
rect 93 40 94 41 
<< m1 >>
rect 94 40 95 41 
<< m1 >>
rect 95 40 96 41 
<< m2 >>
rect 95 40 96 41 
<< m1 >>
rect 96 40 97 41 
<< m1 >>
rect 97 40 98 41 
<< m2 >>
rect 97 40 98 41 
<< m1 >>
rect 98 40 99 41 
<< m1 >>
rect 99 40 100 41 
<< m1 >>
rect 100 40 101 41 
<< m1 >>
rect 101 40 102 41 
<< m1 >>
rect 102 40 103 41 
<< m2 >>
rect 102 40 103 41 
<< m1 >>
rect 103 40 104 41 
<< m2 >>
rect 103 40 104 41 
<< m2 >>
rect 104 40 105 41 
<< m1 >>
rect 109 40 110 41 
<< m1 >>
rect 111 40 112 41 
<< m1 >>
rect 127 40 128 41 
<< m2 >>
rect 127 40 128 41 
<< m1 >>
rect 146 40 147 41 
<< m1 >>
rect 154 40 155 41 
<< m1 >>
rect 160 40 161 41 
<< m1 >>
rect 163 40 164 41 
<< m1 >>
rect 169 40 170 41 
<< m2 >>
rect 169 40 170 41 
<< m1 >>
rect 171 40 172 41 
<< m1 >>
rect 19 41 20 42 
<< m1 >>
rect 37 41 38 42 
<< m2 >>
rect 37 41 38 42 
<< m1 >>
rect 42 41 43 42 
<< m2 >>
rect 42 41 43 42 
<< m2c >>
rect 42 41 43 42 
<< m1 >>
rect 42 41 43 42 
<< m2 >>
rect 42 41 43 42 
<< m2 >>
rect 43 41 44 42 
<< m1 >>
rect 44 41 45 42 
<< m2 >>
rect 44 41 45 42 
<< m2 >>
rect 45 41 46 42 
<< m1 >>
rect 46 41 47 42 
<< m2 >>
rect 46 41 47 42 
<< m2 >>
rect 47 41 48 42 
<< m1 >>
rect 48 41 49 42 
<< m2 >>
rect 48 41 49 42 
<< m2c >>
rect 48 41 49 42 
<< m1 >>
rect 48 41 49 42 
<< m2 >>
rect 48 41 49 42 
<< m1 >>
rect 49 41 50 42 
<< m1 >>
rect 50 41 51 42 
<< m1 >>
rect 51 41 52 42 
<< m1 >>
rect 52 41 53 42 
<< m1 >>
rect 53 41 54 42 
<< m2 >>
rect 53 41 54 42 
<< m2 >>
rect 54 41 55 42 
<< m2 >>
rect 56 41 57 42 
<< m2 >>
rect 57 41 58 42 
<< m2 >>
rect 58 41 59 42 
<< m2 >>
rect 59 41 60 42 
<< m2 >>
rect 60 41 61 42 
<< m2 >>
rect 61 41 62 42 
<< m2 >>
rect 62 41 63 42 
<< m2 >>
rect 63 41 64 42 
<< m2 >>
rect 64 41 65 42 
<< m2 >>
rect 66 41 67 42 
<< m2 >>
rect 73 41 74 42 
<< m2 >>
rect 84 41 85 42 
<< m2 >>
rect 85 41 86 42 
<< m2 >>
rect 86 41 87 42 
<< m2 >>
rect 87 41 88 42 
<< m2 >>
rect 88 41 89 42 
<< m2 >>
rect 89 41 90 42 
<< m2 >>
rect 90 41 91 42 
<< m2 >>
rect 91 41 92 42 
<< m2 >>
rect 93 41 94 42 
<< m2 >>
rect 95 41 96 42 
<< m2 >>
rect 97 41 98 42 
<< m1 >>
rect 103 41 104 42 
<< m1 >>
rect 109 41 110 42 
<< m1 >>
rect 111 41 112 42 
<< m1 >>
rect 127 41 128 42 
<< m2 >>
rect 127 41 128 42 
<< m1 >>
rect 146 41 147 42 
<< m1 >>
rect 154 41 155 42 
<< m1 >>
rect 160 41 161 42 
<< m1 >>
rect 161 41 162 42 
<< m2 >>
rect 161 41 162 42 
<< m2c >>
rect 161 41 162 42 
<< m1 >>
rect 161 41 162 42 
<< m2 >>
rect 161 41 162 42 
<< m2 >>
rect 162 41 163 42 
<< m1 >>
rect 163 41 164 42 
<< m2 >>
rect 163 41 164 42 
<< m2 >>
rect 164 41 165 42 
<< m1 >>
rect 169 41 170 42 
<< m2 >>
rect 169 41 170 42 
<< m1 >>
rect 171 41 172 42 
<< m1 >>
rect 19 42 20 43 
<< m1 >>
rect 37 42 38 43 
<< m2 >>
rect 37 42 38 43 
<< m1 >>
rect 44 42 45 43 
<< m1 >>
rect 46 42 47 43 
<< m1 >>
rect 54 42 55 43 
<< m2 >>
rect 54 42 55 43 
<< m2c >>
rect 54 42 55 43 
<< m1 >>
rect 54 42 55 43 
<< m2 >>
rect 54 42 55 43 
<< m1 >>
rect 64 42 65 43 
<< m2 >>
rect 64 42 65 43 
<< m2c >>
rect 64 42 65 43 
<< m1 >>
rect 64 42 65 43 
<< m2 >>
rect 64 42 65 43 
<< m1 >>
rect 66 42 67 43 
<< m2 >>
rect 66 42 67 43 
<< m2c >>
rect 66 42 67 43 
<< m1 >>
rect 66 42 67 43 
<< m2 >>
rect 66 42 67 43 
<< m1 >>
rect 73 42 74 43 
<< m2 >>
rect 73 42 74 43 
<< m2c >>
rect 73 42 74 43 
<< m1 >>
rect 73 42 74 43 
<< m2 >>
rect 73 42 74 43 
<< m1 >>
rect 91 42 92 43 
<< m2 >>
rect 91 42 92 43 
<< m2c >>
rect 91 42 92 43 
<< m1 >>
rect 91 42 92 43 
<< m2 >>
rect 91 42 92 43 
<< m1 >>
rect 93 42 94 43 
<< m2 >>
rect 93 42 94 43 
<< m2c >>
rect 93 42 94 43 
<< m1 >>
rect 93 42 94 43 
<< m2 >>
rect 93 42 94 43 
<< m1 >>
rect 95 42 96 43 
<< m2 >>
rect 95 42 96 43 
<< m2c >>
rect 95 42 96 43 
<< m1 >>
rect 95 42 96 43 
<< m2 >>
rect 95 42 96 43 
<< m1 >>
rect 97 42 98 43 
<< m2 >>
rect 97 42 98 43 
<< m2c >>
rect 97 42 98 43 
<< m1 >>
rect 97 42 98 43 
<< m2 >>
rect 97 42 98 43 
<< m1 >>
rect 98 42 99 43 
<< m1 >>
rect 99 42 100 43 
<< m1 >>
rect 100 42 101 43 
<< m1 >>
rect 101 42 102 43 
<< m2 >>
rect 101 42 102 43 
<< m2c >>
rect 101 42 102 43 
<< m1 >>
rect 101 42 102 43 
<< m2 >>
rect 101 42 102 43 
<< m2 >>
rect 102 42 103 43 
<< m1 >>
rect 103 42 104 43 
<< m2 >>
rect 103 42 104 43 
<< m2 >>
rect 104 42 105 43 
<< m1 >>
rect 105 42 106 43 
<< m2 >>
rect 105 42 106 43 
<< m2c >>
rect 105 42 106 43 
<< m1 >>
rect 105 42 106 43 
<< m2 >>
rect 105 42 106 43 
<< m1 >>
rect 106 42 107 43 
<< m1 >>
rect 109 42 110 43 
<< m1 >>
rect 111 42 112 43 
<< m1 >>
rect 127 42 128 43 
<< m2 >>
rect 127 42 128 43 
<< m1 >>
rect 146 42 147 43 
<< m1 >>
rect 154 42 155 43 
<< m1 >>
rect 163 42 164 43 
<< m2 >>
rect 164 42 165 43 
<< m1 >>
rect 169 42 170 43 
<< m2 >>
rect 169 42 170 43 
<< m1 >>
rect 171 42 172 43 
<< m1 >>
rect 19 43 20 44 
<< m1 >>
rect 37 43 38 44 
<< m2 >>
rect 37 43 38 44 
<< m1 >>
rect 44 43 45 44 
<< m2 >>
rect 44 43 45 44 
<< m2c >>
rect 44 43 45 44 
<< m1 >>
rect 44 43 45 44 
<< m2 >>
rect 44 43 45 44 
<< m2 >>
rect 45 43 46 44 
<< m1 >>
rect 46 43 47 44 
<< m2 >>
rect 46 43 47 44 
<< m2 >>
rect 47 43 48 44 
<< m1 >>
rect 48 43 49 44 
<< m2 >>
rect 48 43 49 44 
<< m2c >>
rect 48 43 49 44 
<< m1 >>
rect 48 43 49 44 
<< m2 >>
rect 48 43 49 44 
<< m1 >>
rect 49 43 50 44 
<< m1 >>
rect 50 43 51 44 
<< m1 >>
rect 51 43 52 44 
<< m1 >>
rect 52 43 53 44 
<< m1 >>
rect 54 43 55 44 
<< m1 >>
rect 64 43 65 44 
<< m1 >>
rect 66 43 67 44 
<< m1 >>
rect 73 43 74 44 
<< m1 >>
rect 91 43 92 44 
<< m1 >>
rect 93 43 94 44 
<< m1 >>
rect 95 43 96 44 
<< m1 >>
rect 103 43 104 44 
<< m1 >>
rect 106 43 107 44 
<< m1 >>
rect 109 43 110 44 
<< m1 >>
rect 111 43 112 44 
<< m1 >>
rect 113 43 114 44 
<< m1 >>
rect 114 43 115 44 
<< m1 >>
rect 115 43 116 44 
<< m1 >>
rect 116 43 117 44 
<< m1 >>
rect 117 43 118 44 
<< m1 >>
rect 118 43 119 44 
<< m1 >>
rect 119 43 120 44 
<< m1 >>
rect 120 43 121 44 
<< m1 >>
rect 121 43 122 44 
<< m1 >>
rect 122 43 123 44 
<< m1 >>
rect 123 43 124 44 
<< m1 >>
rect 124 43 125 44 
<< m1 >>
rect 127 43 128 44 
<< m2 >>
rect 127 43 128 44 
<< m1 >>
rect 146 43 147 44 
<< m1 >>
rect 154 43 155 44 
<< m1 >>
rect 155 43 156 44 
<< m1 >>
rect 156 43 157 44 
<< m1 >>
rect 157 43 158 44 
<< m1 >>
rect 158 43 159 44 
<< m1 >>
rect 159 43 160 44 
<< m1 >>
rect 160 43 161 44 
<< m1 >>
rect 163 43 164 44 
<< m2 >>
rect 164 43 165 44 
<< m1 >>
rect 169 43 170 44 
<< m2 >>
rect 169 43 170 44 
<< m1 >>
rect 171 43 172 44 
<< m1 >>
rect 19 44 20 45 
<< m1 >>
rect 37 44 38 45 
<< m2 >>
rect 37 44 38 45 
<< m1 >>
rect 46 44 47 45 
<< m1 >>
rect 52 44 53 45 
<< m1 >>
rect 54 44 55 45 
<< m1 >>
rect 64 44 65 45 
<< m1 >>
rect 66 44 67 45 
<< m1 >>
rect 73 44 74 45 
<< m1 >>
rect 91 44 92 45 
<< m1 >>
rect 93 44 94 45 
<< m1 >>
rect 95 44 96 45 
<< m1 >>
rect 103 44 104 45 
<< m1 >>
rect 106 44 107 45 
<< m1 >>
rect 109 44 110 45 
<< m1 >>
rect 111 44 112 45 
<< m1 >>
rect 113 44 114 45 
<< m1 >>
rect 124 44 125 45 
<< m1 >>
rect 127 44 128 45 
<< m2 >>
rect 127 44 128 45 
<< m1 >>
rect 146 44 147 45 
<< m1 >>
rect 160 44 161 45 
<< m1 >>
rect 163 44 164 45 
<< m2 >>
rect 164 44 165 45 
<< m1 >>
rect 169 44 170 45 
<< m2 >>
rect 169 44 170 45 
<< m1 >>
rect 171 44 172 45 
<< m1 >>
rect 13 45 14 46 
<< m1 >>
rect 14 45 15 46 
<< m1 >>
rect 15 45 16 46 
<< m1 >>
rect 16 45 17 46 
<< m1 >>
rect 17 45 18 46 
<< m2 >>
rect 17 45 18 46 
<< m2c >>
rect 17 45 18 46 
<< m1 >>
rect 17 45 18 46 
<< m2 >>
rect 17 45 18 46 
<< m2 >>
rect 18 45 19 46 
<< m1 >>
rect 19 45 20 46 
<< m2 >>
rect 19 45 20 46 
<< m2 >>
rect 20 45 21 46 
<< m1 >>
rect 21 45 22 46 
<< m2 >>
rect 21 45 22 46 
<< m2c >>
rect 21 45 22 46 
<< m1 >>
rect 21 45 22 46 
<< m2 >>
rect 21 45 22 46 
<< m1 >>
rect 22 45 23 46 
<< m1 >>
rect 23 45 24 46 
<< m1 >>
rect 37 45 38 46 
<< m2 >>
rect 37 45 38 46 
<< m1 >>
rect 46 45 47 46 
<< m1 >>
rect 52 45 53 46 
<< m1 >>
rect 54 45 55 46 
<< m1 >>
rect 64 45 65 46 
<< m1 >>
rect 66 45 67 46 
<< m1 >>
rect 73 45 74 46 
<< m1 >>
rect 85 45 86 46 
<< m1 >>
rect 86 45 87 46 
<< m1 >>
rect 87 45 88 46 
<< m1 >>
rect 88 45 89 46 
<< m1 >>
rect 89 45 90 46 
<< m2 >>
rect 89 45 90 46 
<< m2c >>
rect 89 45 90 46 
<< m1 >>
rect 89 45 90 46 
<< m2 >>
rect 89 45 90 46 
<< m2 >>
rect 90 45 91 46 
<< m1 >>
rect 91 45 92 46 
<< m2 >>
rect 91 45 92 46 
<< m2 >>
rect 92 45 93 46 
<< m1 >>
rect 93 45 94 46 
<< m2 >>
rect 93 45 94 46 
<< m2 >>
rect 94 45 95 46 
<< m1 >>
rect 95 45 96 46 
<< m2 >>
rect 95 45 96 46 
<< m2c >>
rect 95 45 96 46 
<< m1 >>
rect 95 45 96 46 
<< m2 >>
rect 95 45 96 46 
<< m1 >>
rect 103 45 104 46 
<< m1 >>
rect 106 45 107 46 
<< m1 >>
rect 109 45 110 46 
<< m1 >>
rect 111 45 112 46 
<< m1 >>
rect 113 45 114 46 
<< m1 >>
rect 124 45 125 46 
<< m1 >>
rect 127 45 128 46 
<< m2 >>
rect 127 45 128 46 
<< m1 >>
rect 146 45 147 46 
<< m1 >>
rect 160 45 161 46 
<< m1 >>
rect 163 45 164 46 
<< m2 >>
rect 164 45 165 46 
<< m1 >>
rect 169 45 170 46 
<< m2 >>
rect 169 45 170 46 
<< m1 >>
rect 171 45 172 46 
<< m1 >>
rect 13 46 14 47 
<< m1 >>
rect 19 46 20 47 
<< m1 >>
rect 23 46 24 47 
<< m1 >>
rect 25 46 26 47 
<< m1 >>
rect 26 46 27 47 
<< m1 >>
rect 27 46 28 47 
<< m1 >>
rect 28 46 29 47 
<< m1 >>
rect 29 46 30 47 
<< m1 >>
rect 30 46 31 47 
<< m1 >>
rect 31 46 32 47 
<< m1 >>
rect 37 46 38 47 
<< m2 >>
rect 37 46 38 47 
<< m1 >>
rect 43 46 44 47 
<< m1 >>
rect 44 46 45 47 
<< m2 >>
rect 44 46 45 47 
<< m2c >>
rect 44 46 45 47 
<< m1 >>
rect 44 46 45 47 
<< m2 >>
rect 44 46 45 47 
<< m2 >>
rect 45 46 46 47 
<< m1 >>
rect 46 46 47 47 
<< m2 >>
rect 46 46 47 47 
<< m2 >>
rect 47 46 48 47 
<< m1 >>
rect 48 46 49 47 
<< m2 >>
rect 48 46 49 47 
<< m2c >>
rect 48 46 49 47 
<< m1 >>
rect 48 46 49 47 
<< m2 >>
rect 48 46 49 47 
<< m1 >>
rect 49 46 50 47 
<< m1 >>
rect 52 46 53 47 
<< m1 >>
rect 54 46 55 47 
<< m1 >>
rect 55 46 56 47 
<< m2 >>
rect 63 46 64 47 
<< m1 >>
rect 64 46 65 47 
<< m2 >>
rect 64 46 65 47 
<< m2 >>
rect 65 46 66 47 
<< m1 >>
rect 66 46 67 47 
<< m2 >>
rect 66 46 67 47 
<< m2c >>
rect 66 46 67 47 
<< m1 >>
rect 66 46 67 47 
<< m2 >>
rect 66 46 67 47 
<< m1 >>
rect 73 46 74 47 
<< m1 >>
rect 85 46 86 47 
<< m1 >>
rect 91 46 92 47 
<< m1 >>
rect 93 46 94 47 
<< m1 >>
rect 103 46 104 47 
<< m1 >>
rect 106 46 107 47 
<< m1 >>
rect 109 46 110 47 
<< m1 >>
rect 111 46 112 47 
<< m1 >>
rect 113 46 114 47 
<< m1 >>
rect 124 46 125 47 
<< m1 >>
rect 127 46 128 47 
<< m2 >>
rect 127 46 128 47 
<< m1 >>
rect 142 46 143 47 
<< m1 >>
rect 143 46 144 47 
<< m1 >>
rect 144 46 145 47 
<< m2 >>
rect 144 46 145 47 
<< m2c >>
rect 144 46 145 47 
<< m1 >>
rect 144 46 145 47 
<< m2 >>
rect 144 46 145 47 
<< m2 >>
rect 145 46 146 47 
<< m1 >>
rect 146 46 147 47 
<< m2 >>
rect 146 46 147 47 
<< m2 >>
rect 147 46 148 47 
<< m1 >>
rect 148 46 149 47 
<< m2 >>
rect 148 46 149 47 
<< m2c >>
rect 148 46 149 47 
<< m1 >>
rect 148 46 149 47 
<< m2 >>
rect 148 46 149 47 
<< m1 >>
rect 160 46 161 47 
<< m1 >>
rect 163 46 164 47 
<< m2 >>
rect 164 46 165 47 
<< m1 >>
rect 169 46 170 47 
<< m2 >>
rect 169 46 170 47 
<< m1 >>
rect 171 46 172 47 
<< m1 >>
rect 13 47 14 48 
<< m1 >>
rect 19 47 20 48 
<< m1 >>
rect 23 47 24 48 
<< m1 >>
rect 25 47 26 48 
<< m1 >>
rect 31 47 32 48 
<< m1 >>
rect 37 47 38 48 
<< m2 >>
rect 37 47 38 48 
<< m1 >>
rect 43 47 44 48 
<< m1 >>
rect 46 47 47 48 
<< m1 >>
rect 49 47 50 48 
<< m1 >>
rect 52 47 53 48 
<< m1 >>
rect 55 47 56 48 
<< m2 >>
rect 63 47 64 48 
<< m1 >>
rect 64 47 65 48 
<< m1 >>
rect 73 47 74 48 
<< m1 >>
rect 85 47 86 48 
<< m1 >>
rect 91 47 92 48 
<< m1 >>
rect 93 47 94 48 
<< m1 >>
rect 103 47 104 48 
<< m1 >>
rect 106 47 107 48 
<< m1 >>
rect 109 47 110 48 
<< m1 >>
rect 111 47 112 48 
<< m1 >>
rect 113 47 114 48 
<< m1 >>
rect 124 47 125 48 
<< m1 >>
rect 127 47 128 48 
<< m2 >>
rect 127 47 128 48 
<< m1 >>
rect 142 47 143 48 
<< m1 >>
rect 146 47 147 48 
<< m1 >>
rect 148 47 149 48 
<< m1 >>
rect 160 47 161 48 
<< m1 >>
rect 163 47 164 48 
<< m2 >>
rect 164 47 165 48 
<< m1 >>
rect 169 47 170 48 
<< m2 >>
rect 169 47 170 48 
<< m1 >>
rect 171 47 172 48 
<< pdiffusion >>
rect 12 48 13 49 
<< m1 >>
rect 13 48 14 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< m1 >>
rect 19 48 20 49 
<< m1 >>
rect 23 48 24 49 
<< m1 >>
rect 25 48 26 49 
<< pdiffusion >>
rect 30 48 31 49 
<< m1 >>
rect 31 48 32 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< m1 >>
rect 37 48 38 49 
<< m2 >>
rect 37 48 38 49 
<< m1 >>
rect 43 48 44 49 
<< m1 >>
rect 46 48 47 49 
<< pdiffusion >>
rect 48 48 49 49 
<< m1 >>
rect 49 48 50 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< m1 >>
rect 52 48 53 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 55 48 56 49 
<< m2 >>
rect 63 48 64 49 
<< m1 >>
rect 64 48 65 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< m1 >>
rect 73 48 74 49 
<< pdiffusion >>
rect 84 48 85 49 
<< m1 >>
rect 85 48 86 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< m1 >>
rect 93 48 94 49 
<< pdiffusion >>
rect 102 48 103 49 
<< m1 >>
rect 103 48 104 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< m1 >>
rect 106 48 107 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< m1 >>
rect 109 48 110 49 
<< m1 >>
rect 111 48 112 49 
<< m1 >>
rect 113 48 114 49 
<< pdiffusion >>
rect 120 48 121 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< m1 >>
rect 124 48 125 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< m1 >>
rect 127 48 128 49 
<< m2 >>
rect 127 48 128 49 
<< pdiffusion >>
rect 138 48 139 49 
<< pdiffusion >>
rect 139 48 140 49 
<< pdiffusion >>
rect 140 48 141 49 
<< pdiffusion >>
rect 141 48 142 49 
<< m1 >>
rect 142 48 143 49 
<< pdiffusion >>
rect 142 48 143 49 
<< pdiffusion >>
rect 143 48 144 49 
<< m1 >>
rect 146 48 147 49 
<< m1 >>
rect 148 48 149 49 
<< pdiffusion >>
rect 156 48 157 49 
<< pdiffusion >>
rect 157 48 158 49 
<< pdiffusion >>
rect 158 48 159 49 
<< pdiffusion >>
rect 159 48 160 49 
<< m1 >>
rect 160 48 161 49 
<< pdiffusion >>
rect 160 48 161 49 
<< pdiffusion >>
rect 161 48 162 49 
<< m1 >>
rect 163 48 164 49 
<< m2 >>
rect 164 48 165 49 
<< m1 >>
rect 169 48 170 49 
<< m2 >>
rect 169 48 170 49 
<< m1 >>
rect 171 48 172 49 
<< pdiffusion >>
rect 174 48 175 49 
<< pdiffusion >>
rect 175 48 176 49 
<< pdiffusion >>
rect 176 48 177 49 
<< pdiffusion >>
rect 177 48 178 49 
<< pdiffusion >>
rect 178 48 179 49 
<< pdiffusion >>
rect 179 48 180 49 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< m1 >>
rect 19 49 20 50 
<< m1 >>
rect 23 49 24 50 
<< m1 >>
rect 25 49 26 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< m1 >>
rect 37 49 38 50 
<< m2 >>
rect 37 49 38 50 
<< m1 >>
rect 43 49 44 50 
<< m1 >>
rect 46 49 47 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 55 49 56 50 
<< m2 >>
rect 63 49 64 50 
<< m1 >>
rect 64 49 65 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< m1 >>
rect 73 49 74 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< m1 >>
rect 93 49 94 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< m1 >>
rect 109 49 110 50 
<< m1 >>
rect 111 49 112 50 
<< m1 >>
rect 113 49 114 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< m1 >>
rect 127 49 128 50 
<< m2 >>
rect 127 49 128 50 
<< pdiffusion >>
rect 138 49 139 50 
<< pdiffusion >>
rect 139 49 140 50 
<< pdiffusion >>
rect 140 49 141 50 
<< pdiffusion >>
rect 141 49 142 50 
<< pdiffusion >>
rect 142 49 143 50 
<< pdiffusion >>
rect 143 49 144 50 
<< m1 >>
rect 146 49 147 50 
<< m1 >>
rect 148 49 149 50 
<< pdiffusion >>
rect 156 49 157 50 
<< pdiffusion >>
rect 157 49 158 50 
<< pdiffusion >>
rect 158 49 159 50 
<< pdiffusion >>
rect 159 49 160 50 
<< pdiffusion >>
rect 160 49 161 50 
<< pdiffusion >>
rect 161 49 162 50 
<< m1 >>
rect 163 49 164 50 
<< m2 >>
rect 164 49 165 50 
<< m1 >>
rect 169 49 170 50 
<< m2 >>
rect 169 49 170 50 
<< m1 >>
rect 171 49 172 50 
<< pdiffusion >>
rect 174 49 175 50 
<< pdiffusion >>
rect 175 49 176 50 
<< pdiffusion >>
rect 176 49 177 50 
<< pdiffusion >>
rect 177 49 178 50 
<< pdiffusion >>
rect 178 49 179 50 
<< pdiffusion >>
rect 179 49 180 50 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< m1 >>
rect 19 50 20 51 
<< m1 >>
rect 23 50 24 51 
<< m1 >>
rect 25 50 26 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< m1 >>
rect 37 50 38 51 
<< m2 >>
rect 37 50 38 51 
<< m1 >>
rect 43 50 44 51 
<< m1 >>
rect 46 50 47 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 55 50 56 51 
<< m2 >>
rect 63 50 64 51 
<< m1 >>
rect 64 50 65 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< m1 >>
rect 73 50 74 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< m1 >>
rect 93 50 94 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< m1 >>
rect 109 50 110 51 
<< m1 >>
rect 111 50 112 51 
<< m1 >>
rect 113 50 114 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< m1 >>
rect 127 50 128 51 
<< m2 >>
rect 127 50 128 51 
<< pdiffusion >>
rect 138 50 139 51 
<< pdiffusion >>
rect 139 50 140 51 
<< pdiffusion >>
rect 140 50 141 51 
<< pdiffusion >>
rect 141 50 142 51 
<< pdiffusion >>
rect 142 50 143 51 
<< pdiffusion >>
rect 143 50 144 51 
<< m1 >>
rect 146 50 147 51 
<< m1 >>
rect 148 50 149 51 
<< pdiffusion >>
rect 156 50 157 51 
<< pdiffusion >>
rect 157 50 158 51 
<< pdiffusion >>
rect 158 50 159 51 
<< pdiffusion >>
rect 159 50 160 51 
<< pdiffusion >>
rect 160 50 161 51 
<< pdiffusion >>
rect 161 50 162 51 
<< m1 >>
rect 163 50 164 51 
<< m2 >>
rect 164 50 165 51 
<< m1 >>
rect 169 50 170 51 
<< m2 >>
rect 169 50 170 51 
<< m1 >>
rect 171 50 172 51 
<< pdiffusion >>
rect 174 50 175 51 
<< pdiffusion >>
rect 175 50 176 51 
<< pdiffusion >>
rect 176 50 177 51 
<< pdiffusion >>
rect 177 50 178 51 
<< pdiffusion >>
rect 178 50 179 51 
<< pdiffusion >>
rect 179 50 180 51 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< m1 >>
rect 19 51 20 52 
<< m1 >>
rect 23 51 24 52 
<< m1 >>
rect 25 51 26 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< m1 >>
rect 37 51 38 52 
<< m2 >>
rect 37 51 38 52 
<< m1 >>
rect 43 51 44 52 
<< m1 >>
rect 46 51 47 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 55 51 56 52 
<< m2 >>
rect 63 51 64 52 
<< m1 >>
rect 64 51 65 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< m1 >>
rect 73 51 74 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< m1 >>
rect 93 51 94 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< m1 >>
rect 109 51 110 52 
<< m1 >>
rect 111 51 112 52 
<< m1 >>
rect 113 51 114 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< m1 >>
rect 127 51 128 52 
<< m2 >>
rect 127 51 128 52 
<< pdiffusion >>
rect 138 51 139 52 
<< pdiffusion >>
rect 139 51 140 52 
<< pdiffusion >>
rect 140 51 141 52 
<< pdiffusion >>
rect 141 51 142 52 
<< pdiffusion >>
rect 142 51 143 52 
<< pdiffusion >>
rect 143 51 144 52 
<< m1 >>
rect 146 51 147 52 
<< m1 >>
rect 148 51 149 52 
<< pdiffusion >>
rect 156 51 157 52 
<< pdiffusion >>
rect 157 51 158 52 
<< pdiffusion >>
rect 158 51 159 52 
<< pdiffusion >>
rect 159 51 160 52 
<< pdiffusion >>
rect 160 51 161 52 
<< pdiffusion >>
rect 161 51 162 52 
<< m1 >>
rect 163 51 164 52 
<< m2 >>
rect 164 51 165 52 
<< m1 >>
rect 169 51 170 52 
<< m2 >>
rect 169 51 170 52 
<< m1 >>
rect 171 51 172 52 
<< pdiffusion >>
rect 174 51 175 52 
<< pdiffusion >>
rect 175 51 176 52 
<< pdiffusion >>
rect 176 51 177 52 
<< pdiffusion >>
rect 177 51 178 52 
<< pdiffusion >>
rect 178 51 179 52 
<< pdiffusion >>
rect 179 51 180 52 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< m1 >>
rect 19 52 20 53 
<< m1 >>
rect 23 52 24 53 
<< m1 >>
rect 25 52 26 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< m1 >>
rect 37 52 38 53 
<< m2 >>
rect 37 52 38 53 
<< m1 >>
rect 43 52 44 53 
<< m1 >>
rect 46 52 47 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 55 52 56 53 
<< m2 >>
rect 63 52 64 53 
<< m1 >>
rect 64 52 65 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< m1 >>
rect 73 52 74 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< m1 >>
rect 93 52 94 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< m1 >>
rect 109 52 110 53 
<< m1 >>
rect 111 52 112 53 
<< m1 >>
rect 113 52 114 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< m1 >>
rect 127 52 128 53 
<< m2 >>
rect 127 52 128 53 
<< pdiffusion >>
rect 138 52 139 53 
<< pdiffusion >>
rect 139 52 140 53 
<< pdiffusion >>
rect 140 52 141 53 
<< pdiffusion >>
rect 141 52 142 53 
<< pdiffusion >>
rect 142 52 143 53 
<< pdiffusion >>
rect 143 52 144 53 
<< m1 >>
rect 146 52 147 53 
<< m1 >>
rect 148 52 149 53 
<< pdiffusion >>
rect 156 52 157 53 
<< pdiffusion >>
rect 157 52 158 53 
<< pdiffusion >>
rect 158 52 159 53 
<< pdiffusion >>
rect 159 52 160 53 
<< pdiffusion >>
rect 160 52 161 53 
<< pdiffusion >>
rect 161 52 162 53 
<< m1 >>
rect 163 52 164 53 
<< m2 >>
rect 164 52 165 53 
<< m1 >>
rect 169 52 170 53 
<< m2 >>
rect 169 52 170 53 
<< m1 >>
rect 171 52 172 53 
<< pdiffusion >>
rect 174 52 175 53 
<< pdiffusion >>
rect 175 52 176 53 
<< pdiffusion >>
rect 176 52 177 53 
<< pdiffusion >>
rect 177 52 178 53 
<< pdiffusion >>
rect 178 52 179 53 
<< pdiffusion >>
rect 179 52 180 53 
<< pdiffusion >>
rect 12 53 13 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< m1 >>
rect 19 53 20 54 
<< m1 >>
rect 23 53 24 54 
<< m1 >>
rect 25 53 26 54 
<< pdiffusion >>
rect 30 53 31 54 
<< m1 >>
rect 31 53 32 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< m1 >>
rect 34 53 35 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< m1 >>
rect 37 53 38 54 
<< m2 >>
rect 37 53 38 54 
<< m1 >>
rect 43 53 44 54 
<< m1 >>
rect 46 53 47 54 
<< pdiffusion >>
rect 48 53 49 54 
<< m1 >>
rect 49 53 50 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< m1 >>
rect 52 53 53 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 55 53 56 54 
<< m2 >>
rect 63 53 64 54 
<< m1 >>
rect 64 53 65 54 
<< pdiffusion >>
rect 66 53 67 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< m1 >>
rect 73 53 74 54 
<< pdiffusion >>
rect 84 53 85 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< m1 >>
rect 88 53 89 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< m1 >>
rect 93 53 94 54 
<< pdiffusion >>
rect 102 53 103 54 
<< m1 >>
rect 103 53 104 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< m1 >>
rect 106 53 107 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< m1 >>
rect 109 53 110 54 
<< m1 >>
rect 111 53 112 54 
<< m1 >>
rect 113 53 114 54 
<< pdiffusion >>
rect 120 53 121 54 
<< m1 >>
rect 121 53 122 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< m1 >>
rect 127 53 128 54 
<< m2 >>
rect 127 53 128 54 
<< pdiffusion >>
rect 138 53 139 54 
<< m1 >>
rect 139 53 140 54 
<< pdiffusion >>
rect 139 53 140 54 
<< pdiffusion >>
rect 140 53 141 54 
<< pdiffusion >>
rect 141 53 142 54 
<< m1 >>
rect 142 53 143 54 
<< pdiffusion >>
rect 142 53 143 54 
<< pdiffusion >>
rect 143 53 144 54 
<< m1 >>
rect 146 53 147 54 
<< m1 >>
rect 148 53 149 54 
<< pdiffusion >>
rect 156 53 157 54 
<< m1 >>
rect 157 53 158 54 
<< pdiffusion >>
rect 157 53 158 54 
<< pdiffusion >>
rect 158 53 159 54 
<< pdiffusion >>
rect 159 53 160 54 
<< m1 >>
rect 160 53 161 54 
<< pdiffusion >>
rect 160 53 161 54 
<< pdiffusion >>
rect 161 53 162 54 
<< m1 >>
rect 163 53 164 54 
<< m2 >>
rect 164 53 165 54 
<< m1 >>
rect 169 53 170 54 
<< m2 >>
rect 169 53 170 54 
<< m1 >>
rect 171 53 172 54 
<< pdiffusion >>
rect 174 53 175 54 
<< pdiffusion >>
rect 175 53 176 54 
<< pdiffusion >>
rect 176 53 177 54 
<< pdiffusion >>
rect 177 53 178 54 
<< pdiffusion >>
rect 178 53 179 54 
<< pdiffusion >>
rect 179 53 180 54 
<< m1 >>
rect 19 54 20 55 
<< m1 >>
rect 21 54 22 55 
<< m2 >>
rect 21 54 22 55 
<< m2c >>
rect 21 54 22 55 
<< m1 >>
rect 21 54 22 55 
<< m2 >>
rect 21 54 22 55 
<< m2 >>
rect 22 54 23 55 
<< m1 >>
rect 23 54 24 55 
<< m2 >>
rect 23 54 24 55 
<< m2 >>
rect 24 54 25 55 
<< m1 >>
rect 25 54 26 55 
<< m2 >>
rect 25 54 26 55 
<< m2c >>
rect 25 54 26 55 
<< m1 >>
rect 25 54 26 55 
<< m2 >>
rect 25 54 26 55 
<< m1 >>
rect 31 54 32 55 
<< m1 >>
rect 34 54 35 55 
<< m1 >>
rect 37 54 38 55 
<< m2 >>
rect 37 54 38 55 
<< m1 >>
rect 43 54 44 55 
<< m1 >>
rect 46 54 47 55 
<< m1 >>
rect 49 54 50 55 
<< m1 >>
rect 52 54 53 55 
<< m1 >>
rect 55 54 56 55 
<< m2 >>
rect 63 54 64 55 
<< m1 >>
rect 64 54 65 55 
<< m1 >>
rect 73 54 74 55 
<< m1 >>
rect 88 54 89 55 
<< m1 >>
rect 91 54 92 55 
<< m1 >>
rect 93 54 94 55 
<< m1 >>
rect 103 54 104 55 
<< m1 >>
rect 106 54 107 55 
<< m1 >>
rect 109 54 110 55 
<< m1 >>
rect 111 54 112 55 
<< m1 >>
rect 113 54 114 55 
<< m1 >>
rect 121 54 122 55 
<< m1 >>
rect 127 54 128 55 
<< m2 >>
rect 127 54 128 55 
<< m1 >>
rect 139 54 140 55 
<< m1 >>
rect 142 54 143 55 
<< m1 >>
rect 146 54 147 55 
<< m1 >>
rect 148 54 149 55 
<< m1 >>
rect 157 54 158 55 
<< m1 >>
rect 160 54 161 55 
<< m1 >>
rect 163 54 164 55 
<< m2 >>
rect 164 54 165 55 
<< m1 >>
rect 169 54 170 55 
<< m2 >>
rect 169 54 170 55 
<< m1 >>
rect 171 54 172 55 
<< m1 >>
rect 19 55 20 56 
<< m1 >>
rect 21 55 22 56 
<< m1 >>
rect 23 55 24 56 
<< m1 >>
rect 31 55 32 56 
<< m1 >>
rect 34 55 35 56 
<< m1 >>
rect 37 55 38 56 
<< m2 >>
rect 37 55 38 56 
<< m1 >>
rect 43 55 44 56 
<< m1 >>
rect 46 55 47 56 
<< m1 >>
rect 49 55 50 56 
<< m1 >>
rect 52 55 53 56 
<< m1 >>
rect 53 55 54 56 
<< m1 >>
rect 54 55 55 56 
<< m1 >>
rect 55 55 56 56 
<< m2 >>
rect 63 55 64 56 
<< m1 >>
rect 64 55 65 56 
<< m1 >>
rect 73 55 74 56 
<< m1 >>
rect 74 55 75 56 
<< m1 >>
rect 75 55 76 56 
<< m1 >>
rect 76 55 77 56 
<< m1 >>
rect 77 55 78 56 
<< m1 >>
rect 78 55 79 56 
<< m1 >>
rect 79 55 80 56 
<< m1 >>
rect 80 55 81 56 
<< m1 >>
rect 81 55 82 56 
<< m1 >>
rect 82 55 83 56 
<< m1 >>
rect 83 55 84 56 
<< m1 >>
rect 88 55 89 56 
<< m1 >>
rect 89 55 90 56 
<< m1 >>
rect 90 55 91 56 
<< m1 >>
rect 91 55 92 56 
<< m1 >>
rect 93 55 94 56 
<< m1 >>
rect 94 55 95 56 
<< m1 >>
rect 95 55 96 56 
<< m1 >>
rect 96 55 97 56 
<< m1 >>
rect 97 55 98 56 
<< m1 >>
rect 98 55 99 56 
<< m1 >>
rect 99 55 100 56 
<< m1 >>
rect 100 55 101 56 
<< m1 >>
rect 101 55 102 56 
<< m1 >>
rect 102 55 103 56 
<< m1 >>
rect 103 55 104 56 
<< m1 >>
rect 105 55 106 56 
<< m1 >>
rect 106 55 107 56 
<< m1 >>
rect 109 55 110 56 
<< m1 >>
rect 111 55 112 56 
<< m1 >>
rect 113 55 114 56 
<< m1 >>
rect 118 55 119 56 
<< m1 >>
rect 119 55 120 56 
<< m1 >>
rect 120 55 121 56 
<< m1 >>
rect 121 55 122 56 
<< m1 >>
rect 127 55 128 56 
<< m2 >>
rect 127 55 128 56 
<< m1 >>
rect 128 55 129 56 
<< m1 >>
rect 129 55 130 56 
<< m1 >>
rect 130 55 131 56 
<< m1 >>
rect 131 55 132 56 
<< m1 >>
rect 132 55 133 56 
<< m1 >>
rect 133 55 134 56 
<< m1 >>
rect 134 55 135 56 
<< m1 >>
rect 135 55 136 56 
<< m1 >>
rect 136 55 137 56 
<< m1 >>
rect 137 55 138 56 
<< m1 >>
rect 138 55 139 56 
<< m1 >>
rect 139 55 140 56 
<< m1 >>
rect 142 55 143 56 
<< m1 >>
rect 146 55 147 56 
<< m1 >>
rect 148 55 149 56 
<< m1 >>
rect 157 55 158 56 
<< m1 >>
rect 158 55 159 56 
<< m2 >>
rect 158 55 159 56 
<< m2c >>
rect 158 55 159 56 
<< m1 >>
rect 158 55 159 56 
<< m2 >>
rect 158 55 159 56 
<< m2 >>
rect 159 55 160 56 
<< m1 >>
rect 160 55 161 56 
<< m1 >>
rect 163 55 164 56 
<< m2 >>
rect 164 55 165 56 
<< m1 >>
rect 169 55 170 56 
<< m2 >>
rect 169 55 170 56 
<< m1 >>
rect 171 55 172 56 
<< m2 >>
rect 18 56 19 57 
<< m1 >>
rect 19 56 20 57 
<< m2 >>
rect 19 56 20 57 
<< m2 >>
rect 20 56 21 57 
<< m1 >>
rect 21 56 22 57 
<< m2 >>
rect 21 56 22 57 
<< m2c >>
rect 21 56 22 57 
<< m1 >>
rect 21 56 22 57 
<< m2 >>
rect 21 56 22 57 
<< m1 >>
rect 23 56 24 57 
<< m2 >>
rect 23 56 24 57 
<< m2c >>
rect 23 56 24 57 
<< m1 >>
rect 23 56 24 57 
<< m2 >>
rect 23 56 24 57 
<< m1 >>
rect 31 56 32 57 
<< m2 >>
rect 31 56 32 57 
<< m2c >>
rect 31 56 32 57 
<< m1 >>
rect 31 56 32 57 
<< m2 >>
rect 31 56 32 57 
<< m1 >>
rect 34 56 35 57 
<< m1 >>
rect 37 56 38 57 
<< m2 >>
rect 37 56 38 57 
<< m1 >>
rect 43 56 44 57 
<< m1 >>
rect 46 56 47 57 
<< m1 >>
rect 49 56 50 57 
<< m2 >>
rect 63 56 64 57 
<< m1 >>
rect 64 56 65 57 
<< m1 >>
rect 83 56 84 57 
<< m1 >>
rect 105 56 106 57 
<< m1 >>
rect 109 56 110 57 
<< m1 >>
rect 111 56 112 57 
<< m1 >>
rect 113 56 114 57 
<< m1 >>
rect 118 56 119 57 
<< m2 >>
rect 127 56 128 57 
<< m1 >>
rect 142 56 143 57 
<< m1 >>
rect 146 56 147 57 
<< m2 >>
rect 146 56 147 57 
<< m2c >>
rect 146 56 147 57 
<< m1 >>
rect 146 56 147 57 
<< m2 >>
rect 146 56 147 57 
<< m1 >>
rect 148 56 149 57 
<< m2 >>
rect 148 56 149 57 
<< m2c >>
rect 148 56 149 57 
<< m1 >>
rect 148 56 149 57 
<< m2 >>
rect 148 56 149 57 
<< m2 >>
rect 159 56 160 57 
<< m1 >>
rect 160 56 161 57 
<< m2 >>
rect 160 56 161 57 
<< m2 >>
rect 161 56 162 57 
<< m1 >>
rect 162 56 163 57 
<< m2 >>
rect 162 56 163 57 
<< m2c >>
rect 162 56 163 57 
<< m1 >>
rect 162 56 163 57 
<< m2 >>
rect 162 56 163 57 
<< m1 >>
rect 163 56 164 57 
<< m2 >>
rect 164 56 165 57 
<< m1 >>
rect 169 56 170 57 
<< m2 >>
rect 169 56 170 57 
<< m1 >>
rect 171 56 172 57 
<< m2 >>
rect 18 57 19 58 
<< m1 >>
rect 19 57 20 58 
<< m2 >>
rect 23 57 24 58 
<< m2 >>
rect 31 57 32 58 
<< m1 >>
rect 34 57 35 58 
<< m1 >>
rect 37 57 38 58 
<< m2 >>
rect 37 57 38 58 
<< m1 >>
rect 43 57 44 58 
<< m1 >>
rect 46 57 47 58 
<< m1 >>
rect 49 57 50 58 
<< m2 >>
rect 63 57 64 58 
<< m1 >>
rect 64 57 65 58 
<< m1 >>
rect 83 57 84 58 
<< m1 >>
rect 105 57 106 58 
<< m2 >>
rect 105 57 106 58 
<< m2c >>
rect 105 57 106 58 
<< m1 >>
rect 105 57 106 58 
<< m2 >>
rect 105 57 106 58 
<< m1 >>
rect 109 57 110 58 
<< m1 >>
rect 111 57 112 58 
<< m1 >>
rect 113 57 114 58 
<< m1 >>
rect 118 57 119 58 
<< m1 >>
rect 127 57 128 58 
<< m2 >>
rect 127 57 128 58 
<< m2c >>
rect 127 57 128 58 
<< m1 >>
rect 127 57 128 58 
<< m2 >>
rect 127 57 128 58 
<< m1 >>
rect 142 57 143 58 
<< m2 >>
rect 146 57 147 58 
<< m2 >>
rect 148 57 149 58 
<< m1 >>
rect 160 57 161 58 
<< m2 >>
rect 164 57 165 58 
<< m1 >>
rect 169 57 170 58 
<< m2 >>
rect 169 57 170 58 
<< m1 >>
rect 171 57 172 58 
<< m2 >>
rect 18 58 19 59 
<< m1 >>
rect 19 58 20 59 
<< m2 >>
rect 20 58 21 59 
<< m1 >>
rect 21 58 22 59 
<< m2 >>
rect 21 58 22 59 
<< m2c >>
rect 21 58 22 59 
<< m1 >>
rect 21 58 22 59 
<< m2 >>
rect 21 58 22 59 
<< m1 >>
rect 22 58 23 59 
<< m1 >>
rect 23 58 24 59 
<< m2 >>
rect 23 58 24 59 
<< m1 >>
rect 24 58 25 59 
<< m1 >>
rect 25 58 26 59 
<< m1 >>
rect 26 58 27 59 
<< m1 >>
rect 27 58 28 59 
<< m1 >>
rect 28 58 29 59 
<< m1 >>
rect 29 58 30 59 
<< m1 >>
rect 30 58 31 59 
<< m1 >>
rect 31 58 32 59 
<< m2 >>
rect 31 58 32 59 
<< m1 >>
rect 32 58 33 59 
<< m1 >>
rect 33 58 34 59 
<< m1 >>
rect 34 58 35 59 
<< m1 >>
rect 37 58 38 59 
<< m2 >>
rect 37 58 38 59 
<< m1 >>
rect 43 58 44 59 
<< m1 >>
rect 46 58 47 59 
<< m1 >>
rect 49 58 50 59 
<< m2 >>
rect 63 58 64 59 
<< m1 >>
rect 64 58 65 59 
<< m1 >>
rect 83 58 84 59 
<< m2 >>
rect 105 58 106 59 
<< m1 >>
rect 109 58 110 59 
<< m1 >>
rect 111 58 112 59 
<< m1 >>
rect 113 58 114 59 
<< m1 >>
rect 118 58 119 59 
<< m1 >>
rect 127 58 128 59 
<< m1 >>
rect 128 58 129 59 
<< m1 >>
rect 129 58 130 59 
<< m1 >>
rect 130 58 131 59 
<< m1 >>
rect 131 58 132 59 
<< m1 >>
rect 132 58 133 59 
<< m1 >>
rect 133 58 134 59 
<< m1 >>
rect 134 58 135 59 
<< m1 >>
rect 135 58 136 59 
<< m1 >>
rect 136 58 137 59 
<< m1 >>
rect 137 58 138 59 
<< m1 >>
rect 138 58 139 59 
<< m1 >>
rect 139 58 140 59 
<< m1 >>
rect 140 58 141 59 
<< m1 >>
rect 141 58 142 59 
<< m1 >>
rect 142 58 143 59 
<< m2 >>
rect 143 58 144 59 
<< m1 >>
rect 144 58 145 59 
<< m2 >>
rect 144 58 145 59 
<< m2c >>
rect 144 58 145 59 
<< m1 >>
rect 144 58 145 59 
<< m2 >>
rect 144 58 145 59 
<< m1 >>
rect 145 58 146 59 
<< m1 >>
rect 146 58 147 59 
<< m2 >>
rect 146 58 147 59 
<< m1 >>
rect 147 58 148 59 
<< m1 >>
rect 148 58 149 59 
<< m2 >>
rect 148 58 149 59 
<< m1 >>
rect 149 58 150 59 
<< m1 >>
rect 150 58 151 59 
<< m1 >>
rect 151 58 152 59 
<< m1 >>
rect 152 58 153 59 
<< m1 >>
rect 153 58 154 59 
<< m1 >>
rect 154 58 155 59 
<< m1 >>
rect 155 58 156 59 
<< m1 >>
rect 156 58 157 59 
<< m1 >>
rect 157 58 158 59 
<< m1 >>
rect 158 58 159 59 
<< m1 >>
rect 159 58 160 59 
<< m1 >>
rect 160 58 161 59 
<< m1 >>
rect 164 58 165 59 
<< m2 >>
rect 164 58 165 59 
<< m2c >>
rect 164 58 165 59 
<< m1 >>
rect 164 58 165 59 
<< m2 >>
rect 164 58 165 59 
<< m1 >>
rect 169 58 170 59 
<< m2 >>
rect 169 58 170 59 
<< m1 >>
rect 171 58 172 59 
<< m2 >>
rect 18 59 19 60 
<< m1 >>
rect 19 59 20 60 
<< m2 >>
rect 20 59 21 60 
<< m2 >>
rect 23 59 24 60 
<< m2 >>
rect 31 59 32 60 
<< m1 >>
rect 37 59 38 60 
<< m2 >>
rect 37 59 38 60 
<< m1 >>
rect 43 59 44 60 
<< m1 >>
rect 46 59 47 60 
<< m1 >>
rect 49 59 50 60 
<< m2 >>
rect 49 59 50 60 
<< m2c >>
rect 49 59 50 60 
<< m1 >>
rect 49 59 50 60 
<< m2 >>
rect 49 59 50 60 
<< m2 >>
rect 63 59 64 60 
<< m1 >>
rect 64 59 65 60 
<< m1 >>
rect 83 59 84 60 
<< m2 >>
rect 83 59 84 60 
<< m2c >>
rect 83 59 84 60 
<< m1 >>
rect 83 59 84 60 
<< m2 >>
rect 83 59 84 60 
<< m1 >>
rect 100 59 101 60 
<< m1 >>
rect 101 59 102 60 
<< m1 >>
rect 102 59 103 60 
<< m1 >>
rect 103 59 104 60 
<< m1 >>
rect 104 59 105 60 
<< m1 >>
rect 105 59 106 60 
<< m2 >>
rect 105 59 106 60 
<< m1 >>
rect 106 59 107 60 
<< m1 >>
rect 107 59 108 60 
<< m2 >>
rect 107 59 108 60 
<< m2c >>
rect 107 59 108 60 
<< m1 >>
rect 107 59 108 60 
<< m2 >>
rect 107 59 108 60 
<< m2 >>
rect 108 59 109 60 
<< m1 >>
rect 109 59 110 60 
<< m2 >>
rect 109 59 110 60 
<< m2 >>
rect 110 59 111 60 
<< m1 >>
rect 111 59 112 60 
<< m2 >>
rect 111 59 112 60 
<< m2 >>
rect 112 59 113 60 
<< m1 >>
rect 113 59 114 60 
<< m2 >>
rect 113 59 114 60 
<< m2 >>
rect 114 59 115 60 
<< m1 >>
rect 115 59 116 60 
<< m2 >>
rect 115 59 116 60 
<< m1 >>
rect 116 59 117 60 
<< m2 >>
rect 116 59 117 60 
<< m2c >>
rect 116 59 117 60 
<< m1 >>
rect 116 59 117 60 
<< m2 >>
rect 116 59 117 60 
<< m2 >>
rect 117 59 118 60 
<< m1 >>
rect 118 59 119 60 
<< m2 >>
rect 118 59 119 60 
<< m2 >>
rect 119 59 120 60 
<< m1 >>
rect 120 59 121 60 
<< m2 >>
rect 120 59 121 60 
<< m2c >>
rect 120 59 121 60 
<< m1 >>
rect 120 59 121 60 
<< m2 >>
rect 120 59 121 60 
<< m1 >>
rect 121 59 122 60 
<< m1 >>
rect 122 59 123 60 
<< m1 >>
rect 123 59 124 60 
<< m1 >>
rect 124 59 125 60 
<< m1 >>
rect 125 59 126 60 
<< m2 >>
rect 125 59 126 60 
<< m2c >>
rect 125 59 126 60 
<< m1 >>
rect 125 59 126 60 
<< m2 >>
rect 125 59 126 60 
<< m2 >>
rect 126 59 127 60 
<< m2 >>
rect 127 59 128 60 
<< m2 >>
rect 128 59 129 60 
<< m2 >>
rect 129 59 130 60 
<< m2 >>
rect 130 59 131 60 
<< m2 >>
rect 131 59 132 60 
<< m2 >>
rect 132 59 133 60 
<< m2 >>
rect 133 59 134 60 
<< m2 >>
rect 134 59 135 60 
<< m2 >>
rect 135 59 136 60 
<< m2 >>
rect 136 59 137 60 
<< m2 >>
rect 137 59 138 60 
<< m2 >>
rect 138 59 139 60 
<< m2 >>
rect 139 59 140 60 
<< m2 >>
rect 140 59 141 60 
<< m2 >>
rect 141 59 142 60 
<< m2 >>
rect 142 59 143 60 
<< m2 >>
rect 143 59 144 60 
<< m2 >>
rect 146 59 147 60 
<< m2 >>
rect 148 59 149 60 
<< m1 >>
rect 164 59 165 60 
<< m1 >>
rect 169 59 170 60 
<< m2 >>
rect 169 59 170 60 
<< m1 >>
rect 171 59 172 60 
<< m2 >>
rect 18 60 19 61 
<< m1 >>
rect 19 60 20 61 
<< m2 >>
rect 20 60 21 61 
<< m1 >>
rect 23 60 24 61 
<< m2 >>
rect 23 60 24 61 
<< m2c >>
rect 23 60 24 61 
<< m1 >>
rect 23 60 24 61 
<< m2 >>
rect 23 60 24 61 
<< m1 >>
rect 30 60 31 61 
<< m1 >>
rect 31 60 32 61 
<< m2 >>
rect 31 60 32 61 
<< m2c >>
rect 31 60 32 61 
<< m1 >>
rect 31 60 32 61 
<< m2 >>
rect 31 60 32 61 
<< m1 >>
rect 37 60 38 61 
<< m2 >>
rect 37 60 38 61 
<< m1 >>
rect 43 60 44 61 
<< m1 >>
rect 46 60 47 61 
<< m2 >>
rect 48 60 49 61 
<< m2 >>
rect 49 60 50 61 
<< m2 >>
rect 63 60 64 61 
<< m1 >>
rect 64 60 65 61 
<< m2 >>
rect 83 60 84 61 
<< m2 >>
rect 84 60 85 61 
<< m2 >>
rect 85 60 86 61 
<< m2 >>
rect 86 60 87 61 
<< m1 >>
rect 100 60 101 61 
<< m2 >>
rect 105 60 106 61 
<< m1 >>
rect 109 60 110 61 
<< m1 >>
rect 111 60 112 61 
<< m1 >>
rect 113 60 114 61 
<< m1 >>
rect 118 60 119 61 
<< m1 >>
rect 146 60 147 61 
<< m2 >>
rect 146 60 147 61 
<< m2c >>
rect 146 60 147 61 
<< m1 >>
rect 146 60 147 61 
<< m2 >>
rect 146 60 147 61 
<< m1 >>
rect 148 60 149 61 
<< m2 >>
rect 148 60 149 61 
<< m2c >>
rect 148 60 149 61 
<< m1 >>
rect 148 60 149 61 
<< m2 >>
rect 148 60 149 61 
<< m1 >>
rect 164 60 165 61 
<< m1 >>
rect 169 60 170 61 
<< m2 >>
rect 169 60 170 61 
<< m1 >>
rect 171 60 172 61 
<< m1 >>
rect 10 61 11 62 
<< m1 >>
rect 11 61 12 62 
<< m1 >>
rect 12 61 13 62 
<< m1 >>
rect 13 61 14 62 
<< m1 >>
rect 14 61 15 62 
<< m1 >>
rect 15 61 16 62 
<< m1 >>
rect 16 61 17 62 
<< m1 >>
rect 17 61 18 62 
<< m2 >>
rect 17 61 18 62 
<< m2c >>
rect 17 61 18 62 
<< m1 >>
rect 17 61 18 62 
<< m2 >>
rect 17 61 18 62 
<< m2 >>
rect 18 61 19 62 
<< m1 >>
rect 19 61 20 62 
<< m2 >>
rect 20 61 21 62 
<< m1 >>
rect 23 61 24 62 
<< m1 >>
rect 30 61 31 62 
<< m1 >>
rect 37 61 38 62 
<< m2 >>
rect 37 61 38 62 
<< m1 >>
rect 43 61 44 62 
<< m1 >>
rect 46 61 47 62 
<< m1 >>
rect 47 61 48 62 
<< m1 >>
rect 48 61 49 62 
<< m2 >>
rect 48 61 49 62 
<< m1 >>
rect 49 61 50 62 
<< m1 >>
rect 50 61 51 62 
<< m1 >>
rect 51 61 52 62 
<< m1 >>
rect 52 61 53 62 
<< m2 >>
rect 63 61 64 62 
<< m1 >>
rect 64 61 65 62 
<< m1 >>
rect 84 61 85 62 
<< m1 >>
rect 85 61 86 62 
<< m1 >>
rect 86 61 87 62 
<< m2 >>
rect 86 61 87 62 
<< m1 >>
rect 87 61 88 62 
<< m2 >>
rect 87 61 88 62 
<< m1 >>
rect 88 61 89 62 
<< m2 >>
rect 88 61 89 62 
<< m1 >>
rect 89 61 90 62 
<< m2 >>
rect 89 61 90 62 
<< m1 >>
rect 90 61 91 62 
<< m2 >>
rect 90 61 91 62 
<< m1 >>
rect 91 61 92 62 
<< m2 >>
rect 91 61 92 62 
<< m1 >>
rect 92 61 93 62 
<< m2 >>
rect 92 61 93 62 
<< m1 >>
rect 93 61 94 62 
<< m2 >>
rect 93 61 94 62 
<< m1 >>
rect 94 61 95 62 
<< m2 >>
rect 94 61 95 62 
<< m1 >>
rect 95 61 96 62 
<< m2 >>
rect 95 61 96 62 
<< m1 >>
rect 96 61 97 62 
<< m2 >>
rect 96 61 97 62 
<< m1 >>
rect 97 61 98 62 
<< m2 >>
rect 97 61 98 62 
<< m1 >>
rect 98 61 99 62 
<< m2 >>
rect 98 61 99 62 
<< m2 >>
rect 99 61 100 62 
<< m1 >>
rect 100 61 101 62 
<< m2 >>
rect 100 61 101 62 
<< m2 >>
rect 101 61 102 62 
<< m1 >>
rect 102 61 103 62 
<< m2 >>
rect 102 61 103 62 
<< m2c >>
rect 102 61 103 62 
<< m1 >>
rect 102 61 103 62 
<< m2 >>
rect 102 61 103 62 
<< m1 >>
rect 103 61 104 62 
<< m1 >>
rect 105 61 106 62 
<< m2 >>
rect 105 61 106 62 
<< m2c >>
rect 105 61 106 62 
<< m1 >>
rect 105 61 106 62 
<< m2 >>
rect 105 61 106 62 
<< m1 >>
rect 106 61 107 62 
<< m1 >>
rect 107 61 108 62 
<< m2 >>
rect 107 61 108 62 
<< m2c >>
rect 107 61 108 62 
<< m1 >>
rect 107 61 108 62 
<< m2 >>
rect 107 61 108 62 
<< m2 >>
rect 108 61 109 62 
<< m1 >>
rect 109 61 110 62 
<< m2 >>
rect 109 61 110 62 
<< m2 >>
rect 110 61 111 62 
<< m1 >>
rect 111 61 112 62 
<< m2 >>
rect 111 61 112 62 
<< m2 >>
rect 112 61 113 62 
<< m1 >>
rect 113 61 114 62 
<< m2 >>
rect 113 61 114 62 
<< m2 >>
rect 114 61 115 62 
<< m1 >>
rect 115 61 116 62 
<< m2 >>
rect 115 61 116 62 
<< m2c >>
rect 115 61 116 62 
<< m1 >>
rect 115 61 116 62 
<< m2 >>
rect 115 61 116 62 
<< m1 >>
rect 118 61 119 62 
<< m1 >>
rect 124 61 125 62 
<< m1 >>
rect 125 61 126 62 
<< m1 >>
rect 126 61 127 62 
<< m1 >>
rect 127 61 128 62 
<< m1 >>
rect 128 61 129 62 
<< m1 >>
rect 129 61 130 62 
<< m1 >>
rect 130 61 131 62 
<< m1 >>
rect 131 61 132 62 
<< m1 >>
rect 132 61 133 62 
<< m1 >>
rect 133 61 134 62 
<< m1 >>
rect 134 61 135 62 
<< m1 >>
rect 135 61 136 62 
<< m1 >>
rect 136 61 137 62 
<< m1 >>
rect 137 61 138 62 
<< m1 >>
rect 138 61 139 62 
<< m1 >>
rect 139 61 140 62 
<< m1 >>
rect 140 61 141 62 
<< m1 >>
rect 141 61 142 62 
<< m1 >>
rect 142 61 143 62 
<< m1 >>
rect 143 61 144 62 
<< m1 >>
rect 144 61 145 62 
<< m1 >>
rect 146 61 147 62 
<< m1 >>
rect 148 61 149 62 
<< m1 >>
rect 154 61 155 62 
<< m1 >>
rect 155 61 156 62 
<< m1 >>
rect 156 61 157 62 
<< m1 >>
rect 157 61 158 62 
<< m1 >>
rect 158 61 159 62 
<< m1 >>
rect 159 61 160 62 
<< m1 >>
rect 160 61 161 62 
<< m1 >>
rect 164 61 165 62 
<< m1 >>
rect 169 61 170 62 
<< m2 >>
rect 169 61 170 62 
<< m1 >>
rect 171 61 172 62 
<< m1 >>
rect 10 62 11 63 
<< m1 >>
rect 19 62 20 63 
<< m2 >>
rect 20 62 21 63 
<< m2 >>
rect 22 62 23 63 
<< m1 >>
rect 23 62 24 63 
<< m2 >>
rect 23 62 24 63 
<< m2 >>
rect 24 62 25 63 
<< m1 >>
rect 25 62 26 63 
<< m2 >>
rect 25 62 26 63 
<< m2c >>
rect 25 62 26 63 
<< m1 >>
rect 25 62 26 63 
<< m2 >>
rect 25 62 26 63 
<< m1 >>
rect 26 62 27 63 
<< m1 >>
rect 27 62 28 63 
<< m1 >>
rect 28 62 29 63 
<< m1 >>
rect 29 62 30 63 
<< m1 >>
rect 30 62 31 63 
<< m1 >>
rect 37 62 38 63 
<< m2 >>
rect 37 62 38 63 
<< m1 >>
rect 43 62 44 63 
<< m2 >>
rect 48 62 49 63 
<< m1 >>
rect 52 62 53 63 
<< m2 >>
rect 63 62 64 63 
<< m1 >>
rect 64 62 65 63 
<< m1 >>
rect 84 62 85 63 
<< m2 >>
rect 84 62 85 63 
<< m2c >>
rect 84 62 85 63 
<< m1 >>
rect 84 62 85 63 
<< m2 >>
rect 84 62 85 63 
<< m1 >>
rect 98 62 99 63 
<< m1 >>
rect 100 62 101 63 
<< m1 >>
rect 103 62 104 63 
<< m1 >>
rect 109 62 110 63 
<< m1 >>
rect 111 62 112 63 
<< m1 >>
rect 113 62 114 63 
<< m1 >>
rect 115 62 116 63 
<< m1 >>
rect 118 62 119 63 
<< m1 >>
rect 124 62 125 63 
<< m1 >>
rect 144 62 145 63 
<< m2 >>
rect 144 62 145 63 
<< m2c >>
rect 144 62 145 63 
<< m1 >>
rect 144 62 145 63 
<< m2 >>
rect 144 62 145 63 
<< m2 >>
rect 145 62 146 63 
<< m1 >>
rect 146 62 147 63 
<< m2 >>
rect 146 62 147 63 
<< m2 >>
rect 147 62 148 63 
<< m1 >>
rect 148 62 149 63 
<< m2 >>
rect 148 62 149 63 
<< m2c >>
rect 148 62 149 63 
<< m1 >>
rect 148 62 149 63 
<< m2 >>
rect 148 62 149 63 
<< m1 >>
rect 154 62 155 63 
<< m1 >>
rect 160 62 161 63 
<< m1 >>
rect 164 62 165 63 
<< m1 >>
rect 169 62 170 63 
<< m2 >>
rect 169 62 170 63 
<< m1 >>
rect 171 62 172 63 
<< m1 >>
rect 10 63 11 64 
<< m1 >>
rect 19 63 20 64 
<< m2 >>
rect 20 63 21 64 
<< m2 >>
rect 22 63 23 64 
<< m1 >>
rect 23 63 24 64 
<< m1 >>
rect 37 63 38 64 
<< m2 >>
rect 37 63 38 64 
<< m1 >>
rect 43 63 44 64 
<< m1 >>
rect 46 63 47 64 
<< m1 >>
rect 47 63 48 64 
<< m1 >>
rect 48 63 49 64 
<< m2 >>
rect 48 63 49 64 
<< m2c >>
rect 48 63 49 64 
<< m1 >>
rect 48 63 49 64 
<< m2 >>
rect 48 63 49 64 
<< m1 >>
rect 52 63 53 64 
<< m2 >>
rect 63 63 64 64 
<< m1 >>
rect 64 63 65 64 
<< m2 >>
rect 82 63 83 64 
<< m2 >>
rect 83 63 84 64 
<< m2 >>
rect 84 63 85 64 
<< m1 >>
rect 98 63 99 64 
<< m1 >>
rect 100 63 101 64 
<< m1 >>
rect 103 63 104 64 
<< m1 >>
rect 109 63 110 64 
<< m1 >>
rect 111 63 112 64 
<< m1 >>
rect 113 63 114 64 
<< m1 >>
rect 115 63 116 64 
<< m1 >>
rect 118 63 119 64 
<< m1 >>
rect 124 63 125 64 
<< m1 >>
rect 146 63 147 64 
<< m1 >>
rect 154 63 155 64 
<< m1 >>
rect 160 63 161 64 
<< m1 >>
rect 164 63 165 64 
<< m1 >>
rect 169 63 170 64 
<< m2 >>
rect 169 63 170 64 
<< m1 >>
rect 171 63 172 64 
<< m1 >>
rect 10 64 11 65 
<< m1 >>
rect 19 64 20 65 
<< m2 >>
rect 20 64 21 65 
<< m2 >>
rect 22 64 23 65 
<< m1 >>
rect 23 64 24 65 
<< m1 >>
rect 28 64 29 65 
<< m1 >>
rect 29 64 30 65 
<< m1 >>
rect 30 64 31 65 
<< m1 >>
rect 31 64 32 65 
<< m1 >>
rect 34 64 35 65 
<< m1 >>
rect 35 64 36 65 
<< m2 >>
rect 35 64 36 65 
<< m2c >>
rect 35 64 36 65 
<< m1 >>
rect 35 64 36 65 
<< m2 >>
rect 35 64 36 65 
<< m2 >>
rect 36 64 37 65 
<< m1 >>
rect 37 64 38 65 
<< m2 >>
rect 37 64 38 65 
<< m1 >>
rect 43 64 44 65 
<< m1 >>
rect 46 64 47 65 
<< m1 >>
rect 52 64 53 65 
<< m2 >>
rect 63 64 64 65 
<< m1 >>
rect 64 64 65 65 
<< m1 >>
rect 65 64 66 65 
<< m1 >>
rect 66 64 67 65 
<< m1 >>
rect 67 64 68 65 
<< m1 >>
rect 70 64 71 65 
<< m1 >>
rect 71 64 72 65 
<< m1 >>
rect 72 64 73 65 
<< m1 >>
rect 73 64 74 65 
<< m1 >>
rect 82 64 83 65 
<< m2 >>
rect 82 64 83 65 
<< m1 >>
rect 83 64 84 65 
<< m1 >>
rect 84 64 85 65 
<< m1 >>
rect 85 64 86 65 
<< m1 >>
rect 98 64 99 65 
<< m1 >>
rect 100 64 101 65 
<< m1 >>
rect 103 64 104 65 
<< m1 >>
rect 106 64 107 65 
<< m1 >>
rect 107 64 108 65 
<< m2 >>
rect 107 64 108 65 
<< m2c >>
rect 107 64 108 65 
<< m1 >>
rect 107 64 108 65 
<< m2 >>
rect 107 64 108 65 
<< m2 >>
rect 108 64 109 65 
<< m1 >>
rect 109 64 110 65 
<< m2 >>
rect 109 64 110 65 
<< m2 >>
rect 110 64 111 65 
<< m1 >>
rect 111 64 112 65 
<< m2 >>
rect 111 64 112 65 
<< m2 >>
rect 112 64 113 65 
<< m1 >>
rect 113 64 114 65 
<< m2 >>
rect 113 64 114 65 
<< m2 >>
rect 114 64 115 65 
<< m1 >>
rect 115 64 116 65 
<< m2 >>
rect 115 64 116 65 
<< m2 >>
rect 116 64 117 65 
<< m2 >>
rect 117 64 118 65 
<< m1 >>
rect 118 64 119 65 
<< m2 >>
rect 118 64 119 65 
<< m1 >>
rect 124 64 125 65 
<< m1 >>
rect 146 64 147 65 
<< m1 >>
rect 154 64 155 65 
<< m1 >>
rect 160 64 161 65 
<< m1 >>
rect 164 64 165 65 
<< m1 >>
rect 169 64 170 65 
<< m2 >>
rect 169 64 170 65 
<< m1 >>
rect 171 64 172 65 
<< m1 >>
rect 10 65 11 66 
<< m1 >>
rect 19 65 20 66 
<< m2 >>
rect 20 65 21 66 
<< m2 >>
rect 22 65 23 66 
<< m1 >>
rect 23 65 24 66 
<< m1 >>
rect 28 65 29 66 
<< m1 >>
rect 31 65 32 66 
<< m1 >>
rect 34 65 35 66 
<< m1 >>
rect 37 65 38 66 
<< m1 >>
rect 43 65 44 66 
<< m1 >>
rect 46 65 47 66 
<< m1 >>
rect 52 65 53 66 
<< m2 >>
rect 63 65 64 66 
<< m1 >>
rect 67 65 68 66 
<< m1 >>
rect 70 65 71 66 
<< m1 >>
rect 73 65 74 66 
<< m1 >>
rect 82 65 83 66 
<< m2 >>
rect 82 65 83 66 
<< m1 >>
rect 85 65 86 66 
<< m1 >>
rect 98 65 99 66 
<< m1 >>
rect 100 65 101 66 
<< m1 >>
rect 103 65 104 66 
<< m1 >>
rect 106 65 107 66 
<< m1 >>
rect 109 65 110 66 
<< m1 >>
rect 111 65 112 66 
<< m1 >>
rect 113 65 114 66 
<< m1 >>
rect 115 65 116 66 
<< m1 >>
rect 118 65 119 66 
<< m2 >>
rect 118 65 119 66 
<< m1 >>
rect 124 65 125 66 
<< m1 >>
rect 146 65 147 66 
<< m1 >>
rect 154 65 155 66 
<< m1 >>
rect 160 65 161 66 
<< m1 >>
rect 164 65 165 66 
<< m1 >>
rect 169 65 170 66 
<< m2 >>
rect 169 65 170 66 
<< m1 >>
rect 171 65 172 66 
<< m1 >>
rect 10 66 11 67 
<< pdiffusion >>
rect 12 66 13 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< m1 >>
rect 19 66 20 67 
<< m2 >>
rect 20 66 21 67 
<< m2 >>
rect 22 66 23 67 
<< m1 >>
rect 23 66 24 67 
<< m1 >>
rect 28 66 29 67 
<< pdiffusion >>
rect 30 66 31 67 
<< m1 >>
rect 31 66 32 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< m1 >>
rect 34 66 35 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< m1 >>
rect 37 66 38 67 
<< m1 >>
rect 43 66 44 67 
<< m1 >>
rect 46 66 47 67 
<< pdiffusion >>
rect 48 66 49 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< m1 >>
rect 52 66 53 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 63 66 64 67 
<< m2 >>
rect 63 66 64 67 
<< m2c >>
rect 63 66 64 67 
<< m1 >>
rect 63 66 64 67 
<< m2 >>
rect 63 66 64 67 
<< pdiffusion >>
rect 66 66 67 67 
<< m1 >>
rect 67 66 68 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< m1 >>
rect 70 66 71 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< m1 >>
rect 73 66 74 67 
<< m1 >>
rect 82 66 83 67 
<< m2 >>
rect 82 66 83 67 
<< pdiffusion >>
rect 84 66 85 67 
<< m1 >>
rect 85 66 86 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< m1 >>
rect 98 66 99 67 
<< m1 >>
rect 100 66 101 67 
<< pdiffusion >>
rect 102 66 103 67 
<< m1 >>
rect 103 66 104 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< m1 >>
rect 106 66 107 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< m1 >>
rect 109 66 110 67 
<< m1 >>
rect 111 66 112 67 
<< m1 >>
rect 113 66 114 67 
<< m1 >>
rect 115 66 116 67 
<< m1 >>
rect 118 66 119 67 
<< m2 >>
rect 118 66 119 67 
<< pdiffusion >>
rect 120 66 121 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< m1 >>
rect 124 66 125 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< pdiffusion >>
rect 138 66 139 67 
<< pdiffusion >>
rect 139 66 140 67 
<< pdiffusion >>
rect 140 66 141 67 
<< pdiffusion >>
rect 141 66 142 67 
<< pdiffusion >>
rect 142 66 143 67 
<< pdiffusion >>
rect 143 66 144 67 
<< m1 >>
rect 146 66 147 67 
<< m1 >>
rect 154 66 155 67 
<< pdiffusion >>
rect 156 66 157 67 
<< pdiffusion >>
rect 157 66 158 67 
<< pdiffusion >>
rect 158 66 159 67 
<< pdiffusion >>
rect 159 66 160 67 
<< m1 >>
rect 160 66 161 67 
<< pdiffusion >>
rect 160 66 161 67 
<< pdiffusion >>
rect 161 66 162 67 
<< m1 >>
rect 164 66 165 67 
<< m1 >>
rect 169 66 170 67 
<< m2 >>
rect 169 66 170 67 
<< m1 >>
rect 171 66 172 67 
<< pdiffusion >>
rect 174 66 175 67 
<< pdiffusion >>
rect 175 66 176 67 
<< pdiffusion >>
rect 176 66 177 67 
<< pdiffusion >>
rect 177 66 178 67 
<< pdiffusion >>
rect 178 66 179 67 
<< pdiffusion >>
rect 179 66 180 67 
<< m1 >>
rect 10 67 11 68 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< m1 >>
rect 19 67 20 68 
<< m2 >>
rect 20 67 21 68 
<< m2 >>
rect 22 67 23 68 
<< m1 >>
rect 23 67 24 68 
<< m1 >>
rect 28 67 29 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< m1 >>
rect 37 67 38 68 
<< m1 >>
rect 43 67 44 68 
<< m1 >>
rect 46 67 47 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 63 67 64 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< m1 >>
rect 73 67 74 68 
<< m1 >>
rect 82 67 83 68 
<< m2 >>
rect 82 67 83 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< m1 >>
rect 98 67 99 68 
<< m1 >>
rect 100 67 101 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< m1 >>
rect 109 67 110 68 
<< m1 >>
rect 111 67 112 68 
<< m1 >>
rect 113 67 114 68 
<< m1 >>
rect 115 67 116 68 
<< m1 >>
rect 118 67 119 68 
<< m2 >>
rect 118 67 119 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< pdiffusion >>
rect 138 67 139 68 
<< pdiffusion >>
rect 139 67 140 68 
<< pdiffusion >>
rect 140 67 141 68 
<< pdiffusion >>
rect 141 67 142 68 
<< pdiffusion >>
rect 142 67 143 68 
<< pdiffusion >>
rect 143 67 144 68 
<< m1 >>
rect 146 67 147 68 
<< m1 >>
rect 154 67 155 68 
<< pdiffusion >>
rect 156 67 157 68 
<< pdiffusion >>
rect 157 67 158 68 
<< pdiffusion >>
rect 158 67 159 68 
<< pdiffusion >>
rect 159 67 160 68 
<< pdiffusion >>
rect 160 67 161 68 
<< pdiffusion >>
rect 161 67 162 68 
<< m1 >>
rect 164 67 165 68 
<< m1 >>
rect 169 67 170 68 
<< m2 >>
rect 169 67 170 68 
<< m1 >>
rect 171 67 172 68 
<< pdiffusion >>
rect 174 67 175 68 
<< pdiffusion >>
rect 175 67 176 68 
<< pdiffusion >>
rect 176 67 177 68 
<< pdiffusion >>
rect 177 67 178 68 
<< pdiffusion >>
rect 178 67 179 68 
<< pdiffusion >>
rect 179 67 180 68 
<< m1 >>
rect 10 68 11 69 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< m1 >>
rect 19 68 20 69 
<< m2 >>
rect 20 68 21 69 
<< m2 >>
rect 22 68 23 69 
<< m1 >>
rect 23 68 24 69 
<< m1 >>
rect 28 68 29 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< m1 >>
rect 37 68 38 69 
<< m1 >>
rect 43 68 44 69 
<< m1 >>
rect 46 68 47 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 63 68 64 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< m1 >>
rect 73 68 74 69 
<< m1 >>
rect 82 68 83 69 
<< m2 >>
rect 82 68 83 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< m1 >>
rect 98 68 99 69 
<< m1 >>
rect 100 68 101 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< m1 >>
rect 109 68 110 69 
<< m1 >>
rect 111 68 112 69 
<< m1 >>
rect 113 68 114 69 
<< m1 >>
rect 115 68 116 69 
<< m1 >>
rect 118 68 119 69 
<< m2 >>
rect 118 68 119 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< pdiffusion >>
rect 138 68 139 69 
<< pdiffusion >>
rect 139 68 140 69 
<< pdiffusion >>
rect 140 68 141 69 
<< pdiffusion >>
rect 141 68 142 69 
<< pdiffusion >>
rect 142 68 143 69 
<< pdiffusion >>
rect 143 68 144 69 
<< m1 >>
rect 146 68 147 69 
<< m1 >>
rect 154 68 155 69 
<< pdiffusion >>
rect 156 68 157 69 
<< pdiffusion >>
rect 157 68 158 69 
<< pdiffusion >>
rect 158 68 159 69 
<< pdiffusion >>
rect 159 68 160 69 
<< pdiffusion >>
rect 160 68 161 69 
<< pdiffusion >>
rect 161 68 162 69 
<< m1 >>
rect 164 68 165 69 
<< m1 >>
rect 169 68 170 69 
<< m2 >>
rect 169 68 170 69 
<< m1 >>
rect 171 68 172 69 
<< pdiffusion >>
rect 174 68 175 69 
<< pdiffusion >>
rect 175 68 176 69 
<< pdiffusion >>
rect 176 68 177 69 
<< pdiffusion >>
rect 177 68 178 69 
<< pdiffusion >>
rect 178 68 179 69 
<< pdiffusion >>
rect 179 68 180 69 
<< m1 >>
rect 10 69 11 70 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< m1 >>
rect 19 69 20 70 
<< m2 >>
rect 20 69 21 70 
<< m2 >>
rect 22 69 23 70 
<< m1 >>
rect 23 69 24 70 
<< m1 >>
rect 28 69 29 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< m1 >>
rect 37 69 38 70 
<< m1 >>
rect 43 69 44 70 
<< m1 >>
rect 46 69 47 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 63 69 64 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< m1 >>
rect 73 69 74 70 
<< m1 >>
rect 82 69 83 70 
<< m2 >>
rect 82 69 83 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< m1 >>
rect 98 69 99 70 
<< m1 >>
rect 100 69 101 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< m1 >>
rect 109 69 110 70 
<< m1 >>
rect 111 69 112 70 
<< m1 >>
rect 113 69 114 70 
<< m1 >>
rect 115 69 116 70 
<< m1 >>
rect 118 69 119 70 
<< m2 >>
rect 118 69 119 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< pdiffusion >>
rect 138 69 139 70 
<< pdiffusion >>
rect 139 69 140 70 
<< pdiffusion >>
rect 140 69 141 70 
<< pdiffusion >>
rect 141 69 142 70 
<< pdiffusion >>
rect 142 69 143 70 
<< pdiffusion >>
rect 143 69 144 70 
<< m1 >>
rect 146 69 147 70 
<< m1 >>
rect 154 69 155 70 
<< pdiffusion >>
rect 156 69 157 70 
<< pdiffusion >>
rect 157 69 158 70 
<< pdiffusion >>
rect 158 69 159 70 
<< pdiffusion >>
rect 159 69 160 70 
<< pdiffusion >>
rect 160 69 161 70 
<< pdiffusion >>
rect 161 69 162 70 
<< m1 >>
rect 164 69 165 70 
<< m1 >>
rect 169 69 170 70 
<< m2 >>
rect 169 69 170 70 
<< m1 >>
rect 171 69 172 70 
<< pdiffusion >>
rect 174 69 175 70 
<< pdiffusion >>
rect 175 69 176 70 
<< pdiffusion >>
rect 176 69 177 70 
<< pdiffusion >>
rect 177 69 178 70 
<< pdiffusion >>
rect 178 69 179 70 
<< pdiffusion >>
rect 179 69 180 70 
<< m1 >>
rect 10 70 11 71 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< m1 >>
rect 19 70 20 71 
<< m2 >>
rect 20 70 21 71 
<< m2 >>
rect 22 70 23 71 
<< m1 >>
rect 23 70 24 71 
<< m1 >>
rect 28 70 29 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< m1 >>
rect 37 70 38 71 
<< m1 >>
rect 43 70 44 71 
<< m1 >>
rect 46 70 47 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 63 70 64 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< m1 >>
rect 73 70 74 71 
<< m1 >>
rect 82 70 83 71 
<< m2 >>
rect 82 70 83 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< m1 >>
rect 98 70 99 71 
<< m1 >>
rect 100 70 101 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< m1 >>
rect 109 70 110 71 
<< m1 >>
rect 111 70 112 71 
<< m1 >>
rect 113 70 114 71 
<< m1 >>
rect 115 70 116 71 
<< m1 >>
rect 118 70 119 71 
<< m2 >>
rect 118 70 119 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< pdiffusion >>
rect 138 70 139 71 
<< pdiffusion >>
rect 139 70 140 71 
<< pdiffusion >>
rect 140 70 141 71 
<< pdiffusion >>
rect 141 70 142 71 
<< pdiffusion >>
rect 142 70 143 71 
<< pdiffusion >>
rect 143 70 144 71 
<< m1 >>
rect 146 70 147 71 
<< m1 >>
rect 154 70 155 71 
<< pdiffusion >>
rect 156 70 157 71 
<< pdiffusion >>
rect 157 70 158 71 
<< pdiffusion >>
rect 158 70 159 71 
<< pdiffusion >>
rect 159 70 160 71 
<< pdiffusion >>
rect 160 70 161 71 
<< pdiffusion >>
rect 161 70 162 71 
<< m1 >>
rect 164 70 165 71 
<< m1 >>
rect 169 70 170 71 
<< m2 >>
rect 169 70 170 71 
<< m1 >>
rect 171 70 172 71 
<< pdiffusion >>
rect 174 70 175 71 
<< pdiffusion >>
rect 175 70 176 71 
<< pdiffusion >>
rect 176 70 177 71 
<< pdiffusion >>
rect 177 70 178 71 
<< pdiffusion >>
rect 178 70 179 71 
<< pdiffusion >>
rect 179 70 180 71 
<< m1 >>
rect 10 71 11 72 
<< pdiffusion >>
rect 12 71 13 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< m1 >>
rect 19 71 20 72 
<< m2 >>
rect 20 71 21 72 
<< m2 >>
rect 22 71 23 72 
<< m1 >>
rect 23 71 24 72 
<< m1 >>
rect 28 71 29 72 
<< pdiffusion >>
rect 30 71 31 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< m1 >>
rect 37 71 38 72 
<< m1 >>
rect 43 71 44 72 
<< m1 >>
rect 46 71 47 72 
<< pdiffusion >>
rect 48 71 49 72 
<< m1 >>
rect 49 71 50 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 63 71 64 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< m1 >>
rect 73 71 74 72 
<< m1 >>
rect 82 71 83 72 
<< m2 >>
rect 82 71 83 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< m1 >>
rect 98 71 99 72 
<< m1 >>
rect 100 71 101 72 
<< pdiffusion >>
rect 102 71 103 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< m1 >>
rect 106 71 107 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< m1 >>
rect 109 71 110 72 
<< m1 >>
rect 111 71 112 72 
<< m1 >>
rect 113 71 114 72 
<< m1 >>
rect 115 71 116 72 
<< m1 >>
rect 118 71 119 72 
<< m2 >>
rect 118 71 119 72 
<< pdiffusion >>
rect 120 71 121 72 
<< m1 >>
rect 121 71 122 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< m1 >>
rect 124 71 125 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< pdiffusion >>
rect 138 71 139 72 
<< m1 >>
rect 139 71 140 72 
<< pdiffusion >>
rect 139 71 140 72 
<< pdiffusion >>
rect 140 71 141 72 
<< pdiffusion >>
rect 141 71 142 72 
<< pdiffusion >>
rect 142 71 143 72 
<< pdiffusion >>
rect 143 71 144 72 
<< m1 >>
rect 146 71 147 72 
<< m1 >>
rect 154 71 155 72 
<< pdiffusion >>
rect 156 71 157 72 
<< pdiffusion >>
rect 157 71 158 72 
<< pdiffusion >>
rect 158 71 159 72 
<< pdiffusion >>
rect 159 71 160 72 
<< m1 >>
rect 160 71 161 72 
<< pdiffusion >>
rect 160 71 161 72 
<< pdiffusion >>
rect 161 71 162 72 
<< m1 >>
rect 163 71 164 72 
<< m2 >>
rect 163 71 164 72 
<< m2c >>
rect 163 71 164 72 
<< m1 >>
rect 163 71 164 72 
<< m2 >>
rect 163 71 164 72 
<< m1 >>
rect 164 71 165 72 
<< m1 >>
rect 169 71 170 72 
<< m2 >>
rect 169 71 170 72 
<< m1 >>
rect 171 71 172 72 
<< pdiffusion >>
rect 174 71 175 72 
<< pdiffusion >>
rect 175 71 176 72 
<< pdiffusion >>
rect 176 71 177 72 
<< pdiffusion >>
rect 177 71 178 72 
<< pdiffusion >>
rect 178 71 179 72 
<< pdiffusion >>
rect 179 71 180 72 
<< m1 >>
rect 10 72 11 73 
<< m1 >>
rect 19 72 20 73 
<< m2 >>
rect 20 72 21 73 
<< m2 >>
rect 22 72 23 73 
<< m1 >>
rect 23 72 24 73 
<< m1 >>
rect 28 72 29 73 
<< m1 >>
rect 37 72 38 73 
<< m1 >>
rect 43 72 44 73 
<< m1 >>
rect 46 72 47 73 
<< m1 >>
rect 49 72 50 73 
<< m1 >>
rect 63 72 64 73 
<< m1 >>
rect 73 72 74 73 
<< m1 >>
rect 82 72 83 73 
<< m2 >>
rect 82 72 83 73 
<< m1 >>
rect 98 72 99 73 
<< m1 >>
rect 100 72 101 73 
<< m1 >>
rect 106 72 107 73 
<< m2 >>
rect 106 72 107 73 
<< m2c >>
rect 106 72 107 73 
<< m1 >>
rect 106 72 107 73 
<< m2 >>
rect 106 72 107 73 
<< m1 >>
rect 109 72 110 73 
<< m1 >>
rect 111 72 112 73 
<< m1 >>
rect 113 72 114 73 
<< m1 >>
rect 115 72 116 73 
<< m1 >>
rect 118 72 119 73 
<< m2 >>
rect 118 72 119 73 
<< m1 >>
rect 121 72 122 73 
<< m1 >>
rect 124 72 125 73 
<< m1 >>
rect 139 72 140 73 
<< m1 >>
rect 146 72 147 73 
<< m1 >>
rect 154 72 155 73 
<< m1 >>
rect 160 72 161 73 
<< m2 >>
rect 163 72 164 73 
<< m1 >>
rect 169 72 170 73 
<< m2 >>
rect 169 72 170 73 
<< m1 >>
rect 171 72 172 73 
<< m1 >>
rect 10 73 11 74 
<< m1 >>
rect 17 73 18 74 
<< m2 >>
rect 17 73 18 74 
<< m2c >>
rect 17 73 18 74 
<< m1 >>
rect 17 73 18 74 
<< m2 >>
rect 17 73 18 74 
<< m2 >>
rect 18 73 19 74 
<< m1 >>
rect 19 73 20 74 
<< m2 >>
rect 19 73 20 74 
<< m2 >>
rect 20 73 21 74 
<< m2 >>
rect 22 73 23 74 
<< m1 >>
rect 23 73 24 74 
<< m1 >>
rect 28 73 29 74 
<< m1 >>
rect 37 73 38 74 
<< m1 >>
rect 43 73 44 74 
<< m1 >>
rect 46 73 47 74 
<< m1 >>
rect 49 73 50 74 
<< m1 >>
rect 63 73 64 74 
<< m1 >>
rect 73 73 74 74 
<< m1 >>
rect 82 73 83 74 
<< m2 >>
rect 82 73 83 74 
<< m1 >>
rect 98 73 99 74 
<< m2 >>
rect 98 73 99 74 
<< m2c >>
rect 98 73 99 74 
<< m1 >>
rect 98 73 99 74 
<< m2 >>
rect 98 73 99 74 
<< m2 >>
rect 99 73 100 74 
<< m1 >>
rect 100 73 101 74 
<< m2 >>
rect 100 73 101 74 
<< m2 >>
rect 101 73 102 74 
<< m1 >>
rect 102 73 103 74 
<< m2 >>
rect 102 73 103 74 
<< m2c >>
rect 102 73 103 74 
<< m1 >>
rect 102 73 103 74 
<< m2 >>
rect 102 73 103 74 
<< m2 >>
rect 106 73 107 74 
<< m1 >>
rect 109 73 110 74 
<< m1 >>
rect 111 73 112 74 
<< m1 >>
rect 113 73 114 74 
<< m1 >>
rect 115 73 116 74 
<< m1 >>
rect 118 73 119 74 
<< m2 >>
rect 118 73 119 74 
<< m1 >>
rect 119 73 120 74 
<< m2 >>
rect 119 73 120 74 
<< m1 >>
rect 120 73 121 74 
<< m1 >>
rect 121 73 122 74 
<< m1 >>
rect 124 73 125 74 
<< m1 >>
rect 139 73 140 74 
<< m1 >>
rect 146 73 147 74 
<< m1 >>
rect 154 73 155 74 
<< m1 >>
rect 160 73 161 74 
<< m1 >>
rect 161 73 162 74 
<< m1 >>
rect 162 73 163 74 
<< m1 >>
rect 163 73 164 74 
<< m2 >>
rect 163 73 164 74 
<< m1 >>
rect 164 73 165 74 
<< m1 >>
rect 165 73 166 74 
<< m1 >>
rect 166 73 167 74 
<< m1 >>
rect 167 73 168 74 
<< m1 >>
rect 169 73 170 74 
<< m2 >>
rect 169 73 170 74 
<< m1 >>
rect 171 73 172 74 
<< m1 >>
rect 10 74 11 75 
<< m1 >>
rect 16 74 17 75 
<< m1 >>
rect 17 74 18 75 
<< m1 >>
rect 19 74 20 75 
<< m2 >>
rect 22 74 23 75 
<< m1 >>
rect 23 74 24 75 
<< m1 >>
rect 28 74 29 75 
<< m1 >>
rect 37 74 38 75 
<< m2 >>
rect 37 74 38 75 
<< m2c >>
rect 37 74 38 75 
<< m1 >>
rect 37 74 38 75 
<< m2 >>
rect 37 74 38 75 
<< m1 >>
rect 43 74 44 75 
<< m2 >>
rect 43 74 44 75 
<< m2c >>
rect 43 74 44 75 
<< m1 >>
rect 43 74 44 75 
<< m2 >>
rect 43 74 44 75 
<< m1 >>
rect 46 74 47 75 
<< m2 >>
rect 46 74 47 75 
<< m2c >>
rect 46 74 47 75 
<< m1 >>
rect 46 74 47 75 
<< m2 >>
rect 46 74 47 75 
<< m1 >>
rect 49 74 50 75 
<< m1 >>
rect 58 74 59 75 
<< m1 >>
rect 59 74 60 75 
<< m1 >>
rect 60 74 61 75 
<< m1 >>
rect 61 74 62 75 
<< m1 >>
rect 62 74 63 75 
<< m1 >>
rect 63 74 64 75 
<< m1 >>
rect 73 74 74 75 
<< m2 >>
rect 73 74 74 75 
<< m2c >>
rect 73 74 74 75 
<< m1 >>
rect 73 74 74 75 
<< m2 >>
rect 73 74 74 75 
<< m1 >>
rect 82 74 83 75 
<< m2 >>
rect 82 74 83 75 
<< m1 >>
rect 100 74 101 75 
<< m1 >>
rect 102 74 103 75 
<< m1 >>
rect 106 74 107 75 
<< m2 >>
rect 106 74 107 75 
<< m1 >>
rect 107 74 108 75 
<< m1 >>
rect 108 74 109 75 
<< m1 >>
rect 109 74 110 75 
<< m1 >>
rect 111 74 112 75 
<< m1 >>
rect 113 74 114 75 
<< m1 >>
rect 115 74 116 75 
<< m2 >>
rect 119 74 120 75 
<< m1 >>
rect 124 74 125 75 
<< m1 >>
rect 139 74 140 75 
<< m1 >>
rect 146 74 147 75 
<< m1 >>
rect 154 74 155 75 
<< m2 >>
rect 163 74 164 75 
<< m1 >>
rect 167 74 168 75 
<< m1 >>
rect 169 74 170 75 
<< m2 >>
rect 169 74 170 75 
<< m1 >>
rect 171 74 172 75 
<< m1 >>
rect 10 75 11 76 
<< m1 >>
rect 16 75 17 76 
<< m1 >>
rect 19 75 20 76 
<< m2 >>
rect 22 75 23 76 
<< m1 >>
rect 23 75 24 76 
<< m1 >>
rect 28 75 29 76 
<< m2 >>
rect 37 75 38 76 
<< m2 >>
rect 43 75 44 76 
<< m2 >>
rect 45 75 46 76 
<< m2 >>
rect 46 75 47 76 
<< m1 >>
rect 49 75 50 76 
<< m1 >>
rect 58 75 59 76 
<< m2 >>
rect 73 75 74 76 
<< m1 >>
rect 82 75 83 76 
<< m2 >>
rect 82 75 83 76 
<< m1 >>
rect 100 75 101 76 
<< m2 >>
rect 100 75 101 76 
<< m2c >>
rect 100 75 101 76 
<< m1 >>
rect 100 75 101 76 
<< m2 >>
rect 100 75 101 76 
<< m1 >>
rect 102 75 103 76 
<< m2 >>
rect 102 75 103 76 
<< m2c >>
rect 102 75 103 76 
<< m1 >>
rect 102 75 103 76 
<< m2 >>
rect 102 75 103 76 
<< m1 >>
rect 106 75 107 76 
<< m2 >>
rect 106 75 107 76 
<< m2 >>
rect 107 75 108 76 
<< m2 >>
rect 108 75 109 76 
<< m2 >>
rect 109 75 110 76 
<< m2 >>
rect 110 75 111 76 
<< m1 >>
rect 111 75 112 76 
<< m2 >>
rect 111 75 112 76 
<< m2 >>
rect 112 75 113 76 
<< m1 >>
rect 113 75 114 76 
<< m2 >>
rect 113 75 114 76 
<< m2 >>
rect 114 75 115 76 
<< m1 >>
rect 115 75 116 76 
<< m2 >>
rect 115 75 116 76 
<< m2 >>
rect 116 75 117 76 
<< m1 >>
rect 117 75 118 76 
<< m2 >>
rect 117 75 118 76 
<< m2c >>
rect 117 75 118 76 
<< m1 >>
rect 117 75 118 76 
<< m2 >>
rect 117 75 118 76 
<< m1 >>
rect 118 75 119 76 
<< m1 >>
rect 119 75 120 76 
<< m2 >>
rect 119 75 120 76 
<< m1 >>
rect 120 75 121 76 
<< m1 >>
rect 124 75 125 76 
<< m1 >>
rect 139 75 140 76 
<< m1 >>
rect 146 75 147 76 
<< m1 >>
rect 154 75 155 76 
<< m1 >>
rect 163 75 164 76 
<< m2 >>
rect 163 75 164 76 
<< m2c >>
rect 163 75 164 76 
<< m1 >>
rect 163 75 164 76 
<< m2 >>
rect 163 75 164 76 
<< m1 >>
rect 167 75 168 76 
<< m1 >>
rect 169 75 170 76 
<< m2 >>
rect 169 75 170 76 
<< m1 >>
rect 171 75 172 76 
<< m1 >>
rect 10 76 11 77 
<< m1 >>
rect 16 76 17 77 
<< m1 >>
rect 19 76 20 77 
<< m2 >>
rect 22 76 23 77 
<< m1 >>
rect 23 76 24 77 
<< m1 >>
rect 26 76 27 77 
<< m2 >>
rect 26 76 27 77 
<< m2c >>
rect 26 76 27 77 
<< m1 >>
rect 26 76 27 77 
<< m2 >>
rect 26 76 27 77 
<< m2 >>
rect 27 76 28 77 
<< m1 >>
rect 28 76 29 77 
<< m2 >>
rect 28 76 29 77 
<< m2 >>
rect 29 76 30 77 
<< m1 >>
rect 30 76 31 77 
<< m2 >>
rect 30 76 31 77 
<< m2c >>
rect 30 76 31 77 
<< m1 >>
rect 30 76 31 77 
<< m2 >>
rect 30 76 31 77 
<< m1 >>
rect 31 76 32 77 
<< m1 >>
rect 32 76 33 77 
<< m1 >>
rect 33 76 34 77 
<< m1 >>
rect 34 76 35 77 
<< m1 >>
rect 35 76 36 77 
<< m1 >>
rect 36 76 37 77 
<< m1 >>
rect 37 76 38 77 
<< m2 >>
rect 37 76 38 77 
<< m1 >>
rect 38 76 39 77 
<< m1 >>
rect 39 76 40 77 
<< m1 >>
rect 40 76 41 77 
<< m1 >>
rect 41 76 42 77 
<< m1 >>
rect 42 76 43 77 
<< m1 >>
rect 43 76 44 77 
<< m2 >>
rect 43 76 44 77 
<< m1 >>
rect 44 76 45 77 
<< m1 >>
rect 45 76 46 77 
<< m2 >>
rect 45 76 46 77 
<< m1 >>
rect 46 76 47 77 
<< m1 >>
rect 47 76 48 77 
<< m1 >>
rect 48 76 49 77 
<< m1 >>
rect 49 76 50 77 
<< m1 >>
rect 58 76 59 77 
<< m1 >>
rect 62 76 63 77 
<< m1 >>
rect 63 76 64 77 
<< m1 >>
rect 64 76 65 77 
<< m1 >>
rect 65 76 66 77 
<< m1 >>
rect 66 76 67 77 
<< m1 >>
rect 67 76 68 77 
<< m1 >>
rect 68 76 69 77 
<< m1 >>
rect 69 76 70 77 
<< m1 >>
rect 70 76 71 77 
<< m1 >>
rect 71 76 72 77 
<< m1 >>
rect 72 76 73 77 
<< m1 >>
rect 73 76 74 77 
<< m2 >>
rect 73 76 74 77 
<< m1 >>
rect 74 76 75 77 
<< m1 >>
rect 75 76 76 77 
<< m1 >>
rect 76 76 77 77 
<< m1 >>
rect 77 76 78 77 
<< m1 >>
rect 78 76 79 77 
<< m1 >>
rect 79 76 80 77 
<< m1 >>
rect 80 76 81 77 
<< m1 >>
rect 81 76 82 77 
<< m1 >>
rect 82 76 83 77 
<< m2 >>
rect 82 76 83 77 
<< m2 >>
rect 84 76 85 77 
<< m2 >>
rect 85 76 86 77 
<< m2 >>
rect 86 76 87 77 
<< m2 >>
rect 87 76 88 77 
<< m2 >>
rect 88 76 89 77 
<< m2 >>
rect 89 76 90 77 
<< m2 >>
rect 90 76 91 77 
<< m2 >>
rect 91 76 92 77 
<< m2 >>
rect 92 76 93 77 
<< m2 >>
rect 93 76 94 77 
<< m2 >>
rect 94 76 95 77 
<< m2 >>
rect 95 76 96 77 
<< m2 >>
rect 96 76 97 77 
<< m2 >>
rect 97 76 98 77 
<< m2 >>
rect 98 76 99 77 
<< m2 >>
rect 99 76 100 77 
<< m2 >>
rect 100 76 101 77 
<< m2 >>
rect 102 76 103 77 
<< m1 >>
rect 106 76 107 77 
<< m1 >>
rect 111 76 112 77 
<< m1 >>
rect 113 76 114 77 
<< m1 >>
rect 115 76 116 77 
<< m2 >>
rect 119 76 120 77 
<< m1 >>
rect 120 76 121 77 
<< m1 >>
rect 124 76 125 77 
<< m1 >>
rect 139 76 140 77 
<< m1 >>
rect 146 76 147 77 
<< m1 >>
rect 154 76 155 77 
<< m1 >>
rect 163 76 164 77 
<< m1 >>
rect 167 76 168 77 
<< m1 >>
rect 169 76 170 77 
<< m2 >>
rect 169 76 170 77 
<< m1 >>
rect 171 76 172 77 
<< m1 >>
rect 10 77 11 78 
<< m1 >>
rect 16 77 17 78 
<< m1 >>
rect 19 77 20 78 
<< m2 >>
rect 22 77 23 78 
<< m1 >>
rect 23 77 24 78 
<< m1 >>
rect 26 77 27 78 
<< m1 >>
rect 28 77 29 78 
<< m2 >>
rect 37 77 38 78 
<< m2 >>
rect 43 77 44 78 
<< m2 >>
rect 45 77 46 78 
<< m1 >>
rect 58 77 59 78 
<< m1 >>
rect 62 77 63 78 
<< m2 >>
rect 73 77 74 78 
<< m2 >>
rect 82 77 83 78 
<< m1 >>
rect 84 77 85 78 
<< m2 >>
rect 84 77 85 78 
<< m1 >>
rect 85 77 86 78 
<< m1 >>
rect 86 77 87 78 
<< m1 >>
rect 87 77 88 78 
<< m1 >>
rect 88 77 89 78 
<< m1 >>
rect 89 77 90 78 
<< m1 >>
rect 90 77 91 78 
<< m1 >>
rect 91 77 92 78 
<< m1 >>
rect 92 77 93 78 
<< m1 >>
rect 93 77 94 78 
<< m1 >>
rect 94 77 95 78 
<< m1 >>
rect 95 77 96 78 
<< m1 >>
rect 96 77 97 78 
<< m1 >>
rect 97 77 98 78 
<< m1 >>
rect 98 77 99 78 
<< m1 >>
rect 99 77 100 78 
<< m1 >>
rect 100 77 101 78 
<< m1 >>
rect 101 77 102 78 
<< m1 >>
rect 102 77 103 78 
<< m2 >>
rect 102 77 103 78 
<< m1 >>
rect 103 77 104 78 
<< m1 >>
rect 104 77 105 78 
<< m2 >>
rect 104 77 105 78 
<< m2c >>
rect 104 77 105 78 
<< m1 >>
rect 104 77 105 78 
<< m2 >>
rect 104 77 105 78 
<< m2 >>
rect 105 77 106 78 
<< m1 >>
rect 106 77 107 78 
<< m2 >>
rect 106 77 107 78 
<< m2 >>
rect 107 77 108 78 
<< m1 >>
rect 108 77 109 78 
<< m2 >>
rect 108 77 109 78 
<< m2c >>
rect 108 77 109 78 
<< m1 >>
rect 108 77 109 78 
<< m2 >>
rect 108 77 109 78 
<< m1 >>
rect 109 77 110 78 
<< m2 >>
rect 109 77 110 78 
<< m2 >>
rect 110 77 111 78 
<< m1 >>
rect 111 77 112 78 
<< m2 >>
rect 111 77 112 78 
<< m2 >>
rect 112 77 113 78 
<< m1 >>
rect 113 77 114 78 
<< m2 >>
rect 113 77 114 78 
<< m2c >>
rect 113 77 114 78 
<< m1 >>
rect 113 77 114 78 
<< m2 >>
rect 113 77 114 78 
<< m1 >>
rect 115 77 116 78 
<< m2 >>
rect 115 77 116 78 
<< m2c >>
rect 115 77 116 78 
<< m1 >>
rect 115 77 116 78 
<< m2 >>
rect 115 77 116 78 
<< m2 >>
rect 119 77 120 78 
<< m1 >>
rect 120 77 121 78 
<< m1 >>
rect 121 77 122 78 
<< m1 >>
rect 122 77 123 78 
<< m2 >>
rect 122 77 123 78 
<< m2c >>
rect 122 77 123 78 
<< m1 >>
rect 122 77 123 78 
<< m2 >>
rect 122 77 123 78 
<< m2 >>
rect 123 77 124 78 
<< m1 >>
rect 124 77 125 78 
<< m2 >>
rect 124 77 125 78 
<< m2 >>
rect 125 77 126 78 
<< m1 >>
rect 126 77 127 78 
<< m2 >>
rect 126 77 127 78 
<< m2c >>
rect 126 77 127 78 
<< m1 >>
rect 126 77 127 78 
<< m2 >>
rect 126 77 127 78 
<< m1 >>
rect 127 77 128 78 
<< m1 >>
rect 128 77 129 78 
<< m1 >>
rect 129 77 130 78 
<< m1 >>
rect 130 77 131 78 
<< m1 >>
rect 131 77 132 78 
<< m1 >>
rect 132 77 133 78 
<< m1 >>
rect 133 77 134 78 
<< m1 >>
rect 134 77 135 78 
<< m1 >>
rect 135 77 136 78 
<< m1 >>
rect 136 77 137 78 
<< m1 >>
rect 137 77 138 78 
<< m2 >>
rect 137 77 138 78 
<< m2c >>
rect 137 77 138 78 
<< m1 >>
rect 137 77 138 78 
<< m2 >>
rect 137 77 138 78 
<< m2 >>
rect 138 77 139 78 
<< m1 >>
rect 139 77 140 78 
<< m2 >>
rect 139 77 140 78 
<< m2 >>
rect 140 77 141 78 
<< m1 >>
rect 146 77 147 78 
<< m1 >>
rect 154 77 155 78 
<< m1 >>
rect 163 77 164 78 
<< m1 >>
rect 167 77 168 78 
<< m1 >>
rect 169 77 170 78 
<< m2 >>
rect 169 77 170 78 
<< m1 >>
rect 171 77 172 78 
<< m1 >>
rect 10 78 11 79 
<< m1 >>
rect 16 78 17 79 
<< m1 >>
rect 19 78 20 79 
<< m2 >>
rect 22 78 23 79 
<< m1 >>
rect 23 78 24 79 
<< m1 >>
rect 24 78 25 79 
<< m2 >>
rect 24 78 25 79 
<< m2c >>
rect 24 78 25 79 
<< m1 >>
rect 24 78 25 79 
<< m2 >>
rect 24 78 25 79 
<< m2 >>
rect 25 78 26 79 
<< m1 >>
rect 26 78 27 79 
<< m2 >>
rect 26 78 27 79 
<< m2 >>
rect 27 78 28 79 
<< m1 >>
rect 28 78 29 79 
<< m2 >>
rect 28 78 29 79 
<< m2 >>
rect 29 78 30 79 
<< m1 >>
rect 30 78 31 79 
<< m2 >>
rect 30 78 31 79 
<< m2c >>
rect 30 78 31 79 
<< m1 >>
rect 30 78 31 79 
<< m2 >>
rect 30 78 31 79 
<< m1 >>
rect 31 78 32 79 
<< m1 >>
rect 32 78 33 79 
<< m1 >>
rect 33 78 34 79 
<< m1 >>
rect 34 78 35 79 
<< m1 >>
rect 35 78 36 79 
<< m1 >>
rect 36 78 37 79 
<< m1 >>
rect 37 78 38 79 
<< m2 >>
rect 37 78 38 79 
<< m1 >>
rect 38 78 39 79 
<< m1 >>
rect 39 78 40 79 
<< m1 >>
rect 40 78 41 79 
<< m1 >>
rect 41 78 42 79 
<< m1 >>
rect 42 78 43 79 
<< m1 >>
rect 43 78 44 79 
<< m2 >>
rect 43 78 44 79 
<< m1 >>
rect 44 78 45 79 
<< m1 >>
rect 45 78 46 79 
<< m2 >>
rect 45 78 46 79 
<< m1 >>
rect 46 78 47 79 
<< m1 >>
rect 47 78 48 79 
<< m1 >>
rect 48 78 49 79 
<< m1 >>
rect 49 78 50 79 
<< m1 >>
rect 58 78 59 79 
<< m1 >>
rect 62 78 63 79 
<< m1 >>
rect 73 78 74 79 
<< m2 >>
rect 73 78 74 79 
<< m2c >>
rect 73 78 74 79 
<< m1 >>
rect 73 78 74 79 
<< m2 >>
rect 73 78 74 79 
<< m1 >>
rect 82 78 83 79 
<< m2 >>
rect 82 78 83 79 
<< m2c >>
rect 82 78 83 79 
<< m1 >>
rect 82 78 83 79 
<< m2 >>
rect 82 78 83 79 
<< m1 >>
rect 84 78 85 79 
<< m2 >>
rect 84 78 85 79 
<< m2 >>
rect 102 78 103 79 
<< m1 >>
rect 106 78 107 79 
<< m1 >>
rect 111 78 112 79 
<< m2 >>
rect 115 78 116 79 
<< m2 >>
rect 119 78 120 79 
<< m1 >>
rect 124 78 125 79 
<< m1 >>
rect 139 78 140 79 
<< m2 >>
rect 140 78 141 79 
<< m1 >>
rect 146 78 147 79 
<< m1 >>
rect 154 78 155 79 
<< m1 >>
rect 163 78 164 79 
<< m1 >>
rect 167 78 168 79 
<< m1 >>
rect 169 78 170 79 
<< m2 >>
rect 169 78 170 79 
<< m1 >>
rect 171 78 172 79 
<< m1 >>
rect 10 79 11 80 
<< m1 >>
rect 16 79 17 80 
<< m1 >>
rect 19 79 20 80 
<< m2 >>
rect 22 79 23 80 
<< m1 >>
rect 26 79 27 80 
<< m1 >>
rect 28 79 29 80 
<< m2 >>
rect 37 79 38 80 
<< m2 >>
rect 43 79 44 80 
<< m2 >>
rect 45 79 46 80 
<< m2 >>
rect 48 79 49 80 
<< m1 >>
rect 49 79 50 80 
<< m2 >>
rect 49 79 50 80 
<< m2 >>
rect 50 79 51 80 
<< m1 >>
rect 51 79 52 80 
<< m2 >>
rect 51 79 52 80 
<< m2c >>
rect 51 79 52 80 
<< m1 >>
rect 51 79 52 80 
<< m2 >>
rect 51 79 52 80 
<< m1 >>
rect 52 79 53 80 
<< m1 >>
rect 53 79 54 80 
<< m1 >>
rect 54 79 55 80 
<< m1 >>
rect 55 79 56 80 
<< m1 >>
rect 56 79 57 80 
<< m2 >>
rect 56 79 57 80 
<< m2c >>
rect 56 79 57 80 
<< m1 >>
rect 56 79 57 80 
<< m2 >>
rect 56 79 57 80 
<< m2 >>
rect 57 79 58 80 
<< m1 >>
rect 58 79 59 80 
<< m2 >>
rect 58 79 59 80 
<< m2 >>
rect 59 79 60 80 
<< m1 >>
rect 60 79 61 80 
<< m2 >>
rect 60 79 61 80 
<< m2c >>
rect 60 79 61 80 
<< m1 >>
rect 60 79 61 80 
<< m2 >>
rect 60 79 61 80 
<< m2 >>
rect 61 79 62 80 
<< m1 >>
rect 62 79 63 80 
<< m2 >>
rect 62 79 63 80 
<< m2 >>
rect 63 79 64 80 
<< m1 >>
rect 64 79 65 80 
<< m2 >>
rect 64 79 65 80 
<< m1 >>
rect 65 79 66 80 
<< m2 >>
rect 65 79 66 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m1 >>
rect 67 79 68 80 
<< m2 >>
rect 67 79 68 80 
<< m1 >>
rect 68 79 69 80 
<< m2 >>
rect 68 79 69 80 
<< m2 >>
rect 69 79 70 80 
<< m1 >>
rect 73 79 74 80 
<< m2 >>
rect 82 79 83 80 
<< m1 >>
rect 84 79 85 80 
<< m2 >>
rect 84 79 85 80 
<< m1 >>
rect 88 79 89 80 
<< m1 >>
rect 89 79 90 80 
<< m1 >>
rect 90 79 91 80 
<< m1 >>
rect 91 79 92 80 
<< m1 >>
rect 92 79 93 80 
<< m1 >>
rect 93 79 94 80 
<< m1 >>
rect 94 79 95 80 
<< m1 >>
rect 95 79 96 80 
<< m1 >>
rect 96 79 97 80 
<< m1 >>
rect 97 79 98 80 
<< m1 >>
rect 98 79 99 80 
<< m1 >>
rect 99 79 100 80 
<< m1 >>
rect 100 79 101 80 
<< m1 >>
rect 101 79 102 80 
<< m1 >>
rect 102 79 103 80 
<< m2 >>
rect 102 79 103 80 
<< m1 >>
rect 103 79 104 80 
<< m1 >>
rect 104 79 105 80 
<< m2 >>
rect 104 79 105 80 
<< m2c >>
rect 104 79 105 80 
<< m1 >>
rect 104 79 105 80 
<< m2 >>
rect 104 79 105 80 
<< m2 >>
rect 105 79 106 80 
<< m1 >>
rect 106 79 107 80 
<< m2 >>
rect 106 79 107 80 
<< m2 >>
rect 107 79 108 80 
<< m1 >>
rect 108 79 109 80 
<< m2 >>
rect 108 79 109 80 
<< m2c >>
rect 108 79 109 80 
<< m1 >>
rect 108 79 109 80 
<< m2 >>
rect 108 79 109 80 
<< m1 >>
rect 109 79 110 80 
<< m1 >>
rect 110 79 111 80 
<< m1 >>
rect 111 79 112 80 
<< m1 >>
rect 113 79 114 80 
<< m1 >>
rect 114 79 115 80 
<< m1 >>
rect 115 79 116 80 
<< m2 >>
rect 115 79 116 80 
<< m1 >>
rect 116 79 117 80 
<< m1 >>
rect 117 79 118 80 
<< m1 >>
rect 118 79 119 80 
<< m1 >>
rect 119 79 120 80 
<< m2 >>
rect 119 79 120 80 
<< m1 >>
rect 120 79 121 80 
<< m1 >>
rect 121 79 122 80 
<< m1 >>
rect 122 79 123 80 
<< m2 >>
rect 122 79 123 80 
<< m2c >>
rect 122 79 123 80 
<< m1 >>
rect 122 79 123 80 
<< m2 >>
rect 122 79 123 80 
<< m2 >>
rect 123 79 124 80 
<< m1 >>
rect 124 79 125 80 
<< m2 >>
rect 124 79 125 80 
<< m2 >>
rect 125 79 126 80 
<< m1 >>
rect 126 79 127 80 
<< m2 >>
rect 126 79 127 80 
<< m2c >>
rect 126 79 127 80 
<< m1 >>
rect 126 79 127 80 
<< m2 >>
rect 126 79 127 80 
<< m1 >>
rect 127 79 128 80 
<< m1 >>
rect 128 79 129 80 
<< m1 >>
rect 129 79 130 80 
<< m1 >>
rect 130 79 131 80 
<< m1 >>
rect 131 79 132 80 
<< m1 >>
rect 132 79 133 80 
<< m1 >>
rect 133 79 134 80 
<< m1 >>
rect 134 79 135 80 
<< m1 >>
rect 135 79 136 80 
<< m1 >>
rect 136 79 137 80 
<< m1 >>
rect 137 79 138 80 
<< m1 >>
rect 138 79 139 80 
<< m1 >>
rect 139 79 140 80 
<< m2 >>
rect 140 79 141 80 
<< m1 >>
rect 146 79 147 80 
<< m1 >>
rect 154 79 155 80 
<< m1 >>
rect 163 79 164 80 
<< m1 >>
rect 167 79 168 80 
<< m1 >>
rect 169 79 170 80 
<< m2 >>
rect 169 79 170 80 
<< m1 >>
rect 171 79 172 80 
<< m1 >>
rect 10 80 11 81 
<< m2 >>
rect 10 80 11 81 
<< m2c >>
rect 10 80 11 81 
<< m1 >>
rect 10 80 11 81 
<< m2 >>
rect 10 80 11 81 
<< m1 >>
rect 16 80 17 81 
<< m1 >>
rect 19 80 20 81 
<< m1 >>
rect 22 80 23 81 
<< m2 >>
rect 22 80 23 81 
<< m2c >>
rect 22 80 23 81 
<< m1 >>
rect 22 80 23 81 
<< m2 >>
rect 22 80 23 81 
<< m1 >>
rect 26 80 27 81 
<< m1 >>
rect 28 80 29 81 
<< m1 >>
rect 37 80 38 81 
<< m2 >>
rect 37 80 38 81 
<< m2c >>
rect 37 80 38 81 
<< m1 >>
rect 37 80 38 81 
<< m2 >>
rect 37 80 38 81 
<< m1 >>
rect 43 80 44 81 
<< m2 >>
rect 43 80 44 81 
<< m2c >>
rect 43 80 44 81 
<< m1 >>
rect 43 80 44 81 
<< m2 >>
rect 43 80 44 81 
<< m1 >>
rect 45 80 46 81 
<< m2 >>
rect 45 80 46 81 
<< m2c >>
rect 45 80 46 81 
<< m1 >>
rect 45 80 46 81 
<< m2 >>
rect 45 80 46 81 
<< m1 >>
rect 47 80 48 81 
<< m2 >>
rect 47 80 48 81 
<< m2c >>
rect 47 80 48 81 
<< m1 >>
rect 47 80 48 81 
<< m2 >>
rect 47 80 48 81 
<< m2 >>
rect 48 80 49 81 
<< m1 >>
rect 49 80 50 81 
<< m1 >>
rect 58 80 59 81 
<< m1 >>
rect 62 80 63 81 
<< m1 >>
rect 64 80 65 81 
<< m1 >>
rect 68 80 69 81 
<< m1 >>
rect 69 80 70 81 
<< m2 >>
rect 69 80 70 81 
<< m1 >>
rect 70 80 71 81 
<< m1 >>
rect 71 80 72 81 
<< m2 >>
rect 71 80 72 81 
<< m2c >>
rect 71 80 72 81 
<< m1 >>
rect 71 80 72 81 
<< m2 >>
rect 71 80 72 81 
<< m2 >>
rect 72 80 73 81 
<< m1 >>
rect 73 80 74 81 
<< m2 >>
rect 73 80 74 81 
<< m2 >>
rect 74 80 75 81 
<< m1 >>
rect 75 80 76 81 
<< m2 >>
rect 75 80 76 81 
<< m2c >>
rect 75 80 76 81 
<< m1 >>
rect 75 80 76 81 
<< m2 >>
rect 75 80 76 81 
<< m1 >>
rect 76 80 77 81 
<< m1 >>
rect 77 80 78 81 
<< m1 >>
rect 78 80 79 81 
<< m1 >>
rect 79 80 80 81 
<< m1 >>
rect 80 80 81 81 
<< m1 >>
rect 81 80 82 81 
<< m1 >>
rect 82 80 83 81 
<< m2 >>
rect 82 80 83 81 
<< m1 >>
rect 83 80 84 81 
<< m1 >>
rect 84 80 85 81 
<< m2 >>
rect 84 80 85 81 
<< m1 >>
rect 88 80 89 81 
<< m2 >>
rect 100 80 101 81 
<< m2 >>
rect 101 80 102 81 
<< m2 >>
rect 102 80 103 81 
<< m1 >>
rect 106 80 107 81 
<< m1 >>
rect 113 80 114 81 
<< m2 >>
rect 115 80 116 81 
<< m2 >>
rect 119 80 120 81 
<< m1 >>
rect 124 80 125 81 
<< m2 >>
rect 140 80 141 81 
<< m1 >>
rect 146 80 147 81 
<< m1 >>
rect 154 80 155 81 
<< m2 >>
rect 154 80 155 81 
<< m2c >>
rect 154 80 155 81 
<< m1 >>
rect 154 80 155 81 
<< m2 >>
rect 154 80 155 81 
<< m1 >>
rect 163 80 164 81 
<< m2 >>
rect 163 80 164 81 
<< m2c >>
rect 163 80 164 81 
<< m1 >>
rect 163 80 164 81 
<< m2 >>
rect 163 80 164 81 
<< m1 >>
rect 167 80 168 81 
<< m1 >>
rect 169 80 170 81 
<< m2 >>
rect 169 80 170 81 
<< m1 >>
rect 171 80 172 81 
<< m2 >>
rect 10 81 11 82 
<< m1 >>
rect 16 81 17 82 
<< m1 >>
rect 19 81 20 82 
<< m1 >>
rect 22 81 23 82 
<< m1 >>
rect 26 81 27 82 
<< m1 >>
rect 28 81 29 82 
<< m1 >>
rect 37 81 38 82 
<< m2 >>
rect 43 81 44 82 
<< m2 >>
rect 45 81 46 82 
<< m1 >>
rect 47 81 48 82 
<< m1 >>
rect 49 81 50 82 
<< m1 >>
rect 58 81 59 82 
<< m1 >>
rect 62 81 63 82 
<< m1 >>
rect 64 81 65 82 
<< m2 >>
rect 69 81 70 82 
<< m1 >>
rect 73 81 74 82 
<< m2 >>
rect 82 81 83 82 
<< m2 >>
rect 84 81 85 82 
<< m1 >>
rect 88 81 89 82 
<< m1 >>
rect 100 81 101 82 
<< m2 >>
rect 100 81 101 82 
<< m2c >>
rect 100 81 101 82 
<< m1 >>
rect 100 81 101 82 
<< m2 >>
rect 100 81 101 82 
<< m1 >>
rect 106 81 107 82 
<< m1 >>
rect 113 81 114 82 
<< m1 >>
rect 115 81 116 82 
<< m2 >>
rect 115 81 116 82 
<< m2c >>
rect 115 81 116 82 
<< m1 >>
rect 115 81 116 82 
<< m2 >>
rect 115 81 116 82 
<< m1 >>
rect 116 81 117 82 
<< m1 >>
rect 117 81 118 82 
<< m1 >>
rect 118 81 119 82 
<< m1 >>
rect 119 81 120 82 
<< m2 >>
rect 119 81 120 82 
<< m1 >>
rect 120 81 121 82 
<< m1 >>
rect 121 81 122 82 
<< m1 >>
rect 124 81 125 82 
<< m1 >>
rect 125 81 126 82 
<< m1 >>
rect 126 81 127 82 
<< m1 >>
rect 127 81 128 82 
<< m1 >>
rect 128 81 129 82 
<< m1 >>
rect 129 81 130 82 
<< m1 >>
rect 130 81 131 82 
<< m1 >>
rect 131 81 132 82 
<< m1 >>
rect 132 81 133 82 
<< m1 >>
rect 133 81 134 82 
<< m1 >>
rect 134 81 135 82 
<< m1 >>
rect 135 81 136 82 
<< m1 >>
rect 136 81 137 82 
<< m1 >>
rect 139 81 140 82 
<< m1 >>
rect 140 81 141 82 
<< m2 >>
rect 140 81 141 82 
<< m1 >>
rect 141 81 142 82 
<< m2 >>
rect 141 81 142 82 
<< m1 >>
rect 142 81 143 82 
<< m2 >>
rect 142 81 143 82 
<< m1 >>
rect 143 81 144 82 
<< m2 >>
rect 143 81 144 82 
<< m1 >>
rect 144 81 145 82 
<< m2 >>
rect 144 81 145 82 
<< m1 >>
rect 145 81 146 82 
<< m2 >>
rect 145 81 146 82 
<< m1 >>
rect 146 81 147 82 
<< m2 >>
rect 146 81 147 82 
<< m2 >>
rect 147 81 148 82 
<< m2 >>
rect 154 81 155 82 
<< m2 >>
rect 163 81 164 82 
<< m1 >>
rect 167 81 168 82 
<< m1 >>
rect 169 81 170 82 
<< m2 >>
rect 169 81 170 82 
<< m1 >>
rect 171 81 172 82 
<< m1 >>
rect 10 82 11 83 
<< m2 >>
rect 10 82 11 83 
<< m1 >>
rect 11 82 12 83 
<< m1 >>
rect 12 82 13 83 
<< m1 >>
rect 13 82 14 83 
<< m1 >>
rect 16 82 17 83 
<< m1 >>
rect 19 82 20 83 
<< m1 >>
rect 22 82 23 83 
<< m1 >>
rect 26 82 27 83 
<< m1 >>
rect 28 82 29 83 
<< m1 >>
rect 37 82 38 83 
<< m2 >>
rect 38 82 39 83 
<< m1 >>
rect 39 82 40 83 
<< m2 >>
rect 39 82 40 83 
<< m2c >>
rect 39 82 40 83 
<< m1 >>
rect 39 82 40 83 
<< m2 >>
rect 39 82 40 83 
<< m1 >>
rect 40 82 41 83 
<< m1 >>
rect 41 82 42 83 
<< m1 >>
rect 42 82 43 83 
<< m1 >>
rect 43 82 44 83 
<< m2 >>
rect 43 82 44 83 
<< m1 >>
rect 44 82 45 83 
<< m1 >>
rect 45 82 46 83 
<< m2 >>
rect 45 82 46 83 
<< m1 >>
rect 46 82 47 83 
<< m1 >>
rect 47 82 48 83 
<< m1 >>
rect 49 82 50 83 
<< m1 >>
rect 58 82 59 83 
<< m1 >>
rect 62 82 63 83 
<< m1 >>
rect 64 82 65 83 
<< m1 >>
rect 69 82 70 83 
<< m2 >>
rect 69 82 70 83 
<< m2c >>
rect 69 82 70 83 
<< m1 >>
rect 69 82 70 83 
<< m2 >>
rect 69 82 70 83 
<< m1 >>
rect 70 82 71 83 
<< m1 >>
rect 73 82 74 83 
<< m2 >>
rect 74 82 75 83 
<< m1 >>
rect 75 82 76 83 
<< m2 >>
rect 75 82 76 83 
<< m2c >>
rect 75 82 76 83 
<< m1 >>
rect 75 82 76 83 
<< m2 >>
rect 75 82 76 83 
<< m1 >>
rect 76 82 77 83 
<< m1 >>
rect 77 82 78 83 
<< m1 >>
rect 78 82 79 83 
<< m1 >>
rect 79 82 80 83 
<< m1 >>
rect 80 82 81 83 
<< m1 >>
rect 81 82 82 83 
<< m1 >>
rect 82 82 83 83 
<< m2 >>
rect 82 82 83 83 
<< m1 >>
rect 83 82 84 83 
<< m1 >>
rect 84 82 85 83 
<< m2 >>
rect 84 82 85 83 
<< m2c >>
rect 84 82 85 83 
<< m1 >>
rect 84 82 85 83 
<< m2 >>
rect 84 82 85 83 
<< m1 >>
rect 88 82 89 83 
<< m1 >>
rect 100 82 101 83 
<< m1 >>
rect 106 82 107 83 
<< m1 >>
rect 113 82 114 83 
<< m2 >>
rect 117 82 118 83 
<< m2 >>
rect 118 82 119 83 
<< m2 >>
rect 119 82 120 83 
<< m1 >>
rect 121 82 122 83 
<< m1 >>
rect 136 82 137 83 
<< m1 >>
rect 139 82 140 83 
<< m2 >>
rect 147 82 148 83 
<< m1 >>
rect 148 82 149 83 
<< m2 >>
rect 148 82 149 83 
<< m2c >>
rect 148 82 149 83 
<< m1 >>
rect 148 82 149 83 
<< m2 >>
rect 148 82 149 83 
<< m1 >>
rect 149 82 150 83 
<< m1 >>
rect 150 82 151 83 
<< m1 >>
rect 151 82 152 83 
<< m1 >>
rect 152 82 153 83 
<< m1 >>
rect 153 82 154 83 
<< m2 >>
rect 154 82 155 83 
<< m1 >>
rect 160 82 161 83 
<< m1 >>
rect 161 82 162 83 
<< m1 >>
rect 162 82 163 83 
<< m1 >>
rect 163 82 164 83 
<< m2 >>
rect 163 82 164 83 
<< m1 >>
rect 167 82 168 83 
<< m1 >>
rect 169 82 170 83 
<< m2 >>
rect 169 82 170 83 
<< m1 >>
rect 171 82 172 83 
<< m1 >>
rect 10 83 11 84 
<< m2 >>
rect 10 83 11 84 
<< m1 >>
rect 13 83 14 84 
<< m1 >>
rect 16 83 17 84 
<< m1 >>
rect 19 83 20 84 
<< m1 >>
rect 22 83 23 84 
<< m1 >>
rect 26 83 27 84 
<< m1 >>
rect 28 83 29 84 
<< m1 >>
rect 37 83 38 84 
<< m2 >>
rect 38 83 39 84 
<< m2 >>
rect 43 83 44 84 
<< m2 >>
rect 45 83 46 84 
<< m1 >>
rect 49 83 50 84 
<< m1 >>
rect 58 83 59 84 
<< m1 >>
rect 62 83 63 84 
<< m1 >>
rect 64 83 65 84 
<< m1 >>
rect 70 83 71 84 
<< m1 >>
rect 73 83 74 84 
<< m2 >>
rect 74 83 75 84 
<< m2 >>
rect 82 83 83 84 
<< m1 >>
rect 88 83 89 84 
<< m1 >>
rect 100 83 101 84 
<< m1 >>
rect 106 83 107 84 
<< m1 >>
rect 113 83 114 84 
<< m1 >>
rect 117 83 118 84 
<< m2 >>
rect 117 83 118 84 
<< m2c >>
rect 117 83 118 84 
<< m1 >>
rect 117 83 118 84 
<< m2 >>
rect 117 83 118 84 
<< m1 >>
rect 121 83 122 84 
<< m1 >>
rect 136 83 137 84 
<< m1 >>
rect 139 83 140 84 
<< m1 >>
rect 153 83 154 84 
<< m2 >>
rect 154 83 155 84 
<< m1 >>
rect 160 83 161 84 
<< m1 >>
rect 163 83 164 84 
<< m2 >>
rect 163 83 164 84 
<< m1 >>
rect 167 83 168 84 
<< m1 >>
rect 169 83 170 84 
<< m2 >>
rect 169 83 170 84 
<< m1 >>
rect 171 83 172 84 
<< m1 >>
rect 10 84 11 85 
<< m2 >>
rect 10 84 11 85 
<< pdiffusion >>
rect 12 84 13 85 
<< m1 >>
rect 13 84 14 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< m1 >>
rect 16 84 17 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< m1 >>
rect 19 84 20 85 
<< m1 >>
rect 22 84 23 85 
<< m1 >>
rect 26 84 27 85 
<< m1 >>
rect 28 84 29 85 
<< pdiffusion >>
rect 30 84 31 85 
<< pdiffusion >>
rect 31 84 32 85 
<< pdiffusion >>
rect 32 84 33 85 
<< pdiffusion >>
rect 33 84 34 85 
<< pdiffusion >>
rect 34 84 35 85 
<< pdiffusion >>
rect 35 84 36 85 
<< m1 >>
rect 37 84 38 85 
<< m2 >>
rect 38 84 39 85 
<< m1 >>
rect 43 84 44 85 
<< m2 >>
rect 43 84 44 85 
<< m2c >>
rect 43 84 44 85 
<< m1 >>
rect 43 84 44 85 
<< m2 >>
rect 43 84 44 85 
<< m1 >>
rect 45 84 46 85 
<< m2 >>
rect 45 84 46 85 
<< m2c >>
rect 45 84 46 85 
<< m1 >>
rect 45 84 46 85 
<< m2 >>
rect 45 84 46 85 
<< pdiffusion >>
rect 48 84 49 85 
<< m1 >>
rect 49 84 50 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< m1 >>
rect 58 84 59 85 
<< m1 >>
rect 62 84 63 85 
<< m1 >>
rect 64 84 65 85 
<< pdiffusion >>
rect 66 84 67 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< m1 >>
rect 70 84 71 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< m1 >>
rect 73 84 74 85 
<< m2 >>
rect 74 84 75 85 
<< m1 >>
rect 82 84 83 85 
<< m2 >>
rect 82 84 83 85 
<< m2c >>
rect 82 84 83 85 
<< m1 >>
rect 82 84 83 85 
<< m2 >>
rect 82 84 83 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< m1 >>
rect 88 84 89 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 100 84 101 85 
<< pdiffusion >>
rect 102 84 103 85 
<< pdiffusion >>
rect 103 84 104 85 
<< pdiffusion >>
rect 104 84 105 85 
<< pdiffusion >>
rect 105 84 106 85 
<< m1 >>
rect 106 84 107 85 
<< pdiffusion >>
rect 106 84 107 85 
<< pdiffusion >>
rect 107 84 108 85 
<< m1 >>
rect 113 84 114 85 
<< m1 >>
rect 117 84 118 85 
<< pdiffusion >>
rect 120 84 121 85 
<< m1 >>
rect 121 84 122 85 
<< pdiffusion >>
rect 121 84 122 85 
<< pdiffusion >>
rect 122 84 123 85 
<< pdiffusion >>
rect 123 84 124 85 
<< pdiffusion >>
rect 124 84 125 85 
<< pdiffusion >>
rect 125 84 126 85 
<< m1 >>
rect 136 84 137 85 
<< pdiffusion >>
rect 138 84 139 85 
<< m1 >>
rect 139 84 140 85 
<< pdiffusion >>
rect 139 84 140 85 
<< pdiffusion >>
rect 140 84 141 85 
<< pdiffusion >>
rect 141 84 142 85 
<< pdiffusion >>
rect 142 84 143 85 
<< pdiffusion >>
rect 143 84 144 85 
<< m1 >>
rect 151 84 152 85 
<< m2 >>
rect 151 84 152 85 
<< m2c >>
rect 151 84 152 85 
<< m1 >>
rect 151 84 152 85 
<< m2 >>
rect 151 84 152 85 
<< m2 >>
rect 152 84 153 85 
<< m1 >>
rect 153 84 154 85 
<< m2 >>
rect 153 84 154 85 
<< m2 >>
rect 154 84 155 85 
<< pdiffusion >>
rect 156 84 157 85 
<< pdiffusion >>
rect 157 84 158 85 
<< pdiffusion >>
rect 158 84 159 85 
<< pdiffusion >>
rect 159 84 160 85 
<< m1 >>
rect 160 84 161 85 
<< pdiffusion >>
rect 160 84 161 85 
<< pdiffusion >>
rect 161 84 162 85 
<< m1 >>
rect 163 84 164 85 
<< m2 >>
rect 163 84 164 85 
<< m1 >>
rect 167 84 168 85 
<< m1 >>
rect 169 84 170 85 
<< m2 >>
rect 169 84 170 85 
<< m1 >>
rect 171 84 172 85 
<< pdiffusion >>
rect 174 84 175 85 
<< pdiffusion >>
rect 175 84 176 85 
<< pdiffusion >>
rect 176 84 177 85 
<< pdiffusion >>
rect 177 84 178 85 
<< pdiffusion >>
rect 178 84 179 85 
<< pdiffusion >>
rect 179 84 180 85 
<< m1 >>
rect 10 85 11 86 
<< m2 >>
rect 10 85 11 86 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< m1 >>
rect 19 85 20 86 
<< m1 >>
rect 22 85 23 86 
<< m1 >>
rect 26 85 27 86 
<< m1 >>
rect 28 85 29 86 
<< pdiffusion >>
rect 30 85 31 86 
<< pdiffusion >>
rect 31 85 32 86 
<< pdiffusion >>
rect 32 85 33 86 
<< pdiffusion >>
rect 33 85 34 86 
<< pdiffusion >>
rect 34 85 35 86 
<< pdiffusion >>
rect 35 85 36 86 
<< m1 >>
rect 37 85 38 86 
<< m2 >>
rect 38 85 39 86 
<< m1 >>
rect 43 85 44 86 
<< m1 >>
rect 45 85 46 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< m1 >>
rect 58 85 59 86 
<< m1 >>
rect 62 85 63 86 
<< m1 >>
rect 64 85 65 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< m1 >>
rect 73 85 74 86 
<< m2 >>
rect 74 85 75 86 
<< m1 >>
rect 82 85 83 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 100 85 101 86 
<< pdiffusion >>
rect 102 85 103 86 
<< pdiffusion >>
rect 103 85 104 86 
<< pdiffusion >>
rect 104 85 105 86 
<< pdiffusion >>
rect 105 85 106 86 
<< pdiffusion >>
rect 106 85 107 86 
<< pdiffusion >>
rect 107 85 108 86 
<< m1 >>
rect 113 85 114 86 
<< m1 >>
rect 117 85 118 86 
<< pdiffusion >>
rect 120 85 121 86 
<< pdiffusion >>
rect 121 85 122 86 
<< pdiffusion >>
rect 122 85 123 86 
<< pdiffusion >>
rect 123 85 124 86 
<< pdiffusion >>
rect 124 85 125 86 
<< pdiffusion >>
rect 125 85 126 86 
<< m1 >>
rect 136 85 137 86 
<< pdiffusion >>
rect 138 85 139 86 
<< pdiffusion >>
rect 139 85 140 86 
<< pdiffusion >>
rect 140 85 141 86 
<< pdiffusion >>
rect 141 85 142 86 
<< pdiffusion >>
rect 142 85 143 86 
<< pdiffusion >>
rect 143 85 144 86 
<< m1 >>
rect 151 85 152 86 
<< m1 >>
rect 153 85 154 86 
<< pdiffusion >>
rect 156 85 157 86 
<< pdiffusion >>
rect 157 85 158 86 
<< pdiffusion >>
rect 158 85 159 86 
<< pdiffusion >>
rect 159 85 160 86 
<< pdiffusion >>
rect 160 85 161 86 
<< pdiffusion >>
rect 161 85 162 86 
<< m1 >>
rect 163 85 164 86 
<< m2 >>
rect 163 85 164 86 
<< m1 >>
rect 167 85 168 86 
<< m1 >>
rect 169 85 170 86 
<< m2 >>
rect 169 85 170 86 
<< m1 >>
rect 171 85 172 86 
<< pdiffusion >>
rect 174 85 175 86 
<< pdiffusion >>
rect 175 85 176 86 
<< pdiffusion >>
rect 176 85 177 86 
<< pdiffusion >>
rect 177 85 178 86 
<< pdiffusion >>
rect 178 85 179 86 
<< pdiffusion >>
rect 179 85 180 86 
<< m1 >>
rect 10 86 11 87 
<< m2 >>
rect 10 86 11 87 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< m1 >>
rect 19 86 20 87 
<< m1 >>
rect 22 86 23 87 
<< m1 >>
rect 26 86 27 87 
<< m1 >>
rect 28 86 29 87 
<< pdiffusion >>
rect 30 86 31 87 
<< pdiffusion >>
rect 31 86 32 87 
<< pdiffusion >>
rect 32 86 33 87 
<< pdiffusion >>
rect 33 86 34 87 
<< pdiffusion >>
rect 34 86 35 87 
<< pdiffusion >>
rect 35 86 36 87 
<< m1 >>
rect 37 86 38 87 
<< m2 >>
rect 38 86 39 87 
<< m1 >>
rect 43 86 44 87 
<< m1 >>
rect 45 86 46 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< m1 >>
rect 58 86 59 87 
<< m1 >>
rect 62 86 63 87 
<< m1 >>
rect 64 86 65 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< m1 >>
rect 73 86 74 87 
<< m2 >>
rect 74 86 75 87 
<< m1 >>
rect 82 86 83 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 100 86 101 87 
<< pdiffusion >>
rect 102 86 103 87 
<< pdiffusion >>
rect 103 86 104 87 
<< pdiffusion >>
rect 104 86 105 87 
<< pdiffusion >>
rect 105 86 106 87 
<< pdiffusion >>
rect 106 86 107 87 
<< pdiffusion >>
rect 107 86 108 87 
<< m1 >>
rect 113 86 114 87 
<< m1 >>
rect 117 86 118 87 
<< pdiffusion >>
rect 120 86 121 87 
<< pdiffusion >>
rect 121 86 122 87 
<< pdiffusion >>
rect 122 86 123 87 
<< pdiffusion >>
rect 123 86 124 87 
<< pdiffusion >>
rect 124 86 125 87 
<< pdiffusion >>
rect 125 86 126 87 
<< m1 >>
rect 136 86 137 87 
<< pdiffusion >>
rect 138 86 139 87 
<< pdiffusion >>
rect 139 86 140 87 
<< pdiffusion >>
rect 140 86 141 87 
<< pdiffusion >>
rect 141 86 142 87 
<< pdiffusion >>
rect 142 86 143 87 
<< pdiffusion >>
rect 143 86 144 87 
<< m1 >>
rect 151 86 152 87 
<< m1 >>
rect 153 86 154 87 
<< pdiffusion >>
rect 156 86 157 87 
<< pdiffusion >>
rect 157 86 158 87 
<< pdiffusion >>
rect 158 86 159 87 
<< pdiffusion >>
rect 159 86 160 87 
<< pdiffusion >>
rect 160 86 161 87 
<< pdiffusion >>
rect 161 86 162 87 
<< m1 >>
rect 163 86 164 87 
<< m2 >>
rect 163 86 164 87 
<< m1 >>
rect 167 86 168 87 
<< m1 >>
rect 169 86 170 87 
<< m2 >>
rect 169 86 170 87 
<< m1 >>
rect 171 86 172 87 
<< pdiffusion >>
rect 174 86 175 87 
<< pdiffusion >>
rect 175 86 176 87 
<< pdiffusion >>
rect 176 86 177 87 
<< pdiffusion >>
rect 177 86 178 87 
<< pdiffusion >>
rect 178 86 179 87 
<< pdiffusion >>
rect 179 86 180 87 
<< m1 >>
rect 10 87 11 88 
<< m2 >>
rect 10 87 11 88 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< m1 >>
rect 19 87 20 88 
<< m1 >>
rect 22 87 23 88 
<< m1 >>
rect 26 87 27 88 
<< m1 >>
rect 28 87 29 88 
<< pdiffusion >>
rect 30 87 31 88 
<< pdiffusion >>
rect 31 87 32 88 
<< pdiffusion >>
rect 32 87 33 88 
<< pdiffusion >>
rect 33 87 34 88 
<< pdiffusion >>
rect 34 87 35 88 
<< pdiffusion >>
rect 35 87 36 88 
<< m1 >>
rect 37 87 38 88 
<< m2 >>
rect 38 87 39 88 
<< m1 >>
rect 43 87 44 88 
<< m1 >>
rect 45 87 46 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< m1 >>
rect 58 87 59 88 
<< m1 >>
rect 62 87 63 88 
<< m1 >>
rect 64 87 65 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< m1 >>
rect 73 87 74 88 
<< m2 >>
rect 74 87 75 88 
<< m1 >>
rect 82 87 83 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 100 87 101 88 
<< pdiffusion >>
rect 102 87 103 88 
<< pdiffusion >>
rect 103 87 104 88 
<< pdiffusion >>
rect 104 87 105 88 
<< pdiffusion >>
rect 105 87 106 88 
<< pdiffusion >>
rect 106 87 107 88 
<< pdiffusion >>
rect 107 87 108 88 
<< m1 >>
rect 113 87 114 88 
<< m1 >>
rect 117 87 118 88 
<< pdiffusion >>
rect 120 87 121 88 
<< pdiffusion >>
rect 121 87 122 88 
<< pdiffusion >>
rect 122 87 123 88 
<< pdiffusion >>
rect 123 87 124 88 
<< pdiffusion >>
rect 124 87 125 88 
<< pdiffusion >>
rect 125 87 126 88 
<< m1 >>
rect 136 87 137 88 
<< pdiffusion >>
rect 138 87 139 88 
<< pdiffusion >>
rect 139 87 140 88 
<< pdiffusion >>
rect 140 87 141 88 
<< pdiffusion >>
rect 141 87 142 88 
<< pdiffusion >>
rect 142 87 143 88 
<< pdiffusion >>
rect 143 87 144 88 
<< m1 >>
rect 151 87 152 88 
<< m1 >>
rect 153 87 154 88 
<< pdiffusion >>
rect 156 87 157 88 
<< pdiffusion >>
rect 157 87 158 88 
<< pdiffusion >>
rect 158 87 159 88 
<< pdiffusion >>
rect 159 87 160 88 
<< pdiffusion >>
rect 160 87 161 88 
<< pdiffusion >>
rect 161 87 162 88 
<< m1 >>
rect 163 87 164 88 
<< m2 >>
rect 163 87 164 88 
<< m1 >>
rect 167 87 168 88 
<< m1 >>
rect 169 87 170 88 
<< m2 >>
rect 169 87 170 88 
<< m1 >>
rect 171 87 172 88 
<< pdiffusion >>
rect 174 87 175 88 
<< pdiffusion >>
rect 175 87 176 88 
<< pdiffusion >>
rect 176 87 177 88 
<< pdiffusion >>
rect 177 87 178 88 
<< pdiffusion >>
rect 178 87 179 88 
<< pdiffusion >>
rect 179 87 180 88 
<< m1 >>
rect 10 88 11 89 
<< m2 >>
rect 10 88 11 89 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< m1 >>
rect 19 88 20 89 
<< m1 >>
rect 22 88 23 89 
<< m1 >>
rect 26 88 27 89 
<< m1 >>
rect 28 88 29 89 
<< pdiffusion >>
rect 30 88 31 89 
<< pdiffusion >>
rect 31 88 32 89 
<< pdiffusion >>
rect 32 88 33 89 
<< pdiffusion >>
rect 33 88 34 89 
<< pdiffusion >>
rect 34 88 35 89 
<< pdiffusion >>
rect 35 88 36 89 
<< m1 >>
rect 37 88 38 89 
<< m2 >>
rect 38 88 39 89 
<< m1 >>
rect 43 88 44 89 
<< m1 >>
rect 45 88 46 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< m1 >>
rect 58 88 59 89 
<< m1 >>
rect 62 88 63 89 
<< m1 >>
rect 64 88 65 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< m1 >>
rect 73 88 74 89 
<< m2 >>
rect 74 88 75 89 
<< m1 >>
rect 82 88 83 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 100 88 101 89 
<< pdiffusion >>
rect 102 88 103 89 
<< pdiffusion >>
rect 103 88 104 89 
<< pdiffusion >>
rect 104 88 105 89 
<< pdiffusion >>
rect 105 88 106 89 
<< pdiffusion >>
rect 106 88 107 89 
<< pdiffusion >>
rect 107 88 108 89 
<< m1 >>
rect 113 88 114 89 
<< m1 >>
rect 117 88 118 89 
<< pdiffusion >>
rect 120 88 121 89 
<< pdiffusion >>
rect 121 88 122 89 
<< pdiffusion >>
rect 122 88 123 89 
<< pdiffusion >>
rect 123 88 124 89 
<< pdiffusion >>
rect 124 88 125 89 
<< pdiffusion >>
rect 125 88 126 89 
<< m1 >>
rect 136 88 137 89 
<< pdiffusion >>
rect 138 88 139 89 
<< pdiffusion >>
rect 139 88 140 89 
<< pdiffusion >>
rect 140 88 141 89 
<< pdiffusion >>
rect 141 88 142 89 
<< pdiffusion >>
rect 142 88 143 89 
<< pdiffusion >>
rect 143 88 144 89 
<< m1 >>
rect 151 88 152 89 
<< m1 >>
rect 153 88 154 89 
<< pdiffusion >>
rect 156 88 157 89 
<< pdiffusion >>
rect 157 88 158 89 
<< pdiffusion >>
rect 158 88 159 89 
<< pdiffusion >>
rect 159 88 160 89 
<< pdiffusion >>
rect 160 88 161 89 
<< pdiffusion >>
rect 161 88 162 89 
<< m1 >>
rect 163 88 164 89 
<< m2 >>
rect 163 88 164 89 
<< m1 >>
rect 167 88 168 89 
<< m1 >>
rect 169 88 170 89 
<< m2 >>
rect 169 88 170 89 
<< m1 >>
rect 171 88 172 89 
<< pdiffusion >>
rect 174 88 175 89 
<< pdiffusion >>
rect 175 88 176 89 
<< pdiffusion >>
rect 176 88 177 89 
<< pdiffusion >>
rect 177 88 178 89 
<< pdiffusion >>
rect 178 88 179 89 
<< pdiffusion >>
rect 179 88 180 89 
<< m1 >>
rect 10 89 11 90 
<< m2 >>
rect 10 89 11 90 
<< pdiffusion >>
rect 12 89 13 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< m1 >>
rect 19 89 20 90 
<< m1 >>
rect 22 89 23 90 
<< m1 >>
rect 26 89 27 90 
<< m1 >>
rect 28 89 29 90 
<< pdiffusion >>
rect 30 89 31 90 
<< m1 >>
rect 31 89 32 90 
<< pdiffusion >>
rect 31 89 32 90 
<< pdiffusion >>
rect 32 89 33 90 
<< pdiffusion >>
rect 33 89 34 90 
<< pdiffusion >>
rect 34 89 35 90 
<< pdiffusion >>
rect 35 89 36 90 
<< m1 >>
rect 37 89 38 90 
<< m2 >>
rect 38 89 39 90 
<< m1 >>
rect 43 89 44 90 
<< m1 >>
rect 45 89 46 90 
<< pdiffusion >>
rect 48 89 49 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< m1 >>
rect 52 89 53 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< m1 >>
rect 58 89 59 90 
<< m1 >>
rect 62 89 63 90 
<< m1 >>
rect 64 89 65 90 
<< pdiffusion >>
rect 66 89 67 90 
<< m1 >>
rect 67 89 68 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< m1 >>
rect 70 89 71 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< m1 >>
rect 73 89 74 90 
<< m2 >>
rect 74 89 75 90 
<< m1 >>
rect 82 89 83 90 
<< pdiffusion >>
rect 84 89 85 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 100 89 101 90 
<< pdiffusion >>
rect 102 89 103 90 
<< m1 >>
rect 103 89 104 90 
<< pdiffusion >>
rect 103 89 104 90 
<< pdiffusion >>
rect 104 89 105 90 
<< pdiffusion >>
rect 105 89 106 90 
<< m1 >>
rect 106 89 107 90 
<< pdiffusion >>
rect 106 89 107 90 
<< pdiffusion >>
rect 107 89 108 90 
<< m1 >>
rect 113 89 114 90 
<< m1 >>
rect 117 89 118 90 
<< pdiffusion >>
rect 120 89 121 90 
<< pdiffusion >>
rect 121 89 122 90 
<< pdiffusion >>
rect 122 89 123 90 
<< pdiffusion >>
rect 123 89 124 90 
<< pdiffusion >>
rect 124 89 125 90 
<< pdiffusion >>
rect 125 89 126 90 
<< m1 >>
rect 136 89 137 90 
<< pdiffusion >>
rect 138 89 139 90 
<< pdiffusion >>
rect 139 89 140 90 
<< pdiffusion >>
rect 140 89 141 90 
<< pdiffusion >>
rect 141 89 142 90 
<< pdiffusion >>
rect 142 89 143 90 
<< pdiffusion >>
rect 143 89 144 90 
<< m1 >>
rect 151 89 152 90 
<< m1 >>
rect 153 89 154 90 
<< pdiffusion >>
rect 156 89 157 90 
<< pdiffusion >>
rect 157 89 158 90 
<< pdiffusion >>
rect 158 89 159 90 
<< pdiffusion >>
rect 159 89 160 90 
<< pdiffusion >>
rect 160 89 161 90 
<< pdiffusion >>
rect 161 89 162 90 
<< m1 >>
rect 163 89 164 90 
<< m2 >>
rect 163 89 164 90 
<< m1 >>
rect 167 89 168 90 
<< m1 >>
rect 169 89 170 90 
<< m2 >>
rect 169 89 170 90 
<< m1 >>
rect 171 89 172 90 
<< m2 >>
rect 171 89 172 90 
<< m2c >>
rect 171 89 172 90 
<< m1 >>
rect 171 89 172 90 
<< m2 >>
rect 171 89 172 90 
<< pdiffusion >>
rect 174 89 175 90 
<< m1 >>
rect 175 89 176 90 
<< pdiffusion >>
rect 175 89 176 90 
<< pdiffusion >>
rect 176 89 177 90 
<< pdiffusion >>
rect 177 89 178 90 
<< m1 >>
rect 178 89 179 90 
<< pdiffusion >>
rect 178 89 179 90 
<< pdiffusion >>
rect 179 89 180 90 
<< m1 >>
rect 10 90 11 91 
<< m2 >>
rect 10 90 11 91 
<< m1 >>
rect 19 90 20 91 
<< m1 >>
rect 22 90 23 91 
<< m1 >>
rect 26 90 27 91 
<< m1 >>
rect 28 90 29 91 
<< m1 >>
rect 31 90 32 91 
<< m1 >>
rect 37 90 38 91 
<< m2 >>
rect 38 90 39 91 
<< m1 >>
rect 43 90 44 91 
<< m1 >>
rect 45 90 46 91 
<< m1 >>
rect 52 90 53 91 
<< m1 >>
rect 58 90 59 91 
<< m1 >>
rect 62 90 63 91 
<< m1 >>
rect 64 90 65 91 
<< m1 >>
rect 67 90 68 91 
<< m1 >>
rect 70 90 71 91 
<< m1 >>
rect 73 90 74 91 
<< m2 >>
rect 74 90 75 91 
<< m1 >>
rect 82 90 83 91 
<< m1 >>
rect 100 90 101 91 
<< m1 >>
rect 103 90 104 91 
<< m1 >>
rect 106 90 107 91 
<< m1 >>
rect 113 90 114 91 
<< m1 >>
rect 117 90 118 91 
<< m1 >>
rect 136 90 137 91 
<< m1 >>
rect 151 90 152 91 
<< m1 >>
rect 153 90 154 91 
<< m1 >>
rect 163 90 164 91 
<< m2 >>
rect 163 90 164 91 
<< m1 >>
rect 167 90 168 91 
<< m1 >>
rect 169 90 170 91 
<< m2 >>
rect 169 90 170 91 
<< m2 >>
rect 171 90 172 91 
<< m1 >>
rect 175 90 176 91 
<< m1 >>
rect 178 90 179 91 
<< m1 >>
rect 10 91 11 92 
<< m2 >>
rect 10 91 11 92 
<< m1 >>
rect 19 91 20 92 
<< m1 >>
rect 22 91 23 92 
<< m1 >>
rect 26 91 27 92 
<< m1 >>
rect 28 91 29 92 
<< m1 >>
rect 31 91 32 92 
<< m1 >>
rect 35 91 36 92 
<< m2 >>
rect 35 91 36 92 
<< m2c >>
rect 35 91 36 92 
<< m1 >>
rect 35 91 36 92 
<< m2 >>
rect 35 91 36 92 
<< m2 >>
rect 36 91 37 92 
<< m1 >>
rect 37 91 38 92 
<< m2 >>
rect 37 91 38 92 
<< m2 >>
rect 38 91 39 92 
<< m1 >>
rect 43 91 44 92 
<< m1 >>
rect 45 91 46 92 
<< m1 >>
rect 52 91 53 92 
<< m1 >>
rect 58 91 59 92 
<< m1 >>
rect 62 91 63 92 
<< m1 >>
rect 64 91 65 92 
<< m1 >>
rect 67 91 68 92 
<< m1 >>
rect 70 91 71 92 
<< m1 >>
rect 71 91 72 92 
<< m2 >>
rect 71 91 72 92 
<< m2c >>
rect 71 91 72 92 
<< m1 >>
rect 71 91 72 92 
<< m2 >>
rect 71 91 72 92 
<< m2 >>
rect 72 91 73 92 
<< m1 >>
rect 73 91 74 92 
<< m2 >>
rect 73 91 74 92 
<< m2 >>
rect 74 91 75 92 
<< m1 >>
rect 82 91 83 92 
<< m2 >>
rect 82 91 83 92 
<< m2c >>
rect 82 91 83 92 
<< m1 >>
rect 82 91 83 92 
<< m2 >>
rect 82 91 83 92 
<< m1 >>
rect 100 91 101 92 
<< m1 >>
rect 101 91 102 92 
<< m1 >>
rect 102 91 103 92 
<< m1 >>
rect 103 91 104 92 
<< m1 >>
rect 106 91 107 92 
<< m1 >>
rect 113 91 114 92 
<< m1 >>
rect 117 91 118 92 
<< m1 >>
rect 136 91 137 92 
<< m1 >>
rect 151 91 152 92 
<< m1 >>
rect 153 91 154 92 
<< m1 >>
rect 163 91 164 92 
<< m2 >>
rect 163 91 164 92 
<< m1 >>
rect 167 91 168 92 
<< m1 >>
rect 169 91 170 92 
<< m2 >>
rect 169 91 170 92 
<< m1 >>
rect 170 91 171 92 
<< m1 >>
rect 171 91 172 92 
<< m2 >>
rect 171 91 172 92 
<< m1 >>
rect 172 91 173 92 
<< m1 >>
rect 173 91 174 92 
<< m1 >>
rect 174 91 175 92 
<< m1 >>
rect 175 91 176 92 
<< m1 >>
rect 178 91 179 92 
<< m1 >>
rect 10 92 11 93 
<< m2 >>
rect 10 92 11 93 
<< m1 >>
rect 19 92 20 93 
<< m1 >>
rect 22 92 23 93 
<< m1 >>
rect 26 92 27 93 
<< m1 >>
rect 28 92 29 93 
<< m1 >>
rect 31 92 32 93 
<< m1 >>
rect 32 92 33 93 
<< m1 >>
rect 33 92 34 93 
<< m1 >>
rect 34 92 35 93 
<< m1 >>
rect 35 92 36 93 
<< m1 >>
rect 37 92 38 93 
<< m1 >>
rect 43 92 44 93 
<< m1 >>
rect 45 92 46 93 
<< m1 >>
rect 52 92 53 93 
<< m1 >>
rect 54 92 55 93 
<< m1 >>
rect 55 92 56 93 
<< m1 >>
rect 56 92 57 93 
<< m2 >>
rect 56 92 57 93 
<< m2c >>
rect 56 92 57 93 
<< m1 >>
rect 56 92 57 93 
<< m2 >>
rect 56 92 57 93 
<< m2 >>
rect 57 92 58 93 
<< m1 >>
rect 58 92 59 93 
<< m2 >>
rect 58 92 59 93 
<< m2 >>
rect 59 92 60 93 
<< m1 >>
rect 60 92 61 93 
<< m2 >>
rect 60 92 61 93 
<< m2c >>
rect 60 92 61 93 
<< m1 >>
rect 60 92 61 93 
<< m2 >>
rect 60 92 61 93 
<< m2 >>
rect 61 92 62 93 
<< m1 >>
rect 62 92 63 93 
<< m2 >>
rect 62 92 63 93 
<< m2 >>
rect 63 92 64 93 
<< m1 >>
rect 64 92 65 93 
<< m2 >>
rect 64 92 65 93 
<< m2c >>
rect 64 92 65 93 
<< m1 >>
rect 64 92 65 93 
<< m2 >>
rect 64 92 65 93 
<< m1 >>
rect 67 92 68 93 
<< m1 >>
rect 73 92 74 93 
<< m2 >>
rect 81 92 82 93 
<< m2 >>
rect 82 92 83 93 
<< m2 >>
rect 105 92 106 93 
<< m1 >>
rect 106 92 107 93 
<< m2 >>
rect 106 92 107 93 
<< m2 >>
rect 107 92 108 93 
<< m1 >>
rect 108 92 109 93 
<< m2 >>
rect 108 92 109 93 
<< m2c >>
rect 108 92 109 93 
<< m1 >>
rect 108 92 109 93 
<< m2 >>
rect 108 92 109 93 
<< m1 >>
rect 109 92 110 93 
<< m1 >>
rect 110 92 111 93 
<< m2 >>
rect 110 92 111 93 
<< m1 >>
rect 111 92 112 93 
<< m2 >>
rect 111 92 112 93 
<< m1 >>
rect 112 92 113 93 
<< m2 >>
rect 112 92 113 93 
<< m1 >>
rect 113 92 114 93 
<< m2 >>
rect 113 92 114 93 
<< m2 >>
rect 114 92 115 93 
<< m1 >>
rect 115 92 116 93 
<< m2 >>
rect 115 92 116 93 
<< m2c >>
rect 115 92 116 93 
<< m1 >>
rect 115 92 116 93 
<< m2 >>
rect 115 92 116 93 
<< m1 >>
rect 116 92 117 93 
<< m1 >>
rect 117 92 118 93 
<< m1 >>
rect 136 92 137 93 
<< m1 >>
rect 151 92 152 93 
<< m2 >>
rect 151 92 152 93 
<< m2c >>
rect 151 92 152 93 
<< m1 >>
rect 151 92 152 93 
<< m2 >>
rect 151 92 152 93 
<< m1 >>
rect 153 92 154 93 
<< m2 >>
rect 153 92 154 93 
<< m2c >>
rect 153 92 154 93 
<< m1 >>
rect 153 92 154 93 
<< m2 >>
rect 153 92 154 93 
<< m1 >>
rect 159 92 160 93 
<< m2 >>
rect 159 92 160 93 
<< m2c >>
rect 159 92 160 93 
<< m1 >>
rect 159 92 160 93 
<< m2 >>
rect 159 92 160 93 
<< m1 >>
rect 160 92 161 93 
<< m1 >>
rect 161 92 162 93 
<< m2 >>
rect 161 92 162 93 
<< m2c >>
rect 161 92 162 93 
<< m1 >>
rect 161 92 162 93 
<< m2 >>
rect 161 92 162 93 
<< m2 >>
rect 162 92 163 93 
<< m1 >>
rect 163 92 164 93 
<< m2 >>
rect 163 92 164 93 
<< m1 >>
rect 167 92 168 93 
<< m2 >>
rect 167 92 168 93 
<< m2c >>
rect 167 92 168 93 
<< m1 >>
rect 167 92 168 93 
<< m2 >>
rect 167 92 168 93 
<< m2 >>
rect 169 92 170 93 
<< m2 >>
rect 171 92 172 93 
<< m1 >>
rect 178 92 179 93 
<< m1 >>
rect 10 93 11 94 
<< m2 >>
rect 10 93 11 94 
<< m1 >>
rect 19 93 20 94 
<< m1 >>
rect 22 93 23 94 
<< m1 >>
rect 26 93 27 94 
<< m1 >>
rect 28 93 29 94 
<< m1 >>
rect 37 93 38 94 
<< m2 >>
rect 38 93 39 94 
<< m1 >>
rect 39 93 40 94 
<< m2 >>
rect 39 93 40 94 
<< m2c >>
rect 39 93 40 94 
<< m1 >>
rect 39 93 40 94 
<< m2 >>
rect 39 93 40 94 
<< m1 >>
rect 40 93 41 94 
<< m1 >>
rect 41 93 42 94 
<< m1 >>
rect 42 93 43 94 
<< m1 >>
rect 43 93 44 94 
<< m1 >>
rect 45 93 46 94 
<< m1 >>
rect 52 93 53 94 
<< m1 >>
rect 54 93 55 94 
<< m1 >>
rect 58 93 59 94 
<< m1 >>
rect 62 93 63 94 
<< m1 >>
rect 67 93 68 94 
<< m2 >>
rect 68 93 69 94 
<< m1 >>
rect 69 93 70 94 
<< m2 >>
rect 69 93 70 94 
<< m2c >>
rect 69 93 70 94 
<< m1 >>
rect 69 93 70 94 
<< m2 >>
rect 69 93 70 94 
<< m1 >>
rect 70 93 71 94 
<< m1 >>
rect 71 93 72 94 
<< m2 >>
rect 71 93 72 94 
<< m2c >>
rect 71 93 72 94 
<< m1 >>
rect 71 93 72 94 
<< m2 >>
rect 71 93 72 94 
<< m2 >>
rect 72 93 73 94 
<< m1 >>
rect 73 93 74 94 
<< m2 >>
rect 73 93 74 94 
<< m2 >>
rect 74 93 75 94 
<< m1 >>
rect 75 93 76 94 
<< m2 >>
rect 75 93 76 94 
<< m2c >>
rect 75 93 76 94 
<< m1 >>
rect 75 93 76 94 
<< m2 >>
rect 75 93 76 94 
<< m1 >>
rect 76 93 77 94 
<< m1 >>
rect 77 93 78 94 
<< m1 >>
rect 78 93 79 94 
<< m1 >>
rect 79 93 80 94 
<< m1 >>
rect 80 93 81 94 
<< m1 >>
rect 81 93 82 94 
<< m2 >>
rect 81 93 82 94 
<< m1 >>
rect 82 93 83 94 
<< m1 >>
rect 83 93 84 94 
<< m1 >>
rect 84 93 85 94 
<< m2 >>
rect 105 93 106 94 
<< m1 >>
rect 106 93 107 94 
<< m2 >>
rect 110 93 111 94 
<< m1 >>
rect 136 93 137 94 
<< m2 >>
rect 151 93 152 94 
<< m2 >>
rect 153 93 154 94 
<< m2 >>
rect 159 93 160 94 
<< m1 >>
rect 163 93 164 94 
<< m2 >>
rect 167 93 168 94 
<< m2 >>
rect 169 93 170 94 
<< m2 >>
rect 171 93 172 94 
<< m1 >>
rect 178 93 179 94 
<< m1 >>
rect 10 94 11 95 
<< m2 >>
rect 10 94 11 95 
<< m2 >>
rect 11 94 12 95 
<< m1 >>
rect 12 94 13 95 
<< m2 >>
rect 12 94 13 95 
<< m2c >>
rect 12 94 13 95 
<< m1 >>
rect 12 94 13 95 
<< m2 >>
rect 12 94 13 95 
<< m1 >>
rect 13 94 14 95 
<< m1 >>
rect 14 94 15 95 
<< m1 >>
rect 15 94 16 95 
<< m1 >>
rect 16 94 17 95 
<< m1 >>
rect 17 94 18 95 
<< m2 >>
rect 17 94 18 95 
<< m2c >>
rect 17 94 18 95 
<< m1 >>
rect 17 94 18 95 
<< m2 >>
rect 17 94 18 95 
<< m2 >>
rect 18 94 19 95 
<< m1 >>
rect 19 94 20 95 
<< m2 >>
rect 19 94 20 95 
<< m2 >>
rect 20 94 21 95 
<< m2 >>
rect 21 94 22 95 
<< m1 >>
rect 22 94 23 95 
<< m2 >>
rect 22 94 23 95 
<< m2 >>
rect 23 94 24 95 
<< m1 >>
rect 24 94 25 95 
<< m2 >>
rect 24 94 25 95 
<< m2c >>
rect 24 94 25 95 
<< m1 >>
rect 24 94 25 95 
<< m2 >>
rect 24 94 25 95 
<< m2 >>
rect 25 94 26 95 
<< m1 >>
rect 26 94 27 95 
<< m2 >>
rect 26 94 27 95 
<< m2 >>
rect 27 94 28 95 
<< m1 >>
rect 28 94 29 95 
<< m2 >>
rect 28 94 29 95 
<< m2 >>
rect 29 94 30 95 
<< m1 >>
rect 30 94 31 95 
<< m2 >>
rect 30 94 31 95 
<< m2c >>
rect 30 94 31 95 
<< m1 >>
rect 30 94 31 95 
<< m2 >>
rect 30 94 31 95 
<< m1 >>
rect 31 94 32 95 
<< m1 >>
rect 32 94 33 95 
<< m2 >>
rect 32 94 33 95 
<< m2c >>
rect 32 94 33 95 
<< m1 >>
rect 32 94 33 95 
<< m2 >>
rect 32 94 33 95 
<< m2 >>
rect 33 94 34 95 
<< m2 >>
rect 34 94 35 95 
<< m2 >>
rect 35 94 36 95 
<< m2 >>
rect 36 94 37 95 
<< m1 >>
rect 37 94 38 95 
<< m2 >>
rect 37 94 38 95 
<< m2 >>
rect 38 94 39 95 
<< m1 >>
rect 45 94 46 95 
<< m1 >>
rect 52 94 53 95 
<< m1 >>
rect 54 94 55 95 
<< m1 >>
rect 56 94 57 95 
<< m2 >>
rect 56 94 57 95 
<< m2c >>
rect 56 94 57 95 
<< m1 >>
rect 56 94 57 95 
<< m2 >>
rect 56 94 57 95 
<< m2 >>
rect 57 94 58 95 
<< m1 >>
rect 58 94 59 95 
<< m2 >>
rect 58 94 59 95 
<< m2 >>
rect 59 94 60 95 
<< m1 >>
rect 60 94 61 95 
<< m2 >>
rect 60 94 61 95 
<< m2c >>
rect 60 94 61 95 
<< m1 >>
rect 60 94 61 95 
<< m2 >>
rect 60 94 61 95 
<< m2 >>
rect 61 94 62 95 
<< m1 >>
rect 62 94 63 95 
<< m2 >>
rect 62 94 63 95 
<< m2 >>
rect 63 94 64 95 
<< m1 >>
rect 64 94 65 95 
<< m2 >>
rect 64 94 65 95 
<< m1 >>
rect 65 94 66 95 
<< m2 >>
rect 65 94 66 95 
<< m2c >>
rect 65 94 66 95 
<< m1 >>
rect 65 94 66 95 
<< m2 >>
rect 65 94 66 95 
<< m2 >>
rect 66 94 67 95 
<< m1 >>
rect 67 94 68 95 
<< m2 >>
rect 67 94 68 95 
<< m2 >>
rect 68 94 69 95 
<< m1 >>
rect 73 94 74 95 
<< m2 >>
rect 81 94 82 95 
<< m1 >>
rect 84 94 85 95 
<< m2 >>
rect 105 94 106 95 
<< m1 >>
rect 106 94 107 95 
<< m1 >>
rect 107 94 108 95 
<< m1 >>
rect 108 94 109 95 
<< m1 >>
rect 109 94 110 95 
<< m1 >>
rect 110 94 111 95 
<< m2 >>
rect 110 94 111 95 
<< m1 >>
rect 111 94 112 95 
<< m1 >>
rect 112 94 113 95 
<< m1 >>
rect 113 94 114 95 
<< m1 >>
rect 114 94 115 95 
<< m1 >>
rect 115 94 116 95 
<< m1 >>
rect 116 94 117 95 
<< m1 >>
rect 117 94 118 95 
<< m1 >>
rect 118 94 119 95 
<< m1 >>
rect 119 94 120 95 
<< m1 >>
rect 120 94 121 95 
<< m1 >>
rect 121 94 122 95 
<< m1 >>
rect 122 94 123 95 
<< m1 >>
rect 123 94 124 95 
<< m1 >>
rect 124 94 125 95 
<< m1 >>
rect 136 94 137 95 
<< m1 >>
rect 137 94 138 95 
<< m1 >>
rect 138 94 139 95 
<< m1 >>
rect 139 94 140 95 
<< m1 >>
rect 140 94 141 95 
<< m1 >>
rect 141 94 142 95 
<< m1 >>
rect 142 94 143 95 
<< m1 >>
rect 143 94 144 95 
<< m1 >>
rect 144 94 145 95 
<< m1 >>
rect 145 94 146 95 
<< m1 >>
rect 146 94 147 95 
<< m1 >>
rect 147 94 148 95 
<< m1 >>
rect 148 94 149 95 
<< m1 >>
rect 149 94 150 95 
<< m1 >>
rect 150 94 151 95 
<< m1 >>
rect 151 94 152 95 
<< m2 >>
rect 151 94 152 95 
<< m1 >>
rect 152 94 153 95 
<< m1 >>
rect 153 94 154 95 
<< m2 >>
rect 153 94 154 95 
<< m1 >>
rect 154 94 155 95 
<< m1 >>
rect 155 94 156 95 
<< m1 >>
rect 156 94 157 95 
<< m1 >>
rect 157 94 158 95 
<< m1 >>
rect 158 94 159 95 
<< m1 >>
rect 159 94 160 95 
<< m2 >>
rect 159 94 160 95 
<< m1 >>
rect 160 94 161 95 
<< m1 >>
rect 161 94 162 95 
<< m2 >>
rect 161 94 162 95 
<< m2c >>
rect 161 94 162 95 
<< m1 >>
rect 161 94 162 95 
<< m2 >>
rect 161 94 162 95 
<< m2 >>
rect 162 94 163 95 
<< m1 >>
rect 163 94 164 95 
<< m2 >>
rect 163 94 164 95 
<< m2 >>
rect 164 94 165 95 
<< m1 >>
rect 165 94 166 95 
<< m2 >>
rect 165 94 166 95 
<< m2c >>
rect 165 94 166 95 
<< m1 >>
rect 165 94 166 95 
<< m2 >>
rect 165 94 166 95 
<< m1 >>
rect 166 94 167 95 
<< m1 >>
rect 167 94 168 95 
<< m2 >>
rect 167 94 168 95 
<< m1 >>
rect 168 94 169 95 
<< m1 >>
rect 169 94 170 95 
<< m2 >>
rect 169 94 170 95 
<< m1 >>
rect 170 94 171 95 
<< m1 >>
rect 171 94 172 95 
<< m2 >>
rect 171 94 172 95 
<< m1 >>
rect 172 94 173 95 
<< m1 >>
rect 173 94 174 95 
<< m1 >>
rect 174 94 175 95 
<< m1 >>
rect 175 94 176 95 
<< m1 >>
rect 176 94 177 95 
<< m1 >>
rect 177 94 178 95 
<< m1 >>
rect 178 94 179 95 
<< m1 >>
rect 10 95 11 96 
<< m1 >>
rect 19 95 20 96 
<< m1 >>
rect 22 95 23 96 
<< m1 >>
rect 26 95 27 96 
<< m1 >>
rect 28 95 29 96 
<< m1 >>
rect 34 95 35 96 
<< m1 >>
rect 35 95 36 96 
<< m1 >>
rect 36 95 37 96 
<< m1 >>
rect 37 95 38 96 
<< m1 >>
rect 45 95 46 96 
<< m2 >>
rect 45 95 46 96 
<< m2c >>
rect 45 95 46 96 
<< m1 >>
rect 45 95 46 96 
<< m2 >>
rect 45 95 46 96 
<< m1 >>
rect 52 95 53 96 
<< m1 >>
rect 54 95 55 96 
<< m1 >>
rect 56 95 57 96 
<< m1 >>
rect 58 95 59 96 
<< m1 >>
rect 62 95 63 96 
<< m1 >>
rect 67 95 68 96 
<< m1 >>
rect 68 95 69 96 
<< m1 >>
rect 69 95 70 96 
<< m1 >>
rect 70 95 71 96 
<< m2 >>
rect 70 95 71 96 
<< m2c >>
rect 70 95 71 96 
<< m1 >>
rect 70 95 71 96 
<< m2 >>
rect 70 95 71 96 
<< m1 >>
rect 73 95 74 96 
<< m2 >>
rect 73 95 74 96 
<< m2c >>
rect 73 95 74 96 
<< m1 >>
rect 73 95 74 96 
<< m2 >>
rect 73 95 74 96 
<< m1 >>
rect 81 95 82 96 
<< m2 >>
rect 81 95 82 96 
<< m2c >>
rect 81 95 82 96 
<< m1 >>
rect 81 95 82 96 
<< m2 >>
rect 81 95 82 96 
<< m2 >>
rect 83 95 84 96 
<< m1 >>
rect 84 95 85 96 
<< m2 >>
rect 84 95 85 96 
<< m1 >>
rect 85 95 86 96 
<< m2 >>
rect 85 95 86 96 
<< m1 >>
rect 86 95 87 96 
<< m2 >>
rect 86 95 87 96 
<< m1 >>
rect 87 95 88 96 
<< m2 >>
rect 87 95 88 96 
<< m1 >>
rect 88 95 89 96 
<< m2 >>
rect 88 95 89 96 
<< m1 >>
rect 89 95 90 96 
<< m2 >>
rect 89 95 90 96 
<< m1 >>
rect 90 95 91 96 
<< m2 >>
rect 90 95 91 96 
<< m1 >>
rect 91 95 92 96 
<< m2 >>
rect 91 95 92 96 
<< m1 >>
rect 92 95 93 96 
<< m2 >>
rect 92 95 93 96 
<< m1 >>
rect 93 95 94 96 
<< m2 >>
rect 93 95 94 96 
<< m1 >>
rect 94 95 95 96 
<< m2 >>
rect 94 95 95 96 
<< m1 >>
rect 95 95 96 96 
<< m2 >>
rect 95 95 96 96 
<< m1 >>
rect 96 95 97 96 
<< m2 >>
rect 96 95 97 96 
<< m1 >>
rect 97 95 98 96 
<< m2 >>
rect 97 95 98 96 
<< m1 >>
rect 98 95 99 96 
<< m2 >>
rect 98 95 99 96 
<< m1 >>
rect 99 95 100 96 
<< m2 >>
rect 99 95 100 96 
<< m1 >>
rect 100 95 101 96 
<< m2 >>
rect 100 95 101 96 
<< m1 >>
rect 101 95 102 96 
<< m2 >>
rect 101 95 102 96 
<< m1 >>
rect 102 95 103 96 
<< m2 >>
rect 102 95 103 96 
<< m1 >>
rect 103 95 104 96 
<< m2 >>
rect 103 95 104 96 
<< m2 >>
rect 104 95 105 96 
<< m2 >>
rect 105 95 106 96 
<< m2 >>
rect 107 95 108 96 
<< m2 >>
rect 108 95 109 96 
<< m2 >>
rect 109 95 110 96 
<< m2 >>
rect 110 95 111 96 
<< m1 >>
rect 124 95 125 96 
<< m2 >>
rect 151 95 152 96 
<< m2 >>
rect 153 95 154 96 
<< m2 >>
rect 159 95 160 96 
<< m1 >>
rect 163 95 164 96 
<< m2 >>
rect 167 95 168 96 
<< m2 >>
rect 169 95 170 96 
<< m2 >>
rect 171 95 172 96 
<< m1 >>
rect 10 96 11 97 
<< m1 >>
rect 19 96 20 97 
<< m1 >>
rect 22 96 23 97 
<< m1 >>
rect 26 96 27 97 
<< m1 >>
rect 28 96 29 97 
<< m1 >>
rect 34 96 35 97 
<< m2 >>
rect 45 96 46 97 
<< m1 >>
rect 52 96 53 97 
<< m1 >>
rect 54 96 55 97 
<< m1 >>
rect 56 96 57 97 
<< m1 >>
rect 58 96 59 97 
<< m1 >>
rect 62 96 63 97 
<< m2 >>
rect 70 96 71 97 
<< m2 >>
rect 73 96 74 97 
<< m2 >>
rect 75 96 76 97 
<< m2 >>
rect 76 96 77 97 
<< m2 >>
rect 77 96 78 97 
<< m2 >>
rect 78 96 79 97 
<< m2 >>
rect 79 96 80 97 
<< m2 >>
rect 80 96 81 97 
<< m2 >>
rect 81 96 82 97 
<< m2 >>
rect 83 96 84 97 
<< m1 >>
rect 103 96 104 97 
<< m1 >>
rect 107 96 108 97 
<< m2 >>
rect 107 96 108 97 
<< m2c >>
rect 107 96 108 97 
<< m1 >>
rect 107 96 108 97 
<< m2 >>
rect 107 96 108 97 
<< m1 >>
rect 124 96 125 97 
<< m1 >>
rect 151 96 152 97 
<< m2 >>
rect 151 96 152 97 
<< m2c >>
rect 151 96 152 97 
<< m1 >>
rect 151 96 152 97 
<< m2 >>
rect 151 96 152 97 
<< m1 >>
rect 153 96 154 97 
<< m2 >>
rect 153 96 154 97 
<< m2c >>
rect 153 96 154 97 
<< m1 >>
rect 153 96 154 97 
<< m2 >>
rect 153 96 154 97 
<< m1 >>
rect 159 96 160 97 
<< m2 >>
rect 159 96 160 97 
<< m2c >>
rect 159 96 160 97 
<< m1 >>
rect 159 96 160 97 
<< m2 >>
rect 159 96 160 97 
<< m1 >>
rect 163 96 164 97 
<< m1 >>
rect 167 96 168 97 
<< m2 >>
rect 167 96 168 97 
<< m2c >>
rect 167 96 168 97 
<< m1 >>
rect 167 96 168 97 
<< m2 >>
rect 167 96 168 97 
<< m1 >>
rect 169 96 170 97 
<< m2 >>
rect 169 96 170 97 
<< m2c >>
rect 169 96 170 97 
<< m1 >>
rect 169 96 170 97 
<< m2 >>
rect 169 96 170 97 
<< m1 >>
rect 171 96 172 97 
<< m2 >>
rect 171 96 172 97 
<< m2c >>
rect 171 96 172 97 
<< m1 >>
rect 171 96 172 97 
<< m2 >>
rect 171 96 172 97 
<< m1 >>
rect 10 97 11 98 
<< m1 >>
rect 19 97 20 98 
<< m1 >>
rect 22 97 23 98 
<< m1 >>
rect 26 97 27 98 
<< m1 >>
rect 28 97 29 98 
<< m1 >>
rect 34 97 35 98 
<< m1 >>
rect 37 97 38 98 
<< m1 >>
rect 38 97 39 98 
<< m1 >>
rect 39 97 40 98 
<< m1 >>
rect 40 97 41 98 
<< m1 >>
rect 41 97 42 98 
<< m1 >>
rect 42 97 43 98 
<< m1 >>
rect 43 97 44 98 
<< m1 >>
rect 44 97 45 98 
<< m1 >>
rect 45 97 46 98 
<< m2 >>
rect 45 97 46 98 
<< m1 >>
rect 46 97 47 98 
<< m1 >>
rect 47 97 48 98 
<< m1 >>
rect 48 97 49 98 
<< m1 >>
rect 49 97 50 98 
<< m1 >>
rect 50 97 51 98 
<< m2 >>
rect 50 97 51 98 
<< m2c >>
rect 50 97 51 98 
<< m1 >>
rect 50 97 51 98 
<< m2 >>
rect 50 97 51 98 
<< m2 >>
rect 51 97 52 98 
<< m1 >>
rect 52 97 53 98 
<< m2 >>
rect 52 97 53 98 
<< m2 >>
rect 53 97 54 98 
<< m1 >>
rect 54 97 55 98 
<< m2 >>
rect 54 97 55 98 
<< m2c >>
rect 54 97 55 98 
<< m1 >>
rect 54 97 55 98 
<< m2 >>
rect 54 97 55 98 
<< m1 >>
rect 56 97 57 98 
<< m2 >>
rect 56 97 57 98 
<< m2c >>
rect 56 97 57 98 
<< m1 >>
rect 56 97 57 98 
<< m2 >>
rect 56 97 57 98 
<< m1 >>
rect 58 97 59 98 
<< m2 >>
rect 58 97 59 98 
<< m2c >>
rect 58 97 59 98 
<< m1 >>
rect 58 97 59 98 
<< m2 >>
rect 58 97 59 98 
<< m1 >>
rect 62 97 63 98 
<< m1 >>
rect 64 97 65 98 
<< m1 >>
rect 65 97 66 98 
<< m1 >>
rect 66 97 67 98 
<< m1 >>
rect 67 97 68 98 
<< m1 >>
rect 68 97 69 98 
<< m1 >>
rect 69 97 70 98 
<< m1 >>
rect 70 97 71 98 
<< m2 >>
rect 70 97 71 98 
<< m1 >>
rect 71 97 72 98 
<< m1 >>
rect 72 97 73 98 
<< m1 >>
rect 73 97 74 98 
<< m2 >>
rect 73 97 74 98 
<< m1 >>
rect 74 97 75 98 
<< m1 >>
rect 75 97 76 98 
<< m2 >>
rect 75 97 76 98 
<< m1 >>
rect 76 97 77 98 
<< m1 >>
rect 77 97 78 98 
<< m1 >>
rect 78 97 79 98 
<< m1 >>
rect 79 97 80 98 
<< m1 >>
rect 80 97 81 98 
<< m1 >>
rect 81 97 82 98 
<< m1 >>
rect 82 97 83 98 
<< m1 >>
rect 83 97 84 98 
<< m2 >>
rect 83 97 84 98 
<< m1 >>
rect 84 97 85 98 
<< m1 >>
rect 85 97 86 98 
<< m1 >>
rect 86 97 87 98 
<< m1 >>
rect 87 97 88 98 
<< m1 >>
rect 88 97 89 98 
<< m2 >>
rect 102 97 103 98 
<< m1 >>
rect 103 97 104 98 
<< m2 >>
rect 103 97 104 98 
<< m2 >>
rect 104 97 105 98 
<< m1 >>
rect 105 97 106 98 
<< m2 >>
rect 105 97 106 98 
<< m2c >>
rect 105 97 106 98 
<< m1 >>
rect 105 97 106 98 
<< m2 >>
rect 105 97 106 98 
<< m1 >>
rect 106 97 107 98 
<< m1 >>
rect 107 97 108 98 
<< m1 >>
rect 124 97 125 98 
<< m1 >>
rect 151 97 152 98 
<< m1 >>
rect 153 97 154 98 
<< m1 >>
rect 159 97 160 98 
<< m1 >>
rect 163 97 164 98 
<< m1 >>
rect 167 97 168 98 
<< m1 >>
rect 169 97 170 98 
<< m1 >>
rect 171 97 172 98 
<< m1 >>
rect 10 98 11 99 
<< m1 >>
rect 19 98 20 99 
<< m1 >>
rect 22 98 23 99 
<< m1 >>
rect 26 98 27 99 
<< m1 >>
rect 28 98 29 99 
<< m1 >>
rect 34 98 35 99 
<< m1 >>
rect 37 98 38 99 
<< m2 >>
rect 45 98 46 99 
<< m1 >>
rect 52 98 53 99 
<< m2 >>
rect 56 98 57 99 
<< m2 >>
rect 58 98 59 99 
<< m1 >>
rect 62 98 63 99 
<< m1 >>
rect 64 98 65 99 
<< m2 >>
rect 70 98 71 99 
<< m2 >>
rect 73 98 74 99 
<< m2 >>
rect 75 98 76 99 
<< m2 >>
rect 77 98 78 99 
<< m2 >>
rect 78 98 79 99 
<< m2 >>
rect 79 98 80 99 
<< m2 >>
rect 80 98 81 99 
<< m2 >>
rect 81 98 82 99 
<< m2 >>
rect 82 98 83 99 
<< m2 >>
rect 83 98 84 99 
<< m1 >>
rect 88 98 89 99 
<< m2 >>
rect 102 98 103 99 
<< m1 >>
rect 103 98 104 99 
<< m1 >>
rect 124 98 125 99 
<< m1 >>
rect 151 98 152 99 
<< m1 >>
rect 153 98 154 99 
<< m1 >>
rect 159 98 160 99 
<< m1 >>
rect 160 98 161 99 
<< m1 >>
rect 161 98 162 99 
<< m2 >>
rect 161 98 162 99 
<< m2c >>
rect 161 98 162 99 
<< m1 >>
rect 161 98 162 99 
<< m2 >>
rect 161 98 162 99 
<< m2 >>
rect 162 98 163 99 
<< m1 >>
rect 163 98 164 99 
<< m2 >>
rect 163 98 164 99 
<< m2 >>
rect 164 98 165 99 
<< m1 >>
rect 165 98 166 99 
<< m2 >>
rect 165 98 166 99 
<< m2c >>
rect 165 98 166 99 
<< m1 >>
rect 165 98 166 99 
<< m2 >>
rect 165 98 166 99 
<< m2 >>
rect 166 98 167 99 
<< m1 >>
rect 167 98 168 99 
<< m2 >>
rect 167 98 168 99 
<< m2 >>
rect 168 98 169 99 
<< m1 >>
rect 169 98 170 99 
<< m2 >>
rect 169 98 170 99 
<< m2 >>
rect 170 98 171 99 
<< m1 >>
rect 171 98 172 99 
<< m2 >>
rect 171 98 172 99 
<< m2c >>
rect 171 98 172 99 
<< m1 >>
rect 171 98 172 99 
<< m2 >>
rect 171 98 172 99 
<< m1 >>
rect 10 99 11 100 
<< m1 >>
rect 13 99 14 100 
<< m1 >>
rect 14 99 15 100 
<< m1 >>
rect 15 99 16 100 
<< m1 >>
rect 16 99 17 100 
<< m1 >>
rect 17 99 18 100 
<< m1 >>
rect 18 99 19 100 
<< m1 >>
rect 19 99 20 100 
<< m1 >>
rect 22 99 23 100 
<< m1 >>
rect 26 99 27 100 
<< m1 >>
rect 28 99 29 100 
<< m1 >>
rect 34 99 35 100 
<< m1 >>
rect 37 99 38 100 
<< m1 >>
rect 45 99 46 100 
<< m2 >>
rect 45 99 46 100 
<< m2c >>
rect 45 99 46 100 
<< m1 >>
rect 45 99 46 100 
<< m2 >>
rect 45 99 46 100 
<< m1 >>
rect 52 99 53 100 
<< m1 >>
rect 53 99 54 100 
<< m1 >>
rect 54 99 55 100 
<< m1 >>
rect 55 99 56 100 
<< m1 >>
rect 56 99 57 100 
<< m2 >>
rect 56 99 57 100 
<< m1 >>
rect 57 99 58 100 
<< m1 >>
rect 58 99 59 100 
<< m2 >>
rect 58 99 59 100 
<< m1 >>
rect 59 99 60 100 
<< m1 >>
rect 60 99 61 100 
<< m1 >>
rect 62 99 63 100 
<< m1 >>
rect 64 99 65 100 
<< m1 >>
rect 70 99 71 100 
<< m2 >>
rect 70 99 71 100 
<< m2c >>
rect 70 99 71 100 
<< m1 >>
rect 70 99 71 100 
<< m2 >>
rect 70 99 71 100 
<< m1 >>
rect 73 99 74 100 
<< m2 >>
rect 73 99 74 100 
<< m2c >>
rect 73 99 74 100 
<< m1 >>
rect 73 99 74 100 
<< m2 >>
rect 73 99 74 100 
<< m1 >>
rect 75 99 76 100 
<< m2 >>
rect 75 99 76 100 
<< m2c >>
rect 75 99 76 100 
<< m1 >>
rect 75 99 76 100 
<< m2 >>
rect 75 99 76 100 
<< m1 >>
rect 77 99 78 100 
<< m2 >>
rect 77 99 78 100 
<< m2c >>
rect 77 99 78 100 
<< m1 >>
rect 77 99 78 100 
<< m2 >>
rect 77 99 78 100 
<< m1 >>
rect 88 99 89 100 
<< m2 >>
rect 102 99 103 100 
<< m1 >>
rect 103 99 104 100 
<< m1 >>
rect 124 99 125 100 
<< m1 >>
rect 151 99 152 100 
<< m1 >>
rect 153 99 154 100 
<< m1 >>
rect 163 99 164 100 
<< m1 >>
rect 167 99 168 100 
<< m1 >>
rect 169 99 170 100 
<< m1 >>
rect 10 100 11 101 
<< m1 >>
rect 13 100 14 101 
<< m1 >>
rect 22 100 23 101 
<< m2 >>
rect 25 100 26 101 
<< m1 >>
rect 26 100 27 101 
<< m2 >>
rect 26 100 27 101 
<< m2 >>
rect 27 100 28 101 
<< m1 >>
rect 28 100 29 101 
<< m2 >>
rect 28 100 29 101 
<< m2 >>
rect 29 100 30 101 
<< m1 >>
rect 30 100 31 101 
<< m2 >>
rect 30 100 31 101 
<< m2c >>
rect 30 100 31 101 
<< m1 >>
rect 30 100 31 101 
<< m2 >>
rect 30 100 31 101 
<< m1 >>
rect 31 100 32 101 
<< m1 >>
rect 34 100 35 101 
<< m1 >>
rect 37 100 38 101 
<< m1 >>
rect 45 100 46 101 
<< m2 >>
rect 56 100 57 101 
<< m2 >>
rect 58 100 59 101 
<< m1 >>
rect 60 100 61 101 
<< m1 >>
rect 62 100 63 101 
<< m1 >>
rect 64 100 65 101 
<< m1 >>
rect 70 100 71 101 
<< m1 >>
rect 73 100 74 101 
<< m1 >>
rect 75 100 76 101 
<< m1 >>
rect 77 100 78 101 
<< m1 >>
rect 81 100 82 101 
<< m1 >>
rect 82 100 83 101 
<< m1 >>
rect 83 100 84 101 
<< m1 >>
rect 84 100 85 101 
<< m1 >>
rect 85 100 86 101 
<< m1 >>
rect 88 100 89 101 
<< m1 >>
rect 93 100 94 101 
<< m1 >>
rect 94 100 95 101 
<< m1 >>
rect 95 100 96 101 
<< m1 >>
rect 96 100 97 101 
<< m1 >>
rect 97 100 98 101 
<< m1 >>
rect 98 100 99 101 
<< m1 >>
rect 99 100 100 101 
<< m1 >>
rect 100 100 101 101 
<< m1 >>
rect 101 100 102 101 
<< m2 >>
rect 101 100 102 101 
<< m2c >>
rect 101 100 102 101 
<< m1 >>
rect 101 100 102 101 
<< m2 >>
rect 101 100 102 101 
<< m2 >>
rect 102 100 103 101 
<< m1 >>
rect 103 100 104 101 
<< m1 >>
rect 124 100 125 101 
<< m1 >>
rect 151 100 152 101 
<< m1 >>
rect 153 100 154 101 
<< m1 >>
rect 163 100 164 101 
<< m1 >>
rect 167 100 168 101 
<< m1 >>
rect 169 100 170 101 
<< m1 >>
rect 10 101 11 102 
<< m1 >>
rect 13 101 14 102 
<< m1 >>
rect 22 101 23 102 
<< m2 >>
rect 25 101 26 102 
<< m1 >>
rect 26 101 27 102 
<< m1 >>
rect 28 101 29 102 
<< m1 >>
rect 31 101 32 102 
<< m1 >>
rect 34 101 35 102 
<< m1 >>
rect 37 101 38 102 
<< m1 >>
rect 45 101 46 102 
<< m1 >>
rect 56 101 57 102 
<< m2 >>
rect 56 101 57 102 
<< m2c >>
rect 56 101 57 102 
<< m1 >>
rect 56 101 57 102 
<< m2 >>
rect 56 101 57 102 
<< m1 >>
rect 58 101 59 102 
<< m2 >>
rect 58 101 59 102 
<< m2c >>
rect 58 101 59 102 
<< m1 >>
rect 58 101 59 102 
<< m2 >>
rect 58 101 59 102 
<< m1 >>
rect 60 101 61 102 
<< m1 >>
rect 62 101 63 102 
<< m1 >>
rect 64 101 65 102 
<< m1 >>
rect 70 101 71 102 
<< m1 >>
rect 73 101 74 102 
<< m1 >>
rect 75 101 76 102 
<< m2 >>
rect 75 101 76 102 
<< m2c >>
rect 75 101 76 102 
<< m1 >>
rect 75 101 76 102 
<< m2 >>
rect 75 101 76 102 
<< m2 >>
rect 76 101 77 102 
<< m1 >>
rect 77 101 78 102 
<< m2 >>
rect 77 101 78 102 
<< m2 >>
rect 78 101 79 102 
<< m1 >>
rect 79 101 80 102 
<< m2 >>
rect 79 101 80 102 
<< m2c >>
rect 79 101 80 102 
<< m1 >>
rect 79 101 80 102 
<< m2 >>
rect 79 101 80 102 
<< m1 >>
rect 81 101 82 102 
<< m1 >>
rect 85 101 86 102 
<< m1 >>
rect 88 101 89 102 
<< m1 >>
rect 93 101 94 102 
<< m1 >>
rect 103 101 104 102 
<< m1 >>
rect 124 101 125 102 
<< m1 >>
rect 151 101 152 102 
<< m1 >>
rect 153 101 154 102 
<< m1 >>
rect 163 101 164 102 
<< m1 >>
rect 167 101 168 102 
<< m1 >>
rect 169 101 170 102 
<< m1 >>
rect 10 102 11 103 
<< pdiffusion >>
rect 12 102 13 103 
<< m1 >>
rect 13 102 14 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< m1 >>
rect 22 102 23 103 
<< m2 >>
rect 25 102 26 103 
<< m1 >>
rect 26 102 27 103 
<< m1 >>
rect 28 102 29 103 
<< pdiffusion >>
rect 30 102 31 103 
<< m1 >>
rect 31 102 32 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< pdiffusion >>
rect 33 102 34 103 
<< m1 >>
rect 34 102 35 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< m1 >>
rect 37 102 38 103 
<< m1 >>
rect 45 102 46 103 
<< pdiffusion >>
rect 48 102 49 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m1 >>
rect 56 102 57 103 
<< m1 >>
rect 58 102 59 103 
<< m1 >>
rect 60 102 61 103 
<< m1 >>
rect 62 102 63 103 
<< m1 >>
rect 64 102 65 103 
<< pdiffusion >>
rect 66 102 67 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< m1 >>
rect 70 102 71 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< m1 >>
rect 73 102 74 103 
<< m1 >>
rect 77 102 78 103 
<< m1 >>
rect 79 102 80 103 
<< m1 >>
rect 81 102 82 103 
<< pdiffusion >>
rect 84 102 85 103 
<< m1 >>
rect 85 102 86 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< m1 >>
rect 88 102 89 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< m1 >>
rect 93 102 94 103 
<< pdiffusion >>
rect 102 102 103 103 
<< m1 >>
rect 103 102 104 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< pdiffusion >>
rect 120 102 121 103 
<< pdiffusion >>
rect 121 102 122 103 
<< pdiffusion >>
rect 122 102 123 103 
<< pdiffusion >>
rect 123 102 124 103 
<< m1 >>
rect 124 102 125 103 
<< pdiffusion >>
rect 124 102 125 103 
<< pdiffusion >>
rect 125 102 126 103 
<< pdiffusion >>
rect 138 102 139 103 
<< pdiffusion >>
rect 139 102 140 103 
<< pdiffusion >>
rect 140 102 141 103 
<< pdiffusion >>
rect 141 102 142 103 
<< pdiffusion >>
rect 142 102 143 103 
<< pdiffusion >>
rect 143 102 144 103 
<< m1 >>
rect 151 102 152 103 
<< m1 >>
rect 153 102 154 103 
<< pdiffusion >>
rect 156 102 157 103 
<< pdiffusion >>
rect 157 102 158 103 
<< pdiffusion >>
rect 158 102 159 103 
<< pdiffusion >>
rect 159 102 160 103 
<< pdiffusion >>
rect 160 102 161 103 
<< pdiffusion >>
rect 161 102 162 103 
<< m1 >>
rect 163 102 164 103 
<< m1 >>
rect 167 102 168 103 
<< m1 >>
rect 169 102 170 103 
<< pdiffusion >>
rect 174 102 175 103 
<< pdiffusion >>
rect 175 102 176 103 
<< pdiffusion >>
rect 176 102 177 103 
<< pdiffusion >>
rect 177 102 178 103 
<< pdiffusion >>
rect 178 102 179 103 
<< pdiffusion >>
rect 179 102 180 103 
<< m1 >>
rect 10 103 11 104 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< m1 >>
rect 22 103 23 104 
<< m2 >>
rect 25 103 26 104 
<< m1 >>
rect 26 103 27 104 
<< m1 >>
rect 28 103 29 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< m1 >>
rect 37 103 38 104 
<< m1 >>
rect 45 103 46 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m1 >>
rect 56 103 57 104 
<< m1 >>
rect 58 103 59 104 
<< m1 >>
rect 60 103 61 104 
<< m1 >>
rect 62 103 63 104 
<< m1 >>
rect 64 103 65 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< m1 >>
rect 73 103 74 104 
<< m1 >>
rect 77 103 78 104 
<< m1 >>
rect 79 103 80 104 
<< m1 >>
rect 81 103 82 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< m1 >>
rect 93 103 94 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< pdiffusion >>
rect 120 103 121 104 
<< pdiffusion >>
rect 121 103 122 104 
<< pdiffusion >>
rect 122 103 123 104 
<< pdiffusion >>
rect 123 103 124 104 
<< pdiffusion >>
rect 124 103 125 104 
<< pdiffusion >>
rect 125 103 126 104 
<< pdiffusion >>
rect 138 103 139 104 
<< pdiffusion >>
rect 139 103 140 104 
<< pdiffusion >>
rect 140 103 141 104 
<< pdiffusion >>
rect 141 103 142 104 
<< pdiffusion >>
rect 142 103 143 104 
<< pdiffusion >>
rect 143 103 144 104 
<< m1 >>
rect 151 103 152 104 
<< m1 >>
rect 153 103 154 104 
<< pdiffusion >>
rect 156 103 157 104 
<< pdiffusion >>
rect 157 103 158 104 
<< pdiffusion >>
rect 158 103 159 104 
<< pdiffusion >>
rect 159 103 160 104 
<< pdiffusion >>
rect 160 103 161 104 
<< pdiffusion >>
rect 161 103 162 104 
<< m1 >>
rect 163 103 164 104 
<< m1 >>
rect 167 103 168 104 
<< m1 >>
rect 169 103 170 104 
<< pdiffusion >>
rect 174 103 175 104 
<< pdiffusion >>
rect 175 103 176 104 
<< pdiffusion >>
rect 176 103 177 104 
<< pdiffusion >>
rect 177 103 178 104 
<< pdiffusion >>
rect 178 103 179 104 
<< pdiffusion >>
rect 179 103 180 104 
<< m1 >>
rect 10 104 11 105 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< m1 >>
rect 22 104 23 105 
<< m2 >>
rect 25 104 26 105 
<< m1 >>
rect 26 104 27 105 
<< m1 >>
rect 28 104 29 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< m1 >>
rect 37 104 38 105 
<< m1 >>
rect 45 104 46 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m1 >>
rect 56 104 57 105 
<< m1 >>
rect 58 104 59 105 
<< m1 >>
rect 60 104 61 105 
<< m1 >>
rect 62 104 63 105 
<< m1 >>
rect 64 104 65 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< m1 >>
rect 73 104 74 105 
<< m1 >>
rect 77 104 78 105 
<< m1 >>
rect 79 104 80 105 
<< m1 >>
rect 81 104 82 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< m1 >>
rect 93 104 94 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< pdiffusion >>
rect 120 104 121 105 
<< pdiffusion >>
rect 121 104 122 105 
<< pdiffusion >>
rect 122 104 123 105 
<< pdiffusion >>
rect 123 104 124 105 
<< pdiffusion >>
rect 124 104 125 105 
<< pdiffusion >>
rect 125 104 126 105 
<< pdiffusion >>
rect 138 104 139 105 
<< pdiffusion >>
rect 139 104 140 105 
<< pdiffusion >>
rect 140 104 141 105 
<< pdiffusion >>
rect 141 104 142 105 
<< pdiffusion >>
rect 142 104 143 105 
<< pdiffusion >>
rect 143 104 144 105 
<< m1 >>
rect 151 104 152 105 
<< m1 >>
rect 153 104 154 105 
<< pdiffusion >>
rect 156 104 157 105 
<< pdiffusion >>
rect 157 104 158 105 
<< pdiffusion >>
rect 158 104 159 105 
<< pdiffusion >>
rect 159 104 160 105 
<< pdiffusion >>
rect 160 104 161 105 
<< pdiffusion >>
rect 161 104 162 105 
<< m1 >>
rect 163 104 164 105 
<< m1 >>
rect 167 104 168 105 
<< m1 >>
rect 169 104 170 105 
<< pdiffusion >>
rect 174 104 175 105 
<< pdiffusion >>
rect 175 104 176 105 
<< pdiffusion >>
rect 176 104 177 105 
<< pdiffusion >>
rect 177 104 178 105 
<< pdiffusion >>
rect 178 104 179 105 
<< pdiffusion >>
rect 179 104 180 105 
<< m1 >>
rect 10 105 11 106 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< m1 >>
rect 22 105 23 106 
<< m2 >>
rect 25 105 26 106 
<< m1 >>
rect 26 105 27 106 
<< m1 >>
rect 28 105 29 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< m1 >>
rect 37 105 38 106 
<< m1 >>
rect 45 105 46 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m1 >>
rect 56 105 57 106 
<< m1 >>
rect 58 105 59 106 
<< m1 >>
rect 60 105 61 106 
<< m1 >>
rect 62 105 63 106 
<< m1 >>
rect 64 105 65 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< m1 >>
rect 73 105 74 106 
<< m1 >>
rect 77 105 78 106 
<< m1 >>
rect 79 105 80 106 
<< m1 >>
rect 81 105 82 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< m1 >>
rect 93 105 94 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< pdiffusion >>
rect 120 105 121 106 
<< pdiffusion >>
rect 121 105 122 106 
<< pdiffusion >>
rect 122 105 123 106 
<< pdiffusion >>
rect 123 105 124 106 
<< pdiffusion >>
rect 124 105 125 106 
<< pdiffusion >>
rect 125 105 126 106 
<< pdiffusion >>
rect 138 105 139 106 
<< pdiffusion >>
rect 139 105 140 106 
<< pdiffusion >>
rect 140 105 141 106 
<< pdiffusion >>
rect 141 105 142 106 
<< pdiffusion >>
rect 142 105 143 106 
<< pdiffusion >>
rect 143 105 144 106 
<< m1 >>
rect 151 105 152 106 
<< m1 >>
rect 153 105 154 106 
<< pdiffusion >>
rect 156 105 157 106 
<< pdiffusion >>
rect 157 105 158 106 
<< pdiffusion >>
rect 158 105 159 106 
<< pdiffusion >>
rect 159 105 160 106 
<< pdiffusion >>
rect 160 105 161 106 
<< pdiffusion >>
rect 161 105 162 106 
<< m1 >>
rect 163 105 164 106 
<< m1 >>
rect 167 105 168 106 
<< m1 >>
rect 169 105 170 106 
<< pdiffusion >>
rect 174 105 175 106 
<< pdiffusion >>
rect 175 105 176 106 
<< pdiffusion >>
rect 176 105 177 106 
<< pdiffusion >>
rect 177 105 178 106 
<< pdiffusion >>
rect 178 105 179 106 
<< pdiffusion >>
rect 179 105 180 106 
<< m1 >>
rect 10 106 11 107 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< m1 >>
rect 22 106 23 107 
<< m2 >>
rect 25 106 26 107 
<< m1 >>
rect 26 106 27 107 
<< m1 >>
rect 28 106 29 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< m1 >>
rect 37 106 38 107 
<< m1 >>
rect 45 106 46 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m1 >>
rect 56 106 57 107 
<< m1 >>
rect 58 106 59 107 
<< m1 >>
rect 60 106 61 107 
<< m1 >>
rect 62 106 63 107 
<< m1 >>
rect 64 106 65 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< m1 >>
rect 73 106 74 107 
<< m1 >>
rect 77 106 78 107 
<< m1 >>
rect 79 106 80 107 
<< m1 >>
rect 81 106 82 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< m1 >>
rect 93 106 94 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< pdiffusion >>
rect 120 106 121 107 
<< pdiffusion >>
rect 121 106 122 107 
<< pdiffusion >>
rect 122 106 123 107 
<< pdiffusion >>
rect 123 106 124 107 
<< pdiffusion >>
rect 124 106 125 107 
<< pdiffusion >>
rect 125 106 126 107 
<< pdiffusion >>
rect 138 106 139 107 
<< pdiffusion >>
rect 139 106 140 107 
<< pdiffusion >>
rect 140 106 141 107 
<< pdiffusion >>
rect 141 106 142 107 
<< pdiffusion >>
rect 142 106 143 107 
<< pdiffusion >>
rect 143 106 144 107 
<< m1 >>
rect 151 106 152 107 
<< m1 >>
rect 153 106 154 107 
<< pdiffusion >>
rect 156 106 157 107 
<< pdiffusion >>
rect 157 106 158 107 
<< pdiffusion >>
rect 158 106 159 107 
<< pdiffusion >>
rect 159 106 160 107 
<< pdiffusion >>
rect 160 106 161 107 
<< pdiffusion >>
rect 161 106 162 107 
<< m1 >>
rect 163 106 164 107 
<< m1 >>
rect 167 106 168 107 
<< m1 >>
rect 169 106 170 107 
<< pdiffusion >>
rect 174 106 175 107 
<< pdiffusion >>
rect 175 106 176 107 
<< pdiffusion >>
rect 176 106 177 107 
<< pdiffusion >>
rect 177 106 178 107 
<< pdiffusion >>
rect 178 106 179 107 
<< pdiffusion >>
rect 179 106 180 107 
<< m1 >>
rect 10 107 11 108 
<< pdiffusion >>
rect 12 107 13 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< m1 >>
rect 16 107 17 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< m1 >>
rect 22 107 23 108 
<< m2 >>
rect 22 107 23 108 
<< m2c >>
rect 22 107 23 108 
<< m1 >>
rect 22 107 23 108 
<< m2 >>
rect 22 107 23 108 
<< m2 >>
rect 25 107 26 108 
<< m1 >>
rect 26 107 27 108 
<< m1 >>
rect 28 107 29 108 
<< pdiffusion >>
rect 30 107 31 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< m1 >>
rect 34 107 35 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< m1 >>
rect 37 107 38 108 
<< m1 >>
rect 45 107 46 108 
<< pdiffusion >>
rect 48 107 49 108 
<< m1 >>
rect 49 107 50 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m1 >>
rect 56 107 57 108 
<< m1 >>
rect 58 107 59 108 
<< m1 >>
rect 60 107 61 108 
<< m1 >>
rect 62 107 63 108 
<< m1 >>
rect 64 107 65 108 
<< pdiffusion >>
rect 66 107 67 108 
<< m1 >>
rect 67 107 68 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< m1 >>
rect 70 107 71 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< m1 >>
rect 73 107 74 108 
<< m1 >>
rect 77 107 78 108 
<< m1 >>
rect 79 107 80 108 
<< m1 >>
rect 81 107 82 108 
<< pdiffusion >>
rect 84 107 85 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< m1 >>
rect 93 107 94 108 
<< pdiffusion >>
rect 102 107 103 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< m1 >>
rect 106 107 107 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< pdiffusion >>
rect 120 107 121 108 
<< pdiffusion >>
rect 121 107 122 108 
<< pdiffusion >>
rect 122 107 123 108 
<< pdiffusion >>
rect 123 107 124 108 
<< m1 >>
rect 124 107 125 108 
<< pdiffusion >>
rect 124 107 125 108 
<< pdiffusion >>
rect 125 107 126 108 
<< pdiffusion >>
rect 138 107 139 108 
<< pdiffusion >>
rect 139 107 140 108 
<< pdiffusion >>
rect 140 107 141 108 
<< pdiffusion >>
rect 141 107 142 108 
<< pdiffusion >>
rect 142 107 143 108 
<< pdiffusion >>
rect 143 107 144 108 
<< m1 >>
rect 151 107 152 108 
<< m1 >>
rect 153 107 154 108 
<< pdiffusion >>
rect 156 107 157 108 
<< pdiffusion >>
rect 157 107 158 108 
<< pdiffusion >>
rect 158 107 159 108 
<< pdiffusion >>
rect 159 107 160 108 
<< pdiffusion >>
rect 160 107 161 108 
<< pdiffusion >>
rect 161 107 162 108 
<< m1 >>
rect 163 107 164 108 
<< m1 >>
rect 167 107 168 108 
<< m1 >>
rect 169 107 170 108 
<< pdiffusion >>
rect 174 107 175 108 
<< pdiffusion >>
rect 175 107 176 108 
<< pdiffusion >>
rect 176 107 177 108 
<< pdiffusion >>
rect 177 107 178 108 
<< m1 >>
rect 178 107 179 108 
<< pdiffusion >>
rect 178 107 179 108 
<< pdiffusion >>
rect 179 107 180 108 
<< m1 >>
rect 10 108 11 109 
<< m1 >>
rect 16 108 17 109 
<< m2 >>
rect 22 108 23 109 
<< m2 >>
rect 25 108 26 109 
<< m1 >>
rect 26 108 27 109 
<< m1 >>
rect 28 108 29 109 
<< m1 >>
rect 34 108 35 109 
<< m1 >>
rect 37 108 38 109 
<< m1 >>
rect 45 108 46 109 
<< m1 >>
rect 49 108 50 109 
<< m1 >>
rect 56 108 57 109 
<< m2 >>
rect 56 108 57 109 
<< m2c >>
rect 56 108 57 109 
<< m1 >>
rect 56 108 57 109 
<< m2 >>
rect 56 108 57 109 
<< m1 >>
rect 58 108 59 109 
<< m2 >>
rect 58 108 59 109 
<< m2c >>
rect 58 108 59 109 
<< m1 >>
rect 58 108 59 109 
<< m2 >>
rect 58 108 59 109 
<< m1 >>
rect 60 108 61 109 
<< m2 >>
rect 60 108 61 109 
<< m2c >>
rect 60 108 61 109 
<< m1 >>
rect 60 108 61 109 
<< m2 >>
rect 60 108 61 109 
<< m2 >>
rect 61 108 62 109 
<< m1 >>
rect 62 108 63 109 
<< m2 >>
rect 62 108 63 109 
<< m2 >>
rect 63 108 64 109 
<< m1 >>
rect 64 108 65 109 
<< m2 >>
rect 64 108 65 109 
<< m1 >>
rect 67 108 68 109 
<< m1 >>
rect 70 108 71 109 
<< m2 >>
rect 70 108 71 109 
<< m2c >>
rect 70 108 71 109 
<< m1 >>
rect 70 108 71 109 
<< m2 >>
rect 70 108 71 109 
<< m1 >>
rect 73 108 74 109 
<< m1 >>
rect 77 108 78 109 
<< m1 >>
rect 79 108 80 109 
<< m1 >>
rect 81 108 82 109 
<< m1 >>
rect 93 108 94 109 
<< m1 >>
rect 106 108 107 109 
<< m1 >>
rect 124 108 125 109 
<< m1 >>
rect 151 108 152 109 
<< m1 >>
rect 153 108 154 109 
<< m1 >>
rect 163 108 164 109 
<< m1 >>
rect 167 108 168 109 
<< m1 >>
rect 169 108 170 109 
<< m1 >>
rect 178 108 179 109 
<< m1 >>
rect 10 109 11 110 
<< m1 >>
rect 16 109 17 110 
<< m1 >>
rect 17 109 18 110 
<< m1 >>
rect 18 109 19 110 
<< m1 >>
rect 19 109 20 110 
<< m1 >>
rect 20 109 21 110 
<< m1 >>
rect 21 109 22 110 
<< m1 >>
rect 22 109 23 110 
<< m2 >>
rect 22 109 23 110 
<< m1 >>
rect 23 109 24 110 
<< m1 >>
rect 24 109 25 110 
<< m1 >>
rect 25 109 26 110 
<< m2 >>
rect 25 109 26 110 
<< m1 >>
rect 26 109 27 110 
<< m1 >>
rect 28 109 29 110 
<< m1 >>
rect 34 109 35 110 
<< m1 >>
rect 35 109 36 110 
<< m1 >>
rect 36 109 37 110 
<< m1 >>
rect 37 109 38 110 
<< m1 >>
rect 45 109 46 110 
<< m1 >>
rect 49 109 50 110 
<< m2 >>
rect 56 109 57 110 
<< m2 >>
rect 58 109 59 110 
<< m1 >>
rect 62 109 63 110 
<< m1 >>
rect 64 109 65 110 
<< m2 >>
rect 64 109 65 110 
<< m1 >>
rect 67 109 68 110 
<< m2 >>
rect 70 109 71 110 
<< m2 >>
rect 71 109 72 110 
<< m2 >>
rect 72 109 73 110 
<< m1 >>
rect 73 109 74 110 
<< m2 >>
rect 73 109 74 110 
<< m2 >>
rect 74 109 75 110 
<< m1 >>
rect 75 109 76 110 
<< m2 >>
rect 75 109 76 110 
<< m2c >>
rect 75 109 76 110 
<< m1 >>
rect 75 109 76 110 
<< m2 >>
rect 75 109 76 110 
<< m2 >>
rect 76 109 77 110 
<< m1 >>
rect 77 109 78 110 
<< m2 >>
rect 77 109 78 110 
<< m2 >>
rect 78 109 79 110 
<< m1 >>
rect 79 109 80 110 
<< m2 >>
rect 79 109 80 110 
<< m2 >>
rect 80 109 81 110 
<< m1 >>
rect 81 109 82 110 
<< m2 >>
rect 81 109 82 110 
<< m2 >>
rect 82 109 83 110 
<< m1 >>
rect 83 109 84 110 
<< m2 >>
rect 83 109 84 110 
<< m2c >>
rect 83 109 84 110 
<< m1 >>
rect 83 109 84 110 
<< m2 >>
rect 83 109 84 110 
<< m1 >>
rect 84 109 85 110 
<< m1 >>
rect 93 109 94 110 
<< m1 >>
rect 106 109 107 110 
<< m1 >>
rect 124 109 125 110 
<< m1 >>
rect 151 109 152 110 
<< m1 >>
rect 153 109 154 110 
<< m1 >>
rect 163 109 164 110 
<< m1 >>
rect 167 109 168 110 
<< m1 >>
rect 169 109 170 110 
<< m1 >>
rect 178 109 179 110 
<< m1 >>
rect 10 110 11 111 
<< m2 >>
rect 22 110 23 111 
<< m2 >>
rect 25 110 26 111 
<< m1 >>
rect 28 110 29 111 
<< m1 >>
rect 45 110 46 111 
<< m1 >>
rect 49 110 50 111 
<< m1 >>
rect 50 110 51 111 
<< m1 >>
rect 51 110 52 111 
<< m1 >>
rect 52 110 53 111 
<< m1 >>
rect 53 110 54 111 
<< m1 >>
rect 54 110 55 111 
<< m1 >>
rect 55 110 56 111 
<< m1 >>
rect 56 110 57 111 
<< m2 >>
rect 56 110 57 111 
<< m1 >>
rect 57 110 58 111 
<< m1 >>
rect 58 110 59 111 
<< m2 >>
rect 58 110 59 111 
<< m1 >>
rect 59 110 60 111 
<< m1 >>
rect 60 110 61 111 
<< m1 >>
rect 61 110 62 111 
<< m1 >>
rect 62 110 63 111 
<< m1 >>
rect 64 110 65 111 
<< m2 >>
rect 64 110 65 111 
<< m1 >>
rect 67 110 68 111 
<< m1 >>
rect 68 110 69 111 
<< m1 >>
rect 69 110 70 111 
<< m1 >>
rect 70 110 71 111 
<< m1 >>
rect 71 110 72 111 
<< m1 >>
rect 72 110 73 111 
<< m1 >>
rect 73 110 74 111 
<< m1 >>
rect 77 110 78 111 
<< m1 >>
rect 79 110 80 111 
<< m1 >>
rect 81 110 82 111 
<< m1 >>
rect 84 110 85 111 
<< m1 >>
rect 93 110 94 111 
<< m1 >>
rect 106 110 107 111 
<< m1 >>
rect 124 110 125 111 
<< m1 >>
rect 151 110 152 111 
<< m1 >>
rect 153 110 154 111 
<< m1 >>
rect 163 110 164 111 
<< m1 >>
rect 167 110 168 111 
<< m1 >>
rect 169 110 170 111 
<< m2 >>
rect 169 110 170 111 
<< m2c >>
rect 169 110 170 111 
<< m1 >>
rect 169 110 170 111 
<< m2 >>
rect 169 110 170 111 
<< m1 >>
rect 178 110 179 111 
<< m1 >>
rect 10 111 11 112 
<< m1 >>
rect 22 111 23 112 
<< m2 >>
rect 22 111 23 112 
<< m2c >>
rect 22 111 23 112 
<< m1 >>
rect 22 111 23 112 
<< m2 >>
rect 22 111 23 112 
<< m1 >>
rect 25 111 26 112 
<< m2 >>
rect 25 111 26 112 
<< m2c >>
rect 25 111 26 112 
<< m1 >>
rect 25 111 26 112 
<< m2 >>
rect 25 111 26 112 
<< m1 >>
rect 28 111 29 112 
<< m1 >>
rect 45 111 46 112 
<< m2 >>
rect 56 111 57 112 
<< m2 >>
rect 58 111 59 112 
<< m2 >>
rect 59 111 60 112 
<< m2 >>
rect 60 111 61 112 
<< m2 >>
rect 61 111 62 112 
<< m2 >>
rect 62 111 63 112 
<< m1 >>
rect 64 111 65 112 
<< m2 >>
rect 64 111 65 112 
<< m1 >>
rect 75 111 76 112 
<< m2 >>
rect 75 111 76 112 
<< m2c >>
rect 75 111 76 112 
<< m1 >>
rect 75 111 76 112 
<< m2 >>
rect 75 111 76 112 
<< m2 >>
rect 76 111 77 112 
<< m1 >>
rect 77 111 78 112 
<< m2 >>
rect 77 111 78 112 
<< m2 >>
rect 78 111 79 112 
<< m1 >>
rect 79 111 80 112 
<< m2 >>
rect 79 111 80 112 
<< m2 >>
rect 80 111 81 112 
<< m1 >>
rect 81 111 82 112 
<< m2 >>
rect 81 111 82 112 
<< m2c >>
rect 81 111 82 112 
<< m1 >>
rect 81 111 82 112 
<< m2 >>
rect 81 111 82 112 
<< m1 >>
rect 84 111 85 112 
<< m1 >>
rect 93 111 94 112 
<< m2 >>
rect 93 111 94 112 
<< m2c >>
rect 93 111 94 112 
<< m1 >>
rect 93 111 94 112 
<< m2 >>
rect 93 111 94 112 
<< m1 >>
rect 106 111 107 112 
<< m1 >>
rect 124 111 125 112 
<< m1 >>
rect 151 111 152 112 
<< m1 >>
rect 153 111 154 112 
<< m1 >>
rect 163 111 164 112 
<< m1 >>
rect 167 111 168 112 
<< m2 >>
rect 169 111 170 112 
<< m1 >>
rect 178 111 179 112 
<< m1 >>
rect 10 112 11 113 
<< m1 >>
rect 22 112 23 113 
<< m1 >>
rect 25 112 26 113 
<< m1 >>
rect 28 112 29 113 
<< m1 >>
rect 45 112 46 113 
<< m1 >>
rect 56 112 57 113 
<< m2 >>
rect 56 112 57 113 
<< m2c >>
rect 56 112 57 113 
<< m1 >>
rect 56 112 57 113 
<< m2 >>
rect 56 112 57 113 
<< m1 >>
rect 62 112 63 113 
<< m2 >>
rect 62 112 63 113 
<< m2c >>
rect 62 112 63 113 
<< m1 >>
rect 62 112 63 113 
<< m2 >>
rect 62 112 63 113 
<< m1 >>
rect 64 112 65 113 
<< m2 >>
rect 64 112 65 113 
<< m1 >>
rect 75 112 76 113 
<< m1 >>
rect 77 112 78 113 
<< m1 >>
rect 79 112 80 113 
<< m1 >>
rect 84 112 85 113 
<< m2 >>
rect 93 112 94 113 
<< m1 >>
rect 100 112 101 113 
<< m1 >>
rect 101 112 102 113 
<< m1 >>
rect 102 112 103 113 
<< m1 >>
rect 103 112 104 113 
<< m1 >>
rect 104 112 105 113 
<< m1 >>
rect 105 112 106 113 
<< m1 >>
rect 106 112 107 113 
<< m1 >>
rect 124 112 125 113 
<< m1 >>
rect 151 112 152 113 
<< m1 >>
rect 153 112 154 113 
<< m1 >>
rect 163 112 164 113 
<< m1 >>
rect 167 112 168 113 
<< m1 >>
rect 168 112 169 113 
<< m1 >>
rect 169 112 170 113 
<< m2 >>
rect 169 112 170 113 
<< m1 >>
rect 170 112 171 113 
<< m1 >>
rect 171 112 172 113 
<< m1 >>
rect 172 112 173 113 
<< m1 >>
rect 173 112 174 113 
<< m1 >>
rect 174 112 175 113 
<< m1 >>
rect 175 112 176 113 
<< m1 >>
rect 176 112 177 113 
<< m1 >>
rect 177 112 178 113 
<< m1 >>
rect 178 112 179 113 
<< m1 >>
rect 10 113 11 114 
<< m1 >>
rect 22 113 23 114 
<< m1 >>
rect 25 113 26 114 
<< m1 >>
rect 28 113 29 114 
<< m1 >>
rect 45 113 46 114 
<< m1 >>
rect 56 113 57 114 
<< m1 >>
rect 62 113 63 114 
<< m1 >>
rect 64 113 65 114 
<< m2 >>
rect 64 113 65 114 
<< m1 >>
rect 68 113 69 114 
<< m2 >>
rect 68 113 69 114 
<< m2c >>
rect 68 113 69 114 
<< m1 >>
rect 68 113 69 114 
<< m2 >>
rect 68 113 69 114 
<< m1 >>
rect 69 113 70 114 
<< m1 >>
rect 70 113 71 114 
<< m1 >>
rect 71 113 72 114 
<< m1 >>
rect 72 113 73 114 
<< m1 >>
rect 73 113 74 114 
<< m1 >>
rect 74 113 75 114 
<< m1 >>
rect 75 113 76 114 
<< m1 >>
rect 77 113 78 114 
<< m2 >>
rect 77 113 78 114 
<< m2c >>
rect 77 113 78 114 
<< m1 >>
rect 77 113 78 114 
<< m2 >>
rect 77 113 78 114 
<< m1 >>
rect 79 113 80 114 
<< m2 >>
rect 79 113 80 114 
<< m2c >>
rect 79 113 80 114 
<< m1 >>
rect 79 113 80 114 
<< m2 >>
rect 79 113 80 114 
<< m1 >>
rect 84 113 85 114 
<< m1 >>
rect 85 113 86 114 
<< m1 >>
rect 86 113 87 114 
<< m1 >>
rect 87 113 88 114 
<< m1 >>
rect 88 113 89 114 
<< m1 >>
rect 89 113 90 114 
<< m1 >>
rect 90 113 91 114 
<< m1 >>
rect 91 113 92 114 
<< m1 >>
rect 92 113 93 114 
<< m1 >>
rect 93 113 94 114 
<< m2 >>
rect 93 113 94 114 
<< m1 >>
rect 100 113 101 114 
<< m1 >>
rect 124 113 125 114 
<< m1 >>
rect 151 113 152 114 
<< m1 >>
rect 153 113 154 114 
<< m1 >>
rect 163 113 164 114 
<< m2 >>
rect 169 113 170 114 
<< m1 >>
rect 10 114 11 115 
<< m1 >>
rect 22 114 23 115 
<< m1 >>
rect 25 114 26 115 
<< m1 >>
rect 28 114 29 115 
<< m1 >>
rect 45 114 46 115 
<< m1 >>
rect 56 114 57 115 
<< m1 >>
rect 62 114 63 115 
<< m1 >>
rect 64 114 65 115 
<< m2 >>
rect 64 114 65 115 
<< m2 >>
rect 68 114 69 115 
<< m2 >>
rect 77 114 78 115 
<< m2 >>
rect 79 114 80 115 
<< m1 >>
rect 93 114 94 115 
<< m2 >>
rect 93 114 94 115 
<< m1 >>
rect 100 114 101 115 
<< m1 >>
rect 124 114 125 115 
<< m1 >>
rect 151 114 152 115 
<< m1 >>
rect 153 114 154 115 
<< m1 >>
rect 163 114 164 115 
<< m1 >>
rect 169 114 170 115 
<< m2 >>
rect 169 114 170 115 
<< m2c >>
rect 169 114 170 115 
<< m1 >>
rect 169 114 170 115 
<< m2 >>
rect 169 114 170 115 
<< m1 >>
rect 10 115 11 116 
<< m1 >>
rect 22 115 23 116 
<< m1 >>
rect 25 115 26 116 
<< m1 >>
rect 28 115 29 116 
<< m1 >>
rect 45 115 46 116 
<< m1 >>
rect 56 115 57 116 
<< m1 >>
rect 62 115 63 116 
<< m1 >>
rect 64 115 65 116 
<< m2 >>
rect 64 115 65 116 
<< m2 >>
rect 65 115 66 116 
<< m1 >>
rect 66 115 67 116 
<< m2 >>
rect 66 115 67 116 
<< m2c >>
rect 66 115 67 116 
<< m1 >>
rect 66 115 67 116 
<< m2 >>
rect 66 115 67 116 
<< m1 >>
rect 67 115 68 116 
<< m1 >>
rect 68 115 69 116 
<< m2 >>
rect 68 115 69 116 
<< m1 >>
rect 69 115 70 116 
<< m1 >>
rect 70 115 71 116 
<< m1 >>
rect 71 115 72 116 
<< m1 >>
rect 72 115 73 116 
<< m1 >>
rect 73 115 74 116 
<< m1 >>
rect 74 115 75 116 
<< m1 >>
rect 75 115 76 116 
<< m1 >>
rect 76 115 77 116 
<< m1 >>
rect 77 115 78 116 
<< m2 >>
rect 77 115 78 116 
<< m1 >>
rect 78 115 79 116 
<< m1 >>
rect 79 115 80 116 
<< m2 >>
rect 79 115 80 116 
<< m1 >>
rect 80 115 81 116 
<< m1 >>
rect 81 115 82 116 
<< m1 >>
rect 82 115 83 116 
<< m1 >>
rect 83 115 84 116 
<< m1 >>
rect 84 115 85 116 
<< m1 >>
rect 85 115 86 116 
<< m1 >>
rect 86 115 87 116 
<< m1 >>
rect 87 115 88 116 
<< m1 >>
rect 88 115 89 116 
<< m1 >>
rect 89 115 90 116 
<< m1 >>
rect 90 115 91 116 
<< m1 >>
rect 91 115 92 116 
<< m1 >>
rect 93 115 94 116 
<< m2 >>
rect 93 115 94 116 
<< m1 >>
rect 100 115 101 116 
<< m1 >>
rect 124 115 125 116 
<< m1 >>
rect 151 115 152 116 
<< m1 >>
rect 153 115 154 116 
<< m1 >>
rect 163 115 164 116 
<< m1 >>
rect 169 115 170 116 
<< m1 >>
rect 10 116 11 117 
<< m1 >>
rect 22 116 23 117 
<< m1 >>
rect 25 116 26 117 
<< m1 >>
rect 28 116 29 117 
<< m2 >>
rect 28 116 29 117 
<< m2c >>
rect 28 116 29 117 
<< m1 >>
rect 28 116 29 117 
<< m2 >>
rect 28 116 29 117 
<< m1 >>
rect 45 116 46 117 
<< m1 >>
rect 56 116 57 117 
<< m1 >>
rect 62 116 63 117 
<< m1 >>
rect 64 116 65 117 
<< m2 >>
rect 68 116 69 117 
<< m2 >>
rect 77 116 78 117 
<< m2 >>
rect 79 116 80 117 
<< m1 >>
rect 91 116 92 117 
<< m2 >>
rect 91 116 92 117 
<< m2c >>
rect 91 116 92 117 
<< m1 >>
rect 91 116 92 117 
<< m2 >>
rect 91 116 92 117 
<< m1 >>
rect 93 116 94 117 
<< m2 >>
rect 93 116 94 117 
<< m1 >>
rect 100 116 101 117 
<< m1 >>
rect 124 116 125 117 
<< m1 >>
rect 151 116 152 117 
<< m1 >>
rect 153 116 154 117 
<< m1 >>
rect 163 116 164 117 
<< m1 >>
rect 169 116 170 117 
<< m1 >>
rect 10 117 11 118 
<< m1 >>
rect 22 117 23 118 
<< m1 >>
rect 25 117 26 118 
<< m2 >>
rect 27 117 28 118 
<< m2 >>
rect 28 117 29 118 
<< m1 >>
rect 45 117 46 118 
<< m1 >>
rect 56 117 57 118 
<< m1 >>
rect 62 117 63 118 
<< m1 >>
rect 64 117 65 118 
<< m1 >>
rect 68 117 69 118 
<< m2 >>
rect 68 117 69 118 
<< m2c >>
rect 68 117 69 118 
<< m1 >>
rect 68 117 69 118 
<< m2 >>
rect 68 117 69 118 
<< m1 >>
rect 77 117 78 118 
<< m2 >>
rect 77 117 78 118 
<< m2c >>
rect 77 117 78 118 
<< m1 >>
rect 77 117 78 118 
<< m2 >>
rect 77 117 78 118 
<< m1 >>
rect 79 117 80 118 
<< m2 >>
rect 79 117 80 118 
<< m2c >>
rect 79 117 80 118 
<< m1 >>
rect 79 117 80 118 
<< m2 >>
rect 79 117 80 118 
<< m2 >>
rect 91 117 92 118 
<< m1 >>
rect 93 117 94 118 
<< m2 >>
rect 93 117 94 118 
<< m1 >>
rect 100 117 101 118 
<< m1 >>
rect 124 117 125 118 
<< m1 >>
rect 125 117 126 118 
<< m1 >>
rect 126 117 127 118 
<< m1 >>
rect 127 117 128 118 
<< m1 >>
rect 128 117 129 118 
<< m1 >>
rect 129 117 130 118 
<< m1 >>
rect 130 117 131 118 
<< m1 >>
rect 131 117 132 118 
<< m1 >>
rect 132 117 133 118 
<< m1 >>
rect 133 117 134 118 
<< m1 >>
rect 134 117 135 118 
<< m1 >>
rect 135 117 136 118 
<< m1 >>
rect 136 117 137 118 
<< m1 >>
rect 151 117 152 118 
<< m1 >>
rect 153 117 154 118 
<< m1 >>
rect 163 117 164 118 
<< m1 >>
rect 169 117 170 118 
<< m1 >>
rect 10 118 11 119 
<< m1 >>
rect 11 118 12 119 
<< m1 >>
rect 12 118 13 119 
<< m1 >>
rect 13 118 14 119 
<< m1 >>
rect 22 118 23 119 
<< m1 >>
rect 25 118 26 119 
<< m2 >>
rect 27 118 28 119 
<< m1 >>
rect 28 118 29 119 
<< m1 >>
rect 29 118 30 119 
<< m1 >>
rect 30 118 31 119 
<< m1 >>
rect 31 118 32 119 
<< m1 >>
rect 45 118 46 119 
<< m1 >>
rect 56 118 57 119 
<< m1 >>
rect 62 118 63 119 
<< m1 >>
rect 64 118 65 119 
<< m1 >>
rect 67 118 68 119 
<< m1 >>
rect 68 118 69 119 
<< m1 >>
rect 70 118 71 119 
<< m1 >>
rect 71 118 72 119 
<< m1 >>
rect 72 118 73 119 
<< m1 >>
rect 73 118 74 119 
<< m1 >>
rect 77 118 78 119 
<< m1 >>
rect 79 118 80 119 
<< m1 >>
rect 82 118 83 119 
<< m1 >>
rect 83 118 84 119 
<< m1 >>
rect 84 118 85 119 
<< m1 >>
rect 85 118 86 119 
<< m1 >>
rect 88 118 89 119 
<< m1 >>
rect 89 118 90 119 
<< m1 >>
rect 90 118 91 119 
<< m1 >>
rect 91 118 92 119 
<< m2 >>
rect 91 118 92 119 
<< m1 >>
rect 93 118 94 119 
<< m2 >>
rect 93 118 94 119 
<< m1 >>
rect 100 118 101 119 
<< m1 >>
rect 136 118 137 119 
<< m1 >>
rect 142 118 143 119 
<< m1 >>
rect 143 118 144 119 
<< m1 >>
rect 144 118 145 119 
<< m1 >>
rect 145 118 146 119 
<< m1 >>
rect 151 118 152 119 
<< m1 >>
rect 153 118 154 119 
<< m1 >>
rect 163 118 164 119 
<< m1 >>
rect 169 118 170 119 
<< m1 >>
rect 13 119 14 120 
<< m1 >>
rect 22 119 23 120 
<< m1 >>
rect 25 119 26 120 
<< m2 >>
rect 27 119 28 120 
<< m1 >>
rect 28 119 29 120 
<< m1 >>
rect 31 119 32 120 
<< m1 >>
rect 45 119 46 120 
<< m1 >>
rect 56 119 57 120 
<< m1 >>
rect 62 119 63 120 
<< m1 >>
rect 64 119 65 120 
<< m1 >>
rect 67 119 68 120 
<< m1 >>
rect 70 119 71 120 
<< m1 >>
rect 73 119 74 120 
<< m1 >>
rect 77 119 78 120 
<< m1 >>
rect 79 119 80 120 
<< m1 >>
rect 82 119 83 120 
<< m1 >>
rect 85 119 86 120 
<< m1 >>
rect 88 119 89 120 
<< m1 >>
rect 91 119 92 120 
<< m2 >>
rect 91 119 92 120 
<< m1 >>
rect 93 119 94 120 
<< m2 >>
rect 93 119 94 120 
<< m1 >>
rect 100 119 101 120 
<< m1 >>
rect 136 119 137 120 
<< m1 >>
rect 142 119 143 120 
<< m1 >>
rect 145 119 146 120 
<< m1 >>
rect 151 119 152 120 
<< m1 >>
rect 153 119 154 120 
<< m1 >>
rect 163 119 164 120 
<< m1 >>
rect 169 119 170 120 
<< pdiffusion >>
rect 12 120 13 121 
<< m1 >>
rect 13 120 14 121 
<< pdiffusion >>
rect 13 120 14 121 
<< pdiffusion >>
rect 14 120 15 121 
<< pdiffusion >>
rect 15 120 16 121 
<< pdiffusion >>
rect 16 120 17 121 
<< pdiffusion >>
rect 17 120 18 121 
<< m1 >>
rect 22 120 23 121 
<< m1 >>
rect 25 120 26 121 
<< m2 >>
rect 27 120 28 121 
<< m1 >>
rect 28 120 29 121 
<< pdiffusion >>
rect 30 120 31 121 
<< m1 >>
rect 31 120 32 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< m1 >>
rect 45 120 46 121 
<< pdiffusion >>
rect 48 120 49 121 
<< pdiffusion >>
rect 49 120 50 121 
<< pdiffusion >>
rect 50 120 51 121 
<< pdiffusion >>
rect 51 120 52 121 
<< pdiffusion >>
rect 52 120 53 121 
<< pdiffusion >>
rect 53 120 54 121 
<< m1 >>
rect 56 120 57 121 
<< m1 >>
rect 62 120 63 121 
<< m1 >>
rect 64 120 65 121 
<< pdiffusion >>
rect 66 120 67 121 
<< m1 >>
rect 67 120 68 121 
<< pdiffusion >>
rect 67 120 68 121 
<< pdiffusion >>
rect 68 120 69 121 
<< pdiffusion >>
rect 69 120 70 121 
<< m1 >>
rect 70 120 71 121 
<< pdiffusion >>
rect 70 120 71 121 
<< pdiffusion >>
rect 71 120 72 121 
<< m1 >>
rect 73 120 74 121 
<< m1 >>
rect 77 120 78 121 
<< m1 >>
rect 79 120 80 121 
<< m1 >>
rect 82 120 83 121 
<< pdiffusion >>
rect 84 120 85 121 
<< m1 >>
rect 85 120 86 121 
<< pdiffusion >>
rect 85 120 86 121 
<< pdiffusion >>
rect 86 120 87 121 
<< pdiffusion >>
rect 87 120 88 121 
<< m1 >>
rect 88 120 89 121 
<< pdiffusion >>
rect 88 120 89 121 
<< pdiffusion >>
rect 89 120 90 121 
<< m1 >>
rect 91 120 92 121 
<< m2 >>
rect 91 120 92 121 
<< m1 >>
rect 93 120 94 121 
<< m2 >>
rect 93 120 94 121 
<< m1 >>
rect 100 120 101 121 
<< pdiffusion >>
rect 102 120 103 121 
<< pdiffusion >>
rect 103 120 104 121 
<< pdiffusion >>
rect 104 120 105 121 
<< pdiffusion >>
rect 105 120 106 121 
<< pdiffusion >>
rect 106 120 107 121 
<< pdiffusion >>
rect 107 120 108 121 
<< pdiffusion >>
rect 120 120 121 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< m1 >>
rect 136 120 137 121 
<< pdiffusion >>
rect 138 120 139 121 
<< pdiffusion >>
rect 139 120 140 121 
<< pdiffusion >>
rect 140 120 141 121 
<< pdiffusion >>
rect 141 120 142 121 
<< m1 >>
rect 142 120 143 121 
<< pdiffusion >>
rect 142 120 143 121 
<< pdiffusion >>
rect 143 120 144 121 
<< m1 >>
rect 145 120 146 121 
<< m1 >>
rect 151 120 152 121 
<< m1 >>
rect 153 120 154 121 
<< pdiffusion >>
rect 156 120 157 121 
<< pdiffusion >>
rect 157 120 158 121 
<< pdiffusion >>
rect 158 120 159 121 
<< pdiffusion >>
rect 159 120 160 121 
<< pdiffusion >>
rect 160 120 161 121 
<< pdiffusion >>
rect 161 120 162 121 
<< m1 >>
rect 163 120 164 121 
<< m1 >>
rect 169 120 170 121 
<< pdiffusion >>
rect 174 120 175 121 
<< pdiffusion >>
rect 175 120 176 121 
<< pdiffusion >>
rect 176 120 177 121 
<< pdiffusion >>
rect 177 120 178 121 
<< pdiffusion >>
rect 178 120 179 121 
<< pdiffusion >>
rect 179 120 180 121 
<< pdiffusion >>
rect 12 121 13 122 
<< pdiffusion >>
rect 13 121 14 122 
<< pdiffusion >>
rect 14 121 15 122 
<< pdiffusion >>
rect 15 121 16 122 
<< pdiffusion >>
rect 16 121 17 122 
<< pdiffusion >>
rect 17 121 18 122 
<< m1 >>
rect 22 121 23 122 
<< m1 >>
rect 25 121 26 122 
<< m2 >>
rect 27 121 28 122 
<< m1 >>
rect 28 121 29 122 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< m1 >>
rect 45 121 46 122 
<< pdiffusion >>
rect 48 121 49 122 
<< pdiffusion >>
rect 49 121 50 122 
<< pdiffusion >>
rect 50 121 51 122 
<< pdiffusion >>
rect 51 121 52 122 
<< pdiffusion >>
rect 52 121 53 122 
<< pdiffusion >>
rect 53 121 54 122 
<< m1 >>
rect 56 121 57 122 
<< m1 >>
rect 62 121 63 122 
<< m1 >>
rect 64 121 65 122 
<< pdiffusion >>
rect 66 121 67 122 
<< pdiffusion >>
rect 67 121 68 122 
<< pdiffusion >>
rect 68 121 69 122 
<< pdiffusion >>
rect 69 121 70 122 
<< pdiffusion >>
rect 70 121 71 122 
<< pdiffusion >>
rect 71 121 72 122 
<< m1 >>
rect 73 121 74 122 
<< m1 >>
rect 77 121 78 122 
<< m1 >>
rect 79 121 80 122 
<< m1 >>
rect 82 121 83 122 
<< pdiffusion >>
rect 84 121 85 122 
<< pdiffusion >>
rect 85 121 86 122 
<< pdiffusion >>
rect 86 121 87 122 
<< pdiffusion >>
rect 87 121 88 122 
<< pdiffusion >>
rect 88 121 89 122 
<< pdiffusion >>
rect 89 121 90 122 
<< m1 >>
rect 91 121 92 122 
<< m2 >>
rect 91 121 92 122 
<< m1 >>
rect 93 121 94 122 
<< m2 >>
rect 93 121 94 122 
<< m1 >>
rect 100 121 101 122 
<< pdiffusion >>
rect 102 121 103 122 
<< pdiffusion >>
rect 103 121 104 122 
<< pdiffusion >>
rect 104 121 105 122 
<< pdiffusion >>
rect 105 121 106 122 
<< pdiffusion >>
rect 106 121 107 122 
<< pdiffusion >>
rect 107 121 108 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< m1 >>
rect 136 121 137 122 
<< pdiffusion >>
rect 138 121 139 122 
<< pdiffusion >>
rect 139 121 140 122 
<< pdiffusion >>
rect 140 121 141 122 
<< pdiffusion >>
rect 141 121 142 122 
<< pdiffusion >>
rect 142 121 143 122 
<< pdiffusion >>
rect 143 121 144 122 
<< m1 >>
rect 145 121 146 122 
<< m1 >>
rect 151 121 152 122 
<< m1 >>
rect 153 121 154 122 
<< pdiffusion >>
rect 156 121 157 122 
<< pdiffusion >>
rect 157 121 158 122 
<< pdiffusion >>
rect 158 121 159 122 
<< pdiffusion >>
rect 159 121 160 122 
<< pdiffusion >>
rect 160 121 161 122 
<< pdiffusion >>
rect 161 121 162 122 
<< m1 >>
rect 163 121 164 122 
<< m1 >>
rect 169 121 170 122 
<< pdiffusion >>
rect 174 121 175 122 
<< pdiffusion >>
rect 175 121 176 122 
<< pdiffusion >>
rect 176 121 177 122 
<< pdiffusion >>
rect 177 121 178 122 
<< pdiffusion >>
rect 178 121 179 122 
<< pdiffusion >>
rect 179 121 180 122 
<< pdiffusion >>
rect 12 122 13 123 
<< pdiffusion >>
rect 13 122 14 123 
<< pdiffusion >>
rect 14 122 15 123 
<< pdiffusion >>
rect 15 122 16 123 
<< pdiffusion >>
rect 16 122 17 123 
<< pdiffusion >>
rect 17 122 18 123 
<< m1 >>
rect 22 122 23 123 
<< m1 >>
rect 25 122 26 123 
<< m2 >>
rect 27 122 28 123 
<< m1 >>
rect 28 122 29 123 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< m1 >>
rect 45 122 46 123 
<< pdiffusion >>
rect 48 122 49 123 
<< pdiffusion >>
rect 49 122 50 123 
<< pdiffusion >>
rect 50 122 51 123 
<< pdiffusion >>
rect 51 122 52 123 
<< pdiffusion >>
rect 52 122 53 123 
<< pdiffusion >>
rect 53 122 54 123 
<< m1 >>
rect 56 122 57 123 
<< m1 >>
rect 62 122 63 123 
<< m1 >>
rect 64 122 65 123 
<< pdiffusion >>
rect 66 122 67 123 
<< pdiffusion >>
rect 67 122 68 123 
<< pdiffusion >>
rect 68 122 69 123 
<< pdiffusion >>
rect 69 122 70 123 
<< pdiffusion >>
rect 70 122 71 123 
<< pdiffusion >>
rect 71 122 72 123 
<< m1 >>
rect 73 122 74 123 
<< m1 >>
rect 77 122 78 123 
<< m1 >>
rect 79 122 80 123 
<< m1 >>
rect 82 122 83 123 
<< pdiffusion >>
rect 84 122 85 123 
<< pdiffusion >>
rect 85 122 86 123 
<< pdiffusion >>
rect 86 122 87 123 
<< pdiffusion >>
rect 87 122 88 123 
<< pdiffusion >>
rect 88 122 89 123 
<< pdiffusion >>
rect 89 122 90 123 
<< m1 >>
rect 91 122 92 123 
<< m2 >>
rect 91 122 92 123 
<< m1 >>
rect 93 122 94 123 
<< m2 >>
rect 93 122 94 123 
<< m1 >>
rect 100 122 101 123 
<< pdiffusion >>
rect 102 122 103 123 
<< pdiffusion >>
rect 103 122 104 123 
<< pdiffusion >>
rect 104 122 105 123 
<< pdiffusion >>
rect 105 122 106 123 
<< pdiffusion >>
rect 106 122 107 123 
<< pdiffusion >>
rect 107 122 108 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< m1 >>
rect 136 122 137 123 
<< pdiffusion >>
rect 138 122 139 123 
<< pdiffusion >>
rect 139 122 140 123 
<< pdiffusion >>
rect 140 122 141 123 
<< pdiffusion >>
rect 141 122 142 123 
<< pdiffusion >>
rect 142 122 143 123 
<< pdiffusion >>
rect 143 122 144 123 
<< m1 >>
rect 145 122 146 123 
<< m1 >>
rect 151 122 152 123 
<< m1 >>
rect 153 122 154 123 
<< pdiffusion >>
rect 156 122 157 123 
<< pdiffusion >>
rect 157 122 158 123 
<< pdiffusion >>
rect 158 122 159 123 
<< pdiffusion >>
rect 159 122 160 123 
<< pdiffusion >>
rect 160 122 161 123 
<< pdiffusion >>
rect 161 122 162 123 
<< m1 >>
rect 163 122 164 123 
<< m1 >>
rect 169 122 170 123 
<< pdiffusion >>
rect 174 122 175 123 
<< pdiffusion >>
rect 175 122 176 123 
<< pdiffusion >>
rect 176 122 177 123 
<< pdiffusion >>
rect 177 122 178 123 
<< pdiffusion >>
rect 178 122 179 123 
<< pdiffusion >>
rect 179 122 180 123 
<< pdiffusion >>
rect 12 123 13 124 
<< pdiffusion >>
rect 13 123 14 124 
<< pdiffusion >>
rect 14 123 15 124 
<< pdiffusion >>
rect 15 123 16 124 
<< pdiffusion >>
rect 16 123 17 124 
<< pdiffusion >>
rect 17 123 18 124 
<< m1 >>
rect 22 123 23 124 
<< m1 >>
rect 25 123 26 124 
<< m2 >>
rect 27 123 28 124 
<< m1 >>
rect 28 123 29 124 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< m1 >>
rect 45 123 46 124 
<< pdiffusion >>
rect 48 123 49 124 
<< pdiffusion >>
rect 49 123 50 124 
<< pdiffusion >>
rect 50 123 51 124 
<< pdiffusion >>
rect 51 123 52 124 
<< pdiffusion >>
rect 52 123 53 124 
<< pdiffusion >>
rect 53 123 54 124 
<< m1 >>
rect 56 123 57 124 
<< m1 >>
rect 62 123 63 124 
<< m1 >>
rect 64 123 65 124 
<< pdiffusion >>
rect 66 123 67 124 
<< pdiffusion >>
rect 67 123 68 124 
<< pdiffusion >>
rect 68 123 69 124 
<< pdiffusion >>
rect 69 123 70 124 
<< pdiffusion >>
rect 70 123 71 124 
<< pdiffusion >>
rect 71 123 72 124 
<< m1 >>
rect 73 123 74 124 
<< m1 >>
rect 77 123 78 124 
<< m1 >>
rect 79 123 80 124 
<< m1 >>
rect 82 123 83 124 
<< pdiffusion >>
rect 84 123 85 124 
<< pdiffusion >>
rect 85 123 86 124 
<< pdiffusion >>
rect 86 123 87 124 
<< pdiffusion >>
rect 87 123 88 124 
<< pdiffusion >>
rect 88 123 89 124 
<< pdiffusion >>
rect 89 123 90 124 
<< m1 >>
rect 91 123 92 124 
<< m2 >>
rect 91 123 92 124 
<< m1 >>
rect 93 123 94 124 
<< m2 >>
rect 93 123 94 124 
<< m1 >>
rect 100 123 101 124 
<< pdiffusion >>
rect 102 123 103 124 
<< pdiffusion >>
rect 103 123 104 124 
<< pdiffusion >>
rect 104 123 105 124 
<< pdiffusion >>
rect 105 123 106 124 
<< pdiffusion >>
rect 106 123 107 124 
<< pdiffusion >>
rect 107 123 108 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< m1 >>
rect 136 123 137 124 
<< pdiffusion >>
rect 138 123 139 124 
<< pdiffusion >>
rect 139 123 140 124 
<< pdiffusion >>
rect 140 123 141 124 
<< pdiffusion >>
rect 141 123 142 124 
<< pdiffusion >>
rect 142 123 143 124 
<< pdiffusion >>
rect 143 123 144 124 
<< m1 >>
rect 145 123 146 124 
<< m1 >>
rect 151 123 152 124 
<< m1 >>
rect 153 123 154 124 
<< pdiffusion >>
rect 156 123 157 124 
<< pdiffusion >>
rect 157 123 158 124 
<< pdiffusion >>
rect 158 123 159 124 
<< pdiffusion >>
rect 159 123 160 124 
<< pdiffusion >>
rect 160 123 161 124 
<< pdiffusion >>
rect 161 123 162 124 
<< m1 >>
rect 163 123 164 124 
<< m1 >>
rect 169 123 170 124 
<< pdiffusion >>
rect 174 123 175 124 
<< pdiffusion >>
rect 175 123 176 124 
<< pdiffusion >>
rect 176 123 177 124 
<< pdiffusion >>
rect 177 123 178 124 
<< pdiffusion >>
rect 178 123 179 124 
<< pdiffusion >>
rect 179 123 180 124 
<< pdiffusion >>
rect 12 124 13 125 
<< pdiffusion >>
rect 13 124 14 125 
<< pdiffusion >>
rect 14 124 15 125 
<< pdiffusion >>
rect 15 124 16 125 
<< pdiffusion >>
rect 16 124 17 125 
<< pdiffusion >>
rect 17 124 18 125 
<< m1 >>
rect 22 124 23 125 
<< m1 >>
rect 25 124 26 125 
<< m2 >>
rect 27 124 28 125 
<< m1 >>
rect 28 124 29 125 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< m1 >>
rect 45 124 46 125 
<< pdiffusion >>
rect 48 124 49 125 
<< pdiffusion >>
rect 49 124 50 125 
<< pdiffusion >>
rect 50 124 51 125 
<< pdiffusion >>
rect 51 124 52 125 
<< pdiffusion >>
rect 52 124 53 125 
<< pdiffusion >>
rect 53 124 54 125 
<< m1 >>
rect 56 124 57 125 
<< m1 >>
rect 62 124 63 125 
<< m1 >>
rect 64 124 65 125 
<< pdiffusion >>
rect 66 124 67 125 
<< pdiffusion >>
rect 67 124 68 125 
<< pdiffusion >>
rect 68 124 69 125 
<< pdiffusion >>
rect 69 124 70 125 
<< pdiffusion >>
rect 70 124 71 125 
<< pdiffusion >>
rect 71 124 72 125 
<< m1 >>
rect 73 124 74 125 
<< m1 >>
rect 77 124 78 125 
<< m1 >>
rect 79 124 80 125 
<< m1 >>
rect 82 124 83 125 
<< pdiffusion >>
rect 84 124 85 125 
<< pdiffusion >>
rect 85 124 86 125 
<< pdiffusion >>
rect 86 124 87 125 
<< pdiffusion >>
rect 87 124 88 125 
<< pdiffusion >>
rect 88 124 89 125 
<< pdiffusion >>
rect 89 124 90 125 
<< m1 >>
rect 91 124 92 125 
<< m2 >>
rect 91 124 92 125 
<< m1 >>
rect 93 124 94 125 
<< m2 >>
rect 93 124 94 125 
<< m1 >>
rect 100 124 101 125 
<< pdiffusion >>
rect 102 124 103 125 
<< pdiffusion >>
rect 103 124 104 125 
<< pdiffusion >>
rect 104 124 105 125 
<< pdiffusion >>
rect 105 124 106 125 
<< pdiffusion >>
rect 106 124 107 125 
<< pdiffusion >>
rect 107 124 108 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< m1 >>
rect 136 124 137 125 
<< pdiffusion >>
rect 138 124 139 125 
<< pdiffusion >>
rect 139 124 140 125 
<< pdiffusion >>
rect 140 124 141 125 
<< pdiffusion >>
rect 141 124 142 125 
<< pdiffusion >>
rect 142 124 143 125 
<< pdiffusion >>
rect 143 124 144 125 
<< m1 >>
rect 145 124 146 125 
<< m1 >>
rect 151 124 152 125 
<< m1 >>
rect 153 124 154 125 
<< pdiffusion >>
rect 156 124 157 125 
<< pdiffusion >>
rect 157 124 158 125 
<< pdiffusion >>
rect 158 124 159 125 
<< pdiffusion >>
rect 159 124 160 125 
<< pdiffusion >>
rect 160 124 161 125 
<< pdiffusion >>
rect 161 124 162 125 
<< m1 >>
rect 163 124 164 125 
<< m1 >>
rect 169 124 170 125 
<< pdiffusion >>
rect 174 124 175 125 
<< pdiffusion >>
rect 175 124 176 125 
<< pdiffusion >>
rect 176 124 177 125 
<< pdiffusion >>
rect 177 124 178 125 
<< pdiffusion >>
rect 178 124 179 125 
<< pdiffusion >>
rect 179 124 180 125 
<< pdiffusion >>
rect 12 125 13 126 
<< pdiffusion >>
rect 13 125 14 126 
<< pdiffusion >>
rect 14 125 15 126 
<< pdiffusion >>
rect 15 125 16 126 
<< m1 >>
rect 16 125 17 126 
<< pdiffusion >>
rect 16 125 17 126 
<< pdiffusion >>
rect 17 125 18 126 
<< m1 >>
rect 22 125 23 126 
<< m1 >>
rect 25 125 26 126 
<< m2 >>
rect 27 125 28 126 
<< m1 >>
rect 28 125 29 126 
<< pdiffusion >>
rect 30 125 31 126 
<< m1 >>
rect 31 125 32 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< m1 >>
rect 34 125 35 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< m1 >>
rect 45 125 46 126 
<< pdiffusion >>
rect 48 125 49 126 
<< m1 >>
rect 49 125 50 126 
<< pdiffusion >>
rect 49 125 50 126 
<< pdiffusion >>
rect 50 125 51 126 
<< pdiffusion >>
rect 51 125 52 126 
<< m1 >>
rect 52 125 53 126 
<< pdiffusion >>
rect 52 125 53 126 
<< pdiffusion >>
rect 53 125 54 126 
<< m1 >>
rect 56 125 57 126 
<< m1 >>
rect 62 125 63 126 
<< m1 >>
rect 64 125 65 126 
<< pdiffusion >>
rect 66 125 67 126 
<< m1 >>
rect 67 125 68 126 
<< pdiffusion >>
rect 67 125 68 126 
<< pdiffusion >>
rect 68 125 69 126 
<< pdiffusion >>
rect 69 125 70 126 
<< pdiffusion >>
rect 70 125 71 126 
<< pdiffusion >>
rect 71 125 72 126 
<< m1 >>
rect 73 125 74 126 
<< m1 >>
rect 77 125 78 126 
<< m1 >>
rect 79 125 80 126 
<< m1 >>
rect 82 125 83 126 
<< pdiffusion >>
rect 84 125 85 126 
<< pdiffusion >>
rect 85 125 86 126 
<< pdiffusion >>
rect 86 125 87 126 
<< pdiffusion >>
rect 87 125 88 126 
<< m1 >>
rect 88 125 89 126 
<< pdiffusion >>
rect 88 125 89 126 
<< pdiffusion >>
rect 89 125 90 126 
<< m1 >>
rect 91 125 92 126 
<< m2 >>
rect 91 125 92 126 
<< m1 >>
rect 93 125 94 126 
<< m2 >>
rect 93 125 94 126 
<< m1 >>
rect 100 125 101 126 
<< pdiffusion >>
rect 102 125 103 126 
<< pdiffusion >>
rect 103 125 104 126 
<< pdiffusion >>
rect 104 125 105 126 
<< pdiffusion >>
rect 105 125 106 126 
<< m1 >>
rect 106 125 107 126 
<< pdiffusion >>
rect 106 125 107 126 
<< pdiffusion >>
rect 107 125 108 126 
<< pdiffusion >>
rect 120 125 121 126 
<< m1 >>
rect 121 125 122 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< m1 >>
rect 124 125 125 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< m1 >>
rect 136 125 137 126 
<< pdiffusion >>
rect 138 125 139 126 
<< pdiffusion >>
rect 139 125 140 126 
<< pdiffusion >>
rect 140 125 141 126 
<< pdiffusion >>
rect 141 125 142 126 
<< pdiffusion >>
rect 142 125 143 126 
<< pdiffusion >>
rect 143 125 144 126 
<< m1 >>
rect 145 125 146 126 
<< m1 >>
rect 151 125 152 126 
<< m1 >>
rect 153 125 154 126 
<< pdiffusion >>
rect 156 125 157 126 
<< pdiffusion >>
rect 157 125 158 126 
<< pdiffusion >>
rect 158 125 159 126 
<< pdiffusion >>
rect 159 125 160 126 
<< m1 >>
rect 160 125 161 126 
<< pdiffusion >>
rect 160 125 161 126 
<< pdiffusion >>
rect 161 125 162 126 
<< m1 >>
rect 163 125 164 126 
<< m1 >>
rect 169 125 170 126 
<< pdiffusion >>
rect 174 125 175 126 
<< pdiffusion >>
rect 175 125 176 126 
<< pdiffusion >>
rect 176 125 177 126 
<< pdiffusion >>
rect 177 125 178 126 
<< m1 >>
rect 178 125 179 126 
<< pdiffusion >>
rect 178 125 179 126 
<< pdiffusion >>
rect 179 125 180 126 
<< m1 >>
rect 16 126 17 127 
<< m1 >>
rect 22 126 23 127 
<< m1 >>
rect 25 126 26 127 
<< m2 >>
rect 27 126 28 127 
<< m1 >>
rect 28 126 29 127 
<< m1 >>
rect 31 126 32 127 
<< m1 >>
rect 34 126 35 127 
<< m1 >>
rect 45 126 46 127 
<< m1 >>
rect 49 126 50 127 
<< m1 >>
rect 52 126 53 127 
<< m2 >>
rect 52 126 53 127 
<< m2c >>
rect 52 126 53 127 
<< m1 >>
rect 52 126 53 127 
<< m2 >>
rect 52 126 53 127 
<< m1 >>
rect 56 126 57 127 
<< m2 >>
rect 56 126 57 127 
<< m2c >>
rect 56 126 57 127 
<< m1 >>
rect 56 126 57 127 
<< m2 >>
rect 56 126 57 127 
<< m1 >>
rect 62 126 63 127 
<< m2 >>
rect 62 126 63 127 
<< m2c >>
rect 62 126 63 127 
<< m1 >>
rect 62 126 63 127 
<< m2 >>
rect 62 126 63 127 
<< m2 >>
rect 63 126 64 127 
<< m1 >>
rect 64 126 65 127 
<< m2 >>
rect 64 126 65 127 
<< m1 >>
rect 67 126 68 127 
<< m1 >>
rect 73 126 74 127 
<< m1 >>
rect 77 126 78 127 
<< m1 >>
rect 79 126 80 127 
<< m1 >>
rect 82 126 83 127 
<< m1 >>
rect 88 126 89 127 
<< m1 >>
rect 91 126 92 127 
<< m2 >>
rect 91 126 92 127 
<< m1 >>
rect 93 126 94 127 
<< m2 >>
rect 93 126 94 127 
<< m1 >>
rect 100 126 101 127 
<< m1 >>
rect 106 126 107 127 
<< m1 >>
rect 121 126 122 127 
<< m1 >>
rect 124 126 125 127 
<< m1 >>
rect 136 126 137 127 
<< m1 >>
rect 145 126 146 127 
<< m1 >>
rect 151 126 152 127 
<< m1 >>
rect 153 126 154 127 
<< m1 >>
rect 160 126 161 127 
<< m1 >>
rect 163 126 164 127 
<< m1 >>
rect 169 126 170 127 
<< m1 >>
rect 178 126 179 127 
<< m1 >>
rect 16 127 17 128 
<< m1 >>
rect 22 127 23 128 
<< m1 >>
rect 25 127 26 128 
<< m2 >>
rect 27 127 28 128 
<< m1 >>
rect 28 127 29 128 
<< m1 >>
rect 31 127 32 128 
<< m1 >>
rect 34 127 35 128 
<< m1 >>
rect 45 127 46 128 
<< m1 >>
rect 49 127 50 128 
<< m2 >>
rect 52 127 53 128 
<< m2 >>
rect 53 127 54 128 
<< m2 >>
rect 54 127 55 128 
<< m2 >>
rect 55 127 56 128 
<< m2 >>
rect 56 127 57 128 
<< m1 >>
rect 64 127 65 128 
<< m2 >>
rect 64 127 65 128 
<< m2 >>
rect 65 127 66 128 
<< m1 >>
rect 66 127 67 128 
<< m2 >>
rect 66 127 67 128 
<< m2c >>
rect 66 127 67 128 
<< m1 >>
rect 66 127 67 128 
<< m2 >>
rect 66 127 67 128 
<< m1 >>
rect 67 127 68 128 
<< m1 >>
rect 73 127 74 128 
<< m1 >>
rect 77 127 78 128 
<< m1 >>
rect 79 127 80 128 
<< m1 >>
rect 82 127 83 128 
<< m1 >>
rect 88 127 89 128 
<< m1 >>
rect 89 127 90 128 
<< m2 >>
rect 89 127 90 128 
<< m2c >>
rect 89 127 90 128 
<< m1 >>
rect 89 127 90 128 
<< m2 >>
rect 89 127 90 128 
<< m2 >>
rect 90 127 91 128 
<< m1 >>
rect 91 127 92 128 
<< m2 >>
rect 91 127 92 128 
<< m1 >>
rect 93 127 94 128 
<< m2 >>
rect 93 127 94 128 
<< m1 >>
rect 100 127 101 128 
<< m1 >>
rect 106 127 107 128 
<< m1 >>
rect 107 127 108 128 
<< m1 >>
rect 108 127 109 128 
<< m1 >>
rect 109 127 110 128 
<< m1 >>
rect 110 127 111 128 
<< m1 >>
rect 111 127 112 128 
<< m1 >>
rect 112 127 113 128 
<< m1 >>
rect 113 127 114 128 
<< m1 >>
rect 114 127 115 128 
<< m1 >>
rect 115 127 116 128 
<< m1 >>
rect 116 127 117 128 
<< m1 >>
rect 117 127 118 128 
<< m1 >>
rect 118 127 119 128 
<< m1 >>
rect 119 127 120 128 
<< m1 >>
rect 120 127 121 128 
<< m1 >>
rect 121 127 122 128 
<< m1 >>
rect 124 127 125 128 
<< m1 >>
rect 136 127 137 128 
<< m1 >>
rect 145 127 146 128 
<< m1 >>
rect 151 127 152 128 
<< m1 >>
rect 153 127 154 128 
<< m1 >>
rect 160 127 161 128 
<< m1 >>
rect 163 127 164 128 
<< m1 >>
rect 169 127 170 128 
<< m1 >>
rect 178 127 179 128 
<< m1 >>
rect 16 128 17 129 
<< m1 >>
rect 22 128 23 129 
<< m1 >>
rect 25 128 26 129 
<< m2 >>
rect 27 128 28 129 
<< m1 >>
rect 28 128 29 129 
<< m1 >>
rect 31 128 32 129 
<< m1 >>
rect 34 128 35 129 
<< m1 >>
rect 45 128 46 129 
<< m1 >>
rect 49 128 50 129 
<< m1 >>
rect 50 128 51 129 
<< m1 >>
rect 51 128 52 129 
<< m1 >>
rect 52 128 53 129 
<< m1 >>
rect 53 128 54 129 
<< m1 >>
rect 54 128 55 129 
<< m1 >>
rect 55 128 56 129 
<< m1 >>
rect 56 128 57 129 
<< m1 >>
rect 57 128 58 129 
<< m1 >>
rect 58 128 59 129 
<< m1 >>
rect 59 128 60 129 
<< m1 >>
rect 60 128 61 129 
<< m1 >>
rect 61 128 62 129 
<< m1 >>
rect 62 128 63 129 
<< m1 >>
rect 63 128 64 129 
<< m1 >>
rect 64 128 65 129 
<< m1 >>
rect 73 128 74 129 
<< m2 >>
rect 73 128 74 129 
<< m2c >>
rect 73 128 74 129 
<< m1 >>
rect 73 128 74 129 
<< m2 >>
rect 73 128 74 129 
<< m1 >>
rect 77 128 78 129 
<< m2 >>
rect 77 128 78 129 
<< m2c >>
rect 77 128 78 129 
<< m1 >>
rect 77 128 78 129 
<< m2 >>
rect 77 128 78 129 
<< m1 >>
rect 79 128 80 129 
<< m2 >>
rect 79 128 80 129 
<< m2c >>
rect 79 128 80 129 
<< m1 >>
rect 79 128 80 129 
<< m2 >>
rect 79 128 80 129 
<< m1 >>
rect 82 128 83 129 
<< m2 >>
rect 82 128 83 129 
<< m2c >>
rect 82 128 83 129 
<< m1 >>
rect 82 128 83 129 
<< m2 >>
rect 82 128 83 129 
<< m1 >>
rect 91 128 92 129 
<< m1 >>
rect 93 128 94 129 
<< m2 >>
rect 93 128 94 129 
<< m1 >>
rect 100 128 101 129 
<< m1 >>
rect 124 128 125 129 
<< m1 >>
rect 136 128 137 129 
<< m1 >>
rect 137 128 138 129 
<< m1 >>
rect 138 128 139 129 
<< m2 >>
rect 138 128 139 129 
<< m2c >>
rect 138 128 139 129 
<< m1 >>
rect 138 128 139 129 
<< m2 >>
rect 138 128 139 129 
<< m1 >>
rect 145 128 146 129 
<< m2 >>
rect 145 128 146 129 
<< m2c >>
rect 145 128 146 129 
<< m1 >>
rect 145 128 146 129 
<< m2 >>
rect 145 128 146 129 
<< m1 >>
rect 151 128 152 129 
<< m2 >>
rect 151 128 152 129 
<< m2c >>
rect 151 128 152 129 
<< m1 >>
rect 151 128 152 129 
<< m2 >>
rect 151 128 152 129 
<< m1 >>
rect 153 128 154 129 
<< m2 >>
rect 153 128 154 129 
<< m2c >>
rect 153 128 154 129 
<< m1 >>
rect 153 128 154 129 
<< m2 >>
rect 153 128 154 129 
<< m1 >>
rect 160 128 161 129 
<< m1 >>
rect 163 128 164 129 
<< m1 >>
rect 169 128 170 129 
<< m1 >>
rect 178 128 179 129 
<< m1 >>
rect 16 129 17 130 
<< m1 >>
rect 22 129 23 130 
<< m1 >>
rect 25 129 26 130 
<< m2 >>
rect 27 129 28 130 
<< m1 >>
rect 28 129 29 130 
<< m1 >>
rect 31 129 32 130 
<< m1 >>
rect 34 129 35 130 
<< m1 >>
rect 45 129 46 130 
<< m2 >>
rect 73 129 74 130 
<< m2 >>
rect 77 129 78 130 
<< m2 >>
rect 79 129 80 130 
<< m2 >>
rect 82 129 83 130 
<< m2 >>
rect 86 129 87 130 
<< m2 >>
rect 87 129 88 130 
<< m2 >>
rect 88 129 89 130 
<< m2 >>
rect 89 129 90 130 
<< m2 >>
rect 90 129 91 130 
<< m1 >>
rect 91 129 92 130 
<< m2 >>
rect 91 129 92 130 
<< m2 >>
rect 92 129 93 130 
<< m1 >>
rect 93 129 94 130 
<< m2 >>
rect 93 129 94 130 
<< m1 >>
rect 100 129 101 130 
<< m1 >>
rect 124 129 125 130 
<< m2 >>
rect 138 129 139 130 
<< m2 >>
rect 145 129 146 130 
<< m2 >>
rect 146 129 147 130 
<< m2 >>
rect 147 129 148 130 
<< m2 >>
rect 151 129 152 130 
<< m2 >>
rect 153 129 154 130 
<< m2 >>
rect 158 129 159 130 
<< m1 >>
rect 159 129 160 130 
<< m2 >>
rect 159 129 160 130 
<< m2c >>
rect 159 129 160 130 
<< m1 >>
rect 159 129 160 130 
<< m2 >>
rect 159 129 160 130 
<< m1 >>
rect 160 129 161 130 
<< m1 >>
rect 163 129 164 130 
<< m1 >>
rect 169 129 170 130 
<< m1 >>
rect 178 129 179 130 
<< m1 >>
rect 16 130 17 131 
<< m1 >>
rect 22 130 23 131 
<< m1 >>
rect 25 130 26 131 
<< m2 >>
rect 27 130 28 131 
<< m1 >>
rect 28 130 29 131 
<< m1 >>
rect 31 130 32 131 
<< m1 >>
rect 34 130 35 131 
<< m1 >>
rect 45 130 46 131 
<< m2 >>
rect 45 130 46 131 
<< m2c >>
rect 45 130 46 131 
<< m1 >>
rect 45 130 46 131 
<< m2 >>
rect 45 130 46 131 
<< m1 >>
rect 64 130 65 131 
<< m1 >>
rect 65 130 66 131 
<< m1 >>
rect 66 130 67 131 
<< m1 >>
rect 67 130 68 131 
<< m1 >>
rect 68 130 69 131 
<< m1 >>
rect 69 130 70 131 
<< m1 >>
rect 70 130 71 131 
<< m1 >>
rect 71 130 72 131 
<< m1 >>
rect 72 130 73 131 
<< m1 >>
rect 73 130 74 131 
<< m2 >>
rect 73 130 74 131 
<< m1 >>
rect 74 130 75 131 
<< m1 >>
rect 75 130 76 131 
<< m1 >>
rect 76 130 77 131 
<< m1 >>
rect 77 130 78 131 
<< m2 >>
rect 77 130 78 131 
<< m1 >>
rect 78 130 79 131 
<< m1 >>
rect 79 130 80 131 
<< m2 >>
rect 79 130 80 131 
<< m1 >>
rect 80 130 81 131 
<< m1 >>
rect 81 130 82 131 
<< m1 >>
rect 82 130 83 131 
<< m2 >>
rect 82 130 83 131 
<< m1 >>
rect 83 130 84 131 
<< m1 >>
rect 84 130 85 131 
<< m1 >>
rect 85 130 86 131 
<< m1 >>
rect 86 130 87 131 
<< m2 >>
rect 86 130 87 131 
<< m1 >>
rect 87 130 88 131 
<< m1 >>
rect 88 130 89 131 
<< m1 >>
rect 89 130 90 131 
<< m1 >>
rect 90 130 91 131 
<< m1 >>
rect 91 130 92 131 
<< m1 >>
rect 93 130 94 131 
<< m1 >>
rect 100 130 101 131 
<< m1 >>
rect 124 130 125 131 
<< m1 >>
rect 125 130 126 131 
<< m1 >>
rect 126 130 127 131 
<< m1 >>
rect 127 130 128 131 
<< m1 >>
rect 128 130 129 131 
<< m1 >>
rect 129 130 130 131 
<< m1 >>
rect 130 130 131 131 
<< m1 >>
rect 131 130 132 131 
<< m1 >>
rect 132 130 133 131 
<< m1 >>
rect 133 130 134 131 
<< m1 >>
rect 134 130 135 131 
<< m1 >>
rect 135 130 136 131 
<< m1 >>
rect 136 130 137 131 
<< m1 >>
rect 137 130 138 131 
<< m1 >>
rect 138 130 139 131 
<< m2 >>
rect 138 130 139 131 
<< m1 >>
rect 139 130 140 131 
<< m1 >>
rect 140 130 141 131 
<< m1 >>
rect 141 130 142 131 
<< m1 >>
rect 142 130 143 131 
<< m1 >>
rect 143 130 144 131 
<< m1 >>
rect 144 130 145 131 
<< m1 >>
rect 145 130 146 131 
<< m1 >>
rect 146 130 147 131 
<< m1 >>
rect 147 130 148 131 
<< m2 >>
rect 147 130 148 131 
<< m1 >>
rect 148 130 149 131 
<< m1 >>
rect 149 130 150 131 
<< m1 >>
rect 150 130 151 131 
<< m1 >>
rect 151 130 152 131 
<< m2 >>
rect 151 130 152 131 
<< m1 >>
rect 152 130 153 131 
<< m1 >>
rect 153 130 154 131 
<< m2 >>
rect 153 130 154 131 
<< m1 >>
rect 154 130 155 131 
<< m1 >>
rect 155 130 156 131 
<< m1 >>
rect 156 130 157 131 
<< m1 >>
rect 157 130 158 131 
<< m2 >>
rect 158 130 159 131 
<< m1 >>
rect 163 130 164 131 
<< m1 >>
rect 169 130 170 131 
<< m1 >>
rect 170 130 171 131 
<< m1 >>
rect 171 130 172 131 
<< m1 >>
rect 172 130 173 131 
<< m1 >>
rect 173 130 174 131 
<< m1 >>
rect 174 130 175 131 
<< m1 >>
rect 175 130 176 131 
<< m1 >>
rect 176 130 177 131 
<< m1 >>
rect 177 130 178 131 
<< m1 >>
rect 178 130 179 131 
<< m1 >>
rect 10 131 11 132 
<< m1 >>
rect 11 131 12 132 
<< m1 >>
rect 12 131 13 132 
<< m1 >>
rect 13 131 14 132 
<< m1 >>
rect 14 131 15 132 
<< m1 >>
rect 15 131 16 132 
<< m1 >>
rect 16 131 17 132 
<< m1 >>
rect 22 131 23 132 
<< m2 >>
rect 22 131 23 132 
<< m2c >>
rect 22 131 23 132 
<< m1 >>
rect 22 131 23 132 
<< m2 >>
rect 22 131 23 132 
<< m1 >>
rect 25 131 26 132 
<< m2 >>
rect 25 131 26 132 
<< m2c >>
rect 25 131 26 132 
<< m1 >>
rect 25 131 26 132 
<< m2 >>
rect 25 131 26 132 
<< m2 >>
rect 27 131 28 132 
<< m1 >>
rect 28 131 29 132 
<< m1 >>
rect 29 131 30 132 
<< m2 >>
rect 29 131 30 132 
<< m2c >>
rect 29 131 30 132 
<< m1 >>
rect 29 131 30 132 
<< m2 >>
rect 29 131 30 132 
<< m2 >>
rect 30 131 31 132 
<< m1 >>
rect 31 131 32 132 
<< m2 >>
rect 31 131 32 132 
<< m2 >>
rect 32 131 33 132 
<< m1 >>
rect 34 131 35 132 
<< m2 >>
rect 45 131 46 132 
<< m1 >>
rect 64 131 65 132 
<< m2 >>
rect 73 131 74 132 
<< m2 >>
rect 77 131 78 132 
<< m2 >>
rect 79 131 80 132 
<< m2 >>
rect 82 131 83 132 
<< m2 >>
rect 86 131 87 132 
<< m2 >>
rect 88 131 89 132 
<< m2 >>
rect 89 131 90 132 
<< m2 >>
rect 90 131 91 132 
<< m2 >>
rect 91 131 92 132 
<< m2 >>
rect 92 131 93 132 
<< m1 >>
rect 93 131 94 132 
<< m2 >>
rect 93 131 94 132 
<< m2c >>
rect 93 131 94 132 
<< m1 >>
rect 93 131 94 132 
<< m2 >>
rect 93 131 94 132 
<< m1 >>
rect 100 131 101 132 
<< m2 >>
rect 100 131 101 132 
<< m2c >>
rect 100 131 101 132 
<< m1 >>
rect 100 131 101 132 
<< m2 >>
rect 100 131 101 132 
<< m2 >>
rect 138 131 139 132 
<< m2 >>
rect 139 131 140 132 
<< m2 >>
rect 140 131 141 132 
<< m2 >>
rect 141 131 142 132 
<< m2 >>
rect 142 131 143 132 
<< m2 >>
rect 143 131 144 132 
<< m2 >>
rect 144 131 145 132 
<< m2 >>
rect 145 131 146 132 
<< m2 >>
rect 147 131 148 132 
<< m2 >>
rect 151 131 152 132 
<< m2 >>
rect 153 131 154 132 
<< m1 >>
rect 157 131 158 132 
<< m2 >>
rect 158 131 159 132 
<< m1 >>
rect 163 131 164 132 
<< m1 >>
rect 10 132 11 133 
<< m2 >>
rect 22 132 23 133 
<< m2 >>
rect 25 132 26 133 
<< m2 >>
rect 27 132 28 133 
<< m1 >>
rect 31 132 32 133 
<< m2 >>
rect 32 132 33 133 
<< m1 >>
rect 34 132 35 133 
<< m1 >>
rect 35 132 36 133 
<< m1 >>
rect 36 132 37 133 
<< m1 >>
rect 37 132 38 133 
<< m1 >>
rect 38 132 39 133 
<< m1 >>
rect 39 132 40 133 
<< m1 >>
rect 40 132 41 133 
<< m1 >>
rect 41 132 42 133 
<< m1 >>
rect 42 132 43 133 
<< m1 >>
rect 43 132 44 133 
<< m1 >>
rect 44 132 45 133 
<< m1 >>
rect 45 132 46 133 
<< m2 >>
rect 45 132 46 133 
<< m1 >>
rect 64 132 65 133 
<< m1 >>
rect 73 132 74 133 
<< m2 >>
rect 73 132 74 133 
<< m2c >>
rect 73 132 74 133 
<< m1 >>
rect 73 132 74 133 
<< m2 >>
rect 73 132 74 133 
<< m1 >>
rect 77 132 78 133 
<< m2 >>
rect 77 132 78 133 
<< m2c >>
rect 77 132 78 133 
<< m1 >>
rect 77 132 78 133 
<< m2 >>
rect 77 132 78 133 
<< m1 >>
rect 79 132 80 133 
<< m2 >>
rect 79 132 80 133 
<< m2c >>
rect 79 132 80 133 
<< m1 >>
rect 79 132 80 133 
<< m2 >>
rect 79 132 80 133 
<< m1 >>
rect 82 132 83 133 
<< m2 >>
rect 82 132 83 133 
<< m2c >>
rect 82 132 83 133 
<< m1 >>
rect 82 132 83 133 
<< m2 >>
rect 82 132 83 133 
<< m2 >>
rect 86 132 87 133 
<< m2 >>
rect 88 132 89 133 
<< m2 >>
rect 100 132 101 133 
<< m1 >>
rect 145 132 146 133 
<< m2 >>
rect 145 132 146 133 
<< m2c >>
rect 145 132 146 133 
<< m1 >>
rect 145 132 146 133 
<< m2 >>
rect 145 132 146 133 
<< m1 >>
rect 147 132 148 133 
<< m2 >>
rect 147 132 148 133 
<< m2c >>
rect 147 132 148 133 
<< m1 >>
rect 147 132 148 133 
<< m2 >>
rect 147 132 148 133 
<< m1 >>
rect 151 132 152 133 
<< m2 >>
rect 151 132 152 133 
<< m2c >>
rect 151 132 152 133 
<< m1 >>
rect 151 132 152 133 
<< m2 >>
rect 151 132 152 133 
<< m1 >>
rect 153 132 154 133 
<< m2 >>
rect 153 132 154 133 
<< m2c >>
rect 153 132 154 133 
<< m1 >>
rect 153 132 154 133 
<< m2 >>
rect 153 132 154 133 
<< m1 >>
rect 155 132 156 133 
<< m2 >>
rect 155 132 156 133 
<< m2c >>
rect 155 132 156 133 
<< m1 >>
rect 155 132 156 133 
<< m2 >>
rect 155 132 156 133 
<< m2 >>
rect 156 132 157 133 
<< m1 >>
rect 157 132 158 133 
<< m2 >>
rect 157 132 158 133 
<< m2 >>
rect 158 132 159 133 
<< m1 >>
rect 163 132 164 133 
<< m1 >>
rect 10 133 11 134 
<< m1 >>
rect 16 133 17 134 
<< m1 >>
rect 17 133 18 134 
<< m1 >>
rect 18 133 19 134 
<< m1 >>
rect 19 133 20 134 
<< m1 >>
rect 20 133 21 134 
<< m1 >>
rect 21 133 22 134 
<< m1 >>
rect 22 133 23 134 
<< m2 >>
rect 22 133 23 134 
<< m1 >>
rect 23 133 24 134 
<< m1 >>
rect 24 133 25 134 
<< m1 >>
rect 25 133 26 134 
<< m2 >>
rect 25 133 26 134 
<< m1 >>
rect 26 133 27 134 
<< m1 >>
rect 27 133 28 134 
<< m2 >>
rect 27 133 28 134 
<< m1 >>
rect 28 133 29 134 
<< m1 >>
rect 29 133 30 134 
<< m1 >>
rect 30 133 31 134 
<< m1 >>
rect 31 133 32 134 
<< m2 >>
rect 32 133 33 134 
<< m1 >>
rect 45 133 46 134 
<< m2 >>
rect 45 133 46 134 
<< m1 >>
rect 48 133 49 134 
<< m1 >>
rect 49 133 50 134 
<< m1 >>
rect 50 133 51 134 
<< m1 >>
rect 51 133 52 134 
<< m1 >>
rect 52 133 53 134 
<< m1 >>
rect 64 133 65 134 
<< m2 >>
rect 64 133 65 134 
<< m2 >>
rect 65 133 66 134 
<< m1 >>
rect 66 133 67 134 
<< m2 >>
rect 66 133 67 134 
<< m2c >>
rect 66 133 67 134 
<< m1 >>
rect 66 133 67 134 
<< m2 >>
rect 66 133 67 134 
<< m1 >>
rect 67 133 68 134 
<< m1 >>
rect 68 133 69 134 
<< m1 >>
rect 69 133 70 134 
<< m1 >>
rect 70 133 71 134 
<< m1 >>
rect 71 133 72 134 
<< m1 >>
rect 73 133 74 134 
<< m2 >>
rect 77 133 78 134 
<< m2 >>
rect 79 133 80 134 
<< m1 >>
rect 82 133 83 134 
<< m1 >>
rect 84 133 85 134 
<< m2 >>
rect 84 133 85 134 
<< m1 >>
rect 85 133 86 134 
<< m2 >>
rect 85 133 86 134 
<< m1 >>
rect 86 133 87 134 
<< m2 >>
rect 86 133 87 134 
<< m1 >>
rect 87 133 88 134 
<< m1 >>
rect 88 133 89 134 
<< m2 >>
rect 88 133 89 134 
<< m1 >>
rect 89 133 90 134 
<< m1 >>
rect 90 133 91 134 
<< m1 >>
rect 91 133 92 134 
<< m1 >>
rect 92 133 93 134 
<< m1 >>
rect 93 133 94 134 
<< m1 >>
rect 94 133 95 134 
<< m1 >>
rect 95 133 96 134 
<< m1 >>
rect 96 133 97 134 
<< m1 >>
rect 97 133 98 134 
<< m1 >>
rect 98 133 99 134 
<< m1 >>
rect 99 133 100 134 
<< m1 >>
rect 100 133 101 134 
<< m2 >>
rect 100 133 101 134 
<< m1 >>
rect 101 133 102 134 
<< m1 >>
rect 102 133 103 134 
<< m1 >>
rect 103 133 104 134 
<< m1 >>
rect 104 133 105 134 
<< m1 >>
rect 105 133 106 134 
<< m1 >>
rect 106 133 107 134 
<< m1 >>
rect 107 133 108 134 
<< m1 >>
rect 108 133 109 134 
<< m1 >>
rect 109 133 110 134 
<< m1 >>
rect 110 133 111 134 
<< m1 >>
rect 111 133 112 134 
<< m1 >>
rect 112 133 113 134 
<< m1 >>
rect 113 133 114 134 
<< m1 >>
rect 114 133 115 134 
<< m1 >>
rect 115 133 116 134 
<< m1 >>
rect 116 133 117 134 
<< m1 >>
rect 117 133 118 134 
<< m1 >>
rect 118 133 119 134 
<< m1 >>
rect 119 133 120 134 
<< m1 >>
rect 120 133 121 134 
<< m1 >>
rect 121 133 122 134 
<< m1 >>
rect 122 133 123 134 
<< m1 >>
rect 123 133 124 134 
<< m1 >>
rect 124 133 125 134 
<< m1 >>
rect 145 133 146 134 
<< m1 >>
rect 147 133 148 134 
<< m2 >>
rect 151 133 152 134 
<< m2 >>
rect 153 133 154 134 
<< m1 >>
rect 155 133 156 134 
<< m1 >>
rect 157 133 158 134 
<< m1 >>
rect 163 133 164 134 
<< m1 >>
rect 10 134 11 135 
<< m1 >>
rect 16 134 17 135 
<< m2 >>
rect 22 134 23 135 
<< m2 >>
rect 25 134 26 135 
<< m2 >>
rect 27 134 28 135 
<< m2 >>
rect 32 134 33 135 
<< m1 >>
rect 33 134 34 135 
<< m2 >>
rect 33 134 34 135 
<< m2c >>
rect 33 134 34 135 
<< m1 >>
rect 33 134 34 135 
<< m2 >>
rect 33 134 34 135 
<< m1 >>
rect 34 134 35 135 
<< m1 >>
rect 43 134 44 135 
<< m2 >>
rect 43 134 44 135 
<< m2c >>
rect 43 134 44 135 
<< m1 >>
rect 43 134 44 135 
<< m2 >>
rect 43 134 44 135 
<< m2 >>
rect 44 134 45 135 
<< m1 >>
rect 45 134 46 135 
<< m2 >>
rect 45 134 46 135 
<< m1 >>
rect 48 134 49 135 
<< m1 >>
rect 52 134 53 135 
<< m1 >>
rect 64 134 65 135 
<< m2 >>
rect 64 134 65 135 
<< m1 >>
rect 71 134 72 135 
<< m2 >>
rect 71 134 72 135 
<< m2c >>
rect 71 134 72 135 
<< m1 >>
rect 71 134 72 135 
<< m2 >>
rect 71 134 72 135 
<< m2 >>
rect 72 134 73 135 
<< m1 >>
rect 73 134 74 135 
<< m2 >>
rect 73 134 74 135 
<< m2 >>
rect 74 134 75 135 
<< m1 >>
rect 75 134 76 135 
<< m2 >>
rect 75 134 76 135 
<< m2c >>
rect 75 134 76 135 
<< m1 >>
rect 75 134 76 135 
<< m2 >>
rect 75 134 76 135 
<< m1 >>
rect 76 134 77 135 
<< m1 >>
rect 77 134 78 135 
<< m2 >>
rect 77 134 78 135 
<< m1 >>
rect 78 134 79 135 
<< m1 >>
rect 79 134 80 135 
<< m2 >>
rect 79 134 80 135 
<< m1 >>
rect 80 134 81 135 
<< m1 >>
rect 81 134 82 135 
<< m1 >>
rect 82 134 83 135 
<< m1 >>
rect 84 134 85 135 
<< m2 >>
rect 84 134 85 135 
<< m2 >>
rect 88 134 89 135 
<< m2 >>
rect 100 134 101 135 
<< m1 >>
rect 124 134 125 135 
<< m1 >>
rect 145 134 146 135 
<< m2 >>
rect 145 134 146 135 
<< m2 >>
rect 146 134 147 135 
<< m1 >>
rect 147 134 148 135 
<< m2 >>
rect 147 134 148 135 
<< m2 >>
rect 148 134 149 135 
<< m1 >>
rect 149 134 150 135 
<< m2 >>
rect 149 134 150 135 
<< m2c >>
rect 149 134 150 135 
<< m1 >>
rect 149 134 150 135 
<< m2 >>
rect 149 134 150 135 
<< m1 >>
rect 150 134 151 135 
<< m1 >>
rect 151 134 152 135 
<< m2 >>
rect 151 134 152 135 
<< m1 >>
rect 152 134 153 135 
<< m1 >>
rect 153 134 154 135 
<< m2 >>
rect 153 134 154 135 
<< m1 >>
rect 154 134 155 135 
<< m1 >>
rect 155 134 156 135 
<< m1 >>
rect 157 134 158 135 
<< m1 >>
rect 163 134 164 135 
<< m1 >>
rect 10 135 11 136 
<< m1 >>
rect 16 135 17 136 
<< m1 >>
rect 22 135 23 136 
<< m2 >>
rect 22 135 23 136 
<< m2c >>
rect 22 135 23 136 
<< m1 >>
rect 22 135 23 136 
<< m2 >>
rect 22 135 23 136 
<< m1 >>
rect 25 135 26 136 
<< m2 >>
rect 25 135 26 136 
<< m2c >>
rect 25 135 26 136 
<< m1 >>
rect 25 135 26 136 
<< m2 >>
rect 25 135 26 136 
<< m1 >>
rect 27 135 28 136 
<< m2 >>
rect 27 135 28 136 
<< m2c >>
rect 27 135 28 136 
<< m1 >>
rect 27 135 28 136 
<< m2 >>
rect 27 135 28 136 
<< m1 >>
rect 34 135 35 136 
<< m1 >>
rect 43 135 44 136 
<< m1 >>
rect 45 135 46 136 
<< m1 >>
rect 48 135 49 136 
<< m1 >>
rect 52 135 53 136 
<< m1 >>
rect 64 135 65 136 
<< m2 >>
rect 64 135 65 136 
<< m1 >>
rect 73 135 74 136 
<< m2 >>
rect 77 135 78 136 
<< m2 >>
rect 79 135 80 136 
<< m1 >>
rect 84 135 85 136 
<< m2 >>
rect 84 135 85 136 
<< m1 >>
rect 88 135 89 136 
<< m2 >>
rect 88 135 89 136 
<< m2c >>
rect 88 135 89 136 
<< m1 >>
rect 88 135 89 136 
<< m2 >>
rect 88 135 89 136 
<< m1 >>
rect 100 135 101 136 
<< m2 >>
rect 100 135 101 136 
<< m2c >>
rect 100 135 101 136 
<< m1 >>
rect 100 135 101 136 
<< m2 >>
rect 100 135 101 136 
<< m1 >>
rect 124 135 125 136 
<< m1 >>
rect 145 135 146 136 
<< m2 >>
rect 145 135 146 136 
<< m1 >>
rect 147 135 148 136 
<< m2 >>
rect 151 135 152 136 
<< m2 >>
rect 153 135 154 136 
<< m2 >>
rect 154 135 155 136 
<< m1 >>
rect 157 135 158 136 
<< m1 >>
rect 163 135 164 136 
<< m1 >>
rect 10 136 11 137 
<< m1 >>
rect 16 136 17 137 
<< m1 >>
rect 22 136 23 137 
<< m1 >>
rect 25 136 26 137 
<< m1 >>
rect 27 136 28 137 
<< m1 >>
rect 34 136 35 137 
<< m1 >>
rect 41 136 42 137 
<< m2 >>
rect 41 136 42 137 
<< m2c >>
rect 41 136 42 137 
<< m1 >>
rect 41 136 42 137 
<< m2 >>
rect 41 136 42 137 
<< m2 >>
rect 42 136 43 137 
<< m1 >>
rect 43 136 44 137 
<< m2 >>
rect 43 136 44 137 
<< m2 >>
rect 44 136 45 137 
<< m1 >>
rect 45 136 46 137 
<< m2 >>
rect 45 136 46 137 
<< m2 >>
rect 46 136 47 137 
<< m1 >>
rect 47 136 48 137 
<< m2 >>
rect 47 136 48 137 
<< m2c >>
rect 47 136 48 137 
<< m1 >>
rect 47 136 48 137 
<< m2 >>
rect 47 136 48 137 
<< m1 >>
rect 48 136 49 137 
<< m1 >>
rect 52 136 53 137 
<< m1 >>
rect 64 136 65 137 
<< m2 >>
rect 64 136 65 137 
<< m1 >>
rect 70 136 71 137 
<< m1 >>
rect 71 136 72 137 
<< m2 >>
rect 71 136 72 137 
<< m2c >>
rect 71 136 72 137 
<< m1 >>
rect 71 136 72 137 
<< m2 >>
rect 71 136 72 137 
<< m2 >>
rect 72 136 73 137 
<< m1 >>
rect 73 136 74 137 
<< m2 >>
rect 73 136 74 137 
<< m2 >>
rect 74 136 75 137 
<< m1 >>
rect 75 136 76 137 
<< m2 >>
rect 75 136 76 137 
<< m2c >>
rect 75 136 76 137 
<< m1 >>
rect 75 136 76 137 
<< m2 >>
rect 75 136 76 137 
<< m1 >>
rect 76 136 77 137 
<< m1 >>
rect 77 136 78 137 
<< m2 >>
rect 77 136 78 137 
<< m2c >>
rect 77 136 78 137 
<< m1 >>
rect 77 136 78 137 
<< m2 >>
rect 77 136 78 137 
<< m1 >>
rect 79 136 80 137 
<< m2 >>
rect 79 136 80 137 
<< m2c >>
rect 79 136 80 137 
<< m1 >>
rect 79 136 80 137 
<< m2 >>
rect 79 136 80 137 
<< m1 >>
rect 81 136 82 137 
<< m2 >>
rect 81 136 82 137 
<< m1 >>
rect 82 136 83 137 
<< m2 >>
rect 82 136 83 137 
<< m1 >>
rect 83 136 84 137 
<< m2 >>
rect 83 136 84 137 
<< m1 >>
rect 84 136 85 137 
<< m2 >>
rect 84 136 85 137 
<< m1 >>
rect 88 136 89 137 
<< m1 >>
rect 100 136 101 137 
<< m1 >>
rect 124 136 125 137 
<< m1 >>
rect 145 136 146 137 
<< m2 >>
rect 145 136 146 137 
<< m1 >>
rect 147 136 148 137 
<< m1 >>
rect 151 136 152 137 
<< m2 >>
rect 151 136 152 137 
<< m2c >>
rect 151 136 152 137 
<< m1 >>
rect 151 136 152 137 
<< m2 >>
rect 151 136 152 137 
<< m1 >>
rect 154 136 155 137 
<< m2 >>
rect 154 136 155 137 
<< m2c >>
rect 154 136 155 137 
<< m1 >>
rect 154 136 155 137 
<< m2 >>
rect 154 136 155 137 
<< m1 >>
rect 157 136 158 137 
<< m1 >>
rect 163 136 164 137 
<< m1 >>
rect 10 137 11 138 
<< m1 >>
rect 16 137 17 138 
<< m1 >>
rect 22 137 23 138 
<< m1 >>
rect 25 137 26 138 
<< m1 >>
rect 27 137 28 138 
<< m1 >>
rect 34 137 35 138 
<< m1 >>
rect 41 137 42 138 
<< m1 >>
rect 43 137 44 138 
<< m1 >>
rect 45 137 46 138 
<< m1 >>
rect 52 137 53 138 
<< m1 >>
rect 64 137 65 138 
<< m2 >>
rect 64 137 65 138 
<< m1 >>
rect 70 137 71 138 
<< m1 >>
rect 73 137 74 138 
<< m1 >>
rect 79 137 80 138 
<< m1 >>
rect 81 137 82 138 
<< m2 >>
rect 81 137 82 138 
<< m1 >>
rect 88 137 89 138 
<< m1 >>
rect 100 137 101 138 
<< m1 >>
rect 124 137 125 138 
<< m1 >>
rect 145 137 146 138 
<< m2 >>
rect 145 137 146 138 
<< m1 >>
rect 147 137 148 138 
<< m1 >>
rect 151 137 152 138 
<< m1 >>
rect 154 137 155 138 
<< m1 >>
rect 157 137 158 138 
<< m1 >>
rect 163 137 164 138 
<< m1 >>
rect 10 138 11 139 
<< pdiffusion >>
rect 12 138 13 139 
<< pdiffusion >>
rect 13 138 14 139 
<< pdiffusion >>
rect 14 138 15 139 
<< pdiffusion >>
rect 15 138 16 139 
<< m1 >>
rect 16 138 17 139 
<< pdiffusion >>
rect 16 138 17 139 
<< pdiffusion >>
rect 17 138 18 139 
<< m1 >>
rect 22 138 23 139 
<< m1 >>
rect 25 138 26 139 
<< m1 >>
rect 27 138 28 139 
<< pdiffusion >>
rect 30 138 31 139 
<< pdiffusion >>
rect 31 138 32 139 
<< pdiffusion >>
rect 32 138 33 139 
<< pdiffusion >>
rect 33 138 34 139 
<< m1 >>
rect 34 138 35 139 
<< pdiffusion >>
rect 34 138 35 139 
<< pdiffusion >>
rect 35 138 36 139 
<< m1 >>
rect 41 138 42 139 
<< m1 >>
rect 43 138 44 139 
<< m1 >>
rect 45 138 46 139 
<< pdiffusion >>
rect 48 138 49 139 
<< pdiffusion >>
rect 49 138 50 139 
<< pdiffusion >>
rect 50 138 51 139 
<< pdiffusion >>
rect 51 138 52 139 
<< m1 >>
rect 52 138 53 139 
<< pdiffusion >>
rect 52 138 53 139 
<< pdiffusion >>
rect 53 138 54 139 
<< m1 >>
rect 64 138 65 139 
<< m2 >>
rect 64 138 65 139 
<< pdiffusion >>
rect 66 138 67 139 
<< pdiffusion >>
rect 67 138 68 139 
<< pdiffusion >>
rect 68 138 69 139 
<< pdiffusion >>
rect 69 138 70 139 
<< m1 >>
rect 70 138 71 139 
<< pdiffusion >>
rect 70 138 71 139 
<< pdiffusion >>
rect 71 138 72 139 
<< m1 >>
rect 73 138 74 139 
<< m1 >>
rect 79 138 80 139 
<< m1 >>
rect 81 138 82 139 
<< m2 >>
rect 81 138 82 139 
<< pdiffusion >>
rect 84 138 85 139 
<< pdiffusion >>
rect 85 138 86 139 
<< pdiffusion >>
rect 86 138 87 139 
<< pdiffusion >>
rect 87 138 88 139 
<< m1 >>
rect 88 138 89 139 
<< pdiffusion >>
rect 88 138 89 139 
<< pdiffusion >>
rect 89 138 90 139 
<< m1 >>
rect 100 138 101 139 
<< pdiffusion >>
rect 102 138 103 139 
<< pdiffusion >>
rect 103 138 104 139 
<< pdiffusion >>
rect 104 138 105 139 
<< pdiffusion >>
rect 105 138 106 139 
<< pdiffusion >>
rect 106 138 107 139 
<< pdiffusion >>
rect 107 138 108 139 
<< pdiffusion >>
rect 120 138 121 139 
<< pdiffusion >>
rect 121 138 122 139 
<< pdiffusion >>
rect 122 138 123 139 
<< pdiffusion >>
rect 123 138 124 139 
<< m1 >>
rect 124 138 125 139 
<< pdiffusion >>
rect 124 138 125 139 
<< pdiffusion >>
rect 125 138 126 139 
<< pdiffusion >>
rect 138 138 139 139 
<< pdiffusion >>
rect 139 138 140 139 
<< pdiffusion >>
rect 140 138 141 139 
<< pdiffusion >>
rect 141 138 142 139 
<< pdiffusion >>
rect 142 138 143 139 
<< pdiffusion >>
rect 143 138 144 139 
<< m1 >>
rect 145 138 146 139 
<< m2 >>
rect 145 138 146 139 
<< m1 >>
rect 147 138 148 139 
<< m1 >>
rect 151 138 152 139 
<< m1 >>
rect 154 138 155 139 
<< pdiffusion >>
rect 156 138 157 139 
<< m1 >>
rect 157 138 158 139 
<< pdiffusion >>
rect 157 138 158 139 
<< pdiffusion >>
rect 158 138 159 139 
<< pdiffusion >>
rect 159 138 160 139 
<< pdiffusion >>
rect 160 138 161 139 
<< pdiffusion >>
rect 161 138 162 139 
<< m1 >>
rect 163 138 164 139 
<< m1 >>
rect 10 139 11 140 
<< pdiffusion >>
rect 12 139 13 140 
<< pdiffusion >>
rect 13 139 14 140 
<< pdiffusion >>
rect 14 139 15 140 
<< pdiffusion >>
rect 15 139 16 140 
<< pdiffusion >>
rect 16 139 17 140 
<< pdiffusion >>
rect 17 139 18 140 
<< m1 >>
rect 22 139 23 140 
<< m1 >>
rect 25 139 26 140 
<< m1 >>
rect 27 139 28 140 
<< pdiffusion >>
rect 30 139 31 140 
<< pdiffusion >>
rect 31 139 32 140 
<< pdiffusion >>
rect 32 139 33 140 
<< pdiffusion >>
rect 33 139 34 140 
<< pdiffusion >>
rect 34 139 35 140 
<< pdiffusion >>
rect 35 139 36 140 
<< m1 >>
rect 41 139 42 140 
<< m1 >>
rect 43 139 44 140 
<< m1 >>
rect 45 139 46 140 
<< pdiffusion >>
rect 48 139 49 140 
<< pdiffusion >>
rect 49 139 50 140 
<< pdiffusion >>
rect 50 139 51 140 
<< pdiffusion >>
rect 51 139 52 140 
<< pdiffusion >>
rect 52 139 53 140 
<< pdiffusion >>
rect 53 139 54 140 
<< m1 >>
rect 64 139 65 140 
<< m2 >>
rect 64 139 65 140 
<< pdiffusion >>
rect 66 139 67 140 
<< pdiffusion >>
rect 67 139 68 140 
<< pdiffusion >>
rect 68 139 69 140 
<< pdiffusion >>
rect 69 139 70 140 
<< pdiffusion >>
rect 70 139 71 140 
<< pdiffusion >>
rect 71 139 72 140 
<< m1 >>
rect 73 139 74 140 
<< m1 >>
rect 79 139 80 140 
<< m1 >>
rect 81 139 82 140 
<< m2 >>
rect 81 139 82 140 
<< pdiffusion >>
rect 84 139 85 140 
<< pdiffusion >>
rect 85 139 86 140 
<< pdiffusion >>
rect 86 139 87 140 
<< pdiffusion >>
rect 87 139 88 140 
<< pdiffusion >>
rect 88 139 89 140 
<< pdiffusion >>
rect 89 139 90 140 
<< m1 >>
rect 100 139 101 140 
<< pdiffusion >>
rect 102 139 103 140 
<< pdiffusion >>
rect 103 139 104 140 
<< pdiffusion >>
rect 104 139 105 140 
<< pdiffusion >>
rect 105 139 106 140 
<< pdiffusion >>
rect 106 139 107 140 
<< pdiffusion >>
rect 107 139 108 140 
<< pdiffusion >>
rect 120 139 121 140 
<< pdiffusion >>
rect 121 139 122 140 
<< pdiffusion >>
rect 122 139 123 140 
<< pdiffusion >>
rect 123 139 124 140 
<< pdiffusion >>
rect 124 139 125 140 
<< pdiffusion >>
rect 125 139 126 140 
<< pdiffusion >>
rect 138 139 139 140 
<< pdiffusion >>
rect 139 139 140 140 
<< pdiffusion >>
rect 140 139 141 140 
<< pdiffusion >>
rect 141 139 142 140 
<< pdiffusion >>
rect 142 139 143 140 
<< pdiffusion >>
rect 143 139 144 140 
<< m1 >>
rect 145 139 146 140 
<< m2 >>
rect 145 139 146 140 
<< m1 >>
rect 147 139 148 140 
<< m1 >>
rect 151 139 152 140 
<< m1 >>
rect 154 139 155 140 
<< pdiffusion >>
rect 156 139 157 140 
<< pdiffusion >>
rect 157 139 158 140 
<< pdiffusion >>
rect 158 139 159 140 
<< pdiffusion >>
rect 159 139 160 140 
<< pdiffusion >>
rect 160 139 161 140 
<< pdiffusion >>
rect 161 139 162 140 
<< m1 >>
rect 163 139 164 140 
<< m1 >>
rect 10 140 11 141 
<< pdiffusion >>
rect 12 140 13 141 
<< pdiffusion >>
rect 13 140 14 141 
<< pdiffusion >>
rect 14 140 15 141 
<< pdiffusion >>
rect 15 140 16 141 
<< pdiffusion >>
rect 16 140 17 141 
<< pdiffusion >>
rect 17 140 18 141 
<< m1 >>
rect 22 140 23 141 
<< m1 >>
rect 25 140 26 141 
<< m1 >>
rect 27 140 28 141 
<< pdiffusion >>
rect 30 140 31 141 
<< pdiffusion >>
rect 31 140 32 141 
<< pdiffusion >>
rect 32 140 33 141 
<< pdiffusion >>
rect 33 140 34 141 
<< pdiffusion >>
rect 34 140 35 141 
<< pdiffusion >>
rect 35 140 36 141 
<< m1 >>
rect 41 140 42 141 
<< m1 >>
rect 43 140 44 141 
<< m1 >>
rect 45 140 46 141 
<< pdiffusion >>
rect 48 140 49 141 
<< pdiffusion >>
rect 49 140 50 141 
<< pdiffusion >>
rect 50 140 51 141 
<< pdiffusion >>
rect 51 140 52 141 
<< pdiffusion >>
rect 52 140 53 141 
<< pdiffusion >>
rect 53 140 54 141 
<< m1 >>
rect 64 140 65 141 
<< m2 >>
rect 64 140 65 141 
<< pdiffusion >>
rect 66 140 67 141 
<< pdiffusion >>
rect 67 140 68 141 
<< pdiffusion >>
rect 68 140 69 141 
<< pdiffusion >>
rect 69 140 70 141 
<< pdiffusion >>
rect 70 140 71 141 
<< pdiffusion >>
rect 71 140 72 141 
<< m1 >>
rect 73 140 74 141 
<< m1 >>
rect 79 140 80 141 
<< m1 >>
rect 81 140 82 141 
<< m2 >>
rect 81 140 82 141 
<< pdiffusion >>
rect 84 140 85 141 
<< pdiffusion >>
rect 85 140 86 141 
<< pdiffusion >>
rect 86 140 87 141 
<< pdiffusion >>
rect 87 140 88 141 
<< pdiffusion >>
rect 88 140 89 141 
<< pdiffusion >>
rect 89 140 90 141 
<< m1 >>
rect 100 140 101 141 
<< pdiffusion >>
rect 102 140 103 141 
<< pdiffusion >>
rect 103 140 104 141 
<< pdiffusion >>
rect 104 140 105 141 
<< pdiffusion >>
rect 105 140 106 141 
<< pdiffusion >>
rect 106 140 107 141 
<< pdiffusion >>
rect 107 140 108 141 
<< pdiffusion >>
rect 120 140 121 141 
<< pdiffusion >>
rect 121 140 122 141 
<< pdiffusion >>
rect 122 140 123 141 
<< pdiffusion >>
rect 123 140 124 141 
<< pdiffusion >>
rect 124 140 125 141 
<< pdiffusion >>
rect 125 140 126 141 
<< pdiffusion >>
rect 138 140 139 141 
<< pdiffusion >>
rect 139 140 140 141 
<< pdiffusion >>
rect 140 140 141 141 
<< pdiffusion >>
rect 141 140 142 141 
<< pdiffusion >>
rect 142 140 143 141 
<< pdiffusion >>
rect 143 140 144 141 
<< m1 >>
rect 145 140 146 141 
<< m2 >>
rect 145 140 146 141 
<< m1 >>
rect 147 140 148 141 
<< m1 >>
rect 151 140 152 141 
<< m1 >>
rect 154 140 155 141 
<< pdiffusion >>
rect 156 140 157 141 
<< pdiffusion >>
rect 157 140 158 141 
<< pdiffusion >>
rect 158 140 159 141 
<< pdiffusion >>
rect 159 140 160 141 
<< pdiffusion >>
rect 160 140 161 141 
<< pdiffusion >>
rect 161 140 162 141 
<< m1 >>
rect 163 140 164 141 
<< m1 >>
rect 10 141 11 142 
<< pdiffusion >>
rect 12 141 13 142 
<< pdiffusion >>
rect 13 141 14 142 
<< pdiffusion >>
rect 14 141 15 142 
<< pdiffusion >>
rect 15 141 16 142 
<< pdiffusion >>
rect 16 141 17 142 
<< pdiffusion >>
rect 17 141 18 142 
<< m1 >>
rect 22 141 23 142 
<< m1 >>
rect 25 141 26 142 
<< m1 >>
rect 27 141 28 142 
<< pdiffusion >>
rect 30 141 31 142 
<< pdiffusion >>
rect 31 141 32 142 
<< pdiffusion >>
rect 32 141 33 142 
<< pdiffusion >>
rect 33 141 34 142 
<< pdiffusion >>
rect 34 141 35 142 
<< pdiffusion >>
rect 35 141 36 142 
<< m1 >>
rect 41 141 42 142 
<< m1 >>
rect 43 141 44 142 
<< m1 >>
rect 45 141 46 142 
<< pdiffusion >>
rect 48 141 49 142 
<< pdiffusion >>
rect 49 141 50 142 
<< pdiffusion >>
rect 50 141 51 142 
<< pdiffusion >>
rect 51 141 52 142 
<< pdiffusion >>
rect 52 141 53 142 
<< pdiffusion >>
rect 53 141 54 142 
<< m1 >>
rect 64 141 65 142 
<< m2 >>
rect 64 141 65 142 
<< pdiffusion >>
rect 66 141 67 142 
<< pdiffusion >>
rect 67 141 68 142 
<< pdiffusion >>
rect 68 141 69 142 
<< pdiffusion >>
rect 69 141 70 142 
<< pdiffusion >>
rect 70 141 71 142 
<< pdiffusion >>
rect 71 141 72 142 
<< m1 >>
rect 73 141 74 142 
<< m1 >>
rect 79 141 80 142 
<< m1 >>
rect 81 141 82 142 
<< m2 >>
rect 81 141 82 142 
<< pdiffusion >>
rect 84 141 85 142 
<< pdiffusion >>
rect 85 141 86 142 
<< pdiffusion >>
rect 86 141 87 142 
<< pdiffusion >>
rect 87 141 88 142 
<< pdiffusion >>
rect 88 141 89 142 
<< pdiffusion >>
rect 89 141 90 142 
<< m1 >>
rect 100 141 101 142 
<< pdiffusion >>
rect 102 141 103 142 
<< pdiffusion >>
rect 103 141 104 142 
<< pdiffusion >>
rect 104 141 105 142 
<< pdiffusion >>
rect 105 141 106 142 
<< pdiffusion >>
rect 106 141 107 142 
<< pdiffusion >>
rect 107 141 108 142 
<< pdiffusion >>
rect 120 141 121 142 
<< pdiffusion >>
rect 121 141 122 142 
<< pdiffusion >>
rect 122 141 123 142 
<< pdiffusion >>
rect 123 141 124 142 
<< pdiffusion >>
rect 124 141 125 142 
<< pdiffusion >>
rect 125 141 126 142 
<< pdiffusion >>
rect 138 141 139 142 
<< pdiffusion >>
rect 139 141 140 142 
<< pdiffusion >>
rect 140 141 141 142 
<< pdiffusion >>
rect 141 141 142 142 
<< pdiffusion >>
rect 142 141 143 142 
<< pdiffusion >>
rect 143 141 144 142 
<< m1 >>
rect 145 141 146 142 
<< m2 >>
rect 145 141 146 142 
<< m1 >>
rect 147 141 148 142 
<< m1 >>
rect 151 141 152 142 
<< m1 >>
rect 154 141 155 142 
<< pdiffusion >>
rect 156 141 157 142 
<< pdiffusion >>
rect 157 141 158 142 
<< pdiffusion >>
rect 158 141 159 142 
<< pdiffusion >>
rect 159 141 160 142 
<< pdiffusion >>
rect 160 141 161 142 
<< pdiffusion >>
rect 161 141 162 142 
<< m1 >>
rect 163 141 164 142 
<< m1 >>
rect 10 142 11 143 
<< pdiffusion >>
rect 12 142 13 143 
<< pdiffusion >>
rect 13 142 14 143 
<< pdiffusion >>
rect 14 142 15 143 
<< pdiffusion >>
rect 15 142 16 143 
<< pdiffusion >>
rect 16 142 17 143 
<< pdiffusion >>
rect 17 142 18 143 
<< m1 >>
rect 22 142 23 143 
<< m1 >>
rect 25 142 26 143 
<< m1 >>
rect 27 142 28 143 
<< pdiffusion >>
rect 30 142 31 143 
<< pdiffusion >>
rect 31 142 32 143 
<< pdiffusion >>
rect 32 142 33 143 
<< pdiffusion >>
rect 33 142 34 143 
<< pdiffusion >>
rect 34 142 35 143 
<< pdiffusion >>
rect 35 142 36 143 
<< m1 >>
rect 41 142 42 143 
<< m1 >>
rect 43 142 44 143 
<< m1 >>
rect 45 142 46 143 
<< pdiffusion >>
rect 48 142 49 143 
<< pdiffusion >>
rect 49 142 50 143 
<< pdiffusion >>
rect 50 142 51 143 
<< pdiffusion >>
rect 51 142 52 143 
<< pdiffusion >>
rect 52 142 53 143 
<< pdiffusion >>
rect 53 142 54 143 
<< m1 >>
rect 64 142 65 143 
<< m2 >>
rect 64 142 65 143 
<< pdiffusion >>
rect 66 142 67 143 
<< pdiffusion >>
rect 67 142 68 143 
<< pdiffusion >>
rect 68 142 69 143 
<< pdiffusion >>
rect 69 142 70 143 
<< pdiffusion >>
rect 70 142 71 143 
<< pdiffusion >>
rect 71 142 72 143 
<< m1 >>
rect 73 142 74 143 
<< m1 >>
rect 79 142 80 143 
<< m1 >>
rect 81 142 82 143 
<< m2 >>
rect 81 142 82 143 
<< pdiffusion >>
rect 84 142 85 143 
<< pdiffusion >>
rect 85 142 86 143 
<< pdiffusion >>
rect 86 142 87 143 
<< pdiffusion >>
rect 87 142 88 143 
<< pdiffusion >>
rect 88 142 89 143 
<< pdiffusion >>
rect 89 142 90 143 
<< m1 >>
rect 100 142 101 143 
<< pdiffusion >>
rect 102 142 103 143 
<< pdiffusion >>
rect 103 142 104 143 
<< pdiffusion >>
rect 104 142 105 143 
<< pdiffusion >>
rect 105 142 106 143 
<< pdiffusion >>
rect 106 142 107 143 
<< pdiffusion >>
rect 107 142 108 143 
<< pdiffusion >>
rect 120 142 121 143 
<< pdiffusion >>
rect 121 142 122 143 
<< pdiffusion >>
rect 122 142 123 143 
<< pdiffusion >>
rect 123 142 124 143 
<< pdiffusion >>
rect 124 142 125 143 
<< pdiffusion >>
rect 125 142 126 143 
<< pdiffusion >>
rect 138 142 139 143 
<< pdiffusion >>
rect 139 142 140 143 
<< pdiffusion >>
rect 140 142 141 143 
<< pdiffusion >>
rect 141 142 142 143 
<< pdiffusion >>
rect 142 142 143 143 
<< pdiffusion >>
rect 143 142 144 143 
<< m1 >>
rect 145 142 146 143 
<< m2 >>
rect 145 142 146 143 
<< m1 >>
rect 147 142 148 143 
<< m1 >>
rect 151 142 152 143 
<< m1 >>
rect 154 142 155 143 
<< pdiffusion >>
rect 156 142 157 143 
<< pdiffusion >>
rect 157 142 158 143 
<< pdiffusion >>
rect 158 142 159 143 
<< pdiffusion >>
rect 159 142 160 143 
<< pdiffusion >>
rect 160 142 161 143 
<< pdiffusion >>
rect 161 142 162 143 
<< m1 >>
rect 163 142 164 143 
<< m1 >>
rect 10 143 11 144 
<< pdiffusion >>
rect 12 143 13 144 
<< m1 >>
rect 13 143 14 144 
<< pdiffusion >>
rect 13 143 14 144 
<< pdiffusion >>
rect 14 143 15 144 
<< pdiffusion >>
rect 15 143 16 144 
<< pdiffusion >>
rect 16 143 17 144 
<< pdiffusion >>
rect 17 143 18 144 
<< m1 >>
rect 22 143 23 144 
<< m1 >>
rect 25 143 26 144 
<< m1 >>
rect 27 143 28 144 
<< pdiffusion >>
rect 30 143 31 144 
<< pdiffusion >>
rect 31 143 32 144 
<< pdiffusion >>
rect 32 143 33 144 
<< pdiffusion >>
rect 33 143 34 144 
<< m1 >>
rect 34 143 35 144 
<< pdiffusion >>
rect 34 143 35 144 
<< pdiffusion >>
rect 35 143 36 144 
<< m1 >>
rect 41 143 42 144 
<< m1 >>
rect 43 143 44 144 
<< m1 >>
rect 45 143 46 144 
<< pdiffusion >>
rect 48 143 49 144 
<< m1 >>
rect 49 143 50 144 
<< pdiffusion >>
rect 49 143 50 144 
<< pdiffusion >>
rect 50 143 51 144 
<< pdiffusion >>
rect 51 143 52 144 
<< pdiffusion >>
rect 52 143 53 144 
<< pdiffusion >>
rect 53 143 54 144 
<< m1 >>
rect 64 143 65 144 
<< m2 >>
rect 64 143 65 144 
<< pdiffusion >>
rect 66 143 67 144 
<< pdiffusion >>
rect 67 143 68 144 
<< pdiffusion >>
rect 68 143 69 144 
<< pdiffusion >>
rect 69 143 70 144 
<< m1 >>
rect 70 143 71 144 
<< pdiffusion >>
rect 70 143 71 144 
<< pdiffusion >>
rect 71 143 72 144 
<< m1 >>
rect 73 143 74 144 
<< m1 >>
rect 79 143 80 144 
<< m1 >>
rect 81 143 82 144 
<< m2 >>
rect 81 143 82 144 
<< pdiffusion >>
rect 84 143 85 144 
<< pdiffusion >>
rect 85 143 86 144 
<< pdiffusion >>
rect 86 143 87 144 
<< pdiffusion >>
rect 87 143 88 144 
<< pdiffusion >>
rect 88 143 89 144 
<< pdiffusion >>
rect 89 143 90 144 
<< m1 >>
rect 100 143 101 144 
<< pdiffusion >>
rect 102 143 103 144 
<< m1 >>
rect 103 143 104 144 
<< pdiffusion >>
rect 103 143 104 144 
<< pdiffusion >>
rect 104 143 105 144 
<< pdiffusion >>
rect 105 143 106 144 
<< pdiffusion >>
rect 106 143 107 144 
<< pdiffusion >>
rect 107 143 108 144 
<< pdiffusion >>
rect 120 143 121 144 
<< pdiffusion >>
rect 121 143 122 144 
<< pdiffusion >>
rect 122 143 123 144 
<< pdiffusion >>
rect 123 143 124 144 
<< pdiffusion >>
rect 124 143 125 144 
<< pdiffusion >>
rect 125 143 126 144 
<< pdiffusion >>
rect 138 143 139 144 
<< m1 >>
rect 139 143 140 144 
<< pdiffusion >>
rect 139 143 140 144 
<< pdiffusion >>
rect 140 143 141 144 
<< pdiffusion >>
rect 141 143 142 144 
<< m1 >>
rect 142 143 143 144 
<< pdiffusion >>
rect 142 143 143 144 
<< pdiffusion >>
rect 143 143 144 144 
<< m1 >>
rect 145 143 146 144 
<< m2 >>
rect 145 143 146 144 
<< m1 >>
rect 147 143 148 144 
<< m1 >>
rect 151 143 152 144 
<< m1 >>
rect 154 143 155 144 
<< pdiffusion >>
rect 156 143 157 144 
<< pdiffusion >>
rect 157 143 158 144 
<< pdiffusion >>
rect 158 143 159 144 
<< pdiffusion >>
rect 159 143 160 144 
<< pdiffusion >>
rect 160 143 161 144 
<< pdiffusion >>
rect 161 143 162 144 
<< m1 >>
rect 163 143 164 144 
<< m1 >>
rect 10 144 11 145 
<< m1 >>
rect 13 144 14 145 
<< m1 >>
rect 22 144 23 145 
<< m1 >>
rect 25 144 26 145 
<< m1 >>
rect 27 144 28 145 
<< m1 >>
rect 34 144 35 145 
<< m1 >>
rect 41 144 42 145 
<< m1 >>
rect 43 144 44 145 
<< m1 >>
rect 45 144 46 145 
<< m1 >>
rect 49 144 50 145 
<< m1 >>
rect 64 144 65 145 
<< m2 >>
rect 64 144 65 145 
<< m1 >>
rect 70 144 71 145 
<< m1 >>
rect 73 144 74 145 
<< m1 >>
rect 77 144 78 145 
<< m2 >>
rect 77 144 78 145 
<< m2c >>
rect 77 144 78 145 
<< m1 >>
rect 77 144 78 145 
<< m2 >>
rect 77 144 78 145 
<< m2 >>
rect 78 144 79 145 
<< m1 >>
rect 79 144 80 145 
<< m2 >>
rect 79 144 80 145 
<< m2 >>
rect 80 144 81 145 
<< m1 >>
rect 81 144 82 145 
<< m2 >>
rect 81 144 82 145 
<< m1 >>
rect 100 144 101 145 
<< m1 >>
rect 103 144 104 145 
<< m1 >>
rect 139 144 140 145 
<< m1 >>
rect 142 144 143 145 
<< m1 >>
rect 145 144 146 145 
<< m2 >>
rect 145 144 146 145 
<< m1 >>
rect 147 144 148 145 
<< m1 >>
rect 151 144 152 145 
<< m1 >>
rect 154 144 155 145 
<< m1 >>
rect 163 144 164 145 
<< m1 >>
rect 10 145 11 146 
<< m2 >>
rect 10 145 11 146 
<< m2 >>
rect 11 145 12 146 
<< m1 >>
rect 12 145 13 146 
<< m2 >>
rect 12 145 13 146 
<< m2c >>
rect 12 145 13 146 
<< m1 >>
rect 12 145 13 146 
<< m2 >>
rect 12 145 13 146 
<< m1 >>
rect 13 145 14 146 
<< m1 >>
rect 22 145 23 146 
<< m1 >>
rect 25 145 26 146 
<< m1 >>
rect 27 145 28 146 
<< m1 >>
rect 34 145 35 146 
<< m1 >>
rect 41 145 42 146 
<< m1 >>
rect 43 145 44 146 
<< m1 >>
rect 45 145 46 146 
<< m1 >>
rect 49 145 50 146 
<< m1 >>
rect 64 145 65 146 
<< m2 >>
rect 64 145 65 146 
<< m1 >>
rect 70 145 71 146 
<< m1 >>
rect 73 145 74 146 
<< m1 >>
rect 77 145 78 146 
<< m1 >>
rect 79 145 80 146 
<< m1 >>
rect 81 145 82 146 
<< m1 >>
rect 100 145 101 146 
<< m1 >>
rect 103 145 104 146 
<< m1 >>
rect 139 145 140 146 
<< m1 >>
rect 142 145 143 146 
<< m1 >>
rect 143 145 144 146 
<< m1 >>
rect 144 145 145 146 
<< m1 >>
rect 145 145 146 146 
<< m2 >>
rect 145 145 146 146 
<< m1 >>
rect 147 145 148 146 
<< m1 >>
rect 151 145 152 146 
<< m1 >>
rect 154 145 155 146 
<< m1 >>
rect 163 145 164 146 
<< m1 >>
rect 10 146 11 147 
<< m2 >>
rect 10 146 11 147 
<< m1 >>
rect 22 146 23 147 
<< m2 >>
rect 22 146 23 147 
<< m2c >>
rect 22 146 23 147 
<< m1 >>
rect 22 146 23 147 
<< m2 >>
rect 22 146 23 147 
<< m1 >>
rect 25 146 26 147 
<< m2 >>
rect 25 146 26 147 
<< m2c >>
rect 25 146 26 147 
<< m1 >>
rect 25 146 26 147 
<< m2 >>
rect 25 146 26 147 
<< m1 >>
rect 27 146 28 147 
<< m2 >>
rect 27 146 28 147 
<< m2c >>
rect 27 146 28 147 
<< m1 >>
rect 27 146 28 147 
<< m2 >>
rect 27 146 28 147 
<< m1 >>
rect 34 146 35 147 
<< m2 >>
rect 34 146 35 147 
<< m2c >>
rect 34 146 35 147 
<< m1 >>
rect 34 146 35 147 
<< m2 >>
rect 34 146 35 147 
<< m1 >>
rect 41 146 42 147 
<< m2 >>
rect 41 146 42 147 
<< m2c >>
rect 41 146 42 147 
<< m1 >>
rect 41 146 42 147 
<< m2 >>
rect 41 146 42 147 
<< m1 >>
rect 43 146 44 147 
<< m2 >>
rect 43 146 44 147 
<< m2c >>
rect 43 146 44 147 
<< m1 >>
rect 43 146 44 147 
<< m2 >>
rect 43 146 44 147 
<< m1 >>
rect 45 146 46 147 
<< m2 >>
rect 45 146 46 147 
<< m2c >>
rect 45 146 46 147 
<< m1 >>
rect 45 146 46 147 
<< m2 >>
rect 45 146 46 147 
<< m1 >>
rect 49 146 50 147 
<< m1 >>
rect 50 146 51 147 
<< m1 >>
rect 51 146 52 147 
<< m1 >>
rect 52 146 53 147 
<< m1 >>
rect 53 146 54 147 
<< m1 >>
rect 54 146 55 147 
<< m1 >>
rect 55 146 56 147 
<< m1 >>
rect 56 146 57 147 
<< m1 >>
rect 57 146 58 147 
<< m1 >>
rect 58 146 59 147 
<< m1 >>
rect 59 146 60 147 
<< m1 >>
rect 60 146 61 147 
<< m1 >>
rect 61 146 62 147 
<< m1 >>
rect 62 146 63 147 
<< m1 >>
rect 63 146 64 147 
<< m1 >>
rect 64 146 65 147 
<< m2 >>
rect 64 146 65 147 
<< m1 >>
rect 70 146 71 147 
<< m2 >>
rect 70 146 71 147 
<< m2c >>
rect 70 146 71 147 
<< m1 >>
rect 70 146 71 147 
<< m2 >>
rect 70 146 71 147 
<< m1 >>
rect 73 146 74 147 
<< m2 >>
rect 73 146 74 147 
<< m2c >>
rect 73 146 74 147 
<< m1 >>
rect 73 146 74 147 
<< m2 >>
rect 73 146 74 147 
<< m1 >>
rect 77 146 78 147 
<< m2 >>
rect 77 146 78 147 
<< m2c >>
rect 77 146 78 147 
<< m1 >>
rect 77 146 78 147 
<< m2 >>
rect 77 146 78 147 
<< m1 >>
rect 79 146 80 147 
<< m2 >>
rect 79 146 80 147 
<< m2c >>
rect 79 146 80 147 
<< m1 >>
rect 79 146 80 147 
<< m2 >>
rect 79 146 80 147 
<< m1 >>
rect 81 146 82 147 
<< m2 >>
rect 81 146 82 147 
<< m2c >>
rect 81 146 82 147 
<< m1 >>
rect 81 146 82 147 
<< m2 >>
rect 81 146 82 147 
<< m1 >>
rect 100 146 101 147 
<< m2 >>
rect 100 146 101 147 
<< m2c >>
rect 100 146 101 147 
<< m1 >>
rect 100 146 101 147 
<< m2 >>
rect 100 146 101 147 
<< m1 >>
rect 102 146 103 147 
<< m2 >>
rect 102 146 103 147 
<< m2c >>
rect 102 146 103 147 
<< m1 >>
rect 102 146 103 147 
<< m2 >>
rect 102 146 103 147 
<< m1 >>
rect 103 146 104 147 
<< m1 >>
rect 139 146 140 147 
<< m1 >>
rect 140 146 141 147 
<< m2 >>
rect 140 146 141 147 
<< m2c >>
rect 140 146 141 147 
<< m1 >>
rect 140 146 141 147 
<< m2 >>
rect 140 146 141 147 
<< m2 >>
rect 141 146 142 147 
<< m2 >>
rect 142 146 143 147 
<< m2 >>
rect 143 146 144 147 
<< m2 >>
rect 144 146 145 147 
<< m2 >>
rect 145 146 146 147 
<< m1 >>
rect 147 146 148 147 
<< m2 >>
rect 147 146 148 147 
<< m2c >>
rect 147 146 148 147 
<< m1 >>
rect 147 146 148 147 
<< m2 >>
rect 147 146 148 147 
<< m1 >>
rect 151 146 152 147 
<< m2 >>
rect 151 146 152 147 
<< m2c >>
rect 151 146 152 147 
<< m1 >>
rect 151 146 152 147 
<< m2 >>
rect 151 146 152 147 
<< m1 >>
rect 154 146 155 147 
<< m1 >>
rect 155 146 156 147 
<< m1 >>
rect 156 146 157 147 
<< m2 >>
rect 156 146 157 147 
<< m2c >>
rect 156 146 157 147 
<< m1 >>
rect 156 146 157 147 
<< m2 >>
rect 156 146 157 147 
<< m1 >>
rect 163 146 164 147 
<< m1 >>
rect 10 147 11 148 
<< m2 >>
rect 10 147 11 148 
<< m2 >>
rect 22 147 23 148 
<< m2 >>
rect 25 147 26 148 
<< m2 >>
rect 27 147 28 148 
<< m2 >>
rect 34 147 35 148 
<< m2 >>
rect 38 147 39 148 
<< m2 >>
rect 39 147 40 148 
<< m2 >>
rect 40 147 41 148 
<< m2 >>
rect 41 147 42 148 
<< m2 >>
rect 43 147 44 148 
<< m2 >>
rect 45 147 46 148 
<< m2 >>
rect 64 147 65 148 
<< m2 >>
rect 70 147 71 148 
<< m2 >>
rect 73 147 74 148 
<< m2 >>
rect 77 147 78 148 
<< m2 >>
rect 79 147 80 148 
<< m2 >>
rect 81 147 82 148 
<< m2 >>
rect 100 147 101 148 
<< m2 >>
rect 102 147 103 148 
<< m2 >>
rect 147 147 148 148 
<< m2 >>
rect 151 147 152 148 
<< m2 >>
rect 156 147 157 148 
<< m1 >>
rect 163 147 164 148 
<< m1 >>
rect 10 148 11 149 
<< m2 >>
rect 10 148 11 149 
<< m1 >>
rect 13 148 14 149 
<< m1 >>
rect 14 148 15 149 
<< m1 >>
rect 15 148 16 149 
<< m1 >>
rect 16 148 17 149 
<< m1 >>
rect 17 148 18 149 
<< m1 >>
rect 18 148 19 149 
<< m1 >>
rect 19 148 20 149 
<< m1 >>
rect 20 148 21 149 
<< m1 >>
rect 21 148 22 149 
<< m1 >>
rect 22 148 23 149 
<< m2 >>
rect 22 148 23 149 
<< m1 >>
rect 23 148 24 149 
<< m1 >>
rect 24 148 25 149 
<< m1 >>
rect 25 148 26 149 
<< m2 >>
rect 25 148 26 149 
<< m1 >>
rect 26 148 27 149 
<< m1 >>
rect 27 148 28 149 
<< m2 >>
rect 27 148 28 149 
<< m1 >>
rect 28 148 29 149 
<< m1 >>
rect 29 148 30 149 
<< m1 >>
rect 30 148 31 149 
<< m1 >>
rect 31 148 32 149 
<< m1 >>
rect 32 148 33 149 
<< m1 >>
rect 33 148 34 149 
<< m1 >>
rect 34 148 35 149 
<< m2 >>
rect 34 148 35 149 
<< m1 >>
rect 35 148 36 149 
<< m1 >>
rect 36 148 37 149 
<< m1 >>
rect 37 148 38 149 
<< m1 >>
rect 38 148 39 149 
<< m2 >>
rect 38 148 39 149 
<< m1 >>
rect 39 148 40 149 
<< m1 >>
rect 40 148 41 149 
<< m1 >>
rect 41 148 42 149 
<< m1 >>
rect 42 148 43 149 
<< m1 >>
rect 43 148 44 149 
<< m2 >>
rect 43 148 44 149 
<< m1 >>
rect 44 148 45 149 
<< m1 >>
rect 45 148 46 149 
<< m2 >>
rect 45 148 46 149 
<< m1 >>
rect 46 148 47 149 
<< m1 >>
rect 47 148 48 149 
<< m1 >>
rect 48 148 49 149 
<< m1 >>
rect 49 148 50 149 
<< m1 >>
rect 50 148 51 149 
<< m1 >>
rect 51 148 52 149 
<< m1 >>
rect 52 148 53 149 
<< m1 >>
rect 53 148 54 149 
<< m1 >>
rect 54 148 55 149 
<< m1 >>
rect 55 148 56 149 
<< m1 >>
rect 56 148 57 149 
<< m1 >>
rect 57 148 58 149 
<< m1 >>
rect 58 148 59 149 
<< m1 >>
rect 59 148 60 149 
<< m1 >>
rect 60 148 61 149 
<< m1 >>
rect 61 148 62 149 
<< m1 >>
rect 62 148 63 149 
<< m1 >>
rect 63 148 64 149 
<< m1 >>
rect 64 148 65 149 
<< m2 >>
rect 64 148 65 149 
<< m1 >>
rect 65 148 66 149 
<< m1 >>
rect 66 148 67 149 
<< m2 >>
rect 66 148 67 149 
<< m1 >>
rect 67 148 68 149 
<< m2 >>
rect 67 148 68 149 
<< m1 >>
rect 68 148 69 149 
<< m2 >>
rect 68 148 69 149 
<< m1 >>
rect 69 148 70 149 
<< m2 >>
rect 69 148 70 149 
<< m1 >>
rect 70 148 71 149 
<< m2 >>
rect 70 148 71 149 
<< m1 >>
rect 71 148 72 149 
<< m1 >>
rect 72 148 73 149 
<< m1 >>
rect 73 148 74 149 
<< m2 >>
rect 73 148 74 149 
<< m1 >>
rect 74 148 75 149 
<< m1 >>
rect 75 148 76 149 
<< m1 >>
rect 76 148 77 149 
<< m1 >>
rect 77 148 78 149 
<< m2 >>
rect 77 148 78 149 
<< m1 >>
rect 78 148 79 149 
<< m1 >>
rect 79 148 80 149 
<< m2 >>
rect 79 148 80 149 
<< m1 >>
rect 80 148 81 149 
<< m1 >>
rect 81 148 82 149 
<< m2 >>
rect 81 148 82 149 
<< m1 >>
rect 82 148 83 149 
<< m1 >>
rect 83 148 84 149 
<< m1 >>
rect 84 148 85 149 
<< m1 >>
rect 85 148 86 149 
<< m1 >>
rect 86 148 87 149 
<< m1 >>
rect 87 148 88 149 
<< m1 >>
rect 88 148 89 149 
<< m1 >>
rect 89 148 90 149 
<< m1 >>
rect 90 148 91 149 
<< m1 >>
rect 91 148 92 149 
<< m1 >>
rect 92 148 93 149 
<< m1 >>
rect 93 148 94 149 
<< m1 >>
rect 94 148 95 149 
<< m1 >>
rect 95 148 96 149 
<< m1 >>
rect 96 148 97 149 
<< m1 >>
rect 97 148 98 149 
<< m1 >>
rect 98 148 99 149 
<< m1 >>
rect 99 148 100 149 
<< m1 >>
rect 100 148 101 149 
<< m2 >>
rect 100 148 101 149 
<< m1 >>
rect 101 148 102 149 
<< m1 >>
rect 102 148 103 149 
<< m2 >>
rect 102 148 103 149 
<< m1 >>
rect 103 148 104 149 
<< m1 >>
rect 104 148 105 149 
<< m1 >>
rect 105 148 106 149 
<< m1 >>
rect 106 148 107 149 
<< m1 >>
rect 107 148 108 149 
<< m1 >>
rect 108 148 109 149 
<< m1 >>
rect 109 148 110 149 
<< m1 >>
rect 110 148 111 149 
<< m1 >>
rect 111 148 112 149 
<< m1 >>
rect 112 148 113 149 
<< m1 >>
rect 113 148 114 149 
<< m1 >>
rect 114 148 115 149 
<< m1 >>
rect 115 148 116 149 
<< m1 >>
rect 116 148 117 149 
<< m1 >>
rect 117 148 118 149 
<< m1 >>
rect 118 148 119 149 
<< m1 >>
rect 119 148 120 149 
<< m1 >>
rect 120 148 121 149 
<< m1 >>
rect 121 148 122 149 
<< m1 >>
rect 122 148 123 149 
<< m1 >>
rect 123 148 124 149 
<< m1 >>
rect 124 148 125 149 
<< m1 >>
rect 125 148 126 149 
<< m1 >>
rect 126 148 127 149 
<< m1 >>
rect 127 148 128 149 
<< m1 >>
rect 128 148 129 149 
<< m1 >>
rect 129 148 130 149 
<< m1 >>
rect 130 148 131 149 
<< m1 >>
rect 131 148 132 149 
<< m1 >>
rect 132 148 133 149 
<< m1 >>
rect 133 148 134 149 
<< m1 >>
rect 134 148 135 149 
<< m1 >>
rect 135 148 136 149 
<< m1 >>
rect 136 148 137 149 
<< m1 >>
rect 137 148 138 149 
<< m1 >>
rect 138 148 139 149 
<< m1 >>
rect 139 148 140 149 
<< m1 >>
rect 140 148 141 149 
<< m1 >>
rect 141 148 142 149 
<< m1 >>
rect 142 148 143 149 
<< m1 >>
rect 143 148 144 149 
<< m1 >>
rect 144 148 145 149 
<< m1 >>
rect 145 148 146 149 
<< m1 >>
rect 146 148 147 149 
<< m1 >>
rect 147 148 148 149 
<< m2 >>
rect 147 148 148 149 
<< m1 >>
rect 148 148 149 149 
<< m1 >>
rect 149 148 150 149 
<< m1 >>
rect 150 148 151 149 
<< m1 >>
rect 151 148 152 149 
<< m2 >>
rect 151 148 152 149 
<< m1 >>
rect 152 148 153 149 
<< m1 >>
rect 153 148 154 149 
<< m1 >>
rect 154 148 155 149 
<< m1 >>
rect 155 148 156 149 
<< m1 >>
rect 156 148 157 149 
<< m2 >>
rect 156 148 157 149 
<< m1 >>
rect 157 148 158 149 
<< m1 >>
rect 158 148 159 149 
<< m1 >>
rect 159 148 160 149 
<< m1 >>
rect 160 148 161 149 
<< m1 >>
rect 161 148 162 149 
<< m1 >>
rect 162 148 163 149 
<< m1 >>
rect 163 148 164 149 
<< m1 >>
rect 10 149 11 150 
<< m2 >>
rect 10 149 11 150 
<< m1 >>
rect 13 149 14 150 
<< m2 >>
rect 22 149 23 150 
<< m2 >>
rect 25 149 26 150 
<< m2 >>
rect 27 149 28 150 
<< m2 >>
rect 34 149 35 150 
<< m2 >>
rect 38 149 39 150 
<< m2 >>
rect 43 149 44 150 
<< m2 >>
rect 45 149 46 150 
<< m2 >>
rect 64 149 65 150 
<< m2 >>
rect 66 149 67 150 
<< m2 >>
rect 73 149 74 150 
<< m2 >>
rect 77 149 78 150 
<< m2 >>
rect 79 149 80 150 
<< m2 >>
rect 81 149 82 150 
<< m2 >>
rect 100 149 101 150 
<< m2 >>
rect 102 149 103 150 
<< m2 >>
rect 147 149 148 150 
<< m2 >>
rect 151 149 152 150 
<< m2 >>
rect 156 149 157 150 
<< m1 >>
rect 10 150 11 151 
<< m2 >>
rect 10 150 11 151 
<< m1 >>
rect 13 150 14 151 
<< m1 >>
rect 22 150 23 151 
<< m2 >>
rect 22 150 23 151 
<< m2c >>
rect 22 150 23 151 
<< m1 >>
rect 22 150 23 151 
<< m2 >>
rect 22 150 23 151 
<< m1 >>
rect 25 150 26 151 
<< m2 >>
rect 25 150 26 151 
<< m2c >>
rect 25 150 26 151 
<< m1 >>
rect 25 150 26 151 
<< m2 >>
rect 25 150 26 151 
<< m1 >>
rect 27 150 28 151 
<< m2 >>
rect 27 150 28 151 
<< m2c >>
rect 27 150 28 151 
<< m1 >>
rect 27 150 28 151 
<< m2 >>
rect 27 150 28 151 
<< m2 >>
rect 34 150 35 151 
<< m2 >>
rect 38 150 39 151 
<< m2 >>
rect 43 150 44 151 
<< m2 >>
rect 45 150 46 151 
<< m1 >>
rect 49 150 50 151 
<< m1 >>
rect 50 150 51 151 
<< m1 >>
rect 51 150 52 151 
<< m1 >>
rect 52 150 53 151 
<< m1 >>
rect 53 150 54 151 
<< m1 >>
rect 54 150 55 151 
<< m1 >>
rect 55 150 56 151 
<< m1 >>
rect 56 150 57 151 
<< m1 >>
rect 57 150 58 151 
<< m1 >>
rect 58 150 59 151 
<< m1 >>
rect 59 150 60 151 
<< m1 >>
rect 60 150 61 151 
<< m1 >>
rect 61 150 62 151 
<< m1 >>
rect 62 150 63 151 
<< m1 >>
rect 63 150 64 151 
<< m1 >>
rect 64 150 65 151 
<< m2 >>
rect 64 150 65 151 
<< m2c >>
rect 64 150 65 151 
<< m1 >>
rect 64 150 65 151 
<< m2 >>
rect 64 150 65 151 
<< m2 >>
rect 66 150 67 151 
<< m1 >>
rect 73 150 74 151 
<< m2 >>
rect 73 150 74 151 
<< m2c >>
rect 73 150 74 151 
<< m1 >>
rect 73 150 74 151 
<< m2 >>
rect 73 150 74 151 
<< m1 >>
rect 77 150 78 151 
<< m2 >>
rect 77 150 78 151 
<< m2c >>
rect 77 150 78 151 
<< m1 >>
rect 77 150 78 151 
<< m2 >>
rect 77 150 78 151 
<< m1 >>
rect 79 150 80 151 
<< m2 >>
rect 79 150 80 151 
<< m2c >>
rect 79 150 80 151 
<< m1 >>
rect 79 150 80 151 
<< m2 >>
rect 79 150 80 151 
<< m1 >>
rect 81 150 82 151 
<< m2 >>
rect 81 150 82 151 
<< m2c >>
rect 81 150 82 151 
<< m1 >>
rect 81 150 82 151 
<< m2 >>
rect 81 150 82 151 
<< m1 >>
rect 100 150 101 151 
<< m2 >>
rect 100 150 101 151 
<< m2c >>
rect 100 150 101 151 
<< m1 >>
rect 100 150 101 151 
<< m2 >>
rect 100 150 101 151 
<< m1 >>
rect 102 150 103 151 
<< m2 >>
rect 102 150 103 151 
<< m2c >>
rect 102 150 103 151 
<< m1 >>
rect 102 150 103 151 
<< m2 >>
rect 102 150 103 151 
<< m1 >>
rect 147 150 148 151 
<< m2 >>
rect 147 150 148 151 
<< m2c >>
rect 147 150 148 151 
<< m1 >>
rect 147 150 148 151 
<< m2 >>
rect 147 150 148 151 
<< m1 >>
rect 148 150 149 151 
<< m1 >>
rect 149 150 150 151 
<< m1 >>
rect 150 150 151 151 
<< m1 >>
rect 151 150 152 151 
<< m2 >>
rect 151 150 152 151 
<< m1 >>
rect 152 150 153 151 
<< m1 >>
rect 153 150 154 151 
<< m1 >>
rect 154 150 155 151 
<< m1 >>
rect 155 150 156 151 
<< m1 >>
rect 156 150 157 151 
<< m2 >>
rect 156 150 157 151 
<< m1 >>
rect 157 150 158 151 
<< m1 >>
rect 158 150 159 151 
<< m1 >>
rect 159 150 160 151 
<< m1 >>
rect 160 150 161 151 
<< m1 >>
rect 161 150 162 151 
<< m1 >>
rect 162 150 163 151 
<< m1 >>
rect 163 150 164 151 
<< m1 >>
rect 10 151 11 152 
<< m2 >>
rect 10 151 11 152 
<< m1 >>
rect 13 151 14 152 
<< m1 >>
rect 22 151 23 152 
<< m1 >>
rect 25 151 26 152 
<< m1 >>
rect 27 151 28 152 
<< m1 >>
rect 31 151 32 152 
<< m1 >>
rect 32 151 33 152 
<< m1 >>
rect 33 151 34 152 
<< m1 >>
rect 34 151 35 152 
<< m2 >>
rect 34 151 35 152 
<< m1 >>
rect 35 151 36 152 
<< m1 >>
rect 36 151 37 152 
<< m1 >>
rect 37 151 38 152 
<< m1 >>
rect 38 151 39 152 
<< m2 >>
rect 38 151 39 152 
<< m1 >>
rect 39 151 40 152 
<< m1 >>
rect 40 151 41 152 
<< m1 >>
rect 41 151 42 152 
<< m1 >>
rect 42 151 43 152 
<< m1 >>
rect 43 151 44 152 
<< m2 >>
rect 43 151 44 152 
<< m1 >>
rect 44 151 45 152 
<< m1 >>
rect 45 151 46 152 
<< m2 >>
rect 45 151 46 152 
<< m1 >>
rect 46 151 47 152 
<< m1 >>
rect 47 151 48 152 
<< m2 >>
rect 47 151 48 152 
<< m2c >>
rect 47 151 48 152 
<< m1 >>
rect 47 151 48 152 
<< m2 >>
rect 47 151 48 152 
<< m2 >>
rect 48 151 49 152 
<< m1 >>
rect 49 151 50 152 
<< m2 >>
rect 49 151 50 152 
<< m2 >>
rect 50 151 51 152 
<< m2 >>
rect 51 151 52 152 
<< m2 >>
rect 52 151 53 152 
<< m2 >>
rect 53 151 54 152 
<< m2 >>
rect 54 151 55 152 
<< m2 >>
rect 55 151 56 152 
<< m2 >>
rect 56 151 57 152 
<< m2 >>
rect 57 151 58 152 
<< m2 >>
rect 58 151 59 152 
<< m2 >>
rect 59 151 60 152 
<< m2 >>
rect 60 151 61 152 
<< m2 >>
rect 61 151 62 152 
<< m2 >>
rect 62 151 63 152 
<< m1 >>
rect 66 151 67 152 
<< m2 >>
rect 66 151 67 152 
<< m1 >>
rect 67 151 68 152 
<< m1 >>
rect 68 151 69 152 
<< m1 >>
rect 69 151 70 152 
<< m1 >>
rect 70 151 71 152 
<< m1 >>
rect 71 151 72 152 
<< m1 >>
rect 73 151 74 152 
<< m2 >>
rect 77 151 78 152 
<< m1 >>
rect 79 151 80 152 
<< m1 >>
rect 81 151 82 152 
<< m1 >>
rect 100 151 101 152 
<< m1 >>
rect 102 151 103 152 
<< m2 >>
rect 151 151 152 152 
<< m2 >>
rect 156 151 157 152 
<< m2 >>
rect 157 151 158 152 
<< m1 >>
rect 163 151 164 152 
<< m1 >>
rect 10 152 11 153 
<< m2 >>
rect 10 152 11 153 
<< m1 >>
rect 13 152 14 153 
<< m1 >>
rect 22 152 23 153 
<< m1 >>
rect 25 152 26 153 
<< m1 >>
rect 27 152 28 153 
<< m1 >>
rect 31 152 32 153 
<< m2 >>
rect 34 152 35 153 
<< m2 >>
rect 38 152 39 153 
<< m2 >>
rect 43 152 44 153 
<< m2 >>
rect 45 152 46 153 
<< m1 >>
rect 49 152 50 153 
<< m1 >>
rect 62 152 63 153 
<< m2 >>
rect 62 152 63 153 
<< m2c >>
rect 62 152 63 153 
<< m1 >>
rect 62 152 63 153 
<< m2 >>
rect 62 152 63 153 
<< m1 >>
rect 63 152 64 153 
<< m1 >>
rect 64 152 65 153 
<< m1 >>
rect 65 152 66 153 
<< m1 >>
rect 66 152 67 153 
<< m2 >>
rect 66 152 67 153 
<< m1 >>
rect 71 152 72 153 
<< m2 >>
rect 71 152 72 153 
<< m2c >>
rect 71 152 72 153 
<< m1 >>
rect 71 152 72 153 
<< m2 >>
rect 71 152 72 153 
<< m2 >>
rect 72 152 73 153 
<< m1 >>
rect 73 152 74 153 
<< m2 >>
rect 73 152 74 153 
<< m2 >>
rect 74 152 75 153 
<< m1 >>
rect 75 152 76 153 
<< m2 >>
rect 75 152 76 153 
<< m2c >>
rect 75 152 76 153 
<< m1 >>
rect 75 152 76 153 
<< m2 >>
rect 75 152 76 153 
<< m1 >>
rect 76 152 77 153 
<< m1 >>
rect 77 152 78 153 
<< m2 >>
rect 77 152 78 153 
<< m1 >>
rect 78 152 79 153 
<< m1 >>
rect 79 152 80 153 
<< m1 >>
rect 81 152 82 153 
<< m2 >>
rect 82 152 83 153 
<< m1 >>
rect 83 152 84 153 
<< m2 >>
rect 83 152 84 153 
<< m2c >>
rect 83 152 84 153 
<< m1 >>
rect 83 152 84 153 
<< m2 >>
rect 83 152 84 153 
<< m1 >>
rect 84 152 85 153 
<< m1 >>
rect 85 152 86 153 
<< m1 >>
rect 86 152 87 153 
<< m1 >>
rect 87 152 88 153 
<< m1 >>
rect 88 152 89 153 
<< m1 >>
rect 89 152 90 153 
<< m1 >>
rect 90 152 91 153 
<< m1 >>
rect 91 152 92 153 
<< m1 >>
rect 92 152 93 153 
<< m1 >>
rect 93 152 94 153 
<< m1 >>
rect 94 152 95 153 
<< m1 >>
rect 95 152 96 153 
<< m1 >>
rect 96 152 97 153 
<< m1 >>
rect 97 152 98 153 
<< m1 >>
rect 98 152 99 153 
<< m1 >>
rect 99 152 100 153 
<< m1 >>
rect 100 152 101 153 
<< m1 >>
rect 102 152 103 153 
<< m1 >>
rect 151 152 152 153 
<< m2 >>
rect 151 152 152 153 
<< m2c >>
rect 151 152 152 153 
<< m1 >>
rect 151 152 152 153 
<< m2 >>
rect 151 152 152 153 
<< m1 >>
rect 157 152 158 153 
<< m2 >>
rect 157 152 158 153 
<< m2c >>
rect 157 152 158 153 
<< m1 >>
rect 157 152 158 153 
<< m2 >>
rect 157 152 158 153 
<< m1 >>
rect 163 152 164 153 
<< m1 >>
rect 10 153 11 154 
<< m2 >>
rect 10 153 11 154 
<< m1 >>
rect 13 153 14 154 
<< m1 >>
rect 22 153 23 154 
<< m1 >>
rect 25 153 26 154 
<< m1 >>
rect 27 153 28 154 
<< m1 >>
rect 31 153 32 154 
<< m1 >>
rect 34 153 35 154 
<< m2 >>
rect 34 153 35 154 
<< m2c >>
rect 34 153 35 154 
<< m1 >>
rect 34 153 35 154 
<< m2 >>
rect 34 153 35 154 
<< m1 >>
rect 35 153 36 154 
<< m1 >>
rect 36 153 37 154 
<< m1 >>
rect 37 153 38 154 
<< m2 >>
rect 38 153 39 154 
<< m1 >>
rect 43 153 44 154 
<< m2 >>
rect 43 153 44 154 
<< m2c >>
rect 43 153 44 154 
<< m1 >>
rect 43 153 44 154 
<< m2 >>
rect 43 153 44 154 
<< m1 >>
rect 45 153 46 154 
<< m2 >>
rect 45 153 46 154 
<< m2c >>
rect 45 153 46 154 
<< m1 >>
rect 45 153 46 154 
<< m2 >>
rect 45 153 46 154 
<< m1 >>
rect 49 153 50 154 
<< m2 >>
rect 66 153 67 154 
<< m1 >>
rect 73 153 74 154 
<< m2 >>
rect 77 153 78 154 
<< m1 >>
rect 81 153 82 154 
<< m2 >>
rect 82 153 83 154 
<< m1 >>
rect 102 153 103 154 
<< m1 >>
rect 151 153 152 154 
<< m1 >>
rect 157 153 158 154 
<< m1 >>
rect 163 153 164 154 
<< m1 >>
rect 10 154 11 155 
<< m2 >>
rect 10 154 11 155 
<< m1 >>
rect 13 154 14 155 
<< m1 >>
rect 22 154 23 155 
<< m1 >>
rect 25 154 26 155 
<< m1 >>
rect 27 154 28 155 
<< m1 >>
rect 31 154 32 155 
<< m1 >>
rect 37 154 38 155 
<< m2 >>
rect 38 154 39 155 
<< m1 >>
rect 43 154 44 155 
<< m1 >>
rect 45 154 46 155 
<< m1 >>
rect 49 154 50 155 
<< m1 >>
rect 64 154 65 155 
<< m1 >>
rect 65 154 66 155 
<< m1 >>
rect 66 154 67 155 
<< m2 >>
rect 66 154 67 155 
<< m2c >>
rect 66 154 67 155 
<< m1 >>
rect 66 154 67 155 
<< m2 >>
rect 66 154 67 155 
<< m1 >>
rect 73 154 74 155 
<< m2 >>
rect 74 154 75 155 
<< m1 >>
rect 75 154 76 155 
<< m2 >>
rect 75 154 76 155 
<< m2c >>
rect 75 154 76 155 
<< m1 >>
rect 75 154 76 155 
<< m2 >>
rect 75 154 76 155 
<< m1 >>
rect 76 154 77 155 
<< m1 >>
rect 77 154 78 155 
<< m2 >>
rect 77 154 78 155 
<< m1 >>
rect 78 154 79 155 
<< m1 >>
rect 79 154 80 155 
<< m2 >>
rect 79 154 80 155 
<< m2c >>
rect 79 154 80 155 
<< m1 >>
rect 79 154 80 155 
<< m2 >>
rect 79 154 80 155 
<< m2 >>
rect 80 154 81 155 
<< m1 >>
rect 81 154 82 155 
<< m2 >>
rect 81 154 82 155 
<< m2 >>
rect 82 154 83 155 
<< m1 >>
rect 102 154 103 155 
<< m1 >>
rect 118 154 119 155 
<< m1 >>
rect 119 154 120 155 
<< m1 >>
rect 120 154 121 155 
<< m1 >>
rect 121 154 122 155 
<< m1 >>
rect 124 154 125 155 
<< m1 >>
rect 125 154 126 155 
<< m1 >>
rect 126 154 127 155 
<< m1 >>
rect 127 154 128 155 
<< m1 >>
rect 128 154 129 155 
<< m1 >>
rect 129 154 130 155 
<< m1 >>
rect 130 154 131 155 
<< m1 >>
rect 131 154 132 155 
<< m1 >>
rect 132 154 133 155 
<< m1 >>
rect 133 154 134 155 
<< m1 >>
rect 134 154 135 155 
<< m1 >>
rect 135 154 136 155 
<< m1 >>
rect 136 154 137 155 
<< m1 >>
rect 137 154 138 155 
<< m1 >>
rect 138 154 139 155 
<< m1 >>
rect 139 154 140 155 
<< m1 >>
rect 140 154 141 155 
<< m1 >>
rect 141 154 142 155 
<< m1 >>
rect 142 154 143 155 
<< m1 >>
rect 151 154 152 155 
<< m1 >>
rect 157 154 158 155 
<< m1 >>
rect 163 154 164 155 
<< m1 >>
rect 10 155 11 156 
<< m2 >>
rect 10 155 11 156 
<< m1 >>
rect 13 155 14 156 
<< m1 >>
rect 22 155 23 156 
<< m1 >>
rect 25 155 26 156 
<< m1 >>
rect 27 155 28 156 
<< m1 >>
rect 31 155 32 156 
<< m1 >>
rect 37 155 38 156 
<< m2 >>
rect 38 155 39 156 
<< m1 >>
rect 43 155 44 156 
<< m1 >>
rect 45 155 46 156 
<< m1 >>
rect 49 155 50 156 
<< m1 >>
rect 64 155 65 156 
<< m1 >>
rect 73 155 74 156 
<< m2 >>
rect 74 155 75 156 
<< m2 >>
rect 77 155 78 156 
<< m1 >>
rect 81 155 82 156 
<< m1 >>
rect 102 155 103 156 
<< m1 >>
rect 118 155 119 156 
<< m1 >>
rect 121 155 122 156 
<< m1 >>
rect 124 155 125 156 
<< m1 >>
rect 142 155 143 156 
<< m1 >>
rect 151 155 152 156 
<< m1 >>
rect 157 155 158 156 
<< m1 >>
rect 163 155 164 156 
<< m1 >>
rect 10 156 11 157 
<< m2 >>
rect 10 156 11 157 
<< pdiffusion >>
rect 12 156 13 157 
<< m1 >>
rect 13 156 14 157 
<< pdiffusion >>
rect 13 156 14 157 
<< pdiffusion >>
rect 14 156 15 157 
<< pdiffusion >>
rect 15 156 16 157 
<< pdiffusion >>
rect 16 156 17 157 
<< pdiffusion >>
rect 17 156 18 157 
<< m1 >>
rect 22 156 23 157 
<< m1 >>
rect 25 156 26 157 
<< m1 >>
rect 27 156 28 157 
<< pdiffusion >>
rect 30 156 31 157 
<< m1 >>
rect 31 156 32 157 
<< pdiffusion >>
rect 31 156 32 157 
<< pdiffusion >>
rect 32 156 33 157 
<< pdiffusion >>
rect 33 156 34 157 
<< pdiffusion >>
rect 34 156 35 157 
<< pdiffusion >>
rect 35 156 36 157 
<< m1 >>
rect 37 156 38 157 
<< m2 >>
rect 38 156 39 157 
<< m1 >>
rect 43 156 44 157 
<< m1 >>
rect 45 156 46 157 
<< pdiffusion >>
rect 48 156 49 157 
<< m1 >>
rect 49 156 50 157 
<< pdiffusion >>
rect 49 156 50 157 
<< pdiffusion >>
rect 50 156 51 157 
<< pdiffusion >>
rect 51 156 52 157 
<< pdiffusion >>
rect 52 156 53 157 
<< pdiffusion >>
rect 53 156 54 157 
<< m1 >>
rect 64 156 65 157 
<< pdiffusion >>
rect 66 156 67 157 
<< pdiffusion >>
rect 67 156 68 157 
<< pdiffusion >>
rect 68 156 69 157 
<< pdiffusion >>
rect 69 156 70 157 
<< pdiffusion >>
rect 70 156 71 157 
<< pdiffusion >>
rect 71 156 72 157 
<< m1 >>
rect 73 156 74 157 
<< m2 >>
rect 74 156 75 157 
<< m1 >>
rect 77 156 78 157 
<< m2 >>
rect 77 156 78 157 
<< m2c >>
rect 77 156 78 157 
<< m1 >>
rect 77 156 78 157 
<< m2 >>
rect 77 156 78 157 
<< m1 >>
rect 81 156 82 157 
<< m1 >>
rect 102 156 103 157 
<< m1 >>
rect 118 156 119 157 
<< pdiffusion >>
rect 120 156 121 157 
<< m1 >>
rect 121 156 122 157 
<< pdiffusion >>
rect 121 156 122 157 
<< pdiffusion >>
rect 122 156 123 157 
<< pdiffusion >>
rect 123 156 124 157 
<< m1 >>
rect 124 156 125 157 
<< pdiffusion >>
rect 124 156 125 157 
<< pdiffusion >>
rect 125 156 126 157 
<< m1 >>
rect 142 156 143 157 
<< m1 >>
rect 151 156 152 157 
<< pdiffusion >>
rect 156 156 157 157 
<< m1 >>
rect 157 156 158 157 
<< pdiffusion >>
rect 157 156 158 157 
<< pdiffusion >>
rect 158 156 159 157 
<< pdiffusion >>
rect 159 156 160 157 
<< pdiffusion >>
rect 160 156 161 157 
<< pdiffusion >>
rect 161 156 162 157 
<< m1 >>
rect 163 156 164 157 
<< pdiffusion >>
rect 174 156 175 157 
<< pdiffusion >>
rect 175 156 176 157 
<< pdiffusion >>
rect 176 156 177 157 
<< pdiffusion >>
rect 177 156 178 157 
<< pdiffusion >>
rect 178 156 179 157 
<< pdiffusion >>
rect 179 156 180 157 
<< m1 >>
rect 10 157 11 158 
<< m2 >>
rect 10 157 11 158 
<< pdiffusion >>
rect 12 157 13 158 
<< pdiffusion >>
rect 13 157 14 158 
<< pdiffusion >>
rect 14 157 15 158 
<< pdiffusion >>
rect 15 157 16 158 
<< pdiffusion >>
rect 16 157 17 158 
<< pdiffusion >>
rect 17 157 18 158 
<< m1 >>
rect 22 157 23 158 
<< m1 >>
rect 25 157 26 158 
<< m1 >>
rect 27 157 28 158 
<< pdiffusion >>
rect 30 157 31 158 
<< pdiffusion >>
rect 31 157 32 158 
<< pdiffusion >>
rect 32 157 33 158 
<< pdiffusion >>
rect 33 157 34 158 
<< pdiffusion >>
rect 34 157 35 158 
<< pdiffusion >>
rect 35 157 36 158 
<< m1 >>
rect 37 157 38 158 
<< m2 >>
rect 38 157 39 158 
<< m1 >>
rect 43 157 44 158 
<< m1 >>
rect 45 157 46 158 
<< pdiffusion >>
rect 48 157 49 158 
<< pdiffusion >>
rect 49 157 50 158 
<< pdiffusion >>
rect 50 157 51 158 
<< pdiffusion >>
rect 51 157 52 158 
<< pdiffusion >>
rect 52 157 53 158 
<< pdiffusion >>
rect 53 157 54 158 
<< m1 >>
rect 64 157 65 158 
<< pdiffusion >>
rect 66 157 67 158 
<< pdiffusion >>
rect 67 157 68 158 
<< pdiffusion >>
rect 68 157 69 158 
<< pdiffusion >>
rect 69 157 70 158 
<< pdiffusion >>
rect 70 157 71 158 
<< pdiffusion >>
rect 71 157 72 158 
<< m1 >>
rect 73 157 74 158 
<< m2 >>
rect 74 157 75 158 
<< m1 >>
rect 77 157 78 158 
<< m1 >>
rect 81 157 82 158 
<< m1 >>
rect 102 157 103 158 
<< m1 >>
rect 118 157 119 158 
<< pdiffusion >>
rect 120 157 121 158 
<< pdiffusion >>
rect 121 157 122 158 
<< pdiffusion >>
rect 122 157 123 158 
<< pdiffusion >>
rect 123 157 124 158 
<< pdiffusion >>
rect 124 157 125 158 
<< pdiffusion >>
rect 125 157 126 158 
<< m1 >>
rect 142 157 143 158 
<< m1 >>
rect 151 157 152 158 
<< pdiffusion >>
rect 156 157 157 158 
<< pdiffusion >>
rect 157 157 158 158 
<< pdiffusion >>
rect 158 157 159 158 
<< pdiffusion >>
rect 159 157 160 158 
<< pdiffusion >>
rect 160 157 161 158 
<< pdiffusion >>
rect 161 157 162 158 
<< m1 >>
rect 163 157 164 158 
<< pdiffusion >>
rect 174 157 175 158 
<< pdiffusion >>
rect 175 157 176 158 
<< pdiffusion >>
rect 176 157 177 158 
<< pdiffusion >>
rect 177 157 178 158 
<< pdiffusion >>
rect 178 157 179 158 
<< pdiffusion >>
rect 179 157 180 158 
<< m1 >>
rect 10 158 11 159 
<< m2 >>
rect 10 158 11 159 
<< pdiffusion >>
rect 12 158 13 159 
<< pdiffusion >>
rect 13 158 14 159 
<< pdiffusion >>
rect 14 158 15 159 
<< pdiffusion >>
rect 15 158 16 159 
<< pdiffusion >>
rect 16 158 17 159 
<< pdiffusion >>
rect 17 158 18 159 
<< m1 >>
rect 22 158 23 159 
<< m1 >>
rect 25 158 26 159 
<< m1 >>
rect 27 158 28 159 
<< pdiffusion >>
rect 30 158 31 159 
<< pdiffusion >>
rect 31 158 32 159 
<< pdiffusion >>
rect 32 158 33 159 
<< pdiffusion >>
rect 33 158 34 159 
<< pdiffusion >>
rect 34 158 35 159 
<< pdiffusion >>
rect 35 158 36 159 
<< m1 >>
rect 37 158 38 159 
<< m2 >>
rect 38 158 39 159 
<< m1 >>
rect 43 158 44 159 
<< m1 >>
rect 45 158 46 159 
<< pdiffusion >>
rect 48 158 49 159 
<< pdiffusion >>
rect 49 158 50 159 
<< pdiffusion >>
rect 50 158 51 159 
<< pdiffusion >>
rect 51 158 52 159 
<< pdiffusion >>
rect 52 158 53 159 
<< pdiffusion >>
rect 53 158 54 159 
<< m1 >>
rect 64 158 65 159 
<< pdiffusion >>
rect 66 158 67 159 
<< pdiffusion >>
rect 67 158 68 159 
<< pdiffusion >>
rect 68 158 69 159 
<< pdiffusion >>
rect 69 158 70 159 
<< pdiffusion >>
rect 70 158 71 159 
<< pdiffusion >>
rect 71 158 72 159 
<< m1 >>
rect 73 158 74 159 
<< m2 >>
rect 74 158 75 159 
<< m1 >>
rect 77 158 78 159 
<< m1 >>
rect 81 158 82 159 
<< m1 >>
rect 102 158 103 159 
<< m1 >>
rect 118 158 119 159 
<< pdiffusion >>
rect 120 158 121 159 
<< pdiffusion >>
rect 121 158 122 159 
<< pdiffusion >>
rect 122 158 123 159 
<< pdiffusion >>
rect 123 158 124 159 
<< pdiffusion >>
rect 124 158 125 159 
<< pdiffusion >>
rect 125 158 126 159 
<< m1 >>
rect 142 158 143 159 
<< m1 >>
rect 151 158 152 159 
<< pdiffusion >>
rect 156 158 157 159 
<< pdiffusion >>
rect 157 158 158 159 
<< pdiffusion >>
rect 158 158 159 159 
<< pdiffusion >>
rect 159 158 160 159 
<< pdiffusion >>
rect 160 158 161 159 
<< pdiffusion >>
rect 161 158 162 159 
<< m1 >>
rect 163 158 164 159 
<< pdiffusion >>
rect 174 158 175 159 
<< pdiffusion >>
rect 175 158 176 159 
<< pdiffusion >>
rect 176 158 177 159 
<< pdiffusion >>
rect 177 158 178 159 
<< pdiffusion >>
rect 178 158 179 159 
<< pdiffusion >>
rect 179 158 180 159 
<< m1 >>
rect 10 159 11 160 
<< m2 >>
rect 10 159 11 160 
<< pdiffusion >>
rect 12 159 13 160 
<< pdiffusion >>
rect 13 159 14 160 
<< pdiffusion >>
rect 14 159 15 160 
<< pdiffusion >>
rect 15 159 16 160 
<< pdiffusion >>
rect 16 159 17 160 
<< pdiffusion >>
rect 17 159 18 160 
<< m1 >>
rect 22 159 23 160 
<< m1 >>
rect 25 159 26 160 
<< m1 >>
rect 27 159 28 160 
<< pdiffusion >>
rect 30 159 31 160 
<< pdiffusion >>
rect 31 159 32 160 
<< pdiffusion >>
rect 32 159 33 160 
<< pdiffusion >>
rect 33 159 34 160 
<< pdiffusion >>
rect 34 159 35 160 
<< pdiffusion >>
rect 35 159 36 160 
<< m1 >>
rect 37 159 38 160 
<< m2 >>
rect 38 159 39 160 
<< m1 >>
rect 43 159 44 160 
<< m1 >>
rect 45 159 46 160 
<< pdiffusion >>
rect 48 159 49 160 
<< pdiffusion >>
rect 49 159 50 160 
<< pdiffusion >>
rect 50 159 51 160 
<< pdiffusion >>
rect 51 159 52 160 
<< pdiffusion >>
rect 52 159 53 160 
<< pdiffusion >>
rect 53 159 54 160 
<< m1 >>
rect 64 159 65 160 
<< pdiffusion >>
rect 66 159 67 160 
<< pdiffusion >>
rect 67 159 68 160 
<< pdiffusion >>
rect 68 159 69 160 
<< pdiffusion >>
rect 69 159 70 160 
<< pdiffusion >>
rect 70 159 71 160 
<< pdiffusion >>
rect 71 159 72 160 
<< m1 >>
rect 73 159 74 160 
<< m2 >>
rect 74 159 75 160 
<< m1 >>
rect 77 159 78 160 
<< m1 >>
rect 81 159 82 160 
<< m1 >>
rect 102 159 103 160 
<< m1 >>
rect 118 159 119 160 
<< pdiffusion >>
rect 120 159 121 160 
<< pdiffusion >>
rect 121 159 122 160 
<< pdiffusion >>
rect 122 159 123 160 
<< pdiffusion >>
rect 123 159 124 160 
<< pdiffusion >>
rect 124 159 125 160 
<< pdiffusion >>
rect 125 159 126 160 
<< m1 >>
rect 142 159 143 160 
<< m1 >>
rect 151 159 152 160 
<< pdiffusion >>
rect 156 159 157 160 
<< pdiffusion >>
rect 157 159 158 160 
<< pdiffusion >>
rect 158 159 159 160 
<< pdiffusion >>
rect 159 159 160 160 
<< pdiffusion >>
rect 160 159 161 160 
<< pdiffusion >>
rect 161 159 162 160 
<< m1 >>
rect 163 159 164 160 
<< pdiffusion >>
rect 174 159 175 160 
<< pdiffusion >>
rect 175 159 176 160 
<< pdiffusion >>
rect 176 159 177 160 
<< pdiffusion >>
rect 177 159 178 160 
<< pdiffusion >>
rect 178 159 179 160 
<< pdiffusion >>
rect 179 159 180 160 
<< m1 >>
rect 10 160 11 161 
<< m2 >>
rect 10 160 11 161 
<< pdiffusion >>
rect 12 160 13 161 
<< pdiffusion >>
rect 13 160 14 161 
<< pdiffusion >>
rect 14 160 15 161 
<< pdiffusion >>
rect 15 160 16 161 
<< pdiffusion >>
rect 16 160 17 161 
<< pdiffusion >>
rect 17 160 18 161 
<< m1 >>
rect 22 160 23 161 
<< m1 >>
rect 25 160 26 161 
<< m1 >>
rect 27 160 28 161 
<< pdiffusion >>
rect 30 160 31 161 
<< pdiffusion >>
rect 31 160 32 161 
<< pdiffusion >>
rect 32 160 33 161 
<< pdiffusion >>
rect 33 160 34 161 
<< pdiffusion >>
rect 34 160 35 161 
<< pdiffusion >>
rect 35 160 36 161 
<< m1 >>
rect 37 160 38 161 
<< m2 >>
rect 38 160 39 161 
<< m1 >>
rect 43 160 44 161 
<< m1 >>
rect 45 160 46 161 
<< pdiffusion >>
rect 48 160 49 161 
<< pdiffusion >>
rect 49 160 50 161 
<< pdiffusion >>
rect 50 160 51 161 
<< pdiffusion >>
rect 51 160 52 161 
<< pdiffusion >>
rect 52 160 53 161 
<< pdiffusion >>
rect 53 160 54 161 
<< m1 >>
rect 64 160 65 161 
<< pdiffusion >>
rect 66 160 67 161 
<< pdiffusion >>
rect 67 160 68 161 
<< pdiffusion >>
rect 68 160 69 161 
<< pdiffusion >>
rect 69 160 70 161 
<< pdiffusion >>
rect 70 160 71 161 
<< pdiffusion >>
rect 71 160 72 161 
<< m1 >>
rect 73 160 74 161 
<< m2 >>
rect 74 160 75 161 
<< m1 >>
rect 77 160 78 161 
<< m1 >>
rect 81 160 82 161 
<< m1 >>
rect 102 160 103 161 
<< m1 >>
rect 118 160 119 161 
<< pdiffusion >>
rect 120 160 121 161 
<< pdiffusion >>
rect 121 160 122 161 
<< pdiffusion >>
rect 122 160 123 161 
<< pdiffusion >>
rect 123 160 124 161 
<< pdiffusion >>
rect 124 160 125 161 
<< pdiffusion >>
rect 125 160 126 161 
<< m1 >>
rect 142 160 143 161 
<< m1 >>
rect 151 160 152 161 
<< pdiffusion >>
rect 156 160 157 161 
<< pdiffusion >>
rect 157 160 158 161 
<< pdiffusion >>
rect 158 160 159 161 
<< pdiffusion >>
rect 159 160 160 161 
<< pdiffusion >>
rect 160 160 161 161 
<< pdiffusion >>
rect 161 160 162 161 
<< m1 >>
rect 163 160 164 161 
<< pdiffusion >>
rect 174 160 175 161 
<< pdiffusion >>
rect 175 160 176 161 
<< pdiffusion >>
rect 176 160 177 161 
<< pdiffusion >>
rect 177 160 178 161 
<< pdiffusion >>
rect 178 160 179 161 
<< pdiffusion >>
rect 179 160 180 161 
<< m1 >>
rect 10 161 11 162 
<< m2 >>
rect 10 161 11 162 
<< pdiffusion >>
rect 12 161 13 162 
<< m1 >>
rect 13 161 14 162 
<< pdiffusion >>
rect 13 161 14 162 
<< pdiffusion >>
rect 14 161 15 162 
<< pdiffusion >>
rect 15 161 16 162 
<< m1 >>
rect 16 161 17 162 
<< pdiffusion >>
rect 16 161 17 162 
<< pdiffusion >>
rect 17 161 18 162 
<< m1 >>
rect 22 161 23 162 
<< m2 >>
rect 22 161 23 162 
<< m2c >>
rect 22 161 23 162 
<< m1 >>
rect 22 161 23 162 
<< m2 >>
rect 22 161 23 162 
<< m1 >>
rect 25 161 26 162 
<< m2 >>
rect 25 161 26 162 
<< m2c >>
rect 25 161 26 162 
<< m1 >>
rect 25 161 26 162 
<< m2 >>
rect 25 161 26 162 
<< m2 >>
rect 26 161 27 162 
<< m1 >>
rect 27 161 28 162 
<< m2 >>
rect 27 161 28 162 
<< m2 >>
rect 28 161 29 162 
<< pdiffusion >>
rect 30 161 31 162 
<< pdiffusion >>
rect 31 161 32 162 
<< pdiffusion >>
rect 32 161 33 162 
<< pdiffusion >>
rect 33 161 34 162 
<< pdiffusion >>
rect 34 161 35 162 
<< pdiffusion >>
rect 35 161 36 162 
<< m1 >>
rect 37 161 38 162 
<< m2 >>
rect 38 161 39 162 
<< m1 >>
rect 43 161 44 162 
<< m1 >>
rect 45 161 46 162 
<< pdiffusion >>
rect 48 161 49 162 
<< pdiffusion >>
rect 49 161 50 162 
<< pdiffusion >>
rect 50 161 51 162 
<< pdiffusion >>
rect 51 161 52 162 
<< pdiffusion >>
rect 52 161 53 162 
<< pdiffusion >>
rect 53 161 54 162 
<< m1 >>
rect 64 161 65 162 
<< pdiffusion >>
rect 66 161 67 162 
<< pdiffusion >>
rect 67 161 68 162 
<< pdiffusion >>
rect 68 161 69 162 
<< pdiffusion >>
rect 69 161 70 162 
<< pdiffusion >>
rect 70 161 71 162 
<< pdiffusion >>
rect 71 161 72 162 
<< m1 >>
rect 73 161 74 162 
<< m2 >>
rect 74 161 75 162 
<< m1 >>
rect 77 161 78 162 
<< m1 >>
rect 81 161 82 162 
<< m1 >>
rect 102 161 103 162 
<< m1 >>
rect 118 161 119 162 
<< pdiffusion >>
rect 120 161 121 162 
<< pdiffusion >>
rect 121 161 122 162 
<< pdiffusion >>
rect 122 161 123 162 
<< pdiffusion >>
rect 123 161 124 162 
<< pdiffusion >>
rect 124 161 125 162 
<< pdiffusion >>
rect 125 161 126 162 
<< m1 >>
rect 142 161 143 162 
<< m1 >>
rect 151 161 152 162 
<< pdiffusion >>
rect 156 161 157 162 
<< pdiffusion >>
rect 157 161 158 162 
<< pdiffusion >>
rect 158 161 159 162 
<< pdiffusion >>
rect 159 161 160 162 
<< pdiffusion >>
rect 160 161 161 162 
<< pdiffusion >>
rect 161 161 162 162 
<< m1 >>
rect 163 161 164 162 
<< pdiffusion >>
rect 174 161 175 162 
<< m1 >>
rect 175 161 176 162 
<< pdiffusion >>
rect 175 161 176 162 
<< pdiffusion >>
rect 176 161 177 162 
<< pdiffusion >>
rect 177 161 178 162 
<< pdiffusion >>
rect 178 161 179 162 
<< pdiffusion >>
rect 179 161 180 162 
<< m1 >>
rect 10 162 11 163 
<< m2 >>
rect 10 162 11 163 
<< m1 >>
rect 13 162 14 163 
<< m1 >>
rect 16 162 17 163 
<< m2 >>
rect 22 162 23 163 
<< m1 >>
rect 27 162 28 163 
<< m2 >>
rect 28 162 29 163 
<< m1 >>
rect 37 162 38 163 
<< m2 >>
rect 38 162 39 163 
<< m1 >>
rect 43 162 44 163 
<< m1 >>
rect 45 162 46 163 
<< m1 >>
rect 64 162 65 163 
<< m1 >>
rect 73 162 74 163 
<< m2 >>
rect 74 162 75 163 
<< m1 >>
rect 77 162 78 163 
<< m1 >>
rect 81 162 82 163 
<< m1 >>
rect 102 162 103 163 
<< m1 >>
rect 118 162 119 163 
<< m1 >>
rect 142 162 143 163 
<< m1 >>
rect 151 162 152 163 
<< m1 >>
rect 163 162 164 163 
<< m1 >>
rect 175 162 176 163 
<< m1 >>
rect 10 163 11 164 
<< m2 >>
rect 10 163 11 164 
<< m1 >>
rect 13 163 14 164 
<< m1 >>
rect 16 163 17 164 
<< m1 >>
rect 17 163 18 164 
<< m1 >>
rect 18 163 19 164 
<< m1 >>
rect 19 163 20 164 
<< m1 >>
rect 20 163 21 164 
<< m1 >>
rect 21 163 22 164 
<< m1 >>
rect 22 163 23 164 
<< m2 >>
rect 22 163 23 164 
<< m1 >>
rect 23 163 24 164 
<< m1 >>
rect 24 163 25 164 
<< m1 >>
rect 25 163 26 164 
<< m1 >>
rect 26 163 27 164 
<< m1 >>
rect 27 163 28 164 
<< m2 >>
rect 28 163 29 164 
<< m1 >>
rect 37 163 38 164 
<< m2 >>
rect 38 163 39 164 
<< m1 >>
rect 43 163 44 164 
<< m1 >>
rect 45 163 46 164 
<< m1 >>
rect 64 163 65 164 
<< m1 >>
rect 71 163 72 164 
<< m2 >>
rect 71 163 72 164 
<< m2c >>
rect 71 163 72 164 
<< m1 >>
rect 71 163 72 164 
<< m2 >>
rect 71 163 72 164 
<< m2 >>
rect 72 163 73 164 
<< m1 >>
rect 73 163 74 164 
<< m2 >>
rect 73 163 74 164 
<< m2 >>
rect 74 163 75 164 
<< m1 >>
rect 77 163 78 164 
<< m1 >>
rect 81 163 82 164 
<< m1 >>
rect 102 163 103 164 
<< m1 >>
rect 118 163 119 164 
<< m1 >>
rect 142 163 143 164 
<< m1 >>
rect 151 163 152 164 
<< m1 >>
rect 163 163 164 164 
<< m1 >>
rect 164 163 165 164 
<< m1 >>
rect 165 163 166 164 
<< m1 >>
rect 166 163 167 164 
<< m1 >>
rect 167 163 168 164 
<< m1 >>
rect 168 163 169 164 
<< m1 >>
rect 169 163 170 164 
<< m1 >>
rect 170 163 171 164 
<< m1 >>
rect 171 163 172 164 
<< m1 >>
rect 172 163 173 164 
<< m1 >>
rect 173 163 174 164 
<< m1 >>
rect 174 163 175 164 
<< m1 >>
rect 175 163 176 164 
<< m1 >>
rect 10 164 11 165 
<< m2 >>
rect 10 164 11 165 
<< m1 >>
rect 13 164 14 165 
<< m2 >>
rect 22 164 23 165 
<< m2 >>
rect 28 164 29 165 
<< m1 >>
rect 37 164 38 165 
<< m2 >>
rect 38 164 39 165 
<< m1 >>
rect 43 164 44 165 
<< m1 >>
rect 45 164 46 165 
<< m1 >>
rect 64 164 65 165 
<< m1 >>
rect 69 164 70 165 
<< m2 >>
rect 69 164 70 165 
<< m2c >>
rect 69 164 70 165 
<< m1 >>
rect 69 164 70 165 
<< m2 >>
rect 69 164 70 165 
<< m1 >>
rect 70 164 71 165 
<< m1 >>
rect 71 164 72 165 
<< m1 >>
rect 73 164 74 165 
<< m1 >>
rect 77 164 78 165 
<< m2 >>
rect 77 164 78 165 
<< m2c >>
rect 77 164 78 165 
<< m1 >>
rect 77 164 78 165 
<< m2 >>
rect 77 164 78 165 
<< m1 >>
rect 81 164 82 165 
<< m1 >>
rect 102 164 103 165 
<< m1 >>
rect 118 164 119 165 
<< m1 >>
rect 142 164 143 165 
<< m1 >>
rect 151 164 152 165 
<< m1 >>
rect 10 165 11 166 
<< m2 >>
rect 10 165 11 166 
<< m1 >>
rect 13 165 14 166 
<< m1 >>
rect 22 165 23 166 
<< m2 >>
rect 22 165 23 166 
<< m2c >>
rect 22 165 23 166 
<< m1 >>
rect 22 165 23 166 
<< m2 >>
rect 22 165 23 166 
<< m1 >>
rect 28 165 29 166 
<< m2 >>
rect 28 165 29 166 
<< m2c >>
rect 28 165 29 166 
<< m1 >>
rect 28 165 29 166 
<< m2 >>
rect 28 165 29 166 
<< m1 >>
rect 37 165 38 166 
<< m2 >>
rect 38 165 39 166 
<< m1 >>
rect 43 165 44 166 
<< m1 >>
rect 45 165 46 166 
<< m1 >>
rect 64 165 65 166 
<< m2 >>
rect 69 165 70 166 
<< m1 >>
rect 73 165 74 166 
<< m2 >>
rect 77 165 78 166 
<< m1 >>
rect 81 165 82 166 
<< m1 >>
rect 102 165 103 166 
<< m1 >>
rect 118 165 119 166 
<< m1 >>
rect 142 165 143 166 
<< m1 >>
rect 151 165 152 166 
<< m1 >>
rect 10 166 11 167 
<< m2 >>
rect 10 166 11 167 
<< m1 >>
rect 13 166 14 167 
<< m1 >>
rect 22 166 23 167 
<< m1 >>
rect 28 166 29 167 
<< m1 >>
rect 37 166 38 167 
<< m2 >>
rect 38 166 39 167 
<< m1 >>
rect 43 166 44 167 
<< m1 >>
rect 45 166 46 167 
<< m1 >>
rect 46 166 47 167 
<< m1 >>
rect 47 166 48 167 
<< m1 >>
rect 48 166 49 167 
<< m1 >>
rect 49 166 50 167 
<< m1 >>
rect 50 166 51 167 
<< m1 >>
rect 51 166 52 167 
<< m1 >>
rect 52 166 53 167 
<< m1 >>
rect 53 166 54 167 
<< m1 >>
rect 54 166 55 167 
<< m1 >>
rect 55 166 56 167 
<< m1 >>
rect 56 166 57 167 
<< m1 >>
rect 57 166 58 167 
<< m1 >>
rect 58 166 59 167 
<< m1 >>
rect 59 166 60 167 
<< m1 >>
rect 60 166 61 167 
<< m1 >>
rect 61 166 62 167 
<< m1 >>
rect 62 166 63 167 
<< m2 >>
rect 62 166 63 167 
<< m2c >>
rect 62 166 63 167 
<< m1 >>
rect 62 166 63 167 
<< m2 >>
rect 62 166 63 167 
<< m2 >>
rect 63 166 64 167 
<< m1 >>
rect 64 166 65 167 
<< m2 >>
rect 64 166 65 167 
<< m1 >>
rect 65 166 66 167 
<< m2 >>
rect 65 166 66 167 
<< m1 >>
rect 66 166 67 167 
<< m2 >>
rect 66 166 67 167 
<< m1 >>
rect 67 166 68 167 
<< m2 >>
rect 67 166 68 167 
<< m1 >>
rect 68 166 69 167 
<< m2 >>
rect 68 166 69 167 
<< m1 >>
rect 69 166 70 167 
<< m2 >>
rect 69 166 70 167 
<< m1 >>
rect 70 166 71 167 
<< m1 >>
rect 71 166 72 167 
<< m2 >>
rect 71 166 72 167 
<< m2c >>
rect 71 166 72 167 
<< m1 >>
rect 71 166 72 167 
<< m2 >>
rect 71 166 72 167 
<< m2 >>
rect 72 166 73 167 
<< m1 >>
rect 73 166 74 167 
<< m2 >>
rect 73 166 74 167 
<< m2 >>
rect 74 166 75 167 
<< m1 >>
rect 75 166 76 167 
<< m2 >>
rect 75 166 76 167 
<< m2c >>
rect 75 166 76 167 
<< m1 >>
rect 75 166 76 167 
<< m2 >>
rect 75 166 76 167 
<< m1 >>
rect 76 166 77 167 
<< m1 >>
rect 77 166 78 167 
<< m2 >>
rect 77 166 78 167 
<< m1 >>
rect 78 166 79 167 
<< m1 >>
rect 79 166 80 167 
<< m1 >>
rect 80 166 81 167 
<< m1 >>
rect 81 166 82 167 
<< m1 >>
rect 102 166 103 167 
<< m1 >>
rect 118 166 119 167 
<< m1 >>
rect 142 166 143 167 
<< m1 >>
rect 151 166 152 167 
<< m1 >>
rect 10 167 11 168 
<< m2 >>
rect 10 167 11 168 
<< m1 >>
rect 13 167 14 168 
<< m1 >>
rect 22 167 23 168 
<< m2 >>
rect 22 167 23 168 
<< m2c >>
rect 22 167 23 168 
<< m1 >>
rect 22 167 23 168 
<< m2 >>
rect 22 167 23 168 
<< m1 >>
rect 28 167 29 168 
<< m2 >>
rect 28 167 29 168 
<< m2c >>
rect 28 167 29 168 
<< m1 >>
rect 28 167 29 168 
<< m2 >>
rect 28 167 29 168 
<< m1 >>
rect 37 167 38 168 
<< m2 >>
rect 38 167 39 168 
<< m1 >>
rect 43 167 44 168 
<< m1 >>
rect 73 167 74 168 
<< m2 >>
rect 77 167 78 168 
<< m1 >>
rect 102 167 103 168 
<< m1 >>
rect 118 167 119 168 
<< m1 >>
rect 142 167 143 168 
<< m1 >>
rect 151 167 152 168 
<< m1 >>
rect 10 168 11 169 
<< m2 >>
rect 10 168 11 169 
<< m1 >>
rect 13 168 14 169 
<< m2 >>
rect 22 168 23 169 
<< m2 >>
rect 28 168 29 169 
<< m1 >>
rect 37 168 38 169 
<< m2 >>
rect 38 168 39 169 
<< m1 >>
rect 43 168 44 169 
<< m1 >>
rect 44 168 45 169 
<< m1 >>
rect 45 168 46 169 
<< m1 >>
rect 46 168 47 169 
<< m1 >>
rect 47 168 48 169 
<< m1 >>
rect 48 168 49 169 
<< m1 >>
rect 49 168 50 169 
<< m1 >>
rect 50 168 51 169 
<< m1 >>
rect 51 168 52 169 
<< m1 >>
rect 52 168 53 169 
<< m1 >>
rect 53 168 54 169 
<< m1 >>
rect 54 168 55 169 
<< m1 >>
rect 55 168 56 169 
<< m1 >>
rect 56 168 57 169 
<< m1 >>
rect 57 168 58 169 
<< m1 >>
rect 58 168 59 169 
<< m1 >>
rect 59 168 60 169 
<< m1 >>
rect 60 168 61 169 
<< m1 >>
rect 61 168 62 169 
<< m1 >>
rect 62 168 63 169 
<< m1 >>
rect 63 168 64 169 
<< m1 >>
rect 64 168 65 169 
<< m1 >>
rect 65 168 66 169 
<< m1 >>
rect 66 168 67 169 
<< m1 >>
rect 67 168 68 169 
<< m1 >>
rect 68 168 69 169 
<< m1 >>
rect 69 168 70 169 
<< m1 >>
rect 70 168 71 169 
<< m1 >>
rect 71 168 72 169 
<< m2 >>
rect 71 168 72 169 
<< m2c >>
rect 71 168 72 169 
<< m1 >>
rect 71 168 72 169 
<< m2 >>
rect 71 168 72 169 
<< m2 >>
rect 72 168 73 169 
<< m1 >>
rect 73 168 74 169 
<< m2 >>
rect 73 168 74 169 
<< m2 >>
rect 74 168 75 169 
<< m1 >>
rect 75 168 76 169 
<< m2 >>
rect 75 168 76 169 
<< m2c >>
rect 75 168 76 169 
<< m1 >>
rect 75 168 76 169 
<< m2 >>
rect 75 168 76 169 
<< m1 >>
rect 76 168 77 169 
<< m1 >>
rect 77 168 78 169 
<< m2 >>
rect 77 168 78 169 
<< m1 >>
rect 78 168 79 169 
<< m1 >>
rect 79 168 80 169 
<< m1 >>
rect 80 168 81 169 
<< m1 >>
rect 81 168 82 169 
<< m1 >>
rect 82 168 83 169 
<< m1 >>
rect 83 168 84 169 
<< m1 >>
rect 84 168 85 169 
<< m1 >>
rect 85 168 86 169 
<< m1 >>
rect 86 168 87 169 
<< m1 >>
rect 87 168 88 169 
<< m1 >>
rect 88 168 89 169 
<< m1 >>
rect 89 168 90 169 
<< m1 >>
rect 90 168 91 169 
<< m1 >>
rect 91 168 92 169 
<< m1 >>
rect 92 168 93 169 
<< m1 >>
rect 93 168 94 169 
<< m1 >>
rect 94 168 95 169 
<< m1 >>
rect 95 168 96 169 
<< m1 >>
rect 96 168 97 169 
<< m1 >>
rect 97 168 98 169 
<< m1 >>
rect 98 168 99 169 
<< m1 >>
rect 99 168 100 169 
<< m1 >>
rect 100 168 101 169 
<< m1 >>
rect 101 168 102 169 
<< m1 >>
rect 102 168 103 169 
<< m1 >>
rect 118 168 119 169 
<< m1 >>
rect 142 168 143 169 
<< m1 >>
rect 151 168 152 169 
<< m1 >>
rect 10 169 11 170 
<< m2 >>
rect 10 169 11 170 
<< m1 >>
rect 13 169 14 170 
<< m1 >>
rect 14 169 15 170 
<< m1 >>
rect 15 169 16 170 
<< m1 >>
rect 16 169 17 170 
<< m1 >>
rect 17 169 18 170 
<< m1 >>
rect 18 169 19 170 
<< m1 >>
rect 19 169 20 170 
<< m1 >>
rect 20 169 21 170 
<< m1 >>
rect 21 169 22 170 
<< m1 >>
rect 22 169 23 170 
<< m2 >>
rect 22 169 23 170 
<< m1 >>
rect 23 169 24 170 
<< m1 >>
rect 24 169 25 170 
<< m1 >>
rect 25 169 26 170 
<< m1 >>
rect 26 169 27 170 
<< m1 >>
rect 27 169 28 170 
<< m1 >>
rect 28 169 29 170 
<< m2 >>
rect 28 169 29 170 
<< m1 >>
rect 29 169 30 170 
<< m1 >>
rect 30 169 31 170 
<< m1 >>
rect 31 169 32 170 
<< m1 >>
rect 37 169 38 170 
<< m2 >>
rect 38 169 39 170 
<< m1 >>
rect 73 169 74 170 
<< m2 >>
rect 77 169 78 170 
<< m1 >>
rect 118 169 119 170 
<< m1 >>
rect 142 169 143 170 
<< m1 >>
rect 151 169 152 170 
<< m1 >>
rect 10 170 11 171 
<< m2 >>
rect 10 170 11 171 
<< m2 >>
rect 22 170 23 171 
<< m2 >>
rect 28 170 29 171 
<< m1 >>
rect 31 170 32 171 
<< m1 >>
rect 37 170 38 171 
<< m2 >>
rect 38 170 39 171 
<< m1 >>
rect 73 170 74 171 
<< m1 >>
rect 77 170 78 171 
<< m2 >>
rect 77 170 78 171 
<< m2c >>
rect 77 170 78 171 
<< m1 >>
rect 77 170 78 171 
<< m2 >>
rect 77 170 78 171 
<< m1 >>
rect 118 170 119 171 
<< m1 >>
rect 142 170 143 171 
<< m1 >>
rect 151 170 152 171 
<< m1 >>
rect 10 171 11 172 
<< m2 >>
rect 10 171 11 172 
<< m1 >>
rect 22 171 23 172 
<< m2 >>
rect 22 171 23 172 
<< m2c >>
rect 22 171 23 172 
<< m1 >>
rect 22 171 23 172 
<< m2 >>
rect 22 171 23 172 
<< m1 >>
rect 28 171 29 172 
<< m2 >>
rect 28 171 29 172 
<< m2c >>
rect 28 171 29 172 
<< m1 >>
rect 28 171 29 172 
<< m2 >>
rect 28 171 29 172 
<< m1 >>
rect 31 171 32 172 
<< m1 >>
rect 37 171 38 172 
<< m2 >>
rect 38 171 39 172 
<< m1 >>
rect 73 171 74 172 
<< m1 >>
rect 77 171 78 172 
<< m1 >>
rect 118 171 119 172 
<< m1 >>
rect 142 171 143 172 
<< m1 >>
rect 151 171 152 172 
<< m1 >>
rect 10 172 11 173 
<< m2 >>
rect 10 172 11 173 
<< m1 >>
rect 11 172 12 173 
<< m1 >>
rect 12 172 13 173 
<< m1 >>
rect 13 172 14 173 
<< m1 >>
rect 22 172 23 173 
<< m1 >>
rect 28 172 29 173 
<< m1 >>
rect 31 172 32 173 
<< m1 >>
rect 37 172 38 173 
<< m2 >>
rect 38 172 39 173 
<< m1 >>
rect 73 172 74 173 
<< m1 >>
rect 77 172 78 173 
<< m1 >>
rect 118 172 119 173 
<< m1 >>
rect 142 172 143 173 
<< m1 >>
rect 151 172 152 173 
<< m2 >>
rect 10 173 11 174 
<< m1 >>
rect 13 173 14 174 
<< m1 >>
rect 22 173 23 174 
<< m1 >>
rect 28 173 29 174 
<< m1 >>
rect 31 173 32 174 
<< m1 >>
rect 37 173 38 174 
<< m2 >>
rect 38 173 39 174 
<< m1 >>
rect 73 173 74 174 
<< m1 >>
rect 77 173 78 174 
<< m1 >>
rect 118 173 119 174 
<< m1 >>
rect 142 173 143 174 
<< m1 >>
rect 151 173 152 174 
<< m1 >>
rect 10 174 11 175 
<< m2 >>
rect 10 174 11 175 
<< m2c >>
rect 10 174 11 175 
<< m1 >>
rect 10 174 11 175 
<< m2 >>
rect 10 174 11 175 
<< pdiffusion >>
rect 12 174 13 175 
<< m1 >>
rect 13 174 14 175 
<< pdiffusion >>
rect 13 174 14 175 
<< pdiffusion >>
rect 14 174 15 175 
<< pdiffusion >>
rect 15 174 16 175 
<< pdiffusion >>
rect 16 174 17 175 
<< pdiffusion >>
rect 17 174 18 175 
<< m1 >>
rect 22 174 23 175 
<< m1 >>
rect 28 174 29 175 
<< pdiffusion >>
rect 30 174 31 175 
<< m1 >>
rect 31 174 32 175 
<< pdiffusion >>
rect 31 174 32 175 
<< pdiffusion >>
rect 32 174 33 175 
<< pdiffusion >>
rect 33 174 34 175 
<< pdiffusion >>
rect 34 174 35 175 
<< pdiffusion >>
rect 35 174 36 175 
<< m1 >>
rect 37 174 38 175 
<< m2 >>
rect 38 174 39 175 
<< m1 >>
rect 73 174 74 175 
<< m1 >>
rect 77 174 78 175 
<< pdiffusion >>
rect 84 174 85 175 
<< pdiffusion >>
rect 85 174 86 175 
<< pdiffusion >>
rect 86 174 87 175 
<< pdiffusion >>
rect 87 174 88 175 
<< pdiffusion >>
rect 88 174 89 175 
<< pdiffusion >>
rect 89 174 90 175 
<< pdiffusion >>
rect 102 174 103 175 
<< pdiffusion >>
rect 103 174 104 175 
<< pdiffusion >>
rect 104 174 105 175 
<< pdiffusion >>
rect 105 174 106 175 
<< pdiffusion >>
rect 106 174 107 175 
<< pdiffusion >>
rect 107 174 108 175 
<< m1 >>
rect 118 174 119 175 
<< pdiffusion >>
rect 120 174 121 175 
<< pdiffusion >>
rect 121 174 122 175 
<< pdiffusion >>
rect 122 174 123 175 
<< pdiffusion >>
rect 123 174 124 175 
<< pdiffusion >>
rect 124 174 125 175 
<< pdiffusion >>
rect 125 174 126 175 
<< pdiffusion >>
rect 138 174 139 175 
<< pdiffusion >>
rect 139 174 140 175 
<< pdiffusion >>
rect 140 174 141 175 
<< pdiffusion >>
rect 141 174 142 175 
<< m1 >>
rect 142 174 143 175 
<< pdiffusion >>
rect 142 174 143 175 
<< pdiffusion >>
rect 143 174 144 175 
<< m1 >>
rect 151 174 152 175 
<< m1 >>
rect 10 175 11 176 
<< pdiffusion >>
rect 12 175 13 176 
<< pdiffusion >>
rect 13 175 14 176 
<< pdiffusion >>
rect 14 175 15 176 
<< pdiffusion >>
rect 15 175 16 176 
<< pdiffusion >>
rect 16 175 17 176 
<< pdiffusion >>
rect 17 175 18 176 
<< m1 >>
rect 22 175 23 176 
<< m1 >>
rect 28 175 29 176 
<< pdiffusion >>
rect 30 175 31 176 
<< pdiffusion >>
rect 31 175 32 176 
<< pdiffusion >>
rect 32 175 33 176 
<< pdiffusion >>
rect 33 175 34 176 
<< pdiffusion >>
rect 34 175 35 176 
<< pdiffusion >>
rect 35 175 36 176 
<< m1 >>
rect 37 175 38 176 
<< m2 >>
rect 38 175 39 176 
<< m1 >>
rect 73 175 74 176 
<< m1 >>
rect 77 175 78 176 
<< pdiffusion >>
rect 84 175 85 176 
<< pdiffusion >>
rect 85 175 86 176 
<< pdiffusion >>
rect 86 175 87 176 
<< pdiffusion >>
rect 87 175 88 176 
<< pdiffusion >>
rect 88 175 89 176 
<< pdiffusion >>
rect 89 175 90 176 
<< pdiffusion >>
rect 102 175 103 176 
<< pdiffusion >>
rect 103 175 104 176 
<< pdiffusion >>
rect 104 175 105 176 
<< pdiffusion >>
rect 105 175 106 176 
<< pdiffusion >>
rect 106 175 107 176 
<< pdiffusion >>
rect 107 175 108 176 
<< m1 >>
rect 118 175 119 176 
<< pdiffusion >>
rect 120 175 121 176 
<< pdiffusion >>
rect 121 175 122 176 
<< pdiffusion >>
rect 122 175 123 176 
<< pdiffusion >>
rect 123 175 124 176 
<< pdiffusion >>
rect 124 175 125 176 
<< pdiffusion >>
rect 125 175 126 176 
<< pdiffusion >>
rect 138 175 139 176 
<< pdiffusion >>
rect 139 175 140 176 
<< pdiffusion >>
rect 140 175 141 176 
<< pdiffusion >>
rect 141 175 142 176 
<< pdiffusion >>
rect 142 175 143 176 
<< pdiffusion >>
rect 143 175 144 176 
<< m1 >>
rect 151 175 152 176 
<< m1 >>
rect 10 176 11 177 
<< pdiffusion >>
rect 12 176 13 177 
<< pdiffusion >>
rect 13 176 14 177 
<< pdiffusion >>
rect 14 176 15 177 
<< pdiffusion >>
rect 15 176 16 177 
<< pdiffusion >>
rect 16 176 17 177 
<< pdiffusion >>
rect 17 176 18 177 
<< m1 >>
rect 22 176 23 177 
<< m1 >>
rect 28 176 29 177 
<< pdiffusion >>
rect 30 176 31 177 
<< pdiffusion >>
rect 31 176 32 177 
<< pdiffusion >>
rect 32 176 33 177 
<< pdiffusion >>
rect 33 176 34 177 
<< pdiffusion >>
rect 34 176 35 177 
<< pdiffusion >>
rect 35 176 36 177 
<< m1 >>
rect 37 176 38 177 
<< m2 >>
rect 38 176 39 177 
<< m1 >>
rect 73 176 74 177 
<< m1 >>
rect 77 176 78 177 
<< pdiffusion >>
rect 84 176 85 177 
<< pdiffusion >>
rect 85 176 86 177 
<< pdiffusion >>
rect 86 176 87 177 
<< pdiffusion >>
rect 87 176 88 177 
<< pdiffusion >>
rect 88 176 89 177 
<< pdiffusion >>
rect 89 176 90 177 
<< pdiffusion >>
rect 102 176 103 177 
<< pdiffusion >>
rect 103 176 104 177 
<< pdiffusion >>
rect 104 176 105 177 
<< pdiffusion >>
rect 105 176 106 177 
<< pdiffusion >>
rect 106 176 107 177 
<< pdiffusion >>
rect 107 176 108 177 
<< m1 >>
rect 118 176 119 177 
<< pdiffusion >>
rect 120 176 121 177 
<< pdiffusion >>
rect 121 176 122 177 
<< pdiffusion >>
rect 122 176 123 177 
<< pdiffusion >>
rect 123 176 124 177 
<< pdiffusion >>
rect 124 176 125 177 
<< pdiffusion >>
rect 125 176 126 177 
<< pdiffusion >>
rect 138 176 139 177 
<< pdiffusion >>
rect 139 176 140 177 
<< pdiffusion >>
rect 140 176 141 177 
<< pdiffusion >>
rect 141 176 142 177 
<< pdiffusion >>
rect 142 176 143 177 
<< pdiffusion >>
rect 143 176 144 177 
<< m1 >>
rect 151 176 152 177 
<< m1 >>
rect 10 177 11 178 
<< pdiffusion >>
rect 12 177 13 178 
<< pdiffusion >>
rect 13 177 14 178 
<< pdiffusion >>
rect 14 177 15 178 
<< pdiffusion >>
rect 15 177 16 178 
<< pdiffusion >>
rect 16 177 17 178 
<< pdiffusion >>
rect 17 177 18 178 
<< m1 >>
rect 22 177 23 178 
<< m1 >>
rect 28 177 29 178 
<< pdiffusion >>
rect 30 177 31 178 
<< pdiffusion >>
rect 31 177 32 178 
<< pdiffusion >>
rect 32 177 33 178 
<< pdiffusion >>
rect 33 177 34 178 
<< pdiffusion >>
rect 34 177 35 178 
<< pdiffusion >>
rect 35 177 36 178 
<< m1 >>
rect 37 177 38 178 
<< m2 >>
rect 38 177 39 178 
<< m1 >>
rect 73 177 74 178 
<< m1 >>
rect 77 177 78 178 
<< pdiffusion >>
rect 84 177 85 178 
<< pdiffusion >>
rect 85 177 86 178 
<< pdiffusion >>
rect 86 177 87 178 
<< pdiffusion >>
rect 87 177 88 178 
<< pdiffusion >>
rect 88 177 89 178 
<< pdiffusion >>
rect 89 177 90 178 
<< pdiffusion >>
rect 102 177 103 178 
<< pdiffusion >>
rect 103 177 104 178 
<< pdiffusion >>
rect 104 177 105 178 
<< pdiffusion >>
rect 105 177 106 178 
<< pdiffusion >>
rect 106 177 107 178 
<< pdiffusion >>
rect 107 177 108 178 
<< m1 >>
rect 118 177 119 178 
<< pdiffusion >>
rect 120 177 121 178 
<< pdiffusion >>
rect 121 177 122 178 
<< pdiffusion >>
rect 122 177 123 178 
<< pdiffusion >>
rect 123 177 124 178 
<< pdiffusion >>
rect 124 177 125 178 
<< pdiffusion >>
rect 125 177 126 178 
<< pdiffusion >>
rect 138 177 139 178 
<< pdiffusion >>
rect 139 177 140 178 
<< pdiffusion >>
rect 140 177 141 178 
<< pdiffusion >>
rect 141 177 142 178 
<< pdiffusion >>
rect 142 177 143 178 
<< pdiffusion >>
rect 143 177 144 178 
<< m1 >>
rect 151 177 152 178 
<< m1 >>
rect 10 178 11 179 
<< pdiffusion >>
rect 12 178 13 179 
<< pdiffusion >>
rect 13 178 14 179 
<< pdiffusion >>
rect 14 178 15 179 
<< pdiffusion >>
rect 15 178 16 179 
<< pdiffusion >>
rect 16 178 17 179 
<< pdiffusion >>
rect 17 178 18 179 
<< m1 >>
rect 22 178 23 179 
<< m1 >>
rect 28 178 29 179 
<< pdiffusion >>
rect 30 178 31 179 
<< pdiffusion >>
rect 31 178 32 179 
<< pdiffusion >>
rect 32 178 33 179 
<< pdiffusion >>
rect 33 178 34 179 
<< pdiffusion >>
rect 34 178 35 179 
<< pdiffusion >>
rect 35 178 36 179 
<< m1 >>
rect 37 178 38 179 
<< m2 >>
rect 38 178 39 179 
<< m1 >>
rect 73 178 74 179 
<< m1 >>
rect 77 178 78 179 
<< pdiffusion >>
rect 84 178 85 179 
<< pdiffusion >>
rect 85 178 86 179 
<< pdiffusion >>
rect 86 178 87 179 
<< pdiffusion >>
rect 87 178 88 179 
<< pdiffusion >>
rect 88 178 89 179 
<< pdiffusion >>
rect 89 178 90 179 
<< pdiffusion >>
rect 102 178 103 179 
<< pdiffusion >>
rect 103 178 104 179 
<< pdiffusion >>
rect 104 178 105 179 
<< pdiffusion >>
rect 105 178 106 179 
<< pdiffusion >>
rect 106 178 107 179 
<< pdiffusion >>
rect 107 178 108 179 
<< m1 >>
rect 118 178 119 179 
<< pdiffusion >>
rect 120 178 121 179 
<< pdiffusion >>
rect 121 178 122 179 
<< pdiffusion >>
rect 122 178 123 179 
<< pdiffusion >>
rect 123 178 124 179 
<< pdiffusion >>
rect 124 178 125 179 
<< pdiffusion >>
rect 125 178 126 179 
<< pdiffusion >>
rect 138 178 139 179 
<< pdiffusion >>
rect 139 178 140 179 
<< pdiffusion >>
rect 140 178 141 179 
<< pdiffusion >>
rect 141 178 142 179 
<< pdiffusion >>
rect 142 178 143 179 
<< pdiffusion >>
rect 143 178 144 179 
<< m1 >>
rect 151 178 152 179 
<< m1 >>
rect 10 179 11 180 
<< pdiffusion >>
rect 12 179 13 180 
<< m1 >>
rect 13 179 14 180 
<< pdiffusion >>
rect 13 179 14 180 
<< pdiffusion >>
rect 14 179 15 180 
<< pdiffusion >>
rect 15 179 16 180 
<< pdiffusion >>
rect 16 179 17 180 
<< pdiffusion >>
rect 17 179 18 180 
<< m1 >>
rect 22 179 23 180 
<< m1 >>
rect 28 179 29 180 
<< pdiffusion >>
rect 30 179 31 180 
<< pdiffusion >>
rect 31 179 32 180 
<< pdiffusion >>
rect 32 179 33 180 
<< pdiffusion >>
rect 33 179 34 180 
<< m1 >>
rect 34 179 35 180 
<< pdiffusion >>
rect 34 179 35 180 
<< pdiffusion >>
rect 35 179 36 180 
<< m1 >>
rect 37 179 38 180 
<< m2 >>
rect 38 179 39 180 
<< m2 >>
rect 72 179 73 180 
<< m1 >>
rect 73 179 74 180 
<< m2 >>
rect 73 179 74 180 
<< m2 >>
rect 74 179 75 180 
<< m1 >>
rect 75 179 76 180 
<< m2 >>
rect 75 179 76 180 
<< m2c >>
rect 75 179 76 180 
<< m1 >>
rect 75 179 76 180 
<< m2 >>
rect 75 179 76 180 
<< m1 >>
rect 76 179 77 180 
<< m1 >>
rect 77 179 78 180 
<< pdiffusion >>
rect 84 179 85 180 
<< m1 >>
rect 85 179 86 180 
<< pdiffusion >>
rect 85 179 86 180 
<< pdiffusion >>
rect 86 179 87 180 
<< pdiffusion >>
rect 87 179 88 180 
<< pdiffusion >>
rect 88 179 89 180 
<< pdiffusion >>
rect 89 179 90 180 
<< pdiffusion >>
rect 102 179 103 180 
<< pdiffusion >>
rect 103 179 104 180 
<< pdiffusion >>
rect 104 179 105 180 
<< pdiffusion >>
rect 105 179 106 180 
<< m1 >>
rect 106 179 107 180 
<< pdiffusion >>
rect 106 179 107 180 
<< pdiffusion >>
rect 107 179 108 180 
<< m1 >>
rect 118 179 119 180 
<< pdiffusion >>
rect 120 179 121 180 
<< pdiffusion >>
rect 121 179 122 180 
<< pdiffusion >>
rect 122 179 123 180 
<< pdiffusion >>
rect 123 179 124 180 
<< m1 >>
rect 124 179 125 180 
<< pdiffusion >>
rect 124 179 125 180 
<< pdiffusion >>
rect 125 179 126 180 
<< pdiffusion >>
rect 138 179 139 180 
<< pdiffusion >>
rect 139 179 140 180 
<< pdiffusion >>
rect 140 179 141 180 
<< pdiffusion >>
rect 141 179 142 180 
<< pdiffusion >>
rect 142 179 143 180 
<< pdiffusion >>
rect 143 179 144 180 
<< m1 >>
rect 151 179 152 180 
<< m1 >>
rect 10 180 11 181 
<< m1 >>
rect 13 180 14 181 
<< m1 >>
rect 22 180 23 181 
<< m1 >>
rect 28 180 29 181 
<< m1 >>
rect 34 180 35 181 
<< m1 >>
rect 37 180 38 181 
<< m2 >>
rect 38 180 39 181 
<< m2 >>
rect 72 180 73 181 
<< m1 >>
rect 73 180 74 181 
<< m1 >>
rect 85 180 86 181 
<< m1 >>
rect 106 180 107 181 
<< m1 >>
rect 118 180 119 181 
<< m1 >>
rect 124 180 125 181 
<< m1 >>
rect 151 180 152 181 
<< m1 >>
rect 10 181 11 182 
<< m1 >>
rect 11 181 12 182 
<< m1 >>
rect 12 181 13 182 
<< m1 >>
rect 13 181 14 182 
<< m1 >>
rect 22 181 23 182 
<< m1 >>
rect 28 181 29 182 
<< m1 >>
rect 34 181 35 182 
<< m1 >>
rect 35 181 36 182 
<< m2 >>
rect 35 181 36 182 
<< m2c >>
rect 35 181 36 182 
<< m1 >>
rect 35 181 36 182 
<< m2 >>
rect 35 181 36 182 
<< m2 >>
rect 36 181 37 182 
<< m1 >>
rect 37 181 38 182 
<< m2 >>
rect 37 181 38 182 
<< m2 >>
rect 38 181 39 182 
<< m2 >>
rect 72 181 73 182 
<< m1 >>
rect 73 181 74 182 
<< m1 >>
rect 74 181 75 182 
<< m1 >>
rect 75 181 76 182 
<< m1 >>
rect 76 181 77 182 
<< m1 >>
rect 77 181 78 182 
<< m1 >>
rect 78 181 79 182 
<< m1 >>
rect 79 181 80 182 
<< m1 >>
rect 80 181 81 182 
<< m1 >>
rect 81 181 82 182 
<< m1 >>
rect 82 181 83 182 
<< m1 >>
rect 83 181 84 182 
<< m1 >>
rect 84 181 85 182 
<< m1 >>
rect 85 181 86 182 
<< m1 >>
rect 106 181 107 182 
<< m1 >>
rect 107 181 108 182 
<< m1 >>
rect 108 181 109 182 
<< m1 >>
rect 109 181 110 182 
<< m1 >>
rect 110 181 111 182 
<< m1 >>
rect 111 181 112 182 
<< m1 >>
rect 112 181 113 182 
<< m1 >>
rect 113 181 114 182 
<< m1 >>
rect 114 181 115 182 
<< m1 >>
rect 115 181 116 182 
<< m1 >>
rect 116 181 117 182 
<< m1 >>
rect 117 181 118 182 
<< m1 >>
rect 118 181 119 182 
<< m1 >>
rect 124 181 125 182 
<< m1 >>
rect 151 181 152 182 
<< m1 >>
rect 22 182 23 183 
<< m1 >>
rect 28 182 29 183 
<< m1 >>
rect 29 182 30 183 
<< m1 >>
rect 30 182 31 183 
<< m2 >>
rect 30 182 31 183 
<< m2c >>
rect 30 182 31 183 
<< m1 >>
rect 30 182 31 183 
<< m2 >>
rect 30 182 31 183 
<< m1 >>
rect 37 182 38 183 
<< m2 >>
rect 72 182 73 183 
<< m1 >>
rect 124 182 125 183 
<< m1 >>
rect 151 182 152 183 
<< m1 >>
rect 22 183 23 184 
<< m2 >>
rect 30 183 31 184 
<< m1 >>
rect 37 183 38 184 
<< m2 >>
rect 72 183 73 184 
<< m1 >>
rect 124 183 125 184 
<< m1 >>
rect 151 183 152 184 
<< m1 >>
rect 22 184 23 185 
<< m1 >>
rect 23 184 24 185 
<< m1 >>
rect 24 184 25 185 
<< m1 >>
rect 25 184 26 185 
<< m1 >>
rect 26 184 27 185 
<< m1 >>
rect 27 184 28 185 
<< m1 >>
rect 28 184 29 185 
<< m1 >>
rect 29 184 30 185 
<< m1 >>
rect 30 184 31 185 
<< m2 >>
rect 30 184 31 185 
<< m1 >>
rect 31 184 32 185 
<< m1 >>
rect 32 184 33 185 
<< m1 >>
rect 33 184 34 185 
<< m1 >>
rect 34 184 35 185 
<< m1 >>
rect 35 184 36 185 
<< m2 >>
rect 35 184 36 185 
<< m2c >>
rect 35 184 36 185 
<< m1 >>
rect 35 184 36 185 
<< m2 >>
rect 35 184 36 185 
<< m2 >>
rect 36 184 37 185 
<< m1 >>
rect 37 184 38 185 
<< m2 >>
rect 37 184 38 185 
<< m1 >>
rect 38 184 39 185 
<< m2 >>
rect 38 184 39 185 
<< m1 >>
rect 39 184 40 185 
<< m2 >>
rect 39 184 40 185 
<< m1 >>
rect 40 184 41 185 
<< m2 >>
rect 40 184 41 185 
<< m1 >>
rect 41 184 42 185 
<< m2 >>
rect 41 184 42 185 
<< m1 >>
rect 42 184 43 185 
<< m2 >>
rect 42 184 43 185 
<< m1 >>
rect 43 184 44 185 
<< m2 >>
rect 43 184 44 185 
<< m1 >>
rect 44 184 45 185 
<< m2 >>
rect 44 184 45 185 
<< m1 >>
rect 45 184 46 185 
<< m2 >>
rect 45 184 46 185 
<< m1 >>
rect 46 184 47 185 
<< m2 >>
rect 46 184 47 185 
<< m1 >>
rect 47 184 48 185 
<< m2 >>
rect 47 184 48 185 
<< m1 >>
rect 48 184 49 185 
<< m2 >>
rect 48 184 49 185 
<< m1 >>
rect 49 184 50 185 
<< m2 >>
rect 49 184 50 185 
<< m1 >>
rect 50 184 51 185 
<< m2 >>
rect 50 184 51 185 
<< m1 >>
rect 51 184 52 185 
<< m2 >>
rect 51 184 52 185 
<< m1 >>
rect 52 184 53 185 
<< m2 >>
rect 52 184 53 185 
<< m1 >>
rect 53 184 54 185 
<< m2 >>
rect 53 184 54 185 
<< m1 >>
rect 54 184 55 185 
<< m2 >>
rect 54 184 55 185 
<< m1 >>
rect 55 184 56 185 
<< m2 >>
rect 55 184 56 185 
<< m1 >>
rect 56 184 57 185 
<< m2 >>
rect 56 184 57 185 
<< m1 >>
rect 57 184 58 185 
<< m2 >>
rect 57 184 58 185 
<< m1 >>
rect 58 184 59 185 
<< m2 >>
rect 58 184 59 185 
<< m1 >>
rect 59 184 60 185 
<< m2 >>
rect 59 184 60 185 
<< m1 >>
rect 60 184 61 185 
<< m2 >>
rect 60 184 61 185 
<< m1 >>
rect 61 184 62 185 
<< m2 >>
rect 61 184 62 185 
<< m1 >>
rect 62 184 63 185 
<< m2 >>
rect 62 184 63 185 
<< m1 >>
rect 63 184 64 185 
<< m2 >>
rect 63 184 64 185 
<< m1 >>
rect 64 184 65 185 
<< m2 >>
rect 64 184 65 185 
<< m1 >>
rect 65 184 66 185 
<< m2 >>
rect 65 184 66 185 
<< m1 >>
rect 66 184 67 185 
<< m2 >>
rect 66 184 67 185 
<< m1 >>
rect 67 184 68 185 
<< m2 >>
rect 67 184 68 185 
<< m1 >>
rect 68 184 69 185 
<< m2 >>
rect 68 184 69 185 
<< m1 >>
rect 69 184 70 185 
<< m2 >>
rect 69 184 70 185 
<< m1 >>
rect 70 184 71 185 
<< m2 >>
rect 70 184 71 185 
<< m1 >>
rect 71 184 72 185 
<< m2 >>
rect 71 184 72 185 
<< m1 >>
rect 72 184 73 185 
<< m2 >>
rect 72 184 73 185 
<< m1 >>
rect 73 184 74 185 
<< m1 >>
rect 74 184 75 185 
<< m1 >>
rect 75 184 76 185 
<< m1 >>
rect 76 184 77 185 
<< m1 >>
rect 77 184 78 185 
<< m1 >>
rect 78 184 79 185 
<< m1 >>
rect 79 184 80 185 
<< m1 >>
rect 80 184 81 185 
<< m1 >>
rect 81 184 82 185 
<< m1 >>
rect 82 184 83 185 
<< m1 >>
rect 83 184 84 185 
<< m1 >>
rect 84 184 85 185 
<< m1 >>
rect 85 184 86 185 
<< m1 >>
rect 86 184 87 185 
<< m1 >>
rect 87 184 88 185 
<< m1 >>
rect 88 184 89 185 
<< m1 >>
rect 89 184 90 185 
<< m1 >>
rect 90 184 91 185 
<< m1 >>
rect 91 184 92 185 
<< m1 >>
rect 92 184 93 185 
<< m1 >>
rect 93 184 94 185 
<< m1 >>
rect 94 184 95 185 
<< m1 >>
rect 95 184 96 185 
<< m1 >>
rect 96 184 97 185 
<< m1 >>
rect 97 184 98 185 
<< m1 >>
rect 98 184 99 185 
<< m1 >>
rect 99 184 100 185 
<< m1 >>
rect 100 184 101 185 
<< m1 >>
rect 101 184 102 185 
<< m1 >>
rect 102 184 103 185 
<< m1 >>
rect 103 184 104 185 
<< m1 >>
rect 104 184 105 185 
<< m1 >>
rect 105 184 106 185 
<< m1 >>
rect 106 184 107 185 
<< m1 >>
rect 107 184 108 185 
<< m1 >>
rect 108 184 109 185 
<< m1 >>
rect 109 184 110 185 
<< m1 >>
rect 110 184 111 185 
<< m1 >>
rect 111 184 112 185 
<< m1 >>
rect 112 184 113 185 
<< m1 >>
rect 113 184 114 185 
<< m1 >>
rect 114 184 115 185 
<< m1 >>
rect 115 184 116 185 
<< m1 >>
rect 116 184 117 185 
<< m1 >>
rect 117 184 118 185 
<< m1 >>
rect 118 184 119 185 
<< m1 >>
rect 119 184 120 185 
<< m1 >>
rect 120 184 121 185 
<< m1 >>
rect 121 184 122 185 
<< m1 >>
rect 122 184 123 185 
<< m1 >>
rect 123 184 124 185 
<< m1 >>
rect 124 184 125 185 
<< m1 >>
rect 151 184 152 185 
<< m2 >>
rect 30 185 31 186 
<< m2 >>
rect 31 185 32 186 
<< m2 >>
rect 32 185 33 186 
<< m2 >>
rect 33 185 34 186 
<< m1 >>
rect 151 185 152 186 
<< m1 >>
rect 33 186 34 187 
<< m2 >>
rect 33 186 34 187 
<< m2c >>
rect 33 186 34 187 
<< m1 >>
rect 33 186 34 187 
<< m2 >>
rect 33 186 34 187 
<< m1 >>
rect 34 186 35 187 
<< m1 >>
rect 35 186 36 187 
<< m1 >>
rect 36 186 37 187 
<< m1 >>
rect 37 186 38 187 
<< m1 >>
rect 38 186 39 187 
<< m1 >>
rect 39 186 40 187 
<< m1 >>
rect 40 186 41 187 
<< m1 >>
rect 41 186 42 187 
<< m1 >>
rect 42 186 43 187 
<< m1 >>
rect 43 186 44 187 
<< m1 >>
rect 44 186 45 187 
<< m1 >>
rect 45 186 46 187 
<< m1 >>
rect 46 186 47 187 
<< m1 >>
rect 47 186 48 187 
<< m1 >>
rect 48 186 49 187 
<< m1 >>
rect 49 186 50 187 
<< m1 >>
rect 50 186 51 187 
<< m1 >>
rect 51 186 52 187 
<< m1 >>
rect 52 186 53 187 
<< m1 >>
rect 53 186 54 187 
<< m1 >>
rect 54 186 55 187 
<< m1 >>
rect 55 186 56 187 
<< m1 >>
rect 56 186 57 187 
<< m1 >>
rect 57 186 58 187 
<< m1 >>
rect 58 186 59 187 
<< m1 >>
rect 59 186 60 187 
<< m1 >>
rect 60 186 61 187 
<< m1 >>
rect 61 186 62 187 
<< m1 >>
rect 62 186 63 187 
<< m1 >>
rect 63 186 64 187 
<< m1 >>
rect 64 186 65 187 
<< m1 >>
rect 65 186 66 187 
<< m1 >>
rect 66 186 67 187 
<< m1 >>
rect 67 186 68 187 
<< m1 >>
rect 68 186 69 187 
<< m1 >>
rect 69 186 70 187 
<< m1 >>
rect 70 186 71 187 
<< m1 >>
rect 71 186 72 187 
<< m1 >>
rect 72 186 73 187 
<< m1 >>
rect 73 186 74 187 
<< m1 >>
rect 74 186 75 187 
<< m1 >>
rect 75 186 76 187 
<< m1 >>
rect 76 186 77 187 
<< m1 >>
rect 77 186 78 187 
<< m1 >>
rect 78 186 79 187 
<< m1 >>
rect 79 186 80 187 
<< m1 >>
rect 80 186 81 187 
<< m1 >>
rect 81 186 82 187 
<< m1 >>
rect 82 186 83 187 
<< m1 >>
rect 83 186 84 187 
<< m1 >>
rect 84 186 85 187 
<< m1 >>
rect 85 186 86 187 
<< m1 >>
rect 86 186 87 187 
<< m1 >>
rect 87 186 88 187 
<< m1 >>
rect 88 186 89 187 
<< m1 >>
rect 89 186 90 187 
<< m1 >>
rect 90 186 91 187 
<< m1 >>
rect 91 186 92 187 
<< m1 >>
rect 92 186 93 187 
<< m1 >>
rect 93 186 94 187 
<< m1 >>
rect 94 186 95 187 
<< m1 >>
rect 95 186 96 187 
<< m1 >>
rect 96 186 97 187 
<< m1 >>
rect 97 186 98 187 
<< m1 >>
rect 98 186 99 187 
<< m1 >>
rect 99 186 100 187 
<< m1 >>
rect 100 186 101 187 
<< m1 >>
rect 101 186 102 187 
<< m1 >>
rect 102 186 103 187 
<< m1 >>
rect 103 186 104 187 
<< m1 >>
rect 104 186 105 187 
<< m1 >>
rect 105 186 106 187 
<< m1 >>
rect 106 186 107 187 
<< m1 >>
rect 107 186 108 187 
<< m1 >>
rect 108 186 109 187 
<< m1 >>
rect 109 186 110 187 
<< m1 >>
rect 110 186 111 187 
<< m1 >>
rect 111 186 112 187 
<< m1 >>
rect 112 186 113 187 
<< m1 >>
rect 113 186 114 187 
<< m1 >>
rect 114 186 115 187 
<< m1 >>
rect 115 186 116 187 
<< m1 >>
rect 116 186 117 187 
<< m1 >>
rect 117 186 118 187 
<< m1 >>
rect 118 186 119 187 
<< m1 >>
rect 119 186 120 187 
<< m1 >>
rect 120 186 121 187 
<< m1 >>
rect 121 186 122 187 
<< m1 >>
rect 122 186 123 187 
<< m1 >>
rect 123 186 124 187 
<< m1 >>
rect 124 186 125 187 
<< m1 >>
rect 125 186 126 187 
<< m1 >>
rect 126 186 127 187 
<< m1 >>
rect 127 186 128 187 
<< m1 >>
rect 128 186 129 187 
<< m1 >>
rect 129 186 130 187 
<< m1 >>
rect 130 186 131 187 
<< m1 >>
rect 131 186 132 187 
<< m1 >>
rect 132 186 133 187 
<< m1 >>
rect 133 186 134 187 
<< m1 >>
rect 134 186 135 187 
<< m1 >>
rect 135 186 136 187 
<< m1 >>
rect 136 186 137 187 
<< m1 >>
rect 137 186 138 187 
<< m1 >>
rect 138 186 139 187 
<< m1 >>
rect 139 186 140 187 
<< m1 >>
rect 140 186 141 187 
<< m1 >>
rect 141 186 142 187 
<< m1 >>
rect 142 186 143 187 
<< m1 >>
rect 143 186 144 187 
<< m1 >>
rect 144 186 145 187 
<< m1 >>
rect 145 186 146 187 
<< m1 >>
rect 146 186 147 187 
<< m1 >>
rect 147 186 148 187 
<< m1 >>
rect 148 186 149 187 
<< m1 >>
rect 149 186 150 187 
<< m1 >>
rect 150 186 151 187 
<< m1 >>
rect 151 186 152 187 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 1
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 2
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 3
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 4
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 139 30 140 31  0 t = 1
rlabel pdiffusion 142 30 143 31  0 t = 2
rlabel pdiffusion 139 35 140 36  0 t = 3
rlabel pdiffusion 142 35 143 36  0 t = 4
rlabel pdiffusion 138 30 144 36 0 cell no = 5
<< m1 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2c >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< labels >>
rlabel pdiffusion 67 138 68 139  0 t = 1
rlabel pdiffusion 70 138 71 139  0 t = 2
rlabel pdiffusion 67 143 68 144  0 t = 3
rlabel pdiffusion 70 143 71 144  0 t = 4
rlabel pdiffusion 66 138 72 144 0 cell no = 6
<< m1 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2c >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< labels >>
rlabel pdiffusion 103 138 104 139  0 t = 1
rlabel pdiffusion 106 138 107 139  0 t = 2
rlabel pdiffusion 103 143 104 144  0 t = 3
rlabel pdiffusion 106 143 107 144  0 t = 4
rlabel pdiffusion 102 138 108 144 0 cell no = 7
<< m1 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2c >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 8
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 175 120 176 121  0 t = 1
rlabel pdiffusion 178 120 179 121  0 t = 2
rlabel pdiffusion 175 125 176 126  0 t = 3
rlabel pdiffusion 178 125 179 126  0 t = 4
rlabel pdiffusion 174 120 180 126 0 cell no = 9
<< m1 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2c >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< labels >>
rlabel pdiffusion 67 120 68 121  0 t = 1
rlabel pdiffusion 70 120 71 121  0 t = 2
rlabel pdiffusion 67 125 68 126  0 t = 3
rlabel pdiffusion 70 125 71 126  0 t = 4
rlabel pdiffusion 66 120 72 126 0 cell no = 10
<< m1 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2c >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< labels >>
rlabel pdiffusion 175 12 176 13  0 t = 1
rlabel pdiffusion 178 12 179 13  0 t = 2
rlabel pdiffusion 175 17 176 18  0 t = 3
rlabel pdiffusion 178 17 179 18  0 t = 4
rlabel pdiffusion 174 12 180 18 0 cell no = 11
<< m1 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2c >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< labels >>
rlabel pdiffusion 85 12 86 13  0 t = 1
rlabel pdiffusion 88 12 89 13  0 t = 2
rlabel pdiffusion 85 17 86 18  0 t = 3
rlabel pdiffusion 88 17 89 18  0 t = 4
rlabel pdiffusion 84 12 90 18 0 cell no = 12
<< m1 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2c >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 13
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 13 138 14 139  0 t = 1
rlabel pdiffusion 16 138 17 139  0 t = 2
rlabel pdiffusion 13 143 14 144  0 t = 3
rlabel pdiffusion 16 143 17 144  0 t = 4
rlabel pdiffusion 12 138 18 144 0 cell no = 14
<< m1 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2c >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< labels >>
rlabel pdiffusion 103 30 104 31  0 t = 1
rlabel pdiffusion 106 30 107 31  0 t = 2
rlabel pdiffusion 103 35 104 36  0 t = 3
rlabel pdiffusion 106 35 107 36  0 t = 4
rlabel pdiffusion 102 30 108 36 0 cell no = 15
<< m1 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2c >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< labels >>
rlabel pdiffusion 157 120 158 121  0 t = 1
rlabel pdiffusion 160 120 161 121  0 t = 2
rlabel pdiffusion 157 125 158 126  0 t = 3
rlabel pdiffusion 160 125 161 126  0 t = 4
rlabel pdiffusion 156 120 162 126 0 cell no = 16
<< m1 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2c >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 17
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 157 66 158 67  0 t = 1
rlabel pdiffusion 160 66 161 67  0 t = 2
rlabel pdiffusion 157 71 158 72  0 t = 3
rlabel pdiffusion 160 71 161 72  0 t = 4
rlabel pdiffusion 156 66 162 72 0 cell no = 18
<< m1 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2c >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 19
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 31 138 32 139  0 t = 1
rlabel pdiffusion 34 138 35 139  0 t = 2
rlabel pdiffusion 31 143 32 144  0 t = 3
rlabel pdiffusion 34 143 35 144  0 t = 4
rlabel pdiffusion 30 138 36 144 0 cell no = 20
<< m1 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2c >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 21
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 31 12 32 13  0 t = 1
rlabel pdiffusion 34 12 35 13  0 t = 2
rlabel pdiffusion 31 17 32 18  0 t = 3
rlabel pdiffusion 34 17 35 18  0 t = 4
rlabel pdiffusion 30 12 36 18 0 cell no = 22
<< m1 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2c >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 23
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 24
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 25
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 26
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 27
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 28
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 157 156 158 157  0 t = 1
rlabel pdiffusion 160 156 161 157  0 t = 2
rlabel pdiffusion 157 161 158 162  0 t = 3
rlabel pdiffusion 160 161 161 162  0 t = 4
rlabel pdiffusion 156 156 162 162 0 cell no = 29
<< m1 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2c >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 30
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 31
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 157 48 158 49  0 t = 1
rlabel pdiffusion 160 48 161 49  0 t = 2
rlabel pdiffusion 157 53 158 54  0 t = 3
rlabel pdiffusion 160 53 161 54  0 t = 4
rlabel pdiffusion 156 48 162 54 0 cell no = 32
<< m1 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2c >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< labels >>
rlabel pdiffusion 157 30 158 31  0 t = 1
rlabel pdiffusion 160 30 161 31  0 t = 2
rlabel pdiffusion 157 35 158 36  0 t = 3
rlabel pdiffusion 160 35 161 36  0 t = 4
rlabel pdiffusion 156 30 162 36 0 cell no = 33
<< m1 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2c >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< labels >>
rlabel pdiffusion 139 174 140 175  0 t = 1
rlabel pdiffusion 142 174 143 175  0 t = 2
rlabel pdiffusion 139 179 140 180  0 t = 3
rlabel pdiffusion 142 179 143 180  0 t = 4
rlabel pdiffusion 138 174 144 180 0 cell no = 34
<< m1 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2c >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 35
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 175 48 176 49  0 t = 1
rlabel pdiffusion 178 48 179 49  0 t = 2
rlabel pdiffusion 175 53 176 54  0 t = 3
rlabel pdiffusion 178 53 179 54  0 t = 4
rlabel pdiffusion 174 48 180 54 0 cell no = 36
<< m1 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2c >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< labels >>
rlabel pdiffusion 121 156 122 157  0 t = 1
rlabel pdiffusion 124 156 125 157  0 t = 2
rlabel pdiffusion 121 161 122 162  0 t = 3
rlabel pdiffusion 124 161 125 162  0 t = 4
rlabel pdiffusion 120 156 126 162 0 cell no = 37
<< m1 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2c >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 38
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 85 174 86 175  0 t = 1
rlabel pdiffusion 88 174 89 175  0 t = 2
rlabel pdiffusion 85 179 86 180  0 t = 3
rlabel pdiffusion 88 179 89 180  0 t = 4
rlabel pdiffusion 84 174 90 180 0 cell no = 39
<< m1 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2c >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< labels >>
rlabel pdiffusion 175 66 176 67  0 t = 1
rlabel pdiffusion 178 66 179 67  0 t = 2
rlabel pdiffusion 175 71 176 72  0 t = 3
rlabel pdiffusion 178 71 179 72  0 t = 4
rlabel pdiffusion 174 66 180 72 0 cell no = 40
<< m1 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2c >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< labels >>
rlabel pdiffusion 85 138 86 139  0 t = 1
rlabel pdiffusion 88 138 89 139  0 t = 2
rlabel pdiffusion 85 143 86 144  0 t = 3
rlabel pdiffusion 88 143 89 144  0 t = 4
rlabel pdiffusion 84 138 90 144 0 cell no = 41
<< m1 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2c >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< labels >>
rlabel pdiffusion 157 12 158 13  0 t = 1
rlabel pdiffusion 160 12 161 13  0 t = 2
rlabel pdiffusion 157 17 158 18  0 t = 3
rlabel pdiffusion 160 17 161 18  0 t = 4
rlabel pdiffusion 156 12 162 18 0 cell no = 42
<< m1 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2c >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 43
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 44
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 45
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 139 48 140 49  0 t = 1
rlabel pdiffusion 142 48 143 49  0 t = 2
rlabel pdiffusion 139 53 140 54  0 t = 3
rlabel pdiffusion 142 53 143 54  0 t = 4
rlabel pdiffusion 138 48 144 54 0 cell no = 46
<< m1 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2c >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< labels >>
rlabel pdiffusion 85 120 86 121  0 t = 1
rlabel pdiffusion 88 120 89 121  0 t = 2
rlabel pdiffusion 85 125 86 126  0 t = 3
rlabel pdiffusion 88 125 89 126  0 t = 4
rlabel pdiffusion 84 120 90 126 0 cell no = 47
<< m1 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2c >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 48
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 139 66 140 67  0 t = 1
rlabel pdiffusion 142 66 143 67  0 t = 2
rlabel pdiffusion 139 71 140 72  0 t = 3
rlabel pdiffusion 142 71 143 72  0 t = 4
rlabel pdiffusion 138 66 144 72 0 cell no = 49
<< m1 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2c >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 50
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 139 12 140 13  0 t = 1
rlabel pdiffusion 142 12 143 13  0 t = 2
rlabel pdiffusion 139 17 140 18  0 t = 3
rlabel pdiffusion 142 17 143 18  0 t = 4
rlabel pdiffusion 138 12 144 18 0 cell no = 51
<< m1 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2c >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< labels >>
rlabel pdiffusion 13 174 14 175  0 t = 1
rlabel pdiffusion 16 174 17 175  0 t = 2
rlabel pdiffusion 13 179 14 180  0 t = 3
rlabel pdiffusion 16 179 17 180  0 t = 4
rlabel pdiffusion 12 174 18 180 0 cell no = 52
<< m1 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2c >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< labels >>
rlabel pdiffusion 49 120 50 121  0 t = 1
rlabel pdiffusion 52 120 53 121  0 t = 2
rlabel pdiffusion 49 125 50 126  0 t = 3
rlabel pdiffusion 52 125 53 126  0 t = 4
rlabel pdiffusion 48 120 54 126 0 cell no = 53
<< m1 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2c >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 54
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 103 120 104 121  0 t = 1
rlabel pdiffusion 106 120 107 121  0 t = 2
rlabel pdiffusion 103 125 104 126  0 t = 3
rlabel pdiffusion 106 125 107 126  0 t = 4
rlabel pdiffusion 102 120 108 126 0 cell no = 55
<< m1 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2c >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< labels >>
rlabel pdiffusion 49 138 50 139  0 t = 1
rlabel pdiffusion 52 138 53 139  0 t = 2
rlabel pdiffusion 49 143 50 144  0 t = 3
rlabel pdiffusion 52 143 53 144  0 t = 4
rlabel pdiffusion 48 138 54 144 0 cell no = 56
<< m1 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2c >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< labels >>
rlabel pdiffusion 121 174 122 175  0 t = 1
rlabel pdiffusion 124 174 125 175  0 t = 2
rlabel pdiffusion 121 179 122 180  0 t = 3
rlabel pdiffusion 124 179 125 180  0 t = 4
rlabel pdiffusion 120 174 126 180 0 cell no = 57
<< m1 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2c >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< labels >>
rlabel pdiffusion 139 84 140 85  0 t = 1
rlabel pdiffusion 142 84 143 85  0 t = 2
rlabel pdiffusion 139 89 140 90  0 t = 3
rlabel pdiffusion 142 89 143 90  0 t = 4
rlabel pdiffusion 138 84 144 90 0 cell no = 58
<< m1 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2c >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 59
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 121 84 122 85  0 t = 1
rlabel pdiffusion 124 84 125 85  0 t = 2
rlabel pdiffusion 121 89 122 90  0 t = 3
rlabel pdiffusion 124 89 125 90  0 t = 4
rlabel pdiffusion 120 84 126 90 0 cell no = 60
<< m1 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2c >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< labels >>
rlabel pdiffusion 13 120 14 121  0 t = 1
rlabel pdiffusion 16 120 17 121  0 t = 2
rlabel pdiffusion 13 125 14 126  0 t = 3
rlabel pdiffusion 16 125 17 126  0 t = 4
rlabel pdiffusion 12 120 18 126 0 cell no = 61
<< m1 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2c >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 62
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 63
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 64
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 175 102 176 103  0 t = 1
rlabel pdiffusion 178 102 179 103  0 t = 2
rlabel pdiffusion 175 107 176 108  0 t = 3
rlabel pdiffusion 178 107 179 108  0 t = 4
rlabel pdiffusion 174 102 180 108 0 cell no = 65
<< m1 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2c >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 66
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 175 84 176 85  0 t = 1
rlabel pdiffusion 178 84 179 85  0 t = 2
rlabel pdiffusion 175 89 176 90  0 t = 3
rlabel pdiffusion 178 89 179 90  0 t = 4
rlabel pdiffusion 174 84 180 90 0 cell no = 67
<< m1 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2c >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< labels >>
rlabel pdiffusion 157 84 158 85  0 t = 1
rlabel pdiffusion 160 84 161 85  0 t = 2
rlabel pdiffusion 157 89 158 90  0 t = 3
rlabel pdiffusion 160 89 161 90  0 t = 4
rlabel pdiffusion 156 84 162 90 0 cell no = 68
<< m1 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2c >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 69
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 67 156 68 157  0 t = 1
rlabel pdiffusion 70 156 71 157  0 t = 2
rlabel pdiffusion 67 161 68 162  0 t = 3
rlabel pdiffusion 70 161 71 162  0 t = 4
rlabel pdiffusion 66 156 72 162 0 cell no = 70
<< m1 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2c >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 71
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 139 120 140 121  0 t = 1
rlabel pdiffusion 142 120 143 121  0 t = 2
rlabel pdiffusion 139 125 140 126  0 t = 3
rlabel pdiffusion 142 125 143 126  0 t = 4
rlabel pdiffusion 138 120 144 126 0 cell no = 72
<< m1 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2c >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< labels >>
rlabel pdiffusion 103 174 104 175  0 t = 1
rlabel pdiffusion 106 174 107 175  0 t = 2
rlabel pdiffusion 103 179 104 180  0 t = 3
rlabel pdiffusion 106 179 107 180  0 t = 4
rlabel pdiffusion 102 174 108 180 0 cell no = 73
<< m1 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2c >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 74
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 75
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 76
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 139 138 140 139  0 t = 1
rlabel pdiffusion 142 138 143 139  0 t = 2
rlabel pdiffusion 139 143 140 144  0 t = 3
rlabel pdiffusion 142 143 143 144  0 t = 4
rlabel pdiffusion 138 138 144 144 0 cell no = 77
<< m1 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2c >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< labels >>
rlabel pdiffusion 121 138 122 139  0 t = 1
rlabel pdiffusion 124 138 125 139  0 t = 2
rlabel pdiffusion 121 143 122 144  0 t = 3
rlabel pdiffusion 124 143 125 144  0 t = 4
rlabel pdiffusion 120 138 126 144 0 cell no = 78
<< m1 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2c >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< labels >>
rlabel pdiffusion 157 102 158 103  0 t = 1
rlabel pdiffusion 160 102 161 103  0 t = 2
rlabel pdiffusion 157 107 158 108  0 t = 3
rlabel pdiffusion 160 107 161 108  0 t = 4
rlabel pdiffusion 156 102 162 108 0 cell no = 79
<< m1 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2c >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< labels >>
rlabel pdiffusion 103 84 104 85  0 t = 1
rlabel pdiffusion 106 84 107 85  0 t = 2
rlabel pdiffusion 103 89 104 90  0 t = 3
rlabel pdiffusion 106 89 107 90  0 t = 4
rlabel pdiffusion 102 84 108 90 0 cell no = 80
<< m1 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2c >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< labels >>
rlabel pdiffusion 175 156 176 157  0 t = 1
rlabel pdiffusion 178 156 179 157  0 t = 2
rlabel pdiffusion 175 161 176 162  0 t = 3
rlabel pdiffusion 178 161 179 162  0 t = 4
rlabel pdiffusion 174 156 180 162 0 cell no = 81
<< m1 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2c >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< labels >>
rlabel pdiffusion 31 156 32 157  0 t = 1
rlabel pdiffusion 34 156 35 157  0 t = 2
rlabel pdiffusion 31 161 32 162  0 t = 3
rlabel pdiffusion 34 161 35 162  0 t = 4
rlabel pdiffusion 30 156 36 162 0 cell no = 82
<< m1 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2c >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< labels >>
rlabel pdiffusion 31 174 32 175  0 t = 1
rlabel pdiffusion 34 174 35 175  0 t = 2
rlabel pdiffusion 31 179 32 180  0 t = 3
rlabel pdiffusion 34 179 35 180  0 t = 4
rlabel pdiffusion 30 174 36 180 0 cell no = 83
<< m1 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2c >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< labels >>
rlabel pdiffusion 49 156 50 157  0 t = 1
rlabel pdiffusion 52 156 53 157  0 t = 2
rlabel pdiffusion 49 161 50 162  0 t = 3
rlabel pdiffusion 52 161 53 162  0 t = 4
rlabel pdiffusion 48 156 54 162 0 cell no = 84
<< m1 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2c >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< labels >>
rlabel pdiffusion 31 84 32 85  0 t = 1
rlabel pdiffusion 34 84 35 85  0 t = 2
rlabel pdiffusion 31 89 32 90  0 t = 3
rlabel pdiffusion 34 89 35 90  0 t = 4
rlabel pdiffusion 30 84 36 90 0 cell no = 85
<< m1 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2c >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< labels >>
rlabel pdiffusion 157 138 158 139  0 t = 1
rlabel pdiffusion 160 138 161 139  0 t = 2
rlabel pdiffusion 157 143 158 144  0 t = 3
rlabel pdiffusion 160 143 161 144  0 t = 4
rlabel pdiffusion 156 138 162 144 0 cell no = 86
<< m1 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2c >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< labels >>
rlabel pdiffusion 121 102 122 103  0 t = 1
rlabel pdiffusion 124 102 125 103  0 t = 2
rlabel pdiffusion 121 107 122 108  0 t = 3
rlabel pdiffusion 124 107 125 108  0 t = 4
rlabel pdiffusion 120 102 126 108 0 cell no = 87
<< m1 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2c >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< labels >>
rlabel pdiffusion 139 102 140 103  0 t = 1
rlabel pdiffusion 142 102 143 103  0 t = 2
rlabel pdiffusion 139 107 140 108  0 t = 3
rlabel pdiffusion 142 107 143 108  0 t = 4
rlabel pdiffusion 138 102 144 108 0 cell no = 88
<< m1 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2c >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< labels >>
rlabel pdiffusion 67 30 68 31  0 t = 1
rlabel pdiffusion 70 30 71 31  0 t = 2
rlabel pdiffusion 67 35 68 36  0 t = 3
rlabel pdiffusion 70 35 71 36  0 t = 4
rlabel pdiffusion 66 30 72 36 0 cell no = 89
<< m1 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2c >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< labels >>
rlabel pdiffusion 13 156 14 157  0 t = 1
rlabel pdiffusion 16 156 17 157  0 t = 2
rlabel pdiffusion 13 161 14 162  0 t = 3
rlabel pdiffusion 16 161 17 162  0 t = 4
rlabel pdiffusion 12 156 18 162 0 cell no = 90
<< m1 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2c >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< end >> 
