magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 88 10 89 11 
<< m1 >>
rect 89 10 90 11 
<< m1 >>
rect 90 10 91 11 
<< m1 >>
rect 91 10 92 11 
<< m1 >>
rect 160 10 161 11 
<< m1 >>
rect 161 10 162 11 
<< m1 >>
rect 162 10 163 11 
<< m1 >>
rect 163 10 164 11 
<< m1 >>
rect 250 10 251 11 
<< m1 >>
rect 251 10 252 11 
<< m1 >>
rect 252 10 253 11 
<< m1 >>
rect 253 10 254 11 
<< m1 >>
rect 88 11 89 12 
<< m1 >>
rect 91 11 92 12 
<< m1 >>
rect 160 11 161 12 
<< m1 >>
rect 163 11 164 12 
<< m1 >>
rect 250 11 251 12 
<< m1 >>
rect 253 11 254 12 
<< pdiffusion >>
rect 12 12 13 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< pdiffusion >>
rect 30 12 31 13 
<< pdiffusion >>
rect 31 12 32 13 
<< pdiffusion >>
rect 32 12 33 13 
<< pdiffusion >>
rect 33 12 34 13 
<< pdiffusion >>
rect 34 12 35 13 
<< pdiffusion >>
rect 35 12 36 13 
<< pdiffusion >>
rect 48 12 49 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< pdiffusion >>
rect 51 12 52 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< pdiffusion >>
rect 66 12 67 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< pdiffusion >>
rect 84 12 85 13 
<< pdiffusion >>
rect 85 12 86 13 
<< pdiffusion >>
rect 86 12 87 13 
<< pdiffusion >>
rect 87 12 88 13 
<< m1 >>
rect 88 12 89 13 
<< pdiffusion >>
rect 88 12 89 13 
<< pdiffusion >>
rect 89 12 90 13 
<< m1 >>
rect 91 12 92 13 
<< pdiffusion >>
rect 102 12 103 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< pdiffusion >>
rect 120 12 121 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< pdiffusion >>
rect 138 12 139 13 
<< pdiffusion >>
rect 139 12 140 13 
<< pdiffusion >>
rect 140 12 141 13 
<< pdiffusion >>
rect 141 12 142 13 
<< pdiffusion >>
rect 142 12 143 13 
<< pdiffusion >>
rect 143 12 144 13 
<< pdiffusion >>
rect 156 12 157 13 
<< pdiffusion >>
rect 157 12 158 13 
<< pdiffusion >>
rect 158 12 159 13 
<< pdiffusion >>
rect 159 12 160 13 
<< m1 >>
rect 160 12 161 13 
<< pdiffusion >>
rect 160 12 161 13 
<< pdiffusion >>
rect 161 12 162 13 
<< m1 >>
rect 163 12 164 13 
<< pdiffusion >>
rect 174 12 175 13 
<< pdiffusion >>
rect 175 12 176 13 
<< pdiffusion >>
rect 176 12 177 13 
<< pdiffusion >>
rect 177 12 178 13 
<< pdiffusion >>
rect 178 12 179 13 
<< pdiffusion >>
rect 179 12 180 13 
<< pdiffusion >>
rect 192 12 193 13 
<< pdiffusion >>
rect 193 12 194 13 
<< pdiffusion >>
rect 194 12 195 13 
<< pdiffusion >>
rect 195 12 196 13 
<< pdiffusion >>
rect 196 12 197 13 
<< pdiffusion >>
rect 197 12 198 13 
<< pdiffusion >>
rect 210 12 211 13 
<< pdiffusion >>
rect 211 12 212 13 
<< pdiffusion >>
rect 212 12 213 13 
<< pdiffusion >>
rect 213 12 214 13 
<< pdiffusion >>
rect 214 12 215 13 
<< pdiffusion >>
rect 215 12 216 13 
<< pdiffusion >>
rect 228 12 229 13 
<< pdiffusion >>
rect 229 12 230 13 
<< pdiffusion >>
rect 230 12 231 13 
<< pdiffusion >>
rect 231 12 232 13 
<< pdiffusion >>
rect 232 12 233 13 
<< pdiffusion >>
rect 233 12 234 13 
<< pdiffusion >>
rect 246 12 247 13 
<< pdiffusion >>
rect 247 12 248 13 
<< pdiffusion >>
rect 248 12 249 13 
<< pdiffusion >>
rect 249 12 250 13 
<< m1 >>
rect 250 12 251 13 
<< pdiffusion >>
rect 250 12 251 13 
<< pdiffusion >>
rect 251 12 252 13 
<< m1 >>
rect 253 12 254 13 
<< pdiffusion >>
rect 264 12 265 13 
<< pdiffusion >>
rect 265 12 266 13 
<< pdiffusion >>
rect 266 12 267 13 
<< pdiffusion >>
rect 267 12 268 13 
<< pdiffusion >>
rect 268 12 269 13 
<< pdiffusion >>
rect 269 12 270 13 
<< pdiffusion >>
rect 282 12 283 13 
<< pdiffusion >>
rect 283 12 284 13 
<< pdiffusion >>
rect 284 12 285 13 
<< pdiffusion >>
rect 285 12 286 13 
<< pdiffusion >>
rect 286 12 287 13 
<< pdiffusion >>
rect 287 12 288 13 
<< pdiffusion >>
rect 300 12 301 13 
<< pdiffusion >>
rect 301 12 302 13 
<< pdiffusion >>
rect 302 12 303 13 
<< pdiffusion >>
rect 303 12 304 13 
<< pdiffusion >>
rect 304 12 305 13 
<< pdiffusion >>
rect 305 12 306 13 
<< pdiffusion >>
rect 318 12 319 13 
<< pdiffusion >>
rect 319 12 320 13 
<< pdiffusion >>
rect 320 12 321 13 
<< pdiffusion >>
rect 321 12 322 13 
<< pdiffusion >>
rect 322 12 323 13 
<< pdiffusion >>
rect 323 12 324 13 
<< pdiffusion >>
rect 336 12 337 13 
<< pdiffusion >>
rect 337 12 338 13 
<< pdiffusion >>
rect 338 12 339 13 
<< pdiffusion >>
rect 339 12 340 13 
<< pdiffusion >>
rect 340 12 341 13 
<< pdiffusion >>
rect 341 12 342 13 
<< pdiffusion >>
rect 354 12 355 13 
<< pdiffusion >>
rect 355 12 356 13 
<< pdiffusion >>
rect 356 12 357 13 
<< pdiffusion >>
rect 357 12 358 13 
<< pdiffusion >>
rect 358 12 359 13 
<< pdiffusion >>
rect 359 12 360 13 
<< pdiffusion >>
rect 372 12 373 13 
<< pdiffusion >>
rect 373 12 374 13 
<< pdiffusion >>
rect 374 12 375 13 
<< pdiffusion >>
rect 375 12 376 13 
<< pdiffusion >>
rect 376 12 377 13 
<< pdiffusion >>
rect 377 12 378 13 
<< pdiffusion >>
rect 390 12 391 13 
<< pdiffusion >>
rect 391 12 392 13 
<< pdiffusion >>
rect 392 12 393 13 
<< pdiffusion >>
rect 393 12 394 13 
<< pdiffusion >>
rect 394 12 395 13 
<< pdiffusion >>
rect 395 12 396 13 
<< pdiffusion >>
rect 408 12 409 13 
<< pdiffusion >>
rect 409 12 410 13 
<< pdiffusion >>
rect 410 12 411 13 
<< pdiffusion >>
rect 411 12 412 13 
<< pdiffusion >>
rect 412 12 413 13 
<< pdiffusion >>
rect 413 12 414 13 
<< pdiffusion >>
rect 426 12 427 13 
<< pdiffusion >>
rect 427 12 428 13 
<< pdiffusion >>
rect 428 12 429 13 
<< pdiffusion >>
rect 429 12 430 13 
<< pdiffusion >>
rect 430 12 431 13 
<< pdiffusion >>
rect 431 12 432 13 
<< pdiffusion >>
rect 444 12 445 13 
<< pdiffusion >>
rect 445 12 446 13 
<< pdiffusion >>
rect 446 12 447 13 
<< pdiffusion >>
rect 447 12 448 13 
<< pdiffusion >>
rect 448 12 449 13 
<< pdiffusion >>
rect 449 12 450 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< pdiffusion >>
rect 30 13 31 14 
<< pdiffusion >>
rect 31 13 32 14 
<< pdiffusion >>
rect 32 13 33 14 
<< pdiffusion >>
rect 33 13 34 14 
<< pdiffusion >>
rect 34 13 35 14 
<< pdiffusion >>
rect 35 13 36 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< pdiffusion >>
rect 84 13 85 14 
<< pdiffusion >>
rect 85 13 86 14 
<< pdiffusion >>
rect 86 13 87 14 
<< pdiffusion >>
rect 87 13 88 14 
<< pdiffusion >>
rect 88 13 89 14 
<< pdiffusion >>
rect 89 13 90 14 
<< m1 >>
rect 91 13 92 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< pdiffusion >>
rect 138 13 139 14 
<< pdiffusion >>
rect 139 13 140 14 
<< pdiffusion >>
rect 140 13 141 14 
<< pdiffusion >>
rect 141 13 142 14 
<< pdiffusion >>
rect 142 13 143 14 
<< pdiffusion >>
rect 143 13 144 14 
<< pdiffusion >>
rect 156 13 157 14 
<< pdiffusion >>
rect 157 13 158 14 
<< pdiffusion >>
rect 158 13 159 14 
<< pdiffusion >>
rect 159 13 160 14 
<< pdiffusion >>
rect 160 13 161 14 
<< pdiffusion >>
rect 161 13 162 14 
<< m1 >>
rect 163 13 164 14 
<< pdiffusion >>
rect 174 13 175 14 
<< pdiffusion >>
rect 175 13 176 14 
<< pdiffusion >>
rect 176 13 177 14 
<< pdiffusion >>
rect 177 13 178 14 
<< pdiffusion >>
rect 178 13 179 14 
<< pdiffusion >>
rect 179 13 180 14 
<< pdiffusion >>
rect 192 13 193 14 
<< pdiffusion >>
rect 193 13 194 14 
<< pdiffusion >>
rect 194 13 195 14 
<< pdiffusion >>
rect 195 13 196 14 
<< pdiffusion >>
rect 196 13 197 14 
<< pdiffusion >>
rect 197 13 198 14 
<< pdiffusion >>
rect 210 13 211 14 
<< pdiffusion >>
rect 211 13 212 14 
<< pdiffusion >>
rect 212 13 213 14 
<< pdiffusion >>
rect 213 13 214 14 
<< pdiffusion >>
rect 214 13 215 14 
<< pdiffusion >>
rect 215 13 216 14 
<< pdiffusion >>
rect 228 13 229 14 
<< pdiffusion >>
rect 229 13 230 14 
<< pdiffusion >>
rect 230 13 231 14 
<< pdiffusion >>
rect 231 13 232 14 
<< pdiffusion >>
rect 232 13 233 14 
<< pdiffusion >>
rect 233 13 234 14 
<< pdiffusion >>
rect 246 13 247 14 
<< pdiffusion >>
rect 247 13 248 14 
<< pdiffusion >>
rect 248 13 249 14 
<< pdiffusion >>
rect 249 13 250 14 
<< pdiffusion >>
rect 250 13 251 14 
<< pdiffusion >>
rect 251 13 252 14 
<< m1 >>
rect 253 13 254 14 
<< pdiffusion >>
rect 264 13 265 14 
<< pdiffusion >>
rect 265 13 266 14 
<< pdiffusion >>
rect 266 13 267 14 
<< pdiffusion >>
rect 267 13 268 14 
<< pdiffusion >>
rect 268 13 269 14 
<< pdiffusion >>
rect 269 13 270 14 
<< pdiffusion >>
rect 282 13 283 14 
<< pdiffusion >>
rect 283 13 284 14 
<< pdiffusion >>
rect 284 13 285 14 
<< pdiffusion >>
rect 285 13 286 14 
<< pdiffusion >>
rect 286 13 287 14 
<< pdiffusion >>
rect 287 13 288 14 
<< pdiffusion >>
rect 300 13 301 14 
<< pdiffusion >>
rect 301 13 302 14 
<< pdiffusion >>
rect 302 13 303 14 
<< pdiffusion >>
rect 303 13 304 14 
<< pdiffusion >>
rect 304 13 305 14 
<< pdiffusion >>
rect 305 13 306 14 
<< pdiffusion >>
rect 318 13 319 14 
<< pdiffusion >>
rect 319 13 320 14 
<< pdiffusion >>
rect 320 13 321 14 
<< pdiffusion >>
rect 321 13 322 14 
<< pdiffusion >>
rect 322 13 323 14 
<< pdiffusion >>
rect 323 13 324 14 
<< pdiffusion >>
rect 336 13 337 14 
<< pdiffusion >>
rect 337 13 338 14 
<< pdiffusion >>
rect 338 13 339 14 
<< pdiffusion >>
rect 339 13 340 14 
<< pdiffusion >>
rect 340 13 341 14 
<< pdiffusion >>
rect 341 13 342 14 
<< pdiffusion >>
rect 354 13 355 14 
<< pdiffusion >>
rect 355 13 356 14 
<< pdiffusion >>
rect 356 13 357 14 
<< pdiffusion >>
rect 357 13 358 14 
<< pdiffusion >>
rect 358 13 359 14 
<< pdiffusion >>
rect 359 13 360 14 
<< pdiffusion >>
rect 372 13 373 14 
<< pdiffusion >>
rect 373 13 374 14 
<< pdiffusion >>
rect 374 13 375 14 
<< pdiffusion >>
rect 375 13 376 14 
<< pdiffusion >>
rect 376 13 377 14 
<< pdiffusion >>
rect 377 13 378 14 
<< pdiffusion >>
rect 390 13 391 14 
<< pdiffusion >>
rect 391 13 392 14 
<< pdiffusion >>
rect 392 13 393 14 
<< pdiffusion >>
rect 393 13 394 14 
<< pdiffusion >>
rect 394 13 395 14 
<< pdiffusion >>
rect 395 13 396 14 
<< pdiffusion >>
rect 408 13 409 14 
<< pdiffusion >>
rect 409 13 410 14 
<< pdiffusion >>
rect 410 13 411 14 
<< pdiffusion >>
rect 411 13 412 14 
<< pdiffusion >>
rect 412 13 413 14 
<< pdiffusion >>
rect 413 13 414 14 
<< pdiffusion >>
rect 426 13 427 14 
<< pdiffusion >>
rect 427 13 428 14 
<< pdiffusion >>
rect 428 13 429 14 
<< pdiffusion >>
rect 429 13 430 14 
<< pdiffusion >>
rect 430 13 431 14 
<< pdiffusion >>
rect 431 13 432 14 
<< pdiffusion >>
rect 444 13 445 14 
<< pdiffusion >>
rect 445 13 446 14 
<< pdiffusion >>
rect 446 13 447 14 
<< pdiffusion >>
rect 447 13 448 14 
<< pdiffusion >>
rect 448 13 449 14 
<< pdiffusion >>
rect 449 13 450 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< pdiffusion >>
rect 30 14 31 15 
<< pdiffusion >>
rect 31 14 32 15 
<< pdiffusion >>
rect 32 14 33 15 
<< pdiffusion >>
rect 33 14 34 15 
<< pdiffusion >>
rect 34 14 35 15 
<< pdiffusion >>
rect 35 14 36 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< pdiffusion >>
rect 84 14 85 15 
<< pdiffusion >>
rect 85 14 86 15 
<< pdiffusion >>
rect 86 14 87 15 
<< pdiffusion >>
rect 87 14 88 15 
<< pdiffusion >>
rect 88 14 89 15 
<< pdiffusion >>
rect 89 14 90 15 
<< m1 >>
rect 91 14 92 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< pdiffusion >>
rect 138 14 139 15 
<< pdiffusion >>
rect 139 14 140 15 
<< pdiffusion >>
rect 140 14 141 15 
<< pdiffusion >>
rect 141 14 142 15 
<< pdiffusion >>
rect 142 14 143 15 
<< pdiffusion >>
rect 143 14 144 15 
<< pdiffusion >>
rect 156 14 157 15 
<< pdiffusion >>
rect 157 14 158 15 
<< pdiffusion >>
rect 158 14 159 15 
<< pdiffusion >>
rect 159 14 160 15 
<< pdiffusion >>
rect 160 14 161 15 
<< pdiffusion >>
rect 161 14 162 15 
<< m1 >>
rect 163 14 164 15 
<< pdiffusion >>
rect 174 14 175 15 
<< pdiffusion >>
rect 175 14 176 15 
<< pdiffusion >>
rect 176 14 177 15 
<< pdiffusion >>
rect 177 14 178 15 
<< pdiffusion >>
rect 178 14 179 15 
<< pdiffusion >>
rect 179 14 180 15 
<< pdiffusion >>
rect 192 14 193 15 
<< pdiffusion >>
rect 193 14 194 15 
<< pdiffusion >>
rect 194 14 195 15 
<< pdiffusion >>
rect 195 14 196 15 
<< pdiffusion >>
rect 196 14 197 15 
<< pdiffusion >>
rect 197 14 198 15 
<< pdiffusion >>
rect 210 14 211 15 
<< pdiffusion >>
rect 211 14 212 15 
<< pdiffusion >>
rect 212 14 213 15 
<< pdiffusion >>
rect 213 14 214 15 
<< pdiffusion >>
rect 214 14 215 15 
<< pdiffusion >>
rect 215 14 216 15 
<< pdiffusion >>
rect 228 14 229 15 
<< pdiffusion >>
rect 229 14 230 15 
<< pdiffusion >>
rect 230 14 231 15 
<< pdiffusion >>
rect 231 14 232 15 
<< pdiffusion >>
rect 232 14 233 15 
<< pdiffusion >>
rect 233 14 234 15 
<< pdiffusion >>
rect 246 14 247 15 
<< pdiffusion >>
rect 247 14 248 15 
<< pdiffusion >>
rect 248 14 249 15 
<< pdiffusion >>
rect 249 14 250 15 
<< pdiffusion >>
rect 250 14 251 15 
<< pdiffusion >>
rect 251 14 252 15 
<< m1 >>
rect 253 14 254 15 
<< pdiffusion >>
rect 264 14 265 15 
<< pdiffusion >>
rect 265 14 266 15 
<< pdiffusion >>
rect 266 14 267 15 
<< pdiffusion >>
rect 267 14 268 15 
<< pdiffusion >>
rect 268 14 269 15 
<< pdiffusion >>
rect 269 14 270 15 
<< pdiffusion >>
rect 282 14 283 15 
<< pdiffusion >>
rect 283 14 284 15 
<< pdiffusion >>
rect 284 14 285 15 
<< pdiffusion >>
rect 285 14 286 15 
<< pdiffusion >>
rect 286 14 287 15 
<< pdiffusion >>
rect 287 14 288 15 
<< pdiffusion >>
rect 300 14 301 15 
<< pdiffusion >>
rect 301 14 302 15 
<< pdiffusion >>
rect 302 14 303 15 
<< pdiffusion >>
rect 303 14 304 15 
<< pdiffusion >>
rect 304 14 305 15 
<< pdiffusion >>
rect 305 14 306 15 
<< pdiffusion >>
rect 318 14 319 15 
<< pdiffusion >>
rect 319 14 320 15 
<< pdiffusion >>
rect 320 14 321 15 
<< pdiffusion >>
rect 321 14 322 15 
<< pdiffusion >>
rect 322 14 323 15 
<< pdiffusion >>
rect 323 14 324 15 
<< pdiffusion >>
rect 336 14 337 15 
<< pdiffusion >>
rect 337 14 338 15 
<< pdiffusion >>
rect 338 14 339 15 
<< pdiffusion >>
rect 339 14 340 15 
<< pdiffusion >>
rect 340 14 341 15 
<< pdiffusion >>
rect 341 14 342 15 
<< pdiffusion >>
rect 354 14 355 15 
<< pdiffusion >>
rect 355 14 356 15 
<< pdiffusion >>
rect 356 14 357 15 
<< pdiffusion >>
rect 357 14 358 15 
<< pdiffusion >>
rect 358 14 359 15 
<< pdiffusion >>
rect 359 14 360 15 
<< pdiffusion >>
rect 372 14 373 15 
<< pdiffusion >>
rect 373 14 374 15 
<< pdiffusion >>
rect 374 14 375 15 
<< pdiffusion >>
rect 375 14 376 15 
<< pdiffusion >>
rect 376 14 377 15 
<< pdiffusion >>
rect 377 14 378 15 
<< pdiffusion >>
rect 390 14 391 15 
<< pdiffusion >>
rect 391 14 392 15 
<< pdiffusion >>
rect 392 14 393 15 
<< pdiffusion >>
rect 393 14 394 15 
<< pdiffusion >>
rect 394 14 395 15 
<< pdiffusion >>
rect 395 14 396 15 
<< pdiffusion >>
rect 408 14 409 15 
<< pdiffusion >>
rect 409 14 410 15 
<< pdiffusion >>
rect 410 14 411 15 
<< pdiffusion >>
rect 411 14 412 15 
<< pdiffusion >>
rect 412 14 413 15 
<< pdiffusion >>
rect 413 14 414 15 
<< pdiffusion >>
rect 426 14 427 15 
<< pdiffusion >>
rect 427 14 428 15 
<< pdiffusion >>
rect 428 14 429 15 
<< pdiffusion >>
rect 429 14 430 15 
<< pdiffusion >>
rect 430 14 431 15 
<< pdiffusion >>
rect 431 14 432 15 
<< pdiffusion >>
rect 444 14 445 15 
<< pdiffusion >>
rect 445 14 446 15 
<< pdiffusion >>
rect 446 14 447 15 
<< pdiffusion >>
rect 447 14 448 15 
<< pdiffusion >>
rect 448 14 449 15 
<< pdiffusion >>
rect 449 14 450 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< pdiffusion >>
rect 30 15 31 16 
<< pdiffusion >>
rect 31 15 32 16 
<< pdiffusion >>
rect 32 15 33 16 
<< pdiffusion >>
rect 33 15 34 16 
<< pdiffusion >>
rect 34 15 35 16 
<< pdiffusion >>
rect 35 15 36 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< pdiffusion >>
rect 84 15 85 16 
<< pdiffusion >>
rect 85 15 86 16 
<< pdiffusion >>
rect 86 15 87 16 
<< pdiffusion >>
rect 87 15 88 16 
<< pdiffusion >>
rect 88 15 89 16 
<< pdiffusion >>
rect 89 15 90 16 
<< m1 >>
rect 91 15 92 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< pdiffusion >>
rect 138 15 139 16 
<< pdiffusion >>
rect 139 15 140 16 
<< pdiffusion >>
rect 140 15 141 16 
<< pdiffusion >>
rect 141 15 142 16 
<< pdiffusion >>
rect 142 15 143 16 
<< pdiffusion >>
rect 143 15 144 16 
<< pdiffusion >>
rect 156 15 157 16 
<< pdiffusion >>
rect 157 15 158 16 
<< pdiffusion >>
rect 158 15 159 16 
<< pdiffusion >>
rect 159 15 160 16 
<< pdiffusion >>
rect 160 15 161 16 
<< pdiffusion >>
rect 161 15 162 16 
<< m1 >>
rect 163 15 164 16 
<< pdiffusion >>
rect 174 15 175 16 
<< pdiffusion >>
rect 175 15 176 16 
<< pdiffusion >>
rect 176 15 177 16 
<< pdiffusion >>
rect 177 15 178 16 
<< pdiffusion >>
rect 178 15 179 16 
<< pdiffusion >>
rect 179 15 180 16 
<< pdiffusion >>
rect 192 15 193 16 
<< pdiffusion >>
rect 193 15 194 16 
<< pdiffusion >>
rect 194 15 195 16 
<< pdiffusion >>
rect 195 15 196 16 
<< pdiffusion >>
rect 196 15 197 16 
<< pdiffusion >>
rect 197 15 198 16 
<< pdiffusion >>
rect 210 15 211 16 
<< pdiffusion >>
rect 211 15 212 16 
<< pdiffusion >>
rect 212 15 213 16 
<< pdiffusion >>
rect 213 15 214 16 
<< pdiffusion >>
rect 214 15 215 16 
<< pdiffusion >>
rect 215 15 216 16 
<< pdiffusion >>
rect 228 15 229 16 
<< pdiffusion >>
rect 229 15 230 16 
<< pdiffusion >>
rect 230 15 231 16 
<< pdiffusion >>
rect 231 15 232 16 
<< pdiffusion >>
rect 232 15 233 16 
<< pdiffusion >>
rect 233 15 234 16 
<< pdiffusion >>
rect 246 15 247 16 
<< pdiffusion >>
rect 247 15 248 16 
<< pdiffusion >>
rect 248 15 249 16 
<< pdiffusion >>
rect 249 15 250 16 
<< pdiffusion >>
rect 250 15 251 16 
<< pdiffusion >>
rect 251 15 252 16 
<< m1 >>
rect 253 15 254 16 
<< pdiffusion >>
rect 264 15 265 16 
<< pdiffusion >>
rect 265 15 266 16 
<< pdiffusion >>
rect 266 15 267 16 
<< pdiffusion >>
rect 267 15 268 16 
<< pdiffusion >>
rect 268 15 269 16 
<< pdiffusion >>
rect 269 15 270 16 
<< pdiffusion >>
rect 282 15 283 16 
<< pdiffusion >>
rect 283 15 284 16 
<< pdiffusion >>
rect 284 15 285 16 
<< pdiffusion >>
rect 285 15 286 16 
<< pdiffusion >>
rect 286 15 287 16 
<< pdiffusion >>
rect 287 15 288 16 
<< pdiffusion >>
rect 300 15 301 16 
<< pdiffusion >>
rect 301 15 302 16 
<< pdiffusion >>
rect 302 15 303 16 
<< pdiffusion >>
rect 303 15 304 16 
<< pdiffusion >>
rect 304 15 305 16 
<< pdiffusion >>
rect 305 15 306 16 
<< pdiffusion >>
rect 318 15 319 16 
<< pdiffusion >>
rect 319 15 320 16 
<< pdiffusion >>
rect 320 15 321 16 
<< pdiffusion >>
rect 321 15 322 16 
<< pdiffusion >>
rect 322 15 323 16 
<< pdiffusion >>
rect 323 15 324 16 
<< pdiffusion >>
rect 336 15 337 16 
<< pdiffusion >>
rect 337 15 338 16 
<< pdiffusion >>
rect 338 15 339 16 
<< pdiffusion >>
rect 339 15 340 16 
<< pdiffusion >>
rect 340 15 341 16 
<< pdiffusion >>
rect 341 15 342 16 
<< pdiffusion >>
rect 354 15 355 16 
<< pdiffusion >>
rect 355 15 356 16 
<< pdiffusion >>
rect 356 15 357 16 
<< pdiffusion >>
rect 357 15 358 16 
<< pdiffusion >>
rect 358 15 359 16 
<< pdiffusion >>
rect 359 15 360 16 
<< pdiffusion >>
rect 372 15 373 16 
<< pdiffusion >>
rect 373 15 374 16 
<< pdiffusion >>
rect 374 15 375 16 
<< pdiffusion >>
rect 375 15 376 16 
<< pdiffusion >>
rect 376 15 377 16 
<< pdiffusion >>
rect 377 15 378 16 
<< pdiffusion >>
rect 390 15 391 16 
<< pdiffusion >>
rect 391 15 392 16 
<< pdiffusion >>
rect 392 15 393 16 
<< pdiffusion >>
rect 393 15 394 16 
<< pdiffusion >>
rect 394 15 395 16 
<< pdiffusion >>
rect 395 15 396 16 
<< pdiffusion >>
rect 408 15 409 16 
<< pdiffusion >>
rect 409 15 410 16 
<< pdiffusion >>
rect 410 15 411 16 
<< pdiffusion >>
rect 411 15 412 16 
<< pdiffusion >>
rect 412 15 413 16 
<< pdiffusion >>
rect 413 15 414 16 
<< pdiffusion >>
rect 426 15 427 16 
<< pdiffusion >>
rect 427 15 428 16 
<< pdiffusion >>
rect 428 15 429 16 
<< pdiffusion >>
rect 429 15 430 16 
<< pdiffusion >>
rect 430 15 431 16 
<< pdiffusion >>
rect 431 15 432 16 
<< pdiffusion >>
rect 444 15 445 16 
<< pdiffusion >>
rect 445 15 446 16 
<< pdiffusion >>
rect 446 15 447 16 
<< pdiffusion >>
rect 447 15 448 16 
<< pdiffusion >>
rect 448 15 449 16 
<< pdiffusion >>
rect 449 15 450 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< pdiffusion >>
rect 30 16 31 17 
<< pdiffusion >>
rect 31 16 32 17 
<< pdiffusion >>
rect 32 16 33 17 
<< pdiffusion >>
rect 33 16 34 17 
<< pdiffusion >>
rect 34 16 35 17 
<< pdiffusion >>
rect 35 16 36 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< pdiffusion >>
rect 84 16 85 17 
<< pdiffusion >>
rect 85 16 86 17 
<< pdiffusion >>
rect 86 16 87 17 
<< pdiffusion >>
rect 87 16 88 17 
<< pdiffusion >>
rect 88 16 89 17 
<< pdiffusion >>
rect 89 16 90 17 
<< m1 >>
rect 91 16 92 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< pdiffusion >>
rect 138 16 139 17 
<< pdiffusion >>
rect 139 16 140 17 
<< pdiffusion >>
rect 140 16 141 17 
<< pdiffusion >>
rect 141 16 142 17 
<< pdiffusion >>
rect 142 16 143 17 
<< pdiffusion >>
rect 143 16 144 17 
<< pdiffusion >>
rect 156 16 157 17 
<< pdiffusion >>
rect 157 16 158 17 
<< pdiffusion >>
rect 158 16 159 17 
<< pdiffusion >>
rect 159 16 160 17 
<< pdiffusion >>
rect 160 16 161 17 
<< pdiffusion >>
rect 161 16 162 17 
<< m1 >>
rect 163 16 164 17 
<< pdiffusion >>
rect 174 16 175 17 
<< pdiffusion >>
rect 175 16 176 17 
<< pdiffusion >>
rect 176 16 177 17 
<< pdiffusion >>
rect 177 16 178 17 
<< pdiffusion >>
rect 178 16 179 17 
<< pdiffusion >>
rect 179 16 180 17 
<< pdiffusion >>
rect 192 16 193 17 
<< pdiffusion >>
rect 193 16 194 17 
<< pdiffusion >>
rect 194 16 195 17 
<< pdiffusion >>
rect 195 16 196 17 
<< pdiffusion >>
rect 196 16 197 17 
<< pdiffusion >>
rect 197 16 198 17 
<< pdiffusion >>
rect 210 16 211 17 
<< pdiffusion >>
rect 211 16 212 17 
<< pdiffusion >>
rect 212 16 213 17 
<< pdiffusion >>
rect 213 16 214 17 
<< pdiffusion >>
rect 214 16 215 17 
<< pdiffusion >>
rect 215 16 216 17 
<< pdiffusion >>
rect 228 16 229 17 
<< pdiffusion >>
rect 229 16 230 17 
<< pdiffusion >>
rect 230 16 231 17 
<< pdiffusion >>
rect 231 16 232 17 
<< pdiffusion >>
rect 232 16 233 17 
<< pdiffusion >>
rect 233 16 234 17 
<< pdiffusion >>
rect 246 16 247 17 
<< pdiffusion >>
rect 247 16 248 17 
<< pdiffusion >>
rect 248 16 249 17 
<< pdiffusion >>
rect 249 16 250 17 
<< pdiffusion >>
rect 250 16 251 17 
<< pdiffusion >>
rect 251 16 252 17 
<< m1 >>
rect 253 16 254 17 
<< pdiffusion >>
rect 264 16 265 17 
<< pdiffusion >>
rect 265 16 266 17 
<< pdiffusion >>
rect 266 16 267 17 
<< pdiffusion >>
rect 267 16 268 17 
<< pdiffusion >>
rect 268 16 269 17 
<< pdiffusion >>
rect 269 16 270 17 
<< pdiffusion >>
rect 282 16 283 17 
<< pdiffusion >>
rect 283 16 284 17 
<< pdiffusion >>
rect 284 16 285 17 
<< pdiffusion >>
rect 285 16 286 17 
<< pdiffusion >>
rect 286 16 287 17 
<< pdiffusion >>
rect 287 16 288 17 
<< pdiffusion >>
rect 300 16 301 17 
<< pdiffusion >>
rect 301 16 302 17 
<< pdiffusion >>
rect 302 16 303 17 
<< pdiffusion >>
rect 303 16 304 17 
<< pdiffusion >>
rect 304 16 305 17 
<< pdiffusion >>
rect 305 16 306 17 
<< pdiffusion >>
rect 318 16 319 17 
<< pdiffusion >>
rect 319 16 320 17 
<< pdiffusion >>
rect 320 16 321 17 
<< pdiffusion >>
rect 321 16 322 17 
<< pdiffusion >>
rect 322 16 323 17 
<< pdiffusion >>
rect 323 16 324 17 
<< pdiffusion >>
rect 336 16 337 17 
<< pdiffusion >>
rect 337 16 338 17 
<< pdiffusion >>
rect 338 16 339 17 
<< pdiffusion >>
rect 339 16 340 17 
<< pdiffusion >>
rect 340 16 341 17 
<< pdiffusion >>
rect 341 16 342 17 
<< pdiffusion >>
rect 354 16 355 17 
<< pdiffusion >>
rect 355 16 356 17 
<< pdiffusion >>
rect 356 16 357 17 
<< pdiffusion >>
rect 357 16 358 17 
<< pdiffusion >>
rect 358 16 359 17 
<< pdiffusion >>
rect 359 16 360 17 
<< pdiffusion >>
rect 372 16 373 17 
<< pdiffusion >>
rect 373 16 374 17 
<< pdiffusion >>
rect 374 16 375 17 
<< pdiffusion >>
rect 375 16 376 17 
<< pdiffusion >>
rect 376 16 377 17 
<< pdiffusion >>
rect 377 16 378 17 
<< pdiffusion >>
rect 390 16 391 17 
<< pdiffusion >>
rect 391 16 392 17 
<< pdiffusion >>
rect 392 16 393 17 
<< pdiffusion >>
rect 393 16 394 17 
<< pdiffusion >>
rect 394 16 395 17 
<< pdiffusion >>
rect 395 16 396 17 
<< pdiffusion >>
rect 408 16 409 17 
<< pdiffusion >>
rect 409 16 410 17 
<< pdiffusion >>
rect 410 16 411 17 
<< pdiffusion >>
rect 411 16 412 17 
<< pdiffusion >>
rect 412 16 413 17 
<< pdiffusion >>
rect 413 16 414 17 
<< pdiffusion >>
rect 426 16 427 17 
<< pdiffusion >>
rect 427 16 428 17 
<< pdiffusion >>
rect 428 16 429 17 
<< pdiffusion >>
rect 429 16 430 17 
<< pdiffusion >>
rect 430 16 431 17 
<< pdiffusion >>
rect 431 16 432 17 
<< pdiffusion >>
rect 444 16 445 17 
<< pdiffusion >>
rect 445 16 446 17 
<< pdiffusion >>
rect 446 16 447 17 
<< pdiffusion >>
rect 447 16 448 17 
<< pdiffusion >>
rect 448 16 449 17 
<< pdiffusion >>
rect 449 16 450 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< pdiffusion >>
rect 30 17 31 18 
<< pdiffusion >>
rect 31 17 32 18 
<< pdiffusion >>
rect 32 17 33 18 
<< pdiffusion >>
rect 33 17 34 18 
<< pdiffusion >>
rect 34 17 35 18 
<< pdiffusion >>
rect 35 17 36 18 
<< pdiffusion >>
rect 48 17 49 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< pdiffusion >>
rect 66 17 67 18 
<< m1 >>
rect 67 17 68 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< pdiffusion >>
rect 84 17 85 18 
<< pdiffusion >>
rect 85 17 86 18 
<< pdiffusion >>
rect 86 17 87 18 
<< pdiffusion >>
rect 87 17 88 18 
<< pdiffusion >>
rect 88 17 89 18 
<< pdiffusion >>
rect 89 17 90 18 
<< m1 >>
rect 91 17 92 18 
<< pdiffusion >>
rect 102 17 103 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< pdiffusion >>
rect 120 17 121 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< pdiffusion >>
rect 138 17 139 18 
<< pdiffusion >>
rect 139 17 140 18 
<< pdiffusion >>
rect 140 17 141 18 
<< pdiffusion >>
rect 141 17 142 18 
<< pdiffusion >>
rect 142 17 143 18 
<< pdiffusion >>
rect 143 17 144 18 
<< pdiffusion >>
rect 156 17 157 18 
<< pdiffusion >>
rect 157 17 158 18 
<< pdiffusion >>
rect 158 17 159 18 
<< pdiffusion >>
rect 159 17 160 18 
<< pdiffusion >>
rect 160 17 161 18 
<< pdiffusion >>
rect 161 17 162 18 
<< m1 >>
rect 163 17 164 18 
<< pdiffusion >>
rect 174 17 175 18 
<< pdiffusion >>
rect 175 17 176 18 
<< pdiffusion >>
rect 176 17 177 18 
<< pdiffusion >>
rect 177 17 178 18 
<< pdiffusion >>
rect 178 17 179 18 
<< pdiffusion >>
rect 179 17 180 18 
<< pdiffusion >>
rect 192 17 193 18 
<< pdiffusion >>
rect 193 17 194 18 
<< pdiffusion >>
rect 194 17 195 18 
<< pdiffusion >>
rect 195 17 196 18 
<< pdiffusion >>
rect 196 17 197 18 
<< pdiffusion >>
rect 197 17 198 18 
<< pdiffusion >>
rect 210 17 211 18 
<< pdiffusion >>
rect 211 17 212 18 
<< pdiffusion >>
rect 212 17 213 18 
<< pdiffusion >>
rect 213 17 214 18 
<< pdiffusion >>
rect 214 17 215 18 
<< pdiffusion >>
rect 215 17 216 18 
<< pdiffusion >>
rect 228 17 229 18 
<< pdiffusion >>
rect 229 17 230 18 
<< pdiffusion >>
rect 230 17 231 18 
<< pdiffusion >>
rect 231 17 232 18 
<< pdiffusion >>
rect 232 17 233 18 
<< pdiffusion >>
rect 233 17 234 18 
<< pdiffusion >>
rect 246 17 247 18 
<< m1 >>
rect 247 17 248 18 
<< pdiffusion >>
rect 247 17 248 18 
<< pdiffusion >>
rect 248 17 249 18 
<< pdiffusion >>
rect 249 17 250 18 
<< pdiffusion >>
rect 250 17 251 18 
<< pdiffusion >>
rect 251 17 252 18 
<< m1 >>
rect 253 17 254 18 
<< pdiffusion >>
rect 264 17 265 18 
<< pdiffusion >>
rect 265 17 266 18 
<< pdiffusion >>
rect 266 17 267 18 
<< pdiffusion >>
rect 267 17 268 18 
<< m1 >>
rect 268 17 269 18 
<< pdiffusion >>
rect 268 17 269 18 
<< pdiffusion >>
rect 269 17 270 18 
<< pdiffusion >>
rect 282 17 283 18 
<< pdiffusion >>
rect 283 17 284 18 
<< pdiffusion >>
rect 284 17 285 18 
<< pdiffusion >>
rect 285 17 286 18 
<< pdiffusion >>
rect 286 17 287 18 
<< pdiffusion >>
rect 287 17 288 18 
<< pdiffusion >>
rect 300 17 301 18 
<< pdiffusion >>
rect 301 17 302 18 
<< pdiffusion >>
rect 302 17 303 18 
<< pdiffusion >>
rect 303 17 304 18 
<< pdiffusion >>
rect 304 17 305 18 
<< pdiffusion >>
rect 305 17 306 18 
<< pdiffusion >>
rect 318 17 319 18 
<< pdiffusion >>
rect 319 17 320 18 
<< pdiffusion >>
rect 320 17 321 18 
<< pdiffusion >>
rect 321 17 322 18 
<< pdiffusion >>
rect 322 17 323 18 
<< pdiffusion >>
rect 323 17 324 18 
<< pdiffusion >>
rect 336 17 337 18 
<< pdiffusion >>
rect 337 17 338 18 
<< pdiffusion >>
rect 338 17 339 18 
<< pdiffusion >>
rect 339 17 340 18 
<< pdiffusion >>
rect 340 17 341 18 
<< pdiffusion >>
rect 341 17 342 18 
<< pdiffusion >>
rect 354 17 355 18 
<< pdiffusion >>
rect 355 17 356 18 
<< pdiffusion >>
rect 356 17 357 18 
<< pdiffusion >>
rect 357 17 358 18 
<< pdiffusion >>
rect 358 17 359 18 
<< pdiffusion >>
rect 359 17 360 18 
<< pdiffusion >>
rect 372 17 373 18 
<< pdiffusion >>
rect 373 17 374 18 
<< pdiffusion >>
rect 374 17 375 18 
<< pdiffusion >>
rect 375 17 376 18 
<< pdiffusion >>
rect 376 17 377 18 
<< pdiffusion >>
rect 377 17 378 18 
<< pdiffusion >>
rect 390 17 391 18 
<< pdiffusion >>
rect 391 17 392 18 
<< pdiffusion >>
rect 392 17 393 18 
<< pdiffusion >>
rect 393 17 394 18 
<< pdiffusion >>
rect 394 17 395 18 
<< pdiffusion >>
rect 395 17 396 18 
<< pdiffusion >>
rect 408 17 409 18 
<< pdiffusion >>
rect 409 17 410 18 
<< pdiffusion >>
rect 410 17 411 18 
<< pdiffusion >>
rect 411 17 412 18 
<< pdiffusion >>
rect 412 17 413 18 
<< pdiffusion >>
rect 413 17 414 18 
<< pdiffusion >>
rect 426 17 427 18 
<< pdiffusion >>
rect 427 17 428 18 
<< pdiffusion >>
rect 428 17 429 18 
<< pdiffusion >>
rect 429 17 430 18 
<< pdiffusion >>
rect 430 17 431 18 
<< pdiffusion >>
rect 431 17 432 18 
<< pdiffusion >>
rect 444 17 445 18 
<< pdiffusion >>
rect 445 17 446 18 
<< pdiffusion >>
rect 446 17 447 18 
<< pdiffusion >>
rect 447 17 448 18 
<< m1 >>
rect 448 17 449 18 
<< pdiffusion >>
rect 448 17 449 18 
<< pdiffusion >>
rect 449 17 450 18 
<< m1 >>
rect 67 18 68 19 
<< m1 >>
rect 91 18 92 19 
<< m1 >>
rect 163 18 164 19 
<< m1 >>
rect 247 18 248 19 
<< m1 >>
rect 253 18 254 19 
<< m1 >>
rect 268 18 269 19 
<< m1 >>
rect 448 18 449 19 
<< m1 >>
rect 67 19 68 20 
<< m1 >>
rect 91 19 92 20 
<< m1 >>
rect 163 19 164 20 
<< m1 >>
rect 244 19 245 20 
<< m1 >>
rect 245 19 246 20 
<< m1 >>
rect 246 19 247 20 
<< m1 >>
rect 247 19 248 20 
<< m1 >>
rect 253 19 254 20 
<< m1 >>
rect 268 19 269 20 
<< m1 >>
rect 448 19 449 20 
<< m1 >>
rect 67 20 68 21 
<< m1 >>
rect 91 20 92 21 
<< m1 >>
rect 163 20 164 21 
<< m1 >>
rect 244 20 245 21 
<< m1 >>
rect 253 20 254 21 
<< m1 >>
rect 268 20 269 21 
<< m1 >>
rect 448 20 449 21 
<< m1 >>
rect 67 21 68 22 
<< m1 >>
rect 91 21 92 22 
<< m1 >>
rect 163 21 164 22 
<< m1 >>
rect 244 21 245 22 
<< m1 >>
rect 253 21 254 22 
<< m1 >>
rect 268 21 269 22 
<< m1 >>
rect 448 21 449 22 
<< m1 >>
rect 67 22 68 23 
<< m1 >>
rect 91 22 92 23 
<< m1 >>
rect 163 22 164 23 
<< m1 >>
rect 244 22 245 23 
<< m1 >>
rect 253 22 254 23 
<< m1 >>
rect 268 22 269 23 
<< m1 >>
rect 442 22 443 23 
<< m1 >>
rect 443 22 444 23 
<< m1 >>
rect 444 22 445 23 
<< m1 >>
rect 445 22 446 23 
<< m1 >>
rect 446 22 447 23 
<< m1 >>
rect 447 22 448 23 
<< m1 >>
rect 448 22 449 23 
<< m1 >>
rect 67 23 68 24 
<< m1 >>
rect 91 23 92 24 
<< m1 >>
rect 163 23 164 24 
<< m1 >>
rect 244 23 245 24 
<< m1 >>
rect 253 23 254 24 
<< m1 >>
rect 268 23 269 24 
<< m2 >>
rect 268 23 269 24 
<< m2c >>
rect 268 23 269 24 
<< m1 >>
rect 268 23 269 24 
<< m2 >>
rect 268 23 269 24 
<< m1 >>
rect 442 23 443 24 
<< m1 >>
rect 67 24 68 25 
<< m1 >>
rect 91 24 92 25 
<< m1 >>
rect 163 24 164 25 
<< m1 >>
rect 244 24 245 25 
<< m1 >>
rect 253 24 254 25 
<< m2 >>
rect 264 24 265 25 
<< m2 >>
rect 265 24 266 25 
<< m2 >>
rect 266 24 267 25 
<< m2 >>
rect 267 24 268 25 
<< m2 >>
rect 268 24 269 25 
<< m1 >>
rect 442 24 443 25 
<< m1 >>
rect 64 25 65 26 
<< m1 >>
rect 65 25 66 26 
<< m1 >>
rect 66 25 67 26 
<< m1 >>
rect 67 25 68 26 
<< m1 >>
rect 91 25 92 26 
<< m1 >>
rect 163 25 164 26 
<< m1 >>
rect 244 25 245 26 
<< m1 >>
rect 253 25 254 26 
<< m2 >>
rect 254 25 255 26 
<< m1 >>
rect 255 25 256 26 
<< m2 >>
rect 255 25 256 26 
<< m2c >>
rect 255 25 256 26 
<< m1 >>
rect 255 25 256 26 
<< m2 >>
rect 255 25 256 26 
<< m1 >>
rect 256 25 257 26 
<< m1 >>
rect 257 25 258 26 
<< m1 >>
rect 258 25 259 26 
<< m1 >>
rect 259 25 260 26 
<< m1 >>
rect 260 25 261 26 
<< m1 >>
rect 261 25 262 26 
<< m1 >>
rect 262 25 263 26 
<< m1 >>
rect 263 25 264 26 
<< m1 >>
rect 264 25 265 26 
<< m2 >>
rect 264 25 265 26 
<< m1 >>
rect 265 25 266 26 
<< m1 >>
rect 266 25 267 26 
<< m1 >>
rect 267 25 268 26 
<< m1 >>
rect 268 25 269 26 
<< m1 >>
rect 442 25 443 26 
<< m1 >>
rect 64 26 65 27 
<< m1 >>
rect 91 26 92 27 
<< m1 >>
rect 163 26 164 27 
<< m1 >>
rect 244 26 245 27 
<< m1 >>
rect 253 26 254 27 
<< m2 >>
rect 254 26 255 27 
<< m2 >>
rect 264 26 265 27 
<< m1 >>
rect 268 26 269 27 
<< m1 >>
rect 442 26 443 27 
<< m1 >>
rect 64 27 65 28 
<< m1 >>
rect 91 27 92 28 
<< m1 >>
rect 163 27 164 28 
<< m1 >>
rect 244 27 245 28 
<< m1 >>
rect 253 27 254 28 
<< m2 >>
rect 254 27 255 28 
<< m1 >>
rect 258 27 259 28 
<< m1 >>
rect 259 27 260 28 
<< m1 >>
rect 260 27 261 28 
<< m1 >>
rect 261 27 262 28 
<< m1 >>
rect 262 27 263 28 
<< m1 >>
rect 263 27 264 28 
<< m1 >>
rect 264 27 265 28 
<< m2 >>
rect 264 27 265 28 
<< m2c >>
rect 264 27 265 28 
<< m1 >>
rect 264 27 265 28 
<< m2 >>
rect 264 27 265 28 
<< m1 >>
rect 268 27 269 28 
<< m1 >>
rect 442 27 443 28 
<< m1 >>
rect 64 28 65 29 
<< m1 >>
rect 91 28 92 29 
<< m1 >>
rect 100 28 101 29 
<< m1 >>
rect 101 28 102 29 
<< m1 >>
rect 102 28 103 29 
<< m1 >>
rect 103 28 104 29 
<< m1 >>
rect 163 28 164 29 
<< m1 >>
rect 244 28 245 29 
<< m1 >>
rect 253 28 254 29 
<< m2 >>
rect 254 28 255 29 
<< m1 >>
rect 258 28 259 29 
<< m1 >>
rect 268 28 269 29 
<< m1 >>
rect 442 28 443 29 
<< m1 >>
rect 64 29 65 30 
<< m1 >>
rect 91 29 92 30 
<< m1 >>
rect 100 29 101 30 
<< m1 >>
rect 103 29 104 30 
<< m1 >>
rect 163 29 164 30 
<< m1 >>
rect 244 29 245 30 
<< m1 >>
rect 253 29 254 30 
<< m2 >>
rect 254 29 255 30 
<< m1 >>
rect 258 29 259 30 
<< m1 >>
rect 268 29 269 30 
<< m1 >>
rect 442 29 443 30 
<< pdiffusion >>
rect 12 30 13 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< pdiffusion >>
rect 15 30 16 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< pdiffusion >>
rect 30 30 31 31 
<< pdiffusion >>
rect 31 30 32 31 
<< pdiffusion >>
rect 32 30 33 31 
<< pdiffusion >>
rect 33 30 34 31 
<< pdiffusion >>
rect 34 30 35 31 
<< pdiffusion >>
rect 35 30 36 31 
<< pdiffusion >>
rect 48 30 49 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 64 30 65 31 
<< pdiffusion >>
rect 66 30 67 31 
<< pdiffusion >>
rect 67 30 68 31 
<< pdiffusion >>
rect 68 30 69 31 
<< pdiffusion >>
rect 69 30 70 31 
<< pdiffusion >>
rect 70 30 71 31 
<< pdiffusion >>
rect 71 30 72 31 
<< pdiffusion >>
rect 84 30 85 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< m1 >>
rect 91 30 92 31 
<< m1 >>
rect 100 30 101 31 
<< pdiffusion >>
rect 102 30 103 31 
<< m1 >>
rect 103 30 104 31 
<< pdiffusion >>
rect 103 30 104 31 
<< pdiffusion >>
rect 104 30 105 31 
<< pdiffusion >>
rect 105 30 106 31 
<< pdiffusion >>
rect 106 30 107 31 
<< pdiffusion >>
rect 107 30 108 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< pdiffusion >>
rect 156 30 157 31 
<< pdiffusion >>
rect 157 30 158 31 
<< pdiffusion >>
rect 158 30 159 31 
<< pdiffusion >>
rect 159 30 160 31 
<< pdiffusion >>
rect 160 30 161 31 
<< pdiffusion >>
rect 161 30 162 31 
<< m1 >>
rect 163 30 164 31 
<< pdiffusion >>
rect 174 30 175 31 
<< pdiffusion >>
rect 175 30 176 31 
<< pdiffusion >>
rect 176 30 177 31 
<< pdiffusion >>
rect 177 30 178 31 
<< pdiffusion >>
rect 178 30 179 31 
<< pdiffusion >>
rect 179 30 180 31 
<< pdiffusion >>
rect 192 30 193 31 
<< pdiffusion >>
rect 193 30 194 31 
<< pdiffusion >>
rect 194 30 195 31 
<< pdiffusion >>
rect 195 30 196 31 
<< pdiffusion >>
rect 196 30 197 31 
<< pdiffusion >>
rect 197 30 198 31 
<< pdiffusion >>
rect 210 30 211 31 
<< pdiffusion >>
rect 211 30 212 31 
<< pdiffusion >>
rect 212 30 213 31 
<< pdiffusion >>
rect 213 30 214 31 
<< pdiffusion >>
rect 214 30 215 31 
<< pdiffusion >>
rect 215 30 216 31 
<< pdiffusion >>
rect 228 30 229 31 
<< pdiffusion >>
rect 229 30 230 31 
<< pdiffusion >>
rect 230 30 231 31 
<< pdiffusion >>
rect 231 30 232 31 
<< pdiffusion >>
rect 232 30 233 31 
<< pdiffusion >>
rect 233 30 234 31 
<< m1 >>
rect 244 30 245 31 
<< pdiffusion >>
rect 246 30 247 31 
<< pdiffusion >>
rect 247 30 248 31 
<< pdiffusion >>
rect 248 30 249 31 
<< pdiffusion >>
rect 249 30 250 31 
<< pdiffusion >>
rect 250 30 251 31 
<< pdiffusion >>
rect 251 30 252 31 
<< m1 >>
rect 253 30 254 31 
<< m2 >>
rect 254 30 255 31 
<< m1 >>
rect 258 30 259 31 
<< pdiffusion >>
rect 264 30 265 31 
<< pdiffusion >>
rect 265 30 266 31 
<< pdiffusion >>
rect 266 30 267 31 
<< pdiffusion >>
rect 267 30 268 31 
<< m1 >>
rect 268 30 269 31 
<< pdiffusion >>
rect 268 30 269 31 
<< pdiffusion >>
rect 269 30 270 31 
<< pdiffusion >>
rect 282 30 283 31 
<< pdiffusion >>
rect 283 30 284 31 
<< pdiffusion >>
rect 284 30 285 31 
<< pdiffusion >>
rect 285 30 286 31 
<< pdiffusion >>
rect 286 30 287 31 
<< pdiffusion >>
rect 287 30 288 31 
<< pdiffusion >>
rect 300 30 301 31 
<< pdiffusion >>
rect 301 30 302 31 
<< pdiffusion >>
rect 302 30 303 31 
<< pdiffusion >>
rect 303 30 304 31 
<< pdiffusion >>
rect 304 30 305 31 
<< pdiffusion >>
rect 305 30 306 31 
<< pdiffusion >>
rect 318 30 319 31 
<< pdiffusion >>
rect 319 30 320 31 
<< pdiffusion >>
rect 320 30 321 31 
<< pdiffusion >>
rect 321 30 322 31 
<< pdiffusion >>
rect 322 30 323 31 
<< pdiffusion >>
rect 323 30 324 31 
<< pdiffusion >>
rect 336 30 337 31 
<< pdiffusion >>
rect 337 30 338 31 
<< pdiffusion >>
rect 338 30 339 31 
<< pdiffusion >>
rect 339 30 340 31 
<< pdiffusion >>
rect 340 30 341 31 
<< pdiffusion >>
rect 341 30 342 31 
<< pdiffusion >>
rect 354 30 355 31 
<< pdiffusion >>
rect 355 30 356 31 
<< pdiffusion >>
rect 356 30 357 31 
<< pdiffusion >>
rect 357 30 358 31 
<< pdiffusion >>
rect 358 30 359 31 
<< pdiffusion >>
rect 359 30 360 31 
<< pdiffusion >>
rect 372 30 373 31 
<< pdiffusion >>
rect 373 30 374 31 
<< pdiffusion >>
rect 374 30 375 31 
<< pdiffusion >>
rect 375 30 376 31 
<< pdiffusion >>
rect 376 30 377 31 
<< pdiffusion >>
rect 377 30 378 31 
<< pdiffusion >>
rect 390 30 391 31 
<< pdiffusion >>
rect 391 30 392 31 
<< pdiffusion >>
rect 392 30 393 31 
<< pdiffusion >>
rect 393 30 394 31 
<< pdiffusion >>
rect 394 30 395 31 
<< pdiffusion >>
rect 395 30 396 31 
<< pdiffusion >>
rect 408 30 409 31 
<< pdiffusion >>
rect 409 30 410 31 
<< pdiffusion >>
rect 410 30 411 31 
<< pdiffusion >>
rect 411 30 412 31 
<< pdiffusion >>
rect 412 30 413 31 
<< pdiffusion >>
rect 413 30 414 31 
<< pdiffusion >>
rect 426 30 427 31 
<< pdiffusion >>
rect 427 30 428 31 
<< pdiffusion >>
rect 428 30 429 31 
<< pdiffusion >>
rect 429 30 430 31 
<< pdiffusion >>
rect 430 30 431 31 
<< pdiffusion >>
rect 431 30 432 31 
<< m1 >>
rect 442 30 443 31 
<< pdiffusion >>
rect 444 30 445 31 
<< pdiffusion >>
rect 445 30 446 31 
<< pdiffusion >>
rect 446 30 447 31 
<< pdiffusion >>
rect 447 30 448 31 
<< pdiffusion >>
rect 448 30 449 31 
<< pdiffusion >>
rect 449 30 450 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< pdiffusion >>
rect 30 31 31 32 
<< pdiffusion >>
rect 31 31 32 32 
<< pdiffusion >>
rect 32 31 33 32 
<< pdiffusion >>
rect 33 31 34 32 
<< pdiffusion >>
rect 34 31 35 32 
<< pdiffusion >>
rect 35 31 36 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 64 31 65 32 
<< pdiffusion >>
rect 66 31 67 32 
<< pdiffusion >>
rect 67 31 68 32 
<< pdiffusion >>
rect 68 31 69 32 
<< pdiffusion >>
rect 69 31 70 32 
<< pdiffusion >>
rect 70 31 71 32 
<< pdiffusion >>
rect 71 31 72 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< m1 >>
rect 91 31 92 32 
<< m1 >>
rect 100 31 101 32 
<< pdiffusion >>
rect 102 31 103 32 
<< pdiffusion >>
rect 103 31 104 32 
<< pdiffusion >>
rect 104 31 105 32 
<< pdiffusion >>
rect 105 31 106 32 
<< pdiffusion >>
rect 106 31 107 32 
<< pdiffusion >>
rect 107 31 108 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< pdiffusion >>
rect 156 31 157 32 
<< pdiffusion >>
rect 157 31 158 32 
<< pdiffusion >>
rect 158 31 159 32 
<< pdiffusion >>
rect 159 31 160 32 
<< pdiffusion >>
rect 160 31 161 32 
<< pdiffusion >>
rect 161 31 162 32 
<< m1 >>
rect 163 31 164 32 
<< pdiffusion >>
rect 174 31 175 32 
<< pdiffusion >>
rect 175 31 176 32 
<< pdiffusion >>
rect 176 31 177 32 
<< pdiffusion >>
rect 177 31 178 32 
<< pdiffusion >>
rect 178 31 179 32 
<< pdiffusion >>
rect 179 31 180 32 
<< pdiffusion >>
rect 192 31 193 32 
<< pdiffusion >>
rect 193 31 194 32 
<< pdiffusion >>
rect 194 31 195 32 
<< pdiffusion >>
rect 195 31 196 32 
<< pdiffusion >>
rect 196 31 197 32 
<< pdiffusion >>
rect 197 31 198 32 
<< pdiffusion >>
rect 210 31 211 32 
<< pdiffusion >>
rect 211 31 212 32 
<< pdiffusion >>
rect 212 31 213 32 
<< pdiffusion >>
rect 213 31 214 32 
<< pdiffusion >>
rect 214 31 215 32 
<< pdiffusion >>
rect 215 31 216 32 
<< pdiffusion >>
rect 228 31 229 32 
<< pdiffusion >>
rect 229 31 230 32 
<< pdiffusion >>
rect 230 31 231 32 
<< pdiffusion >>
rect 231 31 232 32 
<< pdiffusion >>
rect 232 31 233 32 
<< pdiffusion >>
rect 233 31 234 32 
<< m1 >>
rect 244 31 245 32 
<< pdiffusion >>
rect 246 31 247 32 
<< pdiffusion >>
rect 247 31 248 32 
<< pdiffusion >>
rect 248 31 249 32 
<< pdiffusion >>
rect 249 31 250 32 
<< pdiffusion >>
rect 250 31 251 32 
<< pdiffusion >>
rect 251 31 252 32 
<< m1 >>
rect 253 31 254 32 
<< m2 >>
rect 254 31 255 32 
<< m1 >>
rect 258 31 259 32 
<< pdiffusion >>
rect 264 31 265 32 
<< pdiffusion >>
rect 265 31 266 32 
<< pdiffusion >>
rect 266 31 267 32 
<< pdiffusion >>
rect 267 31 268 32 
<< pdiffusion >>
rect 268 31 269 32 
<< pdiffusion >>
rect 269 31 270 32 
<< pdiffusion >>
rect 282 31 283 32 
<< pdiffusion >>
rect 283 31 284 32 
<< pdiffusion >>
rect 284 31 285 32 
<< pdiffusion >>
rect 285 31 286 32 
<< pdiffusion >>
rect 286 31 287 32 
<< pdiffusion >>
rect 287 31 288 32 
<< pdiffusion >>
rect 300 31 301 32 
<< pdiffusion >>
rect 301 31 302 32 
<< pdiffusion >>
rect 302 31 303 32 
<< pdiffusion >>
rect 303 31 304 32 
<< pdiffusion >>
rect 304 31 305 32 
<< pdiffusion >>
rect 305 31 306 32 
<< pdiffusion >>
rect 318 31 319 32 
<< pdiffusion >>
rect 319 31 320 32 
<< pdiffusion >>
rect 320 31 321 32 
<< pdiffusion >>
rect 321 31 322 32 
<< pdiffusion >>
rect 322 31 323 32 
<< pdiffusion >>
rect 323 31 324 32 
<< pdiffusion >>
rect 336 31 337 32 
<< pdiffusion >>
rect 337 31 338 32 
<< pdiffusion >>
rect 338 31 339 32 
<< pdiffusion >>
rect 339 31 340 32 
<< pdiffusion >>
rect 340 31 341 32 
<< pdiffusion >>
rect 341 31 342 32 
<< pdiffusion >>
rect 354 31 355 32 
<< pdiffusion >>
rect 355 31 356 32 
<< pdiffusion >>
rect 356 31 357 32 
<< pdiffusion >>
rect 357 31 358 32 
<< pdiffusion >>
rect 358 31 359 32 
<< pdiffusion >>
rect 359 31 360 32 
<< pdiffusion >>
rect 372 31 373 32 
<< pdiffusion >>
rect 373 31 374 32 
<< pdiffusion >>
rect 374 31 375 32 
<< pdiffusion >>
rect 375 31 376 32 
<< pdiffusion >>
rect 376 31 377 32 
<< pdiffusion >>
rect 377 31 378 32 
<< pdiffusion >>
rect 390 31 391 32 
<< pdiffusion >>
rect 391 31 392 32 
<< pdiffusion >>
rect 392 31 393 32 
<< pdiffusion >>
rect 393 31 394 32 
<< pdiffusion >>
rect 394 31 395 32 
<< pdiffusion >>
rect 395 31 396 32 
<< pdiffusion >>
rect 408 31 409 32 
<< pdiffusion >>
rect 409 31 410 32 
<< pdiffusion >>
rect 410 31 411 32 
<< pdiffusion >>
rect 411 31 412 32 
<< pdiffusion >>
rect 412 31 413 32 
<< pdiffusion >>
rect 413 31 414 32 
<< pdiffusion >>
rect 426 31 427 32 
<< pdiffusion >>
rect 427 31 428 32 
<< pdiffusion >>
rect 428 31 429 32 
<< pdiffusion >>
rect 429 31 430 32 
<< pdiffusion >>
rect 430 31 431 32 
<< pdiffusion >>
rect 431 31 432 32 
<< m1 >>
rect 442 31 443 32 
<< pdiffusion >>
rect 444 31 445 32 
<< pdiffusion >>
rect 445 31 446 32 
<< pdiffusion >>
rect 446 31 447 32 
<< pdiffusion >>
rect 447 31 448 32 
<< pdiffusion >>
rect 448 31 449 32 
<< pdiffusion >>
rect 449 31 450 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< pdiffusion >>
rect 30 32 31 33 
<< pdiffusion >>
rect 31 32 32 33 
<< pdiffusion >>
rect 32 32 33 33 
<< pdiffusion >>
rect 33 32 34 33 
<< pdiffusion >>
rect 34 32 35 33 
<< pdiffusion >>
rect 35 32 36 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 64 32 65 33 
<< pdiffusion >>
rect 66 32 67 33 
<< pdiffusion >>
rect 67 32 68 33 
<< pdiffusion >>
rect 68 32 69 33 
<< pdiffusion >>
rect 69 32 70 33 
<< pdiffusion >>
rect 70 32 71 33 
<< pdiffusion >>
rect 71 32 72 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< m1 >>
rect 91 32 92 33 
<< m1 >>
rect 100 32 101 33 
<< pdiffusion >>
rect 102 32 103 33 
<< pdiffusion >>
rect 103 32 104 33 
<< pdiffusion >>
rect 104 32 105 33 
<< pdiffusion >>
rect 105 32 106 33 
<< pdiffusion >>
rect 106 32 107 33 
<< pdiffusion >>
rect 107 32 108 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< pdiffusion >>
rect 156 32 157 33 
<< pdiffusion >>
rect 157 32 158 33 
<< pdiffusion >>
rect 158 32 159 33 
<< pdiffusion >>
rect 159 32 160 33 
<< pdiffusion >>
rect 160 32 161 33 
<< pdiffusion >>
rect 161 32 162 33 
<< m1 >>
rect 163 32 164 33 
<< pdiffusion >>
rect 174 32 175 33 
<< pdiffusion >>
rect 175 32 176 33 
<< pdiffusion >>
rect 176 32 177 33 
<< pdiffusion >>
rect 177 32 178 33 
<< pdiffusion >>
rect 178 32 179 33 
<< pdiffusion >>
rect 179 32 180 33 
<< pdiffusion >>
rect 192 32 193 33 
<< pdiffusion >>
rect 193 32 194 33 
<< pdiffusion >>
rect 194 32 195 33 
<< pdiffusion >>
rect 195 32 196 33 
<< pdiffusion >>
rect 196 32 197 33 
<< pdiffusion >>
rect 197 32 198 33 
<< pdiffusion >>
rect 210 32 211 33 
<< pdiffusion >>
rect 211 32 212 33 
<< pdiffusion >>
rect 212 32 213 33 
<< pdiffusion >>
rect 213 32 214 33 
<< pdiffusion >>
rect 214 32 215 33 
<< pdiffusion >>
rect 215 32 216 33 
<< pdiffusion >>
rect 228 32 229 33 
<< pdiffusion >>
rect 229 32 230 33 
<< pdiffusion >>
rect 230 32 231 33 
<< pdiffusion >>
rect 231 32 232 33 
<< pdiffusion >>
rect 232 32 233 33 
<< pdiffusion >>
rect 233 32 234 33 
<< m1 >>
rect 244 32 245 33 
<< pdiffusion >>
rect 246 32 247 33 
<< pdiffusion >>
rect 247 32 248 33 
<< pdiffusion >>
rect 248 32 249 33 
<< pdiffusion >>
rect 249 32 250 33 
<< pdiffusion >>
rect 250 32 251 33 
<< pdiffusion >>
rect 251 32 252 33 
<< m1 >>
rect 253 32 254 33 
<< m2 >>
rect 254 32 255 33 
<< m1 >>
rect 258 32 259 33 
<< pdiffusion >>
rect 264 32 265 33 
<< pdiffusion >>
rect 265 32 266 33 
<< pdiffusion >>
rect 266 32 267 33 
<< pdiffusion >>
rect 267 32 268 33 
<< pdiffusion >>
rect 268 32 269 33 
<< pdiffusion >>
rect 269 32 270 33 
<< pdiffusion >>
rect 282 32 283 33 
<< pdiffusion >>
rect 283 32 284 33 
<< pdiffusion >>
rect 284 32 285 33 
<< pdiffusion >>
rect 285 32 286 33 
<< pdiffusion >>
rect 286 32 287 33 
<< pdiffusion >>
rect 287 32 288 33 
<< pdiffusion >>
rect 300 32 301 33 
<< pdiffusion >>
rect 301 32 302 33 
<< pdiffusion >>
rect 302 32 303 33 
<< pdiffusion >>
rect 303 32 304 33 
<< pdiffusion >>
rect 304 32 305 33 
<< pdiffusion >>
rect 305 32 306 33 
<< pdiffusion >>
rect 318 32 319 33 
<< pdiffusion >>
rect 319 32 320 33 
<< pdiffusion >>
rect 320 32 321 33 
<< pdiffusion >>
rect 321 32 322 33 
<< pdiffusion >>
rect 322 32 323 33 
<< pdiffusion >>
rect 323 32 324 33 
<< pdiffusion >>
rect 336 32 337 33 
<< pdiffusion >>
rect 337 32 338 33 
<< pdiffusion >>
rect 338 32 339 33 
<< pdiffusion >>
rect 339 32 340 33 
<< pdiffusion >>
rect 340 32 341 33 
<< pdiffusion >>
rect 341 32 342 33 
<< pdiffusion >>
rect 354 32 355 33 
<< pdiffusion >>
rect 355 32 356 33 
<< pdiffusion >>
rect 356 32 357 33 
<< pdiffusion >>
rect 357 32 358 33 
<< pdiffusion >>
rect 358 32 359 33 
<< pdiffusion >>
rect 359 32 360 33 
<< pdiffusion >>
rect 372 32 373 33 
<< pdiffusion >>
rect 373 32 374 33 
<< pdiffusion >>
rect 374 32 375 33 
<< pdiffusion >>
rect 375 32 376 33 
<< pdiffusion >>
rect 376 32 377 33 
<< pdiffusion >>
rect 377 32 378 33 
<< pdiffusion >>
rect 390 32 391 33 
<< pdiffusion >>
rect 391 32 392 33 
<< pdiffusion >>
rect 392 32 393 33 
<< pdiffusion >>
rect 393 32 394 33 
<< pdiffusion >>
rect 394 32 395 33 
<< pdiffusion >>
rect 395 32 396 33 
<< pdiffusion >>
rect 408 32 409 33 
<< pdiffusion >>
rect 409 32 410 33 
<< pdiffusion >>
rect 410 32 411 33 
<< pdiffusion >>
rect 411 32 412 33 
<< pdiffusion >>
rect 412 32 413 33 
<< pdiffusion >>
rect 413 32 414 33 
<< pdiffusion >>
rect 426 32 427 33 
<< pdiffusion >>
rect 427 32 428 33 
<< pdiffusion >>
rect 428 32 429 33 
<< pdiffusion >>
rect 429 32 430 33 
<< pdiffusion >>
rect 430 32 431 33 
<< pdiffusion >>
rect 431 32 432 33 
<< m1 >>
rect 442 32 443 33 
<< pdiffusion >>
rect 444 32 445 33 
<< pdiffusion >>
rect 445 32 446 33 
<< pdiffusion >>
rect 446 32 447 33 
<< pdiffusion >>
rect 447 32 448 33 
<< pdiffusion >>
rect 448 32 449 33 
<< pdiffusion >>
rect 449 32 450 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< pdiffusion >>
rect 30 33 31 34 
<< pdiffusion >>
rect 31 33 32 34 
<< pdiffusion >>
rect 32 33 33 34 
<< pdiffusion >>
rect 33 33 34 34 
<< pdiffusion >>
rect 34 33 35 34 
<< pdiffusion >>
rect 35 33 36 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 64 33 65 34 
<< pdiffusion >>
rect 66 33 67 34 
<< pdiffusion >>
rect 67 33 68 34 
<< pdiffusion >>
rect 68 33 69 34 
<< pdiffusion >>
rect 69 33 70 34 
<< pdiffusion >>
rect 70 33 71 34 
<< pdiffusion >>
rect 71 33 72 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< m1 >>
rect 91 33 92 34 
<< m1 >>
rect 100 33 101 34 
<< pdiffusion >>
rect 102 33 103 34 
<< pdiffusion >>
rect 103 33 104 34 
<< pdiffusion >>
rect 104 33 105 34 
<< pdiffusion >>
rect 105 33 106 34 
<< pdiffusion >>
rect 106 33 107 34 
<< pdiffusion >>
rect 107 33 108 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< pdiffusion >>
rect 156 33 157 34 
<< pdiffusion >>
rect 157 33 158 34 
<< pdiffusion >>
rect 158 33 159 34 
<< pdiffusion >>
rect 159 33 160 34 
<< pdiffusion >>
rect 160 33 161 34 
<< pdiffusion >>
rect 161 33 162 34 
<< m1 >>
rect 163 33 164 34 
<< pdiffusion >>
rect 174 33 175 34 
<< pdiffusion >>
rect 175 33 176 34 
<< pdiffusion >>
rect 176 33 177 34 
<< pdiffusion >>
rect 177 33 178 34 
<< pdiffusion >>
rect 178 33 179 34 
<< pdiffusion >>
rect 179 33 180 34 
<< pdiffusion >>
rect 192 33 193 34 
<< pdiffusion >>
rect 193 33 194 34 
<< pdiffusion >>
rect 194 33 195 34 
<< pdiffusion >>
rect 195 33 196 34 
<< pdiffusion >>
rect 196 33 197 34 
<< pdiffusion >>
rect 197 33 198 34 
<< pdiffusion >>
rect 210 33 211 34 
<< pdiffusion >>
rect 211 33 212 34 
<< pdiffusion >>
rect 212 33 213 34 
<< pdiffusion >>
rect 213 33 214 34 
<< pdiffusion >>
rect 214 33 215 34 
<< pdiffusion >>
rect 215 33 216 34 
<< pdiffusion >>
rect 228 33 229 34 
<< pdiffusion >>
rect 229 33 230 34 
<< pdiffusion >>
rect 230 33 231 34 
<< pdiffusion >>
rect 231 33 232 34 
<< pdiffusion >>
rect 232 33 233 34 
<< pdiffusion >>
rect 233 33 234 34 
<< m1 >>
rect 244 33 245 34 
<< pdiffusion >>
rect 246 33 247 34 
<< pdiffusion >>
rect 247 33 248 34 
<< pdiffusion >>
rect 248 33 249 34 
<< pdiffusion >>
rect 249 33 250 34 
<< pdiffusion >>
rect 250 33 251 34 
<< pdiffusion >>
rect 251 33 252 34 
<< m1 >>
rect 253 33 254 34 
<< m2 >>
rect 254 33 255 34 
<< m1 >>
rect 258 33 259 34 
<< pdiffusion >>
rect 264 33 265 34 
<< pdiffusion >>
rect 265 33 266 34 
<< pdiffusion >>
rect 266 33 267 34 
<< pdiffusion >>
rect 267 33 268 34 
<< pdiffusion >>
rect 268 33 269 34 
<< pdiffusion >>
rect 269 33 270 34 
<< pdiffusion >>
rect 282 33 283 34 
<< pdiffusion >>
rect 283 33 284 34 
<< pdiffusion >>
rect 284 33 285 34 
<< pdiffusion >>
rect 285 33 286 34 
<< pdiffusion >>
rect 286 33 287 34 
<< pdiffusion >>
rect 287 33 288 34 
<< pdiffusion >>
rect 300 33 301 34 
<< pdiffusion >>
rect 301 33 302 34 
<< pdiffusion >>
rect 302 33 303 34 
<< pdiffusion >>
rect 303 33 304 34 
<< pdiffusion >>
rect 304 33 305 34 
<< pdiffusion >>
rect 305 33 306 34 
<< pdiffusion >>
rect 318 33 319 34 
<< pdiffusion >>
rect 319 33 320 34 
<< pdiffusion >>
rect 320 33 321 34 
<< pdiffusion >>
rect 321 33 322 34 
<< pdiffusion >>
rect 322 33 323 34 
<< pdiffusion >>
rect 323 33 324 34 
<< pdiffusion >>
rect 336 33 337 34 
<< pdiffusion >>
rect 337 33 338 34 
<< pdiffusion >>
rect 338 33 339 34 
<< pdiffusion >>
rect 339 33 340 34 
<< pdiffusion >>
rect 340 33 341 34 
<< pdiffusion >>
rect 341 33 342 34 
<< pdiffusion >>
rect 354 33 355 34 
<< pdiffusion >>
rect 355 33 356 34 
<< pdiffusion >>
rect 356 33 357 34 
<< pdiffusion >>
rect 357 33 358 34 
<< pdiffusion >>
rect 358 33 359 34 
<< pdiffusion >>
rect 359 33 360 34 
<< pdiffusion >>
rect 372 33 373 34 
<< pdiffusion >>
rect 373 33 374 34 
<< pdiffusion >>
rect 374 33 375 34 
<< pdiffusion >>
rect 375 33 376 34 
<< pdiffusion >>
rect 376 33 377 34 
<< pdiffusion >>
rect 377 33 378 34 
<< pdiffusion >>
rect 390 33 391 34 
<< pdiffusion >>
rect 391 33 392 34 
<< pdiffusion >>
rect 392 33 393 34 
<< pdiffusion >>
rect 393 33 394 34 
<< pdiffusion >>
rect 394 33 395 34 
<< pdiffusion >>
rect 395 33 396 34 
<< pdiffusion >>
rect 408 33 409 34 
<< pdiffusion >>
rect 409 33 410 34 
<< pdiffusion >>
rect 410 33 411 34 
<< pdiffusion >>
rect 411 33 412 34 
<< pdiffusion >>
rect 412 33 413 34 
<< pdiffusion >>
rect 413 33 414 34 
<< pdiffusion >>
rect 426 33 427 34 
<< pdiffusion >>
rect 427 33 428 34 
<< pdiffusion >>
rect 428 33 429 34 
<< pdiffusion >>
rect 429 33 430 34 
<< pdiffusion >>
rect 430 33 431 34 
<< pdiffusion >>
rect 431 33 432 34 
<< m1 >>
rect 442 33 443 34 
<< pdiffusion >>
rect 444 33 445 34 
<< pdiffusion >>
rect 445 33 446 34 
<< pdiffusion >>
rect 446 33 447 34 
<< pdiffusion >>
rect 447 33 448 34 
<< pdiffusion >>
rect 448 33 449 34 
<< pdiffusion >>
rect 449 33 450 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< pdiffusion >>
rect 30 34 31 35 
<< pdiffusion >>
rect 31 34 32 35 
<< pdiffusion >>
rect 32 34 33 35 
<< pdiffusion >>
rect 33 34 34 35 
<< pdiffusion >>
rect 34 34 35 35 
<< pdiffusion >>
rect 35 34 36 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 64 34 65 35 
<< pdiffusion >>
rect 66 34 67 35 
<< pdiffusion >>
rect 67 34 68 35 
<< pdiffusion >>
rect 68 34 69 35 
<< pdiffusion >>
rect 69 34 70 35 
<< pdiffusion >>
rect 70 34 71 35 
<< pdiffusion >>
rect 71 34 72 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< m1 >>
rect 91 34 92 35 
<< m1 >>
rect 100 34 101 35 
<< pdiffusion >>
rect 102 34 103 35 
<< pdiffusion >>
rect 103 34 104 35 
<< pdiffusion >>
rect 104 34 105 35 
<< pdiffusion >>
rect 105 34 106 35 
<< pdiffusion >>
rect 106 34 107 35 
<< pdiffusion >>
rect 107 34 108 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< pdiffusion >>
rect 156 34 157 35 
<< pdiffusion >>
rect 157 34 158 35 
<< pdiffusion >>
rect 158 34 159 35 
<< pdiffusion >>
rect 159 34 160 35 
<< pdiffusion >>
rect 160 34 161 35 
<< pdiffusion >>
rect 161 34 162 35 
<< m1 >>
rect 163 34 164 35 
<< pdiffusion >>
rect 174 34 175 35 
<< pdiffusion >>
rect 175 34 176 35 
<< pdiffusion >>
rect 176 34 177 35 
<< pdiffusion >>
rect 177 34 178 35 
<< pdiffusion >>
rect 178 34 179 35 
<< pdiffusion >>
rect 179 34 180 35 
<< pdiffusion >>
rect 192 34 193 35 
<< pdiffusion >>
rect 193 34 194 35 
<< pdiffusion >>
rect 194 34 195 35 
<< pdiffusion >>
rect 195 34 196 35 
<< pdiffusion >>
rect 196 34 197 35 
<< pdiffusion >>
rect 197 34 198 35 
<< pdiffusion >>
rect 210 34 211 35 
<< pdiffusion >>
rect 211 34 212 35 
<< pdiffusion >>
rect 212 34 213 35 
<< pdiffusion >>
rect 213 34 214 35 
<< pdiffusion >>
rect 214 34 215 35 
<< pdiffusion >>
rect 215 34 216 35 
<< pdiffusion >>
rect 228 34 229 35 
<< pdiffusion >>
rect 229 34 230 35 
<< pdiffusion >>
rect 230 34 231 35 
<< pdiffusion >>
rect 231 34 232 35 
<< pdiffusion >>
rect 232 34 233 35 
<< pdiffusion >>
rect 233 34 234 35 
<< m1 >>
rect 244 34 245 35 
<< pdiffusion >>
rect 246 34 247 35 
<< pdiffusion >>
rect 247 34 248 35 
<< pdiffusion >>
rect 248 34 249 35 
<< pdiffusion >>
rect 249 34 250 35 
<< pdiffusion >>
rect 250 34 251 35 
<< pdiffusion >>
rect 251 34 252 35 
<< m1 >>
rect 253 34 254 35 
<< m2 >>
rect 254 34 255 35 
<< m1 >>
rect 258 34 259 35 
<< pdiffusion >>
rect 264 34 265 35 
<< pdiffusion >>
rect 265 34 266 35 
<< pdiffusion >>
rect 266 34 267 35 
<< pdiffusion >>
rect 267 34 268 35 
<< pdiffusion >>
rect 268 34 269 35 
<< pdiffusion >>
rect 269 34 270 35 
<< pdiffusion >>
rect 282 34 283 35 
<< pdiffusion >>
rect 283 34 284 35 
<< pdiffusion >>
rect 284 34 285 35 
<< pdiffusion >>
rect 285 34 286 35 
<< pdiffusion >>
rect 286 34 287 35 
<< pdiffusion >>
rect 287 34 288 35 
<< pdiffusion >>
rect 300 34 301 35 
<< pdiffusion >>
rect 301 34 302 35 
<< pdiffusion >>
rect 302 34 303 35 
<< pdiffusion >>
rect 303 34 304 35 
<< pdiffusion >>
rect 304 34 305 35 
<< pdiffusion >>
rect 305 34 306 35 
<< pdiffusion >>
rect 318 34 319 35 
<< pdiffusion >>
rect 319 34 320 35 
<< pdiffusion >>
rect 320 34 321 35 
<< pdiffusion >>
rect 321 34 322 35 
<< pdiffusion >>
rect 322 34 323 35 
<< pdiffusion >>
rect 323 34 324 35 
<< pdiffusion >>
rect 336 34 337 35 
<< pdiffusion >>
rect 337 34 338 35 
<< pdiffusion >>
rect 338 34 339 35 
<< pdiffusion >>
rect 339 34 340 35 
<< pdiffusion >>
rect 340 34 341 35 
<< pdiffusion >>
rect 341 34 342 35 
<< pdiffusion >>
rect 354 34 355 35 
<< pdiffusion >>
rect 355 34 356 35 
<< pdiffusion >>
rect 356 34 357 35 
<< pdiffusion >>
rect 357 34 358 35 
<< pdiffusion >>
rect 358 34 359 35 
<< pdiffusion >>
rect 359 34 360 35 
<< pdiffusion >>
rect 372 34 373 35 
<< pdiffusion >>
rect 373 34 374 35 
<< pdiffusion >>
rect 374 34 375 35 
<< pdiffusion >>
rect 375 34 376 35 
<< pdiffusion >>
rect 376 34 377 35 
<< pdiffusion >>
rect 377 34 378 35 
<< pdiffusion >>
rect 390 34 391 35 
<< pdiffusion >>
rect 391 34 392 35 
<< pdiffusion >>
rect 392 34 393 35 
<< pdiffusion >>
rect 393 34 394 35 
<< pdiffusion >>
rect 394 34 395 35 
<< pdiffusion >>
rect 395 34 396 35 
<< pdiffusion >>
rect 408 34 409 35 
<< pdiffusion >>
rect 409 34 410 35 
<< pdiffusion >>
rect 410 34 411 35 
<< pdiffusion >>
rect 411 34 412 35 
<< pdiffusion >>
rect 412 34 413 35 
<< pdiffusion >>
rect 413 34 414 35 
<< pdiffusion >>
rect 426 34 427 35 
<< pdiffusion >>
rect 427 34 428 35 
<< pdiffusion >>
rect 428 34 429 35 
<< pdiffusion >>
rect 429 34 430 35 
<< pdiffusion >>
rect 430 34 431 35 
<< pdiffusion >>
rect 431 34 432 35 
<< m1 >>
rect 442 34 443 35 
<< pdiffusion >>
rect 444 34 445 35 
<< pdiffusion >>
rect 445 34 446 35 
<< pdiffusion >>
rect 446 34 447 35 
<< pdiffusion >>
rect 447 34 448 35 
<< pdiffusion >>
rect 448 34 449 35 
<< pdiffusion >>
rect 449 34 450 35 
<< pdiffusion >>
rect 12 35 13 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< pdiffusion >>
rect 30 35 31 36 
<< pdiffusion >>
rect 31 35 32 36 
<< pdiffusion >>
rect 32 35 33 36 
<< pdiffusion >>
rect 33 35 34 36 
<< pdiffusion >>
rect 34 35 35 36 
<< pdiffusion >>
rect 35 35 36 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 64 35 65 36 
<< pdiffusion >>
rect 66 35 67 36 
<< pdiffusion >>
rect 67 35 68 36 
<< pdiffusion >>
rect 68 35 69 36 
<< pdiffusion >>
rect 69 35 70 36 
<< pdiffusion >>
rect 70 35 71 36 
<< pdiffusion >>
rect 71 35 72 36 
<< pdiffusion >>
rect 84 35 85 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< m1 >>
rect 91 35 92 36 
<< m1 >>
rect 100 35 101 36 
<< pdiffusion >>
rect 102 35 103 36 
<< pdiffusion >>
rect 103 35 104 36 
<< pdiffusion >>
rect 104 35 105 36 
<< pdiffusion >>
rect 105 35 106 36 
<< pdiffusion >>
rect 106 35 107 36 
<< pdiffusion >>
rect 107 35 108 36 
<< pdiffusion >>
rect 120 35 121 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< pdiffusion >>
rect 156 35 157 36 
<< pdiffusion >>
rect 157 35 158 36 
<< pdiffusion >>
rect 158 35 159 36 
<< pdiffusion >>
rect 159 35 160 36 
<< pdiffusion >>
rect 160 35 161 36 
<< pdiffusion >>
rect 161 35 162 36 
<< m1 >>
rect 163 35 164 36 
<< pdiffusion >>
rect 174 35 175 36 
<< pdiffusion >>
rect 175 35 176 36 
<< pdiffusion >>
rect 176 35 177 36 
<< pdiffusion >>
rect 177 35 178 36 
<< m1 >>
rect 178 35 179 36 
<< pdiffusion >>
rect 178 35 179 36 
<< pdiffusion >>
rect 179 35 180 36 
<< pdiffusion >>
rect 192 35 193 36 
<< pdiffusion >>
rect 193 35 194 36 
<< pdiffusion >>
rect 194 35 195 36 
<< pdiffusion >>
rect 195 35 196 36 
<< pdiffusion >>
rect 196 35 197 36 
<< pdiffusion >>
rect 197 35 198 36 
<< pdiffusion >>
rect 210 35 211 36 
<< pdiffusion >>
rect 211 35 212 36 
<< pdiffusion >>
rect 212 35 213 36 
<< pdiffusion >>
rect 213 35 214 36 
<< pdiffusion >>
rect 214 35 215 36 
<< pdiffusion >>
rect 215 35 216 36 
<< pdiffusion >>
rect 228 35 229 36 
<< m1 >>
rect 229 35 230 36 
<< pdiffusion >>
rect 229 35 230 36 
<< pdiffusion >>
rect 230 35 231 36 
<< pdiffusion >>
rect 231 35 232 36 
<< pdiffusion >>
rect 232 35 233 36 
<< pdiffusion >>
rect 233 35 234 36 
<< m1 >>
rect 244 35 245 36 
<< pdiffusion >>
rect 246 35 247 36 
<< m1 >>
rect 247 35 248 36 
<< pdiffusion >>
rect 247 35 248 36 
<< pdiffusion >>
rect 248 35 249 36 
<< pdiffusion >>
rect 249 35 250 36 
<< pdiffusion >>
rect 250 35 251 36 
<< pdiffusion >>
rect 251 35 252 36 
<< m1 >>
rect 253 35 254 36 
<< m2 >>
rect 254 35 255 36 
<< m1 >>
rect 258 35 259 36 
<< pdiffusion >>
rect 264 35 265 36 
<< pdiffusion >>
rect 265 35 266 36 
<< pdiffusion >>
rect 266 35 267 36 
<< pdiffusion >>
rect 267 35 268 36 
<< pdiffusion >>
rect 268 35 269 36 
<< pdiffusion >>
rect 269 35 270 36 
<< pdiffusion >>
rect 282 35 283 36 
<< m1 >>
rect 283 35 284 36 
<< pdiffusion >>
rect 283 35 284 36 
<< pdiffusion >>
rect 284 35 285 36 
<< pdiffusion >>
rect 285 35 286 36 
<< pdiffusion >>
rect 286 35 287 36 
<< pdiffusion >>
rect 287 35 288 36 
<< pdiffusion >>
rect 300 35 301 36 
<< pdiffusion >>
rect 301 35 302 36 
<< pdiffusion >>
rect 302 35 303 36 
<< pdiffusion >>
rect 303 35 304 36 
<< pdiffusion >>
rect 304 35 305 36 
<< pdiffusion >>
rect 305 35 306 36 
<< pdiffusion >>
rect 318 35 319 36 
<< pdiffusion >>
rect 319 35 320 36 
<< pdiffusion >>
rect 320 35 321 36 
<< pdiffusion >>
rect 321 35 322 36 
<< pdiffusion >>
rect 322 35 323 36 
<< pdiffusion >>
rect 323 35 324 36 
<< pdiffusion >>
rect 336 35 337 36 
<< m1 >>
rect 337 35 338 36 
<< pdiffusion >>
rect 337 35 338 36 
<< pdiffusion >>
rect 338 35 339 36 
<< pdiffusion >>
rect 339 35 340 36 
<< pdiffusion >>
rect 340 35 341 36 
<< pdiffusion >>
rect 341 35 342 36 
<< pdiffusion >>
rect 354 35 355 36 
<< pdiffusion >>
rect 355 35 356 36 
<< pdiffusion >>
rect 356 35 357 36 
<< pdiffusion >>
rect 357 35 358 36 
<< pdiffusion >>
rect 358 35 359 36 
<< pdiffusion >>
rect 359 35 360 36 
<< pdiffusion >>
rect 372 35 373 36 
<< pdiffusion >>
rect 373 35 374 36 
<< pdiffusion >>
rect 374 35 375 36 
<< pdiffusion >>
rect 375 35 376 36 
<< m1 >>
rect 376 35 377 36 
<< pdiffusion >>
rect 376 35 377 36 
<< pdiffusion >>
rect 377 35 378 36 
<< pdiffusion >>
rect 390 35 391 36 
<< pdiffusion >>
rect 391 35 392 36 
<< pdiffusion >>
rect 392 35 393 36 
<< pdiffusion >>
rect 393 35 394 36 
<< pdiffusion >>
rect 394 35 395 36 
<< pdiffusion >>
rect 395 35 396 36 
<< pdiffusion >>
rect 408 35 409 36 
<< pdiffusion >>
rect 409 35 410 36 
<< pdiffusion >>
rect 410 35 411 36 
<< pdiffusion >>
rect 411 35 412 36 
<< pdiffusion >>
rect 412 35 413 36 
<< pdiffusion >>
rect 413 35 414 36 
<< pdiffusion >>
rect 426 35 427 36 
<< pdiffusion >>
rect 427 35 428 36 
<< pdiffusion >>
rect 428 35 429 36 
<< pdiffusion >>
rect 429 35 430 36 
<< pdiffusion >>
rect 430 35 431 36 
<< pdiffusion >>
rect 431 35 432 36 
<< m1 >>
rect 442 35 443 36 
<< pdiffusion >>
rect 444 35 445 36 
<< m1 >>
rect 445 35 446 36 
<< pdiffusion >>
rect 445 35 446 36 
<< pdiffusion >>
rect 446 35 447 36 
<< pdiffusion >>
rect 447 35 448 36 
<< pdiffusion >>
rect 448 35 449 36 
<< pdiffusion >>
rect 449 35 450 36 
<< m1 >>
rect 64 36 65 37 
<< m1 >>
rect 91 36 92 37 
<< m1 >>
rect 100 36 101 37 
<< m1 >>
rect 163 36 164 37 
<< m1 >>
rect 178 36 179 37 
<< m1 >>
rect 229 36 230 37 
<< m1 >>
rect 244 36 245 37 
<< m1 >>
rect 247 36 248 37 
<< m1 >>
rect 253 36 254 37 
<< m2 >>
rect 254 36 255 37 
<< m1 >>
rect 258 36 259 37 
<< m1 >>
rect 283 36 284 37 
<< m1 >>
rect 337 36 338 37 
<< m1 >>
rect 376 36 377 37 
<< m1 >>
rect 442 36 443 37 
<< m1 >>
rect 445 36 446 37 
<< m1 >>
rect 64 37 65 38 
<< m1 >>
rect 91 37 92 38 
<< m1 >>
rect 100 37 101 38 
<< m1 >>
rect 163 37 164 38 
<< m1 >>
rect 178 37 179 38 
<< m1 >>
rect 229 37 230 38 
<< m1 >>
rect 244 37 245 38 
<< m1 >>
rect 247 37 248 38 
<< m1 >>
rect 251 37 252 38 
<< m2 >>
rect 251 37 252 38 
<< m2c >>
rect 251 37 252 38 
<< m1 >>
rect 251 37 252 38 
<< m2 >>
rect 251 37 252 38 
<< m2 >>
rect 252 37 253 38 
<< m1 >>
rect 253 37 254 38 
<< m2 >>
rect 253 37 254 38 
<< m2 >>
rect 254 37 255 38 
<< m1 >>
rect 258 37 259 38 
<< m1 >>
rect 283 37 284 38 
<< m1 >>
rect 337 37 338 38 
<< m1 >>
rect 376 37 377 38 
<< m1 >>
rect 442 37 443 38 
<< m1 >>
rect 443 37 444 38 
<< m1 >>
rect 444 37 445 38 
<< m1 >>
rect 445 37 446 38 
<< m1 >>
rect 64 38 65 39 
<< m1 >>
rect 91 38 92 39 
<< m1 >>
rect 100 38 101 39 
<< m1 >>
rect 163 38 164 39 
<< m1 >>
rect 178 38 179 39 
<< m1 >>
rect 229 38 230 39 
<< m1 >>
rect 230 38 231 39 
<< m1 >>
rect 231 38 232 39 
<< m1 >>
rect 232 38 233 39 
<< m1 >>
rect 233 38 234 39 
<< m1 >>
rect 234 38 235 39 
<< m1 >>
rect 235 38 236 39 
<< m1 >>
rect 236 38 237 39 
<< m1 >>
rect 237 38 238 39 
<< m1 >>
rect 238 38 239 39 
<< m1 >>
rect 239 38 240 39 
<< m1 >>
rect 240 38 241 39 
<< m1 >>
rect 241 38 242 39 
<< m1 >>
rect 242 38 243 39 
<< m1 >>
rect 243 38 244 39 
<< m1 >>
rect 244 38 245 39 
<< m1 >>
rect 247 38 248 39 
<< m1 >>
rect 248 38 249 39 
<< m1 >>
rect 249 38 250 39 
<< m2 >>
rect 249 38 250 39 
<< m2c >>
rect 249 38 250 39 
<< m1 >>
rect 249 38 250 39 
<< m2 >>
rect 249 38 250 39 
<< m1 >>
rect 251 38 252 39 
<< m1 >>
rect 253 38 254 39 
<< m1 >>
rect 258 38 259 39 
<< m1 >>
rect 283 38 284 39 
<< m1 >>
rect 337 38 338 39 
<< m1 >>
rect 376 38 377 39 
<< m1 >>
rect 64 39 65 40 
<< m1 >>
rect 91 39 92 40 
<< m1 >>
rect 100 39 101 40 
<< m1 >>
rect 163 39 164 40 
<< m1 >>
rect 178 39 179 40 
<< m2 >>
rect 249 39 250 40 
<< m2 >>
rect 250 39 251 40 
<< m1 >>
rect 251 39 252 40 
<< m2 >>
rect 251 39 252 40 
<< m2 >>
rect 252 39 253 40 
<< m1 >>
rect 253 39 254 40 
<< m2 >>
rect 253 39 254 40 
<< m2 >>
rect 254 39 255 40 
<< m1 >>
rect 255 39 256 40 
<< m2 >>
rect 255 39 256 40 
<< m2c >>
rect 255 39 256 40 
<< m1 >>
rect 255 39 256 40 
<< m2 >>
rect 255 39 256 40 
<< m1 >>
rect 256 39 257 40 
<< m1 >>
rect 257 39 258 40 
<< m1 >>
rect 258 39 259 40 
<< m1 >>
rect 283 39 284 40 
<< m1 >>
rect 337 39 338 40 
<< m1 >>
rect 376 39 377 40 
<< m1 >>
rect 64 40 65 41 
<< m1 >>
rect 91 40 92 41 
<< m1 >>
rect 100 40 101 41 
<< m1 >>
rect 101 40 102 41 
<< m1 >>
rect 102 40 103 41 
<< m1 >>
rect 103 40 104 41 
<< m1 >>
rect 163 40 164 41 
<< m1 >>
rect 164 40 165 41 
<< m1 >>
rect 165 40 166 41 
<< m1 >>
rect 166 40 167 41 
<< m1 >>
rect 167 40 168 41 
<< m1 >>
rect 168 40 169 41 
<< m1 >>
rect 169 40 170 41 
<< m1 >>
rect 170 40 171 41 
<< m1 >>
rect 171 40 172 41 
<< m1 >>
rect 172 40 173 41 
<< m1 >>
rect 173 40 174 41 
<< m1 >>
rect 174 40 175 41 
<< m1 >>
rect 175 40 176 41 
<< m1 >>
rect 176 40 177 41 
<< m1 >>
rect 177 40 178 41 
<< m1 >>
rect 178 40 179 41 
<< m1 >>
rect 228 40 229 41 
<< m1 >>
rect 229 40 230 41 
<< m1 >>
rect 230 40 231 41 
<< m1 >>
rect 231 40 232 41 
<< m1 >>
rect 232 40 233 41 
<< m1 >>
rect 233 40 234 41 
<< m1 >>
rect 234 40 235 41 
<< m1 >>
rect 235 40 236 41 
<< m1 >>
rect 236 40 237 41 
<< m1 >>
rect 237 40 238 41 
<< m1 >>
rect 238 40 239 41 
<< m1 >>
rect 239 40 240 41 
<< m1 >>
rect 240 40 241 41 
<< m1 >>
rect 241 40 242 41 
<< m1 >>
rect 242 40 243 41 
<< m1 >>
rect 243 40 244 41 
<< m1 >>
rect 244 40 245 41 
<< m1 >>
rect 245 40 246 41 
<< m1 >>
rect 246 40 247 41 
<< m1 >>
rect 247 40 248 41 
<< m1 >>
rect 248 40 249 41 
<< m1 >>
rect 249 40 250 41 
<< m1 >>
rect 250 40 251 41 
<< m1 >>
rect 251 40 252 41 
<< m1 >>
rect 253 40 254 41 
<< m1 >>
rect 260 40 261 41 
<< m1 >>
rect 261 40 262 41 
<< m1 >>
rect 262 40 263 41 
<< m1 >>
rect 263 40 264 41 
<< m1 >>
rect 264 40 265 41 
<< m1 >>
rect 265 40 266 41 
<< m1 >>
rect 266 40 267 41 
<< m1 >>
rect 267 40 268 41 
<< m1 >>
rect 268 40 269 41 
<< m1 >>
rect 269 40 270 41 
<< m1 >>
rect 270 40 271 41 
<< m1 >>
rect 271 40 272 41 
<< m1 >>
rect 272 40 273 41 
<< m1 >>
rect 273 40 274 41 
<< m1 >>
rect 274 40 275 41 
<< m1 >>
rect 275 40 276 41 
<< m1 >>
rect 276 40 277 41 
<< m1 >>
rect 277 40 278 41 
<< m1 >>
rect 278 40 279 41 
<< m1 >>
rect 279 40 280 41 
<< m1 >>
rect 280 40 281 41 
<< m1 >>
rect 281 40 282 41 
<< m1 >>
rect 282 40 283 41 
<< m1 >>
rect 283 40 284 41 
<< m1 >>
rect 337 40 338 41 
<< m1 >>
rect 338 40 339 41 
<< m1 >>
rect 339 40 340 41 
<< m1 >>
rect 340 40 341 41 
<< m1 >>
rect 341 40 342 41 
<< m1 >>
rect 342 40 343 41 
<< m1 >>
rect 343 40 344 41 
<< m1 >>
rect 344 40 345 41 
<< m1 >>
rect 345 40 346 41 
<< m1 >>
rect 346 40 347 41 
<< m1 >>
rect 347 40 348 41 
<< m1 >>
rect 348 40 349 41 
<< m1 >>
rect 349 40 350 41 
<< m1 >>
rect 350 40 351 41 
<< m1 >>
rect 351 40 352 41 
<< m1 >>
rect 352 40 353 41 
<< m1 >>
rect 353 40 354 41 
<< m1 >>
rect 354 40 355 41 
<< m1 >>
rect 355 40 356 41 
<< m1 >>
rect 356 40 357 41 
<< m1 >>
rect 357 40 358 41 
<< m1 >>
rect 358 40 359 41 
<< m1 >>
rect 359 40 360 41 
<< m1 >>
rect 360 40 361 41 
<< m1 >>
rect 361 40 362 41 
<< m1 >>
rect 362 40 363 41 
<< m1 >>
rect 363 40 364 41 
<< m1 >>
rect 364 40 365 41 
<< m1 >>
rect 365 40 366 41 
<< m1 >>
rect 366 40 367 41 
<< m1 >>
rect 367 40 368 41 
<< m1 >>
rect 368 40 369 41 
<< m1 >>
rect 369 40 370 41 
<< m1 >>
rect 370 40 371 41 
<< m1 >>
rect 371 40 372 41 
<< m1 >>
rect 372 40 373 41 
<< m1 >>
rect 373 40 374 41 
<< m1 >>
rect 374 40 375 41 
<< m1 >>
rect 375 40 376 41 
<< m1 >>
rect 376 40 377 41 
<< m1 >>
rect 64 41 65 42 
<< m1 >>
rect 91 41 92 42 
<< m1 >>
rect 103 41 104 42 
<< m1 >>
rect 228 41 229 42 
<< m1 >>
rect 253 41 254 42 
<< m1 >>
rect 260 41 261 42 
<< m1 >>
rect 64 42 65 43 
<< m1 >>
rect 91 42 92 43 
<< m1 >>
rect 103 42 104 43 
<< m1 >>
rect 228 42 229 43 
<< m1 >>
rect 253 42 254 43 
<< m1 >>
rect 260 42 261 43 
<< m1 >>
rect 64 43 65 44 
<< m1 >>
rect 91 43 92 44 
<< m1 >>
rect 103 43 104 44 
<< m1 >>
rect 172 43 173 44 
<< m1 >>
rect 173 43 174 44 
<< m1 >>
rect 174 43 175 44 
<< m1 >>
rect 175 43 176 44 
<< m1 >>
rect 176 43 177 44 
<< m1 >>
rect 177 43 178 44 
<< m1 >>
rect 178 43 179 44 
<< m1 >>
rect 179 43 180 44 
<< m1 >>
rect 180 43 181 44 
<< m1 >>
rect 181 43 182 44 
<< m1 >>
rect 182 43 183 44 
<< m1 >>
rect 183 43 184 44 
<< m1 >>
rect 184 43 185 44 
<< m1 >>
rect 185 43 186 44 
<< m1 >>
rect 186 43 187 44 
<< m1 >>
rect 187 43 188 44 
<< m1 >>
rect 188 43 189 44 
<< m1 >>
rect 189 43 190 44 
<< m1 >>
rect 190 43 191 44 
<< m1 >>
rect 191 43 192 44 
<< m1 >>
rect 192 43 193 44 
<< m1 >>
rect 193 43 194 44 
<< m1 >>
rect 194 43 195 44 
<< m1 >>
rect 195 43 196 44 
<< m1 >>
rect 196 43 197 44 
<< m1 >>
rect 228 43 229 44 
<< m1 >>
rect 253 43 254 44 
<< m1 >>
rect 260 43 261 44 
<< m1 >>
rect 64 44 65 45 
<< m1 >>
rect 91 44 92 45 
<< m1 >>
rect 103 44 104 45 
<< m1 >>
rect 172 44 173 45 
<< m1 >>
rect 196 44 197 45 
<< m1 >>
rect 228 44 229 45 
<< m2 >>
rect 228 44 229 45 
<< m2c >>
rect 228 44 229 45 
<< m1 >>
rect 228 44 229 45 
<< m2 >>
rect 228 44 229 45 
<< m1 >>
rect 253 44 254 45 
<< m1 >>
rect 260 44 261 45 
<< m1 >>
rect 64 45 65 46 
<< m1 >>
rect 91 45 92 46 
<< m1 >>
rect 103 45 104 46 
<< m1 >>
rect 172 45 173 46 
<< m1 >>
rect 196 45 197 46 
<< m2 >>
rect 218 45 219 46 
<< m2 >>
rect 219 45 220 46 
<< m2 >>
rect 220 45 221 46 
<< m2 >>
rect 221 45 222 46 
<< m2 >>
rect 222 45 223 46 
<< m2 >>
rect 223 45 224 46 
<< m2 >>
rect 224 45 225 46 
<< m2 >>
rect 225 45 226 46 
<< m2 >>
rect 226 45 227 46 
<< m2 >>
rect 227 45 228 46 
<< m2 >>
rect 228 45 229 46 
<< m1 >>
rect 253 45 254 46 
<< m1 >>
rect 260 45 261 46 
<< m1 >>
rect 64 46 65 47 
<< m1 >>
rect 91 46 92 47 
<< m1 >>
rect 103 46 104 47 
<< m1 >>
rect 145 46 146 47 
<< m1 >>
rect 146 46 147 47 
<< m1 >>
rect 147 46 148 47 
<< m1 >>
rect 148 46 149 47 
<< m1 >>
rect 149 46 150 47 
<< m1 >>
rect 150 46 151 47 
<< m1 >>
rect 151 46 152 47 
<< m1 >>
rect 152 46 153 47 
<< m1 >>
rect 153 46 154 47 
<< m1 >>
rect 154 46 155 47 
<< m1 >>
rect 155 46 156 47 
<< m1 >>
rect 156 46 157 47 
<< m1 >>
rect 157 46 158 47 
<< m1 >>
rect 172 46 173 47 
<< m1 >>
rect 196 46 197 47 
<< m1 >>
rect 217 46 218 47 
<< m1 >>
rect 218 46 219 47 
<< m2 >>
rect 218 46 219 47 
<< m1 >>
rect 219 46 220 47 
<< m1 >>
rect 220 46 221 47 
<< m1 >>
rect 221 46 222 47 
<< m1 >>
rect 222 46 223 47 
<< m1 >>
rect 223 46 224 47 
<< m1 >>
rect 224 46 225 47 
<< m1 >>
rect 225 46 226 47 
<< m1 >>
rect 226 46 227 47 
<< m1 >>
rect 227 46 228 47 
<< m1 >>
rect 228 46 229 47 
<< m1 >>
rect 229 46 230 47 
<< m1 >>
rect 253 46 254 47 
<< m1 >>
rect 260 46 261 47 
<< m1 >>
rect 64 47 65 48 
<< m1 >>
rect 91 47 92 48 
<< m1 >>
rect 103 47 104 48 
<< m1 >>
rect 145 47 146 48 
<< m1 >>
rect 157 47 158 48 
<< m1 >>
rect 172 47 173 48 
<< m1 >>
rect 196 47 197 48 
<< m1 >>
rect 217 47 218 48 
<< m2 >>
rect 218 47 219 48 
<< m1 >>
rect 229 47 230 48 
<< m1 >>
rect 253 47 254 48 
<< m1 >>
rect 260 47 261 48 
<< pdiffusion >>
rect 12 48 13 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< pdiffusion >>
rect 30 48 31 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< pdiffusion >>
rect 48 48 49 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 64 48 65 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< pdiffusion >>
rect 84 48 85 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< pdiffusion >>
rect 102 48 103 49 
<< m1 >>
rect 103 48 104 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< pdiffusion >>
rect 120 48 121 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< pdiffusion >>
rect 138 48 139 49 
<< pdiffusion >>
rect 139 48 140 49 
<< pdiffusion >>
rect 140 48 141 49 
<< pdiffusion >>
rect 141 48 142 49 
<< pdiffusion >>
rect 142 48 143 49 
<< pdiffusion >>
rect 143 48 144 49 
<< m1 >>
rect 145 48 146 49 
<< pdiffusion >>
rect 156 48 157 49 
<< m1 >>
rect 157 48 158 49 
<< pdiffusion >>
rect 157 48 158 49 
<< pdiffusion >>
rect 158 48 159 49 
<< pdiffusion >>
rect 159 48 160 49 
<< pdiffusion >>
rect 160 48 161 49 
<< pdiffusion >>
rect 161 48 162 49 
<< m1 >>
rect 172 48 173 49 
<< pdiffusion >>
rect 174 48 175 49 
<< pdiffusion >>
rect 175 48 176 49 
<< pdiffusion >>
rect 176 48 177 49 
<< pdiffusion >>
rect 177 48 178 49 
<< pdiffusion >>
rect 178 48 179 49 
<< pdiffusion >>
rect 179 48 180 49 
<< pdiffusion >>
rect 192 48 193 49 
<< pdiffusion >>
rect 193 48 194 49 
<< pdiffusion >>
rect 194 48 195 49 
<< pdiffusion >>
rect 195 48 196 49 
<< m1 >>
rect 196 48 197 49 
<< pdiffusion >>
rect 196 48 197 49 
<< pdiffusion >>
rect 197 48 198 49 
<< pdiffusion >>
rect 210 48 211 49 
<< pdiffusion >>
rect 211 48 212 49 
<< pdiffusion >>
rect 212 48 213 49 
<< pdiffusion >>
rect 213 48 214 49 
<< pdiffusion >>
rect 214 48 215 49 
<< pdiffusion >>
rect 215 48 216 49 
<< m1 >>
rect 217 48 218 49 
<< m2 >>
rect 218 48 219 49 
<< pdiffusion >>
rect 228 48 229 49 
<< m1 >>
rect 229 48 230 49 
<< pdiffusion >>
rect 229 48 230 49 
<< pdiffusion >>
rect 230 48 231 49 
<< pdiffusion >>
rect 231 48 232 49 
<< pdiffusion >>
rect 232 48 233 49 
<< pdiffusion >>
rect 233 48 234 49 
<< pdiffusion >>
rect 246 48 247 49 
<< pdiffusion >>
rect 247 48 248 49 
<< pdiffusion >>
rect 248 48 249 49 
<< pdiffusion >>
rect 249 48 250 49 
<< pdiffusion >>
rect 250 48 251 49 
<< pdiffusion >>
rect 251 48 252 49 
<< m1 >>
rect 253 48 254 49 
<< m1 >>
rect 260 48 261 49 
<< pdiffusion >>
rect 264 48 265 49 
<< pdiffusion >>
rect 265 48 266 49 
<< pdiffusion >>
rect 266 48 267 49 
<< pdiffusion >>
rect 267 48 268 49 
<< pdiffusion >>
rect 268 48 269 49 
<< pdiffusion >>
rect 269 48 270 49 
<< pdiffusion >>
rect 282 48 283 49 
<< pdiffusion >>
rect 283 48 284 49 
<< pdiffusion >>
rect 284 48 285 49 
<< pdiffusion >>
rect 285 48 286 49 
<< pdiffusion >>
rect 286 48 287 49 
<< pdiffusion >>
rect 287 48 288 49 
<< pdiffusion >>
rect 300 48 301 49 
<< pdiffusion >>
rect 301 48 302 49 
<< pdiffusion >>
rect 302 48 303 49 
<< pdiffusion >>
rect 303 48 304 49 
<< pdiffusion >>
rect 304 48 305 49 
<< pdiffusion >>
rect 305 48 306 49 
<< pdiffusion >>
rect 318 48 319 49 
<< pdiffusion >>
rect 319 48 320 49 
<< pdiffusion >>
rect 320 48 321 49 
<< pdiffusion >>
rect 321 48 322 49 
<< pdiffusion >>
rect 322 48 323 49 
<< pdiffusion >>
rect 323 48 324 49 
<< pdiffusion >>
rect 336 48 337 49 
<< pdiffusion >>
rect 337 48 338 49 
<< pdiffusion >>
rect 338 48 339 49 
<< pdiffusion >>
rect 339 48 340 49 
<< pdiffusion >>
rect 340 48 341 49 
<< pdiffusion >>
rect 341 48 342 49 
<< pdiffusion >>
rect 354 48 355 49 
<< pdiffusion >>
rect 355 48 356 49 
<< pdiffusion >>
rect 356 48 357 49 
<< pdiffusion >>
rect 357 48 358 49 
<< pdiffusion >>
rect 358 48 359 49 
<< pdiffusion >>
rect 359 48 360 49 
<< pdiffusion >>
rect 390 48 391 49 
<< pdiffusion >>
rect 391 48 392 49 
<< pdiffusion >>
rect 392 48 393 49 
<< pdiffusion >>
rect 393 48 394 49 
<< pdiffusion >>
rect 394 48 395 49 
<< pdiffusion >>
rect 395 48 396 49 
<< pdiffusion >>
rect 408 48 409 49 
<< pdiffusion >>
rect 409 48 410 49 
<< pdiffusion >>
rect 410 48 411 49 
<< pdiffusion >>
rect 411 48 412 49 
<< pdiffusion >>
rect 412 48 413 49 
<< pdiffusion >>
rect 413 48 414 49 
<< pdiffusion >>
rect 426 48 427 49 
<< pdiffusion >>
rect 427 48 428 49 
<< pdiffusion >>
rect 428 48 429 49 
<< pdiffusion >>
rect 429 48 430 49 
<< pdiffusion >>
rect 430 48 431 49 
<< pdiffusion >>
rect 431 48 432 49 
<< pdiffusion >>
rect 444 48 445 49 
<< pdiffusion >>
rect 445 48 446 49 
<< pdiffusion >>
rect 446 48 447 49 
<< pdiffusion >>
rect 447 48 448 49 
<< pdiffusion >>
rect 448 48 449 49 
<< pdiffusion >>
rect 449 48 450 49 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 64 49 65 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< pdiffusion >>
rect 138 49 139 50 
<< pdiffusion >>
rect 139 49 140 50 
<< pdiffusion >>
rect 140 49 141 50 
<< pdiffusion >>
rect 141 49 142 50 
<< pdiffusion >>
rect 142 49 143 50 
<< pdiffusion >>
rect 143 49 144 50 
<< m1 >>
rect 145 49 146 50 
<< pdiffusion >>
rect 156 49 157 50 
<< pdiffusion >>
rect 157 49 158 50 
<< pdiffusion >>
rect 158 49 159 50 
<< pdiffusion >>
rect 159 49 160 50 
<< pdiffusion >>
rect 160 49 161 50 
<< pdiffusion >>
rect 161 49 162 50 
<< m1 >>
rect 172 49 173 50 
<< pdiffusion >>
rect 174 49 175 50 
<< pdiffusion >>
rect 175 49 176 50 
<< pdiffusion >>
rect 176 49 177 50 
<< pdiffusion >>
rect 177 49 178 50 
<< pdiffusion >>
rect 178 49 179 50 
<< pdiffusion >>
rect 179 49 180 50 
<< pdiffusion >>
rect 192 49 193 50 
<< pdiffusion >>
rect 193 49 194 50 
<< pdiffusion >>
rect 194 49 195 50 
<< pdiffusion >>
rect 195 49 196 50 
<< pdiffusion >>
rect 196 49 197 50 
<< pdiffusion >>
rect 197 49 198 50 
<< pdiffusion >>
rect 210 49 211 50 
<< pdiffusion >>
rect 211 49 212 50 
<< pdiffusion >>
rect 212 49 213 50 
<< pdiffusion >>
rect 213 49 214 50 
<< pdiffusion >>
rect 214 49 215 50 
<< pdiffusion >>
rect 215 49 216 50 
<< m1 >>
rect 217 49 218 50 
<< m2 >>
rect 218 49 219 50 
<< pdiffusion >>
rect 228 49 229 50 
<< pdiffusion >>
rect 229 49 230 50 
<< pdiffusion >>
rect 230 49 231 50 
<< pdiffusion >>
rect 231 49 232 50 
<< pdiffusion >>
rect 232 49 233 50 
<< pdiffusion >>
rect 233 49 234 50 
<< pdiffusion >>
rect 246 49 247 50 
<< pdiffusion >>
rect 247 49 248 50 
<< pdiffusion >>
rect 248 49 249 50 
<< pdiffusion >>
rect 249 49 250 50 
<< pdiffusion >>
rect 250 49 251 50 
<< pdiffusion >>
rect 251 49 252 50 
<< m1 >>
rect 253 49 254 50 
<< m1 >>
rect 260 49 261 50 
<< pdiffusion >>
rect 264 49 265 50 
<< pdiffusion >>
rect 265 49 266 50 
<< pdiffusion >>
rect 266 49 267 50 
<< pdiffusion >>
rect 267 49 268 50 
<< pdiffusion >>
rect 268 49 269 50 
<< pdiffusion >>
rect 269 49 270 50 
<< pdiffusion >>
rect 282 49 283 50 
<< pdiffusion >>
rect 283 49 284 50 
<< pdiffusion >>
rect 284 49 285 50 
<< pdiffusion >>
rect 285 49 286 50 
<< pdiffusion >>
rect 286 49 287 50 
<< pdiffusion >>
rect 287 49 288 50 
<< pdiffusion >>
rect 300 49 301 50 
<< pdiffusion >>
rect 301 49 302 50 
<< pdiffusion >>
rect 302 49 303 50 
<< pdiffusion >>
rect 303 49 304 50 
<< pdiffusion >>
rect 304 49 305 50 
<< pdiffusion >>
rect 305 49 306 50 
<< pdiffusion >>
rect 318 49 319 50 
<< pdiffusion >>
rect 319 49 320 50 
<< pdiffusion >>
rect 320 49 321 50 
<< pdiffusion >>
rect 321 49 322 50 
<< pdiffusion >>
rect 322 49 323 50 
<< pdiffusion >>
rect 323 49 324 50 
<< pdiffusion >>
rect 336 49 337 50 
<< pdiffusion >>
rect 337 49 338 50 
<< pdiffusion >>
rect 338 49 339 50 
<< pdiffusion >>
rect 339 49 340 50 
<< pdiffusion >>
rect 340 49 341 50 
<< pdiffusion >>
rect 341 49 342 50 
<< pdiffusion >>
rect 354 49 355 50 
<< pdiffusion >>
rect 355 49 356 50 
<< pdiffusion >>
rect 356 49 357 50 
<< pdiffusion >>
rect 357 49 358 50 
<< pdiffusion >>
rect 358 49 359 50 
<< pdiffusion >>
rect 359 49 360 50 
<< pdiffusion >>
rect 390 49 391 50 
<< pdiffusion >>
rect 391 49 392 50 
<< pdiffusion >>
rect 392 49 393 50 
<< pdiffusion >>
rect 393 49 394 50 
<< pdiffusion >>
rect 394 49 395 50 
<< pdiffusion >>
rect 395 49 396 50 
<< pdiffusion >>
rect 408 49 409 50 
<< pdiffusion >>
rect 409 49 410 50 
<< pdiffusion >>
rect 410 49 411 50 
<< pdiffusion >>
rect 411 49 412 50 
<< pdiffusion >>
rect 412 49 413 50 
<< pdiffusion >>
rect 413 49 414 50 
<< pdiffusion >>
rect 426 49 427 50 
<< pdiffusion >>
rect 427 49 428 50 
<< pdiffusion >>
rect 428 49 429 50 
<< pdiffusion >>
rect 429 49 430 50 
<< pdiffusion >>
rect 430 49 431 50 
<< pdiffusion >>
rect 431 49 432 50 
<< pdiffusion >>
rect 444 49 445 50 
<< pdiffusion >>
rect 445 49 446 50 
<< pdiffusion >>
rect 446 49 447 50 
<< pdiffusion >>
rect 447 49 448 50 
<< pdiffusion >>
rect 448 49 449 50 
<< pdiffusion >>
rect 449 49 450 50 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 64 50 65 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< pdiffusion >>
rect 138 50 139 51 
<< pdiffusion >>
rect 139 50 140 51 
<< pdiffusion >>
rect 140 50 141 51 
<< pdiffusion >>
rect 141 50 142 51 
<< pdiffusion >>
rect 142 50 143 51 
<< pdiffusion >>
rect 143 50 144 51 
<< m1 >>
rect 145 50 146 51 
<< pdiffusion >>
rect 156 50 157 51 
<< pdiffusion >>
rect 157 50 158 51 
<< pdiffusion >>
rect 158 50 159 51 
<< pdiffusion >>
rect 159 50 160 51 
<< pdiffusion >>
rect 160 50 161 51 
<< pdiffusion >>
rect 161 50 162 51 
<< m1 >>
rect 172 50 173 51 
<< pdiffusion >>
rect 174 50 175 51 
<< pdiffusion >>
rect 175 50 176 51 
<< pdiffusion >>
rect 176 50 177 51 
<< pdiffusion >>
rect 177 50 178 51 
<< pdiffusion >>
rect 178 50 179 51 
<< pdiffusion >>
rect 179 50 180 51 
<< pdiffusion >>
rect 192 50 193 51 
<< pdiffusion >>
rect 193 50 194 51 
<< pdiffusion >>
rect 194 50 195 51 
<< pdiffusion >>
rect 195 50 196 51 
<< pdiffusion >>
rect 196 50 197 51 
<< pdiffusion >>
rect 197 50 198 51 
<< pdiffusion >>
rect 210 50 211 51 
<< pdiffusion >>
rect 211 50 212 51 
<< pdiffusion >>
rect 212 50 213 51 
<< pdiffusion >>
rect 213 50 214 51 
<< pdiffusion >>
rect 214 50 215 51 
<< pdiffusion >>
rect 215 50 216 51 
<< m1 >>
rect 217 50 218 51 
<< m2 >>
rect 218 50 219 51 
<< pdiffusion >>
rect 228 50 229 51 
<< pdiffusion >>
rect 229 50 230 51 
<< pdiffusion >>
rect 230 50 231 51 
<< pdiffusion >>
rect 231 50 232 51 
<< pdiffusion >>
rect 232 50 233 51 
<< pdiffusion >>
rect 233 50 234 51 
<< pdiffusion >>
rect 246 50 247 51 
<< pdiffusion >>
rect 247 50 248 51 
<< pdiffusion >>
rect 248 50 249 51 
<< pdiffusion >>
rect 249 50 250 51 
<< pdiffusion >>
rect 250 50 251 51 
<< pdiffusion >>
rect 251 50 252 51 
<< m1 >>
rect 253 50 254 51 
<< m1 >>
rect 260 50 261 51 
<< pdiffusion >>
rect 264 50 265 51 
<< pdiffusion >>
rect 265 50 266 51 
<< pdiffusion >>
rect 266 50 267 51 
<< pdiffusion >>
rect 267 50 268 51 
<< pdiffusion >>
rect 268 50 269 51 
<< pdiffusion >>
rect 269 50 270 51 
<< pdiffusion >>
rect 282 50 283 51 
<< pdiffusion >>
rect 283 50 284 51 
<< pdiffusion >>
rect 284 50 285 51 
<< pdiffusion >>
rect 285 50 286 51 
<< pdiffusion >>
rect 286 50 287 51 
<< pdiffusion >>
rect 287 50 288 51 
<< pdiffusion >>
rect 300 50 301 51 
<< pdiffusion >>
rect 301 50 302 51 
<< pdiffusion >>
rect 302 50 303 51 
<< pdiffusion >>
rect 303 50 304 51 
<< pdiffusion >>
rect 304 50 305 51 
<< pdiffusion >>
rect 305 50 306 51 
<< pdiffusion >>
rect 318 50 319 51 
<< pdiffusion >>
rect 319 50 320 51 
<< pdiffusion >>
rect 320 50 321 51 
<< pdiffusion >>
rect 321 50 322 51 
<< pdiffusion >>
rect 322 50 323 51 
<< pdiffusion >>
rect 323 50 324 51 
<< pdiffusion >>
rect 336 50 337 51 
<< pdiffusion >>
rect 337 50 338 51 
<< pdiffusion >>
rect 338 50 339 51 
<< pdiffusion >>
rect 339 50 340 51 
<< pdiffusion >>
rect 340 50 341 51 
<< pdiffusion >>
rect 341 50 342 51 
<< pdiffusion >>
rect 354 50 355 51 
<< pdiffusion >>
rect 355 50 356 51 
<< pdiffusion >>
rect 356 50 357 51 
<< pdiffusion >>
rect 357 50 358 51 
<< pdiffusion >>
rect 358 50 359 51 
<< pdiffusion >>
rect 359 50 360 51 
<< pdiffusion >>
rect 390 50 391 51 
<< pdiffusion >>
rect 391 50 392 51 
<< pdiffusion >>
rect 392 50 393 51 
<< pdiffusion >>
rect 393 50 394 51 
<< pdiffusion >>
rect 394 50 395 51 
<< pdiffusion >>
rect 395 50 396 51 
<< pdiffusion >>
rect 408 50 409 51 
<< pdiffusion >>
rect 409 50 410 51 
<< pdiffusion >>
rect 410 50 411 51 
<< pdiffusion >>
rect 411 50 412 51 
<< pdiffusion >>
rect 412 50 413 51 
<< pdiffusion >>
rect 413 50 414 51 
<< pdiffusion >>
rect 426 50 427 51 
<< pdiffusion >>
rect 427 50 428 51 
<< pdiffusion >>
rect 428 50 429 51 
<< pdiffusion >>
rect 429 50 430 51 
<< pdiffusion >>
rect 430 50 431 51 
<< pdiffusion >>
rect 431 50 432 51 
<< pdiffusion >>
rect 444 50 445 51 
<< pdiffusion >>
rect 445 50 446 51 
<< pdiffusion >>
rect 446 50 447 51 
<< pdiffusion >>
rect 447 50 448 51 
<< pdiffusion >>
rect 448 50 449 51 
<< pdiffusion >>
rect 449 50 450 51 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 64 51 65 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< pdiffusion >>
rect 138 51 139 52 
<< pdiffusion >>
rect 139 51 140 52 
<< pdiffusion >>
rect 140 51 141 52 
<< pdiffusion >>
rect 141 51 142 52 
<< pdiffusion >>
rect 142 51 143 52 
<< pdiffusion >>
rect 143 51 144 52 
<< m1 >>
rect 145 51 146 52 
<< pdiffusion >>
rect 156 51 157 52 
<< pdiffusion >>
rect 157 51 158 52 
<< pdiffusion >>
rect 158 51 159 52 
<< pdiffusion >>
rect 159 51 160 52 
<< pdiffusion >>
rect 160 51 161 52 
<< pdiffusion >>
rect 161 51 162 52 
<< m1 >>
rect 172 51 173 52 
<< pdiffusion >>
rect 174 51 175 52 
<< pdiffusion >>
rect 175 51 176 52 
<< pdiffusion >>
rect 176 51 177 52 
<< pdiffusion >>
rect 177 51 178 52 
<< pdiffusion >>
rect 178 51 179 52 
<< pdiffusion >>
rect 179 51 180 52 
<< pdiffusion >>
rect 192 51 193 52 
<< pdiffusion >>
rect 193 51 194 52 
<< pdiffusion >>
rect 194 51 195 52 
<< pdiffusion >>
rect 195 51 196 52 
<< pdiffusion >>
rect 196 51 197 52 
<< pdiffusion >>
rect 197 51 198 52 
<< pdiffusion >>
rect 210 51 211 52 
<< pdiffusion >>
rect 211 51 212 52 
<< pdiffusion >>
rect 212 51 213 52 
<< pdiffusion >>
rect 213 51 214 52 
<< pdiffusion >>
rect 214 51 215 52 
<< pdiffusion >>
rect 215 51 216 52 
<< m1 >>
rect 217 51 218 52 
<< m2 >>
rect 218 51 219 52 
<< pdiffusion >>
rect 228 51 229 52 
<< pdiffusion >>
rect 229 51 230 52 
<< pdiffusion >>
rect 230 51 231 52 
<< pdiffusion >>
rect 231 51 232 52 
<< pdiffusion >>
rect 232 51 233 52 
<< pdiffusion >>
rect 233 51 234 52 
<< pdiffusion >>
rect 246 51 247 52 
<< pdiffusion >>
rect 247 51 248 52 
<< pdiffusion >>
rect 248 51 249 52 
<< pdiffusion >>
rect 249 51 250 52 
<< pdiffusion >>
rect 250 51 251 52 
<< pdiffusion >>
rect 251 51 252 52 
<< m1 >>
rect 253 51 254 52 
<< m1 >>
rect 260 51 261 52 
<< pdiffusion >>
rect 264 51 265 52 
<< pdiffusion >>
rect 265 51 266 52 
<< pdiffusion >>
rect 266 51 267 52 
<< pdiffusion >>
rect 267 51 268 52 
<< pdiffusion >>
rect 268 51 269 52 
<< pdiffusion >>
rect 269 51 270 52 
<< pdiffusion >>
rect 282 51 283 52 
<< pdiffusion >>
rect 283 51 284 52 
<< pdiffusion >>
rect 284 51 285 52 
<< pdiffusion >>
rect 285 51 286 52 
<< pdiffusion >>
rect 286 51 287 52 
<< pdiffusion >>
rect 287 51 288 52 
<< pdiffusion >>
rect 300 51 301 52 
<< pdiffusion >>
rect 301 51 302 52 
<< pdiffusion >>
rect 302 51 303 52 
<< pdiffusion >>
rect 303 51 304 52 
<< pdiffusion >>
rect 304 51 305 52 
<< pdiffusion >>
rect 305 51 306 52 
<< pdiffusion >>
rect 318 51 319 52 
<< pdiffusion >>
rect 319 51 320 52 
<< pdiffusion >>
rect 320 51 321 52 
<< pdiffusion >>
rect 321 51 322 52 
<< pdiffusion >>
rect 322 51 323 52 
<< pdiffusion >>
rect 323 51 324 52 
<< pdiffusion >>
rect 336 51 337 52 
<< pdiffusion >>
rect 337 51 338 52 
<< pdiffusion >>
rect 338 51 339 52 
<< pdiffusion >>
rect 339 51 340 52 
<< pdiffusion >>
rect 340 51 341 52 
<< pdiffusion >>
rect 341 51 342 52 
<< pdiffusion >>
rect 354 51 355 52 
<< pdiffusion >>
rect 355 51 356 52 
<< pdiffusion >>
rect 356 51 357 52 
<< pdiffusion >>
rect 357 51 358 52 
<< pdiffusion >>
rect 358 51 359 52 
<< pdiffusion >>
rect 359 51 360 52 
<< pdiffusion >>
rect 390 51 391 52 
<< pdiffusion >>
rect 391 51 392 52 
<< pdiffusion >>
rect 392 51 393 52 
<< pdiffusion >>
rect 393 51 394 52 
<< pdiffusion >>
rect 394 51 395 52 
<< pdiffusion >>
rect 395 51 396 52 
<< pdiffusion >>
rect 408 51 409 52 
<< pdiffusion >>
rect 409 51 410 52 
<< pdiffusion >>
rect 410 51 411 52 
<< pdiffusion >>
rect 411 51 412 52 
<< pdiffusion >>
rect 412 51 413 52 
<< pdiffusion >>
rect 413 51 414 52 
<< pdiffusion >>
rect 426 51 427 52 
<< pdiffusion >>
rect 427 51 428 52 
<< pdiffusion >>
rect 428 51 429 52 
<< pdiffusion >>
rect 429 51 430 52 
<< pdiffusion >>
rect 430 51 431 52 
<< pdiffusion >>
rect 431 51 432 52 
<< pdiffusion >>
rect 444 51 445 52 
<< pdiffusion >>
rect 445 51 446 52 
<< pdiffusion >>
rect 446 51 447 52 
<< pdiffusion >>
rect 447 51 448 52 
<< pdiffusion >>
rect 448 51 449 52 
<< pdiffusion >>
rect 449 51 450 52 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 64 52 65 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< pdiffusion >>
rect 138 52 139 53 
<< pdiffusion >>
rect 139 52 140 53 
<< pdiffusion >>
rect 140 52 141 53 
<< pdiffusion >>
rect 141 52 142 53 
<< pdiffusion >>
rect 142 52 143 53 
<< pdiffusion >>
rect 143 52 144 53 
<< m1 >>
rect 145 52 146 53 
<< pdiffusion >>
rect 156 52 157 53 
<< pdiffusion >>
rect 157 52 158 53 
<< pdiffusion >>
rect 158 52 159 53 
<< pdiffusion >>
rect 159 52 160 53 
<< pdiffusion >>
rect 160 52 161 53 
<< pdiffusion >>
rect 161 52 162 53 
<< m1 >>
rect 172 52 173 53 
<< pdiffusion >>
rect 174 52 175 53 
<< pdiffusion >>
rect 175 52 176 53 
<< pdiffusion >>
rect 176 52 177 53 
<< pdiffusion >>
rect 177 52 178 53 
<< pdiffusion >>
rect 178 52 179 53 
<< pdiffusion >>
rect 179 52 180 53 
<< pdiffusion >>
rect 192 52 193 53 
<< pdiffusion >>
rect 193 52 194 53 
<< pdiffusion >>
rect 194 52 195 53 
<< pdiffusion >>
rect 195 52 196 53 
<< pdiffusion >>
rect 196 52 197 53 
<< pdiffusion >>
rect 197 52 198 53 
<< pdiffusion >>
rect 210 52 211 53 
<< pdiffusion >>
rect 211 52 212 53 
<< pdiffusion >>
rect 212 52 213 53 
<< pdiffusion >>
rect 213 52 214 53 
<< pdiffusion >>
rect 214 52 215 53 
<< pdiffusion >>
rect 215 52 216 53 
<< m1 >>
rect 217 52 218 53 
<< m2 >>
rect 218 52 219 53 
<< pdiffusion >>
rect 228 52 229 53 
<< pdiffusion >>
rect 229 52 230 53 
<< pdiffusion >>
rect 230 52 231 53 
<< pdiffusion >>
rect 231 52 232 53 
<< pdiffusion >>
rect 232 52 233 53 
<< pdiffusion >>
rect 233 52 234 53 
<< pdiffusion >>
rect 246 52 247 53 
<< pdiffusion >>
rect 247 52 248 53 
<< pdiffusion >>
rect 248 52 249 53 
<< pdiffusion >>
rect 249 52 250 53 
<< pdiffusion >>
rect 250 52 251 53 
<< pdiffusion >>
rect 251 52 252 53 
<< m1 >>
rect 253 52 254 53 
<< m1 >>
rect 260 52 261 53 
<< pdiffusion >>
rect 264 52 265 53 
<< pdiffusion >>
rect 265 52 266 53 
<< pdiffusion >>
rect 266 52 267 53 
<< pdiffusion >>
rect 267 52 268 53 
<< pdiffusion >>
rect 268 52 269 53 
<< pdiffusion >>
rect 269 52 270 53 
<< pdiffusion >>
rect 282 52 283 53 
<< pdiffusion >>
rect 283 52 284 53 
<< pdiffusion >>
rect 284 52 285 53 
<< pdiffusion >>
rect 285 52 286 53 
<< pdiffusion >>
rect 286 52 287 53 
<< pdiffusion >>
rect 287 52 288 53 
<< pdiffusion >>
rect 300 52 301 53 
<< pdiffusion >>
rect 301 52 302 53 
<< pdiffusion >>
rect 302 52 303 53 
<< pdiffusion >>
rect 303 52 304 53 
<< pdiffusion >>
rect 304 52 305 53 
<< pdiffusion >>
rect 305 52 306 53 
<< pdiffusion >>
rect 318 52 319 53 
<< pdiffusion >>
rect 319 52 320 53 
<< pdiffusion >>
rect 320 52 321 53 
<< pdiffusion >>
rect 321 52 322 53 
<< pdiffusion >>
rect 322 52 323 53 
<< pdiffusion >>
rect 323 52 324 53 
<< pdiffusion >>
rect 336 52 337 53 
<< pdiffusion >>
rect 337 52 338 53 
<< pdiffusion >>
rect 338 52 339 53 
<< pdiffusion >>
rect 339 52 340 53 
<< pdiffusion >>
rect 340 52 341 53 
<< pdiffusion >>
rect 341 52 342 53 
<< pdiffusion >>
rect 354 52 355 53 
<< pdiffusion >>
rect 355 52 356 53 
<< pdiffusion >>
rect 356 52 357 53 
<< pdiffusion >>
rect 357 52 358 53 
<< pdiffusion >>
rect 358 52 359 53 
<< pdiffusion >>
rect 359 52 360 53 
<< pdiffusion >>
rect 390 52 391 53 
<< pdiffusion >>
rect 391 52 392 53 
<< pdiffusion >>
rect 392 52 393 53 
<< pdiffusion >>
rect 393 52 394 53 
<< pdiffusion >>
rect 394 52 395 53 
<< pdiffusion >>
rect 395 52 396 53 
<< pdiffusion >>
rect 408 52 409 53 
<< pdiffusion >>
rect 409 52 410 53 
<< pdiffusion >>
rect 410 52 411 53 
<< pdiffusion >>
rect 411 52 412 53 
<< pdiffusion >>
rect 412 52 413 53 
<< pdiffusion >>
rect 413 52 414 53 
<< pdiffusion >>
rect 426 52 427 53 
<< pdiffusion >>
rect 427 52 428 53 
<< pdiffusion >>
rect 428 52 429 53 
<< pdiffusion >>
rect 429 52 430 53 
<< pdiffusion >>
rect 430 52 431 53 
<< pdiffusion >>
rect 431 52 432 53 
<< pdiffusion >>
rect 444 52 445 53 
<< pdiffusion >>
rect 445 52 446 53 
<< pdiffusion >>
rect 446 52 447 53 
<< pdiffusion >>
rect 447 52 448 53 
<< pdiffusion >>
rect 448 52 449 53 
<< pdiffusion >>
rect 449 52 450 53 
<< pdiffusion >>
rect 12 53 13 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< pdiffusion >>
rect 30 53 31 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< pdiffusion >>
rect 48 53 49 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 64 53 65 54 
<< pdiffusion >>
rect 66 53 67 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< pdiffusion >>
rect 84 53 85 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< pdiffusion >>
rect 102 53 103 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< pdiffusion >>
rect 120 53 121 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< pdiffusion >>
rect 138 53 139 54 
<< pdiffusion >>
rect 139 53 140 54 
<< pdiffusion >>
rect 140 53 141 54 
<< pdiffusion >>
rect 141 53 142 54 
<< m1 >>
rect 142 53 143 54 
<< pdiffusion >>
rect 142 53 143 54 
<< pdiffusion >>
rect 143 53 144 54 
<< m1 >>
rect 145 53 146 54 
<< pdiffusion >>
rect 156 53 157 54 
<< pdiffusion >>
rect 157 53 158 54 
<< pdiffusion >>
rect 158 53 159 54 
<< pdiffusion >>
rect 159 53 160 54 
<< m1 >>
rect 160 53 161 54 
<< pdiffusion >>
rect 160 53 161 54 
<< pdiffusion >>
rect 161 53 162 54 
<< m1 >>
rect 172 53 173 54 
<< pdiffusion >>
rect 174 53 175 54 
<< pdiffusion >>
rect 175 53 176 54 
<< pdiffusion >>
rect 176 53 177 54 
<< pdiffusion >>
rect 177 53 178 54 
<< pdiffusion >>
rect 178 53 179 54 
<< pdiffusion >>
rect 179 53 180 54 
<< pdiffusion >>
rect 192 53 193 54 
<< pdiffusion >>
rect 193 53 194 54 
<< pdiffusion >>
rect 194 53 195 54 
<< pdiffusion >>
rect 195 53 196 54 
<< m1 >>
rect 196 53 197 54 
<< pdiffusion >>
rect 196 53 197 54 
<< pdiffusion >>
rect 197 53 198 54 
<< pdiffusion >>
rect 210 53 211 54 
<< pdiffusion >>
rect 211 53 212 54 
<< pdiffusion >>
rect 212 53 213 54 
<< pdiffusion >>
rect 213 53 214 54 
<< m1 >>
rect 214 53 215 54 
<< pdiffusion >>
rect 214 53 215 54 
<< pdiffusion >>
rect 215 53 216 54 
<< m1 >>
rect 217 53 218 54 
<< m2 >>
rect 218 53 219 54 
<< pdiffusion >>
rect 228 53 229 54 
<< pdiffusion >>
rect 229 53 230 54 
<< pdiffusion >>
rect 230 53 231 54 
<< pdiffusion >>
rect 231 53 232 54 
<< pdiffusion >>
rect 232 53 233 54 
<< pdiffusion >>
rect 233 53 234 54 
<< pdiffusion >>
rect 246 53 247 54 
<< m1 >>
rect 247 53 248 54 
<< pdiffusion >>
rect 247 53 248 54 
<< pdiffusion >>
rect 248 53 249 54 
<< pdiffusion >>
rect 249 53 250 54 
<< pdiffusion >>
rect 250 53 251 54 
<< pdiffusion >>
rect 251 53 252 54 
<< m1 >>
rect 253 53 254 54 
<< m1 >>
rect 260 53 261 54 
<< pdiffusion >>
rect 264 53 265 54 
<< pdiffusion >>
rect 265 53 266 54 
<< pdiffusion >>
rect 266 53 267 54 
<< pdiffusion >>
rect 267 53 268 54 
<< pdiffusion >>
rect 268 53 269 54 
<< pdiffusion >>
rect 269 53 270 54 
<< pdiffusion >>
rect 282 53 283 54 
<< pdiffusion >>
rect 283 53 284 54 
<< pdiffusion >>
rect 284 53 285 54 
<< pdiffusion >>
rect 285 53 286 54 
<< m1 >>
rect 286 53 287 54 
<< pdiffusion >>
rect 286 53 287 54 
<< pdiffusion >>
rect 287 53 288 54 
<< pdiffusion >>
rect 300 53 301 54 
<< pdiffusion >>
rect 301 53 302 54 
<< pdiffusion >>
rect 302 53 303 54 
<< pdiffusion >>
rect 303 53 304 54 
<< pdiffusion >>
rect 304 53 305 54 
<< pdiffusion >>
rect 305 53 306 54 
<< pdiffusion >>
rect 318 53 319 54 
<< pdiffusion >>
rect 319 53 320 54 
<< pdiffusion >>
rect 320 53 321 54 
<< pdiffusion >>
rect 321 53 322 54 
<< pdiffusion >>
rect 322 53 323 54 
<< pdiffusion >>
rect 323 53 324 54 
<< pdiffusion >>
rect 336 53 337 54 
<< pdiffusion >>
rect 337 53 338 54 
<< pdiffusion >>
rect 338 53 339 54 
<< pdiffusion >>
rect 339 53 340 54 
<< pdiffusion >>
rect 340 53 341 54 
<< pdiffusion >>
rect 341 53 342 54 
<< pdiffusion >>
rect 354 53 355 54 
<< pdiffusion >>
rect 355 53 356 54 
<< pdiffusion >>
rect 356 53 357 54 
<< pdiffusion >>
rect 357 53 358 54 
<< pdiffusion >>
rect 358 53 359 54 
<< pdiffusion >>
rect 359 53 360 54 
<< pdiffusion >>
rect 390 53 391 54 
<< pdiffusion >>
rect 391 53 392 54 
<< pdiffusion >>
rect 392 53 393 54 
<< pdiffusion >>
rect 393 53 394 54 
<< pdiffusion >>
rect 394 53 395 54 
<< pdiffusion >>
rect 395 53 396 54 
<< pdiffusion >>
rect 408 53 409 54 
<< pdiffusion >>
rect 409 53 410 54 
<< pdiffusion >>
rect 410 53 411 54 
<< pdiffusion >>
rect 411 53 412 54 
<< pdiffusion >>
rect 412 53 413 54 
<< pdiffusion >>
rect 413 53 414 54 
<< pdiffusion >>
rect 426 53 427 54 
<< pdiffusion >>
rect 427 53 428 54 
<< pdiffusion >>
rect 428 53 429 54 
<< pdiffusion >>
rect 429 53 430 54 
<< pdiffusion >>
rect 430 53 431 54 
<< pdiffusion >>
rect 431 53 432 54 
<< pdiffusion >>
rect 444 53 445 54 
<< pdiffusion >>
rect 445 53 446 54 
<< pdiffusion >>
rect 446 53 447 54 
<< pdiffusion >>
rect 447 53 448 54 
<< pdiffusion >>
rect 448 53 449 54 
<< pdiffusion >>
rect 449 53 450 54 
<< m1 >>
rect 64 54 65 55 
<< m1 >>
rect 91 54 92 55 
<< m1 >>
rect 142 54 143 55 
<< m1 >>
rect 145 54 146 55 
<< m1 >>
rect 160 54 161 55 
<< m1 >>
rect 172 54 173 55 
<< m1 >>
rect 196 54 197 55 
<< m1 >>
rect 214 54 215 55 
<< m1 >>
rect 217 54 218 55 
<< m2 >>
rect 218 54 219 55 
<< m1 >>
rect 247 54 248 55 
<< m1 >>
rect 253 54 254 55 
<< m1 >>
rect 260 54 261 55 
<< m1 >>
rect 286 54 287 55 
<< m1 >>
rect 64 55 65 56 
<< m1 >>
rect 91 55 92 56 
<< m1 >>
rect 142 55 143 56 
<< m1 >>
rect 145 55 146 56 
<< m1 >>
rect 160 55 161 56 
<< m1 >>
rect 161 55 162 56 
<< m1 >>
rect 162 55 163 56 
<< m1 >>
rect 163 55 164 56 
<< m1 >>
rect 164 55 165 56 
<< m1 >>
rect 165 55 166 56 
<< m1 >>
rect 166 55 167 56 
<< m1 >>
rect 167 55 168 56 
<< m1 >>
rect 168 55 169 56 
<< m1 >>
rect 169 55 170 56 
<< m1 >>
rect 170 55 171 56 
<< m1 >>
rect 171 55 172 56 
<< m1 >>
rect 172 55 173 56 
<< m1 >>
rect 196 55 197 56 
<< m1 >>
rect 214 55 215 56 
<< m1 >>
rect 217 55 218 56 
<< m2 >>
rect 218 55 219 56 
<< m1 >>
rect 247 55 248 56 
<< m1 >>
rect 253 55 254 56 
<< m1 >>
rect 260 55 261 56 
<< m1 >>
rect 286 55 287 56 
<< m1 >>
rect 64 56 65 57 
<< m1 >>
rect 91 56 92 57 
<< m1 >>
rect 142 56 143 57 
<< m1 >>
rect 145 56 146 57 
<< m1 >>
rect 196 56 197 57 
<< m1 >>
rect 214 56 215 57 
<< m1 >>
rect 217 56 218 57 
<< m2 >>
rect 218 56 219 57 
<< m1 >>
rect 247 56 248 57 
<< m1 >>
rect 248 56 249 57 
<< m1 >>
rect 249 56 250 57 
<< m1 >>
rect 250 56 251 57 
<< m1 >>
rect 251 56 252 57 
<< m1 >>
rect 252 56 253 57 
<< m1 >>
rect 253 56 254 57 
<< m1 >>
rect 260 56 261 57 
<< m1 >>
rect 286 56 287 57 
<< m1 >>
rect 64 57 65 58 
<< m1 >>
rect 91 57 92 58 
<< m1 >>
rect 142 57 143 58 
<< m1 >>
rect 145 57 146 58 
<< m1 >>
rect 196 57 197 58 
<< m1 >>
rect 214 57 215 58 
<< m1 >>
rect 217 57 218 58 
<< m2 >>
rect 218 57 219 58 
<< m1 >>
rect 260 57 261 58 
<< m1 >>
rect 286 57 287 58 
<< m1 >>
rect 64 58 65 59 
<< m1 >>
rect 91 58 92 59 
<< m1 >>
rect 142 58 143 59 
<< m1 >>
rect 145 58 146 59 
<< m1 >>
rect 196 58 197 59 
<< m1 >>
rect 214 58 215 59 
<< m1 >>
rect 217 58 218 59 
<< m2 >>
rect 218 58 219 59 
<< m1 >>
rect 260 58 261 59 
<< m1 >>
rect 262 58 263 59 
<< m1 >>
rect 263 58 264 59 
<< m1 >>
rect 264 58 265 59 
<< m1 >>
rect 265 58 266 59 
<< m1 >>
rect 266 58 267 59 
<< m1 >>
rect 267 58 268 59 
<< m1 >>
rect 268 58 269 59 
<< m1 >>
rect 269 58 270 59 
<< m1 >>
rect 270 58 271 59 
<< m1 >>
rect 271 58 272 59 
<< m1 >>
rect 272 58 273 59 
<< m1 >>
rect 273 58 274 59 
<< m1 >>
rect 274 58 275 59 
<< m1 >>
rect 275 58 276 59 
<< m1 >>
rect 276 58 277 59 
<< m1 >>
rect 277 58 278 59 
<< m1 >>
rect 278 58 279 59 
<< m1 >>
rect 279 58 280 59 
<< m1 >>
rect 280 58 281 59 
<< m1 >>
rect 281 58 282 59 
<< m1 >>
rect 282 58 283 59 
<< m1 >>
rect 283 58 284 59 
<< m1 >>
rect 284 58 285 59 
<< m1 >>
rect 285 58 286 59 
<< m1 >>
rect 286 58 287 59 
<< m1 >>
rect 64 59 65 60 
<< m1 >>
rect 91 59 92 60 
<< m1 >>
rect 142 59 143 60 
<< m1 >>
rect 145 59 146 60 
<< m1 >>
rect 196 59 197 60 
<< m2 >>
rect 196 59 197 60 
<< m2c >>
rect 196 59 197 60 
<< m1 >>
rect 196 59 197 60 
<< m2 >>
rect 196 59 197 60 
<< m1 >>
rect 214 59 215 60 
<< m1 >>
rect 217 59 218 60 
<< m2 >>
rect 218 59 219 60 
<< m1 >>
rect 260 59 261 60 
<< m1 >>
rect 262 59 263 60 
<< m1 >>
rect 64 60 65 61 
<< m1 >>
rect 91 60 92 61 
<< m1 >>
rect 142 60 143 61 
<< m1 >>
rect 145 60 146 61 
<< m2 >>
rect 196 60 197 61 
<< m2 >>
rect 210 60 211 61 
<< m2 >>
rect 211 60 212 61 
<< m2 >>
rect 212 60 213 61 
<< m2 >>
rect 213 60 214 61 
<< m1 >>
rect 214 60 215 61 
<< m2 >>
rect 214 60 215 61 
<< m2 >>
rect 215 60 216 61 
<< m2 >>
rect 216 60 217 61 
<< m1 >>
rect 217 60 218 61 
<< m2 >>
rect 217 60 218 61 
<< m2 >>
rect 218 60 219 61 
<< m1 >>
rect 260 60 261 61 
<< m1 >>
rect 262 60 263 61 
<< m1 >>
rect 64 61 65 62 
<< m1 >>
rect 91 61 92 62 
<< m1 >>
rect 142 61 143 62 
<< m1 >>
rect 145 61 146 62 
<< m2 >>
rect 145 61 146 62 
<< m2c >>
rect 145 61 146 62 
<< m1 >>
rect 145 61 146 62 
<< m2 >>
rect 145 61 146 62 
<< m1 >>
rect 181 61 182 62 
<< m1 >>
rect 182 61 183 62 
<< m1 >>
rect 183 61 184 62 
<< m1 >>
rect 184 61 185 62 
<< m1 >>
rect 185 61 186 62 
<< m1 >>
rect 186 61 187 62 
<< m1 >>
rect 187 61 188 62 
<< m1 >>
rect 188 61 189 62 
<< m1 >>
rect 189 61 190 62 
<< m1 >>
rect 190 61 191 62 
<< m1 >>
rect 191 61 192 62 
<< m1 >>
rect 192 61 193 62 
<< m1 >>
rect 193 61 194 62 
<< m1 >>
rect 194 61 195 62 
<< m1 >>
rect 195 61 196 62 
<< m1 >>
rect 196 61 197 62 
<< m2 >>
rect 196 61 197 62 
<< m1 >>
rect 197 61 198 62 
<< m1 >>
rect 198 61 199 62 
<< m1 >>
rect 199 61 200 62 
<< m1 >>
rect 200 61 201 62 
<< m1 >>
rect 201 61 202 62 
<< m1 >>
rect 202 61 203 62 
<< m1 >>
rect 203 61 204 62 
<< m1 >>
rect 204 61 205 62 
<< m1 >>
rect 205 61 206 62 
<< m1 >>
rect 206 61 207 62 
<< m1 >>
rect 207 61 208 62 
<< m1 >>
rect 208 61 209 62 
<< m1 >>
rect 209 61 210 62 
<< m1 >>
rect 210 61 211 62 
<< m2 >>
rect 210 61 211 62 
<< m1 >>
rect 211 61 212 62 
<< m1 >>
rect 212 61 213 62 
<< m1 >>
rect 213 61 214 62 
<< m1 >>
rect 214 61 215 62 
<< m1 >>
rect 217 61 218 62 
<< m1 >>
rect 221 61 222 62 
<< m1 >>
rect 222 61 223 62 
<< m1 >>
rect 223 61 224 62 
<< m1 >>
rect 224 61 225 62 
<< m1 >>
rect 225 61 226 62 
<< m1 >>
rect 226 61 227 62 
<< m1 >>
rect 227 61 228 62 
<< m1 >>
rect 228 61 229 62 
<< m1 >>
rect 229 61 230 62 
<< m1 >>
rect 230 61 231 62 
<< m1 >>
rect 231 61 232 62 
<< m1 >>
rect 232 61 233 62 
<< m1 >>
rect 260 61 261 62 
<< m1 >>
rect 262 61 263 62 
<< m1 >>
rect 64 62 65 63 
<< m1 >>
rect 91 62 92 63 
<< m1 >>
rect 142 62 143 63 
<< m2 >>
rect 145 62 146 63 
<< m1 >>
rect 181 62 182 63 
<< m2 >>
rect 196 62 197 63 
<< m2 >>
rect 210 62 211 63 
<< m1 >>
rect 217 62 218 63 
<< m1 >>
rect 221 62 222 63 
<< m1 >>
rect 232 62 233 63 
<< m1 >>
rect 260 62 261 63 
<< m1 >>
rect 262 62 263 63 
<< m1 >>
rect 64 63 65 64 
<< m1 >>
rect 91 63 92 64 
<< m1 >>
rect 142 63 143 64 
<< m1 >>
rect 143 63 144 64 
<< m1 >>
rect 144 63 145 64 
<< m1 >>
rect 145 63 146 64 
<< m2 >>
rect 145 63 146 64 
<< m1 >>
rect 146 63 147 64 
<< m1 >>
rect 147 63 148 64 
<< m1 >>
rect 148 63 149 64 
<< m1 >>
rect 149 63 150 64 
<< m1 >>
rect 150 63 151 64 
<< m1 >>
rect 151 63 152 64 
<< m1 >>
rect 152 63 153 64 
<< m1 >>
rect 153 63 154 64 
<< m1 >>
rect 154 63 155 64 
<< m1 >>
rect 181 63 182 64 
<< m1 >>
rect 196 63 197 64 
<< m2 >>
rect 196 63 197 64 
<< m2c >>
rect 196 63 197 64 
<< m1 >>
rect 196 63 197 64 
<< m2 >>
rect 196 63 197 64 
<< m1 >>
rect 197 63 198 64 
<< m1 >>
rect 198 63 199 64 
<< m1 >>
rect 199 63 200 64 
<< m1 >>
rect 200 63 201 64 
<< m1 >>
rect 201 63 202 64 
<< m1 >>
rect 202 63 203 64 
<< m1 >>
rect 203 63 204 64 
<< m1 >>
rect 208 63 209 64 
<< m1 >>
rect 209 63 210 64 
<< m1 >>
rect 210 63 211 64 
<< m2 >>
rect 210 63 211 64 
<< m2c >>
rect 210 63 211 64 
<< m1 >>
rect 210 63 211 64 
<< m2 >>
rect 210 63 211 64 
<< m1 >>
rect 217 63 218 64 
<< m1 >>
rect 221 63 222 64 
<< m1 >>
rect 232 63 233 64 
<< m1 >>
rect 260 63 261 64 
<< m1 >>
rect 262 63 263 64 
<< m1 >>
rect 64 64 65 65 
<< m1 >>
rect 91 64 92 65 
<< m2 >>
rect 145 64 146 65 
<< m1 >>
rect 154 64 155 65 
<< m1 >>
rect 181 64 182 65 
<< m1 >>
rect 203 64 204 65 
<< m1 >>
rect 208 64 209 65 
<< m1 >>
rect 217 64 218 65 
<< m1 >>
rect 221 64 222 65 
<< m1 >>
rect 232 64 233 65 
<< m1 >>
rect 260 64 261 65 
<< m1 >>
rect 262 64 263 65 
<< m1 >>
rect 64 65 65 66 
<< m1 >>
rect 91 65 92 66 
<< m1 >>
rect 145 65 146 66 
<< m2 >>
rect 145 65 146 66 
<< m2c >>
rect 145 65 146 66 
<< m1 >>
rect 145 65 146 66 
<< m2 >>
rect 145 65 146 66 
<< m1 >>
rect 154 65 155 66 
<< m1 >>
rect 181 65 182 66 
<< m1 >>
rect 203 65 204 66 
<< m1 >>
rect 208 65 209 66 
<< m1 >>
rect 217 65 218 66 
<< m1 >>
rect 221 65 222 66 
<< m1 >>
rect 232 65 233 66 
<< m1 >>
rect 260 65 261 66 
<< m1 >>
rect 262 65 263 66 
<< pdiffusion >>
rect 12 66 13 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< pdiffusion >>
rect 30 66 31 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< pdiffusion >>
rect 48 66 49 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 64 66 65 67 
<< pdiffusion >>
rect 66 66 67 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< pdiffusion >>
rect 84 66 85 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< m1 >>
rect 91 66 92 67 
<< pdiffusion >>
rect 102 66 103 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< pdiffusion >>
rect 120 66 121 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< pdiffusion >>
rect 138 66 139 67 
<< pdiffusion >>
rect 139 66 140 67 
<< pdiffusion >>
rect 140 66 141 67 
<< pdiffusion >>
rect 141 66 142 67 
<< pdiffusion >>
rect 142 66 143 67 
<< pdiffusion >>
rect 143 66 144 67 
<< m1 >>
rect 145 66 146 67 
<< m1 >>
rect 154 66 155 67 
<< pdiffusion >>
rect 156 66 157 67 
<< pdiffusion >>
rect 157 66 158 67 
<< pdiffusion >>
rect 158 66 159 67 
<< pdiffusion >>
rect 159 66 160 67 
<< pdiffusion >>
rect 160 66 161 67 
<< pdiffusion >>
rect 161 66 162 67 
<< pdiffusion >>
rect 174 66 175 67 
<< pdiffusion >>
rect 175 66 176 67 
<< pdiffusion >>
rect 176 66 177 67 
<< pdiffusion >>
rect 177 66 178 67 
<< pdiffusion >>
rect 178 66 179 67 
<< pdiffusion >>
rect 179 66 180 67 
<< m1 >>
rect 181 66 182 67 
<< pdiffusion >>
rect 192 66 193 67 
<< pdiffusion >>
rect 193 66 194 67 
<< pdiffusion >>
rect 194 66 195 67 
<< pdiffusion >>
rect 195 66 196 67 
<< pdiffusion >>
rect 196 66 197 67 
<< pdiffusion >>
rect 197 66 198 67 
<< m1 >>
rect 203 66 204 67 
<< m1 >>
rect 208 66 209 67 
<< pdiffusion >>
rect 210 66 211 67 
<< pdiffusion >>
rect 211 66 212 67 
<< pdiffusion >>
rect 212 66 213 67 
<< pdiffusion >>
rect 213 66 214 67 
<< pdiffusion >>
rect 214 66 215 67 
<< pdiffusion >>
rect 215 66 216 67 
<< m1 >>
rect 217 66 218 67 
<< m1 >>
rect 221 66 222 67 
<< pdiffusion >>
rect 228 66 229 67 
<< pdiffusion >>
rect 229 66 230 67 
<< pdiffusion >>
rect 230 66 231 67 
<< pdiffusion >>
rect 231 66 232 67 
<< m1 >>
rect 232 66 233 67 
<< pdiffusion >>
rect 232 66 233 67 
<< pdiffusion >>
rect 233 66 234 67 
<< pdiffusion >>
rect 246 66 247 67 
<< pdiffusion >>
rect 247 66 248 67 
<< pdiffusion >>
rect 248 66 249 67 
<< pdiffusion >>
rect 249 66 250 67 
<< pdiffusion >>
rect 250 66 251 67 
<< pdiffusion >>
rect 251 66 252 67 
<< m1 >>
rect 260 66 261 67 
<< m1 >>
rect 262 66 263 67 
<< pdiffusion >>
rect 264 66 265 67 
<< pdiffusion >>
rect 265 66 266 67 
<< pdiffusion >>
rect 266 66 267 67 
<< pdiffusion >>
rect 267 66 268 67 
<< pdiffusion >>
rect 268 66 269 67 
<< pdiffusion >>
rect 269 66 270 67 
<< pdiffusion >>
rect 282 66 283 67 
<< pdiffusion >>
rect 283 66 284 67 
<< pdiffusion >>
rect 284 66 285 67 
<< pdiffusion >>
rect 285 66 286 67 
<< pdiffusion >>
rect 286 66 287 67 
<< pdiffusion >>
rect 287 66 288 67 
<< pdiffusion >>
rect 300 66 301 67 
<< pdiffusion >>
rect 301 66 302 67 
<< pdiffusion >>
rect 302 66 303 67 
<< pdiffusion >>
rect 303 66 304 67 
<< pdiffusion >>
rect 304 66 305 67 
<< pdiffusion >>
rect 305 66 306 67 
<< pdiffusion >>
rect 336 66 337 67 
<< pdiffusion >>
rect 337 66 338 67 
<< pdiffusion >>
rect 338 66 339 67 
<< pdiffusion >>
rect 339 66 340 67 
<< pdiffusion >>
rect 340 66 341 67 
<< pdiffusion >>
rect 341 66 342 67 
<< pdiffusion >>
rect 354 66 355 67 
<< pdiffusion >>
rect 355 66 356 67 
<< pdiffusion >>
rect 356 66 357 67 
<< pdiffusion >>
rect 357 66 358 67 
<< pdiffusion >>
rect 358 66 359 67 
<< pdiffusion >>
rect 359 66 360 67 
<< pdiffusion >>
rect 372 66 373 67 
<< pdiffusion >>
rect 373 66 374 67 
<< pdiffusion >>
rect 374 66 375 67 
<< pdiffusion >>
rect 375 66 376 67 
<< pdiffusion >>
rect 376 66 377 67 
<< pdiffusion >>
rect 377 66 378 67 
<< pdiffusion >>
rect 390 66 391 67 
<< pdiffusion >>
rect 391 66 392 67 
<< pdiffusion >>
rect 392 66 393 67 
<< pdiffusion >>
rect 393 66 394 67 
<< pdiffusion >>
rect 394 66 395 67 
<< pdiffusion >>
rect 395 66 396 67 
<< pdiffusion >>
rect 408 66 409 67 
<< pdiffusion >>
rect 409 66 410 67 
<< pdiffusion >>
rect 410 66 411 67 
<< pdiffusion >>
rect 411 66 412 67 
<< pdiffusion >>
rect 412 66 413 67 
<< pdiffusion >>
rect 413 66 414 67 
<< pdiffusion >>
rect 426 66 427 67 
<< pdiffusion >>
rect 427 66 428 67 
<< pdiffusion >>
rect 428 66 429 67 
<< pdiffusion >>
rect 429 66 430 67 
<< pdiffusion >>
rect 430 66 431 67 
<< pdiffusion >>
rect 431 66 432 67 
<< pdiffusion >>
rect 444 66 445 67 
<< pdiffusion >>
rect 445 66 446 67 
<< pdiffusion >>
rect 446 66 447 67 
<< pdiffusion >>
rect 447 66 448 67 
<< pdiffusion >>
rect 448 66 449 67 
<< pdiffusion >>
rect 449 66 450 67 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 64 67 65 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< m1 >>
rect 91 67 92 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< pdiffusion >>
rect 138 67 139 68 
<< pdiffusion >>
rect 139 67 140 68 
<< pdiffusion >>
rect 140 67 141 68 
<< pdiffusion >>
rect 141 67 142 68 
<< pdiffusion >>
rect 142 67 143 68 
<< pdiffusion >>
rect 143 67 144 68 
<< m1 >>
rect 145 67 146 68 
<< m1 >>
rect 154 67 155 68 
<< pdiffusion >>
rect 156 67 157 68 
<< pdiffusion >>
rect 157 67 158 68 
<< pdiffusion >>
rect 158 67 159 68 
<< pdiffusion >>
rect 159 67 160 68 
<< pdiffusion >>
rect 160 67 161 68 
<< pdiffusion >>
rect 161 67 162 68 
<< pdiffusion >>
rect 174 67 175 68 
<< pdiffusion >>
rect 175 67 176 68 
<< pdiffusion >>
rect 176 67 177 68 
<< pdiffusion >>
rect 177 67 178 68 
<< pdiffusion >>
rect 178 67 179 68 
<< pdiffusion >>
rect 179 67 180 68 
<< m1 >>
rect 181 67 182 68 
<< pdiffusion >>
rect 192 67 193 68 
<< pdiffusion >>
rect 193 67 194 68 
<< pdiffusion >>
rect 194 67 195 68 
<< pdiffusion >>
rect 195 67 196 68 
<< pdiffusion >>
rect 196 67 197 68 
<< pdiffusion >>
rect 197 67 198 68 
<< m1 >>
rect 203 67 204 68 
<< m1 >>
rect 208 67 209 68 
<< pdiffusion >>
rect 210 67 211 68 
<< pdiffusion >>
rect 211 67 212 68 
<< pdiffusion >>
rect 212 67 213 68 
<< pdiffusion >>
rect 213 67 214 68 
<< pdiffusion >>
rect 214 67 215 68 
<< pdiffusion >>
rect 215 67 216 68 
<< m1 >>
rect 217 67 218 68 
<< m1 >>
rect 221 67 222 68 
<< pdiffusion >>
rect 228 67 229 68 
<< pdiffusion >>
rect 229 67 230 68 
<< pdiffusion >>
rect 230 67 231 68 
<< pdiffusion >>
rect 231 67 232 68 
<< pdiffusion >>
rect 232 67 233 68 
<< pdiffusion >>
rect 233 67 234 68 
<< pdiffusion >>
rect 246 67 247 68 
<< pdiffusion >>
rect 247 67 248 68 
<< pdiffusion >>
rect 248 67 249 68 
<< pdiffusion >>
rect 249 67 250 68 
<< pdiffusion >>
rect 250 67 251 68 
<< pdiffusion >>
rect 251 67 252 68 
<< m1 >>
rect 260 67 261 68 
<< m1 >>
rect 262 67 263 68 
<< pdiffusion >>
rect 264 67 265 68 
<< pdiffusion >>
rect 265 67 266 68 
<< pdiffusion >>
rect 266 67 267 68 
<< pdiffusion >>
rect 267 67 268 68 
<< pdiffusion >>
rect 268 67 269 68 
<< pdiffusion >>
rect 269 67 270 68 
<< pdiffusion >>
rect 282 67 283 68 
<< pdiffusion >>
rect 283 67 284 68 
<< pdiffusion >>
rect 284 67 285 68 
<< pdiffusion >>
rect 285 67 286 68 
<< pdiffusion >>
rect 286 67 287 68 
<< pdiffusion >>
rect 287 67 288 68 
<< pdiffusion >>
rect 300 67 301 68 
<< pdiffusion >>
rect 301 67 302 68 
<< pdiffusion >>
rect 302 67 303 68 
<< pdiffusion >>
rect 303 67 304 68 
<< pdiffusion >>
rect 304 67 305 68 
<< pdiffusion >>
rect 305 67 306 68 
<< pdiffusion >>
rect 336 67 337 68 
<< pdiffusion >>
rect 337 67 338 68 
<< pdiffusion >>
rect 338 67 339 68 
<< pdiffusion >>
rect 339 67 340 68 
<< pdiffusion >>
rect 340 67 341 68 
<< pdiffusion >>
rect 341 67 342 68 
<< pdiffusion >>
rect 354 67 355 68 
<< pdiffusion >>
rect 355 67 356 68 
<< pdiffusion >>
rect 356 67 357 68 
<< pdiffusion >>
rect 357 67 358 68 
<< pdiffusion >>
rect 358 67 359 68 
<< pdiffusion >>
rect 359 67 360 68 
<< pdiffusion >>
rect 372 67 373 68 
<< pdiffusion >>
rect 373 67 374 68 
<< pdiffusion >>
rect 374 67 375 68 
<< pdiffusion >>
rect 375 67 376 68 
<< pdiffusion >>
rect 376 67 377 68 
<< pdiffusion >>
rect 377 67 378 68 
<< pdiffusion >>
rect 390 67 391 68 
<< pdiffusion >>
rect 391 67 392 68 
<< pdiffusion >>
rect 392 67 393 68 
<< pdiffusion >>
rect 393 67 394 68 
<< pdiffusion >>
rect 394 67 395 68 
<< pdiffusion >>
rect 395 67 396 68 
<< pdiffusion >>
rect 408 67 409 68 
<< pdiffusion >>
rect 409 67 410 68 
<< pdiffusion >>
rect 410 67 411 68 
<< pdiffusion >>
rect 411 67 412 68 
<< pdiffusion >>
rect 412 67 413 68 
<< pdiffusion >>
rect 413 67 414 68 
<< pdiffusion >>
rect 426 67 427 68 
<< pdiffusion >>
rect 427 67 428 68 
<< pdiffusion >>
rect 428 67 429 68 
<< pdiffusion >>
rect 429 67 430 68 
<< pdiffusion >>
rect 430 67 431 68 
<< pdiffusion >>
rect 431 67 432 68 
<< pdiffusion >>
rect 444 67 445 68 
<< pdiffusion >>
rect 445 67 446 68 
<< pdiffusion >>
rect 446 67 447 68 
<< pdiffusion >>
rect 447 67 448 68 
<< pdiffusion >>
rect 448 67 449 68 
<< pdiffusion >>
rect 449 67 450 68 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 64 68 65 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< m1 >>
rect 91 68 92 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< pdiffusion >>
rect 138 68 139 69 
<< pdiffusion >>
rect 139 68 140 69 
<< pdiffusion >>
rect 140 68 141 69 
<< pdiffusion >>
rect 141 68 142 69 
<< pdiffusion >>
rect 142 68 143 69 
<< pdiffusion >>
rect 143 68 144 69 
<< m1 >>
rect 145 68 146 69 
<< m1 >>
rect 154 68 155 69 
<< pdiffusion >>
rect 156 68 157 69 
<< pdiffusion >>
rect 157 68 158 69 
<< pdiffusion >>
rect 158 68 159 69 
<< pdiffusion >>
rect 159 68 160 69 
<< pdiffusion >>
rect 160 68 161 69 
<< pdiffusion >>
rect 161 68 162 69 
<< pdiffusion >>
rect 174 68 175 69 
<< pdiffusion >>
rect 175 68 176 69 
<< pdiffusion >>
rect 176 68 177 69 
<< pdiffusion >>
rect 177 68 178 69 
<< pdiffusion >>
rect 178 68 179 69 
<< pdiffusion >>
rect 179 68 180 69 
<< m1 >>
rect 181 68 182 69 
<< pdiffusion >>
rect 192 68 193 69 
<< pdiffusion >>
rect 193 68 194 69 
<< pdiffusion >>
rect 194 68 195 69 
<< pdiffusion >>
rect 195 68 196 69 
<< pdiffusion >>
rect 196 68 197 69 
<< pdiffusion >>
rect 197 68 198 69 
<< m1 >>
rect 203 68 204 69 
<< m1 >>
rect 208 68 209 69 
<< pdiffusion >>
rect 210 68 211 69 
<< pdiffusion >>
rect 211 68 212 69 
<< pdiffusion >>
rect 212 68 213 69 
<< pdiffusion >>
rect 213 68 214 69 
<< pdiffusion >>
rect 214 68 215 69 
<< pdiffusion >>
rect 215 68 216 69 
<< m1 >>
rect 217 68 218 69 
<< m1 >>
rect 221 68 222 69 
<< pdiffusion >>
rect 228 68 229 69 
<< pdiffusion >>
rect 229 68 230 69 
<< pdiffusion >>
rect 230 68 231 69 
<< pdiffusion >>
rect 231 68 232 69 
<< pdiffusion >>
rect 232 68 233 69 
<< pdiffusion >>
rect 233 68 234 69 
<< pdiffusion >>
rect 246 68 247 69 
<< pdiffusion >>
rect 247 68 248 69 
<< pdiffusion >>
rect 248 68 249 69 
<< pdiffusion >>
rect 249 68 250 69 
<< pdiffusion >>
rect 250 68 251 69 
<< pdiffusion >>
rect 251 68 252 69 
<< m1 >>
rect 260 68 261 69 
<< m1 >>
rect 262 68 263 69 
<< pdiffusion >>
rect 264 68 265 69 
<< pdiffusion >>
rect 265 68 266 69 
<< pdiffusion >>
rect 266 68 267 69 
<< pdiffusion >>
rect 267 68 268 69 
<< pdiffusion >>
rect 268 68 269 69 
<< pdiffusion >>
rect 269 68 270 69 
<< pdiffusion >>
rect 282 68 283 69 
<< pdiffusion >>
rect 283 68 284 69 
<< pdiffusion >>
rect 284 68 285 69 
<< pdiffusion >>
rect 285 68 286 69 
<< pdiffusion >>
rect 286 68 287 69 
<< pdiffusion >>
rect 287 68 288 69 
<< pdiffusion >>
rect 300 68 301 69 
<< pdiffusion >>
rect 301 68 302 69 
<< pdiffusion >>
rect 302 68 303 69 
<< pdiffusion >>
rect 303 68 304 69 
<< pdiffusion >>
rect 304 68 305 69 
<< pdiffusion >>
rect 305 68 306 69 
<< pdiffusion >>
rect 336 68 337 69 
<< pdiffusion >>
rect 337 68 338 69 
<< pdiffusion >>
rect 338 68 339 69 
<< pdiffusion >>
rect 339 68 340 69 
<< pdiffusion >>
rect 340 68 341 69 
<< pdiffusion >>
rect 341 68 342 69 
<< pdiffusion >>
rect 354 68 355 69 
<< pdiffusion >>
rect 355 68 356 69 
<< pdiffusion >>
rect 356 68 357 69 
<< pdiffusion >>
rect 357 68 358 69 
<< pdiffusion >>
rect 358 68 359 69 
<< pdiffusion >>
rect 359 68 360 69 
<< pdiffusion >>
rect 372 68 373 69 
<< pdiffusion >>
rect 373 68 374 69 
<< pdiffusion >>
rect 374 68 375 69 
<< pdiffusion >>
rect 375 68 376 69 
<< pdiffusion >>
rect 376 68 377 69 
<< pdiffusion >>
rect 377 68 378 69 
<< pdiffusion >>
rect 390 68 391 69 
<< pdiffusion >>
rect 391 68 392 69 
<< pdiffusion >>
rect 392 68 393 69 
<< pdiffusion >>
rect 393 68 394 69 
<< pdiffusion >>
rect 394 68 395 69 
<< pdiffusion >>
rect 395 68 396 69 
<< pdiffusion >>
rect 408 68 409 69 
<< pdiffusion >>
rect 409 68 410 69 
<< pdiffusion >>
rect 410 68 411 69 
<< pdiffusion >>
rect 411 68 412 69 
<< pdiffusion >>
rect 412 68 413 69 
<< pdiffusion >>
rect 413 68 414 69 
<< pdiffusion >>
rect 426 68 427 69 
<< pdiffusion >>
rect 427 68 428 69 
<< pdiffusion >>
rect 428 68 429 69 
<< pdiffusion >>
rect 429 68 430 69 
<< pdiffusion >>
rect 430 68 431 69 
<< pdiffusion >>
rect 431 68 432 69 
<< pdiffusion >>
rect 444 68 445 69 
<< pdiffusion >>
rect 445 68 446 69 
<< pdiffusion >>
rect 446 68 447 69 
<< pdiffusion >>
rect 447 68 448 69 
<< pdiffusion >>
rect 448 68 449 69 
<< pdiffusion >>
rect 449 68 450 69 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 64 69 65 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< m1 >>
rect 91 69 92 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< pdiffusion >>
rect 138 69 139 70 
<< pdiffusion >>
rect 139 69 140 70 
<< pdiffusion >>
rect 140 69 141 70 
<< pdiffusion >>
rect 141 69 142 70 
<< pdiffusion >>
rect 142 69 143 70 
<< pdiffusion >>
rect 143 69 144 70 
<< m1 >>
rect 145 69 146 70 
<< m1 >>
rect 154 69 155 70 
<< pdiffusion >>
rect 156 69 157 70 
<< pdiffusion >>
rect 157 69 158 70 
<< pdiffusion >>
rect 158 69 159 70 
<< pdiffusion >>
rect 159 69 160 70 
<< pdiffusion >>
rect 160 69 161 70 
<< pdiffusion >>
rect 161 69 162 70 
<< pdiffusion >>
rect 174 69 175 70 
<< pdiffusion >>
rect 175 69 176 70 
<< pdiffusion >>
rect 176 69 177 70 
<< pdiffusion >>
rect 177 69 178 70 
<< pdiffusion >>
rect 178 69 179 70 
<< pdiffusion >>
rect 179 69 180 70 
<< m1 >>
rect 181 69 182 70 
<< pdiffusion >>
rect 192 69 193 70 
<< pdiffusion >>
rect 193 69 194 70 
<< pdiffusion >>
rect 194 69 195 70 
<< pdiffusion >>
rect 195 69 196 70 
<< pdiffusion >>
rect 196 69 197 70 
<< pdiffusion >>
rect 197 69 198 70 
<< m1 >>
rect 203 69 204 70 
<< m1 >>
rect 208 69 209 70 
<< pdiffusion >>
rect 210 69 211 70 
<< pdiffusion >>
rect 211 69 212 70 
<< pdiffusion >>
rect 212 69 213 70 
<< pdiffusion >>
rect 213 69 214 70 
<< pdiffusion >>
rect 214 69 215 70 
<< pdiffusion >>
rect 215 69 216 70 
<< m1 >>
rect 217 69 218 70 
<< m1 >>
rect 221 69 222 70 
<< pdiffusion >>
rect 228 69 229 70 
<< pdiffusion >>
rect 229 69 230 70 
<< pdiffusion >>
rect 230 69 231 70 
<< pdiffusion >>
rect 231 69 232 70 
<< pdiffusion >>
rect 232 69 233 70 
<< pdiffusion >>
rect 233 69 234 70 
<< pdiffusion >>
rect 246 69 247 70 
<< pdiffusion >>
rect 247 69 248 70 
<< pdiffusion >>
rect 248 69 249 70 
<< pdiffusion >>
rect 249 69 250 70 
<< pdiffusion >>
rect 250 69 251 70 
<< pdiffusion >>
rect 251 69 252 70 
<< m1 >>
rect 260 69 261 70 
<< m1 >>
rect 262 69 263 70 
<< pdiffusion >>
rect 264 69 265 70 
<< pdiffusion >>
rect 265 69 266 70 
<< pdiffusion >>
rect 266 69 267 70 
<< pdiffusion >>
rect 267 69 268 70 
<< pdiffusion >>
rect 268 69 269 70 
<< pdiffusion >>
rect 269 69 270 70 
<< pdiffusion >>
rect 282 69 283 70 
<< pdiffusion >>
rect 283 69 284 70 
<< pdiffusion >>
rect 284 69 285 70 
<< pdiffusion >>
rect 285 69 286 70 
<< pdiffusion >>
rect 286 69 287 70 
<< pdiffusion >>
rect 287 69 288 70 
<< pdiffusion >>
rect 300 69 301 70 
<< pdiffusion >>
rect 301 69 302 70 
<< pdiffusion >>
rect 302 69 303 70 
<< pdiffusion >>
rect 303 69 304 70 
<< pdiffusion >>
rect 304 69 305 70 
<< pdiffusion >>
rect 305 69 306 70 
<< pdiffusion >>
rect 336 69 337 70 
<< pdiffusion >>
rect 337 69 338 70 
<< pdiffusion >>
rect 338 69 339 70 
<< pdiffusion >>
rect 339 69 340 70 
<< pdiffusion >>
rect 340 69 341 70 
<< pdiffusion >>
rect 341 69 342 70 
<< pdiffusion >>
rect 354 69 355 70 
<< pdiffusion >>
rect 355 69 356 70 
<< pdiffusion >>
rect 356 69 357 70 
<< pdiffusion >>
rect 357 69 358 70 
<< pdiffusion >>
rect 358 69 359 70 
<< pdiffusion >>
rect 359 69 360 70 
<< pdiffusion >>
rect 372 69 373 70 
<< pdiffusion >>
rect 373 69 374 70 
<< pdiffusion >>
rect 374 69 375 70 
<< pdiffusion >>
rect 375 69 376 70 
<< pdiffusion >>
rect 376 69 377 70 
<< pdiffusion >>
rect 377 69 378 70 
<< pdiffusion >>
rect 390 69 391 70 
<< pdiffusion >>
rect 391 69 392 70 
<< pdiffusion >>
rect 392 69 393 70 
<< pdiffusion >>
rect 393 69 394 70 
<< pdiffusion >>
rect 394 69 395 70 
<< pdiffusion >>
rect 395 69 396 70 
<< pdiffusion >>
rect 408 69 409 70 
<< pdiffusion >>
rect 409 69 410 70 
<< pdiffusion >>
rect 410 69 411 70 
<< pdiffusion >>
rect 411 69 412 70 
<< pdiffusion >>
rect 412 69 413 70 
<< pdiffusion >>
rect 413 69 414 70 
<< pdiffusion >>
rect 426 69 427 70 
<< pdiffusion >>
rect 427 69 428 70 
<< pdiffusion >>
rect 428 69 429 70 
<< pdiffusion >>
rect 429 69 430 70 
<< pdiffusion >>
rect 430 69 431 70 
<< pdiffusion >>
rect 431 69 432 70 
<< pdiffusion >>
rect 444 69 445 70 
<< pdiffusion >>
rect 445 69 446 70 
<< pdiffusion >>
rect 446 69 447 70 
<< pdiffusion >>
rect 447 69 448 70 
<< pdiffusion >>
rect 448 69 449 70 
<< pdiffusion >>
rect 449 69 450 70 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 64 70 65 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< m1 >>
rect 91 70 92 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< pdiffusion >>
rect 138 70 139 71 
<< pdiffusion >>
rect 139 70 140 71 
<< pdiffusion >>
rect 140 70 141 71 
<< pdiffusion >>
rect 141 70 142 71 
<< pdiffusion >>
rect 142 70 143 71 
<< pdiffusion >>
rect 143 70 144 71 
<< m1 >>
rect 145 70 146 71 
<< m1 >>
rect 154 70 155 71 
<< pdiffusion >>
rect 156 70 157 71 
<< pdiffusion >>
rect 157 70 158 71 
<< pdiffusion >>
rect 158 70 159 71 
<< pdiffusion >>
rect 159 70 160 71 
<< pdiffusion >>
rect 160 70 161 71 
<< pdiffusion >>
rect 161 70 162 71 
<< pdiffusion >>
rect 174 70 175 71 
<< pdiffusion >>
rect 175 70 176 71 
<< pdiffusion >>
rect 176 70 177 71 
<< pdiffusion >>
rect 177 70 178 71 
<< pdiffusion >>
rect 178 70 179 71 
<< pdiffusion >>
rect 179 70 180 71 
<< m1 >>
rect 181 70 182 71 
<< pdiffusion >>
rect 192 70 193 71 
<< pdiffusion >>
rect 193 70 194 71 
<< pdiffusion >>
rect 194 70 195 71 
<< pdiffusion >>
rect 195 70 196 71 
<< pdiffusion >>
rect 196 70 197 71 
<< pdiffusion >>
rect 197 70 198 71 
<< m1 >>
rect 203 70 204 71 
<< m2 >>
rect 203 70 204 71 
<< m2c >>
rect 203 70 204 71 
<< m1 >>
rect 203 70 204 71 
<< m2 >>
rect 203 70 204 71 
<< m1 >>
rect 208 70 209 71 
<< pdiffusion >>
rect 210 70 211 71 
<< pdiffusion >>
rect 211 70 212 71 
<< pdiffusion >>
rect 212 70 213 71 
<< pdiffusion >>
rect 213 70 214 71 
<< pdiffusion >>
rect 214 70 215 71 
<< pdiffusion >>
rect 215 70 216 71 
<< m1 >>
rect 217 70 218 71 
<< m1 >>
rect 221 70 222 71 
<< pdiffusion >>
rect 228 70 229 71 
<< pdiffusion >>
rect 229 70 230 71 
<< pdiffusion >>
rect 230 70 231 71 
<< pdiffusion >>
rect 231 70 232 71 
<< pdiffusion >>
rect 232 70 233 71 
<< pdiffusion >>
rect 233 70 234 71 
<< pdiffusion >>
rect 246 70 247 71 
<< pdiffusion >>
rect 247 70 248 71 
<< pdiffusion >>
rect 248 70 249 71 
<< pdiffusion >>
rect 249 70 250 71 
<< pdiffusion >>
rect 250 70 251 71 
<< pdiffusion >>
rect 251 70 252 71 
<< m1 >>
rect 260 70 261 71 
<< m1 >>
rect 262 70 263 71 
<< pdiffusion >>
rect 264 70 265 71 
<< pdiffusion >>
rect 265 70 266 71 
<< pdiffusion >>
rect 266 70 267 71 
<< pdiffusion >>
rect 267 70 268 71 
<< pdiffusion >>
rect 268 70 269 71 
<< pdiffusion >>
rect 269 70 270 71 
<< pdiffusion >>
rect 282 70 283 71 
<< pdiffusion >>
rect 283 70 284 71 
<< pdiffusion >>
rect 284 70 285 71 
<< pdiffusion >>
rect 285 70 286 71 
<< pdiffusion >>
rect 286 70 287 71 
<< pdiffusion >>
rect 287 70 288 71 
<< pdiffusion >>
rect 300 70 301 71 
<< pdiffusion >>
rect 301 70 302 71 
<< pdiffusion >>
rect 302 70 303 71 
<< pdiffusion >>
rect 303 70 304 71 
<< pdiffusion >>
rect 304 70 305 71 
<< pdiffusion >>
rect 305 70 306 71 
<< pdiffusion >>
rect 336 70 337 71 
<< pdiffusion >>
rect 337 70 338 71 
<< pdiffusion >>
rect 338 70 339 71 
<< pdiffusion >>
rect 339 70 340 71 
<< pdiffusion >>
rect 340 70 341 71 
<< pdiffusion >>
rect 341 70 342 71 
<< pdiffusion >>
rect 354 70 355 71 
<< pdiffusion >>
rect 355 70 356 71 
<< pdiffusion >>
rect 356 70 357 71 
<< pdiffusion >>
rect 357 70 358 71 
<< pdiffusion >>
rect 358 70 359 71 
<< pdiffusion >>
rect 359 70 360 71 
<< pdiffusion >>
rect 372 70 373 71 
<< pdiffusion >>
rect 373 70 374 71 
<< pdiffusion >>
rect 374 70 375 71 
<< pdiffusion >>
rect 375 70 376 71 
<< pdiffusion >>
rect 376 70 377 71 
<< pdiffusion >>
rect 377 70 378 71 
<< pdiffusion >>
rect 390 70 391 71 
<< pdiffusion >>
rect 391 70 392 71 
<< pdiffusion >>
rect 392 70 393 71 
<< pdiffusion >>
rect 393 70 394 71 
<< pdiffusion >>
rect 394 70 395 71 
<< pdiffusion >>
rect 395 70 396 71 
<< pdiffusion >>
rect 408 70 409 71 
<< pdiffusion >>
rect 409 70 410 71 
<< pdiffusion >>
rect 410 70 411 71 
<< pdiffusion >>
rect 411 70 412 71 
<< pdiffusion >>
rect 412 70 413 71 
<< pdiffusion >>
rect 413 70 414 71 
<< pdiffusion >>
rect 426 70 427 71 
<< pdiffusion >>
rect 427 70 428 71 
<< pdiffusion >>
rect 428 70 429 71 
<< pdiffusion >>
rect 429 70 430 71 
<< pdiffusion >>
rect 430 70 431 71 
<< pdiffusion >>
rect 431 70 432 71 
<< pdiffusion >>
rect 444 70 445 71 
<< pdiffusion >>
rect 445 70 446 71 
<< pdiffusion >>
rect 446 70 447 71 
<< pdiffusion >>
rect 447 70 448 71 
<< pdiffusion >>
rect 448 70 449 71 
<< pdiffusion >>
rect 449 70 450 71 
<< pdiffusion >>
rect 12 71 13 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< pdiffusion >>
rect 30 71 31 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< pdiffusion >>
rect 48 71 49 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 64 71 65 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< m1 >>
rect 91 71 92 72 
<< pdiffusion >>
rect 102 71 103 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< pdiffusion >>
rect 120 71 121 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< pdiffusion >>
rect 138 71 139 72 
<< m1 >>
rect 139 71 140 72 
<< pdiffusion >>
rect 139 71 140 72 
<< pdiffusion >>
rect 140 71 141 72 
<< pdiffusion >>
rect 141 71 142 72 
<< pdiffusion >>
rect 142 71 143 72 
<< pdiffusion >>
rect 143 71 144 72 
<< m1 >>
rect 145 71 146 72 
<< m1 >>
rect 154 71 155 72 
<< pdiffusion >>
rect 156 71 157 72 
<< pdiffusion >>
rect 157 71 158 72 
<< pdiffusion >>
rect 158 71 159 72 
<< pdiffusion >>
rect 159 71 160 72 
<< pdiffusion >>
rect 160 71 161 72 
<< pdiffusion >>
rect 161 71 162 72 
<< pdiffusion >>
rect 174 71 175 72 
<< pdiffusion >>
rect 175 71 176 72 
<< pdiffusion >>
rect 176 71 177 72 
<< pdiffusion >>
rect 177 71 178 72 
<< pdiffusion >>
rect 178 71 179 72 
<< pdiffusion >>
rect 179 71 180 72 
<< m1 >>
rect 181 71 182 72 
<< pdiffusion >>
rect 192 71 193 72 
<< pdiffusion >>
rect 193 71 194 72 
<< pdiffusion >>
rect 194 71 195 72 
<< pdiffusion >>
rect 195 71 196 72 
<< m1 >>
rect 196 71 197 72 
<< pdiffusion >>
rect 196 71 197 72 
<< pdiffusion >>
rect 197 71 198 72 
<< m2 >>
rect 203 71 204 72 
<< m1 >>
rect 208 71 209 72 
<< pdiffusion >>
rect 210 71 211 72 
<< pdiffusion >>
rect 211 71 212 72 
<< pdiffusion >>
rect 212 71 213 72 
<< pdiffusion >>
rect 213 71 214 72 
<< pdiffusion >>
rect 214 71 215 72 
<< pdiffusion >>
rect 215 71 216 72 
<< m1 >>
rect 217 71 218 72 
<< m1 >>
rect 221 71 222 72 
<< pdiffusion >>
rect 228 71 229 72 
<< pdiffusion >>
rect 229 71 230 72 
<< pdiffusion >>
rect 230 71 231 72 
<< pdiffusion >>
rect 231 71 232 72 
<< m1 >>
rect 232 71 233 72 
<< pdiffusion >>
rect 232 71 233 72 
<< pdiffusion >>
rect 233 71 234 72 
<< pdiffusion >>
rect 246 71 247 72 
<< pdiffusion >>
rect 247 71 248 72 
<< pdiffusion >>
rect 248 71 249 72 
<< pdiffusion >>
rect 249 71 250 72 
<< pdiffusion >>
rect 250 71 251 72 
<< pdiffusion >>
rect 251 71 252 72 
<< m1 >>
rect 260 71 261 72 
<< m1 >>
rect 262 71 263 72 
<< pdiffusion >>
rect 264 71 265 72 
<< pdiffusion >>
rect 265 71 266 72 
<< pdiffusion >>
rect 266 71 267 72 
<< pdiffusion >>
rect 267 71 268 72 
<< m1 >>
rect 268 71 269 72 
<< pdiffusion >>
rect 268 71 269 72 
<< pdiffusion >>
rect 269 71 270 72 
<< pdiffusion >>
rect 282 71 283 72 
<< pdiffusion >>
rect 283 71 284 72 
<< pdiffusion >>
rect 284 71 285 72 
<< pdiffusion >>
rect 285 71 286 72 
<< pdiffusion >>
rect 286 71 287 72 
<< pdiffusion >>
rect 287 71 288 72 
<< pdiffusion >>
rect 300 71 301 72 
<< pdiffusion >>
rect 301 71 302 72 
<< pdiffusion >>
rect 302 71 303 72 
<< pdiffusion >>
rect 303 71 304 72 
<< pdiffusion >>
rect 304 71 305 72 
<< pdiffusion >>
rect 305 71 306 72 
<< pdiffusion >>
rect 336 71 337 72 
<< pdiffusion >>
rect 337 71 338 72 
<< pdiffusion >>
rect 338 71 339 72 
<< pdiffusion >>
rect 339 71 340 72 
<< pdiffusion >>
rect 340 71 341 72 
<< pdiffusion >>
rect 341 71 342 72 
<< pdiffusion >>
rect 354 71 355 72 
<< pdiffusion >>
rect 355 71 356 72 
<< pdiffusion >>
rect 356 71 357 72 
<< pdiffusion >>
rect 357 71 358 72 
<< pdiffusion >>
rect 358 71 359 72 
<< pdiffusion >>
rect 359 71 360 72 
<< pdiffusion >>
rect 372 71 373 72 
<< m1 >>
rect 373 71 374 72 
<< pdiffusion >>
rect 373 71 374 72 
<< pdiffusion >>
rect 374 71 375 72 
<< pdiffusion >>
rect 375 71 376 72 
<< pdiffusion >>
rect 376 71 377 72 
<< pdiffusion >>
rect 377 71 378 72 
<< pdiffusion >>
rect 390 71 391 72 
<< m1 >>
rect 391 71 392 72 
<< pdiffusion >>
rect 391 71 392 72 
<< pdiffusion >>
rect 392 71 393 72 
<< pdiffusion >>
rect 393 71 394 72 
<< pdiffusion >>
rect 394 71 395 72 
<< pdiffusion >>
rect 395 71 396 72 
<< pdiffusion >>
rect 408 71 409 72 
<< pdiffusion >>
rect 409 71 410 72 
<< pdiffusion >>
rect 410 71 411 72 
<< pdiffusion >>
rect 411 71 412 72 
<< m1 >>
rect 412 71 413 72 
<< pdiffusion >>
rect 412 71 413 72 
<< pdiffusion >>
rect 413 71 414 72 
<< pdiffusion >>
rect 426 71 427 72 
<< pdiffusion >>
rect 427 71 428 72 
<< pdiffusion >>
rect 428 71 429 72 
<< pdiffusion >>
rect 429 71 430 72 
<< pdiffusion >>
rect 430 71 431 72 
<< pdiffusion >>
rect 431 71 432 72 
<< pdiffusion >>
rect 444 71 445 72 
<< pdiffusion >>
rect 445 71 446 72 
<< pdiffusion >>
rect 446 71 447 72 
<< pdiffusion >>
rect 447 71 448 72 
<< pdiffusion >>
rect 448 71 449 72 
<< pdiffusion >>
rect 449 71 450 72 
<< m1 >>
rect 64 72 65 73 
<< m1 >>
rect 91 72 92 73 
<< m1 >>
rect 139 72 140 73 
<< m1 >>
rect 145 72 146 73 
<< m1 >>
rect 154 72 155 73 
<< m1 >>
rect 181 72 182 73 
<< m1 >>
rect 196 72 197 73 
<< m2 >>
rect 200 72 201 73 
<< m1 >>
rect 201 72 202 73 
<< m2 >>
rect 201 72 202 73 
<< m2c >>
rect 201 72 202 73 
<< m1 >>
rect 201 72 202 73 
<< m2 >>
rect 201 72 202 73 
<< m1 >>
rect 202 72 203 73 
<< m1 >>
rect 203 72 204 73 
<< m2 >>
rect 203 72 204 73 
<< m1 >>
rect 204 72 205 73 
<< m1 >>
rect 205 72 206 73 
<< m1 >>
rect 206 72 207 73 
<< m1 >>
rect 207 72 208 73 
<< m1 >>
rect 208 72 209 73 
<< m1 >>
rect 217 72 218 73 
<< m1 >>
rect 221 72 222 73 
<< m1 >>
rect 232 72 233 73 
<< m1 >>
rect 260 72 261 73 
<< m1 >>
rect 262 72 263 73 
<< m1 >>
rect 268 72 269 73 
<< m1 >>
rect 373 72 374 73 
<< m1 >>
rect 391 72 392 73 
<< m1 >>
rect 412 72 413 73 
<< m1 >>
rect 64 73 65 74 
<< m1 >>
rect 91 73 92 74 
<< m1 >>
rect 139 73 140 74 
<< m1 >>
rect 145 73 146 74 
<< m1 >>
rect 154 73 155 74 
<< m1 >>
rect 181 73 182 74 
<< m1 >>
rect 196 73 197 74 
<< m1 >>
rect 197 73 198 74 
<< m1 >>
rect 198 73 199 74 
<< m1 >>
rect 199 73 200 74 
<< m2 >>
rect 200 73 201 74 
<< m2 >>
rect 203 73 204 74 
<< m1 >>
rect 217 73 218 74 
<< m1 >>
rect 221 73 222 74 
<< m1 >>
rect 232 73 233 74 
<< m1 >>
rect 260 73 261 74 
<< m1 >>
rect 262 73 263 74 
<< m1 >>
rect 268 73 269 74 
<< m1 >>
rect 373 73 374 74 
<< m1 >>
rect 391 73 392 74 
<< m1 >>
rect 412 73 413 74 
<< m1 >>
rect 64 74 65 75 
<< m1 >>
rect 91 74 92 75 
<< m1 >>
rect 139 74 140 75 
<< m1 >>
rect 140 74 141 75 
<< m1 >>
rect 141 74 142 75 
<< m1 >>
rect 142 74 143 75 
<< m1 >>
rect 143 74 144 75 
<< m1 >>
rect 144 74 145 75 
<< m1 >>
rect 145 74 146 75 
<< m1 >>
rect 154 74 155 75 
<< m1 >>
rect 181 74 182 75 
<< m1 >>
rect 199 74 200 75 
<< m2 >>
rect 200 74 201 75 
<< m1 >>
rect 203 74 204 75 
<< m2 >>
rect 203 74 204 75 
<< m2c >>
rect 203 74 204 75 
<< m1 >>
rect 203 74 204 75 
<< m2 >>
rect 203 74 204 75 
<< m1 >>
rect 217 74 218 75 
<< m1 >>
rect 221 74 222 75 
<< m2 >>
rect 221 74 222 75 
<< m2c >>
rect 221 74 222 75 
<< m1 >>
rect 221 74 222 75 
<< m2 >>
rect 221 74 222 75 
<< m1 >>
rect 232 74 233 75 
<< m1 >>
rect 233 74 234 75 
<< m1 >>
rect 234 74 235 75 
<< m1 >>
rect 235 74 236 75 
<< m1 >>
rect 236 74 237 75 
<< m1 >>
rect 237 74 238 75 
<< m1 >>
rect 238 74 239 75 
<< m1 >>
rect 239 74 240 75 
<< m1 >>
rect 240 74 241 75 
<< m1 >>
rect 241 74 242 75 
<< m1 >>
rect 242 74 243 75 
<< m1 >>
rect 243 74 244 75 
<< m1 >>
rect 244 74 245 75 
<< m1 >>
rect 245 74 246 75 
<< m1 >>
rect 246 74 247 75 
<< m2 >>
rect 246 74 247 75 
<< m2c >>
rect 246 74 247 75 
<< m1 >>
rect 246 74 247 75 
<< m2 >>
rect 246 74 247 75 
<< m1 >>
rect 260 74 261 75 
<< m1 >>
rect 262 74 263 75 
<< m1 >>
rect 268 74 269 75 
<< m1 >>
rect 373 74 374 75 
<< m1 >>
rect 391 74 392 75 
<< m1 >>
rect 412 74 413 75 
<< m1 >>
rect 413 74 414 75 
<< m1 >>
rect 414 74 415 75 
<< m1 >>
rect 415 74 416 75 
<< m1 >>
rect 416 74 417 75 
<< m1 >>
rect 417 74 418 75 
<< m1 >>
rect 418 74 419 75 
<< m1 >>
rect 419 74 420 75 
<< m1 >>
rect 420 74 421 75 
<< m1 >>
rect 421 74 422 75 
<< m1 >>
rect 422 74 423 75 
<< m1 >>
rect 423 74 424 75 
<< m1 >>
rect 424 74 425 75 
<< m1 >>
rect 64 75 65 76 
<< m1 >>
rect 91 75 92 76 
<< m1 >>
rect 154 75 155 76 
<< m1 >>
rect 181 75 182 76 
<< m1 >>
rect 197 75 198 76 
<< m2 >>
rect 197 75 198 76 
<< m2c >>
rect 197 75 198 76 
<< m1 >>
rect 197 75 198 76 
<< m2 >>
rect 197 75 198 76 
<< m2 >>
rect 198 75 199 76 
<< m1 >>
rect 199 75 200 76 
<< m2 >>
rect 199 75 200 76 
<< m2 >>
rect 200 75 201 76 
<< m1 >>
rect 203 75 204 76 
<< m1 >>
rect 217 75 218 76 
<< m2 >>
rect 221 75 222 76 
<< m2 >>
rect 246 75 247 76 
<< m1 >>
rect 260 75 261 76 
<< m1 >>
rect 262 75 263 76 
<< m1 >>
rect 268 75 269 76 
<< m1 >>
rect 373 75 374 76 
<< m1 >>
rect 391 75 392 76 
<< m1 >>
rect 424 75 425 76 
<< m1 >>
rect 64 76 65 77 
<< m1 >>
rect 91 76 92 77 
<< m1 >>
rect 154 76 155 77 
<< m1 >>
rect 181 76 182 77 
<< m1 >>
rect 193 76 194 77 
<< m1 >>
rect 194 76 195 77 
<< m1 >>
rect 195 76 196 77 
<< m1 >>
rect 196 76 197 77 
<< m1 >>
rect 197 76 198 77 
<< m1 >>
rect 199 76 200 77 
<< m1 >>
rect 203 76 204 77 
<< m1 >>
rect 204 76 205 77 
<< m1 >>
rect 205 76 206 77 
<< m1 >>
rect 206 76 207 77 
<< m1 >>
rect 207 76 208 77 
<< m1 >>
rect 208 76 209 77 
<< m1 >>
rect 209 76 210 77 
<< m1 >>
rect 210 76 211 77 
<< m1 >>
rect 211 76 212 77 
<< m1 >>
rect 212 76 213 77 
<< m1 >>
rect 213 76 214 77 
<< m1 >>
rect 214 76 215 77 
<< m1 >>
rect 215 76 216 77 
<< m2 >>
rect 215 76 216 77 
<< m2c >>
rect 215 76 216 77 
<< m1 >>
rect 215 76 216 77 
<< m2 >>
rect 215 76 216 77 
<< m2 >>
rect 216 76 217 77 
<< m1 >>
rect 217 76 218 77 
<< m2 >>
rect 217 76 218 77 
<< m2 >>
rect 218 76 219 77 
<< m1 >>
rect 219 76 220 77 
<< m2 >>
rect 219 76 220 77 
<< m2c >>
rect 219 76 220 77 
<< m1 >>
rect 219 76 220 77 
<< m2 >>
rect 219 76 220 77 
<< m1 >>
rect 220 76 221 77 
<< m1 >>
rect 221 76 222 77 
<< m2 >>
rect 221 76 222 77 
<< m1 >>
rect 222 76 223 77 
<< m1 >>
rect 223 76 224 77 
<< m1 >>
rect 224 76 225 77 
<< m1 >>
rect 225 76 226 77 
<< m1 >>
rect 226 76 227 77 
<< m1 >>
rect 227 76 228 77 
<< m1 >>
rect 228 76 229 77 
<< m1 >>
rect 229 76 230 77 
<< m1 >>
rect 230 76 231 77 
<< m1 >>
rect 231 76 232 77 
<< m1 >>
rect 232 76 233 77 
<< m1 >>
rect 233 76 234 77 
<< m1 >>
rect 234 76 235 77 
<< m1 >>
rect 235 76 236 77 
<< m1 >>
rect 236 76 237 77 
<< m1 >>
rect 237 76 238 77 
<< m1 >>
rect 238 76 239 77 
<< m1 >>
rect 239 76 240 77 
<< m1 >>
rect 240 76 241 77 
<< m1 >>
rect 241 76 242 77 
<< m1 >>
rect 242 76 243 77 
<< m1 >>
rect 243 76 244 77 
<< m1 >>
rect 244 76 245 77 
<< m1 >>
rect 245 76 246 77 
<< m1 >>
rect 246 76 247 77 
<< m2 >>
rect 246 76 247 77 
<< m1 >>
rect 247 76 248 77 
<< m1 >>
rect 248 76 249 77 
<< m1 >>
rect 249 76 250 77 
<< m1 >>
rect 250 76 251 77 
<< m1 >>
rect 251 76 252 77 
<< m1 >>
rect 252 76 253 77 
<< m1 >>
rect 253 76 254 77 
<< m1 >>
rect 254 76 255 77 
<< m1 >>
rect 255 76 256 77 
<< m1 >>
rect 256 76 257 77 
<< m1 >>
rect 257 76 258 77 
<< m1 >>
rect 258 76 259 77 
<< m2 >>
rect 258 76 259 77 
<< m2c >>
rect 258 76 259 77 
<< m1 >>
rect 258 76 259 77 
<< m2 >>
rect 258 76 259 77 
<< m2 >>
rect 259 76 260 77 
<< m1 >>
rect 260 76 261 77 
<< m2 >>
rect 260 76 261 77 
<< m2 >>
rect 261 76 262 77 
<< m1 >>
rect 262 76 263 77 
<< m2 >>
rect 262 76 263 77 
<< m2 >>
rect 263 76 264 77 
<< m1 >>
rect 264 76 265 77 
<< m2 >>
rect 264 76 265 77 
<< m2c >>
rect 264 76 265 77 
<< m1 >>
rect 264 76 265 77 
<< m2 >>
rect 264 76 265 77 
<< m1 >>
rect 265 76 266 77 
<< m1 >>
rect 266 76 267 77 
<< m1 >>
rect 267 76 268 77 
<< m1 >>
rect 268 76 269 77 
<< m1 >>
rect 352 76 353 77 
<< m1 >>
rect 353 76 354 77 
<< m1 >>
rect 354 76 355 77 
<< m1 >>
rect 355 76 356 77 
<< m1 >>
rect 356 76 357 77 
<< m1 >>
rect 357 76 358 77 
<< m1 >>
rect 358 76 359 77 
<< m1 >>
rect 359 76 360 77 
<< m1 >>
rect 360 76 361 77 
<< m1 >>
rect 361 76 362 77 
<< m1 >>
rect 362 76 363 77 
<< m1 >>
rect 363 76 364 77 
<< m1 >>
rect 364 76 365 77 
<< m1 >>
rect 365 76 366 77 
<< m1 >>
rect 366 76 367 77 
<< m1 >>
rect 367 76 368 77 
<< m1 >>
rect 368 76 369 77 
<< m1 >>
rect 369 76 370 77 
<< m1 >>
rect 370 76 371 77 
<< m1 >>
rect 371 76 372 77 
<< m1 >>
rect 372 76 373 77 
<< m1 >>
rect 373 76 374 77 
<< m1 >>
rect 391 76 392 77 
<< m1 >>
rect 392 76 393 77 
<< m1 >>
rect 393 76 394 77 
<< m1 >>
rect 394 76 395 77 
<< m1 >>
rect 395 76 396 77 
<< m1 >>
rect 396 76 397 77 
<< m1 >>
rect 397 76 398 77 
<< m1 >>
rect 398 76 399 77 
<< m1 >>
rect 399 76 400 77 
<< m1 >>
rect 400 76 401 77 
<< m1 >>
rect 401 76 402 77 
<< m1 >>
rect 402 76 403 77 
<< m1 >>
rect 403 76 404 77 
<< m1 >>
rect 404 76 405 77 
<< m1 >>
rect 405 76 406 77 
<< m1 >>
rect 406 76 407 77 
<< m1 >>
rect 407 76 408 77 
<< m1 >>
rect 408 76 409 77 
<< m1 >>
rect 409 76 410 77 
<< m1 >>
rect 410 76 411 77 
<< m1 >>
rect 411 76 412 77 
<< m1 >>
rect 412 76 413 77 
<< m1 >>
rect 424 76 425 77 
<< m1 >>
rect 64 77 65 78 
<< m1 >>
rect 91 77 92 78 
<< m1 >>
rect 154 77 155 78 
<< m1 >>
rect 181 77 182 78 
<< m1 >>
rect 193 77 194 78 
<< m1 >>
rect 199 77 200 78 
<< m1 >>
rect 217 77 218 78 
<< m2 >>
rect 221 77 222 78 
<< m2 >>
rect 246 77 247 78 
<< m2 >>
rect 247 77 248 78 
<< m2 >>
rect 248 77 249 78 
<< m2 >>
rect 249 77 250 78 
<< m2 >>
rect 250 77 251 78 
<< m2 >>
rect 251 77 252 78 
<< m2 >>
rect 252 77 253 78 
<< m2 >>
rect 253 77 254 78 
<< m1 >>
rect 260 77 261 78 
<< m1 >>
rect 262 77 263 78 
<< m1 >>
rect 352 77 353 78 
<< m1 >>
rect 412 77 413 78 
<< m1 >>
rect 424 77 425 78 
<< m1 >>
rect 64 78 65 79 
<< m1 >>
rect 91 78 92 79 
<< m1 >>
rect 154 78 155 79 
<< m1 >>
rect 181 78 182 79 
<< m1 >>
rect 193 78 194 79 
<< m1 >>
rect 199 78 200 79 
<< m1 >>
rect 217 78 218 79 
<< m1 >>
rect 221 78 222 79 
<< m2 >>
rect 221 78 222 79 
<< m2c >>
rect 221 78 222 79 
<< m1 >>
rect 221 78 222 79 
<< m2 >>
rect 221 78 222 79 
<< m1 >>
rect 253 78 254 79 
<< m2 >>
rect 253 78 254 79 
<< m2c >>
rect 253 78 254 79 
<< m1 >>
rect 253 78 254 79 
<< m2 >>
rect 253 78 254 79 
<< m1 >>
rect 260 78 261 79 
<< m1 >>
rect 262 78 263 79 
<< m1 >>
rect 352 78 353 79 
<< m1 >>
rect 412 78 413 79 
<< m1 >>
rect 424 78 425 79 
<< m1 >>
rect 64 79 65 80 
<< m1 >>
rect 91 79 92 80 
<< m1 >>
rect 154 79 155 80 
<< m1 >>
rect 155 79 156 80 
<< m1 >>
rect 156 79 157 80 
<< m1 >>
rect 157 79 158 80 
<< m1 >>
rect 158 79 159 80 
<< m1 >>
rect 159 79 160 80 
<< m1 >>
rect 160 79 161 80 
<< m1 >>
rect 181 79 182 80 
<< m1 >>
rect 190 79 191 80 
<< m1 >>
rect 191 79 192 80 
<< m2 >>
rect 191 79 192 80 
<< m2c >>
rect 191 79 192 80 
<< m1 >>
rect 191 79 192 80 
<< m2 >>
rect 191 79 192 80 
<< m2 >>
rect 192 79 193 80 
<< m1 >>
rect 193 79 194 80 
<< m2 >>
rect 193 79 194 80 
<< m2 >>
rect 194 79 195 80 
<< m1 >>
rect 199 79 200 80 
<< m1 >>
rect 217 79 218 80 
<< m1 >>
rect 221 79 222 80 
<< m1 >>
rect 253 79 254 80 
<< m1 >>
rect 260 79 261 80 
<< m1 >>
rect 262 79 263 80 
<< m1 >>
rect 298 79 299 80 
<< m1 >>
rect 299 79 300 80 
<< m1 >>
rect 300 79 301 80 
<< m1 >>
rect 301 79 302 80 
<< m1 >>
rect 302 79 303 80 
<< m1 >>
rect 303 79 304 80 
<< m1 >>
rect 304 79 305 80 
<< m1 >>
rect 352 79 353 80 
<< m1 >>
rect 412 79 413 80 
<< m1 >>
rect 424 79 425 80 
<< m1 >>
rect 64 80 65 81 
<< m1 >>
rect 91 80 92 81 
<< m1 >>
rect 160 80 161 81 
<< m1 >>
rect 181 80 182 81 
<< m1 >>
rect 190 80 191 81 
<< m1 >>
rect 193 80 194 81 
<< m2 >>
rect 194 80 195 81 
<< m1 >>
rect 199 80 200 81 
<< m1 >>
rect 217 80 218 81 
<< m1 >>
rect 221 80 222 81 
<< m1 >>
rect 253 80 254 81 
<< m1 >>
rect 260 80 261 81 
<< m1 >>
rect 262 80 263 81 
<< m1 >>
rect 298 80 299 81 
<< m1 >>
rect 304 80 305 81 
<< m1 >>
rect 352 80 353 81 
<< m1 >>
rect 412 80 413 81 
<< m1 >>
rect 424 80 425 81 
<< m1 >>
rect 64 81 65 82 
<< m1 >>
rect 91 81 92 82 
<< m1 >>
rect 160 81 161 82 
<< m1 >>
rect 175 81 176 82 
<< m1 >>
rect 176 81 177 82 
<< m1 >>
rect 177 81 178 82 
<< m1 >>
rect 178 81 179 82 
<< m1 >>
rect 179 81 180 82 
<< m1 >>
rect 180 81 181 82 
<< m1 >>
rect 181 81 182 82 
<< m1 >>
rect 190 81 191 82 
<< m1 >>
rect 193 81 194 82 
<< m2 >>
rect 194 81 195 82 
<< m1 >>
rect 199 81 200 82 
<< m1 >>
rect 217 81 218 82 
<< m1 >>
rect 221 81 222 82 
<< m1 >>
rect 253 81 254 82 
<< m1 >>
rect 260 81 261 82 
<< m1 >>
rect 262 81 263 82 
<< m1 >>
rect 298 81 299 82 
<< m1 >>
rect 304 81 305 82 
<< m1 >>
rect 352 81 353 82 
<< m1 >>
rect 412 81 413 82 
<< m1 >>
rect 424 81 425 82 
<< m1 >>
rect 64 82 65 83 
<< m1 >>
rect 65 82 66 83 
<< m1 >>
rect 66 82 67 83 
<< m1 >>
rect 67 82 68 83 
<< m1 >>
rect 91 82 92 83 
<< m1 >>
rect 160 82 161 83 
<< m1 >>
rect 175 82 176 83 
<< m1 >>
rect 190 82 191 83 
<< m1 >>
rect 193 82 194 83 
<< m2 >>
rect 194 82 195 83 
<< m1 >>
rect 195 82 196 83 
<< m2 >>
rect 195 82 196 83 
<< m2c >>
rect 195 82 196 83 
<< m1 >>
rect 195 82 196 83 
<< m2 >>
rect 195 82 196 83 
<< m1 >>
rect 196 82 197 83 
<< m1 >>
rect 199 82 200 83 
<< m1 >>
rect 217 82 218 83 
<< m1 >>
rect 221 82 222 83 
<< m1 >>
rect 253 82 254 83 
<< m1 >>
rect 260 82 261 83 
<< m1 >>
rect 262 82 263 83 
<< m1 >>
rect 298 82 299 83 
<< m1 >>
rect 304 82 305 83 
<< m1 >>
rect 352 82 353 83 
<< m1 >>
rect 376 82 377 83 
<< m1 >>
rect 377 82 378 83 
<< m1 >>
rect 378 82 379 83 
<< m1 >>
rect 379 82 380 83 
<< m1 >>
rect 412 82 413 83 
<< m1 >>
rect 424 82 425 83 
<< m1 >>
rect 448 82 449 83 
<< m1 >>
rect 449 82 450 83 
<< m1 >>
rect 450 82 451 83 
<< m1 >>
rect 451 82 452 83 
<< m1 >>
rect 67 83 68 84 
<< m1 >>
rect 91 83 92 84 
<< m1 >>
rect 160 83 161 84 
<< m1 >>
rect 175 83 176 84 
<< m1 >>
rect 190 83 191 84 
<< m1 >>
rect 193 83 194 84 
<< m1 >>
rect 196 83 197 84 
<< m1 >>
rect 199 83 200 84 
<< m1 >>
rect 217 83 218 84 
<< m1 >>
rect 221 83 222 84 
<< m1 >>
rect 253 83 254 84 
<< m1 >>
rect 260 83 261 84 
<< m1 >>
rect 262 83 263 84 
<< m1 >>
rect 298 83 299 84 
<< m1 >>
rect 304 83 305 84 
<< m1 >>
rect 352 83 353 84 
<< m1 >>
rect 376 83 377 84 
<< m1 >>
rect 379 83 380 84 
<< m1 >>
rect 412 83 413 84 
<< m1 >>
rect 424 83 425 84 
<< m1 >>
rect 448 83 449 84 
<< m1 >>
rect 451 83 452 84 
<< pdiffusion >>
rect 12 84 13 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< pdiffusion >>
rect 30 84 31 85 
<< pdiffusion >>
rect 31 84 32 85 
<< pdiffusion >>
rect 32 84 33 85 
<< pdiffusion >>
rect 33 84 34 85 
<< pdiffusion >>
rect 34 84 35 85 
<< pdiffusion >>
rect 35 84 36 85 
<< pdiffusion >>
rect 48 84 49 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< pdiffusion >>
rect 66 84 67 85 
<< m1 >>
rect 67 84 68 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 91 84 92 85 
<< pdiffusion >>
rect 102 84 103 85 
<< pdiffusion >>
rect 103 84 104 85 
<< pdiffusion >>
rect 104 84 105 85 
<< pdiffusion >>
rect 105 84 106 85 
<< pdiffusion >>
rect 106 84 107 85 
<< pdiffusion >>
rect 107 84 108 85 
<< pdiffusion >>
rect 120 84 121 85 
<< pdiffusion >>
rect 121 84 122 85 
<< pdiffusion >>
rect 122 84 123 85 
<< pdiffusion >>
rect 123 84 124 85 
<< pdiffusion >>
rect 124 84 125 85 
<< pdiffusion >>
rect 125 84 126 85 
<< pdiffusion >>
rect 138 84 139 85 
<< pdiffusion >>
rect 139 84 140 85 
<< pdiffusion >>
rect 140 84 141 85 
<< pdiffusion >>
rect 141 84 142 85 
<< pdiffusion >>
rect 142 84 143 85 
<< pdiffusion >>
rect 143 84 144 85 
<< pdiffusion >>
rect 156 84 157 85 
<< pdiffusion >>
rect 157 84 158 85 
<< pdiffusion >>
rect 158 84 159 85 
<< pdiffusion >>
rect 159 84 160 85 
<< m1 >>
rect 160 84 161 85 
<< pdiffusion >>
rect 160 84 161 85 
<< pdiffusion >>
rect 161 84 162 85 
<< pdiffusion >>
rect 174 84 175 85 
<< m1 >>
rect 175 84 176 85 
<< pdiffusion >>
rect 175 84 176 85 
<< pdiffusion >>
rect 176 84 177 85 
<< pdiffusion >>
rect 177 84 178 85 
<< pdiffusion >>
rect 178 84 179 85 
<< pdiffusion >>
rect 179 84 180 85 
<< m1 >>
rect 190 84 191 85 
<< pdiffusion >>
rect 192 84 193 85 
<< m1 >>
rect 193 84 194 85 
<< pdiffusion >>
rect 193 84 194 85 
<< pdiffusion >>
rect 194 84 195 85 
<< pdiffusion >>
rect 195 84 196 85 
<< m1 >>
rect 196 84 197 85 
<< pdiffusion >>
rect 196 84 197 85 
<< pdiffusion >>
rect 197 84 198 85 
<< m1 >>
rect 199 84 200 85 
<< pdiffusion >>
rect 210 84 211 85 
<< pdiffusion >>
rect 211 84 212 85 
<< pdiffusion >>
rect 212 84 213 85 
<< pdiffusion >>
rect 213 84 214 85 
<< pdiffusion >>
rect 214 84 215 85 
<< pdiffusion >>
rect 215 84 216 85 
<< m1 >>
rect 217 84 218 85 
<< m1 >>
rect 221 84 222 85 
<< pdiffusion >>
rect 228 84 229 85 
<< pdiffusion >>
rect 229 84 230 85 
<< pdiffusion >>
rect 230 84 231 85 
<< pdiffusion >>
rect 231 84 232 85 
<< pdiffusion >>
rect 232 84 233 85 
<< pdiffusion >>
rect 233 84 234 85 
<< pdiffusion >>
rect 246 84 247 85 
<< pdiffusion >>
rect 247 84 248 85 
<< pdiffusion >>
rect 248 84 249 85 
<< pdiffusion >>
rect 249 84 250 85 
<< pdiffusion >>
rect 250 84 251 85 
<< pdiffusion >>
rect 251 84 252 85 
<< m1 >>
rect 253 84 254 85 
<< m1 >>
rect 260 84 261 85 
<< m1 >>
rect 262 84 263 85 
<< pdiffusion >>
rect 264 84 265 85 
<< pdiffusion >>
rect 265 84 266 85 
<< pdiffusion >>
rect 266 84 267 85 
<< pdiffusion >>
rect 267 84 268 85 
<< pdiffusion >>
rect 268 84 269 85 
<< pdiffusion >>
rect 269 84 270 85 
<< pdiffusion >>
rect 282 84 283 85 
<< pdiffusion >>
rect 283 84 284 85 
<< pdiffusion >>
rect 284 84 285 85 
<< pdiffusion >>
rect 285 84 286 85 
<< pdiffusion >>
rect 286 84 287 85 
<< pdiffusion >>
rect 287 84 288 85 
<< m1 >>
rect 298 84 299 85 
<< pdiffusion >>
rect 300 84 301 85 
<< pdiffusion >>
rect 301 84 302 85 
<< pdiffusion >>
rect 302 84 303 85 
<< pdiffusion >>
rect 303 84 304 85 
<< m1 >>
rect 304 84 305 85 
<< pdiffusion >>
rect 304 84 305 85 
<< pdiffusion >>
rect 305 84 306 85 
<< pdiffusion >>
rect 318 84 319 85 
<< pdiffusion >>
rect 319 84 320 85 
<< pdiffusion >>
rect 320 84 321 85 
<< pdiffusion >>
rect 321 84 322 85 
<< pdiffusion >>
rect 322 84 323 85 
<< pdiffusion >>
rect 323 84 324 85 
<< pdiffusion >>
rect 336 84 337 85 
<< pdiffusion >>
rect 337 84 338 85 
<< pdiffusion >>
rect 338 84 339 85 
<< pdiffusion >>
rect 339 84 340 85 
<< pdiffusion >>
rect 340 84 341 85 
<< pdiffusion >>
rect 341 84 342 85 
<< m1 >>
rect 352 84 353 85 
<< pdiffusion >>
rect 354 84 355 85 
<< pdiffusion >>
rect 355 84 356 85 
<< pdiffusion >>
rect 356 84 357 85 
<< pdiffusion >>
rect 357 84 358 85 
<< pdiffusion >>
rect 358 84 359 85 
<< pdiffusion >>
rect 359 84 360 85 
<< pdiffusion >>
rect 372 84 373 85 
<< pdiffusion >>
rect 373 84 374 85 
<< pdiffusion >>
rect 374 84 375 85 
<< pdiffusion >>
rect 375 84 376 85 
<< m1 >>
rect 376 84 377 85 
<< pdiffusion >>
rect 376 84 377 85 
<< pdiffusion >>
rect 377 84 378 85 
<< m1 >>
rect 379 84 380 85 
<< pdiffusion >>
rect 390 84 391 85 
<< pdiffusion >>
rect 391 84 392 85 
<< pdiffusion >>
rect 392 84 393 85 
<< pdiffusion >>
rect 393 84 394 85 
<< pdiffusion >>
rect 394 84 395 85 
<< pdiffusion >>
rect 395 84 396 85 
<< pdiffusion >>
rect 408 84 409 85 
<< pdiffusion >>
rect 409 84 410 85 
<< pdiffusion >>
rect 410 84 411 85 
<< pdiffusion >>
rect 411 84 412 85 
<< m1 >>
rect 412 84 413 85 
<< pdiffusion >>
rect 412 84 413 85 
<< pdiffusion >>
rect 413 84 414 85 
<< m1 >>
rect 424 84 425 85 
<< pdiffusion >>
rect 426 84 427 85 
<< pdiffusion >>
rect 427 84 428 85 
<< pdiffusion >>
rect 428 84 429 85 
<< pdiffusion >>
rect 429 84 430 85 
<< pdiffusion >>
rect 430 84 431 85 
<< pdiffusion >>
rect 431 84 432 85 
<< pdiffusion >>
rect 444 84 445 85 
<< pdiffusion >>
rect 445 84 446 85 
<< pdiffusion >>
rect 446 84 447 85 
<< pdiffusion >>
rect 447 84 448 85 
<< m1 >>
rect 448 84 449 85 
<< pdiffusion >>
rect 448 84 449 85 
<< pdiffusion >>
rect 449 84 450 85 
<< m1 >>
rect 451 84 452 85 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< pdiffusion >>
rect 30 85 31 86 
<< pdiffusion >>
rect 31 85 32 86 
<< pdiffusion >>
rect 32 85 33 86 
<< pdiffusion >>
rect 33 85 34 86 
<< pdiffusion >>
rect 34 85 35 86 
<< pdiffusion >>
rect 35 85 36 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 91 85 92 86 
<< pdiffusion >>
rect 102 85 103 86 
<< pdiffusion >>
rect 103 85 104 86 
<< pdiffusion >>
rect 104 85 105 86 
<< pdiffusion >>
rect 105 85 106 86 
<< pdiffusion >>
rect 106 85 107 86 
<< pdiffusion >>
rect 107 85 108 86 
<< pdiffusion >>
rect 120 85 121 86 
<< pdiffusion >>
rect 121 85 122 86 
<< pdiffusion >>
rect 122 85 123 86 
<< pdiffusion >>
rect 123 85 124 86 
<< pdiffusion >>
rect 124 85 125 86 
<< pdiffusion >>
rect 125 85 126 86 
<< pdiffusion >>
rect 138 85 139 86 
<< pdiffusion >>
rect 139 85 140 86 
<< pdiffusion >>
rect 140 85 141 86 
<< pdiffusion >>
rect 141 85 142 86 
<< pdiffusion >>
rect 142 85 143 86 
<< pdiffusion >>
rect 143 85 144 86 
<< pdiffusion >>
rect 156 85 157 86 
<< pdiffusion >>
rect 157 85 158 86 
<< pdiffusion >>
rect 158 85 159 86 
<< pdiffusion >>
rect 159 85 160 86 
<< pdiffusion >>
rect 160 85 161 86 
<< pdiffusion >>
rect 161 85 162 86 
<< pdiffusion >>
rect 174 85 175 86 
<< pdiffusion >>
rect 175 85 176 86 
<< pdiffusion >>
rect 176 85 177 86 
<< pdiffusion >>
rect 177 85 178 86 
<< pdiffusion >>
rect 178 85 179 86 
<< pdiffusion >>
rect 179 85 180 86 
<< m1 >>
rect 190 85 191 86 
<< pdiffusion >>
rect 192 85 193 86 
<< pdiffusion >>
rect 193 85 194 86 
<< pdiffusion >>
rect 194 85 195 86 
<< pdiffusion >>
rect 195 85 196 86 
<< pdiffusion >>
rect 196 85 197 86 
<< pdiffusion >>
rect 197 85 198 86 
<< m1 >>
rect 199 85 200 86 
<< pdiffusion >>
rect 210 85 211 86 
<< pdiffusion >>
rect 211 85 212 86 
<< pdiffusion >>
rect 212 85 213 86 
<< pdiffusion >>
rect 213 85 214 86 
<< pdiffusion >>
rect 214 85 215 86 
<< pdiffusion >>
rect 215 85 216 86 
<< m1 >>
rect 217 85 218 86 
<< m1 >>
rect 221 85 222 86 
<< pdiffusion >>
rect 228 85 229 86 
<< pdiffusion >>
rect 229 85 230 86 
<< pdiffusion >>
rect 230 85 231 86 
<< pdiffusion >>
rect 231 85 232 86 
<< pdiffusion >>
rect 232 85 233 86 
<< pdiffusion >>
rect 233 85 234 86 
<< pdiffusion >>
rect 246 85 247 86 
<< pdiffusion >>
rect 247 85 248 86 
<< pdiffusion >>
rect 248 85 249 86 
<< pdiffusion >>
rect 249 85 250 86 
<< pdiffusion >>
rect 250 85 251 86 
<< pdiffusion >>
rect 251 85 252 86 
<< m1 >>
rect 253 85 254 86 
<< m1 >>
rect 260 85 261 86 
<< m1 >>
rect 262 85 263 86 
<< pdiffusion >>
rect 264 85 265 86 
<< pdiffusion >>
rect 265 85 266 86 
<< pdiffusion >>
rect 266 85 267 86 
<< pdiffusion >>
rect 267 85 268 86 
<< pdiffusion >>
rect 268 85 269 86 
<< pdiffusion >>
rect 269 85 270 86 
<< pdiffusion >>
rect 282 85 283 86 
<< pdiffusion >>
rect 283 85 284 86 
<< pdiffusion >>
rect 284 85 285 86 
<< pdiffusion >>
rect 285 85 286 86 
<< pdiffusion >>
rect 286 85 287 86 
<< pdiffusion >>
rect 287 85 288 86 
<< m1 >>
rect 298 85 299 86 
<< pdiffusion >>
rect 300 85 301 86 
<< pdiffusion >>
rect 301 85 302 86 
<< pdiffusion >>
rect 302 85 303 86 
<< pdiffusion >>
rect 303 85 304 86 
<< pdiffusion >>
rect 304 85 305 86 
<< pdiffusion >>
rect 305 85 306 86 
<< pdiffusion >>
rect 318 85 319 86 
<< pdiffusion >>
rect 319 85 320 86 
<< pdiffusion >>
rect 320 85 321 86 
<< pdiffusion >>
rect 321 85 322 86 
<< pdiffusion >>
rect 322 85 323 86 
<< pdiffusion >>
rect 323 85 324 86 
<< pdiffusion >>
rect 336 85 337 86 
<< pdiffusion >>
rect 337 85 338 86 
<< pdiffusion >>
rect 338 85 339 86 
<< pdiffusion >>
rect 339 85 340 86 
<< pdiffusion >>
rect 340 85 341 86 
<< pdiffusion >>
rect 341 85 342 86 
<< m1 >>
rect 352 85 353 86 
<< pdiffusion >>
rect 354 85 355 86 
<< pdiffusion >>
rect 355 85 356 86 
<< pdiffusion >>
rect 356 85 357 86 
<< pdiffusion >>
rect 357 85 358 86 
<< pdiffusion >>
rect 358 85 359 86 
<< pdiffusion >>
rect 359 85 360 86 
<< pdiffusion >>
rect 372 85 373 86 
<< pdiffusion >>
rect 373 85 374 86 
<< pdiffusion >>
rect 374 85 375 86 
<< pdiffusion >>
rect 375 85 376 86 
<< pdiffusion >>
rect 376 85 377 86 
<< pdiffusion >>
rect 377 85 378 86 
<< m1 >>
rect 379 85 380 86 
<< pdiffusion >>
rect 390 85 391 86 
<< pdiffusion >>
rect 391 85 392 86 
<< pdiffusion >>
rect 392 85 393 86 
<< pdiffusion >>
rect 393 85 394 86 
<< pdiffusion >>
rect 394 85 395 86 
<< pdiffusion >>
rect 395 85 396 86 
<< pdiffusion >>
rect 408 85 409 86 
<< pdiffusion >>
rect 409 85 410 86 
<< pdiffusion >>
rect 410 85 411 86 
<< pdiffusion >>
rect 411 85 412 86 
<< pdiffusion >>
rect 412 85 413 86 
<< pdiffusion >>
rect 413 85 414 86 
<< m1 >>
rect 424 85 425 86 
<< pdiffusion >>
rect 426 85 427 86 
<< pdiffusion >>
rect 427 85 428 86 
<< pdiffusion >>
rect 428 85 429 86 
<< pdiffusion >>
rect 429 85 430 86 
<< pdiffusion >>
rect 430 85 431 86 
<< pdiffusion >>
rect 431 85 432 86 
<< pdiffusion >>
rect 444 85 445 86 
<< pdiffusion >>
rect 445 85 446 86 
<< pdiffusion >>
rect 446 85 447 86 
<< pdiffusion >>
rect 447 85 448 86 
<< pdiffusion >>
rect 448 85 449 86 
<< pdiffusion >>
rect 449 85 450 86 
<< m1 >>
rect 451 85 452 86 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< pdiffusion >>
rect 30 86 31 87 
<< pdiffusion >>
rect 31 86 32 87 
<< pdiffusion >>
rect 32 86 33 87 
<< pdiffusion >>
rect 33 86 34 87 
<< pdiffusion >>
rect 34 86 35 87 
<< pdiffusion >>
rect 35 86 36 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 91 86 92 87 
<< pdiffusion >>
rect 102 86 103 87 
<< pdiffusion >>
rect 103 86 104 87 
<< pdiffusion >>
rect 104 86 105 87 
<< pdiffusion >>
rect 105 86 106 87 
<< pdiffusion >>
rect 106 86 107 87 
<< pdiffusion >>
rect 107 86 108 87 
<< pdiffusion >>
rect 120 86 121 87 
<< pdiffusion >>
rect 121 86 122 87 
<< pdiffusion >>
rect 122 86 123 87 
<< pdiffusion >>
rect 123 86 124 87 
<< pdiffusion >>
rect 124 86 125 87 
<< pdiffusion >>
rect 125 86 126 87 
<< pdiffusion >>
rect 138 86 139 87 
<< pdiffusion >>
rect 139 86 140 87 
<< pdiffusion >>
rect 140 86 141 87 
<< pdiffusion >>
rect 141 86 142 87 
<< pdiffusion >>
rect 142 86 143 87 
<< pdiffusion >>
rect 143 86 144 87 
<< pdiffusion >>
rect 156 86 157 87 
<< pdiffusion >>
rect 157 86 158 87 
<< pdiffusion >>
rect 158 86 159 87 
<< pdiffusion >>
rect 159 86 160 87 
<< pdiffusion >>
rect 160 86 161 87 
<< pdiffusion >>
rect 161 86 162 87 
<< pdiffusion >>
rect 174 86 175 87 
<< pdiffusion >>
rect 175 86 176 87 
<< pdiffusion >>
rect 176 86 177 87 
<< pdiffusion >>
rect 177 86 178 87 
<< pdiffusion >>
rect 178 86 179 87 
<< pdiffusion >>
rect 179 86 180 87 
<< m1 >>
rect 190 86 191 87 
<< pdiffusion >>
rect 192 86 193 87 
<< pdiffusion >>
rect 193 86 194 87 
<< pdiffusion >>
rect 194 86 195 87 
<< pdiffusion >>
rect 195 86 196 87 
<< pdiffusion >>
rect 196 86 197 87 
<< pdiffusion >>
rect 197 86 198 87 
<< m1 >>
rect 199 86 200 87 
<< pdiffusion >>
rect 210 86 211 87 
<< pdiffusion >>
rect 211 86 212 87 
<< pdiffusion >>
rect 212 86 213 87 
<< pdiffusion >>
rect 213 86 214 87 
<< pdiffusion >>
rect 214 86 215 87 
<< pdiffusion >>
rect 215 86 216 87 
<< m1 >>
rect 217 86 218 87 
<< m1 >>
rect 221 86 222 87 
<< pdiffusion >>
rect 228 86 229 87 
<< pdiffusion >>
rect 229 86 230 87 
<< pdiffusion >>
rect 230 86 231 87 
<< pdiffusion >>
rect 231 86 232 87 
<< pdiffusion >>
rect 232 86 233 87 
<< pdiffusion >>
rect 233 86 234 87 
<< pdiffusion >>
rect 246 86 247 87 
<< pdiffusion >>
rect 247 86 248 87 
<< pdiffusion >>
rect 248 86 249 87 
<< pdiffusion >>
rect 249 86 250 87 
<< pdiffusion >>
rect 250 86 251 87 
<< pdiffusion >>
rect 251 86 252 87 
<< m1 >>
rect 253 86 254 87 
<< m1 >>
rect 260 86 261 87 
<< m1 >>
rect 262 86 263 87 
<< pdiffusion >>
rect 264 86 265 87 
<< pdiffusion >>
rect 265 86 266 87 
<< pdiffusion >>
rect 266 86 267 87 
<< pdiffusion >>
rect 267 86 268 87 
<< pdiffusion >>
rect 268 86 269 87 
<< pdiffusion >>
rect 269 86 270 87 
<< pdiffusion >>
rect 282 86 283 87 
<< pdiffusion >>
rect 283 86 284 87 
<< pdiffusion >>
rect 284 86 285 87 
<< pdiffusion >>
rect 285 86 286 87 
<< pdiffusion >>
rect 286 86 287 87 
<< pdiffusion >>
rect 287 86 288 87 
<< m1 >>
rect 298 86 299 87 
<< pdiffusion >>
rect 300 86 301 87 
<< pdiffusion >>
rect 301 86 302 87 
<< pdiffusion >>
rect 302 86 303 87 
<< pdiffusion >>
rect 303 86 304 87 
<< pdiffusion >>
rect 304 86 305 87 
<< pdiffusion >>
rect 305 86 306 87 
<< pdiffusion >>
rect 318 86 319 87 
<< pdiffusion >>
rect 319 86 320 87 
<< pdiffusion >>
rect 320 86 321 87 
<< pdiffusion >>
rect 321 86 322 87 
<< pdiffusion >>
rect 322 86 323 87 
<< pdiffusion >>
rect 323 86 324 87 
<< pdiffusion >>
rect 336 86 337 87 
<< pdiffusion >>
rect 337 86 338 87 
<< pdiffusion >>
rect 338 86 339 87 
<< pdiffusion >>
rect 339 86 340 87 
<< pdiffusion >>
rect 340 86 341 87 
<< pdiffusion >>
rect 341 86 342 87 
<< m1 >>
rect 352 86 353 87 
<< pdiffusion >>
rect 354 86 355 87 
<< pdiffusion >>
rect 355 86 356 87 
<< pdiffusion >>
rect 356 86 357 87 
<< pdiffusion >>
rect 357 86 358 87 
<< pdiffusion >>
rect 358 86 359 87 
<< pdiffusion >>
rect 359 86 360 87 
<< pdiffusion >>
rect 372 86 373 87 
<< pdiffusion >>
rect 373 86 374 87 
<< pdiffusion >>
rect 374 86 375 87 
<< pdiffusion >>
rect 375 86 376 87 
<< pdiffusion >>
rect 376 86 377 87 
<< pdiffusion >>
rect 377 86 378 87 
<< m1 >>
rect 379 86 380 87 
<< pdiffusion >>
rect 390 86 391 87 
<< pdiffusion >>
rect 391 86 392 87 
<< pdiffusion >>
rect 392 86 393 87 
<< pdiffusion >>
rect 393 86 394 87 
<< pdiffusion >>
rect 394 86 395 87 
<< pdiffusion >>
rect 395 86 396 87 
<< pdiffusion >>
rect 408 86 409 87 
<< pdiffusion >>
rect 409 86 410 87 
<< pdiffusion >>
rect 410 86 411 87 
<< pdiffusion >>
rect 411 86 412 87 
<< pdiffusion >>
rect 412 86 413 87 
<< pdiffusion >>
rect 413 86 414 87 
<< m1 >>
rect 424 86 425 87 
<< pdiffusion >>
rect 426 86 427 87 
<< pdiffusion >>
rect 427 86 428 87 
<< pdiffusion >>
rect 428 86 429 87 
<< pdiffusion >>
rect 429 86 430 87 
<< pdiffusion >>
rect 430 86 431 87 
<< pdiffusion >>
rect 431 86 432 87 
<< pdiffusion >>
rect 444 86 445 87 
<< pdiffusion >>
rect 445 86 446 87 
<< pdiffusion >>
rect 446 86 447 87 
<< pdiffusion >>
rect 447 86 448 87 
<< pdiffusion >>
rect 448 86 449 87 
<< pdiffusion >>
rect 449 86 450 87 
<< m1 >>
rect 451 86 452 87 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< pdiffusion >>
rect 30 87 31 88 
<< pdiffusion >>
rect 31 87 32 88 
<< pdiffusion >>
rect 32 87 33 88 
<< pdiffusion >>
rect 33 87 34 88 
<< pdiffusion >>
rect 34 87 35 88 
<< pdiffusion >>
rect 35 87 36 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 91 87 92 88 
<< pdiffusion >>
rect 102 87 103 88 
<< pdiffusion >>
rect 103 87 104 88 
<< pdiffusion >>
rect 104 87 105 88 
<< pdiffusion >>
rect 105 87 106 88 
<< pdiffusion >>
rect 106 87 107 88 
<< pdiffusion >>
rect 107 87 108 88 
<< pdiffusion >>
rect 120 87 121 88 
<< pdiffusion >>
rect 121 87 122 88 
<< pdiffusion >>
rect 122 87 123 88 
<< pdiffusion >>
rect 123 87 124 88 
<< pdiffusion >>
rect 124 87 125 88 
<< pdiffusion >>
rect 125 87 126 88 
<< pdiffusion >>
rect 138 87 139 88 
<< pdiffusion >>
rect 139 87 140 88 
<< pdiffusion >>
rect 140 87 141 88 
<< pdiffusion >>
rect 141 87 142 88 
<< pdiffusion >>
rect 142 87 143 88 
<< pdiffusion >>
rect 143 87 144 88 
<< pdiffusion >>
rect 156 87 157 88 
<< pdiffusion >>
rect 157 87 158 88 
<< pdiffusion >>
rect 158 87 159 88 
<< pdiffusion >>
rect 159 87 160 88 
<< pdiffusion >>
rect 160 87 161 88 
<< pdiffusion >>
rect 161 87 162 88 
<< pdiffusion >>
rect 174 87 175 88 
<< pdiffusion >>
rect 175 87 176 88 
<< pdiffusion >>
rect 176 87 177 88 
<< pdiffusion >>
rect 177 87 178 88 
<< pdiffusion >>
rect 178 87 179 88 
<< pdiffusion >>
rect 179 87 180 88 
<< m1 >>
rect 190 87 191 88 
<< pdiffusion >>
rect 192 87 193 88 
<< pdiffusion >>
rect 193 87 194 88 
<< pdiffusion >>
rect 194 87 195 88 
<< pdiffusion >>
rect 195 87 196 88 
<< pdiffusion >>
rect 196 87 197 88 
<< pdiffusion >>
rect 197 87 198 88 
<< m1 >>
rect 199 87 200 88 
<< pdiffusion >>
rect 210 87 211 88 
<< pdiffusion >>
rect 211 87 212 88 
<< pdiffusion >>
rect 212 87 213 88 
<< pdiffusion >>
rect 213 87 214 88 
<< pdiffusion >>
rect 214 87 215 88 
<< pdiffusion >>
rect 215 87 216 88 
<< m1 >>
rect 217 87 218 88 
<< m1 >>
rect 221 87 222 88 
<< pdiffusion >>
rect 228 87 229 88 
<< pdiffusion >>
rect 229 87 230 88 
<< pdiffusion >>
rect 230 87 231 88 
<< pdiffusion >>
rect 231 87 232 88 
<< pdiffusion >>
rect 232 87 233 88 
<< pdiffusion >>
rect 233 87 234 88 
<< pdiffusion >>
rect 246 87 247 88 
<< pdiffusion >>
rect 247 87 248 88 
<< pdiffusion >>
rect 248 87 249 88 
<< pdiffusion >>
rect 249 87 250 88 
<< pdiffusion >>
rect 250 87 251 88 
<< pdiffusion >>
rect 251 87 252 88 
<< m1 >>
rect 253 87 254 88 
<< m1 >>
rect 260 87 261 88 
<< m1 >>
rect 262 87 263 88 
<< pdiffusion >>
rect 264 87 265 88 
<< pdiffusion >>
rect 265 87 266 88 
<< pdiffusion >>
rect 266 87 267 88 
<< pdiffusion >>
rect 267 87 268 88 
<< pdiffusion >>
rect 268 87 269 88 
<< pdiffusion >>
rect 269 87 270 88 
<< pdiffusion >>
rect 282 87 283 88 
<< pdiffusion >>
rect 283 87 284 88 
<< pdiffusion >>
rect 284 87 285 88 
<< pdiffusion >>
rect 285 87 286 88 
<< pdiffusion >>
rect 286 87 287 88 
<< pdiffusion >>
rect 287 87 288 88 
<< m1 >>
rect 298 87 299 88 
<< pdiffusion >>
rect 300 87 301 88 
<< pdiffusion >>
rect 301 87 302 88 
<< pdiffusion >>
rect 302 87 303 88 
<< pdiffusion >>
rect 303 87 304 88 
<< pdiffusion >>
rect 304 87 305 88 
<< pdiffusion >>
rect 305 87 306 88 
<< pdiffusion >>
rect 318 87 319 88 
<< pdiffusion >>
rect 319 87 320 88 
<< pdiffusion >>
rect 320 87 321 88 
<< pdiffusion >>
rect 321 87 322 88 
<< pdiffusion >>
rect 322 87 323 88 
<< pdiffusion >>
rect 323 87 324 88 
<< pdiffusion >>
rect 336 87 337 88 
<< pdiffusion >>
rect 337 87 338 88 
<< pdiffusion >>
rect 338 87 339 88 
<< pdiffusion >>
rect 339 87 340 88 
<< pdiffusion >>
rect 340 87 341 88 
<< pdiffusion >>
rect 341 87 342 88 
<< m1 >>
rect 352 87 353 88 
<< pdiffusion >>
rect 354 87 355 88 
<< pdiffusion >>
rect 355 87 356 88 
<< pdiffusion >>
rect 356 87 357 88 
<< pdiffusion >>
rect 357 87 358 88 
<< pdiffusion >>
rect 358 87 359 88 
<< pdiffusion >>
rect 359 87 360 88 
<< pdiffusion >>
rect 372 87 373 88 
<< pdiffusion >>
rect 373 87 374 88 
<< pdiffusion >>
rect 374 87 375 88 
<< pdiffusion >>
rect 375 87 376 88 
<< pdiffusion >>
rect 376 87 377 88 
<< pdiffusion >>
rect 377 87 378 88 
<< m1 >>
rect 379 87 380 88 
<< pdiffusion >>
rect 390 87 391 88 
<< pdiffusion >>
rect 391 87 392 88 
<< pdiffusion >>
rect 392 87 393 88 
<< pdiffusion >>
rect 393 87 394 88 
<< pdiffusion >>
rect 394 87 395 88 
<< pdiffusion >>
rect 395 87 396 88 
<< pdiffusion >>
rect 408 87 409 88 
<< pdiffusion >>
rect 409 87 410 88 
<< pdiffusion >>
rect 410 87 411 88 
<< pdiffusion >>
rect 411 87 412 88 
<< pdiffusion >>
rect 412 87 413 88 
<< pdiffusion >>
rect 413 87 414 88 
<< m1 >>
rect 424 87 425 88 
<< pdiffusion >>
rect 426 87 427 88 
<< pdiffusion >>
rect 427 87 428 88 
<< pdiffusion >>
rect 428 87 429 88 
<< pdiffusion >>
rect 429 87 430 88 
<< pdiffusion >>
rect 430 87 431 88 
<< pdiffusion >>
rect 431 87 432 88 
<< pdiffusion >>
rect 444 87 445 88 
<< pdiffusion >>
rect 445 87 446 88 
<< pdiffusion >>
rect 446 87 447 88 
<< pdiffusion >>
rect 447 87 448 88 
<< pdiffusion >>
rect 448 87 449 88 
<< pdiffusion >>
rect 449 87 450 88 
<< m1 >>
rect 451 87 452 88 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< pdiffusion >>
rect 30 88 31 89 
<< pdiffusion >>
rect 31 88 32 89 
<< pdiffusion >>
rect 32 88 33 89 
<< pdiffusion >>
rect 33 88 34 89 
<< pdiffusion >>
rect 34 88 35 89 
<< pdiffusion >>
rect 35 88 36 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 91 88 92 89 
<< pdiffusion >>
rect 102 88 103 89 
<< pdiffusion >>
rect 103 88 104 89 
<< pdiffusion >>
rect 104 88 105 89 
<< pdiffusion >>
rect 105 88 106 89 
<< pdiffusion >>
rect 106 88 107 89 
<< pdiffusion >>
rect 107 88 108 89 
<< pdiffusion >>
rect 120 88 121 89 
<< pdiffusion >>
rect 121 88 122 89 
<< pdiffusion >>
rect 122 88 123 89 
<< pdiffusion >>
rect 123 88 124 89 
<< pdiffusion >>
rect 124 88 125 89 
<< pdiffusion >>
rect 125 88 126 89 
<< pdiffusion >>
rect 138 88 139 89 
<< pdiffusion >>
rect 139 88 140 89 
<< pdiffusion >>
rect 140 88 141 89 
<< pdiffusion >>
rect 141 88 142 89 
<< pdiffusion >>
rect 142 88 143 89 
<< pdiffusion >>
rect 143 88 144 89 
<< pdiffusion >>
rect 156 88 157 89 
<< pdiffusion >>
rect 157 88 158 89 
<< pdiffusion >>
rect 158 88 159 89 
<< pdiffusion >>
rect 159 88 160 89 
<< pdiffusion >>
rect 160 88 161 89 
<< pdiffusion >>
rect 161 88 162 89 
<< pdiffusion >>
rect 174 88 175 89 
<< pdiffusion >>
rect 175 88 176 89 
<< pdiffusion >>
rect 176 88 177 89 
<< pdiffusion >>
rect 177 88 178 89 
<< pdiffusion >>
rect 178 88 179 89 
<< pdiffusion >>
rect 179 88 180 89 
<< m1 >>
rect 190 88 191 89 
<< pdiffusion >>
rect 192 88 193 89 
<< pdiffusion >>
rect 193 88 194 89 
<< pdiffusion >>
rect 194 88 195 89 
<< pdiffusion >>
rect 195 88 196 89 
<< pdiffusion >>
rect 196 88 197 89 
<< pdiffusion >>
rect 197 88 198 89 
<< m1 >>
rect 199 88 200 89 
<< pdiffusion >>
rect 210 88 211 89 
<< pdiffusion >>
rect 211 88 212 89 
<< pdiffusion >>
rect 212 88 213 89 
<< pdiffusion >>
rect 213 88 214 89 
<< pdiffusion >>
rect 214 88 215 89 
<< pdiffusion >>
rect 215 88 216 89 
<< m1 >>
rect 217 88 218 89 
<< m1 >>
rect 221 88 222 89 
<< pdiffusion >>
rect 228 88 229 89 
<< pdiffusion >>
rect 229 88 230 89 
<< pdiffusion >>
rect 230 88 231 89 
<< pdiffusion >>
rect 231 88 232 89 
<< pdiffusion >>
rect 232 88 233 89 
<< pdiffusion >>
rect 233 88 234 89 
<< pdiffusion >>
rect 246 88 247 89 
<< pdiffusion >>
rect 247 88 248 89 
<< pdiffusion >>
rect 248 88 249 89 
<< pdiffusion >>
rect 249 88 250 89 
<< pdiffusion >>
rect 250 88 251 89 
<< pdiffusion >>
rect 251 88 252 89 
<< m1 >>
rect 253 88 254 89 
<< m1 >>
rect 260 88 261 89 
<< m1 >>
rect 262 88 263 89 
<< pdiffusion >>
rect 264 88 265 89 
<< pdiffusion >>
rect 265 88 266 89 
<< pdiffusion >>
rect 266 88 267 89 
<< pdiffusion >>
rect 267 88 268 89 
<< pdiffusion >>
rect 268 88 269 89 
<< pdiffusion >>
rect 269 88 270 89 
<< pdiffusion >>
rect 282 88 283 89 
<< pdiffusion >>
rect 283 88 284 89 
<< pdiffusion >>
rect 284 88 285 89 
<< pdiffusion >>
rect 285 88 286 89 
<< pdiffusion >>
rect 286 88 287 89 
<< pdiffusion >>
rect 287 88 288 89 
<< m1 >>
rect 298 88 299 89 
<< pdiffusion >>
rect 300 88 301 89 
<< pdiffusion >>
rect 301 88 302 89 
<< pdiffusion >>
rect 302 88 303 89 
<< pdiffusion >>
rect 303 88 304 89 
<< pdiffusion >>
rect 304 88 305 89 
<< pdiffusion >>
rect 305 88 306 89 
<< pdiffusion >>
rect 318 88 319 89 
<< pdiffusion >>
rect 319 88 320 89 
<< pdiffusion >>
rect 320 88 321 89 
<< pdiffusion >>
rect 321 88 322 89 
<< pdiffusion >>
rect 322 88 323 89 
<< pdiffusion >>
rect 323 88 324 89 
<< pdiffusion >>
rect 336 88 337 89 
<< pdiffusion >>
rect 337 88 338 89 
<< pdiffusion >>
rect 338 88 339 89 
<< pdiffusion >>
rect 339 88 340 89 
<< pdiffusion >>
rect 340 88 341 89 
<< pdiffusion >>
rect 341 88 342 89 
<< m1 >>
rect 352 88 353 89 
<< pdiffusion >>
rect 354 88 355 89 
<< pdiffusion >>
rect 355 88 356 89 
<< pdiffusion >>
rect 356 88 357 89 
<< pdiffusion >>
rect 357 88 358 89 
<< pdiffusion >>
rect 358 88 359 89 
<< pdiffusion >>
rect 359 88 360 89 
<< pdiffusion >>
rect 372 88 373 89 
<< pdiffusion >>
rect 373 88 374 89 
<< pdiffusion >>
rect 374 88 375 89 
<< pdiffusion >>
rect 375 88 376 89 
<< pdiffusion >>
rect 376 88 377 89 
<< pdiffusion >>
rect 377 88 378 89 
<< m1 >>
rect 379 88 380 89 
<< pdiffusion >>
rect 390 88 391 89 
<< pdiffusion >>
rect 391 88 392 89 
<< pdiffusion >>
rect 392 88 393 89 
<< pdiffusion >>
rect 393 88 394 89 
<< pdiffusion >>
rect 394 88 395 89 
<< pdiffusion >>
rect 395 88 396 89 
<< pdiffusion >>
rect 408 88 409 89 
<< pdiffusion >>
rect 409 88 410 89 
<< pdiffusion >>
rect 410 88 411 89 
<< pdiffusion >>
rect 411 88 412 89 
<< pdiffusion >>
rect 412 88 413 89 
<< pdiffusion >>
rect 413 88 414 89 
<< m1 >>
rect 424 88 425 89 
<< pdiffusion >>
rect 426 88 427 89 
<< pdiffusion >>
rect 427 88 428 89 
<< pdiffusion >>
rect 428 88 429 89 
<< pdiffusion >>
rect 429 88 430 89 
<< pdiffusion >>
rect 430 88 431 89 
<< pdiffusion >>
rect 431 88 432 89 
<< pdiffusion >>
rect 444 88 445 89 
<< pdiffusion >>
rect 445 88 446 89 
<< pdiffusion >>
rect 446 88 447 89 
<< pdiffusion >>
rect 447 88 448 89 
<< pdiffusion >>
rect 448 88 449 89 
<< pdiffusion >>
rect 449 88 450 89 
<< m1 >>
rect 451 88 452 89 
<< pdiffusion >>
rect 12 89 13 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< m1 >>
rect 16 89 17 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< pdiffusion >>
rect 30 89 31 90 
<< pdiffusion >>
rect 31 89 32 90 
<< pdiffusion >>
rect 32 89 33 90 
<< pdiffusion >>
rect 33 89 34 90 
<< m1 >>
rect 34 89 35 90 
<< pdiffusion >>
rect 34 89 35 90 
<< pdiffusion >>
rect 35 89 36 90 
<< pdiffusion >>
rect 48 89 49 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< pdiffusion >>
rect 66 89 67 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< m1 >>
rect 70 89 71 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< pdiffusion >>
rect 84 89 85 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 91 89 92 90 
<< pdiffusion >>
rect 102 89 103 90 
<< pdiffusion >>
rect 103 89 104 90 
<< pdiffusion >>
rect 104 89 105 90 
<< pdiffusion >>
rect 105 89 106 90 
<< pdiffusion >>
rect 106 89 107 90 
<< pdiffusion >>
rect 107 89 108 90 
<< pdiffusion >>
rect 120 89 121 90 
<< pdiffusion >>
rect 121 89 122 90 
<< pdiffusion >>
rect 122 89 123 90 
<< pdiffusion >>
rect 123 89 124 90 
<< pdiffusion >>
rect 124 89 125 90 
<< pdiffusion >>
rect 125 89 126 90 
<< pdiffusion >>
rect 138 89 139 90 
<< pdiffusion >>
rect 139 89 140 90 
<< pdiffusion >>
rect 140 89 141 90 
<< pdiffusion >>
rect 141 89 142 90 
<< pdiffusion >>
rect 142 89 143 90 
<< pdiffusion >>
rect 143 89 144 90 
<< pdiffusion >>
rect 156 89 157 90 
<< pdiffusion >>
rect 157 89 158 90 
<< pdiffusion >>
rect 158 89 159 90 
<< pdiffusion >>
rect 159 89 160 90 
<< pdiffusion >>
rect 160 89 161 90 
<< pdiffusion >>
rect 161 89 162 90 
<< pdiffusion >>
rect 174 89 175 90 
<< pdiffusion >>
rect 175 89 176 90 
<< pdiffusion >>
rect 176 89 177 90 
<< pdiffusion >>
rect 177 89 178 90 
<< pdiffusion >>
rect 178 89 179 90 
<< pdiffusion >>
rect 179 89 180 90 
<< m1 >>
rect 190 89 191 90 
<< pdiffusion >>
rect 192 89 193 90 
<< pdiffusion >>
rect 193 89 194 90 
<< pdiffusion >>
rect 194 89 195 90 
<< pdiffusion >>
rect 195 89 196 90 
<< pdiffusion >>
rect 196 89 197 90 
<< pdiffusion >>
rect 197 89 198 90 
<< m1 >>
rect 199 89 200 90 
<< pdiffusion >>
rect 210 89 211 90 
<< pdiffusion >>
rect 211 89 212 90 
<< pdiffusion >>
rect 212 89 213 90 
<< pdiffusion >>
rect 213 89 214 90 
<< m1 >>
rect 214 89 215 90 
<< pdiffusion >>
rect 214 89 215 90 
<< pdiffusion >>
rect 215 89 216 90 
<< m1 >>
rect 217 89 218 90 
<< m1 >>
rect 221 89 222 90 
<< pdiffusion >>
rect 228 89 229 90 
<< pdiffusion >>
rect 229 89 230 90 
<< pdiffusion >>
rect 230 89 231 90 
<< pdiffusion >>
rect 231 89 232 90 
<< pdiffusion >>
rect 232 89 233 90 
<< pdiffusion >>
rect 233 89 234 90 
<< pdiffusion >>
rect 246 89 247 90 
<< pdiffusion >>
rect 247 89 248 90 
<< pdiffusion >>
rect 248 89 249 90 
<< pdiffusion >>
rect 249 89 250 90 
<< m1 >>
rect 250 89 251 90 
<< pdiffusion >>
rect 250 89 251 90 
<< pdiffusion >>
rect 251 89 252 90 
<< m1 >>
rect 253 89 254 90 
<< m1 >>
rect 260 89 261 90 
<< m1 >>
rect 262 89 263 90 
<< pdiffusion >>
rect 264 89 265 90 
<< pdiffusion >>
rect 265 89 266 90 
<< pdiffusion >>
rect 266 89 267 90 
<< pdiffusion >>
rect 267 89 268 90 
<< pdiffusion >>
rect 268 89 269 90 
<< pdiffusion >>
rect 269 89 270 90 
<< pdiffusion >>
rect 282 89 283 90 
<< pdiffusion >>
rect 283 89 284 90 
<< pdiffusion >>
rect 284 89 285 90 
<< pdiffusion >>
rect 285 89 286 90 
<< pdiffusion >>
rect 286 89 287 90 
<< pdiffusion >>
rect 287 89 288 90 
<< m1 >>
rect 298 89 299 90 
<< pdiffusion >>
rect 300 89 301 90 
<< pdiffusion >>
rect 301 89 302 90 
<< pdiffusion >>
rect 302 89 303 90 
<< pdiffusion >>
rect 303 89 304 90 
<< pdiffusion >>
rect 304 89 305 90 
<< pdiffusion >>
rect 305 89 306 90 
<< pdiffusion >>
rect 318 89 319 90 
<< pdiffusion >>
rect 319 89 320 90 
<< pdiffusion >>
rect 320 89 321 90 
<< pdiffusion >>
rect 321 89 322 90 
<< pdiffusion >>
rect 322 89 323 90 
<< pdiffusion >>
rect 323 89 324 90 
<< pdiffusion >>
rect 336 89 337 90 
<< m1 >>
rect 337 89 338 90 
<< pdiffusion >>
rect 337 89 338 90 
<< pdiffusion >>
rect 338 89 339 90 
<< pdiffusion >>
rect 339 89 340 90 
<< pdiffusion >>
rect 340 89 341 90 
<< pdiffusion >>
rect 341 89 342 90 
<< m1 >>
rect 352 89 353 90 
<< pdiffusion >>
rect 354 89 355 90 
<< pdiffusion >>
rect 355 89 356 90 
<< pdiffusion >>
rect 356 89 357 90 
<< pdiffusion >>
rect 357 89 358 90 
<< pdiffusion >>
rect 358 89 359 90 
<< pdiffusion >>
rect 359 89 360 90 
<< pdiffusion >>
rect 372 89 373 90 
<< pdiffusion >>
rect 373 89 374 90 
<< pdiffusion >>
rect 374 89 375 90 
<< pdiffusion >>
rect 375 89 376 90 
<< pdiffusion >>
rect 376 89 377 90 
<< pdiffusion >>
rect 377 89 378 90 
<< m1 >>
rect 379 89 380 90 
<< pdiffusion >>
rect 390 89 391 90 
<< pdiffusion >>
rect 391 89 392 90 
<< pdiffusion >>
rect 392 89 393 90 
<< pdiffusion >>
rect 393 89 394 90 
<< pdiffusion >>
rect 394 89 395 90 
<< pdiffusion >>
rect 395 89 396 90 
<< pdiffusion >>
rect 408 89 409 90 
<< pdiffusion >>
rect 409 89 410 90 
<< pdiffusion >>
rect 410 89 411 90 
<< pdiffusion >>
rect 411 89 412 90 
<< pdiffusion >>
rect 412 89 413 90 
<< pdiffusion >>
rect 413 89 414 90 
<< m1 >>
rect 424 89 425 90 
<< pdiffusion >>
rect 426 89 427 90 
<< m1 >>
rect 427 89 428 90 
<< pdiffusion >>
rect 427 89 428 90 
<< pdiffusion >>
rect 428 89 429 90 
<< pdiffusion >>
rect 429 89 430 90 
<< pdiffusion >>
rect 430 89 431 90 
<< pdiffusion >>
rect 431 89 432 90 
<< pdiffusion >>
rect 444 89 445 90 
<< pdiffusion >>
rect 445 89 446 90 
<< pdiffusion >>
rect 446 89 447 90 
<< pdiffusion >>
rect 447 89 448 90 
<< pdiffusion >>
rect 448 89 449 90 
<< pdiffusion >>
rect 449 89 450 90 
<< m1 >>
rect 451 89 452 90 
<< m1 >>
rect 16 90 17 91 
<< m1 >>
rect 34 90 35 91 
<< m1 >>
rect 70 90 71 91 
<< m1 >>
rect 91 90 92 91 
<< m1 >>
rect 190 90 191 91 
<< m1 >>
rect 199 90 200 91 
<< m1 >>
rect 214 90 215 91 
<< m1 >>
rect 217 90 218 91 
<< m1 >>
rect 221 90 222 91 
<< m1 >>
rect 250 90 251 91 
<< m1 >>
rect 253 90 254 91 
<< m1 >>
rect 260 90 261 91 
<< m1 >>
rect 262 90 263 91 
<< m1 >>
rect 298 90 299 91 
<< m1 >>
rect 337 90 338 91 
<< m1 >>
rect 352 90 353 91 
<< m1 >>
rect 379 90 380 91 
<< m1 >>
rect 424 90 425 91 
<< m1 >>
rect 427 90 428 91 
<< m1 >>
rect 451 90 452 91 
<< m1 >>
rect 16 91 17 92 
<< m1 >>
rect 34 91 35 92 
<< m1 >>
rect 70 91 71 92 
<< m1 >>
rect 91 91 92 92 
<< m1 >>
rect 190 91 191 92 
<< m1 >>
rect 199 91 200 92 
<< m1 >>
rect 214 91 215 92 
<< m1 >>
rect 215 91 216 92 
<< m2 >>
rect 215 91 216 92 
<< m2c >>
rect 215 91 216 92 
<< m1 >>
rect 215 91 216 92 
<< m2 >>
rect 215 91 216 92 
<< m2 >>
rect 216 91 217 92 
<< m1 >>
rect 217 91 218 92 
<< m2 >>
rect 217 91 218 92 
<< m2 >>
rect 218 91 219 92 
<< m1 >>
rect 219 91 220 92 
<< m2 >>
rect 219 91 220 92 
<< m2c >>
rect 219 91 220 92 
<< m1 >>
rect 219 91 220 92 
<< m2 >>
rect 219 91 220 92 
<< m1 >>
rect 220 91 221 92 
<< m1 >>
rect 221 91 222 92 
<< m1 >>
rect 250 91 251 92 
<< m1 >>
rect 251 91 252 92 
<< m1 >>
rect 252 91 253 92 
<< m1 >>
rect 253 91 254 92 
<< m1 >>
rect 260 91 261 92 
<< m1 >>
rect 262 91 263 92 
<< m1 >>
rect 298 91 299 92 
<< m1 >>
rect 337 91 338 92 
<< m1 >>
rect 352 91 353 92 
<< m1 >>
rect 379 91 380 92 
<< m1 >>
rect 424 91 425 92 
<< m1 >>
rect 425 91 426 92 
<< m1 >>
rect 426 91 427 92 
<< m1 >>
rect 427 91 428 92 
<< m1 >>
rect 451 91 452 92 
<< m1 >>
rect 16 92 17 93 
<< m1 >>
rect 34 92 35 93 
<< m1 >>
rect 70 92 71 93 
<< m1 >>
rect 91 92 92 93 
<< m1 >>
rect 190 92 191 93 
<< m1 >>
rect 199 92 200 93 
<< m1 >>
rect 217 92 218 93 
<< m1 >>
rect 260 92 261 93 
<< m1 >>
rect 262 92 263 93 
<< m1 >>
rect 298 92 299 93 
<< m1 >>
rect 337 92 338 93 
<< m1 >>
rect 338 92 339 93 
<< m1 >>
rect 339 92 340 93 
<< m1 >>
rect 340 92 341 93 
<< m1 >>
rect 341 92 342 93 
<< m1 >>
rect 342 92 343 93 
<< m1 >>
rect 343 92 344 93 
<< m1 >>
rect 344 92 345 93 
<< m1 >>
rect 345 92 346 93 
<< m1 >>
rect 346 92 347 93 
<< m1 >>
rect 347 92 348 93 
<< m1 >>
rect 348 92 349 93 
<< m1 >>
rect 349 92 350 93 
<< m1 >>
rect 350 92 351 93 
<< m1 >>
rect 351 92 352 93 
<< m1 >>
rect 352 92 353 93 
<< m1 >>
rect 379 92 380 93 
<< m1 >>
rect 451 92 452 93 
<< m1 >>
rect 16 93 17 94 
<< m1 >>
rect 34 93 35 94 
<< m1 >>
rect 70 93 71 94 
<< m1 >>
rect 91 93 92 94 
<< m1 >>
rect 190 93 191 94 
<< m1 >>
rect 199 93 200 94 
<< m1 >>
rect 217 93 218 94 
<< m1 >>
rect 260 93 261 94 
<< m1 >>
rect 262 93 263 94 
<< m1 >>
rect 298 93 299 94 
<< m1 >>
rect 379 93 380 94 
<< m1 >>
rect 451 93 452 94 
<< m1 >>
rect 16 94 17 95 
<< m1 >>
rect 34 94 35 95 
<< m1 >>
rect 64 94 65 95 
<< m1 >>
rect 65 94 66 95 
<< m1 >>
rect 66 94 67 95 
<< m1 >>
rect 67 94 68 95 
<< m1 >>
rect 68 94 69 95 
<< m1 >>
rect 69 94 70 95 
<< m1 >>
rect 70 94 71 95 
<< m1 >>
rect 91 94 92 95 
<< m1 >>
rect 190 94 191 95 
<< m1 >>
rect 199 94 200 95 
<< m1 >>
rect 217 94 218 95 
<< m1 >>
rect 260 94 261 95 
<< m1 >>
rect 262 94 263 95 
<< m1 >>
rect 298 94 299 95 
<< m1 >>
rect 379 94 380 95 
<< m1 >>
rect 451 94 452 95 
<< m1 >>
rect 16 95 17 96 
<< m1 >>
rect 34 95 35 96 
<< m1 >>
rect 64 95 65 96 
<< m1 >>
rect 91 95 92 96 
<< m1 >>
rect 190 95 191 96 
<< m1 >>
rect 199 95 200 96 
<< m1 >>
rect 217 95 218 96 
<< m1 >>
rect 260 95 261 96 
<< m1 >>
rect 262 95 263 96 
<< m1 >>
rect 298 95 299 96 
<< m1 >>
rect 379 95 380 96 
<< m1 >>
rect 451 95 452 96 
<< m1 >>
rect 16 96 17 97 
<< m1 >>
rect 34 96 35 97 
<< m1 >>
rect 64 96 65 97 
<< m1 >>
rect 91 96 92 97 
<< m1 >>
rect 190 96 191 97 
<< m1 >>
rect 199 96 200 97 
<< m1 >>
rect 217 96 218 97 
<< m1 >>
rect 260 96 261 97 
<< m1 >>
rect 262 96 263 97 
<< m1 >>
rect 298 96 299 97 
<< m1 >>
rect 379 96 380 97 
<< m1 >>
rect 451 96 452 97 
<< m1 >>
rect 16 97 17 98 
<< m1 >>
rect 34 97 35 98 
<< m1 >>
rect 64 97 65 98 
<< m1 >>
rect 91 97 92 98 
<< m1 >>
rect 190 97 191 98 
<< m1 >>
rect 199 97 200 98 
<< m1 >>
rect 217 97 218 98 
<< m1 >>
rect 232 97 233 98 
<< m1 >>
rect 233 97 234 98 
<< m1 >>
rect 234 97 235 98 
<< m1 >>
rect 235 97 236 98 
<< m1 >>
rect 236 97 237 98 
<< m1 >>
rect 237 97 238 98 
<< m1 >>
rect 238 97 239 98 
<< m1 >>
rect 239 97 240 98 
<< m1 >>
rect 240 97 241 98 
<< m1 >>
rect 241 97 242 98 
<< m1 >>
rect 242 97 243 98 
<< m1 >>
rect 243 97 244 98 
<< m1 >>
rect 244 97 245 98 
<< m1 >>
rect 245 97 246 98 
<< m1 >>
rect 246 97 247 98 
<< m1 >>
rect 247 97 248 98 
<< m1 >>
rect 248 97 249 98 
<< m1 >>
rect 249 97 250 98 
<< m1 >>
rect 250 97 251 98 
<< m1 >>
rect 251 97 252 98 
<< m1 >>
rect 252 97 253 98 
<< m1 >>
rect 253 97 254 98 
<< m1 >>
rect 254 97 255 98 
<< m1 >>
rect 255 97 256 98 
<< m1 >>
rect 256 97 257 98 
<< m1 >>
rect 257 97 258 98 
<< m1 >>
rect 258 97 259 98 
<< m2 >>
rect 258 97 259 98 
<< m2c >>
rect 258 97 259 98 
<< m1 >>
rect 258 97 259 98 
<< m2 >>
rect 258 97 259 98 
<< m2 >>
rect 259 97 260 98 
<< m1 >>
rect 260 97 261 98 
<< m2 >>
rect 260 97 261 98 
<< m2 >>
rect 261 97 262 98 
<< m1 >>
rect 262 97 263 98 
<< m2 >>
rect 262 97 263 98 
<< m2 >>
rect 263 97 264 98 
<< m1 >>
rect 264 97 265 98 
<< m2 >>
rect 264 97 265 98 
<< m2c >>
rect 264 97 265 98 
<< m1 >>
rect 264 97 265 98 
<< m2 >>
rect 264 97 265 98 
<< m1 >>
rect 265 97 266 98 
<< m1 >>
rect 266 97 267 98 
<< m1 >>
rect 267 97 268 98 
<< m1 >>
rect 268 97 269 98 
<< m1 >>
rect 269 97 270 98 
<< m1 >>
rect 270 97 271 98 
<< m1 >>
rect 271 97 272 98 
<< m1 >>
rect 272 97 273 98 
<< m1 >>
rect 273 97 274 98 
<< m1 >>
rect 274 97 275 98 
<< m1 >>
rect 275 97 276 98 
<< m1 >>
rect 276 97 277 98 
<< m1 >>
rect 277 97 278 98 
<< m1 >>
rect 278 97 279 98 
<< m1 >>
rect 279 97 280 98 
<< m1 >>
rect 280 97 281 98 
<< m1 >>
rect 281 97 282 98 
<< m1 >>
rect 282 97 283 98 
<< m1 >>
rect 283 97 284 98 
<< m1 >>
rect 298 97 299 98 
<< m1 >>
rect 379 97 380 98 
<< m1 >>
rect 451 97 452 98 
<< m1 >>
rect 16 98 17 99 
<< m1 >>
rect 34 98 35 99 
<< m1 >>
rect 64 98 65 99 
<< m1 >>
rect 91 98 92 99 
<< m1 >>
rect 190 98 191 99 
<< m1 >>
rect 199 98 200 99 
<< m1 >>
rect 217 98 218 99 
<< m1 >>
rect 232 98 233 99 
<< m1 >>
rect 260 98 261 99 
<< m1 >>
rect 262 98 263 99 
<< m1 >>
rect 283 98 284 99 
<< m1 >>
rect 298 98 299 99 
<< m1 >>
rect 379 98 380 99 
<< m1 >>
rect 451 98 452 99 
<< m1 >>
rect 16 99 17 100 
<< m1 >>
rect 17 99 18 100 
<< m1 >>
rect 18 99 19 100 
<< m1 >>
rect 19 99 20 100 
<< m1 >>
rect 20 99 21 100 
<< m1 >>
rect 21 99 22 100 
<< m1 >>
rect 22 99 23 100 
<< m1 >>
rect 23 99 24 100 
<< m1 >>
rect 24 99 25 100 
<< m1 >>
rect 25 99 26 100 
<< m1 >>
rect 26 99 27 100 
<< m1 >>
rect 27 99 28 100 
<< m1 >>
rect 28 99 29 100 
<< m1 >>
rect 34 99 35 100 
<< m1 >>
rect 64 99 65 100 
<< m1 >>
rect 91 99 92 100 
<< m1 >>
rect 190 99 191 100 
<< m1 >>
rect 199 99 200 100 
<< m1 >>
rect 217 99 218 100 
<< m1 >>
rect 232 99 233 100 
<< m1 >>
rect 260 99 261 100 
<< m1 >>
rect 262 99 263 100 
<< m1 >>
rect 283 99 284 100 
<< m1 >>
rect 298 99 299 100 
<< m1 >>
rect 379 99 380 100 
<< m1 >>
rect 451 99 452 100 
<< m1 >>
rect 28 100 29 101 
<< m1 >>
rect 34 100 35 101 
<< m1 >>
rect 64 100 65 101 
<< m1 >>
rect 91 100 92 101 
<< m1 >>
rect 118 100 119 101 
<< m1 >>
rect 119 100 120 101 
<< m1 >>
rect 120 100 121 101 
<< m1 >>
rect 121 100 122 101 
<< m1 >>
rect 142 100 143 101 
<< m1 >>
rect 143 100 144 101 
<< m1 >>
rect 144 100 145 101 
<< m1 >>
rect 145 100 146 101 
<< m1 >>
rect 146 100 147 101 
<< m1 >>
rect 147 100 148 101 
<< m1 >>
rect 148 100 149 101 
<< m1 >>
rect 149 100 150 101 
<< m1 >>
rect 150 100 151 101 
<< m1 >>
rect 151 100 152 101 
<< m1 >>
rect 152 100 153 101 
<< m1 >>
rect 153 100 154 101 
<< m1 >>
rect 154 100 155 101 
<< m1 >>
rect 190 100 191 101 
<< m1 >>
rect 199 100 200 101 
<< m1 >>
rect 217 100 218 101 
<< m1 >>
rect 232 100 233 101 
<< m1 >>
rect 260 100 261 101 
<< m1 >>
rect 262 100 263 101 
<< m1 >>
rect 283 100 284 101 
<< m1 >>
rect 298 100 299 101 
<< m1 >>
rect 379 100 380 101 
<< m1 >>
rect 451 100 452 101 
<< m1 >>
rect 28 101 29 102 
<< m1 >>
rect 34 101 35 102 
<< m1 >>
rect 64 101 65 102 
<< m1 >>
rect 91 101 92 102 
<< m1 >>
rect 118 101 119 102 
<< m1 >>
rect 121 101 122 102 
<< m1 >>
rect 142 101 143 102 
<< m1 >>
rect 154 101 155 102 
<< m1 >>
rect 190 101 191 102 
<< m1 >>
rect 199 101 200 102 
<< m1 >>
rect 217 101 218 102 
<< m1 >>
rect 232 101 233 102 
<< m1 >>
rect 260 101 261 102 
<< m1 >>
rect 262 101 263 102 
<< m1 >>
rect 283 101 284 102 
<< m1 >>
rect 298 101 299 102 
<< m1 >>
rect 379 101 380 102 
<< m1 >>
rect 451 101 452 102 
<< pdiffusion >>
rect 12 102 13 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< m1 >>
rect 28 102 29 103 
<< pdiffusion >>
rect 30 102 31 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< pdiffusion >>
rect 33 102 34 103 
<< m1 >>
rect 34 102 35 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< pdiffusion >>
rect 48 102 49 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m1 >>
rect 64 102 65 103 
<< pdiffusion >>
rect 66 102 67 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< pdiffusion >>
rect 84 102 85 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< m1 >>
rect 91 102 92 103 
<< pdiffusion >>
rect 102 102 103 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< m1 >>
rect 118 102 119 103 
<< pdiffusion >>
rect 120 102 121 103 
<< m1 >>
rect 121 102 122 103 
<< pdiffusion >>
rect 121 102 122 103 
<< pdiffusion >>
rect 122 102 123 103 
<< pdiffusion >>
rect 123 102 124 103 
<< pdiffusion >>
rect 124 102 125 103 
<< pdiffusion >>
rect 125 102 126 103 
<< pdiffusion >>
rect 138 102 139 103 
<< pdiffusion >>
rect 139 102 140 103 
<< pdiffusion >>
rect 140 102 141 103 
<< pdiffusion >>
rect 141 102 142 103 
<< m1 >>
rect 142 102 143 103 
<< pdiffusion >>
rect 142 102 143 103 
<< pdiffusion >>
rect 143 102 144 103 
<< m1 >>
rect 154 102 155 103 
<< pdiffusion >>
rect 156 102 157 103 
<< pdiffusion >>
rect 157 102 158 103 
<< pdiffusion >>
rect 158 102 159 103 
<< pdiffusion >>
rect 159 102 160 103 
<< pdiffusion >>
rect 160 102 161 103 
<< pdiffusion >>
rect 161 102 162 103 
<< pdiffusion >>
rect 174 102 175 103 
<< pdiffusion >>
rect 175 102 176 103 
<< pdiffusion >>
rect 176 102 177 103 
<< pdiffusion >>
rect 177 102 178 103 
<< pdiffusion >>
rect 178 102 179 103 
<< pdiffusion >>
rect 179 102 180 103 
<< m1 >>
rect 190 102 191 103 
<< pdiffusion >>
rect 192 102 193 103 
<< pdiffusion >>
rect 193 102 194 103 
<< pdiffusion >>
rect 194 102 195 103 
<< pdiffusion >>
rect 195 102 196 103 
<< pdiffusion >>
rect 196 102 197 103 
<< pdiffusion >>
rect 197 102 198 103 
<< m1 >>
rect 199 102 200 103 
<< pdiffusion >>
rect 210 102 211 103 
<< pdiffusion >>
rect 211 102 212 103 
<< pdiffusion >>
rect 212 102 213 103 
<< pdiffusion >>
rect 213 102 214 103 
<< pdiffusion >>
rect 214 102 215 103 
<< pdiffusion >>
rect 215 102 216 103 
<< m1 >>
rect 217 102 218 103 
<< pdiffusion >>
rect 228 102 229 103 
<< pdiffusion >>
rect 229 102 230 103 
<< pdiffusion >>
rect 230 102 231 103 
<< pdiffusion >>
rect 231 102 232 103 
<< m1 >>
rect 232 102 233 103 
<< pdiffusion >>
rect 232 102 233 103 
<< pdiffusion >>
rect 233 102 234 103 
<< pdiffusion >>
rect 246 102 247 103 
<< pdiffusion >>
rect 247 102 248 103 
<< pdiffusion >>
rect 248 102 249 103 
<< pdiffusion >>
rect 249 102 250 103 
<< pdiffusion >>
rect 250 102 251 103 
<< pdiffusion >>
rect 251 102 252 103 
<< m1 >>
rect 260 102 261 103 
<< m1 >>
rect 262 102 263 103 
<< pdiffusion >>
rect 264 102 265 103 
<< pdiffusion >>
rect 265 102 266 103 
<< pdiffusion >>
rect 266 102 267 103 
<< pdiffusion >>
rect 267 102 268 103 
<< pdiffusion >>
rect 268 102 269 103 
<< pdiffusion >>
rect 269 102 270 103 
<< pdiffusion >>
rect 282 102 283 103 
<< m1 >>
rect 283 102 284 103 
<< pdiffusion >>
rect 283 102 284 103 
<< pdiffusion >>
rect 284 102 285 103 
<< pdiffusion >>
rect 285 102 286 103 
<< pdiffusion >>
rect 286 102 287 103 
<< pdiffusion >>
rect 287 102 288 103 
<< m1 >>
rect 298 102 299 103 
<< pdiffusion >>
rect 300 102 301 103 
<< pdiffusion >>
rect 301 102 302 103 
<< pdiffusion >>
rect 302 102 303 103 
<< pdiffusion >>
rect 303 102 304 103 
<< pdiffusion >>
rect 304 102 305 103 
<< pdiffusion >>
rect 305 102 306 103 
<< pdiffusion >>
rect 318 102 319 103 
<< pdiffusion >>
rect 319 102 320 103 
<< pdiffusion >>
rect 320 102 321 103 
<< pdiffusion >>
rect 321 102 322 103 
<< pdiffusion >>
rect 322 102 323 103 
<< pdiffusion >>
rect 323 102 324 103 
<< pdiffusion >>
rect 336 102 337 103 
<< pdiffusion >>
rect 337 102 338 103 
<< pdiffusion >>
rect 338 102 339 103 
<< pdiffusion >>
rect 339 102 340 103 
<< pdiffusion >>
rect 340 102 341 103 
<< pdiffusion >>
rect 341 102 342 103 
<< pdiffusion >>
rect 354 102 355 103 
<< pdiffusion >>
rect 355 102 356 103 
<< pdiffusion >>
rect 356 102 357 103 
<< pdiffusion >>
rect 357 102 358 103 
<< pdiffusion >>
rect 358 102 359 103 
<< pdiffusion >>
rect 359 102 360 103 
<< pdiffusion >>
rect 372 102 373 103 
<< pdiffusion >>
rect 373 102 374 103 
<< pdiffusion >>
rect 374 102 375 103 
<< pdiffusion >>
rect 375 102 376 103 
<< pdiffusion >>
rect 376 102 377 103 
<< pdiffusion >>
rect 377 102 378 103 
<< m1 >>
rect 379 102 380 103 
<< pdiffusion >>
rect 390 102 391 103 
<< pdiffusion >>
rect 391 102 392 103 
<< pdiffusion >>
rect 392 102 393 103 
<< pdiffusion >>
rect 393 102 394 103 
<< pdiffusion >>
rect 394 102 395 103 
<< pdiffusion >>
rect 395 102 396 103 
<< pdiffusion >>
rect 408 102 409 103 
<< pdiffusion >>
rect 409 102 410 103 
<< pdiffusion >>
rect 410 102 411 103 
<< pdiffusion >>
rect 411 102 412 103 
<< pdiffusion >>
rect 412 102 413 103 
<< pdiffusion >>
rect 413 102 414 103 
<< pdiffusion >>
rect 426 102 427 103 
<< pdiffusion >>
rect 427 102 428 103 
<< pdiffusion >>
rect 428 102 429 103 
<< pdiffusion >>
rect 429 102 430 103 
<< pdiffusion >>
rect 430 102 431 103 
<< pdiffusion >>
rect 431 102 432 103 
<< pdiffusion >>
rect 444 102 445 103 
<< pdiffusion >>
rect 445 102 446 103 
<< pdiffusion >>
rect 446 102 447 103 
<< pdiffusion >>
rect 447 102 448 103 
<< pdiffusion >>
rect 448 102 449 103 
<< pdiffusion >>
rect 449 102 450 103 
<< m1 >>
rect 451 102 452 103 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< m1 >>
rect 28 103 29 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m1 >>
rect 64 103 65 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< m1 >>
rect 91 103 92 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< m1 >>
rect 118 103 119 104 
<< pdiffusion >>
rect 120 103 121 104 
<< pdiffusion >>
rect 121 103 122 104 
<< pdiffusion >>
rect 122 103 123 104 
<< pdiffusion >>
rect 123 103 124 104 
<< pdiffusion >>
rect 124 103 125 104 
<< pdiffusion >>
rect 125 103 126 104 
<< pdiffusion >>
rect 138 103 139 104 
<< pdiffusion >>
rect 139 103 140 104 
<< pdiffusion >>
rect 140 103 141 104 
<< pdiffusion >>
rect 141 103 142 104 
<< pdiffusion >>
rect 142 103 143 104 
<< pdiffusion >>
rect 143 103 144 104 
<< m1 >>
rect 154 103 155 104 
<< pdiffusion >>
rect 156 103 157 104 
<< pdiffusion >>
rect 157 103 158 104 
<< pdiffusion >>
rect 158 103 159 104 
<< pdiffusion >>
rect 159 103 160 104 
<< pdiffusion >>
rect 160 103 161 104 
<< pdiffusion >>
rect 161 103 162 104 
<< pdiffusion >>
rect 174 103 175 104 
<< pdiffusion >>
rect 175 103 176 104 
<< pdiffusion >>
rect 176 103 177 104 
<< pdiffusion >>
rect 177 103 178 104 
<< pdiffusion >>
rect 178 103 179 104 
<< pdiffusion >>
rect 179 103 180 104 
<< m1 >>
rect 190 103 191 104 
<< pdiffusion >>
rect 192 103 193 104 
<< pdiffusion >>
rect 193 103 194 104 
<< pdiffusion >>
rect 194 103 195 104 
<< pdiffusion >>
rect 195 103 196 104 
<< pdiffusion >>
rect 196 103 197 104 
<< pdiffusion >>
rect 197 103 198 104 
<< m1 >>
rect 199 103 200 104 
<< pdiffusion >>
rect 210 103 211 104 
<< pdiffusion >>
rect 211 103 212 104 
<< pdiffusion >>
rect 212 103 213 104 
<< pdiffusion >>
rect 213 103 214 104 
<< pdiffusion >>
rect 214 103 215 104 
<< pdiffusion >>
rect 215 103 216 104 
<< m1 >>
rect 217 103 218 104 
<< pdiffusion >>
rect 228 103 229 104 
<< pdiffusion >>
rect 229 103 230 104 
<< pdiffusion >>
rect 230 103 231 104 
<< pdiffusion >>
rect 231 103 232 104 
<< pdiffusion >>
rect 232 103 233 104 
<< pdiffusion >>
rect 233 103 234 104 
<< pdiffusion >>
rect 246 103 247 104 
<< pdiffusion >>
rect 247 103 248 104 
<< pdiffusion >>
rect 248 103 249 104 
<< pdiffusion >>
rect 249 103 250 104 
<< pdiffusion >>
rect 250 103 251 104 
<< pdiffusion >>
rect 251 103 252 104 
<< m1 >>
rect 260 103 261 104 
<< m1 >>
rect 262 103 263 104 
<< pdiffusion >>
rect 264 103 265 104 
<< pdiffusion >>
rect 265 103 266 104 
<< pdiffusion >>
rect 266 103 267 104 
<< pdiffusion >>
rect 267 103 268 104 
<< pdiffusion >>
rect 268 103 269 104 
<< pdiffusion >>
rect 269 103 270 104 
<< pdiffusion >>
rect 282 103 283 104 
<< pdiffusion >>
rect 283 103 284 104 
<< pdiffusion >>
rect 284 103 285 104 
<< pdiffusion >>
rect 285 103 286 104 
<< pdiffusion >>
rect 286 103 287 104 
<< pdiffusion >>
rect 287 103 288 104 
<< m1 >>
rect 298 103 299 104 
<< pdiffusion >>
rect 300 103 301 104 
<< pdiffusion >>
rect 301 103 302 104 
<< pdiffusion >>
rect 302 103 303 104 
<< pdiffusion >>
rect 303 103 304 104 
<< pdiffusion >>
rect 304 103 305 104 
<< pdiffusion >>
rect 305 103 306 104 
<< pdiffusion >>
rect 318 103 319 104 
<< pdiffusion >>
rect 319 103 320 104 
<< pdiffusion >>
rect 320 103 321 104 
<< pdiffusion >>
rect 321 103 322 104 
<< pdiffusion >>
rect 322 103 323 104 
<< pdiffusion >>
rect 323 103 324 104 
<< pdiffusion >>
rect 336 103 337 104 
<< pdiffusion >>
rect 337 103 338 104 
<< pdiffusion >>
rect 338 103 339 104 
<< pdiffusion >>
rect 339 103 340 104 
<< pdiffusion >>
rect 340 103 341 104 
<< pdiffusion >>
rect 341 103 342 104 
<< pdiffusion >>
rect 354 103 355 104 
<< pdiffusion >>
rect 355 103 356 104 
<< pdiffusion >>
rect 356 103 357 104 
<< pdiffusion >>
rect 357 103 358 104 
<< pdiffusion >>
rect 358 103 359 104 
<< pdiffusion >>
rect 359 103 360 104 
<< pdiffusion >>
rect 372 103 373 104 
<< pdiffusion >>
rect 373 103 374 104 
<< pdiffusion >>
rect 374 103 375 104 
<< pdiffusion >>
rect 375 103 376 104 
<< pdiffusion >>
rect 376 103 377 104 
<< pdiffusion >>
rect 377 103 378 104 
<< m1 >>
rect 379 103 380 104 
<< pdiffusion >>
rect 390 103 391 104 
<< pdiffusion >>
rect 391 103 392 104 
<< pdiffusion >>
rect 392 103 393 104 
<< pdiffusion >>
rect 393 103 394 104 
<< pdiffusion >>
rect 394 103 395 104 
<< pdiffusion >>
rect 395 103 396 104 
<< pdiffusion >>
rect 408 103 409 104 
<< pdiffusion >>
rect 409 103 410 104 
<< pdiffusion >>
rect 410 103 411 104 
<< pdiffusion >>
rect 411 103 412 104 
<< pdiffusion >>
rect 412 103 413 104 
<< pdiffusion >>
rect 413 103 414 104 
<< pdiffusion >>
rect 426 103 427 104 
<< pdiffusion >>
rect 427 103 428 104 
<< pdiffusion >>
rect 428 103 429 104 
<< pdiffusion >>
rect 429 103 430 104 
<< pdiffusion >>
rect 430 103 431 104 
<< pdiffusion >>
rect 431 103 432 104 
<< pdiffusion >>
rect 444 103 445 104 
<< pdiffusion >>
rect 445 103 446 104 
<< pdiffusion >>
rect 446 103 447 104 
<< pdiffusion >>
rect 447 103 448 104 
<< pdiffusion >>
rect 448 103 449 104 
<< pdiffusion >>
rect 449 103 450 104 
<< m1 >>
rect 451 103 452 104 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< m1 >>
rect 28 104 29 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m1 >>
rect 64 104 65 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< m1 >>
rect 91 104 92 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< m1 >>
rect 118 104 119 105 
<< pdiffusion >>
rect 120 104 121 105 
<< pdiffusion >>
rect 121 104 122 105 
<< pdiffusion >>
rect 122 104 123 105 
<< pdiffusion >>
rect 123 104 124 105 
<< pdiffusion >>
rect 124 104 125 105 
<< pdiffusion >>
rect 125 104 126 105 
<< pdiffusion >>
rect 138 104 139 105 
<< pdiffusion >>
rect 139 104 140 105 
<< pdiffusion >>
rect 140 104 141 105 
<< pdiffusion >>
rect 141 104 142 105 
<< pdiffusion >>
rect 142 104 143 105 
<< pdiffusion >>
rect 143 104 144 105 
<< m1 >>
rect 154 104 155 105 
<< pdiffusion >>
rect 156 104 157 105 
<< pdiffusion >>
rect 157 104 158 105 
<< pdiffusion >>
rect 158 104 159 105 
<< pdiffusion >>
rect 159 104 160 105 
<< pdiffusion >>
rect 160 104 161 105 
<< pdiffusion >>
rect 161 104 162 105 
<< pdiffusion >>
rect 174 104 175 105 
<< pdiffusion >>
rect 175 104 176 105 
<< pdiffusion >>
rect 176 104 177 105 
<< pdiffusion >>
rect 177 104 178 105 
<< pdiffusion >>
rect 178 104 179 105 
<< pdiffusion >>
rect 179 104 180 105 
<< m1 >>
rect 190 104 191 105 
<< pdiffusion >>
rect 192 104 193 105 
<< pdiffusion >>
rect 193 104 194 105 
<< pdiffusion >>
rect 194 104 195 105 
<< pdiffusion >>
rect 195 104 196 105 
<< pdiffusion >>
rect 196 104 197 105 
<< pdiffusion >>
rect 197 104 198 105 
<< m1 >>
rect 199 104 200 105 
<< pdiffusion >>
rect 210 104 211 105 
<< pdiffusion >>
rect 211 104 212 105 
<< pdiffusion >>
rect 212 104 213 105 
<< pdiffusion >>
rect 213 104 214 105 
<< pdiffusion >>
rect 214 104 215 105 
<< pdiffusion >>
rect 215 104 216 105 
<< m1 >>
rect 217 104 218 105 
<< pdiffusion >>
rect 228 104 229 105 
<< pdiffusion >>
rect 229 104 230 105 
<< pdiffusion >>
rect 230 104 231 105 
<< pdiffusion >>
rect 231 104 232 105 
<< pdiffusion >>
rect 232 104 233 105 
<< pdiffusion >>
rect 233 104 234 105 
<< pdiffusion >>
rect 246 104 247 105 
<< pdiffusion >>
rect 247 104 248 105 
<< pdiffusion >>
rect 248 104 249 105 
<< pdiffusion >>
rect 249 104 250 105 
<< pdiffusion >>
rect 250 104 251 105 
<< pdiffusion >>
rect 251 104 252 105 
<< m1 >>
rect 260 104 261 105 
<< m1 >>
rect 262 104 263 105 
<< pdiffusion >>
rect 264 104 265 105 
<< pdiffusion >>
rect 265 104 266 105 
<< pdiffusion >>
rect 266 104 267 105 
<< pdiffusion >>
rect 267 104 268 105 
<< pdiffusion >>
rect 268 104 269 105 
<< pdiffusion >>
rect 269 104 270 105 
<< pdiffusion >>
rect 282 104 283 105 
<< pdiffusion >>
rect 283 104 284 105 
<< pdiffusion >>
rect 284 104 285 105 
<< pdiffusion >>
rect 285 104 286 105 
<< pdiffusion >>
rect 286 104 287 105 
<< pdiffusion >>
rect 287 104 288 105 
<< m1 >>
rect 298 104 299 105 
<< pdiffusion >>
rect 300 104 301 105 
<< pdiffusion >>
rect 301 104 302 105 
<< pdiffusion >>
rect 302 104 303 105 
<< pdiffusion >>
rect 303 104 304 105 
<< pdiffusion >>
rect 304 104 305 105 
<< pdiffusion >>
rect 305 104 306 105 
<< pdiffusion >>
rect 318 104 319 105 
<< pdiffusion >>
rect 319 104 320 105 
<< pdiffusion >>
rect 320 104 321 105 
<< pdiffusion >>
rect 321 104 322 105 
<< pdiffusion >>
rect 322 104 323 105 
<< pdiffusion >>
rect 323 104 324 105 
<< pdiffusion >>
rect 336 104 337 105 
<< pdiffusion >>
rect 337 104 338 105 
<< pdiffusion >>
rect 338 104 339 105 
<< pdiffusion >>
rect 339 104 340 105 
<< pdiffusion >>
rect 340 104 341 105 
<< pdiffusion >>
rect 341 104 342 105 
<< pdiffusion >>
rect 354 104 355 105 
<< pdiffusion >>
rect 355 104 356 105 
<< pdiffusion >>
rect 356 104 357 105 
<< pdiffusion >>
rect 357 104 358 105 
<< pdiffusion >>
rect 358 104 359 105 
<< pdiffusion >>
rect 359 104 360 105 
<< pdiffusion >>
rect 372 104 373 105 
<< pdiffusion >>
rect 373 104 374 105 
<< pdiffusion >>
rect 374 104 375 105 
<< pdiffusion >>
rect 375 104 376 105 
<< pdiffusion >>
rect 376 104 377 105 
<< pdiffusion >>
rect 377 104 378 105 
<< m1 >>
rect 379 104 380 105 
<< pdiffusion >>
rect 390 104 391 105 
<< pdiffusion >>
rect 391 104 392 105 
<< pdiffusion >>
rect 392 104 393 105 
<< pdiffusion >>
rect 393 104 394 105 
<< pdiffusion >>
rect 394 104 395 105 
<< pdiffusion >>
rect 395 104 396 105 
<< pdiffusion >>
rect 408 104 409 105 
<< pdiffusion >>
rect 409 104 410 105 
<< pdiffusion >>
rect 410 104 411 105 
<< pdiffusion >>
rect 411 104 412 105 
<< pdiffusion >>
rect 412 104 413 105 
<< pdiffusion >>
rect 413 104 414 105 
<< pdiffusion >>
rect 426 104 427 105 
<< pdiffusion >>
rect 427 104 428 105 
<< pdiffusion >>
rect 428 104 429 105 
<< pdiffusion >>
rect 429 104 430 105 
<< pdiffusion >>
rect 430 104 431 105 
<< pdiffusion >>
rect 431 104 432 105 
<< pdiffusion >>
rect 444 104 445 105 
<< pdiffusion >>
rect 445 104 446 105 
<< pdiffusion >>
rect 446 104 447 105 
<< pdiffusion >>
rect 447 104 448 105 
<< pdiffusion >>
rect 448 104 449 105 
<< pdiffusion >>
rect 449 104 450 105 
<< m1 >>
rect 451 104 452 105 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< m1 >>
rect 28 105 29 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m1 >>
rect 64 105 65 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< m1 >>
rect 91 105 92 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< m1 >>
rect 118 105 119 106 
<< pdiffusion >>
rect 120 105 121 106 
<< pdiffusion >>
rect 121 105 122 106 
<< pdiffusion >>
rect 122 105 123 106 
<< pdiffusion >>
rect 123 105 124 106 
<< pdiffusion >>
rect 124 105 125 106 
<< pdiffusion >>
rect 125 105 126 106 
<< pdiffusion >>
rect 138 105 139 106 
<< pdiffusion >>
rect 139 105 140 106 
<< pdiffusion >>
rect 140 105 141 106 
<< pdiffusion >>
rect 141 105 142 106 
<< pdiffusion >>
rect 142 105 143 106 
<< pdiffusion >>
rect 143 105 144 106 
<< m1 >>
rect 154 105 155 106 
<< pdiffusion >>
rect 156 105 157 106 
<< pdiffusion >>
rect 157 105 158 106 
<< pdiffusion >>
rect 158 105 159 106 
<< pdiffusion >>
rect 159 105 160 106 
<< pdiffusion >>
rect 160 105 161 106 
<< pdiffusion >>
rect 161 105 162 106 
<< pdiffusion >>
rect 174 105 175 106 
<< pdiffusion >>
rect 175 105 176 106 
<< pdiffusion >>
rect 176 105 177 106 
<< pdiffusion >>
rect 177 105 178 106 
<< pdiffusion >>
rect 178 105 179 106 
<< pdiffusion >>
rect 179 105 180 106 
<< m1 >>
rect 190 105 191 106 
<< pdiffusion >>
rect 192 105 193 106 
<< pdiffusion >>
rect 193 105 194 106 
<< pdiffusion >>
rect 194 105 195 106 
<< pdiffusion >>
rect 195 105 196 106 
<< pdiffusion >>
rect 196 105 197 106 
<< pdiffusion >>
rect 197 105 198 106 
<< m1 >>
rect 199 105 200 106 
<< pdiffusion >>
rect 210 105 211 106 
<< pdiffusion >>
rect 211 105 212 106 
<< pdiffusion >>
rect 212 105 213 106 
<< pdiffusion >>
rect 213 105 214 106 
<< pdiffusion >>
rect 214 105 215 106 
<< pdiffusion >>
rect 215 105 216 106 
<< m1 >>
rect 217 105 218 106 
<< pdiffusion >>
rect 228 105 229 106 
<< pdiffusion >>
rect 229 105 230 106 
<< pdiffusion >>
rect 230 105 231 106 
<< pdiffusion >>
rect 231 105 232 106 
<< pdiffusion >>
rect 232 105 233 106 
<< pdiffusion >>
rect 233 105 234 106 
<< pdiffusion >>
rect 246 105 247 106 
<< pdiffusion >>
rect 247 105 248 106 
<< pdiffusion >>
rect 248 105 249 106 
<< pdiffusion >>
rect 249 105 250 106 
<< pdiffusion >>
rect 250 105 251 106 
<< pdiffusion >>
rect 251 105 252 106 
<< m1 >>
rect 260 105 261 106 
<< m1 >>
rect 262 105 263 106 
<< pdiffusion >>
rect 264 105 265 106 
<< pdiffusion >>
rect 265 105 266 106 
<< pdiffusion >>
rect 266 105 267 106 
<< pdiffusion >>
rect 267 105 268 106 
<< pdiffusion >>
rect 268 105 269 106 
<< pdiffusion >>
rect 269 105 270 106 
<< pdiffusion >>
rect 282 105 283 106 
<< pdiffusion >>
rect 283 105 284 106 
<< pdiffusion >>
rect 284 105 285 106 
<< pdiffusion >>
rect 285 105 286 106 
<< pdiffusion >>
rect 286 105 287 106 
<< pdiffusion >>
rect 287 105 288 106 
<< m1 >>
rect 298 105 299 106 
<< pdiffusion >>
rect 300 105 301 106 
<< pdiffusion >>
rect 301 105 302 106 
<< pdiffusion >>
rect 302 105 303 106 
<< pdiffusion >>
rect 303 105 304 106 
<< pdiffusion >>
rect 304 105 305 106 
<< pdiffusion >>
rect 305 105 306 106 
<< pdiffusion >>
rect 318 105 319 106 
<< pdiffusion >>
rect 319 105 320 106 
<< pdiffusion >>
rect 320 105 321 106 
<< pdiffusion >>
rect 321 105 322 106 
<< pdiffusion >>
rect 322 105 323 106 
<< pdiffusion >>
rect 323 105 324 106 
<< pdiffusion >>
rect 336 105 337 106 
<< pdiffusion >>
rect 337 105 338 106 
<< pdiffusion >>
rect 338 105 339 106 
<< pdiffusion >>
rect 339 105 340 106 
<< pdiffusion >>
rect 340 105 341 106 
<< pdiffusion >>
rect 341 105 342 106 
<< pdiffusion >>
rect 354 105 355 106 
<< pdiffusion >>
rect 355 105 356 106 
<< pdiffusion >>
rect 356 105 357 106 
<< pdiffusion >>
rect 357 105 358 106 
<< pdiffusion >>
rect 358 105 359 106 
<< pdiffusion >>
rect 359 105 360 106 
<< pdiffusion >>
rect 372 105 373 106 
<< pdiffusion >>
rect 373 105 374 106 
<< pdiffusion >>
rect 374 105 375 106 
<< pdiffusion >>
rect 375 105 376 106 
<< pdiffusion >>
rect 376 105 377 106 
<< pdiffusion >>
rect 377 105 378 106 
<< m1 >>
rect 379 105 380 106 
<< pdiffusion >>
rect 390 105 391 106 
<< pdiffusion >>
rect 391 105 392 106 
<< pdiffusion >>
rect 392 105 393 106 
<< pdiffusion >>
rect 393 105 394 106 
<< pdiffusion >>
rect 394 105 395 106 
<< pdiffusion >>
rect 395 105 396 106 
<< pdiffusion >>
rect 408 105 409 106 
<< pdiffusion >>
rect 409 105 410 106 
<< pdiffusion >>
rect 410 105 411 106 
<< pdiffusion >>
rect 411 105 412 106 
<< pdiffusion >>
rect 412 105 413 106 
<< pdiffusion >>
rect 413 105 414 106 
<< pdiffusion >>
rect 426 105 427 106 
<< pdiffusion >>
rect 427 105 428 106 
<< pdiffusion >>
rect 428 105 429 106 
<< pdiffusion >>
rect 429 105 430 106 
<< pdiffusion >>
rect 430 105 431 106 
<< pdiffusion >>
rect 431 105 432 106 
<< pdiffusion >>
rect 444 105 445 106 
<< pdiffusion >>
rect 445 105 446 106 
<< pdiffusion >>
rect 446 105 447 106 
<< pdiffusion >>
rect 447 105 448 106 
<< pdiffusion >>
rect 448 105 449 106 
<< pdiffusion >>
rect 449 105 450 106 
<< m1 >>
rect 451 105 452 106 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< m1 >>
rect 28 106 29 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m1 >>
rect 64 106 65 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< m1 >>
rect 91 106 92 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< m1 >>
rect 118 106 119 107 
<< pdiffusion >>
rect 120 106 121 107 
<< pdiffusion >>
rect 121 106 122 107 
<< pdiffusion >>
rect 122 106 123 107 
<< pdiffusion >>
rect 123 106 124 107 
<< pdiffusion >>
rect 124 106 125 107 
<< pdiffusion >>
rect 125 106 126 107 
<< pdiffusion >>
rect 138 106 139 107 
<< pdiffusion >>
rect 139 106 140 107 
<< pdiffusion >>
rect 140 106 141 107 
<< pdiffusion >>
rect 141 106 142 107 
<< pdiffusion >>
rect 142 106 143 107 
<< pdiffusion >>
rect 143 106 144 107 
<< m1 >>
rect 154 106 155 107 
<< pdiffusion >>
rect 156 106 157 107 
<< pdiffusion >>
rect 157 106 158 107 
<< pdiffusion >>
rect 158 106 159 107 
<< pdiffusion >>
rect 159 106 160 107 
<< pdiffusion >>
rect 160 106 161 107 
<< pdiffusion >>
rect 161 106 162 107 
<< pdiffusion >>
rect 174 106 175 107 
<< pdiffusion >>
rect 175 106 176 107 
<< pdiffusion >>
rect 176 106 177 107 
<< pdiffusion >>
rect 177 106 178 107 
<< pdiffusion >>
rect 178 106 179 107 
<< pdiffusion >>
rect 179 106 180 107 
<< m1 >>
rect 190 106 191 107 
<< pdiffusion >>
rect 192 106 193 107 
<< pdiffusion >>
rect 193 106 194 107 
<< pdiffusion >>
rect 194 106 195 107 
<< pdiffusion >>
rect 195 106 196 107 
<< pdiffusion >>
rect 196 106 197 107 
<< pdiffusion >>
rect 197 106 198 107 
<< m1 >>
rect 199 106 200 107 
<< pdiffusion >>
rect 210 106 211 107 
<< pdiffusion >>
rect 211 106 212 107 
<< pdiffusion >>
rect 212 106 213 107 
<< pdiffusion >>
rect 213 106 214 107 
<< pdiffusion >>
rect 214 106 215 107 
<< pdiffusion >>
rect 215 106 216 107 
<< m1 >>
rect 217 106 218 107 
<< pdiffusion >>
rect 228 106 229 107 
<< pdiffusion >>
rect 229 106 230 107 
<< pdiffusion >>
rect 230 106 231 107 
<< pdiffusion >>
rect 231 106 232 107 
<< pdiffusion >>
rect 232 106 233 107 
<< pdiffusion >>
rect 233 106 234 107 
<< pdiffusion >>
rect 246 106 247 107 
<< pdiffusion >>
rect 247 106 248 107 
<< pdiffusion >>
rect 248 106 249 107 
<< pdiffusion >>
rect 249 106 250 107 
<< pdiffusion >>
rect 250 106 251 107 
<< pdiffusion >>
rect 251 106 252 107 
<< m1 >>
rect 260 106 261 107 
<< m1 >>
rect 262 106 263 107 
<< pdiffusion >>
rect 264 106 265 107 
<< pdiffusion >>
rect 265 106 266 107 
<< pdiffusion >>
rect 266 106 267 107 
<< pdiffusion >>
rect 267 106 268 107 
<< pdiffusion >>
rect 268 106 269 107 
<< pdiffusion >>
rect 269 106 270 107 
<< pdiffusion >>
rect 282 106 283 107 
<< pdiffusion >>
rect 283 106 284 107 
<< pdiffusion >>
rect 284 106 285 107 
<< pdiffusion >>
rect 285 106 286 107 
<< pdiffusion >>
rect 286 106 287 107 
<< pdiffusion >>
rect 287 106 288 107 
<< m1 >>
rect 298 106 299 107 
<< pdiffusion >>
rect 300 106 301 107 
<< pdiffusion >>
rect 301 106 302 107 
<< pdiffusion >>
rect 302 106 303 107 
<< pdiffusion >>
rect 303 106 304 107 
<< pdiffusion >>
rect 304 106 305 107 
<< pdiffusion >>
rect 305 106 306 107 
<< pdiffusion >>
rect 318 106 319 107 
<< pdiffusion >>
rect 319 106 320 107 
<< pdiffusion >>
rect 320 106 321 107 
<< pdiffusion >>
rect 321 106 322 107 
<< pdiffusion >>
rect 322 106 323 107 
<< pdiffusion >>
rect 323 106 324 107 
<< pdiffusion >>
rect 336 106 337 107 
<< pdiffusion >>
rect 337 106 338 107 
<< pdiffusion >>
rect 338 106 339 107 
<< pdiffusion >>
rect 339 106 340 107 
<< pdiffusion >>
rect 340 106 341 107 
<< pdiffusion >>
rect 341 106 342 107 
<< pdiffusion >>
rect 354 106 355 107 
<< pdiffusion >>
rect 355 106 356 107 
<< pdiffusion >>
rect 356 106 357 107 
<< pdiffusion >>
rect 357 106 358 107 
<< pdiffusion >>
rect 358 106 359 107 
<< pdiffusion >>
rect 359 106 360 107 
<< pdiffusion >>
rect 372 106 373 107 
<< pdiffusion >>
rect 373 106 374 107 
<< pdiffusion >>
rect 374 106 375 107 
<< pdiffusion >>
rect 375 106 376 107 
<< pdiffusion >>
rect 376 106 377 107 
<< pdiffusion >>
rect 377 106 378 107 
<< m1 >>
rect 379 106 380 107 
<< pdiffusion >>
rect 390 106 391 107 
<< pdiffusion >>
rect 391 106 392 107 
<< pdiffusion >>
rect 392 106 393 107 
<< pdiffusion >>
rect 393 106 394 107 
<< pdiffusion >>
rect 394 106 395 107 
<< pdiffusion >>
rect 395 106 396 107 
<< pdiffusion >>
rect 408 106 409 107 
<< pdiffusion >>
rect 409 106 410 107 
<< pdiffusion >>
rect 410 106 411 107 
<< pdiffusion >>
rect 411 106 412 107 
<< pdiffusion >>
rect 412 106 413 107 
<< pdiffusion >>
rect 413 106 414 107 
<< pdiffusion >>
rect 426 106 427 107 
<< pdiffusion >>
rect 427 106 428 107 
<< pdiffusion >>
rect 428 106 429 107 
<< pdiffusion >>
rect 429 106 430 107 
<< pdiffusion >>
rect 430 106 431 107 
<< pdiffusion >>
rect 431 106 432 107 
<< pdiffusion >>
rect 444 106 445 107 
<< pdiffusion >>
rect 445 106 446 107 
<< pdiffusion >>
rect 446 106 447 107 
<< pdiffusion >>
rect 447 106 448 107 
<< pdiffusion >>
rect 448 106 449 107 
<< pdiffusion >>
rect 449 106 450 107 
<< m1 >>
rect 451 106 452 107 
<< pdiffusion >>
rect 12 107 13 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< m1 >>
rect 28 107 29 108 
<< pdiffusion >>
rect 30 107 31 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< pdiffusion >>
rect 48 107 49 108 
<< m1 >>
rect 49 107 50 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m1 >>
rect 64 107 65 108 
<< pdiffusion >>
rect 66 107 67 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< m1 >>
rect 70 107 71 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< pdiffusion >>
rect 84 107 85 108 
<< m1 >>
rect 85 107 86 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< m1 >>
rect 91 107 92 108 
<< pdiffusion >>
rect 102 107 103 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< m1 >>
rect 118 107 119 108 
<< pdiffusion >>
rect 120 107 121 108 
<< pdiffusion >>
rect 121 107 122 108 
<< pdiffusion >>
rect 122 107 123 108 
<< pdiffusion >>
rect 123 107 124 108 
<< pdiffusion >>
rect 124 107 125 108 
<< pdiffusion >>
rect 125 107 126 108 
<< pdiffusion >>
rect 138 107 139 108 
<< m1 >>
rect 139 107 140 108 
<< pdiffusion >>
rect 139 107 140 108 
<< pdiffusion >>
rect 140 107 141 108 
<< pdiffusion >>
rect 141 107 142 108 
<< m1 >>
rect 142 107 143 108 
<< pdiffusion >>
rect 142 107 143 108 
<< pdiffusion >>
rect 143 107 144 108 
<< m1 >>
rect 154 107 155 108 
<< pdiffusion >>
rect 156 107 157 108 
<< pdiffusion >>
rect 157 107 158 108 
<< pdiffusion >>
rect 158 107 159 108 
<< pdiffusion >>
rect 159 107 160 108 
<< pdiffusion >>
rect 160 107 161 108 
<< pdiffusion >>
rect 161 107 162 108 
<< pdiffusion >>
rect 174 107 175 108 
<< pdiffusion >>
rect 175 107 176 108 
<< pdiffusion >>
rect 176 107 177 108 
<< pdiffusion >>
rect 177 107 178 108 
<< pdiffusion >>
rect 178 107 179 108 
<< pdiffusion >>
rect 179 107 180 108 
<< m1 >>
rect 190 107 191 108 
<< pdiffusion >>
rect 192 107 193 108 
<< pdiffusion >>
rect 193 107 194 108 
<< pdiffusion >>
rect 194 107 195 108 
<< pdiffusion >>
rect 195 107 196 108 
<< pdiffusion >>
rect 196 107 197 108 
<< pdiffusion >>
rect 197 107 198 108 
<< m1 >>
rect 199 107 200 108 
<< pdiffusion >>
rect 210 107 211 108 
<< pdiffusion >>
rect 211 107 212 108 
<< pdiffusion >>
rect 212 107 213 108 
<< pdiffusion >>
rect 213 107 214 108 
<< pdiffusion >>
rect 214 107 215 108 
<< pdiffusion >>
rect 215 107 216 108 
<< m1 >>
rect 217 107 218 108 
<< pdiffusion >>
rect 228 107 229 108 
<< pdiffusion >>
rect 229 107 230 108 
<< pdiffusion >>
rect 230 107 231 108 
<< pdiffusion >>
rect 231 107 232 108 
<< pdiffusion >>
rect 232 107 233 108 
<< pdiffusion >>
rect 233 107 234 108 
<< pdiffusion >>
rect 246 107 247 108 
<< pdiffusion >>
rect 247 107 248 108 
<< pdiffusion >>
rect 248 107 249 108 
<< pdiffusion >>
rect 249 107 250 108 
<< pdiffusion >>
rect 250 107 251 108 
<< pdiffusion >>
rect 251 107 252 108 
<< m1 >>
rect 260 107 261 108 
<< m1 >>
rect 262 107 263 108 
<< pdiffusion >>
rect 264 107 265 108 
<< pdiffusion >>
rect 265 107 266 108 
<< pdiffusion >>
rect 266 107 267 108 
<< pdiffusion >>
rect 267 107 268 108 
<< m1 >>
rect 268 107 269 108 
<< pdiffusion >>
rect 268 107 269 108 
<< pdiffusion >>
rect 269 107 270 108 
<< pdiffusion >>
rect 282 107 283 108 
<< pdiffusion >>
rect 283 107 284 108 
<< pdiffusion >>
rect 284 107 285 108 
<< pdiffusion >>
rect 285 107 286 108 
<< m1 >>
rect 286 107 287 108 
<< pdiffusion >>
rect 286 107 287 108 
<< pdiffusion >>
rect 287 107 288 108 
<< m1 >>
rect 298 107 299 108 
<< pdiffusion >>
rect 300 107 301 108 
<< pdiffusion >>
rect 301 107 302 108 
<< pdiffusion >>
rect 302 107 303 108 
<< pdiffusion >>
rect 303 107 304 108 
<< pdiffusion >>
rect 304 107 305 108 
<< pdiffusion >>
rect 305 107 306 108 
<< pdiffusion >>
rect 318 107 319 108 
<< m1 >>
rect 319 107 320 108 
<< pdiffusion >>
rect 319 107 320 108 
<< pdiffusion >>
rect 320 107 321 108 
<< pdiffusion >>
rect 321 107 322 108 
<< pdiffusion >>
rect 322 107 323 108 
<< pdiffusion >>
rect 323 107 324 108 
<< pdiffusion >>
rect 336 107 337 108 
<< pdiffusion >>
rect 337 107 338 108 
<< pdiffusion >>
rect 338 107 339 108 
<< pdiffusion >>
rect 339 107 340 108 
<< pdiffusion >>
rect 340 107 341 108 
<< pdiffusion >>
rect 341 107 342 108 
<< pdiffusion >>
rect 354 107 355 108 
<< pdiffusion >>
rect 355 107 356 108 
<< pdiffusion >>
rect 356 107 357 108 
<< pdiffusion >>
rect 357 107 358 108 
<< pdiffusion >>
rect 358 107 359 108 
<< pdiffusion >>
rect 359 107 360 108 
<< pdiffusion >>
rect 372 107 373 108 
<< m1 >>
rect 373 107 374 108 
<< pdiffusion >>
rect 373 107 374 108 
<< pdiffusion >>
rect 374 107 375 108 
<< pdiffusion >>
rect 375 107 376 108 
<< pdiffusion >>
rect 376 107 377 108 
<< pdiffusion >>
rect 377 107 378 108 
<< m1 >>
rect 379 107 380 108 
<< pdiffusion >>
rect 390 107 391 108 
<< m1 >>
rect 391 107 392 108 
<< pdiffusion >>
rect 391 107 392 108 
<< pdiffusion >>
rect 392 107 393 108 
<< pdiffusion >>
rect 393 107 394 108 
<< pdiffusion >>
rect 394 107 395 108 
<< pdiffusion >>
rect 395 107 396 108 
<< pdiffusion >>
rect 408 107 409 108 
<< pdiffusion >>
rect 409 107 410 108 
<< pdiffusion >>
rect 410 107 411 108 
<< pdiffusion >>
rect 411 107 412 108 
<< pdiffusion >>
rect 412 107 413 108 
<< pdiffusion >>
rect 413 107 414 108 
<< pdiffusion >>
rect 426 107 427 108 
<< pdiffusion >>
rect 427 107 428 108 
<< pdiffusion >>
rect 428 107 429 108 
<< pdiffusion >>
rect 429 107 430 108 
<< pdiffusion >>
rect 430 107 431 108 
<< pdiffusion >>
rect 431 107 432 108 
<< pdiffusion >>
rect 444 107 445 108 
<< pdiffusion >>
rect 445 107 446 108 
<< pdiffusion >>
rect 446 107 447 108 
<< pdiffusion >>
rect 447 107 448 108 
<< pdiffusion >>
rect 448 107 449 108 
<< pdiffusion >>
rect 449 107 450 108 
<< m1 >>
rect 451 107 452 108 
<< m1 >>
rect 28 108 29 109 
<< m1 >>
rect 49 108 50 109 
<< m1 >>
rect 64 108 65 109 
<< m1 >>
rect 70 108 71 109 
<< m1 >>
rect 85 108 86 109 
<< m1 >>
rect 91 108 92 109 
<< m1 >>
rect 118 108 119 109 
<< m1 >>
rect 139 108 140 109 
<< m1 >>
rect 142 108 143 109 
<< m1 >>
rect 154 108 155 109 
<< m1 >>
rect 190 108 191 109 
<< m1 >>
rect 199 108 200 109 
<< m1 >>
rect 217 108 218 109 
<< m1 >>
rect 260 108 261 109 
<< m1 >>
rect 262 108 263 109 
<< m1 >>
rect 268 108 269 109 
<< m1 >>
rect 286 108 287 109 
<< m1 >>
rect 298 108 299 109 
<< m1 >>
rect 319 108 320 109 
<< m1 >>
rect 373 108 374 109 
<< m1 >>
rect 379 108 380 109 
<< m2 >>
rect 379 108 380 109 
<< m2c >>
rect 379 108 380 109 
<< m1 >>
rect 379 108 380 109 
<< m2 >>
rect 379 108 380 109 
<< m1 >>
rect 391 108 392 109 
<< m1 >>
rect 451 108 452 109 
<< m1 >>
rect 28 109 29 110 
<< m1 >>
rect 49 109 50 110 
<< m1 >>
rect 64 109 65 110 
<< m1 >>
rect 70 109 71 110 
<< m1 >>
rect 85 109 86 110 
<< m1 >>
rect 91 109 92 110 
<< m1 >>
rect 118 109 119 110 
<< m1 >>
rect 139 109 140 110 
<< m1 >>
rect 142 109 143 110 
<< m1 >>
rect 154 109 155 110 
<< m1 >>
rect 190 109 191 110 
<< m1 >>
rect 199 109 200 110 
<< m1 >>
rect 217 109 218 110 
<< m1 >>
rect 260 109 261 110 
<< m1 >>
rect 262 109 263 110 
<< m1 >>
rect 268 109 269 110 
<< m1 >>
rect 269 109 270 110 
<< m1 >>
rect 270 109 271 110 
<< m1 >>
rect 271 109 272 110 
<< m1 >>
rect 286 109 287 110 
<< m1 >>
rect 298 109 299 110 
<< m1 >>
rect 319 109 320 110 
<< m1 >>
rect 373 109 374 110 
<< m1 >>
rect 374 109 375 110 
<< m2 >>
rect 374 109 375 110 
<< m2c >>
rect 374 109 375 110 
<< m1 >>
rect 374 109 375 110 
<< m2 >>
rect 374 109 375 110 
<< m2 >>
rect 375 109 376 110 
<< m2 >>
rect 379 109 380 110 
<< m1 >>
rect 391 109 392 110 
<< m1 >>
rect 451 109 452 110 
<< m1 >>
rect 28 110 29 111 
<< m1 >>
rect 49 110 50 111 
<< m1 >>
rect 64 110 65 111 
<< m1 >>
rect 70 110 71 111 
<< m1 >>
rect 85 110 86 111 
<< m1 >>
rect 91 110 92 111 
<< m1 >>
rect 118 110 119 111 
<< m1 >>
rect 139 110 140 111 
<< m1 >>
rect 142 110 143 111 
<< m1 >>
rect 154 110 155 111 
<< m1 >>
rect 176 110 177 111 
<< m1 >>
rect 177 110 178 111 
<< m1 >>
rect 178 110 179 111 
<< m1 >>
rect 179 110 180 111 
<< m1 >>
rect 180 110 181 111 
<< m1 >>
rect 181 110 182 111 
<< m1 >>
rect 182 110 183 111 
<< m1 >>
rect 183 110 184 111 
<< m1 >>
rect 184 110 185 111 
<< m1 >>
rect 185 110 186 111 
<< m1 >>
rect 186 110 187 111 
<< m1 >>
rect 187 110 188 111 
<< m1 >>
rect 188 110 189 111 
<< m1 >>
rect 189 110 190 111 
<< m1 >>
rect 190 110 191 111 
<< m1 >>
rect 199 110 200 111 
<< m1 >>
rect 217 110 218 111 
<< m1 >>
rect 260 110 261 111 
<< m1 >>
rect 262 110 263 111 
<< m1 >>
rect 271 110 272 111 
<< m1 >>
rect 286 110 287 111 
<< m1 >>
rect 298 110 299 111 
<< m1 >>
rect 319 110 320 111 
<< m2 >>
rect 375 110 376 111 
<< m1 >>
rect 376 110 377 111 
<< m2 >>
rect 376 110 377 111 
<< m1 >>
rect 377 110 378 111 
<< m2 >>
rect 377 110 378 111 
<< m1 >>
rect 378 110 379 111 
<< m2 >>
rect 378 110 379 111 
<< m1 >>
rect 379 110 380 111 
<< m2 >>
rect 379 110 380 111 
<< m1 >>
rect 380 110 381 111 
<< m1 >>
rect 381 110 382 111 
<< m1 >>
rect 382 110 383 111 
<< m1 >>
rect 383 110 384 111 
<< m1 >>
rect 384 110 385 111 
<< m1 >>
rect 385 110 386 111 
<< m1 >>
rect 386 110 387 111 
<< m1 >>
rect 387 110 388 111 
<< m1 >>
rect 388 110 389 111 
<< m1 >>
rect 389 110 390 111 
<< m1 >>
rect 390 110 391 111 
<< m1 >>
rect 391 110 392 111 
<< m1 >>
rect 451 110 452 111 
<< m1 >>
rect 28 111 29 112 
<< m1 >>
rect 49 111 50 112 
<< m1 >>
rect 64 111 65 112 
<< m1 >>
rect 70 111 71 112 
<< m1 >>
rect 85 111 86 112 
<< m1 >>
rect 91 111 92 112 
<< m1 >>
rect 118 111 119 112 
<< m1 >>
rect 139 111 140 112 
<< m1 >>
rect 142 111 143 112 
<< m1 >>
rect 154 111 155 112 
<< m1 >>
rect 176 111 177 112 
<< m1 >>
rect 199 111 200 112 
<< m1 >>
rect 217 111 218 112 
<< m1 >>
rect 260 111 261 112 
<< m1 >>
rect 262 111 263 112 
<< m1 >>
rect 271 111 272 112 
<< m1 >>
rect 286 111 287 112 
<< m1 >>
rect 298 111 299 112 
<< m1 >>
rect 319 111 320 112 
<< m1 >>
rect 376 111 377 112 
<< m1 >>
rect 451 111 452 112 
<< m1 >>
rect 28 112 29 113 
<< m1 >>
rect 29 112 30 113 
<< m1 >>
rect 30 112 31 113 
<< m1 >>
rect 31 112 32 113 
<< m1 >>
rect 32 112 33 113 
<< m1 >>
rect 33 112 34 113 
<< m1 >>
rect 34 112 35 113 
<< m1 >>
rect 35 112 36 113 
<< m1 >>
rect 36 112 37 113 
<< m1 >>
rect 37 112 38 113 
<< m1 >>
rect 38 112 39 113 
<< m1 >>
rect 39 112 40 113 
<< m1 >>
rect 40 112 41 113 
<< m1 >>
rect 41 112 42 113 
<< m1 >>
rect 42 112 43 113 
<< m1 >>
rect 43 112 44 113 
<< m1 >>
rect 44 112 45 113 
<< m1 >>
rect 45 112 46 113 
<< m1 >>
rect 46 112 47 113 
<< m1 >>
rect 47 112 48 113 
<< m2 >>
rect 47 112 48 113 
<< m2c >>
rect 47 112 48 113 
<< m1 >>
rect 47 112 48 113 
<< m2 >>
rect 47 112 48 113 
<< m2 >>
rect 48 112 49 113 
<< m1 >>
rect 49 112 50 113 
<< m2 >>
rect 49 112 50 113 
<< m2 >>
rect 50 112 51 113 
<< m1 >>
rect 51 112 52 113 
<< m2 >>
rect 51 112 52 113 
<< m2c >>
rect 51 112 52 113 
<< m1 >>
rect 51 112 52 113 
<< m2 >>
rect 51 112 52 113 
<< m1 >>
rect 52 112 53 113 
<< m1 >>
rect 53 112 54 113 
<< m1 >>
rect 54 112 55 113 
<< m1 >>
rect 55 112 56 113 
<< m1 >>
rect 56 112 57 113 
<< m1 >>
rect 57 112 58 113 
<< m1 >>
rect 58 112 59 113 
<< m1 >>
rect 59 112 60 113 
<< m1 >>
rect 60 112 61 113 
<< m1 >>
rect 61 112 62 113 
<< m1 >>
rect 62 112 63 113 
<< m2 >>
rect 62 112 63 113 
<< m2c >>
rect 62 112 63 113 
<< m1 >>
rect 62 112 63 113 
<< m2 >>
rect 62 112 63 113 
<< m2 >>
rect 63 112 64 113 
<< m1 >>
rect 64 112 65 113 
<< m2 >>
rect 64 112 65 113 
<< m2 >>
rect 65 112 66 113 
<< m1 >>
rect 66 112 67 113 
<< m2 >>
rect 66 112 67 113 
<< m2c >>
rect 66 112 67 113 
<< m1 >>
rect 66 112 67 113 
<< m2 >>
rect 66 112 67 113 
<< m1 >>
rect 67 112 68 113 
<< m1 >>
rect 68 112 69 113 
<< m1 >>
rect 69 112 70 113 
<< m1 >>
rect 70 112 71 113 
<< m1 >>
rect 85 112 86 113 
<< m1 >>
rect 91 112 92 113 
<< m1 >>
rect 118 112 119 113 
<< m1 >>
rect 139 112 140 113 
<< m1 >>
rect 142 112 143 113 
<< m1 >>
rect 154 112 155 113 
<< m1 >>
rect 176 112 177 113 
<< m1 >>
rect 199 112 200 113 
<< m1 >>
rect 217 112 218 113 
<< m1 >>
rect 228 112 229 113 
<< m1 >>
rect 229 112 230 113 
<< m1 >>
rect 230 112 231 113 
<< m1 >>
rect 231 112 232 113 
<< m1 >>
rect 232 112 233 113 
<< m1 >>
rect 233 112 234 113 
<< m1 >>
rect 234 112 235 113 
<< m1 >>
rect 235 112 236 113 
<< m1 >>
rect 236 112 237 113 
<< m1 >>
rect 237 112 238 113 
<< m1 >>
rect 238 112 239 113 
<< m1 >>
rect 239 112 240 113 
<< m1 >>
rect 240 112 241 113 
<< m1 >>
rect 241 112 242 113 
<< m1 >>
rect 242 112 243 113 
<< m1 >>
rect 243 112 244 113 
<< m1 >>
rect 244 112 245 113 
<< m1 >>
rect 245 112 246 113 
<< m1 >>
rect 246 112 247 113 
<< m1 >>
rect 247 112 248 113 
<< m1 >>
rect 248 112 249 113 
<< m1 >>
rect 249 112 250 113 
<< m1 >>
rect 250 112 251 113 
<< m1 >>
rect 251 112 252 113 
<< m1 >>
rect 252 112 253 113 
<< m1 >>
rect 253 112 254 113 
<< m1 >>
rect 254 112 255 113 
<< m1 >>
rect 255 112 256 113 
<< m1 >>
rect 256 112 257 113 
<< m1 >>
rect 257 112 258 113 
<< m1 >>
rect 258 112 259 113 
<< m1 >>
rect 259 112 260 113 
<< m1 >>
rect 260 112 261 113 
<< m1 >>
rect 262 112 263 113 
<< m1 >>
rect 271 112 272 113 
<< m1 >>
rect 280 112 281 113 
<< m1 >>
rect 281 112 282 113 
<< m1 >>
rect 282 112 283 113 
<< m1 >>
rect 283 112 284 113 
<< m1 >>
rect 284 112 285 113 
<< m1 >>
rect 285 112 286 113 
<< m1 >>
rect 286 112 287 113 
<< m1 >>
rect 298 112 299 113 
<< m1 >>
rect 319 112 320 113 
<< m1 >>
rect 376 112 377 113 
<< m1 >>
rect 451 112 452 113 
<< m1 >>
rect 49 113 50 114 
<< m1 >>
rect 64 113 65 114 
<< m1 >>
rect 85 113 86 114 
<< m1 >>
rect 91 113 92 114 
<< m2 >>
rect 91 113 92 114 
<< m2c >>
rect 91 113 92 114 
<< m1 >>
rect 91 113 92 114 
<< m2 >>
rect 91 113 92 114 
<< m1 >>
rect 118 113 119 114 
<< m1 >>
rect 139 113 140 114 
<< m1 >>
rect 142 113 143 114 
<< m1 >>
rect 154 113 155 114 
<< m1 >>
rect 176 113 177 114 
<< m2 >>
rect 176 113 177 114 
<< m2c >>
rect 176 113 177 114 
<< m1 >>
rect 176 113 177 114 
<< m2 >>
rect 176 113 177 114 
<< m1 >>
rect 199 113 200 114 
<< m1 >>
rect 217 113 218 114 
<< m1 >>
rect 228 113 229 114 
<< m1 >>
rect 262 113 263 114 
<< m1 >>
rect 271 113 272 114 
<< m1 >>
rect 280 113 281 114 
<< m1 >>
rect 298 113 299 114 
<< m1 >>
rect 319 113 320 114 
<< m1 >>
rect 376 113 377 114 
<< m1 >>
rect 451 113 452 114 
<< m1 >>
rect 49 114 50 115 
<< m1 >>
rect 64 114 65 115 
<< m1 >>
rect 85 114 86 115 
<< m2 >>
rect 91 114 92 115 
<< m1 >>
rect 118 114 119 115 
<< m1 >>
rect 139 114 140 115 
<< m1 >>
rect 142 114 143 115 
<< m1 >>
rect 154 114 155 115 
<< m2 >>
rect 174 114 175 115 
<< m2 >>
rect 175 114 176 115 
<< m2 >>
rect 176 114 177 115 
<< m1 >>
rect 199 114 200 115 
<< m1 >>
rect 217 114 218 115 
<< m1 >>
rect 228 114 229 115 
<< m1 >>
rect 262 114 263 115 
<< m1 >>
rect 271 114 272 115 
<< m1 >>
rect 280 114 281 115 
<< m1 >>
rect 298 114 299 115 
<< m1 >>
rect 319 114 320 115 
<< m1 >>
rect 376 114 377 115 
<< m1 >>
rect 451 114 452 115 
<< m1 >>
rect 49 115 50 116 
<< m1 >>
rect 50 115 51 116 
<< m1 >>
rect 51 115 52 116 
<< m1 >>
rect 52 115 53 116 
<< m1 >>
rect 53 115 54 116 
<< m1 >>
rect 54 115 55 116 
<< m1 >>
rect 55 115 56 116 
<< m1 >>
rect 56 115 57 116 
<< m1 >>
rect 57 115 58 116 
<< m1 >>
rect 58 115 59 116 
<< m1 >>
rect 59 115 60 116 
<< m1 >>
rect 60 115 61 116 
<< m1 >>
rect 61 115 62 116 
<< m1 >>
rect 62 115 63 116 
<< m1 >>
rect 64 115 65 116 
<< m1 >>
rect 85 115 86 116 
<< m1 >>
rect 86 115 87 116 
<< m1 >>
rect 87 115 88 116 
<< m1 >>
rect 88 115 89 116 
<< m1 >>
rect 89 115 90 116 
<< m1 >>
rect 90 115 91 116 
<< m1 >>
rect 91 115 92 116 
<< m2 >>
rect 91 115 92 116 
<< m1 >>
rect 92 115 93 116 
<< m1 >>
rect 93 115 94 116 
<< m1 >>
rect 94 115 95 116 
<< m1 >>
rect 95 115 96 116 
<< m1 >>
rect 96 115 97 116 
<< m1 >>
rect 97 115 98 116 
<< m1 >>
rect 98 115 99 116 
<< m1 >>
rect 99 115 100 116 
<< m1 >>
rect 100 115 101 116 
<< m1 >>
rect 101 115 102 116 
<< m1 >>
rect 102 115 103 116 
<< m1 >>
rect 103 115 104 116 
<< m1 >>
rect 104 115 105 116 
<< m1 >>
rect 105 115 106 116 
<< m1 >>
rect 106 115 107 116 
<< m1 >>
rect 107 115 108 116 
<< m1 >>
rect 108 115 109 116 
<< m1 >>
rect 109 115 110 116 
<< m1 >>
rect 110 115 111 116 
<< m1 >>
rect 111 115 112 116 
<< m1 >>
rect 112 115 113 116 
<< m1 >>
rect 113 115 114 116 
<< m1 >>
rect 114 115 115 116 
<< m1 >>
rect 115 115 116 116 
<< m1 >>
rect 116 115 117 116 
<< m1 >>
rect 118 115 119 116 
<< m1 >>
rect 120 115 121 116 
<< m1 >>
rect 121 115 122 116 
<< m1 >>
rect 122 115 123 116 
<< m1 >>
rect 123 115 124 116 
<< m1 >>
rect 124 115 125 116 
<< m1 >>
rect 125 115 126 116 
<< m1 >>
rect 126 115 127 116 
<< m1 >>
rect 127 115 128 116 
<< m1 >>
rect 128 115 129 116 
<< m1 >>
rect 129 115 130 116 
<< m1 >>
rect 130 115 131 116 
<< m1 >>
rect 131 115 132 116 
<< m1 >>
rect 132 115 133 116 
<< m1 >>
rect 133 115 134 116 
<< m1 >>
rect 134 115 135 116 
<< m1 >>
rect 135 115 136 116 
<< m1 >>
rect 136 115 137 116 
<< m1 >>
rect 137 115 138 116 
<< m1 >>
rect 138 115 139 116 
<< m1 >>
rect 139 115 140 116 
<< m1 >>
rect 142 115 143 116 
<< m1 >>
rect 143 115 144 116 
<< m1 >>
rect 144 115 145 116 
<< m1 >>
rect 145 115 146 116 
<< m2 >>
rect 145 115 146 116 
<< m2c >>
rect 145 115 146 116 
<< m1 >>
rect 145 115 146 116 
<< m2 >>
rect 145 115 146 116 
<< m1 >>
rect 154 115 155 116 
<< m1 >>
rect 155 115 156 116 
<< m1 >>
rect 156 115 157 116 
<< m1 >>
rect 157 115 158 116 
<< m1 >>
rect 158 115 159 116 
<< m1 >>
rect 159 115 160 116 
<< m1 >>
rect 160 115 161 116 
<< m1 >>
rect 161 115 162 116 
<< m1 >>
rect 162 115 163 116 
<< m1 >>
rect 163 115 164 116 
<< m1 >>
rect 164 115 165 116 
<< m1 >>
rect 165 115 166 116 
<< m1 >>
rect 166 115 167 116 
<< m1 >>
rect 167 115 168 116 
<< m1 >>
rect 168 115 169 116 
<< m1 >>
rect 169 115 170 116 
<< m1 >>
rect 170 115 171 116 
<< m1 >>
rect 171 115 172 116 
<< m1 >>
rect 172 115 173 116 
<< m1 >>
rect 173 115 174 116 
<< m1 >>
rect 174 115 175 116 
<< m2 >>
rect 174 115 175 116 
<< m1 >>
rect 175 115 176 116 
<< m1 >>
rect 176 115 177 116 
<< m1 >>
rect 177 115 178 116 
<< m1 >>
rect 178 115 179 116 
<< m2 >>
rect 178 115 179 116 
<< m1 >>
rect 179 115 180 116 
<< m2 >>
rect 179 115 180 116 
<< m1 >>
rect 180 115 181 116 
<< m2 >>
rect 180 115 181 116 
<< m1 >>
rect 181 115 182 116 
<< m2 >>
rect 181 115 182 116 
<< m1 >>
rect 182 115 183 116 
<< m2 >>
rect 182 115 183 116 
<< m1 >>
rect 183 115 184 116 
<< m2 >>
rect 183 115 184 116 
<< m1 >>
rect 184 115 185 116 
<< m2 >>
rect 184 115 185 116 
<< m1 >>
rect 185 115 186 116 
<< m2 >>
rect 185 115 186 116 
<< m1 >>
rect 186 115 187 116 
<< m2 >>
rect 186 115 187 116 
<< m1 >>
rect 187 115 188 116 
<< m2 >>
rect 187 115 188 116 
<< m1 >>
rect 188 115 189 116 
<< m2 >>
rect 188 115 189 116 
<< m1 >>
rect 189 115 190 116 
<< m2 >>
rect 189 115 190 116 
<< m1 >>
rect 190 115 191 116 
<< m2 >>
rect 190 115 191 116 
<< m1 >>
rect 191 115 192 116 
<< m2 >>
rect 191 115 192 116 
<< m1 >>
rect 192 115 193 116 
<< m2 >>
rect 192 115 193 116 
<< m1 >>
rect 193 115 194 116 
<< m2 >>
rect 193 115 194 116 
<< m2 >>
rect 194 115 195 116 
<< m1 >>
rect 195 115 196 116 
<< m2 >>
rect 195 115 196 116 
<< m2c >>
rect 195 115 196 116 
<< m1 >>
rect 195 115 196 116 
<< m2 >>
rect 195 115 196 116 
<< m1 >>
rect 196 115 197 116 
<< m1 >>
rect 197 115 198 116 
<< m2 >>
rect 197 115 198 116 
<< m2c >>
rect 197 115 198 116 
<< m1 >>
rect 197 115 198 116 
<< m2 >>
rect 197 115 198 116 
<< m2 >>
rect 198 115 199 116 
<< m1 >>
rect 199 115 200 116 
<< m2 >>
rect 199 115 200 116 
<< m2 >>
rect 200 115 201 116 
<< m1 >>
rect 201 115 202 116 
<< m2 >>
rect 201 115 202 116 
<< m2c >>
rect 201 115 202 116 
<< m1 >>
rect 201 115 202 116 
<< m2 >>
rect 201 115 202 116 
<< m1 >>
rect 202 115 203 116 
<< m1 >>
rect 203 115 204 116 
<< m1 >>
rect 204 115 205 116 
<< m1 >>
rect 205 115 206 116 
<< m1 >>
rect 206 115 207 116 
<< m1 >>
rect 207 115 208 116 
<< m1 >>
rect 208 115 209 116 
<< m1 >>
rect 209 115 210 116 
<< m1 >>
rect 210 115 211 116 
<< m1 >>
rect 211 115 212 116 
<< m1 >>
rect 212 115 213 116 
<< m1 >>
rect 213 115 214 116 
<< m1 >>
rect 214 115 215 116 
<< m1 >>
rect 215 115 216 116 
<< m1 >>
rect 216 115 217 116 
<< m1 >>
rect 217 115 218 116 
<< m1 >>
rect 228 115 229 116 
<< m1 >>
rect 262 115 263 116 
<< m1 >>
rect 271 115 272 116 
<< m1 >>
rect 280 115 281 116 
<< m1 >>
rect 298 115 299 116 
<< m1 >>
rect 319 115 320 116 
<< m1 >>
rect 376 115 377 116 
<< m1 >>
rect 388 115 389 116 
<< m1 >>
rect 389 115 390 116 
<< m1 >>
rect 390 115 391 116 
<< m1 >>
rect 391 115 392 116 
<< m1 >>
rect 392 115 393 116 
<< m1 >>
rect 393 115 394 116 
<< m1 >>
rect 394 115 395 116 
<< m1 >>
rect 395 115 396 116 
<< m1 >>
rect 396 115 397 116 
<< m1 >>
rect 397 115 398 116 
<< m1 >>
rect 398 115 399 116 
<< m1 >>
rect 399 115 400 116 
<< m1 >>
rect 400 115 401 116 
<< m1 >>
rect 401 115 402 116 
<< m1 >>
rect 402 115 403 116 
<< m1 >>
rect 403 115 404 116 
<< m1 >>
rect 404 115 405 116 
<< m1 >>
rect 405 115 406 116 
<< m1 >>
rect 406 115 407 116 
<< m1 >>
rect 407 115 408 116 
<< m1 >>
rect 408 115 409 116 
<< m1 >>
rect 409 115 410 116 
<< m1 >>
rect 410 115 411 116 
<< m1 >>
rect 411 115 412 116 
<< m1 >>
rect 412 115 413 116 
<< m1 >>
rect 451 115 452 116 
<< m1 >>
rect 62 116 63 117 
<< m1 >>
rect 64 116 65 117 
<< m2 >>
rect 91 116 92 117 
<< m1 >>
rect 116 116 117 117 
<< m1 >>
rect 118 116 119 117 
<< m1 >>
rect 120 116 121 117 
<< m2 >>
rect 145 116 146 117 
<< m2 >>
rect 174 116 175 117 
<< m2 >>
rect 178 116 179 117 
<< m1 >>
rect 193 116 194 117 
<< m1 >>
rect 199 116 200 117 
<< m1 >>
rect 228 116 229 117 
<< m1 >>
rect 262 116 263 117 
<< m1 >>
rect 271 116 272 117 
<< m1 >>
rect 280 116 281 117 
<< m1 >>
rect 298 116 299 117 
<< m1 >>
rect 319 116 320 117 
<< m1 >>
rect 376 116 377 117 
<< m1 >>
rect 388 116 389 117 
<< m1 >>
rect 412 116 413 117 
<< m1 >>
rect 451 116 452 117 
<< m1 >>
rect 62 117 63 118 
<< m1 >>
rect 64 117 65 118 
<< m1 >>
rect 91 117 92 118 
<< m2 >>
rect 91 117 92 118 
<< m2c >>
rect 91 117 92 118 
<< m1 >>
rect 91 117 92 118 
<< m2 >>
rect 91 117 92 118 
<< m1 >>
rect 92 117 93 118 
<< m1 >>
rect 93 117 94 118 
<< m1 >>
rect 116 117 117 118 
<< m1 >>
rect 118 117 119 118 
<< m1 >>
rect 120 117 121 118 
<< m1 >>
rect 139 117 140 118 
<< m1 >>
rect 140 117 141 118 
<< m1 >>
rect 141 117 142 118 
<< m1 >>
rect 142 117 143 118 
<< m1 >>
rect 143 117 144 118 
<< m1 >>
rect 144 117 145 118 
<< m1 >>
rect 145 117 146 118 
<< m2 >>
rect 145 117 146 118 
<< m1 >>
rect 157 117 158 118 
<< m1 >>
rect 158 117 159 118 
<< m1 >>
rect 159 117 160 118 
<< m1 >>
rect 160 117 161 118 
<< m1 >>
rect 161 117 162 118 
<< m1 >>
rect 162 117 163 118 
<< m1 >>
rect 163 117 164 118 
<< m1 >>
rect 164 117 165 118 
<< m1 >>
rect 165 117 166 118 
<< m1 >>
rect 166 117 167 118 
<< m1 >>
rect 167 117 168 118 
<< m1 >>
rect 168 117 169 118 
<< m1 >>
rect 169 117 170 118 
<< m1 >>
rect 170 117 171 118 
<< m1 >>
rect 171 117 172 118 
<< m1 >>
rect 172 117 173 118 
<< m1 >>
rect 173 117 174 118 
<< m1 >>
rect 174 117 175 118 
<< m2 >>
rect 174 117 175 118 
<< m2c >>
rect 174 117 175 118 
<< m1 >>
rect 174 117 175 118 
<< m2 >>
rect 174 117 175 118 
<< m1 >>
rect 178 117 179 118 
<< m2 >>
rect 178 117 179 118 
<< m2c >>
rect 178 117 179 118 
<< m1 >>
rect 178 117 179 118 
<< m2 >>
rect 178 117 179 118 
<< m1 >>
rect 193 117 194 118 
<< m1 >>
rect 199 117 200 118 
<< m2 >>
rect 226 117 227 118 
<< m2 >>
rect 227 117 228 118 
<< m1 >>
rect 228 117 229 118 
<< m2 >>
rect 228 117 229 118 
<< m2c >>
rect 228 117 229 118 
<< m1 >>
rect 228 117 229 118 
<< m2 >>
rect 228 117 229 118 
<< m1 >>
rect 262 117 263 118 
<< m1 >>
rect 271 117 272 118 
<< m1 >>
rect 280 117 281 118 
<< m1 >>
rect 298 117 299 118 
<< m1 >>
rect 319 117 320 118 
<< m1 >>
rect 376 117 377 118 
<< m1 >>
rect 388 117 389 118 
<< m1 >>
rect 412 117 413 118 
<< m1 >>
rect 451 117 452 118 
<< m1 >>
rect 62 118 63 119 
<< m1 >>
rect 64 118 65 119 
<< m1 >>
rect 73 118 74 119 
<< m1 >>
rect 74 118 75 119 
<< m1 >>
rect 75 118 76 119 
<< m1 >>
rect 76 118 77 119 
<< m1 >>
rect 77 118 78 119 
<< m1 >>
rect 78 118 79 119 
<< m1 >>
rect 79 118 80 119 
<< m1 >>
rect 80 118 81 119 
<< m1 >>
rect 81 118 82 119 
<< m1 >>
rect 82 118 83 119 
<< m1 >>
rect 83 118 84 119 
<< m1 >>
rect 84 118 85 119 
<< m1 >>
rect 85 118 86 119 
<< m1 >>
rect 93 118 94 119 
<< m2 >>
rect 115 118 116 119 
<< m1 >>
rect 116 118 117 119 
<< m2 >>
rect 116 118 117 119 
<< m2 >>
rect 117 118 118 119 
<< m1 >>
rect 118 118 119 119 
<< m2 >>
rect 118 118 119 119 
<< m2 >>
rect 119 118 120 119 
<< m1 >>
rect 120 118 121 119 
<< m2 >>
rect 120 118 121 119 
<< m2c >>
rect 120 118 121 119 
<< m1 >>
rect 120 118 121 119 
<< m2 >>
rect 120 118 121 119 
<< m1 >>
rect 139 118 140 119 
<< m1 >>
rect 145 118 146 119 
<< m2 >>
rect 145 118 146 119 
<< m1 >>
rect 157 118 158 119 
<< m1 >>
rect 178 118 179 119 
<< m1 >>
rect 193 118 194 119 
<< m1 >>
rect 199 118 200 119 
<< m1 >>
rect 214 118 215 119 
<< m1 >>
rect 215 118 216 119 
<< m1 >>
rect 216 118 217 119 
<< m1 >>
rect 217 118 218 119 
<< m1 >>
rect 218 118 219 119 
<< m1 >>
rect 219 118 220 119 
<< m1 >>
rect 220 118 221 119 
<< m1 >>
rect 221 118 222 119 
<< m1 >>
rect 222 118 223 119 
<< m1 >>
rect 223 118 224 119 
<< m1 >>
rect 224 118 225 119 
<< m1 >>
rect 225 118 226 119 
<< m1 >>
rect 226 118 227 119 
<< m2 >>
rect 226 118 227 119 
<< m1 >>
rect 262 118 263 119 
<< m1 >>
rect 271 118 272 119 
<< m1 >>
rect 280 118 281 119 
<< m1 >>
rect 298 118 299 119 
<< m1 >>
rect 304 118 305 119 
<< m1 >>
rect 305 118 306 119 
<< m1 >>
rect 306 118 307 119 
<< m1 >>
rect 307 118 308 119 
<< m1 >>
rect 319 118 320 119 
<< m1 >>
rect 334 118 335 119 
<< m1 >>
rect 335 118 336 119 
<< m1 >>
rect 336 118 337 119 
<< m1 >>
rect 337 118 338 119 
<< m1 >>
rect 376 118 377 119 
<< m1 >>
rect 388 118 389 119 
<< m1 >>
rect 412 118 413 119 
<< m1 >>
rect 451 118 452 119 
<< m1 >>
rect 62 119 63 120 
<< m1 >>
rect 64 119 65 120 
<< m1 >>
rect 73 119 74 120 
<< m1 >>
rect 85 119 86 120 
<< m1 >>
rect 93 119 94 120 
<< m2 >>
rect 115 119 116 120 
<< m1 >>
rect 116 119 117 120 
<< m1 >>
rect 118 119 119 120 
<< m1 >>
rect 139 119 140 120 
<< m1 >>
rect 145 119 146 120 
<< m2 >>
rect 145 119 146 120 
<< m1 >>
rect 157 119 158 120 
<< m1 >>
rect 178 119 179 120 
<< m1 >>
rect 193 119 194 120 
<< m1 >>
rect 199 119 200 120 
<< m1 >>
rect 214 119 215 120 
<< m1 >>
rect 226 119 227 120 
<< m2 >>
rect 226 119 227 120 
<< m1 >>
rect 262 119 263 120 
<< m1 >>
rect 271 119 272 120 
<< m1 >>
rect 280 119 281 120 
<< m1 >>
rect 298 119 299 120 
<< m1 >>
rect 304 119 305 120 
<< m1 >>
rect 307 119 308 120 
<< m1 >>
rect 319 119 320 120 
<< m1 >>
rect 334 119 335 120 
<< m1 >>
rect 337 119 338 120 
<< m1 >>
rect 376 119 377 120 
<< m1 >>
rect 388 119 389 120 
<< m1 >>
rect 412 119 413 120 
<< m1 >>
rect 451 119 452 120 
<< pdiffusion >>
rect 12 120 13 121 
<< pdiffusion >>
rect 13 120 14 121 
<< pdiffusion >>
rect 14 120 15 121 
<< pdiffusion >>
rect 15 120 16 121 
<< pdiffusion >>
rect 16 120 17 121 
<< pdiffusion >>
rect 17 120 18 121 
<< pdiffusion >>
rect 30 120 31 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< pdiffusion >>
rect 48 120 49 121 
<< pdiffusion >>
rect 49 120 50 121 
<< pdiffusion >>
rect 50 120 51 121 
<< pdiffusion >>
rect 51 120 52 121 
<< pdiffusion >>
rect 52 120 53 121 
<< pdiffusion >>
rect 53 120 54 121 
<< m1 >>
rect 62 120 63 121 
<< m1 >>
rect 64 120 65 121 
<< pdiffusion >>
rect 66 120 67 121 
<< pdiffusion >>
rect 67 120 68 121 
<< pdiffusion >>
rect 68 120 69 121 
<< pdiffusion >>
rect 69 120 70 121 
<< pdiffusion >>
rect 70 120 71 121 
<< pdiffusion >>
rect 71 120 72 121 
<< m1 >>
rect 73 120 74 121 
<< pdiffusion >>
rect 84 120 85 121 
<< m1 >>
rect 85 120 86 121 
<< pdiffusion >>
rect 85 120 86 121 
<< pdiffusion >>
rect 86 120 87 121 
<< pdiffusion >>
rect 87 120 88 121 
<< pdiffusion >>
rect 88 120 89 121 
<< pdiffusion >>
rect 89 120 90 121 
<< m1 >>
rect 93 120 94 121 
<< m2 >>
rect 115 120 116 121 
<< m1 >>
rect 116 120 117 121 
<< m1 >>
rect 118 120 119 121 
<< pdiffusion >>
rect 120 120 121 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< pdiffusion >>
rect 138 120 139 121 
<< m1 >>
rect 139 120 140 121 
<< pdiffusion >>
rect 139 120 140 121 
<< pdiffusion >>
rect 140 120 141 121 
<< pdiffusion >>
rect 141 120 142 121 
<< pdiffusion >>
rect 142 120 143 121 
<< pdiffusion >>
rect 143 120 144 121 
<< m1 >>
rect 145 120 146 121 
<< m2 >>
rect 145 120 146 121 
<< pdiffusion >>
rect 156 120 157 121 
<< m1 >>
rect 157 120 158 121 
<< pdiffusion >>
rect 157 120 158 121 
<< pdiffusion >>
rect 158 120 159 121 
<< pdiffusion >>
rect 159 120 160 121 
<< pdiffusion >>
rect 160 120 161 121 
<< pdiffusion >>
rect 161 120 162 121 
<< pdiffusion >>
rect 174 120 175 121 
<< pdiffusion >>
rect 175 120 176 121 
<< pdiffusion >>
rect 176 120 177 121 
<< pdiffusion >>
rect 177 120 178 121 
<< m1 >>
rect 178 120 179 121 
<< pdiffusion >>
rect 178 120 179 121 
<< pdiffusion >>
rect 179 120 180 121 
<< pdiffusion >>
rect 192 120 193 121 
<< m1 >>
rect 193 120 194 121 
<< pdiffusion >>
rect 193 120 194 121 
<< pdiffusion >>
rect 194 120 195 121 
<< pdiffusion >>
rect 195 120 196 121 
<< pdiffusion >>
rect 196 120 197 121 
<< pdiffusion >>
rect 197 120 198 121 
<< m1 >>
rect 199 120 200 121 
<< pdiffusion >>
rect 210 120 211 121 
<< pdiffusion >>
rect 211 120 212 121 
<< pdiffusion >>
rect 212 120 213 121 
<< pdiffusion >>
rect 213 120 214 121 
<< m1 >>
rect 214 120 215 121 
<< pdiffusion >>
rect 214 120 215 121 
<< pdiffusion >>
rect 215 120 216 121 
<< m1 >>
rect 222 120 223 121 
<< m1 >>
rect 223 120 224 121 
<< m1 >>
rect 224 120 225 121 
<< m2 >>
rect 224 120 225 121 
<< m2c >>
rect 224 120 225 121 
<< m1 >>
rect 224 120 225 121 
<< m2 >>
rect 224 120 225 121 
<< m2 >>
rect 225 120 226 121 
<< m1 >>
rect 226 120 227 121 
<< m2 >>
rect 226 120 227 121 
<< pdiffusion >>
rect 228 120 229 121 
<< pdiffusion >>
rect 229 120 230 121 
<< pdiffusion >>
rect 230 120 231 121 
<< pdiffusion >>
rect 231 120 232 121 
<< pdiffusion >>
rect 232 120 233 121 
<< pdiffusion >>
rect 233 120 234 121 
<< m1 >>
rect 262 120 263 121 
<< pdiffusion >>
rect 264 120 265 121 
<< pdiffusion >>
rect 265 120 266 121 
<< pdiffusion >>
rect 266 120 267 121 
<< pdiffusion >>
rect 267 120 268 121 
<< pdiffusion >>
rect 268 120 269 121 
<< pdiffusion >>
rect 269 120 270 121 
<< m1 >>
rect 271 120 272 121 
<< m1 >>
rect 280 120 281 121 
<< pdiffusion >>
rect 282 120 283 121 
<< pdiffusion >>
rect 283 120 284 121 
<< pdiffusion >>
rect 284 120 285 121 
<< pdiffusion >>
rect 285 120 286 121 
<< pdiffusion >>
rect 286 120 287 121 
<< pdiffusion >>
rect 287 120 288 121 
<< m1 >>
rect 298 120 299 121 
<< pdiffusion >>
rect 300 120 301 121 
<< pdiffusion >>
rect 301 120 302 121 
<< pdiffusion >>
rect 302 120 303 121 
<< pdiffusion >>
rect 303 120 304 121 
<< m1 >>
rect 304 120 305 121 
<< pdiffusion >>
rect 304 120 305 121 
<< pdiffusion >>
rect 305 120 306 121 
<< m1 >>
rect 307 120 308 121 
<< m1 >>
rect 319 120 320 121 
<< m1 >>
rect 334 120 335 121 
<< pdiffusion >>
rect 336 120 337 121 
<< m1 >>
rect 337 120 338 121 
<< pdiffusion >>
rect 337 120 338 121 
<< pdiffusion >>
rect 338 120 339 121 
<< pdiffusion >>
rect 339 120 340 121 
<< pdiffusion >>
rect 340 120 341 121 
<< pdiffusion >>
rect 341 120 342 121 
<< pdiffusion >>
rect 354 120 355 121 
<< pdiffusion >>
rect 355 120 356 121 
<< pdiffusion >>
rect 356 120 357 121 
<< pdiffusion >>
rect 357 120 358 121 
<< pdiffusion >>
rect 358 120 359 121 
<< pdiffusion >>
rect 359 120 360 121 
<< pdiffusion >>
rect 372 120 373 121 
<< pdiffusion >>
rect 373 120 374 121 
<< pdiffusion >>
rect 374 120 375 121 
<< pdiffusion >>
rect 375 120 376 121 
<< m1 >>
rect 376 120 377 121 
<< pdiffusion >>
rect 376 120 377 121 
<< pdiffusion >>
rect 377 120 378 121 
<< m1 >>
rect 388 120 389 121 
<< pdiffusion >>
rect 390 120 391 121 
<< pdiffusion >>
rect 391 120 392 121 
<< pdiffusion >>
rect 392 120 393 121 
<< pdiffusion >>
rect 393 120 394 121 
<< pdiffusion >>
rect 394 120 395 121 
<< pdiffusion >>
rect 395 120 396 121 
<< pdiffusion >>
rect 408 120 409 121 
<< pdiffusion >>
rect 409 120 410 121 
<< pdiffusion >>
rect 410 120 411 121 
<< pdiffusion >>
rect 411 120 412 121 
<< m1 >>
rect 412 120 413 121 
<< pdiffusion >>
rect 412 120 413 121 
<< pdiffusion >>
rect 413 120 414 121 
<< pdiffusion >>
rect 426 120 427 121 
<< pdiffusion >>
rect 427 120 428 121 
<< pdiffusion >>
rect 428 120 429 121 
<< pdiffusion >>
rect 429 120 430 121 
<< pdiffusion >>
rect 430 120 431 121 
<< pdiffusion >>
rect 431 120 432 121 
<< pdiffusion >>
rect 444 120 445 121 
<< pdiffusion >>
rect 445 120 446 121 
<< pdiffusion >>
rect 446 120 447 121 
<< pdiffusion >>
rect 447 120 448 121 
<< pdiffusion >>
rect 448 120 449 121 
<< pdiffusion >>
rect 449 120 450 121 
<< m1 >>
rect 451 120 452 121 
<< pdiffusion >>
rect 12 121 13 122 
<< pdiffusion >>
rect 13 121 14 122 
<< pdiffusion >>
rect 14 121 15 122 
<< pdiffusion >>
rect 15 121 16 122 
<< pdiffusion >>
rect 16 121 17 122 
<< pdiffusion >>
rect 17 121 18 122 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< pdiffusion >>
rect 48 121 49 122 
<< pdiffusion >>
rect 49 121 50 122 
<< pdiffusion >>
rect 50 121 51 122 
<< pdiffusion >>
rect 51 121 52 122 
<< pdiffusion >>
rect 52 121 53 122 
<< pdiffusion >>
rect 53 121 54 122 
<< m1 >>
rect 62 121 63 122 
<< m1 >>
rect 64 121 65 122 
<< pdiffusion >>
rect 66 121 67 122 
<< pdiffusion >>
rect 67 121 68 122 
<< pdiffusion >>
rect 68 121 69 122 
<< pdiffusion >>
rect 69 121 70 122 
<< pdiffusion >>
rect 70 121 71 122 
<< pdiffusion >>
rect 71 121 72 122 
<< m1 >>
rect 73 121 74 122 
<< pdiffusion >>
rect 84 121 85 122 
<< pdiffusion >>
rect 85 121 86 122 
<< pdiffusion >>
rect 86 121 87 122 
<< pdiffusion >>
rect 87 121 88 122 
<< pdiffusion >>
rect 88 121 89 122 
<< pdiffusion >>
rect 89 121 90 122 
<< m1 >>
rect 93 121 94 122 
<< m2 >>
rect 115 121 116 122 
<< m1 >>
rect 116 121 117 122 
<< m1 >>
rect 118 121 119 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< pdiffusion >>
rect 138 121 139 122 
<< pdiffusion >>
rect 139 121 140 122 
<< pdiffusion >>
rect 140 121 141 122 
<< pdiffusion >>
rect 141 121 142 122 
<< pdiffusion >>
rect 142 121 143 122 
<< pdiffusion >>
rect 143 121 144 122 
<< m1 >>
rect 145 121 146 122 
<< m2 >>
rect 145 121 146 122 
<< pdiffusion >>
rect 156 121 157 122 
<< pdiffusion >>
rect 157 121 158 122 
<< pdiffusion >>
rect 158 121 159 122 
<< pdiffusion >>
rect 159 121 160 122 
<< pdiffusion >>
rect 160 121 161 122 
<< pdiffusion >>
rect 161 121 162 122 
<< pdiffusion >>
rect 174 121 175 122 
<< pdiffusion >>
rect 175 121 176 122 
<< pdiffusion >>
rect 176 121 177 122 
<< pdiffusion >>
rect 177 121 178 122 
<< pdiffusion >>
rect 178 121 179 122 
<< pdiffusion >>
rect 179 121 180 122 
<< pdiffusion >>
rect 192 121 193 122 
<< pdiffusion >>
rect 193 121 194 122 
<< pdiffusion >>
rect 194 121 195 122 
<< pdiffusion >>
rect 195 121 196 122 
<< pdiffusion >>
rect 196 121 197 122 
<< pdiffusion >>
rect 197 121 198 122 
<< m1 >>
rect 199 121 200 122 
<< pdiffusion >>
rect 210 121 211 122 
<< pdiffusion >>
rect 211 121 212 122 
<< pdiffusion >>
rect 212 121 213 122 
<< pdiffusion >>
rect 213 121 214 122 
<< pdiffusion >>
rect 214 121 215 122 
<< pdiffusion >>
rect 215 121 216 122 
<< m1 >>
rect 222 121 223 122 
<< m1 >>
rect 226 121 227 122 
<< pdiffusion >>
rect 228 121 229 122 
<< pdiffusion >>
rect 229 121 230 122 
<< pdiffusion >>
rect 230 121 231 122 
<< pdiffusion >>
rect 231 121 232 122 
<< pdiffusion >>
rect 232 121 233 122 
<< pdiffusion >>
rect 233 121 234 122 
<< m1 >>
rect 262 121 263 122 
<< pdiffusion >>
rect 264 121 265 122 
<< pdiffusion >>
rect 265 121 266 122 
<< pdiffusion >>
rect 266 121 267 122 
<< pdiffusion >>
rect 267 121 268 122 
<< pdiffusion >>
rect 268 121 269 122 
<< pdiffusion >>
rect 269 121 270 122 
<< m1 >>
rect 271 121 272 122 
<< m1 >>
rect 280 121 281 122 
<< pdiffusion >>
rect 282 121 283 122 
<< pdiffusion >>
rect 283 121 284 122 
<< pdiffusion >>
rect 284 121 285 122 
<< pdiffusion >>
rect 285 121 286 122 
<< pdiffusion >>
rect 286 121 287 122 
<< pdiffusion >>
rect 287 121 288 122 
<< m1 >>
rect 298 121 299 122 
<< pdiffusion >>
rect 300 121 301 122 
<< pdiffusion >>
rect 301 121 302 122 
<< pdiffusion >>
rect 302 121 303 122 
<< pdiffusion >>
rect 303 121 304 122 
<< pdiffusion >>
rect 304 121 305 122 
<< pdiffusion >>
rect 305 121 306 122 
<< m1 >>
rect 307 121 308 122 
<< m1 >>
rect 319 121 320 122 
<< m1 >>
rect 334 121 335 122 
<< pdiffusion >>
rect 336 121 337 122 
<< pdiffusion >>
rect 337 121 338 122 
<< pdiffusion >>
rect 338 121 339 122 
<< pdiffusion >>
rect 339 121 340 122 
<< pdiffusion >>
rect 340 121 341 122 
<< pdiffusion >>
rect 341 121 342 122 
<< pdiffusion >>
rect 354 121 355 122 
<< pdiffusion >>
rect 355 121 356 122 
<< pdiffusion >>
rect 356 121 357 122 
<< pdiffusion >>
rect 357 121 358 122 
<< pdiffusion >>
rect 358 121 359 122 
<< pdiffusion >>
rect 359 121 360 122 
<< pdiffusion >>
rect 372 121 373 122 
<< pdiffusion >>
rect 373 121 374 122 
<< pdiffusion >>
rect 374 121 375 122 
<< pdiffusion >>
rect 375 121 376 122 
<< pdiffusion >>
rect 376 121 377 122 
<< pdiffusion >>
rect 377 121 378 122 
<< m1 >>
rect 388 121 389 122 
<< pdiffusion >>
rect 390 121 391 122 
<< pdiffusion >>
rect 391 121 392 122 
<< pdiffusion >>
rect 392 121 393 122 
<< pdiffusion >>
rect 393 121 394 122 
<< pdiffusion >>
rect 394 121 395 122 
<< pdiffusion >>
rect 395 121 396 122 
<< pdiffusion >>
rect 408 121 409 122 
<< pdiffusion >>
rect 409 121 410 122 
<< pdiffusion >>
rect 410 121 411 122 
<< pdiffusion >>
rect 411 121 412 122 
<< pdiffusion >>
rect 412 121 413 122 
<< pdiffusion >>
rect 413 121 414 122 
<< pdiffusion >>
rect 426 121 427 122 
<< pdiffusion >>
rect 427 121 428 122 
<< pdiffusion >>
rect 428 121 429 122 
<< pdiffusion >>
rect 429 121 430 122 
<< pdiffusion >>
rect 430 121 431 122 
<< pdiffusion >>
rect 431 121 432 122 
<< pdiffusion >>
rect 444 121 445 122 
<< pdiffusion >>
rect 445 121 446 122 
<< pdiffusion >>
rect 446 121 447 122 
<< pdiffusion >>
rect 447 121 448 122 
<< pdiffusion >>
rect 448 121 449 122 
<< pdiffusion >>
rect 449 121 450 122 
<< m1 >>
rect 451 121 452 122 
<< pdiffusion >>
rect 12 122 13 123 
<< pdiffusion >>
rect 13 122 14 123 
<< pdiffusion >>
rect 14 122 15 123 
<< pdiffusion >>
rect 15 122 16 123 
<< pdiffusion >>
rect 16 122 17 123 
<< pdiffusion >>
rect 17 122 18 123 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< pdiffusion >>
rect 48 122 49 123 
<< pdiffusion >>
rect 49 122 50 123 
<< pdiffusion >>
rect 50 122 51 123 
<< pdiffusion >>
rect 51 122 52 123 
<< pdiffusion >>
rect 52 122 53 123 
<< pdiffusion >>
rect 53 122 54 123 
<< m1 >>
rect 62 122 63 123 
<< m1 >>
rect 64 122 65 123 
<< pdiffusion >>
rect 66 122 67 123 
<< pdiffusion >>
rect 67 122 68 123 
<< pdiffusion >>
rect 68 122 69 123 
<< pdiffusion >>
rect 69 122 70 123 
<< pdiffusion >>
rect 70 122 71 123 
<< pdiffusion >>
rect 71 122 72 123 
<< m1 >>
rect 73 122 74 123 
<< pdiffusion >>
rect 84 122 85 123 
<< pdiffusion >>
rect 85 122 86 123 
<< pdiffusion >>
rect 86 122 87 123 
<< pdiffusion >>
rect 87 122 88 123 
<< pdiffusion >>
rect 88 122 89 123 
<< pdiffusion >>
rect 89 122 90 123 
<< m1 >>
rect 93 122 94 123 
<< m2 >>
rect 115 122 116 123 
<< m1 >>
rect 116 122 117 123 
<< m1 >>
rect 118 122 119 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< pdiffusion >>
rect 138 122 139 123 
<< pdiffusion >>
rect 139 122 140 123 
<< pdiffusion >>
rect 140 122 141 123 
<< pdiffusion >>
rect 141 122 142 123 
<< pdiffusion >>
rect 142 122 143 123 
<< pdiffusion >>
rect 143 122 144 123 
<< m1 >>
rect 145 122 146 123 
<< m2 >>
rect 145 122 146 123 
<< pdiffusion >>
rect 156 122 157 123 
<< pdiffusion >>
rect 157 122 158 123 
<< pdiffusion >>
rect 158 122 159 123 
<< pdiffusion >>
rect 159 122 160 123 
<< pdiffusion >>
rect 160 122 161 123 
<< pdiffusion >>
rect 161 122 162 123 
<< pdiffusion >>
rect 174 122 175 123 
<< pdiffusion >>
rect 175 122 176 123 
<< pdiffusion >>
rect 176 122 177 123 
<< pdiffusion >>
rect 177 122 178 123 
<< pdiffusion >>
rect 178 122 179 123 
<< pdiffusion >>
rect 179 122 180 123 
<< pdiffusion >>
rect 192 122 193 123 
<< pdiffusion >>
rect 193 122 194 123 
<< pdiffusion >>
rect 194 122 195 123 
<< pdiffusion >>
rect 195 122 196 123 
<< pdiffusion >>
rect 196 122 197 123 
<< pdiffusion >>
rect 197 122 198 123 
<< m1 >>
rect 199 122 200 123 
<< pdiffusion >>
rect 210 122 211 123 
<< pdiffusion >>
rect 211 122 212 123 
<< pdiffusion >>
rect 212 122 213 123 
<< pdiffusion >>
rect 213 122 214 123 
<< pdiffusion >>
rect 214 122 215 123 
<< pdiffusion >>
rect 215 122 216 123 
<< m1 >>
rect 222 122 223 123 
<< m1 >>
rect 226 122 227 123 
<< pdiffusion >>
rect 228 122 229 123 
<< pdiffusion >>
rect 229 122 230 123 
<< pdiffusion >>
rect 230 122 231 123 
<< pdiffusion >>
rect 231 122 232 123 
<< pdiffusion >>
rect 232 122 233 123 
<< pdiffusion >>
rect 233 122 234 123 
<< m1 >>
rect 262 122 263 123 
<< pdiffusion >>
rect 264 122 265 123 
<< pdiffusion >>
rect 265 122 266 123 
<< pdiffusion >>
rect 266 122 267 123 
<< pdiffusion >>
rect 267 122 268 123 
<< pdiffusion >>
rect 268 122 269 123 
<< pdiffusion >>
rect 269 122 270 123 
<< m1 >>
rect 271 122 272 123 
<< m1 >>
rect 280 122 281 123 
<< pdiffusion >>
rect 282 122 283 123 
<< pdiffusion >>
rect 283 122 284 123 
<< pdiffusion >>
rect 284 122 285 123 
<< pdiffusion >>
rect 285 122 286 123 
<< pdiffusion >>
rect 286 122 287 123 
<< pdiffusion >>
rect 287 122 288 123 
<< m1 >>
rect 298 122 299 123 
<< pdiffusion >>
rect 300 122 301 123 
<< pdiffusion >>
rect 301 122 302 123 
<< pdiffusion >>
rect 302 122 303 123 
<< pdiffusion >>
rect 303 122 304 123 
<< pdiffusion >>
rect 304 122 305 123 
<< pdiffusion >>
rect 305 122 306 123 
<< m1 >>
rect 307 122 308 123 
<< m1 >>
rect 319 122 320 123 
<< m1 >>
rect 334 122 335 123 
<< pdiffusion >>
rect 336 122 337 123 
<< pdiffusion >>
rect 337 122 338 123 
<< pdiffusion >>
rect 338 122 339 123 
<< pdiffusion >>
rect 339 122 340 123 
<< pdiffusion >>
rect 340 122 341 123 
<< pdiffusion >>
rect 341 122 342 123 
<< pdiffusion >>
rect 354 122 355 123 
<< pdiffusion >>
rect 355 122 356 123 
<< pdiffusion >>
rect 356 122 357 123 
<< pdiffusion >>
rect 357 122 358 123 
<< pdiffusion >>
rect 358 122 359 123 
<< pdiffusion >>
rect 359 122 360 123 
<< pdiffusion >>
rect 372 122 373 123 
<< pdiffusion >>
rect 373 122 374 123 
<< pdiffusion >>
rect 374 122 375 123 
<< pdiffusion >>
rect 375 122 376 123 
<< pdiffusion >>
rect 376 122 377 123 
<< pdiffusion >>
rect 377 122 378 123 
<< m1 >>
rect 388 122 389 123 
<< pdiffusion >>
rect 390 122 391 123 
<< pdiffusion >>
rect 391 122 392 123 
<< pdiffusion >>
rect 392 122 393 123 
<< pdiffusion >>
rect 393 122 394 123 
<< pdiffusion >>
rect 394 122 395 123 
<< pdiffusion >>
rect 395 122 396 123 
<< pdiffusion >>
rect 408 122 409 123 
<< pdiffusion >>
rect 409 122 410 123 
<< pdiffusion >>
rect 410 122 411 123 
<< pdiffusion >>
rect 411 122 412 123 
<< pdiffusion >>
rect 412 122 413 123 
<< pdiffusion >>
rect 413 122 414 123 
<< pdiffusion >>
rect 426 122 427 123 
<< pdiffusion >>
rect 427 122 428 123 
<< pdiffusion >>
rect 428 122 429 123 
<< pdiffusion >>
rect 429 122 430 123 
<< pdiffusion >>
rect 430 122 431 123 
<< pdiffusion >>
rect 431 122 432 123 
<< pdiffusion >>
rect 444 122 445 123 
<< pdiffusion >>
rect 445 122 446 123 
<< pdiffusion >>
rect 446 122 447 123 
<< pdiffusion >>
rect 447 122 448 123 
<< pdiffusion >>
rect 448 122 449 123 
<< pdiffusion >>
rect 449 122 450 123 
<< m1 >>
rect 451 122 452 123 
<< pdiffusion >>
rect 12 123 13 124 
<< pdiffusion >>
rect 13 123 14 124 
<< pdiffusion >>
rect 14 123 15 124 
<< pdiffusion >>
rect 15 123 16 124 
<< pdiffusion >>
rect 16 123 17 124 
<< pdiffusion >>
rect 17 123 18 124 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< pdiffusion >>
rect 48 123 49 124 
<< pdiffusion >>
rect 49 123 50 124 
<< pdiffusion >>
rect 50 123 51 124 
<< pdiffusion >>
rect 51 123 52 124 
<< pdiffusion >>
rect 52 123 53 124 
<< pdiffusion >>
rect 53 123 54 124 
<< m1 >>
rect 62 123 63 124 
<< m1 >>
rect 64 123 65 124 
<< pdiffusion >>
rect 66 123 67 124 
<< pdiffusion >>
rect 67 123 68 124 
<< pdiffusion >>
rect 68 123 69 124 
<< pdiffusion >>
rect 69 123 70 124 
<< pdiffusion >>
rect 70 123 71 124 
<< pdiffusion >>
rect 71 123 72 124 
<< m1 >>
rect 73 123 74 124 
<< pdiffusion >>
rect 84 123 85 124 
<< pdiffusion >>
rect 85 123 86 124 
<< pdiffusion >>
rect 86 123 87 124 
<< pdiffusion >>
rect 87 123 88 124 
<< pdiffusion >>
rect 88 123 89 124 
<< pdiffusion >>
rect 89 123 90 124 
<< m1 >>
rect 93 123 94 124 
<< m2 >>
rect 115 123 116 124 
<< m1 >>
rect 116 123 117 124 
<< m1 >>
rect 118 123 119 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< pdiffusion >>
rect 138 123 139 124 
<< pdiffusion >>
rect 139 123 140 124 
<< pdiffusion >>
rect 140 123 141 124 
<< pdiffusion >>
rect 141 123 142 124 
<< pdiffusion >>
rect 142 123 143 124 
<< pdiffusion >>
rect 143 123 144 124 
<< m1 >>
rect 145 123 146 124 
<< m2 >>
rect 145 123 146 124 
<< pdiffusion >>
rect 156 123 157 124 
<< pdiffusion >>
rect 157 123 158 124 
<< pdiffusion >>
rect 158 123 159 124 
<< pdiffusion >>
rect 159 123 160 124 
<< pdiffusion >>
rect 160 123 161 124 
<< pdiffusion >>
rect 161 123 162 124 
<< pdiffusion >>
rect 174 123 175 124 
<< pdiffusion >>
rect 175 123 176 124 
<< pdiffusion >>
rect 176 123 177 124 
<< pdiffusion >>
rect 177 123 178 124 
<< pdiffusion >>
rect 178 123 179 124 
<< pdiffusion >>
rect 179 123 180 124 
<< pdiffusion >>
rect 192 123 193 124 
<< pdiffusion >>
rect 193 123 194 124 
<< pdiffusion >>
rect 194 123 195 124 
<< pdiffusion >>
rect 195 123 196 124 
<< pdiffusion >>
rect 196 123 197 124 
<< pdiffusion >>
rect 197 123 198 124 
<< m1 >>
rect 199 123 200 124 
<< pdiffusion >>
rect 210 123 211 124 
<< pdiffusion >>
rect 211 123 212 124 
<< pdiffusion >>
rect 212 123 213 124 
<< pdiffusion >>
rect 213 123 214 124 
<< pdiffusion >>
rect 214 123 215 124 
<< pdiffusion >>
rect 215 123 216 124 
<< m1 >>
rect 222 123 223 124 
<< m1 >>
rect 226 123 227 124 
<< pdiffusion >>
rect 228 123 229 124 
<< pdiffusion >>
rect 229 123 230 124 
<< pdiffusion >>
rect 230 123 231 124 
<< pdiffusion >>
rect 231 123 232 124 
<< pdiffusion >>
rect 232 123 233 124 
<< pdiffusion >>
rect 233 123 234 124 
<< m1 >>
rect 262 123 263 124 
<< pdiffusion >>
rect 264 123 265 124 
<< pdiffusion >>
rect 265 123 266 124 
<< pdiffusion >>
rect 266 123 267 124 
<< pdiffusion >>
rect 267 123 268 124 
<< pdiffusion >>
rect 268 123 269 124 
<< pdiffusion >>
rect 269 123 270 124 
<< m1 >>
rect 271 123 272 124 
<< m1 >>
rect 280 123 281 124 
<< pdiffusion >>
rect 282 123 283 124 
<< pdiffusion >>
rect 283 123 284 124 
<< pdiffusion >>
rect 284 123 285 124 
<< pdiffusion >>
rect 285 123 286 124 
<< pdiffusion >>
rect 286 123 287 124 
<< pdiffusion >>
rect 287 123 288 124 
<< m1 >>
rect 298 123 299 124 
<< pdiffusion >>
rect 300 123 301 124 
<< pdiffusion >>
rect 301 123 302 124 
<< pdiffusion >>
rect 302 123 303 124 
<< pdiffusion >>
rect 303 123 304 124 
<< pdiffusion >>
rect 304 123 305 124 
<< pdiffusion >>
rect 305 123 306 124 
<< m1 >>
rect 307 123 308 124 
<< m1 >>
rect 319 123 320 124 
<< m1 >>
rect 334 123 335 124 
<< pdiffusion >>
rect 336 123 337 124 
<< pdiffusion >>
rect 337 123 338 124 
<< pdiffusion >>
rect 338 123 339 124 
<< pdiffusion >>
rect 339 123 340 124 
<< pdiffusion >>
rect 340 123 341 124 
<< pdiffusion >>
rect 341 123 342 124 
<< pdiffusion >>
rect 354 123 355 124 
<< pdiffusion >>
rect 355 123 356 124 
<< pdiffusion >>
rect 356 123 357 124 
<< pdiffusion >>
rect 357 123 358 124 
<< pdiffusion >>
rect 358 123 359 124 
<< pdiffusion >>
rect 359 123 360 124 
<< pdiffusion >>
rect 372 123 373 124 
<< pdiffusion >>
rect 373 123 374 124 
<< pdiffusion >>
rect 374 123 375 124 
<< pdiffusion >>
rect 375 123 376 124 
<< pdiffusion >>
rect 376 123 377 124 
<< pdiffusion >>
rect 377 123 378 124 
<< m1 >>
rect 388 123 389 124 
<< pdiffusion >>
rect 390 123 391 124 
<< pdiffusion >>
rect 391 123 392 124 
<< pdiffusion >>
rect 392 123 393 124 
<< pdiffusion >>
rect 393 123 394 124 
<< pdiffusion >>
rect 394 123 395 124 
<< pdiffusion >>
rect 395 123 396 124 
<< pdiffusion >>
rect 408 123 409 124 
<< pdiffusion >>
rect 409 123 410 124 
<< pdiffusion >>
rect 410 123 411 124 
<< pdiffusion >>
rect 411 123 412 124 
<< pdiffusion >>
rect 412 123 413 124 
<< pdiffusion >>
rect 413 123 414 124 
<< pdiffusion >>
rect 426 123 427 124 
<< pdiffusion >>
rect 427 123 428 124 
<< pdiffusion >>
rect 428 123 429 124 
<< pdiffusion >>
rect 429 123 430 124 
<< pdiffusion >>
rect 430 123 431 124 
<< pdiffusion >>
rect 431 123 432 124 
<< pdiffusion >>
rect 444 123 445 124 
<< pdiffusion >>
rect 445 123 446 124 
<< pdiffusion >>
rect 446 123 447 124 
<< pdiffusion >>
rect 447 123 448 124 
<< pdiffusion >>
rect 448 123 449 124 
<< pdiffusion >>
rect 449 123 450 124 
<< m1 >>
rect 451 123 452 124 
<< pdiffusion >>
rect 12 124 13 125 
<< pdiffusion >>
rect 13 124 14 125 
<< pdiffusion >>
rect 14 124 15 125 
<< pdiffusion >>
rect 15 124 16 125 
<< pdiffusion >>
rect 16 124 17 125 
<< pdiffusion >>
rect 17 124 18 125 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< pdiffusion >>
rect 48 124 49 125 
<< pdiffusion >>
rect 49 124 50 125 
<< pdiffusion >>
rect 50 124 51 125 
<< pdiffusion >>
rect 51 124 52 125 
<< pdiffusion >>
rect 52 124 53 125 
<< pdiffusion >>
rect 53 124 54 125 
<< m1 >>
rect 62 124 63 125 
<< m1 >>
rect 64 124 65 125 
<< pdiffusion >>
rect 66 124 67 125 
<< pdiffusion >>
rect 67 124 68 125 
<< pdiffusion >>
rect 68 124 69 125 
<< pdiffusion >>
rect 69 124 70 125 
<< pdiffusion >>
rect 70 124 71 125 
<< pdiffusion >>
rect 71 124 72 125 
<< m1 >>
rect 73 124 74 125 
<< pdiffusion >>
rect 84 124 85 125 
<< pdiffusion >>
rect 85 124 86 125 
<< pdiffusion >>
rect 86 124 87 125 
<< pdiffusion >>
rect 87 124 88 125 
<< pdiffusion >>
rect 88 124 89 125 
<< pdiffusion >>
rect 89 124 90 125 
<< m1 >>
rect 93 124 94 125 
<< m2 >>
rect 115 124 116 125 
<< m1 >>
rect 116 124 117 125 
<< m1 >>
rect 118 124 119 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< pdiffusion >>
rect 138 124 139 125 
<< pdiffusion >>
rect 139 124 140 125 
<< pdiffusion >>
rect 140 124 141 125 
<< pdiffusion >>
rect 141 124 142 125 
<< pdiffusion >>
rect 142 124 143 125 
<< pdiffusion >>
rect 143 124 144 125 
<< m1 >>
rect 145 124 146 125 
<< m2 >>
rect 145 124 146 125 
<< pdiffusion >>
rect 156 124 157 125 
<< pdiffusion >>
rect 157 124 158 125 
<< pdiffusion >>
rect 158 124 159 125 
<< pdiffusion >>
rect 159 124 160 125 
<< pdiffusion >>
rect 160 124 161 125 
<< pdiffusion >>
rect 161 124 162 125 
<< pdiffusion >>
rect 174 124 175 125 
<< pdiffusion >>
rect 175 124 176 125 
<< pdiffusion >>
rect 176 124 177 125 
<< pdiffusion >>
rect 177 124 178 125 
<< pdiffusion >>
rect 178 124 179 125 
<< pdiffusion >>
rect 179 124 180 125 
<< pdiffusion >>
rect 192 124 193 125 
<< pdiffusion >>
rect 193 124 194 125 
<< pdiffusion >>
rect 194 124 195 125 
<< pdiffusion >>
rect 195 124 196 125 
<< pdiffusion >>
rect 196 124 197 125 
<< pdiffusion >>
rect 197 124 198 125 
<< m1 >>
rect 199 124 200 125 
<< pdiffusion >>
rect 210 124 211 125 
<< pdiffusion >>
rect 211 124 212 125 
<< pdiffusion >>
rect 212 124 213 125 
<< pdiffusion >>
rect 213 124 214 125 
<< pdiffusion >>
rect 214 124 215 125 
<< pdiffusion >>
rect 215 124 216 125 
<< m1 >>
rect 222 124 223 125 
<< m1 >>
rect 226 124 227 125 
<< pdiffusion >>
rect 228 124 229 125 
<< pdiffusion >>
rect 229 124 230 125 
<< pdiffusion >>
rect 230 124 231 125 
<< pdiffusion >>
rect 231 124 232 125 
<< pdiffusion >>
rect 232 124 233 125 
<< pdiffusion >>
rect 233 124 234 125 
<< m1 >>
rect 262 124 263 125 
<< pdiffusion >>
rect 264 124 265 125 
<< pdiffusion >>
rect 265 124 266 125 
<< pdiffusion >>
rect 266 124 267 125 
<< pdiffusion >>
rect 267 124 268 125 
<< pdiffusion >>
rect 268 124 269 125 
<< pdiffusion >>
rect 269 124 270 125 
<< m1 >>
rect 271 124 272 125 
<< m1 >>
rect 280 124 281 125 
<< pdiffusion >>
rect 282 124 283 125 
<< pdiffusion >>
rect 283 124 284 125 
<< pdiffusion >>
rect 284 124 285 125 
<< pdiffusion >>
rect 285 124 286 125 
<< pdiffusion >>
rect 286 124 287 125 
<< pdiffusion >>
rect 287 124 288 125 
<< m1 >>
rect 298 124 299 125 
<< pdiffusion >>
rect 300 124 301 125 
<< pdiffusion >>
rect 301 124 302 125 
<< pdiffusion >>
rect 302 124 303 125 
<< pdiffusion >>
rect 303 124 304 125 
<< pdiffusion >>
rect 304 124 305 125 
<< pdiffusion >>
rect 305 124 306 125 
<< m1 >>
rect 307 124 308 125 
<< m1 >>
rect 319 124 320 125 
<< m1 >>
rect 334 124 335 125 
<< pdiffusion >>
rect 336 124 337 125 
<< pdiffusion >>
rect 337 124 338 125 
<< pdiffusion >>
rect 338 124 339 125 
<< pdiffusion >>
rect 339 124 340 125 
<< pdiffusion >>
rect 340 124 341 125 
<< pdiffusion >>
rect 341 124 342 125 
<< pdiffusion >>
rect 354 124 355 125 
<< pdiffusion >>
rect 355 124 356 125 
<< pdiffusion >>
rect 356 124 357 125 
<< pdiffusion >>
rect 357 124 358 125 
<< pdiffusion >>
rect 358 124 359 125 
<< pdiffusion >>
rect 359 124 360 125 
<< pdiffusion >>
rect 372 124 373 125 
<< pdiffusion >>
rect 373 124 374 125 
<< pdiffusion >>
rect 374 124 375 125 
<< pdiffusion >>
rect 375 124 376 125 
<< pdiffusion >>
rect 376 124 377 125 
<< pdiffusion >>
rect 377 124 378 125 
<< m1 >>
rect 388 124 389 125 
<< pdiffusion >>
rect 390 124 391 125 
<< pdiffusion >>
rect 391 124 392 125 
<< pdiffusion >>
rect 392 124 393 125 
<< pdiffusion >>
rect 393 124 394 125 
<< pdiffusion >>
rect 394 124 395 125 
<< pdiffusion >>
rect 395 124 396 125 
<< pdiffusion >>
rect 408 124 409 125 
<< pdiffusion >>
rect 409 124 410 125 
<< pdiffusion >>
rect 410 124 411 125 
<< pdiffusion >>
rect 411 124 412 125 
<< pdiffusion >>
rect 412 124 413 125 
<< pdiffusion >>
rect 413 124 414 125 
<< pdiffusion >>
rect 426 124 427 125 
<< pdiffusion >>
rect 427 124 428 125 
<< pdiffusion >>
rect 428 124 429 125 
<< pdiffusion >>
rect 429 124 430 125 
<< pdiffusion >>
rect 430 124 431 125 
<< pdiffusion >>
rect 431 124 432 125 
<< pdiffusion >>
rect 444 124 445 125 
<< pdiffusion >>
rect 445 124 446 125 
<< pdiffusion >>
rect 446 124 447 125 
<< pdiffusion >>
rect 447 124 448 125 
<< pdiffusion >>
rect 448 124 449 125 
<< pdiffusion >>
rect 449 124 450 125 
<< m1 >>
rect 451 124 452 125 
<< pdiffusion >>
rect 12 125 13 126 
<< pdiffusion >>
rect 13 125 14 126 
<< pdiffusion >>
rect 14 125 15 126 
<< pdiffusion >>
rect 15 125 16 126 
<< pdiffusion >>
rect 16 125 17 126 
<< pdiffusion >>
rect 17 125 18 126 
<< pdiffusion >>
rect 30 125 31 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< pdiffusion >>
rect 48 125 49 126 
<< pdiffusion >>
rect 49 125 50 126 
<< pdiffusion >>
rect 50 125 51 126 
<< pdiffusion >>
rect 51 125 52 126 
<< pdiffusion >>
rect 52 125 53 126 
<< pdiffusion >>
rect 53 125 54 126 
<< m1 >>
rect 62 125 63 126 
<< m1 >>
rect 64 125 65 126 
<< pdiffusion >>
rect 66 125 67 126 
<< m1 >>
rect 67 125 68 126 
<< pdiffusion >>
rect 67 125 68 126 
<< pdiffusion >>
rect 68 125 69 126 
<< pdiffusion >>
rect 69 125 70 126 
<< pdiffusion >>
rect 70 125 71 126 
<< pdiffusion >>
rect 71 125 72 126 
<< m1 >>
rect 73 125 74 126 
<< pdiffusion >>
rect 84 125 85 126 
<< pdiffusion >>
rect 85 125 86 126 
<< pdiffusion >>
rect 86 125 87 126 
<< pdiffusion >>
rect 87 125 88 126 
<< pdiffusion >>
rect 88 125 89 126 
<< pdiffusion >>
rect 89 125 90 126 
<< m1 >>
rect 93 125 94 126 
<< m2 >>
rect 115 125 116 126 
<< m1 >>
rect 116 125 117 126 
<< m1 >>
rect 118 125 119 126 
<< pdiffusion >>
rect 120 125 121 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< m1 >>
rect 124 125 125 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< pdiffusion >>
rect 138 125 139 126 
<< pdiffusion >>
rect 139 125 140 126 
<< pdiffusion >>
rect 140 125 141 126 
<< pdiffusion >>
rect 141 125 142 126 
<< m1 >>
rect 142 125 143 126 
<< pdiffusion >>
rect 142 125 143 126 
<< pdiffusion >>
rect 143 125 144 126 
<< m1 >>
rect 145 125 146 126 
<< m2 >>
rect 145 125 146 126 
<< pdiffusion >>
rect 156 125 157 126 
<< pdiffusion >>
rect 157 125 158 126 
<< pdiffusion >>
rect 158 125 159 126 
<< pdiffusion >>
rect 159 125 160 126 
<< pdiffusion >>
rect 160 125 161 126 
<< pdiffusion >>
rect 161 125 162 126 
<< pdiffusion >>
rect 174 125 175 126 
<< pdiffusion >>
rect 175 125 176 126 
<< pdiffusion >>
rect 176 125 177 126 
<< pdiffusion >>
rect 177 125 178 126 
<< m1 >>
rect 178 125 179 126 
<< pdiffusion >>
rect 178 125 179 126 
<< pdiffusion >>
rect 179 125 180 126 
<< pdiffusion >>
rect 192 125 193 126 
<< m1 >>
rect 193 125 194 126 
<< pdiffusion >>
rect 193 125 194 126 
<< pdiffusion >>
rect 194 125 195 126 
<< pdiffusion >>
rect 195 125 196 126 
<< pdiffusion >>
rect 196 125 197 126 
<< pdiffusion >>
rect 197 125 198 126 
<< m1 >>
rect 199 125 200 126 
<< pdiffusion >>
rect 210 125 211 126 
<< pdiffusion >>
rect 211 125 212 126 
<< pdiffusion >>
rect 212 125 213 126 
<< pdiffusion >>
rect 213 125 214 126 
<< m1 >>
rect 214 125 215 126 
<< pdiffusion >>
rect 214 125 215 126 
<< pdiffusion >>
rect 215 125 216 126 
<< m1 >>
rect 222 125 223 126 
<< m1 >>
rect 226 125 227 126 
<< pdiffusion >>
rect 228 125 229 126 
<< pdiffusion >>
rect 229 125 230 126 
<< pdiffusion >>
rect 230 125 231 126 
<< pdiffusion >>
rect 231 125 232 126 
<< pdiffusion >>
rect 232 125 233 126 
<< pdiffusion >>
rect 233 125 234 126 
<< m1 >>
rect 262 125 263 126 
<< pdiffusion >>
rect 264 125 265 126 
<< pdiffusion >>
rect 265 125 266 126 
<< pdiffusion >>
rect 266 125 267 126 
<< pdiffusion >>
rect 267 125 268 126 
<< pdiffusion >>
rect 268 125 269 126 
<< pdiffusion >>
rect 269 125 270 126 
<< m1 >>
rect 271 125 272 126 
<< m1 >>
rect 280 125 281 126 
<< m2 >>
rect 280 125 281 126 
<< m2c >>
rect 280 125 281 126 
<< m1 >>
rect 280 125 281 126 
<< m2 >>
rect 280 125 281 126 
<< pdiffusion >>
rect 282 125 283 126 
<< m1 >>
rect 283 125 284 126 
<< pdiffusion >>
rect 283 125 284 126 
<< pdiffusion >>
rect 284 125 285 126 
<< pdiffusion >>
rect 285 125 286 126 
<< m1 >>
rect 286 125 287 126 
<< pdiffusion >>
rect 286 125 287 126 
<< pdiffusion >>
rect 287 125 288 126 
<< m1 >>
rect 298 125 299 126 
<< pdiffusion >>
rect 300 125 301 126 
<< pdiffusion >>
rect 301 125 302 126 
<< pdiffusion >>
rect 302 125 303 126 
<< pdiffusion >>
rect 303 125 304 126 
<< pdiffusion >>
rect 304 125 305 126 
<< pdiffusion >>
rect 305 125 306 126 
<< m1 >>
rect 307 125 308 126 
<< m1 >>
rect 319 125 320 126 
<< m1 >>
rect 334 125 335 126 
<< pdiffusion >>
rect 336 125 337 126 
<< pdiffusion >>
rect 337 125 338 126 
<< pdiffusion >>
rect 338 125 339 126 
<< pdiffusion >>
rect 339 125 340 126 
<< pdiffusion >>
rect 340 125 341 126 
<< pdiffusion >>
rect 341 125 342 126 
<< pdiffusion >>
rect 354 125 355 126 
<< pdiffusion >>
rect 355 125 356 126 
<< pdiffusion >>
rect 356 125 357 126 
<< pdiffusion >>
rect 357 125 358 126 
<< pdiffusion >>
rect 358 125 359 126 
<< pdiffusion >>
rect 359 125 360 126 
<< pdiffusion >>
rect 372 125 373 126 
<< pdiffusion >>
rect 373 125 374 126 
<< pdiffusion >>
rect 374 125 375 126 
<< pdiffusion >>
rect 375 125 376 126 
<< pdiffusion >>
rect 376 125 377 126 
<< pdiffusion >>
rect 377 125 378 126 
<< m1 >>
rect 388 125 389 126 
<< pdiffusion >>
rect 390 125 391 126 
<< pdiffusion >>
rect 391 125 392 126 
<< pdiffusion >>
rect 392 125 393 126 
<< pdiffusion >>
rect 393 125 394 126 
<< m1 >>
rect 394 125 395 126 
<< pdiffusion >>
rect 394 125 395 126 
<< pdiffusion >>
rect 395 125 396 126 
<< pdiffusion >>
rect 408 125 409 126 
<< pdiffusion >>
rect 409 125 410 126 
<< pdiffusion >>
rect 410 125 411 126 
<< pdiffusion >>
rect 411 125 412 126 
<< pdiffusion >>
rect 412 125 413 126 
<< pdiffusion >>
rect 413 125 414 126 
<< pdiffusion >>
rect 426 125 427 126 
<< pdiffusion >>
rect 427 125 428 126 
<< pdiffusion >>
rect 428 125 429 126 
<< pdiffusion >>
rect 429 125 430 126 
<< m1 >>
rect 430 125 431 126 
<< pdiffusion >>
rect 430 125 431 126 
<< pdiffusion >>
rect 431 125 432 126 
<< pdiffusion >>
rect 444 125 445 126 
<< m1 >>
rect 445 125 446 126 
<< pdiffusion >>
rect 445 125 446 126 
<< pdiffusion >>
rect 446 125 447 126 
<< pdiffusion >>
rect 447 125 448 126 
<< pdiffusion >>
rect 448 125 449 126 
<< pdiffusion >>
rect 449 125 450 126 
<< m1 >>
rect 451 125 452 126 
<< m1 >>
rect 62 126 63 127 
<< m1 >>
rect 64 126 65 127 
<< m1 >>
rect 67 126 68 127 
<< m1 >>
rect 73 126 74 127 
<< m1 >>
rect 93 126 94 127 
<< m2 >>
rect 115 126 116 127 
<< m1 >>
rect 116 126 117 127 
<< m1 >>
rect 118 126 119 127 
<< m1 >>
rect 124 126 125 127 
<< m1 >>
rect 142 126 143 127 
<< m1 >>
rect 145 126 146 127 
<< m2 >>
rect 145 126 146 127 
<< m1 >>
rect 178 126 179 127 
<< m1 >>
rect 193 126 194 127 
<< m1 >>
rect 199 126 200 127 
<< m1 >>
rect 214 126 215 127 
<< m1 >>
rect 222 126 223 127 
<< m1 >>
rect 226 126 227 127 
<< m1 >>
rect 262 126 263 127 
<< m1 >>
rect 271 126 272 127 
<< m2 >>
rect 280 126 281 127 
<< m1 >>
rect 283 126 284 127 
<< m1 >>
rect 286 126 287 127 
<< m1 >>
rect 298 126 299 127 
<< m1 >>
rect 307 126 308 127 
<< m1 >>
rect 319 126 320 127 
<< m1 >>
rect 334 126 335 127 
<< m1 >>
rect 388 126 389 127 
<< m1 >>
rect 394 126 395 127 
<< m1 >>
rect 430 126 431 127 
<< m1 >>
rect 445 126 446 127 
<< m1 >>
rect 451 126 452 127 
<< m1 >>
rect 62 127 63 128 
<< m2 >>
rect 62 127 63 128 
<< m2c >>
rect 62 127 63 128 
<< m1 >>
rect 62 127 63 128 
<< m2 >>
rect 62 127 63 128 
<< m2 >>
rect 63 127 64 128 
<< m1 >>
rect 64 127 65 128 
<< m2 >>
rect 64 127 65 128 
<< m2 >>
rect 65 127 66 128 
<< m1 >>
rect 66 127 67 128 
<< m2 >>
rect 66 127 67 128 
<< m2c >>
rect 66 127 67 128 
<< m1 >>
rect 66 127 67 128 
<< m2 >>
rect 66 127 67 128 
<< m1 >>
rect 67 127 68 128 
<< m1 >>
rect 73 127 74 128 
<< m1 >>
rect 93 127 94 128 
<< m2 >>
rect 115 127 116 128 
<< m1 >>
rect 116 127 117 128 
<< m1 >>
rect 118 127 119 128 
<< m1 >>
rect 124 127 125 128 
<< m1 >>
rect 142 127 143 128 
<< m1 >>
rect 143 127 144 128 
<< m2 >>
rect 143 127 144 128 
<< m2c >>
rect 143 127 144 128 
<< m1 >>
rect 143 127 144 128 
<< m2 >>
rect 143 127 144 128 
<< m2 >>
rect 144 127 145 128 
<< m1 >>
rect 145 127 146 128 
<< m2 >>
rect 145 127 146 128 
<< m1 >>
rect 178 127 179 128 
<< m1 >>
rect 193 127 194 128 
<< m1 >>
rect 199 127 200 128 
<< m1 >>
rect 214 127 215 128 
<< m1 >>
rect 222 127 223 128 
<< m1 >>
rect 226 127 227 128 
<< m1 >>
rect 262 127 263 128 
<< m1 >>
rect 271 127 272 128 
<< m2 >>
rect 272 127 273 128 
<< m1 >>
rect 273 127 274 128 
<< m2 >>
rect 273 127 274 128 
<< m2c >>
rect 273 127 274 128 
<< m1 >>
rect 273 127 274 128 
<< m2 >>
rect 273 127 274 128 
<< m1 >>
rect 274 127 275 128 
<< m1 >>
rect 275 127 276 128 
<< m1 >>
rect 276 127 277 128 
<< m1 >>
rect 277 127 278 128 
<< m1 >>
rect 278 127 279 128 
<< m1 >>
rect 279 127 280 128 
<< m1 >>
rect 280 127 281 128 
<< m2 >>
rect 280 127 281 128 
<< m1 >>
rect 281 127 282 128 
<< m1 >>
rect 282 127 283 128 
<< m1 >>
rect 283 127 284 128 
<< m1 >>
rect 286 127 287 128 
<< m1 >>
rect 287 127 288 128 
<< m1 >>
rect 288 127 289 128 
<< m1 >>
rect 289 127 290 128 
<< m1 >>
rect 290 127 291 128 
<< m1 >>
rect 291 127 292 128 
<< m1 >>
rect 292 127 293 128 
<< m1 >>
rect 293 127 294 128 
<< m1 >>
rect 294 127 295 128 
<< m1 >>
rect 295 127 296 128 
<< m1 >>
rect 296 127 297 128 
<< m1 >>
rect 297 127 298 128 
<< m1 >>
rect 298 127 299 128 
<< m1 >>
rect 307 127 308 128 
<< m1 >>
rect 319 127 320 128 
<< m1 >>
rect 334 127 335 128 
<< m1 >>
rect 388 127 389 128 
<< m1 >>
rect 394 127 395 128 
<< m1 >>
rect 430 127 431 128 
<< m1 >>
rect 445 127 446 128 
<< m1 >>
rect 451 127 452 128 
<< m1 >>
rect 64 128 65 129 
<< m1 >>
rect 73 128 74 129 
<< m1 >>
rect 93 128 94 129 
<< m1 >>
rect 95 128 96 129 
<< m1 >>
rect 96 128 97 129 
<< m1 >>
rect 97 128 98 129 
<< m1 >>
rect 98 128 99 129 
<< m1 >>
rect 99 128 100 129 
<< m1 >>
rect 100 128 101 129 
<< m1 >>
rect 101 128 102 129 
<< m1 >>
rect 102 128 103 129 
<< m1 >>
rect 103 128 104 129 
<< m1 >>
rect 104 128 105 129 
<< m1 >>
rect 105 128 106 129 
<< m1 >>
rect 106 128 107 129 
<< m1 >>
rect 107 128 108 129 
<< m1 >>
rect 108 128 109 129 
<< m1 >>
rect 109 128 110 129 
<< m1 >>
rect 110 128 111 129 
<< m1 >>
rect 111 128 112 129 
<< m1 >>
rect 112 128 113 129 
<< m1 >>
rect 113 128 114 129 
<< m1 >>
rect 114 128 115 129 
<< m2 >>
rect 114 128 115 129 
<< m2c >>
rect 114 128 115 129 
<< m1 >>
rect 114 128 115 129 
<< m2 >>
rect 114 128 115 129 
<< m2 >>
rect 115 128 116 129 
<< m1 >>
rect 116 128 117 129 
<< m1 >>
rect 118 128 119 129 
<< m1 >>
rect 124 128 125 129 
<< m1 >>
rect 145 128 146 129 
<< m1 >>
rect 178 128 179 129 
<< m1 >>
rect 193 128 194 129 
<< m1 >>
rect 194 128 195 129 
<< m1 >>
rect 195 128 196 129 
<< m1 >>
rect 196 128 197 129 
<< m1 >>
rect 197 128 198 129 
<< m2 >>
rect 197 128 198 129 
<< m2c >>
rect 197 128 198 129 
<< m1 >>
rect 197 128 198 129 
<< m2 >>
rect 197 128 198 129 
<< m2 >>
rect 198 128 199 129 
<< m1 >>
rect 199 128 200 129 
<< m1 >>
rect 214 128 215 129 
<< m1 >>
rect 222 128 223 129 
<< m2 >>
rect 222 128 223 129 
<< m2c >>
rect 222 128 223 129 
<< m1 >>
rect 222 128 223 129 
<< m2 >>
rect 222 128 223 129 
<< m1 >>
rect 226 128 227 129 
<< m1 >>
rect 262 128 263 129 
<< m2 >>
rect 262 128 263 129 
<< m2c >>
rect 262 128 263 129 
<< m1 >>
rect 262 128 263 129 
<< m2 >>
rect 262 128 263 129 
<< m1 >>
rect 266 128 267 129 
<< m2 >>
rect 266 128 267 129 
<< m2c >>
rect 266 128 267 129 
<< m1 >>
rect 266 128 267 129 
<< m2 >>
rect 266 128 267 129 
<< m2 >>
rect 267 128 268 129 
<< m1 >>
rect 268 128 269 129 
<< m2 >>
rect 268 128 269 129 
<< m1 >>
rect 269 128 270 129 
<< m2 >>
rect 269 128 270 129 
<< m1 >>
rect 270 128 271 129 
<< m2 >>
rect 270 128 271 129 
<< m1 >>
rect 271 128 272 129 
<< m2 >>
rect 271 128 272 129 
<< m2 >>
rect 272 128 273 129 
<< m2 >>
rect 280 128 281 129 
<< m1 >>
rect 307 128 308 129 
<< m1 >>
rect 319 128 320 129 
<< m1 >>
rect 334 128 335 129 
<< m1 >>
rect 376 128 377 129 
<< m1 >>
rect 377 128 378 129 
<< m1 >>
rect 378 128 379 129 
<< m1 >>
rect 379 128 380 129 
<< m1 >>
rect 380 128 381 129 
<< m1 >>
rect 381 128 382 129 
<< m1 >>
rect 382 128 383 129 
<< m1 >>
rect 383 128 384 129 
<< m1 >>
rect 384 128 385 129 
<< m1 >>
rect 385 128 386 129 
<< m1 >>
rect 386 128 387 129 
<< m1 >>
rect 387 128 388 129 
<< m1 >>
rect 388 128 389 129 
<< m1 >>
rect 394 128 395 129 
<< m1 >>
rect 430 128 431 129 
<< m1 >>
rect 445 128 446 129 
<< m1 >>
rect 446 128 447 129 
<< m1 >>
rect 447 128 448 129 
<< m1 >>
rect 448 128 449 129 
<< m1 >>
rect 449 128 450 129 
<< m1 >>
rect 450 128 451 129 
<< m1 >>
rect 451 128 452 129 
<< m1 >>
rect 64 129 65 130 
<< m1 >>
rect 73 129 74 130 
<< m1 >>
rect 93 129 94 130 
<< m1 >>
rect 95 129 96 130 
<< m1 >>
rect 116 129 117 130 
<< m1 >>
rect 118 129 119 130 
<< m1 >>
rect 124 129 125 130 
<< m1 >>
rect 145 129 146 130 
<< m1 >>
rect 178 129 179 130 
<< m2 >>
rect 198 129 199 130 
<< m1 >>
rect 199 129 200 130 
<< m1 >>
rect 214 129 215 130 
<< m2 >>
rect 222 129 223 130 
<< m1 >>
rect 226 129 227 130 
<< m2 >>
rect 254 129 255 130 
<< m2 >>
rect 255 129 256 130 
<< m2 >>
rect 256 129 257 130 
<< m2 >>
rect 257 129 258 130 
<< m2 >>
rect 258 129 259 130 
<< m2 >>
rect 259 129 260 130 
<< m2 >>
rect 260 129 261 130 
<< m2 >>
rect 261 129 262 130 
<< m2 >>
rect 262 129 263 130 
<< m1 >>
rect 266 129 267 130 
<< m1 >>
rect 268 129 269 130 
<< m1 >>
rect 280 129 281 130 
<< m2 >>
rect 280 129 281 130 
<< m2c >>
rect 280 129 281 130 
<< m1 >>
rect 280 129 281 130 
<< m2 >>
rect 280 129 281 130 
<< m1 >>
rect 307 129 308 130 
<< m1 >>
rect 319 129 320 130 
<< m1 >>
rect 334 129 335 130 
<< m1 >>
rect 376 129 377 130 
<< m1 >>
rect 394 129 395 130 
<< m1 >>
rect 430 129 431 130 
<< m1 >>
rect 64 130 65 131 
<< m1 >>
rect 73 130 74 131 
<< m1 >>
rect 93 130 94 131 
<< m1 >>
rect 95 130 96 131 
<< m1 >>
rect 116 130 117 131 
<< m2 >>
rect 116 130 117 131 
<< m2c >>
rect 116 130 117 131 
<< m1 >>
rect 116 130 117 131 
<< m2 >>
rect 116 130 117 131 
<< m2 >>
rect 117 130 118 131 
<< m1 >>
rect 118 130 119 131 
<< m2 >>
rect 118 130 119 131 
<< m2 >>
rect 119 130 120 131 
<< m1 >>
rect 120 130 121 131 
<< m2 >>
rect 120 130 121 131 
<< m2c >>
rect 120 130 121 131 
<< m1 >>
rect 120 130 121 131 
<< m2 >>
rect 120 130 121 131 
<< m1 >>
rect 121 130 122 131 
<< m1 >>
rect 122 130 123 131 
<< m1 >>
rect 123 130 124 131 
<< m1 >>
rect 124 130 125 131 
<< m1 >>
rect 145 130 146 131 
<< m1 >>
rect 170 130 171 131 
<< m1 >>
rect 171 130 172 131 
<< m1 >>
rect 172 130 173 131 
<< m1 >>
rect 173 130 174 131 
<< m1 >>
rect 174 130 175 131 
<< m1 >>
rect 175 130 176 131 
<< m1 >>
rect 176 130 177 131 
<< m1 >>
rect 177 130 178 131 
<< m1 >>
rect 178 130 179 131 
<< m2 >>
rect 198 130 199 131 
<< m1 >>
rect 199 130 200 131 
<< m2 >>
rect 199 130 200 131 
<< m1 >>
rect 200 130 201 131 
<< m2 >>
rect 200 130 201 131 
<< m1 >>
rect 201 130 202 131 
<< m2 >>
rect 201 130 202 131 
<< m1 >>
rect 202 130 203 131 
<< m2 >>
rect 202 130 203 131 
<< m1 >>
rect 203 130 204 131 
<< m2 >>
rect 203 130 204 131 
<< m1 >>
rect 204 130 205 131 
<< m2 >>
rect 204 130 205 131 
<< m1 >>
rect 205 130 206 131 
<< m2 >>
rect 205 130 206 131 
<< m1 >>
rect 206 130 207 131 
<< m2 >>
rect 206 130 207 131 
<< m1 >>
rect 207 130 208 131 
<< m2 >>
rect 207 130 208 131 
<< m1 >>
rect 208 130 209 131 
<< m2 >>
rect 208 130 209 131 
<< m1 >>
rect 209 130 210 131 
<< m2 >>
rect 209 130 210 131 
<< m1 >>
rect 210 130 211 131 
<< m2 >>
rect 210 130 211 131 
<< m1 >>
rect 211 130 212 131 
<< m2 >>
rect 211 130 212 131 
<< m1 >>
rect 212 130 213 131 
<< m2 >>
rect 212 130 213 131 
<< m1 >>
rect 213 130 214 131 
<< m2 >>
rect 213 130 214 131 
<< m1 >>
rect 214 130 215 131 
<< m2 >>
rect 214 130 215 131 
<< m2 >>
rect 215 130 216 131 
<< m1 >>
rect 216 130 217 131 
<< m2 >>
rect 216 130 217 131 
<< m2c >>
rect 216 130 217 131 
<< m1 >>
rect 216 130 217 131 
<< m2 >>
rect 216 130 217 131 
<< m1 >>
rect 217 130 218 131 
<< m1 >>
rect 218 130 219 131 
<< m1 >>
rect 219 130 220 131 
<< m1 >>
rect 220 130 221 131 
<< m1 >>
rect 221 130 222 131 
<< m1 >>
rect 222 130 223 131 
<< m2 >>
rect 222 130 223 131 
<< m1 >>
rect 223 130 224 131 
<< m1 >>
rect 224 130 225 131 
<< m2 >>
rect 224 130 225 131 
<< m2c >>
rect 224 130 225 131 
<< m1 >>
rect 224 130 225 131 
<< m2 >>
rect 224 130 225 131 
<< m2 >>
rect 225 130 226 131 
<< m1 >>
rect 226 130 227 131 
<< m1 >>
rect 229 130 230 131 
<< m1 >>
rect 230 130 231 131 
<< m1 >>
rect 231 130 232 131 
<< m1 >>
rect 232 130 233 131 
<< m1 >>
rect 233 130 234 131 
<< m1 >>
rect 234 130 235 131 
<< m1 >>
rect 235 130 236 131 
<< m1 >>
rect 236 130 237 131 
<< m1 >>
rect 237 130 238 131 
<< m1 >>
rect 238 130 239 131 
<< m1 >>
rect 239 130 240 131 
<< m1 >>
rect 240 130 241 131 
<< m1 >>
rect 241 130 242 131 
<< m1 >>
rect 242 130 243 131 
<< m1 >>
rect 243 130 244 131 
<< m1 >>
rect 244 130 245 131 
<< m1 >>
rect 245 130 246 131 
<< m1 >>
rect 246 130 247 131 
<< m1 >>
rect 247 130 248 131 
<< m1 >>
rect 248 130 249 131 
<< m1 >>
rect 249 130 250 131 
<< m1 >>
rect 250 130 251 131 
<< m1 >>
rect 251 130 252 131 
<< m1 >>
rect 252 130 253 131 
<< m1 >>
rect 253 130 254 131 
<< m1 >>
rect 254 130 255 131 
<< m2 >>
rect 254 130 255 131 
<< m1 >>
rect 255 130 256 131 
<< m1 >>
rect 256 130 257 131 
<< m1 >>
rect 257 130 258 131 
<< m1 >>
rect 258 130 259 131 
<< m1 >>
rect 259 130 260 131 
<< m1 >>
rect 260 130 261 131 
<< m1 >>
rect 261 130 262 131 
<< m1 >>
rect 262 130 263 131 
<< m1 >>
rect 263 130 264 131 
<< m1 >>
rect 264 130 265 131 
<< m1 >>
rect 265 130 266 131 
<< m1 >>
rect 266 130 267 131 
<< m1 >>
rect 268 130 269 131 
<< m1 >>
rect 280 130 281 131 
<< m1 >>
rect 307 130 308 131 
<< m1 >>
rect 319 130 320 131 
<< m1 >>
rect 334 130 335 131 
<< m1 >>
rect 376 130 377 131 
<< m1 >>
rect 394 130 395 131 
<< m1 >>
rect 395 130 396 131 
<< m1 >>
rect 396 130 397 131 
<< m1 >>
rect 397 130 398 131 
<< m1 >>
rect 398 130 399 131 
<< m1 >>
rect 399 130 400 131 
<< m1 >>
rect 400 130 401 131 
<< m1 >>
rect 401 130 402 131 
<< m1 >>
rect 402 130 403 131 
<< m1 >>
rect 403 130 404 131 
<< m1 >>
rect 404 130 405 131 
<< m1 >>
rect 405 130 406 131 
<< m1 >>
rect 406 130 407 131 
<< m1 >>
rect 407 130 408 131 
<< m1 >>
rect 408 130 409 131 
<< m1 >>
rect 409 130 410 131 
<< m1 >>
rect 410 130 411 131 
<< m1 >>
rect 411 130 412 131 
<< m1 >>
rect 412 130 413 131 
<< m1 >>
rect 413 130 414 131 
<< m1 >>
rect 414 130 415 131 
<< m1 >>
rect 415 130 416 131 
<< m1 >>
rect 416 130 417 131 
<< m1 >>
rect 417 130 418 131 
<< m1 >>
rect 418 130 419 131 
<< m1 >>
rect 419 130 420 131 
<< m1 >>
rect 420 130 421 131 
<< m1 >>
rect 421 130 422 131 
<< m1 >>
rect 422 130 423 131 
<< m1 >>
rect 423 130 424 131 
<< m1 >>
rect 424 130 425 131 
<< m1 >>
rect 425 130 426 131 
<< m1 >>
rect 426 130 427 131 
<< m1 >>
rect 427 130 428 131 
<< m1 >>
rect 428 130 429 131 
<< m1 >>
rect 429 130 430 131 
<< m1 >>
rect 430 130 431 131 
<< m1 >>
rect 64 131 65 132 
<< m1 >>
rect 73 131 74 132 
<< m1 >>
rect 93 131 94 132 
<< m1 >>
rect 95 131 96 132 
<< m1 >>
rect 118 131 119 132 
<< m1 >>
rect 145 131 146 132 
<< m1 >>
rect 170 131 171 132 
<< m2 >>
rect 222 131 223 132 
<< m2 >>
rect 225 131 226 132 
<< m1 >>
rect 226 131 227 132 
<< m1 >>
rect 229 131 230 132 
<< m2 >>
rect 254 131 255 132 
<< m1 >>
rect 268 131 269 132 
<< m1 >>
rect 280 131 281 132 
<< m2 >>
rect 280 131 281 132 
<< m2c >>
rect 280 131 281 132 
<< m1 >>
rect 280 131 281 132 
<< m2 >>
rect 280 131 281 132 
<< m1 >>
rect 307 131 308 132 
<< m1 >>
rect 319 131 320 132 
<< m1 >>
rect 334 131 335 132 
<< m1 >>
rect 376 131 377 132 
<< m1 >>
rect 64 132 65 133 
<< m1 >>
rect 73 132 74 133 
<< m1 >>
rect 93 132 94 133 
<< m1 >>
rect 95 132 96 133 
<< m1 >>
rect 118 132 119 133 
<< m1 >>
rect 145 132 146 133 
<< m1 >>
rect 170 132 171 133 
<< m1 >>
rect 208 132 209 133 
<< m1 >>
rect 209 132 210 133 
<< m1 >>
rect 210 132 211 133 
<< m1 >>
rect 211 132 212 133 
<< m1 >>
rect 212 132 213 133 
<< m1 >>
rect 213 132 214 133 
<< m1 >>
rect 214 132 215 133 
<< m1 >>
rect 215 132 216 133 
<< m1 >>
rect 216 132 217 133 
<< m1 >>
rect 217 132 218 133 
<< m1 >>
rect 218 132 219 133 
<< m1 >>
rect 219 132 220 133 
<< m1 >>
rect 220 132 221 133 
<< m1 >>
rect 221 132 222 133 
<< m1 >>
rect 222 132 223 133 
<< m2 >>
rect 222 132 223 133 
<< m2c >>
rect 222 132 223 133 
<< m1 >>
rect 222 132 223 133 
<< m2 >>
rect 222 132 223 133 
<< m2 >>
rect 225 132 226 133 
<< m1 >>
rect 226 132 227 133 
<< m1 >>
rect 229 132 230 133 
<< m2 >>
rect 254 132 255 133 
<< m1 >>
rect 268 132 269 133 
<< m2 >>
rect 280 132 281 133 
<< m1 >>
rect 307 132 308 133 
<< m1 >>
rect 319 132 320 133 
<< m1 >>
rect 334 132 335 133 
<< m1 >>
rect 376 132 377 133 
<< m1 >>
rect 28 133 29 134 
<< m1 >>
rect 29 133 30 134 
<< m1 >>
rect 30 133 31 134 
<< m1 >>
rect 31 133 32 134 
<< m1 >>
rect 32 133 33 134 
<< m1 >>
rect 33 133 34 134 
<< m1 >>
rect 34 133 35 134 
<< m1 >>
rect 64 133 65 134 
<< m1 >>
rect 73 133 74 134 
<< m1 >>
rect 93 133 94 134 
<< m1 >>
rect 95 133 96 134 
<< m1 >>
rect 118 133 119 134 
<< m1 >>
rect 145 133 146 134 
<< m1 >>
rect 170 133 171 134 
<< m1 >>
rect 208 133 209 134 
<< m2 >>
rect 225 133 226 134 
<< m1 >>
rect 226 133 227 134 
<< m1 >>
rect 229 133 230 134 
<< m1 >>
rect 244 133 245 134 
<< m1 >>
rect 245 133 246 134 
<< m1 >>
rect 246 133 247 134 
<< m1 >>
rect 247 133 248 134 
<< m1 >>
rect 248 133 249 134 
<< m1 >>
rect 249 133 250 134 
<< m1 >>
rect 250 133 251 134 
<< m1 >>
rect 251 133 252 134 
<< m1 >>
rect 252 133 253 134 
<< m1 >>
rect 253 133 254 134 
<< m1 >>
rect 254 133 255 134 
<< m2 >>
rect 254 133 255 134 
<< m1 >>
rect 255 133 256 134 
<< m1 >>
rect 256 133 257 134 
<< m1 >>
rect 257 133 258 134 
<< m1 >>
rect 258 133 259 134 
<< m1 >>
rect 259 133 260 134 
<< m1 >>
rect 260 133 261 134 
<< m1 >>
rect 261 133 262 134 
<< m1 >>
rect 262 133 263 134 
<< m1 >>
rect 263 133 264 134 
<< m1 >>
rect 264 133 265 134 
<< m1 >>
rect 265 133 266 134 
<< m1 >>
rect 266 133 267 134 
<< m2 >>
rect 266 133 267 134 
<< m2c >>
rect 266 133 267 134 
<< m1 >>
rect 266 133 267 134 
<< m2 >>
rect 266 133 267 134 
<< m2 >>
rect 267 133 268 134 
<< m1 >>
rect 268 133 269 134 
<< m2 >>
rect 268 133 269 134 
<< m2 >>
rect 269 133 270 134 
<< m1 >>
rect 270 133 271 134 
<< m2 >>
rect 270 133 271 134 
<< m2c >>
rect 270 133 271 134 
<< m1 >>
rect 270 133 271 134 
<< m2 >>
rect 270 133 271 134 
<< m1 >>
rect 271 133 272 134 
<< m1 >>
rect 272 133 273 134 
<< m1 >>
rect 273 133 274 134 
<< m1 >>
rect 274 133 275 134 
<< m1 >>
rect 275 133 276 134 
<< m1 >>
rect 276 133 277 134 
<< m1 >>
rect 277 133 278 134 
<< m1 >>
rect 278 133 279 134 
<< m1 >>
rect 279 133 280 134 
<< m1 >>
rect 280 133 281 134 
<< m2 >>
rect 280 133 281 134 
<< m1 >>
rect 281 133 282 134 
<< m1 >>
rect 282 133 283 134 
<< m1 >>
rect 283 133 284 134 
<< m1 >>
rect 284 133 285 134 
<< m1 >>
rect 285 133 286 134 
<< m1 >>
rect 286 133 287 134 
<< m1 >>
rect 287 133 288 134 
<< m1 >>
rect 288 133 289 134 
<< m1 >>
rect 289 133 290 134 
<< m1 >>
rect 290 133 291 134 
<< m1 >>
rect 291 133 292 134 
<< m1 >>
rect 292 133 293 134 
<< m1 >>
rect 293 133 294 134 
<< m1 >>
rect 294 133 295 134 
<< m1 >>
rect 295 133 296 134 
<< m1 >>
rect 296 133 297 134 
<< m1 >>
rect 297 133 298 134 
<< m1 >>
rect 298 133 299 134 
<< m1 >>
rect 299 133 300 134 
<< m1 >>
rect 300 133 301 134 
<< m1 >>
rect 301 133 302 134 
<< m1 >>
rect 302 133 303 134 
<< m1 >>
rect 303 133 304 134 
<< m1 >>
rect 304 133 305 134 
<< m1 >>
rect 307 133 308 134 
<< m1 >>
rect 311 133 312 134 
<< m1 >>
rect 312 133 313 134 
<< m1 >>
rect 313 133 314 134 
<< m1 >>
rect 314 133 315 134 
<< m1 >>
rect 315 133 316 134 
<< m1 >>
rect 316 133 317 134 
<< m1 >>
rect 317 133 318 134 
<< m1 >>
rect 318 133 319 134 
<< m1 >>
rect 319 133 320 134 
<< m1 >>
rect 334 133 335 134 
<< m1 >>
rect 335 133 336 134 
<< m1 >>
rect 336 133 337 134 
<< m1 >>
rect 337 133 338 134 
<< m1 >>
rect 338 133 339 134 
<< m1 >>
rect 339 133 340 134 
<< m1 >>
rect 340 133 341 134 
<< m1 >>
rect 343 133 344 134 
<< m1 >>
rect 344 133 345 134 
<< m1 >>
rect 345 133 346 134 
<< m1 >>
rect 346 133 347 134 
<< m1 >>
rect 347 133 348 134 
<< m1 >>
rect 348 133 349 134 
<< m1 >>
rect 349 133 350 134 
<< m1 >>
rect 350 133 351 134 
<< m1 >>
rect 351 133 352 134 
<< m1 >>
rect 352 133 353 134 
<< m1 >>
rect 353 133 354 134 
<< m1 >>
rect 354 133 355 134 
<< m1 >>
rect 355 133 356 134 
<< m1 >>
rect 356 133 357 134 
<< m1 >>
rect 357 133 358 134 
<< m1 >>
rect 358 133 359 134 
<< m1 >>
rect 376 133 377 134 
<< m1 >>
rect 28 134 29 135 
<< m1 >>
rect 34 134 35 135 
<< m1 >>
rect 64 134 65 135 
<< m1 >>
rect 73 134 74 135 
<< m1 >>
rect 93 134 94 135 
<< m1 >>
rect 95 134 96 135 
<< m1 >>
rect 118 134 119 135 
<< m1 >>
rect 145 134 146 135 
<< m1 >>
rect 170 134 171 135 
<< m1 >>
rect 208 134 209 135 
<< m2 >>
rect 225 134 226 135 
<< m1 >>
rect 226 134 227 135 
<< m1 >>
rect 229 134 230 135 
<< m1 >>
rect 244 134 245 135 
<< m2 >>
rect 254 134 255 135 
<< m1 >>
rect 268 134 269 135 
<< m2 >>
rect 280 134 281 135 
<< m1 >>
rect 304 134 305 135 
<< m1 >>
rect 307 134 308 135 
<< m1 >>
rect 311 134 312 135 
<< m1 >>
rect 340 134 341 135 
<< m1 >>
rect 343 134 344 135 
<< m1 >>
rect 358 134 359 135 
<< m1 >>
rect 376 134 377 135 
<< m1 >>
rect 28 135 29 136 
<< m1 >>
rect 34 135 35 136 
<< m1 >>
rect 64 135 65 136 
<< m1 >>
rect 67 135 68 136 
<< m1 >>
rect 68 135 69 136 
<< m1 >>
rect 69 135 70 136 
<< m1 >>
rect 70 135 71 136 
<< m1 >>
rect 71 135 72 136 
<< m1 >>
rect 72 135 73 136 
<< m1 >>
rect 73 135 74 136 
<< m1 >>
rect 93 135 94 136 
<< m1 >>
rect 95 135 96 136 
<< m1 >>
rect 118 135 119 136 
<< m1 >>
rect 145 135 146 136 
<< m1 >>
rect 170 135 171 136 
<< m1 >>
rect 208 135 209 136 
<< m2 >>
rect 225 135 226 136 
<< m1 >>
rect 226 135 227 136 
<< m1 >>
rect 229 135 230 136 
<< m1 >>
rect 244 135 245 136 
<< m2 >>
rect 254 135 255 136 
<< m1 >>
rect 268 135 269 136 
<< m1 >>
rect 280 135 281 136 
<< m2 >>
rect 280 135 281 136 
<< m2c >>
rect 280 135 281 136 
<< m1 >>
rect 280 135 281 136 
<< m2 >>
rect 280 135 281 136 
<< m1 >>
rect 281 135 282 136 
<< m1 >>
rect 282 135 283 136 
<< m1 >>
rect 283 135 284 136 
<< m1 >>
rect 304 135 305 136 
<< m1 >>
rect 307 135 308 136 
<< m1 >>
rect 311 135 312 136 
<< m1 >>
rect 340 135 341 136 
<< m1 >>
rect 343 135 344 136 
<< m1 >>
rect 358 135 359 136 
<< m1 >>
rect 376 135 377 136 
<< m1 >>
rect 28 136 29 137 
<< m1 >>
rect 34 136 35 137 
<< m1 >>
rect 64 136 65 137 
<< m1 >>
rect 67 136 68 137 
<< m1 >>
rect 93 136 94 137 
<< m1 >>
rect 95 136 96 137 
<< m1 >>
rect 106 136 107 137 
<< m1 >>
rect 107 136 108 137 
<< m1 >>
rect 108 136 109 137 
<< m1 >>
rect 109 136 110 137 
<< m1 >>
rect 110 136 111 137 
<< m1 >>
rect 111 136 112 137 
<< m1 >>
rect 112 136 113 137 
<< m1 >>
rect 113 136 114 137 
<< m1 >>
rect 114 136 115 137 
<< m1 >>
rect 115 136 116 137 
<< m1 >>
rect 116 136 117 137 
<< m1 >>
rect 118 136 119 137 
<< m1 >>
rect 145 136 146 137 
<< m1 >>
rect 170 136 171 137 
<< m1 >>
rect 172 136 173 137 
<< m1 >>
rect 173 136 174 137 
<< m1 >>
rect 174 136 175 137 
<< m1 >>
rect 175 136 176 137 
<< m1 >>
rect 208 136 209 137 
<< m2 >>
rect 225 136 226 137 
<< m1 >>
rect 226 136 227 137 
<< m1 >>
rect 229 136 230 137 
<< m1 >>
rect 244 136 245 137 
<< m1 >>
rect 253 136 254 137 
<< m1 >>
rect 254 136 255 137 
<< m2 >>
rect 254 136 255 137 
<< m1 >>
rect 255 136 256 137 
<< m1 >>
rect 256 136 257 137 
<< m1 >>
rect 257 136 258 137 
<< m1 >>
rect 258 136 259 137 
<< m1 >>
rect 259 136 260 137 
<< m1 >>
rect 260 136 261 137 
<< m1 >>
rect 261 136 262 137 
<< m1 >>
rect 262 136 263 137 
<< m1 >>
rect 263 136 264 137 
<< m1 >>
rect 264 136 265 137 
<< m1 >>
rect 265 136 266 137 
<< m1 >>
rect 268 136 269 137 
<< m1 >>
rect 283 136 284 137 
<< m1 >>
rect 304 136 305 137 
<< m1 >>
rect 307 136 308 137 
<< m1 >>
rect 311 136 312 137 
<< m1 >>
rect 340 136 341 137 
<< m1 >>
rect 343 136 344 137 
<< m1 >>
rect 358 136 359 137 
<< m1 >>
rect 376 136 377 137 
<< m1 >>
rect 406 136 407 137 
<< m1 >>
rect 407 136 408 137 
<< m1 >>
rect 408 136 409 137 
<< m1 >>
rect 409 136 410 137 
<< m1 >>
rect 28 137 29 138 
<< m1 >>
rect 34 137 35 138 
<< m1 >>
rect 64 137 65 138 
<< m1 >>
rect 67 137 68 138 
<< m1 >>
rect 93 137 94 138 
<< m1 >>
rect 95 137 96 138 
<< m1 >>
rect 106 137 107 138 
<< m1 >>
rect 116 137 117 138 
<< m1 >>
rect 118 137 119 138 
<< m1 >>
rect 145 137 146 138 
<< m1 >>
rect 170 137 171 138 
<< m1 >>
rect 172 137 173 138 
<< m1 >>
rect 175 137 176 138 
<< m1 >>
rect 208 137 209 138 
<< m2 >>
rect 225 137 226 138 
<< m1 >>
rect 226 137 227 138 
<< m1 >>
rect 229 137 230 138 
<< m1 >>
rect 244 137 245 138 
<< m1 >>
rect 253 137 254 138 
<< m2 >>
rect 254 137 255 138 
<< m1 >>
rect 265 137 266 138 
<< m1 >>
rect 268 137 269 138 
<< m1 >>
rect 283 137 284 138 
<< m1 >>
rect 304 137 305 138 
<< m1 >>
rect 307 137 308 138 
<< m1 >>
rect 311 137 312 138 
<< m1 >>
rect 340 137 341 138 
<< m1 >>
rect 343 137 344 138 
<< m1 >>
rect 358 137 359 138 
<< m1 >>
rect 376 137 377 138 
<< m1 >>
rect 406 137 407 138 
<< m1 >>
rect 409 137 410 138 
<< pdiffusion >>
rect 12 138 13 139 
<< pdiffusion >>
rect 13 138 14 139 
<< pdiffusion >>
rect 14 138 15 139 
<< pdiffusion >>
rect 15 138 16 139 
<< pdiffusion >>
rect 16 138 17 139 
<< pdiffusion >>
rect 17 138 18 139 
<< m1 >>
rect 28 138 29 139 
<< pdiffusion >>
rect 30 138 31 139 
<< pdiffusion >>
rect 31 138 32 139 
<< pdiffusion >>
rect 32 138 33 139 
<< pdiffusion >>
rect 33 138 34 139 
<< m1 >>
rect 34 138 35 139 
<< pdiffusion >>
rect 34 138 35 139 
<< pdiffusion >>
rect 35 138 36 139 
<< pdiffusion >>
rect 48 138 49 139 
<< pdiffusion >>
rect 49 138 50 139 
<< pdiffusion >>
rect 50 138 51 139 
<< pdiffusion >>
rect 51 138 52 139 
<< pdiffusion >>
rect 52 138 53 139 
<< pdiffusion >>
rect 53 138 54 139 
<< m1 >>
rect 64 138 65 139 
<< pdiffusion >>
rect 66 138 67 139 
<< m1 >>
rect 67 138 68 139 
<< pdiffusion >>
rect 67 138 68 139 
<< pdiffusion >>
rect 68 138 69 139 
<< pdiffusion >>
rect 69 138 70 139 
<< pdiffusion >>
rect 70 138 71 139 
<< pdiffusion >>
rect 71 138 72 139 
<< pdiffusion >>
rect 84 138 85 139 
<< pdiffusion >>
rect 85 138 86 139 
<< pdiffusion >>
rect 86 138 87 139 
<< pdiffusion >>
rect 87 138 88 139 
<< pdiffusion >>
rect 88 138 89 139 
<< pdiffusion >>
rect 89 138 90 139 
<< m1 >>
rect 93 138 94 139 
<< m1 >>
rect 95 138 96 139 
<< pdiffusion >>
rect 102 138 103 139 
<< pdiffusion >>
rect 103 138 104 139 
<< pdiffusion >>
rect 104 138 105 139 
<< pdiffusion >>
rect 105 138 106 139 
<< m1 >>
rect 106 138 107 139 
<< pdiffusion >>
rect 106 138 107 139 
<< pdiffusion >>
rect 107 138 108 139 
<< m1 >>
rect 116 138 117 139 
<< m1 >>
rect 118 138 119 139 
<< pdiffusion >>
rect 120 138 121 139 
<< pdiffusion >>
rect 121 138 122 139 
<< pdiffusion >>
rect 122 138 123 139 
<< pdiffusion >>
rect 123 138 124 139 
<< pdiffusion >>
rect 124 138 125 139 
<< pdiffusion >>
rect 125 138 126 139 
<< m1 >>
rect 145 138 146 139 
<< pdiffusion >>
rect 156 138 157 139 
<< pdiffusion >>
rect 157 138 158 139 
<< pdiffusion >>
rect 158 138 159 139 
<< pdiffusion >>
rect 159 138 160 139 
<< pdiffusion >>
rect 160 138 161 139 
<< pdiffusion >>
rect 161 138 162 139 
<< m1 >>
rect 170 138 171 139 
<< m1 >>
rect 172 138 173 139 
<< pdiffusion >>
rect 174 138 175 139 
<< m1 >>
rect 175 138 176 139 
<< pdiffusion >>
rect 175 138 176 139 
<< pdiffusion >>
rect 176 138 177 139 
<< pdiffusion >>
rect 177 138 178 139 
<< pdiffusion >>
rect 178 138 179 139 
<< pdiffusion >>
rect 179 138 180 139 
<< pdiffusion >>
rect 192 138 193 139 
<< pdiffusion >>
rect 193 138 194 139 
<< pdiffusion >>
rect 194 138 195 139 
<< pdiffusion >>
rect 195 138 196 139 
<< pdiffusion >>
rect 196 138 197 139 
<< pdiffusion >>
rect 197 138 198 139 
<< m1 >>
rect 208 138 209 139 
<< pdiffusion >>
rect 210 138 211 139 
<< pdiffusion >>
rect 211 138 212 139 
<< pdiffusion >>
rect 212 138 213 139 
<< pdiffusion >>
rect 213 138 214 139 
<< pdiffusion >>
rect 214 138 215 139 
<< pdiffusion >>
rect 215 138 216 139 
<< m2 >>
rect 225 138 226 139 
<< m1 >>
rect 226 138 227 139 
<< pdiffusion >>
rect 228 138 229 139 
<< m1 >>
rect 229 138 230 139 
<< pdiffusion >>
rect 229 138 230 139 
<< pdiffusion >>
rect 230 138 231 139 
<< pdiffusion >>
rect 231 138 232 139 
<< pdiffusion >>
rect 232 138 233 139 
<< pdiffusion >>
rect 233 138 234 139 
<< m1 >>
rect 244 138 245 139 
<< pdiffusion >>
rect 246 138 247 139 
<< pdiffusion >>
rect 247 138 248 139 
<< pdiffusion >>
rect 248 138 249 139 
<< pdiffusion >>
rect 249 138 250 139 
<< pdiffusion >>
rect 250 138 251 139 
<< pdiffusion >>
rect 251 138 252 139 
<< m1 >>
rect 253 138 254 139 
<< m2 >>
rect 254 138 255 139 
<< pdiffusion >>
rect 264 138 265 139 
<< m1 >>
rect 265 138 266 139 
<< pdiffusion >>
rect 265 138 266 139 
<< pdiffusion >>
rect 266 138 267 139 
<< pdiffusion >>
rect 267 138 268 139 
<< m1 >>
rect 268 138 269 139 
<< pdiffusion >>
rect 268 138 269 139 
<< pdiffusion >>
rect 269 138 270 139 
<< pdiffusion >>
rect 282 138 283 139 
<< m1 >>
rect 283 138 284 139 
<< pdiffusion >>
rect 283 138 284 139 
<< pdiffusion >>
rect 284 138 285 139 
<< pdiffusion >>
rect 285 138 286 139 
<< pdiffusion >>
rect 286 138 287 139 
<< pdiffusion >>
rect 287 138 288 139 
<< pdiffusion >>
rect 300 138 301 139 
<< pdiffusion >>
rect 301 138 302 139 
<< pdiffusion >>
rect 302 138 303 139 
<< pdiffusion >>
rect 303 138 304 139 
<< m1 >>
rect 304 138 305 139 
<< pdiffusion >>
rect 304 138 305 139 
<< pdiffusion >>
rect 305 138 306 139 
<< m1 >>
rect 307 138 308 139 
<< m1 >>
rect 311 138 312 139 
<< pdiffusion >>
rect 318 138 319 139 
<< pdiffusion >>
rect 319 138 320 139 
<< pdiffusion >>
rect 320 138 321 139 
<< pdiffusion >>
rect 321 138 322 139 
<< pdiffusion >>
rect 322 138 323 139 
<< pdiffusion >>
rect 323 138 324 139 
<< pdiffusion >>
rect 336 138 337 139 
<< pdiffusion >>
rect 337 138 338 139 
<< pdiffusion >>
rect 338 138 339 139 
<< pdiffusion >>
rect 339 138 340 139 
<< m1 >>
rect 340 138 341 139 
<< pdiffusion >>
rect 340 138 341 139 
<< pdiffusion >>
rect 341 138 342 139 
<< m1 >>
rect 343 138 344 139 
<< pdiffusion >>
rect 354 138 355 139 
<< pdiffusion >>
rect 355 138 356 139 
<< pdiffusion >>
rect 356 138 357 139 
<< pdiffusion >>
rect 357 138 358 139 
<< m1 >>
rect 358 138 359 139 
<< pdiffusion >>
rect 358 138 359 139 
<< pdiffusion >>
rect 359 138 360 139 
<< pdiffusion >>
rect 372 138 373 139 
<< pdiffusion >>
rect 373 138 374 139 
<< pdiffusion >>
rect 374 138 375 139 
<< pdiffusion >>
rect 375 138 376 139 
<< m1 >>
rect 376 138 377 139 
<< pdiffusion >>
rect 376 138 377 139 
<< pdiffusion >>
rect 377 138 378 139 
<< m1 >>
rect 406 138 407 139 
<< pdiffusion >>
rect 408 138 409 139 
<< m1 >>
rect 409 138 410 139 
<< pdiffusion >>
rect 409 138 410 139 
<< pdiffusion >>
rect 410 138 411 139 
<< pdiffusion >>
rect 411 138 412 139 
<< pdiffusion >>
rect 412 138 413 139 
<< pdiffusion >>
rect 413 138 414 139 
<< pdiffusion >>
rect 426 138 427 139 
<< pdiffusion >>
rect 427 138 428 139 
<< pdiffusion >>
rect 428 138 429 139 
<< pdiffusion >>
rect 429 138 430 139 
<< pdiffusion >>
rect 430 138 431 139 
<< pdiffusion >>
rect 431 138 432 139 
<< pdiffusion >>
rect 444 138 445 139 
<< pdiffusion >>
rect 445 138 446 139 
<< pdiffusion >>
rect 446 138 447 139 
<< pdiffusion >>
rect 447 138 448 139 
<< pdiffusion >>
rect 448 138 449 139 
<< pdiffusion >>
rect 449 138 450 139 
<< pdiffusion >>
rect 12 139 13 140 
<< pdiffusion >>
rect 13 139 14 140 
<< pdiffusion >>
rect 14 139 15 140 
<< pdiffusion >>
rect 15 139 16 140 
<< pdiffusion >>
rect 16 139 17 140 
<< pdiffusion >>
rect 17 139 18 140 
<< m1 >>
rect 28 139 29 140 
<< pdiffusion >>
rect 30 139 31 140 
<< pdiffusion >>
rect 31 139 32 140 
<< pdiffusion >>
rect 32 139 33 140 
<< pdiffusion >>
rect 33 139 34 140 
<< pdiffusion >>
rect 34 139 35 140 
<< pdiffusion >>
rect 35 139 36 140 
<< pdiffusion >>
rect 48 139 49 140 
<< pdiffusion >>
rect 49 139 50 140 
<< pdiffusion >>
rect 50 139 51 140 
<< pdiffusion >>
rect 51 139 52 140 
<< pdiffusion >>
rect 52 139 53 140 
<< pdiffusion >>
rect 53 139 54 140 
<< m1 >>
rect 64 139 65 140 
<< pdiffusion >>
rect 66 139 67 140 
<< pdiffusion >>
rect 67 139 68 140 
<< pdiffusion >>
rect 68 139 69 140 
<< pdiffusion >>
rect 69 139 70 140 
<< pdiffusion >>
rect 70 139 71 140 
<< pdiffusion >>
rect 71 139 72 140 
<< pdiffusion >>
rect 84 139 85 140 
<< pdiffusion >>
rect 85 139 86 140 
<< pdiffusion >>
rect 86 139 87 140 
<< pdiffusion >>
rect 87 139 88 140 
<< pdiffusion >>
rect 88 139 89 140 
<< pdiffusion >>
rect 89 139 90 140 
<< m1 >>
rect 93 139 94 140 
<< m1 >>
rect 95 139 96 140 
<< pdiffusion >>
rect 102 139 103 140 
<< pdiffusion >>
rect 103 139 104 140 
<< pdiffusion >>
rect 104 139 105 140 
<< pdiffusion >>
rect 105 139 106 140 
<< pdiffusion >>
rect 106 139 107 140 
<< pdiffusion >>
rect 107 139 108 140 
<< m1 >>
rect 116 139 117 140 
<< m1 >>
rect 118 139 119 140 
<< pdiffusion >>
rect 120 139 121 140 
<< pdiffusion >>
rect 121 139 122 140 
<< pdiffusion >>
rect 122 139 123 140 
<< pdiffusion >>
rect 123 139 124 140 
<< pdiffusion >>
rect 124 139 125 140 
<< pdiffusion >>
rect 125 139 126 140 
<< m1 >>
rect 145 139 146 140 
<< pdiffusion >>
rect 156 139 157 140 
<< pdiffusion >>
rect 157 139 158 140 
<< pdiffusion >>
rect 158 139 159 140 
<< pdiffusion >>
rect 159 139 160 140 
<< pdiffusion >>
rect 160 139 161 140 
<< pdiffusion >>
rect 161 139 162 140 
<< m1 >>
rect 170 139 171 140 
<< m1 >>
rect 172 139 173 140 
<< pdiffusion >>
rect 174 139 175 140 
<< pdiffusion >>
rect 175 139 176 140 
<< pdiffusion >>
rect 176 139 177 140 
<< pdiffusion >>
rect 177 139 178 140 
<< pdiffusion >>
rect 178 139 179 140 
<< pdiffusion >>
rect 179 139 180 140 
<< pdiffusion >>
rect 192 139 193 140 
<< pdiffusion >>
rect 193 139 194 140 
<< pdiffusion >>
rect 194 139 195 140 
<< pdiffusion >>
rect 195 139 196 140 
<< pdiffusion >>
rect 196 139 197 140 
<< pdiffusion >>
rect 197 139 198 140 
<< m1 >>
rect 208 139 209 140 
<< pdiffusion >>
rect 210 139 211 140 
<< pdiffusion >>
rect 211 139 212 140 
<< pdiffusion >>
rect 212 139 213 140 
<< pdiffusion >>
rect 213 139 214 140 
<< pdiffusion >>
rect 214 139 215 140 
<< pdiffusion >>
rect 215 139 216 140 
<< m2 >>
rect 225 139 226 140 
<< m1 >>
rect 226 139 227 140 
<< pdiffusion >>
rect 228 139 229 140 
<< pdiffusion >>
rect 229 139 230 140 
<< pdiffusion >>
rect 230 139 231 140 
<< pdiffusion >>
rect 231 139 232 140 
<< pdiffusion >>
rect 232 139 233 140 
<< pdiffusion >>
rect 233 139 234 140 
<< m1 >>
rect 244 139 245 140 
<< pdiffusion >>
rect 246 139 247 140 
<< pdiffusion >>
rect 247 139 248 140 
<< pdiffusion >>
rect 248 139 249 140 
<< pdiffusion >>
rect 249 139 250 140 
<< pdiffusion >>
rect 250 139 251 140 
<< pdiffusion >>
rect 251 139 252 140 
<< m1 >>
rect 253 139 254 140 
<< m2 >>
rect 254 139 255 140 
<< pdiffusion >>
rect 264 139 265 140 
<< pdiffusion >>
rect 265 139 266 140 
<< pdiffusion >>
rect 266 139 267 140 
<< pdiffusion >>
rect 267 139 268 140 
<< pdiffusion >>
rect 268 139 269 140 
<< pdiffusion >>
rect 269 139 270 140 
<< pdiffusion >>
rect 282 139 283 140 
<< pdiffusion >>
rect 283 139 284 140 
<< pdiffusion >>
rect 284 139 285 140 
<< pdiffusion >>
rect 285 139 286 140 
<< pdiffusion >>
rect 286 139 287 140 
<< pdiffusion >>
rect 287 139 288 140 
<< pdiffusion >>
rect 300 139 301 140 
<< pdiffusion >>
rect 301 139 302 140 
<< pdiffusion >>
rect 302 139 303 140 
<< pdiffusion >>
rect 303 139 304 140 
<< pdiffusion >>
rect 304 139 305 140 
<< pdiffusion >>
rect 305 139 306 140 
<< m1 >>
rect 307 139 308 140 
<< m1 >>
rect 311 139 312 140 
<< pdiffusion >>
rect 318 139 319 140 
<< pdiffusion >>
rect 319 139 320 140 
<< pdiffusion >>
rect 320 139 321 140 
<< pdiffusion >>
rect 321 139 322 140 
<< pdiffusion >>
rect 322 139 323 140 
<< pdiffusion >>
rect 323 139 324 140 
<< pdiffusion >>
rect 336 139 337 140 
<< pdiffusion >>
rect 337 139 338 140 
<< pdiffusion >>
rect 338 139 339 140 
<< pdiffusion >>
rect 339 139 340 140 
<< pdiffusion >>
rect 340 139 341 140 
<< pdiffusion >>
rect 341 139 342 140 
<< m1 >>
rect 343 139 344 140 
<< pdiffusion >>
rect 354 139 355 140 
<< pdiffusion >>
rect 355 139 356 140 
<< pdiffusion >>
rect 356 139 357 140 
<< pdiffusion >>
rect 357 139 358 140 
<< pdiffusion >>
rect 358 139 359 140 
<< pdiffusion >>
rect 359 139 360 140 
<< pdiffusion >>
rect 372 139 373 140 
<< pdiffusion >>
rect 373 139 374 140 
<< pdiffusion >>
rect 374 139 375 140 
<< pdiffusion >>
rect 375 139 376 140 
<< pdiffusion >>
rect 376 139 377 140 
<< pdiffusion >>
rect 377 139 378 140 
<< m1 >>
rect 406 139 407 140 
<< pdiffusion >>
rect 408 139 409 140 
<< pdiffusion >>
rect 409 139 410 140 
<< pdiffusion >>
rect 410 139 411 140 
<< pdiffusion >>
rect 411 139 412 140 
<< pdiffusion >>
rect 412 139 413 140 
<< pdiffusion >>
rect 413 139 414 140 
<< pdiffusion >>
rect 426 139 427 140 
<< pdiffusion >>
rect 427 139 428 140 
<< pdiffusion >>
rect 428 139 429 140 
<< pdiffusion >>
rect 429 139 430 140 
<< pdiffusion >>
rect 430 139 431 140 
<< pdiffusion >>
rect 431 139 432 140 
<< pdiffusion >>
rect 444 139 445 140 
<< pdiffusion >>
rect 445 139 446 140 
<< pdiffusion >>
rect 446 139 447 140 
<< pdiffusion >>
rect 447 139 448 140 
<< pdiffusion >>
rect 448 139 449 140 
<< pdiffusion >>
rect 449 139 450 140 
<< pdiffusion >>
rect 12 140 13 141 
<< pdiffusion >>
rect 13 140 14 141 
<< pdiffusion >>
rect 14 140 15 141 
<< pdiffusion >>
rect 15 140 16 141 
<< pdiffusion >>
rect 16 140 17 141 
<< pdiffusion >>
rect 17 140 18 141 
<< m1 >>
rect 28 140 29 141 
<< pdiffusion >>
rect 30 140 31 141 
<< pdiffusion >>
rect 31 140 32 141 
<< pdiffusion >>
rect 32 140 33 141 
<< pdiffusion >>
rect 33 140 34 141 
<< pdiffusion >>
rect 34 140 35 141 
<< pdiffusion >>
rect 35 140 36 141 
<< pdiffusion >>
rect 48 140 49 141 
<< pdiffusion >>
rect 49 140 50 141 
<< pdiffusion >>
rect 50 140 51 141 
<< pdiffusion >>
rect 51 140 52 141 
<< pdiffusion >>
rect 52 140 53 141 
<< pdiffusion >>
rect 53 140 54 141 
<< m1 >>
rect 64 140 65 141 
<< pdiffusion >>
rect 66 140 67 141 
<< pdiffusion >>
rect 67 140 68 141 
<< pdiffusion >>
rect 68 140 69 141 
<< pdiffusion >>
rect 69 140 70 141 
<< pdiffusion >>
rect 70 140 71 141 
<< pdiffusion >>
rect 71 140 72 141 
<< pdiffusion >>
rect 84 140 85 141 
<< pdiffusion >>
rect 85 140 86 141 
<< pdiffusion >>
rect 86 140 87 141 
<< pdiffusion >>
rect 87 140 88 141 
<< pdiffusion >>
rect 88 140 89 141 
<< pdiffusion >>
rect 89 140 90 141 
<< m1 >>
rect 93 140 94 141 
<< m1 >>
rect 95 140 96 141 
<< pdiffusion >>
rect 102 140 103 141 
<< pdiffusion >>
rect 103 140 104 141 
<< pdiffusion >>
rect 104 140 105 141 
<< pdiffusion >>
rect 105 140 106 141 
<< pdiffusion >>
rect 106 140 107 141 
<< pdiffusion >>
rect 107 140 108 141 
<< m1 >>
rect 116 140 117 141 
<< m1 >>
rect 118 140 119 141 
<< pdiffusion >>
rect 120 140 121 141 
<< pdiffusion >>
rect 121 140 122 141 
<< pdiffusion >>
rect 122 140 123 141 
<< pdiffusion >>
rect 123 140 124 141 
<< pdiffusion >>
rect 124 140 125 141 
<< pdiffusion >>
rect 125 140 126 141 
<< m1 >>
rect 145 140 146 141 
<< pdiffusion >>
rect 156 140 157 141 
<< pdiffusion >>
rect 157 140 158 141 
<< pdiffusion >>
rect 158 140 159 141 
<< pdiffusion >>
rect 159 140 160 141 
<< pdiffusion >>
rect 160 140 161 141 
<< pdiffusion >>
rect 161 140 162 141 
<< m1 >>
rect 170 140 171 141 
<< m1 >>
rect 172 140 173 141 
<< pdiffusion >>
rect 174 140 175 141 
<< pdiffusion >>
rect 175 140 176 141 
<< pdiffusion >>
rect 176 140 177 141 
<< pdiffusion >>
rect 177 140 178 141 
<< pdiffusion >>
rect 178 140 179 141 
<< pdiffusion >>
rect 179 140 180 141 
<< pdiffusion >>
rect 192 140 193 141 
<< pdiffusion >>
rect 193 140 194 141 
<< pdiffusion >>
rect 194 140 195 141 
<< pdiffusion >>
rect 195 140 196 141 
<< pdiffusion >>
rect 196 140 197 141 
<< pdiffusion >>
rect 197 140 198 141 
<< m1 >>
rect 208 140 209 141 
<< pdiffusion >>
rect 210 140 211 141 
<< pdiffusion >>
rect 211 140 212 141 
<< pdiffusion >>
rect 212 140 213 141 
<< pdiffusion >>
rect 213 140 214 141 
<< pdiffusion >>
rect 214 140 215 141 
<< pdiffusion >>
rect 215 140 216 141 
<< m2 >>
rect 225 140 226 141 
<< m1 >>
rect 226 140 227 141 
<< pdiffusion >>
rect 228 140 229 141 
<< pdiffusion >>
rect 229 140 230 141 
<< pdiffusion >>
rect 230 140 231 141 
<< pdiffusion >>
rect 231 140 232 141 
<< pdiffusion >>
rect 232 140 233 141 
<< pdiffusion >>
rect 233 140 234 141 
<< m1 >>
rect 244 140 245 141 
<< pdiffusion >>
rect 246 140 247 141 
<< pdiffusion >>
rect 247 140 248 141 
<< pdiffusion >>
rect 248 140 249 141 
<< pdiffusion >>
rect 249 140 250 141 
<< pdiffusion >>
rect 250 140 251 141 
<< pdiffusion >>
rect 251 140 252 141 
<< m1 >>
rect 253 140 254 141 
<< m2 >>
rect 254 140 255 141 
<< pdiffusion >>
rect 264 140 265 141 
<< pdiffusion >>
rect 265 140 266 141 
<< pdiffusion >>
rect 266 140 267 141 
<< pdiffusion >>
rect 267 140 268 141 
<< pdiffusion >>
rect 268 140 269 141 
<< pdiffusion >>
rect 269 140 270 141 
<< pdiffusion >>
rect 282 140 283 141 
<< pdiffusion >>
rect 283 140 284 141 
<< pdiffusion >>
rect 284 140 285 141 
<< pdiffusion >>
rect 285 140 286 141 
<< pdiffusion >>
rect 286 140 287 141 
<< pdiffusion >>
rect 287 140 288 141 
<< pdiffusion >>
rect 300 140 301 141 
<< pdiffusion >>
rect 301 140 302 141 
<< pdiffusion >>
rect 302 140 303 141 
<< pdiffusion >>
rect 303 140 304 141 
<< pdiffusion >>
rect 304 140 305 141 
<< pdiffusion >>
rect 305 140 306 141 
<< m1 >>
rect 307 140 308 141 
<< m1 >>
rect 311 140 312 141 
<< pdiffusion >>
rect 318 140 319 141 
<< pdiffusion >>
rect 319 140 320 141 
<< pdiffusion >>
rect 320 140 321 141 
<< pdiffusion >>
rect 321 140 322 141 
<< pdiffusion >>
rect 322 140 323 141 
<< pdiffusion >>
rect 323 140 324 141 
<< pdiffusion >>
rect 336 140 337 141 
<< pdiffusion >>
rect 337 140 338 141 
<< pdiffusion >>
rect 338 140 339 141 
<< pdiffusion >>
rect 339 140 340 141 
<< pdiffusion >>
rect 340 140 341 141 
<< pdiffusion >>
rect 341 140 342 141 
<< m1 >>
rect 343 140 344 141 
<< pdiffusion >>
rect 354 140 355 141 
<< pdiffusion >>
rect 355 140 356 141 
<< pdiffusion >>
rect 356 140 357 141 
<< pdiffusion >>
rect 357 140 358 141 
<< pdiffusion >>
rect 358 140 359 141 
<< pdiffusion >>
rect 359 140 360 141 
<< pdiffusion >>
rect 372 140 373 141 
<< pdiffusion >>
rect 373 140 374 141 
<< pdiffusion >>
rect 374 140 375 141 
<< pdiffusion >>
rect 375 140 376 141 
<< pdiffusion >>
rect 376 140 377 141 
<< pdiffusion >>
rect 377 140 378 141 
<< m1 >>
rect 406 140 407 141 
<< pdiffusion >>
rect 408 140 409 141 
<< pdiffusion >>
rect 409 140 410 141 
<< pdiffusion >>
rect 410 140 411 141 
<< pdiffusion >>
rect 411 140 412 141 
<< pdiffusion >>
rect 412 140 413 141 
<< pdiffusion >>
rect 413 140 414 141 
<< pdiffusion >>
rect 426 140 427 141 
<< pdiffusion >>
rect 427 140 428 141 
<< pdiffusion >>
rect 428 140 429 141 
<< pdiffusion >>
rect 429 140 430 141 
<< pdiffusion >>
rect 430 140 431 141 
<< pdiffusion >>
rect 431 140 432 141 
<< pdiffusion >>
rect 444 140 445 141 
<< pdiffusion >>
rect 445 140 446 141 
<< pdiffusion >>
rect 446 140 447 141 
<< pdiffusion >>
rect 447 140 448 141 
<< pdiffusion >>
rect 448 140 449 141 
<< pdiffusion >>
rect 449 140 450 141 
<< pdiffusion >>
rect 12 141 13 142 
<< pdiffusion >>
rect 13 141 14 142 
<< pdiffusion >>
rect 14 141 15 142 
<< pdiffusion >>
rect 15 141 16 142 
<< pdiffusion >>
rect 16 141 17 142 
<< pdiffusion >>
rect 17 141 18 142 
<< m1 >>
rect 28 141 29 142 
<< pdiffusion >>
rect 30 141 31 142 
<< pdiffusion >>
rect 31 141 32 142 
<< pdiffusion >>
rect 32 141 33 142 
<< pdiffusion >>
rect 33 141 34 142 
<< pdiffusion >>
rect 34 141 35 142 
<< pdiffusion >>
rect 35 141 36 142 
<< pdiffusion >>
rect 48 141 49 142 
<< pdiffusion >>
rect 49 141 50 142 
<< pdiffusion >>
rect 50 141 51 142 
<< pdiffusion >>
rect 51 141 52 142 
<< pdiffusion >>
rect 52 141 53 142 
<< pdiffusion >>
rect 53 141 54 142 
<< m1 >>
rect 64 141 65 142 
<< pdiffusion >>
rect 66 141 67 142 
<< pdiffusion >>
rect 67 141 68 142 
<< pdiffusion >>
rect 68 141 69 142 
<< pdiffusion >>
rect 69 141 70 142 
<< pdiffusion >>
rect 70 141 71 142 
<< pdiffusion >>
rect 71 141 72 142 
<< pdiffusion >>
rect 84 141 85 142 
<< pdiffusion >>
rect 85 141 86 142 
<< pdiffusion >>
rect 86 141 87 142 
<< pdiffusion >>
rect 87 141 88 142 
<< pdiffusion >>
rect 88 141 89 142 
<< pdiffusion >>
rect 89 141 90 142 
<< m1 >>
rect 93 141 94 142 
<< m1 >>
rect 95 141 96 142 
<< pdiffusion >>
rect 102 141 103 142 
<< pdiffusion >>
rect 103 141 104 142 
<< pdiffusion >>
rect 104 141 105 142 
<< pdiffusion >>
rect 105 141 106 142 
<< pdiffusion >>
rect 106 141 107 142 
<< pdiffusion >>
rect 107 141 108 142 
<< m1 >>
rect 116 141 117 142 
<< m1 >>
rect 118 141 119 142 
<< pdiffusion >>
rect 120 141 121 142 
<< pdiffusion >>
rect 121 141 122 142 
<< pdiffusion >>
rect 122 141 123 142 
<< pdiffusion >>
rect 123 141 124 142 
<< pdiffusion >>
rect 124 141 125 142 
<< pdiffusion >>
rect 125 141 126 142 
<< m1 >>
rect 145 141 146 142 
<< pdiffusion >>
rect 156 141 157 142 
<< pdiffusion >>
rect 157 141 158 142 
<< pdiffusion >>
rect 158 141 159 142 
<< pdiffusion >>
rect 159 141 160 142 
<< pdiffusion >>
rect 160 141 161 142 
<< pdiffusion >>
rect 161 141 162 142 
<< m1 >>
rect 170 141 171 142 
<< m1 >>
rect 172 141 173 142 
<< pdiffusion >>
rect 174 141 175 142 
<< pdiffusion >>
rect 175 141 176 142 
<< pdiffusion >>
rect 176 141 177 142 
<< pdiffusion >>
rect 177 141 178 142 
<< pdiffusion >>
rect 178 141 179 142 
<< pdiffusion >>
rect 179 141 180 142 
<< pdiffusion >>
rect 192 141 193 142 
<< pdiffusion >>
rect 193 141 194 142 
<< pdiffusion >>
rect 194 141 195 142 
<< pdiffusion >>
rect 195 141 196 142 
<< pdiffusion >>
rect 196 141 197 142 
<< pdiffusion >>
rect 197 141 198 142 
<< m1 >>
rect 208 141 209 142 
<< pdiffusion >>
rect 210 141 211 142 
<< pdiffusion >>
rect 211 141 212 142 
<< pdiffusion >>
rect 212 141 213 142 
<< pdiffusion >>
rect 213 141 214 142 
<< pdiffusion >>
rect 214 141 215 142 
<< pdiffusion >>
rect 215 141 216 142 
<< m2 >>
rect 225 141 226 142 
<< m1 >>
rect 226 141 227 142 
<< pdiffusion >>
rect 228 141 229 142 
<< pdiffusion >>
rect 229 141 230 142 
<< pdiffusion >>
rect 230 141 231 142 
<< pdiffusion >>
rect 231 141 232 142 
<< pdiffusion >>
rect 232 141 233 142 
<< pdiffusion >>
rect 233 141 234 142 
<< m1 >>
rect 244 141 245 142 
<< pdiffusion >>
rect 246 141 247 142 
<< pdiffusion >>
rect 247 141 248 142 
<< pdiffusion >>
rect 248 141 249 142 
<< pdiffusion >>
rect 249 141 250 142 
<< pdiffusion >>
rect 250 141 251 142 
<< pdiffusion >>
rect 251 141 252 142 
<< m1 >>
rect 253 141 254 142 
<< m2 >>
rect 254 141 255 142 
<< pdiffusion >>
rect 264 141 265 142 
<< pdiffusion >>
rect 265 141 266 142 
<< pdiffusion >>
rect 266 141 267 142 
<< pdiffusion >>
rect 267 141 268 142 
<< pdiffusion >>
rect 268 141 269 142 
<< pdiffusion >>
rect 269 141 270 142 
<< pdiffusion >>
rect 282 141 283 142 
<< pdiffusion >>
rect 283 141 284 142 
<< pdiffusion >>
rect 284 141 285 142 
<< pdiffusion >>
rect 285 141 286 142 
<< pdiffusion >>
rect 286 141 287 142 
<< pdiffusion >>
rect 287 141 288 142 
<< pdiffusion >>
rect 300 141 301 142 
<< pdiffusion >>
rect 301 141 302 142 
<< pdiffusion >>
rect 302 141 303 142 
<< pdiffusion >>
rect 303 141 304 142 
<< pdiffusion >>
rect 304 141 305 142 
<< pdiffusion >>
rect 305 141 306 142 
<< m1 >>
rect 307 141 308 142 
<< m1 >>
rect 311 141 312 142 
<< pdiffusion >>
rect 318 141 319 142 
<< pdiffusion >>
rect 319 141 320 142 
<< pdiffusion >>
rect 320 141 321 142 
<< pdiffusion >>
rect 321 141 322 142 
<< pdiffusion >>
rect 322 141 323 142 
<< pdiffusion >>
rect 323 141 324 142 
<< pdiffusion >>
rect 336 141 337 142 
<< pdiffusion >>
rect 337 141 338 142 
<< pdiffusion >>
rect 338 141 339 142 
<< pdiffusion >>
rect 339 141 340 142 
<< pdiffusion >>
rect 340 141 341 142 
<< pdiffusion >>
rect 341 141 342 142 
<< m1 >>
rect 343 141 344 142 
<< pdiffusion >>
rect 354 141 355 142 
<< pdiffusion >>
rect 355 141 356 142 
<< pdiffusion >>
rect 356 141 357 142 
<< pdiffusion >>
rect 357 141 358 142 
<< pdiffusion >>
rect 358 141 359 142 
<< pdiffusion >>
rect 359 141 360 142 
<< pdiffusion >>
rect 372 141 373 142 
<< pdiffusion >>
rect 373 141 374 142 
<< pdiffusion >>
rect 374 141 375 142 
<< pdiffusion >>
rect 375 141 376 142 
<< pdiffusion >>
rect 376 141 377 142 
<< pdiffusion >>
rect 377 141 378 142 
<< m1 >>
rect 406 141 407 142 
<< pdiffusion >>
rect 408 141 409 142 
<< pdiffusion >>
rect 409 141 410 142 
<< pdiffusion >>
rect 410 141 411 142 
<< pdiffusion >>
rect 411 141 412 142 
<< pdiffusion >>
rect 412 141 413 142 
<< pdiffusion >>
rect 413 141 414 142 
<< pdiffusion >>
rect 426 141 427 142 
<< pdiffusion >>
rect 427 141 428 142 
<< pdiffusion >>
rect 428 141 429 142 
<< pdiffusion >>
rect 429 141 430 142 
<< pdiffusion >>
rect 430 141 431 142 
<< pdiffusion >>
rect 431 141 432 142 
<< pdiffusion >>
rect 444 141 445 142 
<< pdiffusion >>
rect 445 141 446 142 
<< pdiffusion >>
rect 446 141 447 142 
<< pdiffusion >>
rect 447 141 448 142 
<< pdiffusion >>
rect 448 141 449 142 
<< pdiffusion >>
rect 449 141 450 142 
<< pdiffusion >>
rect 12 142 13 143 
<< pdiffusion >>
rect 13 142 14 143 
<< pdiffusion >>
rect 14 142 15 143 
<< pdiffusion >>
rect 15 142 16 143 
<< pdiffusion >>
rect 16 142 17 143 
<< pdiffusion >>
rect 17 142 18 143 
<< m1 >>
rect 28 142 29 143 
<< pdiffusion >>
rect 30 142 31 143 
<< pdiffusion >>
rect 31 142 32 143 
<< pdiffusion >>
rect 32 142 33 143 
<< pdiffusion >>
rect 33 142 34 143 
<< pdiffusion >>
rect 34 142 35 143 
<< pdiffusion >>
rect 35 142 36 143 
<< pdiffusion >>
rect 48 142 49 143 
<< pdiffusion >>
rect 49 142 50 143 
<< pdiffusion >>
rect 50 142 51 143 
<< pdiffusion >>
rect 51 142 52 143 
<< pdiffusion >>
rect 52 142 53 143 
<< pdiffusion >>
rect 53 142 54 143 
<< m1 >>
rect 64 142 65 143 
<< pdiffusion >>
rect 66 142 67 143 
<< pdiffusion >>
rect 67 142 68 143 
<< pdiffusion >>
rect 68 142 69 143 
<< pdiffusion >>
rect 69 142 70 143 
<< pdiffusion >>
rect 70 142 71 143 
<< pdiffusion >>
rect 71 142 72 143 
<< pdiffusion >>
rect 84 142 85 143 
<< pdiffusion >>
rect 85 142 86 143 
<< pdiffusion >>
rect 86 142 87 143 
<< pdiffusion >>
rect 87 142 88 143 
<< pdiffusion >>
rect 88 142 89 143 
<< pdiffusion >>
rect 89 142 90 143 
<< m1 >>
rect 93 142 94 143 
<< m1 >>
rect 95 142 96 143 
<< pdiffusion >>
rect 102 142 103 143 
<< pdiffusion >>
rect 103 142 104 143 
<< pdiffusion >>
rect 104 142 105 143 
<< pdiffusion >>
rect 105 142 106 143 
<< pdiffusion >>
rect 106 142 107 143 
<< pdiffusion >>
rect 107 142 108 143 
<< m1 >>
rect 116 142 117 143 
<< m1 >>
rect 118 142 119 143 
<< pdiffusion >>
rect 120 142 121 143 
<< pdiffusion >>
rect 121 142 122 143 
<< pdiffusion >>
rect 122 142 123 143 
<< pdiffusion >>
rect 123 142 124 143 
<< pdiffusion >>
rect 124 142 125 143 
<< pdiffusion >>
rect 125 142 126 143 
<< m1 >>
rect 145 142 146 143 
<< pdiffusion >>
rect 156 142 157 143 
<< pdiffusion >>
rect 157 142 158 143 
<< pdiffusion >>
rect 158 142 159 143 
<< pdiffusion >>
rect 159 142 160 143 
<< pdiffusion >>
rect 160 142 161 143 
<< pdiffusion >>
rect 161 142 162 143 
<< m1 >>
rect 170 142 171 143 
<< m1 >>
rect 172 142 173 143 
<< pdiffusion >>
rect 174 142 175 143 
<< pdiffusion >>
rect 175 142 176 143 
<< pdiffusion >>
rect 176 142 177 143 
<< pdiffusion >>
rect 177 142 178 143 
<< pdiffusion >>
rect 178 142 179 143 
<< pdiffusion >>
rect 179 142 180 143 
<< pdiffusion >>
rect 192 142 193 143 
<< pdiffusion >>
rect 193 142 194 143 
<< pdiffusion >>
rect 194 142 195 143 
<< pdiffusion >>
rect 195 142 196 143 
<< pdiffusion >>
rect 196 142 197 143 
<< pdiffusion >>
rect 197 142 198 143 
<< m1 >>
rect 208 142 209 143 
<< pdiffusion >>
rect 210 142 211 143 
<< pdiffusion >>
rect 211 142 212 143 
<< pdiffusion >>
rect 212 142 213 143 
<< pdiffusion >>
rect 213 142 214 143 
<< pdiffusion >>
rect 214 142 215 143 
<< pdiffusion >>
rect 215 142 216 143 
<< m2 >>
rect 225 142 226 143 
<< m1 >>
rect 226 142 227 143 
<< pdiffusion >>
rect 228 142 229 143 
<< pdiffusion >>
rect 229 142 230 143 
<< pdiffusion >>
rect 230 142 231 143 
<< pdiffusion >>
rect 231 142 232 143 
<< pdiffusion >>
rect 232 142 233 143 
<< pdiffusion >>
rect 233 142 234 143 
<< m1 >>
rect 244 142 245 143 
<< pdiffusion >>
rect 246 142 247 143 
<< pdiffusion >>
rect 247 142 248 143 
<< pdiffusion >>
rect 248 142 249 143 
<< pdiffusion >>
rect 249 142 250 143 
<< pdiffusion >>
rect 250 142 251 143 
<< pdiffusion >>
rect 251 142 252 143 
<< m1 >>
rect 253 142 254 143 
<< m2 >>
rect 254 142 255 143 
<< pdiffusion >>
rect 264 142 265 143 
<< pdiffusion >>
rect 265 142 266 143 
<< pdiffusion >>
rect 266 142 267 143 
<< pdiffusion >>
rect 267 142 268 143 
<< pdiffusion >>
rect 268 142 269 143 
<< pdiffusion >>
rect 269 142 270 143 
<< pdiffusion >>
rect 282 142 283 143 
<< pdiffusion >>
rect 283 142 284 143 
<< pdiffusion >>
rect 284 142 285 143 
<< pdiffusion >>
rect 285 142 286 143 
<< pdiffusion >>
rect 286 142 287 143 
<< pdiffusion >>
rect 287 142 288 143 
<< pdiffusion >>
rect 300 142 301 143 
<< pdiffusion >>
rect 301 142 302 143 
<< pdiffusion >>
rect 302 142 303 143 
<< pdiffusion >>
rect 303 142 304 143 
<< pdiffusion >>
rect 304 142 305 143 
<< pdiffusion >>
rect 305 142 306 143 
<< m1 >>
rect 307 142 308 143 
<< m1 >>
rect 311 142 312 143 
<< pdiffusion >>
rect 318 142 319 143 
<< pdiffusion >>
rect 319 142 320 143 
<< pdiffusion >>
rect 320 142 321 143 
<< pdiffusion >>
rect 321 142 322 143 
<< pdiffusion >>
rect 322 142 323 143 
<< pdiffusion >>
rect 323 142 324 143 
<< pdiffusion >>
rect 336 142 337 143 
<< pdiffusion >>
rect 337 142 338 143 
<< pdiffusion >>
rect 338 142 339 143 
<< pdiffusion >>
rect 339 142 340 143 
<< pdiffusion >>
rect 340 142 341 143 
<< pdiffusion >>
rect 341 142 342 143 
<< m1 >>
rect 343 142 344 143 
<< pdiffusion >>
rect 354 142 355 143 
<< pdiffusion >>
rect 355 142 356 143 
<< pdiffusion >>
rect 356 142 357 143 
<< pdiffusion >>
rect 357 142 358 143 
<< pdiffusion >>
rect 358 142 359 143 
<< pdiffusion >>
rect 359 142 360 143 
<< pdiffusion >>
rect 372 142 373 143 
<< pdiffusion >>
rect 373 142 374 143 
<< pdiffusion >>
rect 374 142 375 143 
<< pdiffusion >>
rect 375 142 376 143 
<< pdiffusion >>
rect 376 142 377 143 
<< pdiffusion >>
rect 377 142 378 143 
<< m1 >>
rect 406 142 407 143 
<< pdiffusion >>
rect 408 142 409 143 
<< pdiffusion >>
rect 409 142 410 143 
<< pdiffusion >>
rect 410 142 411 143 
<< pdiffusion >>
rect 411 142 412 143 
<< pdiffusion >>
rect 412 142 413 143 
<< pdiffusion >>
rect 413 142 414 143 
<< pdiffusion >>
rect 426 142 427 143 
<< pdiffusion >>
rect 427 142 428 143 
<< pdiffusion >>
rect 428 142 429 143 
<< pdiffusion >>
rect 429 142 430 143 
<< pdiffusion >>
rect 430 142 431 143 
<< pdiffusion >>
rect 431 142 432 143 
<< pdiffusion >>
rect 444 142 445 143 
<< pdiffusion >>
rect 445 142 446 143 
<< pdiffusion >>
rect 446 142 447 143 
<< pdiffusion >>
rect 447 142 448 143 
<< pdiffusion >>
rect 448 142 449 143 
<< pdiffusion >>
rect 449 142 450 143 
<< pdiffusion >>
rect 12 143 13 144 
<< pdiffusion >>
rect 13 143 14 144 
<< pdiffusion >>
rect 14 143 15 144 
<< pdiffusion >>
rect 15 143 16 144 
<< m1 >>
rect 16 143 17 144 
<< pdiffusion >>
rect 16 143 17 144 
<< pdiffusion >>
rect 17 143 18 144 
<< m1 >>
rect 28 143 29 144 
<< pdiffusion >>
rect 30 143 31 144 
<< pdiffusion >>
rect 31 143 32 144 
<< pdiffusion >>
rect 32 143 33 144 
<< pdiffusion >>
rect 33 143 34 144 
<< pdiffusion >>
rect 34 143 35 144 
<< pdiffusion >>
rect 35 143 36 144 
<< pdiffusion >>
rect 48 143 49 144 
<< pdiffusion >>
rect 49 143 50 144 
<< pdiffusion >>
rect 50 143 51 144 
<< pdiffusion >>
rect 51 143 52 144 
<< pdiffusion >>
rect 52 143 53 144 
<< pdiffusion >>
rect 53 143 54 144 
<< m1 >>
rect 64 143 65 144 
<< pdiffusion >>
rect 66 143 67 144 
<< pdiffusion >>
rect 67 143 68 144 
<< pdiffusion >>
rect 68 143 69 144 
<< pdiffusion >>
rect 69 143 70 144 
<< pdiffusion >>
rect 70 143 71 144 
<< pdiffusion >>
rect 71 143 72 144 
<< pdiffusion >>
rect 84 143 85 144 
<< pdiffusion >>
rect 85 143 86 144 
<< pdiffusion >>
rect 86 143 87 144 
<< pdiffusion >>
rect 87 143 88 144 
<< pdiffusion >>
rect 88 143 89 144 
<< pdiffusion >>
rect 89 143 90 144 
<< m1 >>
rect 93 143 94 144 
<< m1 >>
rect 95 143 96 144 
<< pdiffusion >>
rect 102 143 103 144 
<< m1 >>
rect 103 143 104 144 
<< pdiffusion >>
rect 103 143 104 144 
<< pdiffusion >>
rect 104 143 105 144 
<< pdiffusion >>
rect 105 143 106 144 
<< pdiffusion >>
rect 106 143 107 144 
<< pdiffusion >>
rect 107 143 108 144 
<< m1 >>
rect 116 143 117 144 
<< m1 >>
rect 118 143 119 144 
<< pdiffusion >>
rect 120 143 121 144 
<< pdiffusion >>
rect 121 143 122 144 
<< pdiffusion >>
rect 122 143 123 144 
<< pdiffusion >>
rect 123 143 124 144 
<< pdiffusion >>
rect 124 143 125 144 
<< pdiffusion >>
rect 125 143 126 144 
<< m1 >>
rect 145 143 146 144 
<< pdiffusion >>
rect 156 143 157 144 
<< pdiffusion >>
rect 157 143 158 144 
<< pdiffusion >>
rect 158 143 159 144 
<< pdiffusion >>
rect 159 143 160 144 
<< pdiffusion >>
rect 160 143 161 144 
<< pdiffusion >>
rect 161 143 162 144 
<< m1 >>
rect 170 143 171 144 
<< m1 >>
rect 172 143 173 144 
<< pdiffusion >>
rect 174 143 175 144 
<< pdiffusion >>
rect 175 143 176 144 
<< pdiffusion >>
rect 176 143 177 144 
<< pdiffusion >>
rect 177 143 178 144 
<< pdiffusion >>
rect 178 143 179 144 
<< pdiffusion >>
rect 179 143 180 144 
<< pdiffusion >>
rect 192 143 193 144 
<< pdiffusion >>
rect 193 143 194 144 
<< pdiffusion >>
rect 194 143 195 144 
<< pdiffusion >>
rect 195 143 196 144 
<< pdiffusion >>
rect 196 143 197 144 
<< pdiffusion >>
rect 197 143 198 144 
<< m1 >>
rect 208 143 209 144 
<< pdiffusion >>
rect 210 143 211 144 
<< pdiffusion >>
rect 211 143 212 144 
<< pdiffusion >>
rect 212 143 213 144 
<< pdiffusion >>
rect 213 143 214 144 
<< pdiffusion >>
rect 214 143 215 144 
<< pdiffusion >>
rect 215 143 216 144 
<< m2 >>
rect 225 143 226 144 
<< m1 >>
rect 226 143 227 144 
<< pdiffusion >>
rect 228 143 229 144 
<< m1 >>
rect 229 143 230 144 
<< pdiffusion >>
rect 229 143 230 144 
<< pdiffusion >>
rect 230 143 231 144 
<< pdiffusion >>
rect 231 143 232 144 
<< pdiffusion >>
rect 232 143 233 144 
<< pdiffusion >>
rect 233 143 234 144 
<< m1 >>
rect 244 143 245 144 
<< pdiffusion >>
rect 246 143 247 144 
<< pdiffusion >>
rect 247 143 248 144 
<< pdiffusion >>
rect 248 143 249 144 
<< pdiffusion >>
rect 249 143 250 144 
<< pdiffusion >>
rect 250 143 251 144 
<< pdiffusion >>
rect 251 143 252 144 
<< m1 >>
rect 253 143 254 144 
<< m2 >>
rect 254 143 255 144 
<< pdiffusion >>
rect 264 143 265 144 
<< pdiffusion >>
rect 265 143 266 144 
<< pdiffusion >>
rect 266 143 267 144 
<< pdiffusion >>
rect 267 143 268 144 
<< pdiffusion >>
rect 268 143 269 144 
<< pdiffusion >>
rect 269 143 270 144 
<< pdiffusion >>
rect 282 143 283 144 
<< pdiffusion >>
rect 283 143 284 144 
<< pdiffusion >>
rect 284 143 285 144 
<< pdiffusion >>
rect 285 143 286 144 
<< pdiffusion >>
rect 286 143 287 144 
<< pdiffusion >>
rect 287 143 288 144 
<< pdiffusion >>
rect 300 143 301 144 
<< pdiffusion >>
rect 301 143 302 144 
<< pdiffusion >>
rect 302 143 303 144 
<< pdiffusion >>
rect 303 143 304 144 
<< m1 >>
rect 304 143 305 144 
<< pdiffusion >>
rect 304 143 305 144 
<< pdiffusion >>
rect 305 143 306 144 
<< m1 >>
rect 307 143 308 144 
<< m1 >>
rect 311 143 312 144 
<< pdiffusion >>
rect 318 143 319 144 
<< m1 >>
rect 319 143 320 144 
<< pdiffusion >>
rect 319 143 320 144 
<< pdiffusion >>
rect 320 143 321 144 
<< pdiffusion >>
rect 321 143 322 144 
<< m1 >>
rect 322 143 323 144 
<< pdiffusion >>
rect 322 143 323 144 
<< pdiffusion >>
rect 323 143 324 144 
<< pdiffusion >>
rect 336 143 337 144 
<< pdiffusion >>
rect 337 143 338 144 
<< pdiffusion >>
rect 338 143 339 144 
<< pdiffusion >>
rect 339 143 340 144 
<< pdiffusion >>
rect 340 143 341 144 
<< pdiffusion >>
rect 341 143 342 144 
<< m1 >>
rect 343 143 344 144 
<< pdiffusion >>
rect 354 143 355 144 
<< pdiffusion >>
rect 355 143 356 144 
<< pdiffusion >>
rect 356 143 357 144 
<< pdiffusion >>
rect 357 143 358 144 
<< pdiffusion >>
rect 358 143 359 144 
<< pdiffusion >>
rect 359 143 360 144 
<< pdiffusion >>
rect 372 143 373 144 
<< pdiffusion >>
rect 373 143 374 144 
<< pdiffusion >>
rect 374 143 375 144 
<< pdiffusion >>
rect 375 143 376 144 
<< pdiffusion >>
rect 376 143 377 144 
<< pdiffusion >>
rect 377 143 378 144 
<< m1 >>
rect 406 143 407 144 
<< pdiffusion >>
rect 408 143 409 144 
<< pdiffusion >>
rect 409 143 410 144 
<< pdiffusion >>
rect 410 143 411 144 
<< pdiffusion >>
rect 411 143 412 144 
<< pdiffusion >>
rect 412 143 413 144 
<< pdiffusion >>
rect 413 143 414 144 
<< pdiffusion >>
rect 426 143 427 144 
<< pdiffusion >>
rect 427 143 428 144 
<< pdiffusion >>
rect 428 143 429 144 
<< pdiffusion >>
rect 429 143 430 144 
<< pdiffusion >>
rect 430 143 431 144 
<< pdiffusion >>
rect 431 143 432 144 
<< pdiffusion >>
rect 444 143 445 144 
<< pdiffusion >>
rect 445 143 446 144 
<< pdiffusion >>
rect 446 143 447 144 
<< pdiffusion >>
rect 447 143 448 144 
<< pdiffusion >>
rect 448 143 449 144 
<< pdiffusion >>
rect 449 143 450 144 
<< m1 >>
rect 16 144 17 145 
<< m1 >>
rect 28 144 29 145 
<< m1 >>
rect 64 144 65 145 
<< m1 >>
rect 93 144 94 145 
<< m1 >>
rect 95 144 96 145 
<< m1 >>
rect 103 144 104 145 
<< m1 >>
rect 116 144 117 145 
<< m2 >>
rect 116 144 117 145 
<< m2c >>
rect 116 144 117 145 
<< m1 >>
rect 116 144 117 145 
<< m2 >>
rect 116 144 117 145 
<< m2 >>
rect 117 144 118 145 
<< m1 >>
rect 118 144 119 145 
<< m2 >>
rect 118 144 119 145 
<< m1 >>
rect 145 144 146 145 
<< m1 >>
rect 170 144 171 145 
<< m1 >>
rect 172 144 173 145 
<< m1 >>
rect 208 144 209 145 
<< m2 >>
rect 225 144 226 145 
<< m1 >>
rect 226 144 227 145 
<< m1 >>
rect 229 144 230 145 
<< m1 >>
rect 244 144 245 145 
<< m1 >>
rect 253 144 254 145 
<< m2 >>
rect 254 144 255 145 
<< m1 >>
rect 304 144 305 145 
<< m1 >>
rect 307 144 308 145 
<< m1 >>
rect 311 144 312 145 
<< m1 >>
rect 319 144 320 145 
<< m1 >>
rect 322 144 323 145 
<< m1 >>
rect 343 144 344 145 
<< m1 >>
rect 406 144 407 145 
<< m1 >>
rect 16 145 17 146 
<< m1 >>
rect 17 145 18 146 
<< m1 >>
rect 18 145 19 146 
<< m1 >>
rect 19 145 20 146 
<< m1 >>
rect 20 145 21 146 
<< m1 >>
rect 21 145 22 146 
<< m1 >>
rect 22 145 23 146 
<< m1 >>
rect 23 145 24 146 
<< m1 >>
rect 24 145 25 146 
<< m1 >>
rect 25 145 26 146 
<< m1 >>
rect 26 145 27 146 
<< m1 >>
rect 27 145 28 146 
<< m1 >>
rect 28 145 29 146 
<< m1 >>
rect 64 145 65 146 
<< m1 >>
rect 93 145 94 146 
<< m1 >>
rect 95 145 96 146 
<< m1 >>
rect 103 145 104 146 
<< m1 >>
rect 118 145 119 146 
<< m2 >>
rect 118 145 119 146 
<< m1 >>
rect 145 145 146 146 
<< m1 >>
rect 170 145 171 146 
<< m1 >>
rect 172 145 173 146 
<< m1 >>
rect 208 145 209 146 
<< m2 >>
rect 225 145 226 146 
<< m1 >>
rect 226 145 227 146 
<< m1 >>
rect 229 145 230 146 
<< m1 >>
rect 244 145 245 146 
<< m1 >>
rect 253 145 254 146 
<< m2 >>
rect 254 145 255 146 
<< m1 >>
rect 304 145 305 146 
<< m1 >>
rect 305 145 306 146 
<< m2 >>
rect 305 145 306 146 
<< m2c >>
rect 305 145 306 146 
<< m1 >>
rect 305 145 306 146 
<< m2 >>
rect 305 145 306 146 
<< m2 >>
rect 306 145 307 146 
<< m1 >>
rect 307 145 308 146 
<< m2 >>
rect 307 145 308 146 
<< m2 >>
rect 308 145 309 146 
<< m1 >>
rect 309 145 310 146 
<< m2 >>
rect 309 145 310 146 
<< m2c >>
rect 309 145 310 146 
<< m1 >>
rect 309 145 310 146 
<< m2 >>
rect 309 145 310 146 
<< m2 >>
rect 310 145 311 146 
<< m1 >>
rect 311 145 312 146 
<< m2 >>
rect 311 145 312 146 
<< m2 >>
rect 312 145 313 146 
<< m1 >>
rect 313 145 314 146 
<< m2 >>
rect 313 145 314 146 
<< m2c >>
rect 313 145 314 146 
<< m1 >>
rect 313 145 314 146 
<< m2 >>
rect 313 145 314 146 
<< m1 >>
rect 314 145 315 146 
<< m1 >>
rect 315 145 316 146 
<< m1 >>
rect 316 145 317 146 
<< m1 >>
rect 317 145 318 146 
<< m1 >>
rect 318 145 319 146 
<< m1 >>
rect 319 145 320 146 
<< m1 >>
rect 322 145 323 146 
<< m1 >>
rect 343 145 344 146 
<< m1 >>
rect 406 145 407 146 
<< m1 >>
rect 64 146 65 147 
<< m1 >>
rect 93 146 94 147 
<< m1 >>
rect 95 146 96 147 
<< m1 >>
rect 103 146 104 147 
<< m1 >>
rect 104 146 105 147 
<< m1 >>
rect 105 146 106 147 
<< m1 >>
rect 106 146 107 147 
<< m1 >>
rect 107 146 108 147 
<< m1 >>
rect 108 146 109 147 
<< m1 >>
rect 109 146 110 147 
<< m1 >>
rect 110 146 111 147 
<< m1 >>
rect 111 146 112 147 
<< m1 >>
rect 112 146 113 147 
<< m1 >>
rect 113 146 114 147 
<< m1 >>
rect 114 146 115 147 
<< m1 >>
rect 115 146 116 147 
<< m1 >>
rect 116 146 117 147 
<< m1 >>
rect 117 146 118 147 
<< m1 >>
rect 118 146 119 147 
<< m2 >>
rect 118 146 119 147 
<< m1 >>
rect 145 146 146 147 
<< m1 >>
rect 170 146 171 147 
<< m1 >>
rect 172 146 173 147 
<< m1 >>
rect 208 146 209 147 
<< m2 >>
rect 225 146 226 147 
<< m1 >>
rect 226 146 227 147 
<< m1 >>
rect 229 146 230 147 
<< m1 >>
rect 230 146 231 147 
<< m1 >>
rect 231 146 232 147 
<< m1 >>
rect 232 146 233 147 
<< m1 >>
rect 233 146 234 147 
<< m1 >>
rect 234 146 235 147 
<< m1 >>
rect 235 146 236 147 
<< m1 >>
rect 236 146 237 147 
<< m1 >>
rect 237 146 238 147 
<< m1 >>
rect 238 146 239 147 
<< m1 >>
rect 239 146 240 147 
<< m1 >>
rect 240 146 241 147 
<< m1 >>
rect 241 146 242 147 
<< m1 >>
rect 242 146 243 147 
<< m1 >>
rect 243 146 244 147 
<< m1 >>
rect 244 146 245 147 
<< m1 >>
rect 253 146 254 147 
<< m2 >>
rect 254 146 255 147 
<< m1 >>
rect 307 146 308 147 
<< m1 >>
rect 311 146 312 147 
<< m1 >>
rect 322 146 323 147 
<< m1 >>
rect 343 146 344 147 
<< m1 >>
rect 406 146 407 147 
<< m1 >>
rect 64 147 65 148 
<< m1 >>
rect 93 147 94 148 
<< m1 >>
rect 95 147 96 148 
<< m2 >>
rect 118 147 119 148 
<< m1 >>
rect 145 147 146 148 
<< m1 >>
rect 170 147 171 148 
<< m1 >>
rect 172 147 173 148 
<< m1 >>
rect 208 147 209 148 
<< m2 >>
rect 225 147 226 148 
<< m1 >>
rect 226 147 227 148 
<< m1 >>
rect 253 147 254 148 
<< m2 >>
rect 254 147 255 148 
<< m1 >>
rect 307 147 308 148 
<< m1 >>
rect 311 147 312 148 
<< m1 >>
rect 322 147 323 148 
<< m1 >>
rect 343 147 344 148 
<< m1 >>
rect 406 147 407 148 
<< m1 >>
rect 64 148 65 149 
<< m1 >>
rect 93 148 94 149 
<< m1 >>
rect 95 148 96 149 
<< m1 >>
rect 118 148 119 149 
<< m2 >>
rect 118 148 119 149 
<< m2c >>
rect 118 148 119 149 
<< m1 >>
rect 118 148 119 149 
<< m2 >>
rect 118 148 119 149 
<< m1 >>
rect 145 148 146 149 
<< m1 >>
rect 146 148 147 149 
<< m1 >>
rect 147 148 148 149 
<< m1 >>
rect 148 148 149 149 
<< m1 >>
rect 149 148 150 149 
<< m1 >>
rect 150 148 151 149 
<< m1 >>
rect 151 148 152 149 
<< m1 >>
rect 152 148 153 149 
<< m1 >>
rect 153 148 154 149 
<< m1 >>
rect 154 148 155 149 
<< m1 >>
rect 155 148 156 149 
<< m1 >>
rect 156 148 157 149 
<< m1 >>
rect 157 148 158 149 
<< m1 >>
rect 170 148 171 149 
<< m1 >>
rect 172 148 173 149 
<< m1 >>
rect 173 148 174 149 
<< m1 >>
rect 174 148 175 149 
<< m1 >>
rect 175 148 176 149 
<< m1 >>
rect 176 148 177 149 
<< m1 >>
rect 177 148 178 149 
<< m1 >>
rect 178 148 179 149 
<< m1 >>
rect 208 148 209 149 
<< m2 >>
rect 225 148 226 149 
<< m1 >>
rect 226 148 227 149 
<< m2 >>
rect 226 148 227 149 
<< m2 >>
rect 227 148 228 149 
<< m1 >>
rect 228 148 229 149 
<< m2 >>
rect 228 148 229 149 
<< m2c >>
rect 228 148 229 149 
<< m1 >>
rect 228 148 229 149 
<< m2 >>
rect 228 148 229 149 
<< m1 >>
rect 229 148 230 149 
<< m1 >>
rect 230 148 231 149 
<< m1 >>
rect 231 148 232 149 
<< m1 >>
rect 232 148 233 149 
<< m1 >>
rect 233 148 234 149 
<< m1 >>
rect 234 148 235 149 
<< m1 >>
rect 235 148 236 149 
<< m1 >>
rect 236 148 237 149 
<< m1 >>
rect 237 148 238 149 
<< m1 >>
rect 238 148 239 149 
<< m1 >>
rect 239 148 240 149 
<< m1 >>
rect 240 148 241 149 
<< m1 >>
rect 241 148 242 149 
<< m1 >>
rect 242 148 243 149 
<< m1 >>
rect 243 148 244 149 
<< m1 >>
rect 244 148 245 149 
<< m1 >>
rect 245 148 246 149 
<< m1 >>
rect 246 148 247 149 
<< m1 >>
rect 247 148 248 149 
<< m1 >>
rect 248 148 249 149 
<< m1 >>
rect 249 148 250 149 
<< m1 >>
rect 250 148 251 149 
<< m1 >>
rect 253 148 254 149 
<< m2 >>
rect 254 148 255 149 
<< m1 >>
rect 307 148 308 149 
<< m1 >>
rect 311 148 312 149 
<< m1 >>
rect 322 148 323 149 
<< m1 >>
rect 343 148 344 149 
<< m1 >>
rect 406 148 407 149 
<< m1 >>
rect 64 149 65 150 
<< m1 >>
rect 93 149 94 150 
<< m1 >>
rect 95 149 96 150 
<< m1 >>
rect 118 149 119 150 
<< m1 >>
rect 157 149 158 150 
<< m1 >>
rect 170 149 171 150 
<< m1 >>
rect 178 149 179 150 
<< m1 >>
rect 208 149 209 150 
<< m1 >>
rect 226 149 227 150 
<< m1 >>
rect 250 149 251 150 
<< m1 >>
rect 253 149 254 150 
<< m2 >>
rect 254 149 255 150 
<< m1 >>
rect 307 149 308 150 
<< m1 >>
rect 311 149 312 150 
<< m1 >>
rect 322 149 323 150 
<< m1 >>
rect 343 149 344 150 
<< m1 >>
rect 406 149 407 150 
<< m1 >>
rect 64 150 65 151 
<< m1 >>
rect 93 150 94 151 
<< m1 >>
rect 95 150 96 151 
<< m1 >>
rect 118 150 119 151 
<< m1 >>
rect 157 150 158 151 
<< m1 >>
rect 170 150 171 151 
<< m1 >>
rect 178 150 179 151 
<< m1 >>
rect 208 150 209 151 
<< m1 >>
rect 226 150 227 151 
<< m2 >>
rect 226 150 227 151 
<< m2 >>
rect 227 150 228 151 
<< m1 >>
rect 228 150 229 151 
<< m2 >>
rect 228 150 229 151 
<< m2c >>
rect 228 150 229 151 
<< m1 >>
rect 228 150 229 151 
<< m2 >>
rect 228 150 229 151 
<< m1 >>
rect 229 150 230 151 
<< m1 >>
rect 230 150 231 151 
<< m1 >>
rect 231 150 232 151 
<< m1 >>
rect 232 150 233 151 
<< m1 >>
rect 233 150 234 151 
<< m1 >>
rect 234 150 235 151 
<< m1 >>
rect 235 150 236 151 
<< m1 >>
rect 236 150 237 151 
<< m1 >>
rect 237 150 238 151 
<< m1 >>
rect 238 150 239 151 
<< m1 >>
rect 239 150 240 151 
<< m1 >>
rect 240 150 241 151 
<< m1 >>
rect 241 150 242 151 
<< m1 >>
rect 242 150 243 151 
<< m1 >>
rect 243 150 244 151 
<< m1 >>
rect 244 150 245 151 
<< m1 >>
rect 245 150 246 151 
<< m1 >>
rect 246 150 247 151 
<< m1 >>
rect 247 150 248 151 
<< m1 >>
rect 248 150 249 151 
<< m2 >>
rect 248 150 249 151 
<< m2c >>
rect 248 150 249 151 
<< m1 >>
rect 248 150 249 151 
<< m2 >>
rect 248 150 249 151 
<< m2 >>
rect 249 150 250 151 
<< m1 >>
rect 250 150 251 151 
<< m2 >>
rect 250 150 251 151 
<< m2 >>
rect 251 150 252 151 
<< m2 >>
rect 252 150 253 151 
<< m1 >>
rect 253 150 254 151 
<< m2 >>
rect 253 150 254 151 
<< m2 >>
rect 254 150 255 151 
<< m1 >>
rect 307 150 308 151 
<< m1 >>
rect 311 150 312 151 
<< m1 >>
rect 322 150 323 151 
<< m1 >>
rect 343 150 344 151 
<< m1 >>
rect 406 150 407 151 
<< m1 >>
rect 64 151 65 152 
<< m1 >>
rect 66 151 67 152 
<< m1 >>
rect 67 151 68 152 
<< m1 >>
rect 68 151 69 152 
<< m1 >>
rect 69 151 70 152 
<< m1 >>
rect 70 151 71 152 
<< m1 >>
rect 71 151 72 152 
<< m1 >>
rect 72 151 73 152 
<< m1 >>
rect 73 151 74 152 
<< m1 >>
rect 74 151 75 152 
<< m1 >>
rect 75 151 76 152 
<< m1 >>
rect 76 151 77 152 
<< m1 >>
rect 77 151 78 152 
<< m1 >>
rect 78 151 79 152 
<< m1 >>
rect 79 151 80 152 
<< m1 >>
rect 80 151 81 152 
<< m1 >>
rect 81 151 82 152 
<< m1 >>
rect 82 151 83 152 
<< m1 >>
rect 83 151 84 152 
<< m1 >>
rect 84 151 85 152 
<< m1 >>
rect 85 151 86 152 
<< m1 >>
rect 86 151 87 152 
<< m1 >>
rect 87 151 88 152 
<< m1 >>
rect 88 151 89 152 
<< m1 >>
rect 89 151 90 152 
<< m1 >>
rect 90 151 91 152 
<< m1 >>
rect 91 151 92 152 
<< m2 >>
rect 91 151 92 152 
<< m2c >>
rect 91 151 92 152 
<< m1 >>
rect 91 151 92 152 
<< m2 >>
rect 91 151 92 152 
<< m2 >>
rect 92 151 93 152 
<< m1 >>
rect 93 151 94 152 
<< m2 >>
rect 93 151 94 152 
<< m2 >>
rect 94 151 95 152 
<< m1 >>
rect 95 151 96 152 
<< m2 >>
rect 95 151 96 152 
<< m2c >>
rect 95 151 96 152 
<< m1 >>
rect 95 151 96 152 
<< m2 >>
rect 95 151 96 152 
<< m1 >>
rect 118 151 119 152 
<< m1 >>
rect 157 151 158 152 
<< m1 >>
rect 170 151 171 152 
<< m1 >>
rect 172 151 173 152 
<< m1 >>
rect 173 151 174 152 
<< m1 >>
rect 174 151 175 152 
<< m1 >>
rect 175 151 176 152 
<< m1 >>
rect 176 151 177 152 
<< m2 >>
rect 176 151 177 152 
<< m2c >>
rect 176 151 177 152 
<< m1 >>
rect 176 151 177 152 
<< m2 >>
rect 176 151 177 152 
<< m2 >>
rect 177 151 178 152 
<< m1 >>
rect 178 151 179 152 
<< m2 >>
rect 178 151 179 152 
<< m2 >>
rect 179 151 180 152 
<< m1 >>
rect 180 151 181 152 
<< m2 >>
rect 180 151 181 152 
<< m2c >>
rect 180 151 181 152 
<< m1 >>
rect 180 151 181 152 
<< m2 >>
rect 180 151 181 152 
<< m1 >>
rect 181 151 182 152 
<< m1 >>
rect 182 151 183 152 
<< m1 >>
rect 183 151 184 152 
<< m1 >>
rect 184 151 185 152 
<< m1 >>
rect 185 151 186 152 
<< m1 >>
rect 186 151 187 152 
<< m1 >>
rect 187 151 188 152 
<< m1 >>
rect 188 151 189 152 
<< m1 >>
rect 189 151 190 152 
<< m1 >>
rect 190 151 191 152 
<< m1 >>
rect 191 151 192 152 
<< m1 >>
rect 192 151 193 152 
<< m1 >>
rect 193 151 194 152 
<< m1 >>
rect 194 151 195 152 
<< m1 >>
rect 195 151 196 152 
<< m1 >>
rect 196 151 197 152 
<< m1 >>
rect 208 151 209 152 
<< m1 >>
rect 226 151 227 152 
<< m2 >>
rect 226 151 227 152 
<< m1 >>
rect 250 151 251 152 
<< m1 >>
rect 253 151 254 152 
<< m1 >>
rect 307 151 308 152 
<< m1 >>
rect 311 151 312 152 
<< m1 >>
rect 322 151 323 152 
<< m1 >>
rect 343 151 344 152 
<< m1 >>
rect 406 151 407 152 
<< m1 >>
rect 64 152 65 153 
<< m1 >>
rect 66 152 67 153 
<< m1 >>
rect 93 152 94 153 
<< m1 >>
rect 118 152 119 153 
<< m1 >>
rect 157 152 158 153 
<< m1 >>
rect 170 152 171 153 
<< m1 >>
rect 172 152 173 153 
<< m1 >>
rect 178 152 179 153 
<< m1 >>
rect 196 152 197 153 
<< m1 >>
rect 208 152 209 153 
<< m1 >>
rect 226 152 227 153 
<< m2 >>
rect 226 152 227 153 
<< m1 >>
rect 250 152 251 153 
<< m1 >>
rect 253 152 254 153 
<< m1 >>
rect 307 152 308 153 
<< m1 >>
rect 311 152 312 153 
<< m1 >>
rect 322 152 323 153 
<< m1 >>
rect 343 152 344 153 
<< m1 >>
rect 406 152 407 153 
<< m1 >>
rect 64 153 65 154 
<< m1 >>
rect 66 153 67 154 
<< m1 >>
rect 93 153 94 154 
<< m1 >>
rect 118 153 119 154 
<< m1 >>
rect 157 153 158 154 
<< m1 >>
rect 170 153 171 154 
<< m1 >>
rect 172 153 173 154 
<< m2 >>
rect 177 153 178 154 
<< m1 >>
rect 178 153 179 154 
<< m2 >>
rect 178 153 179 154 
<< m2 >>
rect 179 153 180 154 
<< m1 >>
rect 180 153 181 154 
<< m2 >>
rect 180 153 181 154 
<< m2c >>
rect 180 153 181 154 
<< m1 >>
rect 180 153 181 154 
<< m2 >>
rect 180 153 181 154 
<< m1 >>
rect 181 153 182 154 
<< m1 >>
rect 196 153 197 154 
<< m1 >>
rect 208 153 209 154 
<< m1 >>
rect 226 153 227 154 
<< m2 >>
rect 226 153 227 154 
<< m1 >>
rect 229 153 230 154 
<< m1 >>
rect 230 153 231 154 
<< m1 >>
rect 231 153 232 154 
<< m1 >>
rect 232 153 233 154 
<< m1 >>
rect 233 153 234 154 
<< m1 >>
rect 234 153 235 154 
<< m1 >>
rect 235 153 236 154 
<< m1 >>
rect 236 153 237 154 
<< m1 >>
rect 237 153 238 154 
<< m1 >>
rect 238 153 239 154 
<< m1 >>
rect 239 153 240 154 
<< m1 >>
rect 240 153 241 154 
<< m1 >>
rect 241 153 242 154 
<< m1 >>
rect 242 153 243 154 
<< m1 >>
rect 243 153 244 154 
<< m1 >>
rect 244 153 245 154 
<< m1 >>
rect 250 153 251 154 
<< m1 >>
rect 253 153 254 154 
<< m1 >>
rect 265 153 266 154 
<< m1 >>
rect 266 153 267 154 
<< m1 >>
rect 267 153 268 154 
<< m1 >>
rect 268 153 269 154 
<< m1 >>
rect 269 153 270 154 
<< m1 >>
rect 270 153 271 154 
<< m1 >>
rect 271 153 272 154 
<< m1 >>
rect 307 153 308 154 
<< m1 >>
rect 311 153 312 154 
<< m1 >>
rect 319 153 320 154 
<< m1 >>
rect 320 153 321 154 
<< m1 >>
rect 321 153 322 154 
<< m1 >>
rect 322 153 323 154 
<< m1 >>
rect 343 153 344 154 
<< m1 >>
rect 406 153 407 154 
<< m2 >>
rect 63 154 64 155 
<< m1 >>
rect 64 154 65 155 
<< m2 >>
rect 64 154 65 155 
<< m2 >>
rect 65 154 66 155 
<< m1 >>
rect 66 154 67 155 
<< m2 >>
rect 66 154 67 155 
<< m2c >>
rect 66 154 67 155 
<< m1 >>
rect 66 154 67 155 
<< m2 >>
rect 66 154 67 155 
<< m1 >>
rect 88 154 89 155 
<< m1 >>
rect 89 154 90 155 
<< m1 >>
rect 90 154 91 155 
<< m1 >>
rect 91 154 92 155 
<< m1 >>
rect 93 154 94 155 
<< m1 >>
rect 118 154 119 155 
<< m1 >>
rect 157 154 158 155 
<< m1 >>
rect 170 154 171 155 
<< m1 >>
rect 172 154 173 155 
<< m1 >>
rect 175 154 176 155 
<< m1 >>
rect 176 154 177 155 
<< m2 >>
rect 176 154 177 155 
<< m2c >>
rect 176 154 177 155 
<< m1 >>
rect 176 154 177 155 
<< m2 >>
rect 176 154 177 155 
<< m2 >>
rect 177 154 178 155 
<< m1 >>
rect 178 154 179 155 
<< m1 >>
rect 181 154 182 155 
<< m1 >>
rect 196 154 197 155 
<< m1 >>
rect 208 154 209 155 
<< m1 >>
rect 226 154 227 155 
<< m2 >>
rect 226 154 227 155 
<< m1 >>
rect 229 154 230 155 
<< m2 >>
rect 235 154 236 155 
<< m2 >>
rect 236 154 237 155 
<< m2 >>
rect 237 154 238 155 
<< m2 >>
rect 238 154 239 155 
<< m2 >>
rect 239 154 240 155 
<< m2 >>
rect 240 154 241 155 
<< m2 >>
rect 241 154 242 155 
<< m2 >>
rect 242 154 243 155 
<< m2 >>
rect 243 154 244 155 
<< m1 >>
rect 244 154 245 155 
<< m2 >>
rect 244 154 245 155 
<< m2 >>
rect 245 154 246 155 
<< m1 >>
rect 246 154 247 155 
<< m2 >>
rect 246 154 247 155 
<< m2c >>
rect 246 154 247 155 
<< m1 >>
rect 246 154 247 155 
<< m2 >>
rect 246 154 247 155 
<< m1 >>
rect 247 154 248 155 
<< m1 >>
rect 250 154 251 155 
<< m1 >>
rect 253 154 254 155 
<< m1 >>
rect 265 154 266 155 
<< m1 >>
rect 271 154 272 155 
<< m1 >>
rect 298 154 299 155 
<< m1 >>
rect 299 154 300 155 
<< m1 >>
rect 300 154 301 155 
<< m1 >>
rect 301 154 302 155 
<< m1 >>
rect 307 154 308 155 
<< m1 >>
rect 311 154 312 155 
<< m1 >>
rect 319 154 320 155 
<< m1 >>
rect 340 154 341 155 
<< m1 >>
rect 341 154 342 155 
<< m2 >>
rect 341 154 342 155 
<< m2c >>
rect 341 154 342 155 
<< m1 >>
rect 341 154 342 155 
<< m2 >>
rect 341 154 342 155 
<< m2 >>
rect 342 154 343 155 
<< m1 >>
rect 343 154 344 155 
<< m2 >>
rect 343 154 344 155 
<< m2 >>
rect 344 154 345 155 
<< m1 >>
rect 345 154 346 155 
<< m2 >>
rect 345 154 346 155 
<< m2c >>
rect 345 154 346 155 
<< m1 >>
rect 345 154 346 155 
<< m2 >>
rect 345 154 346 155 
<< m1 >>
rect 346 154 347 155 
<< m1 >>
rect 347 154 348 155 
<< m1 >>
rect 406 154 407 155 
<< m2 >>
rect 63 155 64 156 
<< m1 >>
rect 64 155 65 156 
<< m1 >>
rect 88 155 89 156 
<< m1 >>
rect 91 155 92 156 
<< m1 >>
rect 93 155 94 156 
<< m1 >>
rect 118 155 119 156 
<< m1 >>
rect 157 155 158 156 
<< m1 >>
rect 170 155 171 156 
<< m1 >>
rect 172 155 173 156 
<< m1 >>
rect 175 155 176 156 
<< m1 >>
rect 178 155 179 156 
<< m1 >>
rect 181 155 182 156 
<< m1 >>
rect 196 155 197 156 
<< m1 >>
rect 208 155 209 156 
<< m1 >>
rect 226 155 227 156 
<< m2 >>
rect 226 155 227 156 
<< m1 >>
rect 229 155 230 156 
<< m1 >>
rect 235 155 236 156 
<< m2 >>
rect 235 155 236 156 
<< m2c >>
rect 235 155 236 156 
<< m1 >>
rect 235 155 236 156 
<< m2 >>
rect 235 155 236 156 
<< m1 >>
rect 244 155 245 156 
<< m1 >>
rect 247 155 248 156 
<< m1 >>
rect 250 155 251 156 
<< m1 >>
rect 253 155 254 156 
<< m1 >>
rect 265 155 266 156 
<< m1 >>
rect 271 155 272 156 
<< m1 >>
rect 298 155 299 156 
<< m1 >>
rect 301 155 302 156 
<< m1 >>
rect 307 155 308 156 
<< m1 >>
rect 311 155 312 156 
<< m1 >>
rect 319 155 320 156 
<< m1 >>
rect 340 155 341 156 
<< m1 >>
rect 343 155 344 156 
<< m1 >>
rect 347 155 348 156 
<< m1 >>
rect 406 155 407 156 
<< pdiffusion >>
rect 12 156 13 157 
<< pdiffusion >>
rect 13 156 14 157 
<< pdiffusion >>
rect 14 156 15 157 
<< pdiffusion >>
rect 15 156 16 157 
<< pdiffusion >>
rect 16 156 17 157 
<< pdiffusion >>
rect 17 156 18 157 
<< pdiffusion >>
rect 48 156 49 157 
<< pdiffusion >>
rect 49 156 50 157 
<< pdiffusion >>
rect 50 156 51 157 
<< pdiffusion >>
rect 51 156 52 157 
<< pdiffusion >>
rect 52 156 53 157 
<< pdiffusion >>
rect 53 156 54 157 
<< m2 >>
rect 63 156 64 157 
<< m1 >>
rect 64 156 65 157 
<< pdiffusion >>
rect 66 156 67 157 
<< pdiffusion >>
rect 67 156 68 157 
<< pdiffusion >>
rect 68 156 69 157 
<< pdiffusion >>
rect 69 156 70 157 
<< pdiffusion >>
rect 70 156 71 157 
<< pdiffusion >>
rect 71 156 72 157 
<< pdiffusion >>
rect 84 156 85 157 
<< pdiffusion >>
rect 85 156 86 157 
<< pdiffusion >>
rect 86 156 87 157 
<< pdiffusion >>
rect 87 156 88 157 
<< m1 >>
rect 88 156 89 157 
<< pdiffusion >>
rect 88 156 89 157 
<< pdiffusion >>
rect 89 156 90 157 
<< m1 >>
rect 91 156 92 157 
<< m1 >>
rect 93 156 94 157 
<< pdiffusion >>
rect 102 156 103 157 
<< pdiffusion >>
rect 103 156 104 157 
<< pdiffusion >>
rect 104 156 105 157 
<< pdiffusion >>
rect 105 156 106 157 
<< pdiffusion >>
rect 106 156 107 157 
<< pdiffusion >>
rect 107 156 108 157 
<< m1 >>
rect 118 156 119 157 
<< pdiffusion >>
rect 120 156 121 157 
<< pdiffusion >>
rect 121 156 122 157 
<< pdiffusion >>
rect 122 156 123 157 
<< pdiffusion >>
rect 123 156 124 157 
<< pdiffusion >>
rect 124 156 125 157 
<< pdiffusion >>
rect 125 156 126 157 
<< pdiffusion >>
rect 138 156 139 157 
<< pdiffusion >>
rect 139 156 140 157 
<< pdiffusion >>
rect 140 156 141 157 
<< pdiffusion >>
rect 141 156 142 157 
<< pdiffusion >>
rect 142 156 143 157 
<< pdiffusion >>
rect 143 156 144 157 
<< pdiffusion >>
rect 156 156 157 157 
<< m1 >>
rect 157 156 158 157 
<< pdiffusion >>
rect 157 156 158 157 
<< pdiffusion >>
rect 158 156 159 157 
<< pdiffusion >>
rect 159 156 160 157 
<< pdiffusion >>
rect 160 156 161 157 
<< pdiffusion >>
rect 161 156 162 157 
<< m1 >>
rect 170 156 171 157 
<< m1 >>
rect 172 156 173 157 
<< pdiffusion >>
rect 174 156 175 157 
<< m1 >>
rect 175 156 176 157 
<< pdiffusion >>
rect 175 156 176 157 
<< pdiffusion >>
rect 176 156 177 157 
<< pdiffusion >>
rect 177 156 178 157 
<< m1 >>
rect 178 156 179 157 
<< pdiffusion >>
rect 178 156 179 157 
<< pdiffusion >>
rect 179 156 180 157 
<< m1 >>
rect 181 156 182 157 
<< pdiffusion >>
rect 192 156 193 157 
<< pdiffusion >>
rect 193 156 194 157 
<< pdiffusion >>
rect 194 156 195 157 
<< pdiffusion >>
rect 195 156 196 157 
<< m1 >>
rect 196 156 197 157 
<< pdiffusion >>
rect 196 156 197 157 
<< pdiffusion >>
rect 197 156 198 157 
<< m1 >>
rect 208 156 209 157 
<< pdiffusion >>
rect 210 156 211 157 
<< pdiffusion >>
rect 211 156 212 157 
<< pdiffusion >>
rect 212 156 213 157 
<< pdiffusion >>
rect 213 156 214 157 
<< pdiffusion >>
rect 214 156 215 157 
<< pdiffusion >>
rect 215 156 216 157 
<< m1 >>
rect 226 156 227 157 
<< m2 >>
rect 226 156 227 157 
<< pdiffusion >>
rect 228 156 229 157 
<< m1 >>
rect 229 156 230 157 
<< pdiffusion >>
rect 229 156 230 157 
<< pdiffusion >>
rect 230 156 231 157 
<< pdiffusion >>
rect 231 156 232 157 
<< pdiffusion >>
rect 232 156 233 157 
<< pdiffusion >>
rect 233 156 234 157 
<< m1 >>
rect 235 156 236 157 
<< m1 >>
rect 244 156 245 157 
<< pdiffusion >>
rect 246 156 247 157 
<< m1 >>
rect 247 156 248 157 
<< pdiffusion >>
rect 247 156 248 157 
<< pdiffusion >>
rect 248 156 249 157 
<< pdiffusion >>
rect 249 156 250 157 
<< m1 >>
rect 250 156 251 157 
<< pdiffusion >>
rect 250 156 251 157 
<< pdiffusion >>
rect 251 156 252 157 
<< m1 >>
rect 253 156 254 157 
<< pdiffusion >>
rect 264 156 265 157 
<< m1 >>
rect 265 156 266 157 
<< pdiffusion >>
rect 265 156 266 157 
<< pdiffusion >>
rect 266 156 267 157 
<< pdiffusion >>
rect 267 156 268 157 
<< pdiffusion >>
rect 268 156 269 157 
<< pdiffusion >>
rect 269 156 270 157 
<< m1 >>
rect 271 156 272 157 
<< pdiffusion >>
rect 282 156 283 157 
<< pdiffusion >>
rect 283 156 284 157 
<< pdiffusion >>
rect 284 156 285 157 
<< pdiffusion >>
rect 285 156 286 157 
<< pdiffusion >>
rect 286 156 287 157 
<< pdiffusion >>
rect 287 156 288 157 
<< m1 >>
rect 298 156 299 157 
<< pdiffusion >>
rect 300 156 301 157 
<< m1 >>
rect 301 156 302 157 
<< pdiffusion >>
rect 301 156 302 157 
<< pdiffusion >>
rect 302 156 303 157 
<< pdiffusion >>
rect 303 156 304 157 
<< pdiffusion >>
rect 304 156 305 157 
<< pdiffusion >>
rect 305 156 306 157 
<< m1 >>
rect 307 156 308 157 
<< m1 >>
rect 311 156 312 157 
<< pdiffusion >>
rect 318 156 319 157 
<< m1 >>
rect 319 156 320 157 
<< pdiffusion >>
rect 319 156 320 157 
<< pdiffusion >>
rect 320 156 321 157 
<< pdiffusion >>
rect 321 156 322 157 
<< pdiffusion >>
rect 322 156 323 157 
<< pdiffusion >>
rect 323 156 324 157 
<< pdiffusion >>
rect 336 156 337 157 
<< pdiffusion >>
rect 337 156 338 157 
<< pdiffusion >>
rect 338 156 339 157 
<< pdiffusion >>
rect 339 156 340 157 
<< m1 >>
rect 340 156 341 157 
<< pdiffusion >>
rect 340 156 341 157 
<< pdiffusion >>
rect 341 156 342 157 
<< m1 >>
rect 343 156 344 157 
<< m1 >>
rect 347 156 348 157 
<< pdiffusion >>
rect 354 156 355 157 
<< pdiffusion >>
rect 355 156 356 157 
<< pdiffusion >>
rect 356 156 357 157 
<< pdiffusion >>
rect 357 156 358 157 
<< pdiffusion >>
rect 358 156 359 157 
<< pdiffusion >>
rect 359 156 360 157 
<< pdiffusion >>
rect 372 156 373 157 
<< pdiffusion >>
rect 373 156 374 157 
<< pdiffusion >>
rect 374 156 375 157 
<< pdiffusion >>
rect 375 156 376 157 
<< pdiffusion >>
rect 376 156 377 157 
<< pdiffusion >>
rect 377 156 378 157 
<< pdiffusion >>
rect 390 156 391 157 
<< pdiffusion >>
rect 391 156 392 157 
<< pdiffusion >>
rect 392 156 393 157 
<< pdiffusion >>
rect 393 156 394 157 
<< pdiffusion >>
rect 394 156 395 157 
<< pdiffusion >>
rect 395 156 396 157 
<< m1 >>
rect 406 156 407 157 
<< pdiffusion >>
rect 408 156 409 157 
<< pdiffusion >>
rect 409 156 410 157 
<< pdiffusion >>
rect 410 156 411 157 
<< pdiffusion >>
rect 411 156 412 157 
<< pdiffusion >>
rect 412 156 413 157 
<< pdiffusion >>
rect 413 156 414 157 
<< pdiffusion >>
rect 426 156 427 157 
<< pdiffusion >>
rect 427 156 428 157 
<< pdiffusion >>
rect 428 156 429 157 
<< pdiffusion >>
rect 429 156 430 157 
<< pdiffusion >>
rect 430 156 431 157 
<< pdiffusion >>
rect 431 156 432 157 
<< pdiffusion >>
rect 444 156 445 157 
<< pdiffusion >>
rect 445 156 446 157 
<< pdiffusion >>
rect 446 156 447 157 
<< pdiffusion >>
rect 447 156 448 157 
<< pdiffusion >>
rect 448 156 449 157 
<< pdiffusion >>
rect 449 156 450 157 
<< pdiffusion >>
rect 12 157 13 158 
<< pdiffusion >>
rect 13 157 14 158 
<< pdiffusion >>
rect 14 157 15 158 
<< pdiffusion >>
rect 15 157 16 158 
<< pdiffusion >>
rect 16 157 17 158 
<< pdiffusion >>
rect 17 157 18 158 
<< pdiffusion >>
rect 48 157 49 158 
<< pdiffusion >>
rect 49 157 50 158 
<< pdiffusion >>
rect 50 157 51 158 
<< pdiffusion >>
rect 51 157 52 158 
<< pdiffusion >>
rect 52 157 53 158 
<< pdiffusion >>
rect 53 157 54 158 
<< m2 >>
rect 63 157 64 158 
<< m1 >>
rect 64 157 65 158 
<< pdiffusion >>
rect 66 157 67 158 
<< pdiffusion >>
rect 67 157 68 158 
<< pdiffusion >>
rect 68 157 69 158 
<< pdiffusion >>
rect 69 157 70 158 
<< pdiffusion >>
rect 70 157 71 158 
<< pdiffusion >>
rect 71 157 72 158 
<< pdiffusion >>
rect 84 157 85 158 
<< pdiffusion >>
rect 85 157 86 158 
<< pdiffusion >>
rect 86 157 87 158 
<< pdiffusion >>
rect 87 157 88 158 
<< pdiffusion >>
rect 88 157 89 158 
<< pdiffusion >>
rect 89 157 90 158 
<< m1 >>
rect 91 157 92 158 
<< m1 >>
rect 93 157 94 158 
<< pdiffusion >>
rect 102 157 103 158 
<< pdiffusion >>
rect 103 157 104 158 
<< pdiffusion >>
rect 104 157 105 158 
<< pdiffusion >>
rect 105 157 106 158 
<< pdiffusion >>
rect 106 157 107 158 
<< pdiffusion >>
rect 107 157 108 158 
<< m1 >>
rect 118 157 119 158 
<< pdiffusion >>
rect 120 157 121 158 
<< pdiffusion >>
rect 121 157 122 158 
<< pdiffusion >>
rect 122 157 123 158 
<< pdiffusion >>
rect 123 157 124 158 
<< pdiffusion >>
rect 124 157 125 158 
<< pdiffusion >>
rect 125 157 126 158 
<< pdiffusion >>
rect 138 157 139 158 
<< pdiffusion >>
rect 139 157 140 158 
<< pdiffusion >>
rect 140 157 141 158 
<< pdiffusion >>
rect 141 157 142 158 
<< pdiffusion >>
rect 142 157 143 158 
<< pdiffusion >>
rect 143 157 144 158 
<< pdiffusion >>
rect 156 157 157 158 
<< pdiffusion >>
rect 157 157 158 158 
<< pdiffusion >>
rect 158 157 159 158 
<< pdiffusion >>
rect 159 157 160 158 
<< pdiffusion >>
rect 160 157 161 158 
<< pdiffusion >>
rect 161 157 162 158 
<< m1 >>
rect 170 157 171 158 
<< m1 >>
rect 172 157 173 158 
<< pdiffusion >>
rect 174 157 175 158 
<< pdiffusion >>
rect 175 157 176 158 
<< pdiffusion >>
rect 176 157 177 158 
<< pdiffusion >>
rect 177 157 178 158 
<< pdiffusion >>
rect 178 157 179 158 
<< pdiffusion >>
rect 179 157 180 158 
<< m1 >>
rect 181 157 182 158 
<< pdiffusion >>
rect 192 157 193 158 
<< pdiffusion >>
rect 193 157 194 158 
<< pdiffusion >>
rect 194 157 195 158 
<< pdiffusion >>
rect 195 157 196 158 
<< pdiffusion >>
rect 196 157 197 158 
<< pdiffusion >>
rect 197 157 198 158 
<< m1 >>
rect 208 157 209 158 
<< pdiffusion >>
rect 210 157 211 158 
<< pdiffusion >>
rect 211 157 212 158 
<< pdiffusion >>
rect 212 157 213 158 
<< pdiffusion >>
rect 213 157 214 158 
<< pdiffusion >>
rect 214 157 215 158 
<< pdiffusion >>
rect 215 157 216 158 
<< m1 >>
rect 226 157 227 158 
<< m2 >>
rect 226 157 227 158 
<< pdiffusion >>
rect 228 157 229 158 
<< pdiffusion >>
rect 229 157 230 158 
<< pdiffusion >>
rect 230 157 231 158 
<< pdiffusion >>
rect 231 157 232 158 
<< pdiffusion >>
rect 232 157 233 158 
<< pdiffusion >>
rect 233 157 234 158 
<< m1 >>
rect 235 157 236 158 
<< m1 >>
rect 244 157 245 158 
<< pdiffusion >>
rect 246 157 247 158 
<< pdiffusion >>
rect 247 157 248 158 
<< pdiffusion >>
rect 248 157 249 158 
<< pdiffusion >>
rect 249 157 250 158 
<< pdiffusion >>
rect 250 157 251 158 
<< pdiffusion >>
rect 251 157 252 158 
<< m1 >>
rect 253 157 254 158 
<< pdiffusion >>
rect 264 157 265 158 
<< pdiffusion >>
rect 265 157 266 158 
<< pdiffusion >>
rect 266 157 267 158 
<< pdiffusion >>
rect 267 157 268 158 
<< pdiffusion >>
rect 268 157 269 158 
<< pdiffusion >>
rect 269 157 270 158 
<< m1 >>
rect 271 157 272 158 
<< pdiffusion >>
rect 282 157 283 158 
<< pdiffusion >>
rect 283 157 284 158 
<< pdiffusion >>
rect 284 157 285 158 
<< pdiffusion >>
rect 285 157 286 158 
<< pdiffusion >>
rect 286 157 287 158 
<< pdiffusion >>
rect 287 157 288 158 
<< m1 >>
rect 298 157 299 158 
<< pdiffusion >>
rect 300 157 301 158 
<< pdiffusion >>
rect 301 157 302 158 
<< pdiffusion >>
rect 302 157 303 158 
<< pdiffusion >>
rect 303 157 304 158 
<< pdiffusion >>
rect 304 157 305 158 
<< pdiffusion >>
rect 305 157 306 158 
<< m1 >>
rect 307 157 308 158 
<< m1 >>
rect 311 157 312 158 
<< pdiffusion >>
rect 318 157 319 158 
<< pdiffusion >>
rect 319 157 320 158 
<< pdiffusion >>
rect 320 157 321 158 
<< pdiffusion >>
rect 321 157 322 158 
<< pdiffusion >>
rect 322 157 323 158 
<< pdiffusion >>
rect 323 157 324 158 
<< pdiffusion >>
rect 336 157 337 158 
<< pdiffusion >>
rect 337 157 338 158 
<< pdiffusion >>
rect 338 157 339 158 
<< pdiffusion >>
rect 339 157 340 158 
<< pdiffusion >>
rect 340 157 341 158 
<< pdiffusion >>
rect 341 157 342 158 
<< m1 >>
rect 343 157 344 158 
<< m1 >>
rect 347 157 348 158 
<< pdiffusion >>
rect 354 157 355 158 
<< pdiffusion >>
rect 355 157 356 158 
<< pdiffusion >>
rect 356 157 357 158 
<< pdiffusion >>
rect 357 157 358 158 
<< pdiffusion >>
rect 358 157 359 158 
<< pdiffusion >>
rect 359 157 360 158 
<< pdiffusion >>
rect 372 157 373 158 
<< pdiffusion >>
rect 373 157 374 158 
<< pdiffusion >>
rect 374 157 375 158 
<< pdiffusion >>
rect 375 157 376 158 
<< pdiffusion >>
rect 376 157 377 158 
<< pdiffusion >>
rect 377 157 378 158 
<< pdiffusion >>
rect 390 157 391 158 
<< pdiffusion >>
rect 391 157 392 158 
<< pdiffusion >>
rect 392 157 393 158 
<< pdiffusion >>
rect 393 157 394 158 
<< pdiffusion >>
rect 394 157 395 158 
<< pdiffusion >>
rect 395 157 396 158 
<< m1 >>
rect 406 157 407 158 
<< pdiffusion >>
rect 408 157 409 158 
<< pdiffusion >>
rect 409 157 410 158 
<< pdiffusion >>
rect 410 157 411 158 
<< pdiffusion >>
rect 411 157 412 158 
<< pdiffusion >>
rect 412 157 413 158 
<< pdiffusion >>
rect 413 157 414 158 
<< pdiffusion >>
rect 426 157 427 158 
<< pdiffusion >>
rect 427 157 428 158 
<< pdiffusion >>
rect 428 157 429 158 
<< pdiffusion >>
rect 429 157 430 158 
<< pdiffusion >>
rect 430 157 431 158 
<< pdiffusion >>
rect 431 157 432 158 
<< pdiffusion >>
rect 444 157 445 158 
<< pdiffusion >>
rect 445 157 446 158 
<< pdiffusion >>
rect 446 157 447 158 
<< pdiffusion >>
rect 447 157 448 158 
<< pdiffusion >>
rect 448 157 449 158 
<< pdiffusion >>
rect 449 157 450 158 
<< pdiffusion >>
rect 12 158 13 159 
<< pdiffusion >>
rect 13 158 14 159 
<< pdiffusion >>
rect 14 158 15 159 
<< pdiffusion >>
rect 15 158 16 159 
<< pdiffusion >>
rect 16 158 17 159 
<< pdiffusion >>
rect 17 158 18 159 
<< pdiffusion >>
rect 48 158 49 159 
<< pdiffusion >>
rect 49 158 50 159 
<< pdiffusion >>
rect 50 158 51 159 
<< pdiffusion >>
rect 51 158 52 159 
<< pdiffusion >>
rect 52 158 53 159 
<< pdiffusion >>
rect 53 158 54 159 
<< m2 >>
rect 63 158 64 159 
<< m1 >>
rect 64 158 65 159 
<< pdiffusion >>
rect 66 158 67 159 
<< pdiffusion >>
rect 67 158 68 159 
<< pdiffusion >>
rect 68 158 69 159 
<< pdiffusion >>
rect 69 158 70 159 
<< pdiffusion >>
rect 70 158 71 159 
<< pdiffusion >>
rect 71 158 72 159 
<< pdiffusion >>
rect 84 158 85 159 
<< pdiffusion >>
rect 85 158 86 159 
<< pdiffusion >>
rect 86 158 87 159 
<< pdiffusion >>
rect 87 158 88 159 
<< pdiffusion >>
rect 88 158 89 159 
<< pdiffusion >>
rect 89 158 90 159 
<< m1 >>
rect 91 158 92 159 
<< m1 >>
rect 93 158 94 159 
<< pdiffusion >>
rect 102 158 103 159 
<< pdiffusion >>
rect 103 158 104 159 
<< pdiffusion >>
rect 104 158 105 159 
<< pdiffusion >>
rect 105 158 106 159 
<< pdiffusion >>
rect 106 158 107 159 
<< pdiffusion >>
rect 107 158 108 159 
<< m1 >>
rect 118 158 119 159 
<< pdiffusion >>
rect 120 158 121 159 
<< pdiffusion >>
rect 121 158 122 159 
<< pdiffusion >>
rect 122 158 123 159 
<< pdiffusion >>
rect 123 158 124 159 
<< pdiffusion >>
rect 124 158 125 159 
<< pdiffusion >>
rect 125 158 126 159 
<< pdiffusion >>
rect 138 158 139 159 
<< pdiffusion >>
rect 139 158 140 159 
<< pdiffusion >>
rect 140 158 141 159 
<< pdiffusion >>
rect 141 158 142 159 
<< pdiffusion >>
rect 142 158 143 159 
<< pdiffusion >>
rect 143 158 144 159 
<< pdiffusion >>
rect 156 158 157 159 
<< pdiffusion >>
rect 157 158 158 159 
<< pdiffusion >>
rect 158 158 159 159 
<< pdiffusion >>
rect 159 158 160 159 
<< pdiffusion >>
rect 160 158 161 159 
<< pdiffusion >>
rect 161 158 162 159 
<< m1 >>
rect 170 158 171 159 
<< m1 >>
rect 172 158 173 159 
<< pdiffusion >>
rect 174 158 175 159 
<< pdiffusion >>
rect 175 158 176 159 
<< pdiffusion >>
rect 176 158 177 159 
<< pdiffusion >>
rect 177 158 178 159 
<< pdiffusion >>
rect 178 158 179 159 
<< pdiffusion >>
rect 179 158 180 159 
<< m1 >>
rect 181 158 182 159 
<< pdiffusion >>
rect 192 158 193 159 
<< pdiffusion >>
rect 193 158 194 159 
<< pdiffusion >>
rect 194 158 195 159 
<< pdiffusion >>
rect 195 158 196 159 
<< pdiffusion >>
rect 196 158 197 159 
<< pdiffusion >>
rect 197 158 198 159 
<< m1 >>
rect 208 158 209 159 
<< pdiffusion >>
rect 210 158 211 159 
<< pdiffusion >>
rect 211 158 212 159 
<< pdiffusion >>
rect 212 158 213 159 
<< pdiffusion >>
rect 213 158 214 159 
<< pdiffusion >>
rect 214 158 215 159 
<< pdiffusion >>
rect 215 158 216 159 
<< m1 >>
rect 226 158 227 159 
<< m2 >>
rect 226 158 227 159 
<< pdiffusion >>
rect 228 158 229 159 
<< pdiffusion >>
rect 229 158 230 159 
<< pdiffusion >>
rect 230 158 231 159 
<< pdiffusion >>
rect 231 158 232 159 
<< pdiffusion >>
rect 232 158 233 159 
<< pdiffusion >>
rect 233 158 234 159 
<< m1 >>
rect 235 158 236 159 
<< m1 >>
rect 244 158 245 159 
<< pdiffusion >>
rect 246 158 247 159 
<< pdiffusion >>
rect 247 158 248 159 
<< pdiffusion >>
rect 248 158 249 159 
<< pdiffusion >>
rect 249 158 250 159 
<< pdiffusion >>
rect 250 158 251 159 
<< pdiffusion >>
rect 251 158 252 159 
<< m1 >>
rect 253 158 254 159 
<< pdiffusion >>
rect 264 158 265 159 
<< pdiffusion >>
rect 265 158 266 159 
<< pdiffusion >>
rect 266 158 267 159 
<< pdiffusion >>
rect 267 158 268 159 
<< pdiffusion >>
rect 268 158 269 159 
<< pdiffusion >>
rect 269 158 270 159 
<< m1 >>
rect 271 158 272 159 
<< pdiffusion >>
rect 282 158 283 159 
<< pdiffusion >>
rect 283 158 284 159 
<< pdiffusion >>
rect 284 158 285 159 
<< pdiffusion >>
rect 285 158 286 159 
<< pdiffusion >>
rect 286 158 287 159 
<< pdiffusion >>
rect 287 158 288 159 
<< m1 >>
rect 298 158 299 159 
<< pdiffusion >>
rect 300 158 301 159 
<< pdiffusion >>
rect 301 158 302 159 
<< pdiffusion >>
rect 302 158 303 159 
<< pdiffusion >>
rect 303 158 304 159 
<< pdiffusion >>
rect 304 158 305 159 
<< pdiffusion >>
rect 305 158 306 159 
<< m1 >>
rect 307 158 308 159 
<< m1 >>
rect 311 158 312 159 
<< pdiffusion >>
rect 318 158 319 159 
<< pdiffusion >>
rect 319 158 320 159 
<< pdiffusion >>
rect 320 158 321 159 
<< pdiffusion >>
rect 321 158 322 159 
<< pdiffusion >>
rect 322 158 323 159 
<< pdiffusion >>
rect 323 158 324 159 
<< pdiffusion >>
rect 336 158 337 159 
<< pdiffusion >>
rect 337 158 338 159 
<< pdiffusion >>
rect 338 158 339 159 
<< pdiffusion >>
rect 339 158 340 159 
<< pdiffusion >>
rect 340 158 341 159 
<< pdiffusion >>
rect 341 158 342 159 
<< m1 >>
rect 343 158 344 159 
<< m1 >>
rect 347 158 348 159 
<< pdiffusion >>
rect 354 158 355 159 
<< pdiffusion >>
rect 355 158 356 159 
<< pdiffusion >>
rect 356 158 357 159 
<< pdiffusion >>
rect 357 158 358 159 
<< pdiffusion >>
rect 358 158 359 159 
<< pdiffusion >>
rect 359 158 360 159 
<< pdiffusion >>
rect 372 158 373 159 
<< pdiffusion >>
rect 373 158 374 159 
<< pdiffusion >>
rect 374 158 375 159 
<< pdiffusion >>
rect 375 158 376 159 
<< pdiffusion >>
rect 376 158 377 159 
<< pdiffusion >>
rect 377 158 378 159 
<< pdiffusion >>
rect 390 158 391 159 
<< pdiffusion >>
rect 391 158 392 159 
<< pdiffusion >>
rect 392 158 393 159 
<< pdiffusion >>
rect 393 158 394 159 
<< pdiffusion >>
rect 394 158 395 159 
<< pdiffusion >>
rect 395 158 396 159 
<< m1 >>
rect 406 158 407 159 
<< pdiffusion >>
rect 408 158 409 159 
<< pdiffusion >>
rect 409 158 410 159 
<< pdiffusion >>
rect 410 158 411 159 
<< pdiffusion >>
rect 411 158 412 159 
<< pdiffusion >>
rect 412 158 413 159 
<< pdiffusion >>
rect 413 158 414 159 
<< pdiffusion >>
rect 426 158 427 159 
<< pdiffusion >>
rect 427 158 428 159 
<< pdiffusion >>
rect 428 158 429 159 
<< pdiffusion >>
rect 429 158 430 159 
<< pdiffusion >>
rect 430 158 431 159 
<< pdiffusion >>
rect 431 158 432 159 
<< pdiffusion >>
rect 444 158 445 159 
<< pdiffusion >>
rect 445 158 446 159 
<< pdiffusion >>
rect 446 158 447 159 
<< pdiffusion >>
rect 447 158 448 159 
<< pdiffusion >>
rect 448 158 449 159 
<< pdiffusion >>
rect 449 158 450 159 
<< pdiffusion >>
rect 12 159 13 160 
<< pdiffusion >>
rect 13 159 14 160 
<< pdiffusion >>
rect 14 159 15 160 
<< pdiffusion >>
rect 15 159 16 160 
<< pdiffusion >>
rect 16 159 17 160 
<< pdiffusion >>
rect 17 159 18 160 
<< pdiffusion >>
rect 48 159 49 160 
<< pdiffusion >>
rect 49 159 50 160 
<< pdiffusion >>
rect 50 159 51 160 
<< pdiffusion >>
rect 51 159 52 160 
<< pdiffusion >>
rect 52 159 53 160 
<< pdiffusion >>
rect 53 159 54 160 
<< m2 >>
rect 63 159 64 160 
<< m1 >>
rect 64 159 65 160 
<< pdiffusion >>
rect 66 159 67 160 
<< pdiffusion >>
rect 67 159 68 160 
<< pdiffusion >>
rect 68 159 69 160 
<< pdiffusion >>
rect 69 159 70 160 
<< pdiffusion >>
rect 70 159 71 160 
<< pdiffusion >>
rect 71 159 72 160 
<< pdiffusion >>
rect 84 159 85 160 
<< pdiffusion >>
rect 85 159 86 160 
<< pdiffusion >>
rect 86 159 87 160 
<< pdiffusion >>
rect 87 159 88 160 
<< pdiffusion >>
rect 88 159 89 160 
<< pdiffusion >>
rect 89 159 90 160 
<< m1 >>
rect 91 159 92 160 
<< m1 >>
rect 93 159 94 160 
<< pdiffusion >>
rect 102 159 103 160 
<< pdiffusion >>
rect 103 159 104 160 
<< pdiffusion >>
rect 104 159 105 160 
<< pdiffusion >>
rect 105 159 106 160 
<< pdiffusion >>
rect 106 159 107 160 
<< pdiffusion >>
rect 107 159 108 160 
<< m1 >>
rect 118 159 119 160 
<< pdiffusion >>
rect 120 159 121 160 
<< pdiffusion >>
rect 121 159 122 160 
<< pdiffusion >>
rect 122 159 123 160 
<< pdiffusion >>
rect 123 159 124 160 
<< pdiffusion >>
rect 124 159 125 160 
<< pdiffusion >>
rect 125 159 126 160 
<< pdiffusion >>
rect 138 159 139 160 
<< pdiffusion >>
rect 139 159 140 160 
<< pdiffusion >>
rect 140 159 141 160 
<< pdiffusion >>
rect 141 159 142 160 
<< pdiffusion >>
rect 142 159 143 160 
<< pdiffusion >>
rect 143 159 144 160 
<< pdiffusion >>
rect 156 159 157 160 
<< pdiffusion >>
rect 157 159 158 160 
<< pdiffusion >>
rect 158 159 159 160 
<< pdiffusion >>
rect 159 159 160 160 
<< pdiffusion >>
rect 160 159 161 160 
<< pdiffusion >>
rect 161 159 162 160 
<< m1 >>
rect 170 159 171 160 
<< m1 >>
rect 172 159 173 160 
<< pdiffusion >>
rect 174 159 175 160 
<< pdiffusion >>
rect 175 159 176 160 
<< pdiffusion >>
rect 176 159 177 160 
<< pdiffusion >>
rect 177 159 178 160 
<< pdiffusion >>
rect 178 159 179 160 
<< pdiffusion >>
rect 179 159 180 160 
<< m1 >>
rect 181 159 182 160 
<< pdiffusion >>
rect 192 159 193 160 
<< pdiffusion >>
rect 193 159 194 160 
<< pdiffusion >>
rect 194 159 195 160 
<< pdiffusion >>
rect 195 159 196 160 
<< pdiffusion >>
rect 196 159 197 160 
<< pdiffusion >>
rect 197 159 198 160 
<< m1 >>
rect 208 159 209 160 
<< pdiffusion >>
rect 210 159 211 160 
<< pdiffusion >>
rect 211 159 212 160 
<< pdiffusion >>
rect 212 159 213 160 
<< pdiffusion >>
rect 213 159 214 160 
<< pdiffusion >>
rect 214 159 215 160 
<< pdiffusion >>
rect 215 159 216 160 
<< m1 >>
rect 226 159 227 160 
<< m2 >>
rect 226 159 227 160 
<< pdiffusion >>
rect 228 159 229 160 
<< pdiffusion >>
rect 229 159 230 160 
<< pdiffusion >>
rect 230 159 231 160 
<< pdiffusion >>
rect 231 159 232 160 
<< pdiffusion >>
rect 232 159 233 160 
<< pdiffusion >>
rect 233 159 234 160 
<< m1 >>
rect 235 159 236 160 
<< m1 >>
rect 244 159 245 160 
<< pdiffusion >>
rect 246 159 247 160 
<< pdiffusion >>
rect 247 159 248 160 
<< pdiffusion >>
rect 248 159 249 160 
<< pdiffusion >>
rect 249 159 250 160 
<< pdiffusion >>
rect 250 159 251 160 
<< pdiffusion >>
rect 251 159 252 160 
<< m1 >>
rect 253 159 254 160 
<< pdiffusion >>
rect 264 159 265 160 
<< pdiffusion >>
rect 265 159 266 160 
<< pdiffusion >>
rect 266 159 267 160 
<< pdiffusion >>
rect 267 159 268 160 
<< pdiffusion >>
rect 268 159 269 160 
<< pdiffusion >>
rect 269 159 270 160 
<< m1 >>
rect 271 159 272 160 
<< pdiffusion >>
rect 282 159 283 160 
<< pdiffusion >>
rect 283 159 284 160 
<< pdiffusion >>
rect 284 159 285 160 
<< pdiffusion >>
rect 285 159 286 160 
<< pdiffusion >>
rect 286 159 287 160 
<< pdiffusion >>
rect 287 159 288 160 
<< m1 >>
rect 298 159 299 160 
<< pdiffusion >>
rect 300 159 301 160 
<< pdiffusion >>
rect 301 159 302 160 
<< pdiffusion >>
rect 302 159 303 160 
<< pdiffusion >>
rect 303 159 304 160 
<< pdiffusion >>
rect 304 159 305 160 
<< pdiffusion >>
rect 305 159 306 160 
<< m1 >>
rect 307 159 308 160 
<< m1 >>
rect 311 159 312 160 
<< pdiffusion >>
rect 318 159 319 160 
<< pdiffusion >>
rect 319 159 320 160 
<< pdiffusion >>
rect 320 159 321 160 
<< pdiffusion >>
rect 321 159 322 160 
<< pdiffusion >>
rect 322 159 323 160 
<< pdiffusion >>
rect 323 159 324 160 
<< pdiffusion >>
rect 336 159 337 160 
<< pdiffusion >>
rect 337 159 338 160 
<< pdiffusion >>
rect 338 159 339 160 
<< pdiffusion >>
rect 339 159 340 160 
<< pdiffusion >>
rect 340 159 341 160 
<< pdiffusion >>
rect 341 159 342 160 
<< m1 >>
rect 343 159 344 160 
<< m1 >>
rect 347 159 348 160 
<< pdiffusion >>
rect 354 159 355 160 
<< pdiffusion >>
rect 355 159 356 160 
<< pdiffusion >>
rect 356 159 357 160 
<< pdiffusion >>
rect 357 159 358 160 
<< pdiffusion >>
rect 358 159 359 160 
<< pdiffusion >>
rect 359 159 360 160 
<< pdiffusion >>
rect 372 159 373 160 
<< pdiffusion >>
rect 373 159 374 160 
<< pdiffusion >>
rect 374 159 375 160 
<< pdiffusion >>
rect 375 159 376 160 
<< pdiffusion >>
rect 376 159 377 160 
<< pdiffusion >>
rect 377 159 378 160 
<< pdiffusion >>
rect 390 159 391 160 
<< pdiffusion >>
rect 391 159 392 160 
<< pdiffusion >>
rect 392 159 393 160 
<< pdiffusion >>
rect 393 159 394 160 
<< pdiffusion >>
rect 394 159 395 160 
<< pdiffusion >>
rect 395 159 396 160 
<< m1 >>
rect 406 159 407 160 
<< pdiffusion >>
rect 408 159 409 160 
<< pdiffusion >>
rect 409 159 410 160 
<< pdiffusion >>
rect 410 159 411 160 
<< pdiffusion >>
rect 411 159 412 160 
<< pdiffusion >>
rect 412 159 413 160 
<< pdiffusion >>
rect 413 159 414 160 
<< pdiffusion >>
rect 426 159 427 160 
<< pdiffusion >>
rect 427 159 428 160 
<< pdiffusion >>
rect 428 159 429 160 
<< pdiffusion >>
rect 429 159 430 160 
<< pdiffusion >>
rect 430 159 431 160 
<< pdiffusion >>
rect 431 159 432 160 
<< pdiffusion >>
rect 444 159 445 160 
<< pdiffusion >>
rect 445 159 446 160 
<< pdiffusion >>
rect 446 159 447 160 
<< pdiffusion >>
rect 447 159 448 160 
<< pdiffusion >>
rect 448 159 449 160 
<< pdiffusion >>
rect 449 159 450 160 
<< pdiffusion >>
rect 12 160 13 161 
<< pdiffusion >>
rect 13 160 14 161 
<< pdiffusion >>
rect 14 160 15 161 
<< pdiffusion >>
rect 15 160 16 161 
<< pdiffusion >>
rect 16 160 17 161 
<< pdiffusion >>
rect 17 160 18 161 
<< pdiffusion >>
rect 48 160 49 161 
<< pdiffusion >>
rect 49 160 50 161 
<< pdiffusion >>
rect 50 160 51 161 
<< pdiffusion >>
rect 51 160 52 161 
<< pdiffusion >>
rect 52 160 53 161 
<< pdiffusion >>
rect 53 160 54 161 
<< m2 >>
rect 63 160 64 161 
<< m1 >>
rect 64 160 65 161 
<< pdiffusion >>
rect 66 160 67 161 
<< pdiffusion >>
rect 67 160 68 161 
<< pdiffusion >>
rect 68 160 69 161 
<< pdiffusion >>
rect 69 160 70 161 
<< pdiffusion >>
rect 70 160 71 161 
<< pdiffusion >>
rect 71 160 72 161 
<< pdiffusion >>
rect 84 160 85 161 
<< pdiffusion >>
rect 85 160 86 161 
<< pdiffusion >>
rect 86 160 87 161 
<< pdiffusion >>
rect 87 160 88 161 
<< pdiffusion >>
rect 88 160 89 161 
<< pdiffusion >>
rect 89 160 90 161 
<< m1 >>
rect 91 160 92 161 
<< m1 >>
rect 93 160 94 161 
<< pdiffusion >>
rect 102 160 103 161 
<< pdiffusion >>
rect 103 160 104 161 
<< pdiffusion >>
rect 104 160 105 161 
<< pdiffusion >>
rect 105 160 106 161 
<< pdiffusion >>
rect 106 160 107 161 
<< pdiffusion >>
rect 107 160 108 161 
<< m1 >>
rect 118 160 119 161 
<< pdiffusion >>
rect 120 160 121 161 
<< pdiffusion >>
rect 121 160 122 161 
<< pdiffusion >>
rect 122 160 123 161 
<< pdiffusion >>
rect 123 160 124 161 
<< pdiffusion >>
rect 124 160 125 161 
<< pdiffusion >>
rect 125 160 126 161 
<< pdiffusion >>
rect 138 160 139 161 
<< pdiffusion >>
rect 139 160 140 161 
<< pdiffusion >>
rect 140 160 141 161 
<< pdiffusion >>
rect 141 160 142 161 
<< pdiffusion >>
rect 142 160 143 161 
<< pdiffusion >>
rect 143 160 144 161 
<< pdiffusion >>
rect 156 160 157 161 
<< pdiffusion >>
rect 157 160 158 161 
<< pdiffusion >>
rect 158 160 159 161 
<< pdiffusion >>
rect 159 160 160 161 
<< pdiffusion >>
rect 160 160 161 161 
<< pdiffusion >>
rect 161 160 162 161 
<< m1 >>
rect 170 160 171 161 
<< m1 >>
rect 172 160 173 161 
<< pdiffusion >>
rect 174 160 175 161 
<< pdiffusion >>
rect 175 160 176 161 
<< pdiffusion >>
rect 176 160 177 161 
<< pdiffusion >>
rect 177 160 178 161 
<< pdiffusion >>
rect 178 160 179 161 
<< pdiffusion >>
rect 179 160 180 161 
<< m1 >>
rect 181 160 182 161 
<< pdiffusion >>
rect 192 160 193 161 
<< pdiffusion >>
rect 193 160 194 161 
<< pdiffusion >>
rect 194 160 195 161 
<< pdiffusion >>
rect 195 160 196 161 
<< pdiffusion >>
rect 196 160 197 161 
<< pdiffusion >>
rect 197 160 198 161 
<< m1 >>
rect 208 160 209 161 
<< pdiffusion >>
rect 210 160 211 161 
<< pdiffusion >>
rect 211 160 212 161 
<< pdiffusion >>
rect 212 160 213 161 
<< pdiffusion >>
rect 213 160 214 161 
<< pdiffusion >>
rect 214 160 215 161 
<< pdiffusion >>
rect 215 160 216 161 
<< m1 >>
rect 226 160 227 161 
<< m2 >>
rect 226 160 227 161 
<< pdiffusion >>
rect 228 160 229 161 
<< pdiffusion >>
rect 229 160 230 161 
<< pdiffusion >>
rect 230 160 231 161 
<< pdiffusion >>
rect 231 160 232 161 
<< pdiffusion >>
rect 232 160 233 161 
<< pdiffusion >>
rect 233 160 234 161 
<< m1 >>
rect 235 160 236 161 
<< m1 >>
rect 244 160 245 161 
<< pdiffusion >>
rect 246 160 247 161 
<< pdiffusion >>
rect 247 160 248 161 
<< pdiffusion >>
rect 248 160 249 161 
<< pdiffusion >>
rect 249 160 250 161 
<< pdiffusion >>
rect 250 160 251 161 
<< pdiffusion >>
rect 251 160 252 161 
<< m1 >>
rect 253 160 254 161 
<< pdiffusion >>
rect 264 160 265 161 
<< pdiffusion >>
rect 265 160 266 161 
<< pdiffusion >>
rect 266 160 267 161 
<< pdiffusion >>
rect 267 160 268 161 
<< pdiffusion >>
rect 268 160 269 161 
<< pdiffusion >>
rect 269 160 270 161 
<< m1 >>
rect 271 160 272 161 
<< pdiffusion >>
rect 282 160 283 161 
<< pdiffusion >>
rect 283 160 284 161 
<< pdiffusion >>
rect 284 160 285 161 
<< pdiffusion >>
rect 285 160 286 161 
<< pdiffusion >>
rect 286 160 287 161 
<< pdiffusion >>
rect 287 160 288 161 
<< m1 >>
rect 298 160 299 161 
<< pdiffusion >>
rect 300 160 301 161 
<< pdiffusion >>
rect 301 160 302 161 
<< pdiffusion >>
rect 302 160 303 161 
<< pdiffusion >>
rect 303 160 304 161 
<< pdiffusion >>
rect 304 160 305 161 
<< pdiffusion >>
rect 305 160 306 161 
<< m1 >>
rect 307 160 308 161 
<< m1 >>
rect 311 160 312 161 
<< pdiffusion >>
rect 318 160 319 161 
<< pdiffusion >>
rect 319 160 320 161 
<< pdiffusion >>
rect 320 160 321 161 
<< pdiffusion >>
rect 321 160 322 161 
<< pdiffusion >>
rect 322 160 323 161 
<< pdiffusion >>
rect 323 160 324 161 
<< pdiffusion >>
rect 336 160 337 161 
<< pdiffusion >>
rect 337 160 338 161 
<< pdiffusion >>
rect 338 160 339 161 
<< pdiffusion >>
rect 339 160 340 161 
<< pdiffusion >>
rect 340 160 341 161 
<< pdiffusion >>
rect 341 160 342 161 
<< m1 >>
rect 343 160 344 161 
<< m1 >>
rect 347 160 348 161 
<< pdiffusion >>
rect 354 160 355 161 
<< pdiffusion >>
rect 355 160 356 161 
<< pdiffusion >>
rect 356 160 357 161 
<< pdiffusion >>
rect 357 160 358 161 
<< pdiffusion >>
rect 358 160 359 161 
<< pdiffusion >>
rect 359 160 360 161 
<< pdiffusion >>
rect 372 160 373 161 
<< pdiffusion >>
rect 373 160 374 161 
<< pdiffusion >>
rect 374 160 375 161 
<< pdiffusion >>
rect 375 160 376 161 
<< pdiffusion >>
rect 376 160 377 161 
<< pdiffusion >>
rect 377 160 378 161 
<< pdiffusion >>
rect 390 160 391 161 
<< pdiffusion >>
rect 391 160 392 161 
<< pdiffusion >>
rect 392 160 393 161 
<< pdiffusion >>
rect 393 160 394 161 
<< pdiffusion >>
rect 394 160 395 161 
<< pdiffusion >>
rect 395 160 396 161 
<< m1 >>
rect 406 160 407 161 
<< pdiffusion >>
rect 408 160 409 161 
<< pdiffusion >>
rect 409 160 410 161 
<< pdiffusion >>
rect 410 160 411 161 
<< pdiffusion >>
rect 411 160 412 161 
<< pdiffusion >>
rect 412 160 413 161 
<< pdiffusion >>
rect 413 160 414 161 
<< pdiffusion >>
rect 426 160 427 161 
<< pdiffusion >>
rect 427 160 428 161 
<< pdiffusion >>
rect 428 160 429 161 
<< pdiffusion >>
rect 429 160 430 161 
<< pdiffusion >>
rect 430 160 431 161 
<< pdiffusion >>
rect 431 160 432 161 
<< pdiffusion >>
rect 444 160 445 161 
<< pdiffusion >>
rect 445 160 446 161 
<< pdiffusion >>
rect 446 160 447 161 
<< pdiffusion >>
rect 447 160 448 161 
<< pdiffusion >>
rect 448 160 449 161 
<< pdiffusion >>
rect 449 160 450 161 
<< pdiffusion >>
rect 12 161 13 162 
<< pdiffusion >>
rect 13 161 14 162 
<< pdiffusion >>
rect 14 161 15 162 
<< pdiffusion >>
rect 15 161 16 162 
<< pdiffusion >>
rect 16 161 17 162 
<< pdiffusion >>
rect 17 161 18 162 
<< pdiffusion >>
rect 48 161 49 162 
<< m1 >>
rect 49 161 50 162 
<< pdiffusion >>
rect 49 161 50 162 
<< pdiffusion >>
rect 50 161 51 162 
<< pdiffusion >>
rect 51 161 52 162 
<< pdiffusion >>
rect 52 161 53 162 
<< pdiffusion >>
rect 53 161 54 162 
<< m2 >>
rect 63 161 64 162 
<< m1 >>
rect 64 161 65 162 
<< pdiffusion >>
rect 66 161 67 162 
<< pdiffusion >>
rect 67 161 68 162 
<< pdiffusion >>
rect 68 161 69 162 
<< pdiffusion >>
rect 69 161 70 162 
<< pdiffusion >>
rect 70 161 71 162 
<< pdiffusion >>
rect 71 161 72 162 
<< pdiffusion >>
rect 84 161 85 162 
<< pdiffusion >>
rect 85 161 86 162 
<< pdiffusion >>
rect 86 161 87 162 
<< pdiffusion >>
rect 87 161 88 162 
<< pdiffusion >>
rect 88 161 89 162 
<< pdiffusion >>
rect 89 161 90 162 
<< m1 >>
rect 91 161 92 162 
<< m1 >>
rect 93 161 94 162 
<< pdiffusion >>
rect 102 161 103 162 
<< pdiffusion >>
rect 103 161 104 162 
<< pdiffusion >>
rect 104 161 105 162 
<< pdiffusion >>
rect 105 161 106 162 
<< m1 >>
rect 106 161 107 162 
<< pdiffusion >>
rect 106 161 107 162 
<< pdiffusion >>
rect 107 161 108 162 
<< m1 >>
rect 118 161 119 162 
<< pdiffusion >>
rect 120 161 121 162 
<< m1 >>
rect 121 161 122 162 
<< pdiffusion >>
rect 121 161 122 162 
<< pdiffusion >>
rect 122 161 123 162 
<< pdiffusion >>
rect 123 161 124 162 
<< pdiffusion >>
rect 124 161 125 162 
<< pdiffusion >>
rect 125 161 126 162 
<< pdiffusion >>
rect 138 161 139 162 
<< pdiffusion >>
rect 139 161 140 162 
<< pdiffusion >>
rect 140 161 141 162 
<< pdiffusion >>
rect 141 161 142 162 
<< pdiffusion >>
rect 142 161 143 162 
<< pdiffusion >>
rect 143 161 144 162 
<< pdiffusion >>
rect 156 161 157 162 
<< pdiffusion >>
rect 157 161 158 162 
<< pdiffusion >>
rect 158 161 159 162 
<< pdiffusion >>
rect 159 161 160 162 
<< m1 >>
rect 160 161 161 162 
<< pdiffusion >>
rect 160 161 161 162 
<< pdiffusion >>
rect 161 161 162 162 
<< m1 >>
rect 170 161 171 162 
<< m1 >>
rect 172 161 173 162 
<< pdiffusion >>
rect 174 161 175 162 
<< pdiffusion >>
rect 175 161 176 162 
<< pdiffusion >>
rect 176 161 177 162 
<< pdiffusion >>
rect 177 161 178 162 
<< pdiffusion >>
rect 178 161 179 162 
<< pdiffusion >>
rect 179 161 180 162 
<< m1 >>
rect 181 161 182 162 
<< pdiffusion >>
rect 192 161 193 162 
<< m1 >>
rect 193 161 194 162 
<< pdiffusion >>
rect 193 161 194 162 
<< pdiffusion >>
rect 194 161 195 162 
<< pdiffusion >>
rect 195 161 196 162 
<< pdiffusion >>
rect 196 161 197 162 
<< pdiffusion >>
rect 197 161 198 162 
<< m1 >>
rect 208 161 209 162 
<< pdiffusion >>
rect 210 161 211 162 
<< pdiffusion >>
rect 211 161 212 162 
<< pdiffusion >>
rect 212 161 213 162 
<< pdiffusion >>
rect 213 161 214 162 
<< pdiffusion >>
rect 214 161 215 162 
<< pdiffusion >>
rect 215 161 216 162 
<< m1 >>
rect 226 161 227 162 
<< m2 >>
rect 226 161 227 162 
<< pdiffusion >>
rect 228 161 229 162 
<< pdiffusion >>
rect 229 161 230 162 
<< pdiffusion >>
rect 230 161 231 162 
<< pdiffusion >>
rect 231 161 232 162 
<< m1 >>
rect 232 161 233 162 
<< pdiffusion >>
rect 232 161 233 162 
<< pdiffusion >>
rect 233 161 234 162 
<< m1 >>
rect 235 161 236 162 
<< m1 >>
rect 244 161 245 162 
<< pdiffusion >>
rect 246 161 247 162 
<< m1 >>
rect 247 161 248 162 
<< pdiffusion >>
rect 247 161 248 162 
<< pdiffusion >>
rect 248 161 249 162 
<< pdiffusion >>
rect 249 161 250 162 
<< pdiffusion >>
rect 250 161 251 162 
<< pdiffusion >>
rect 251 161 252 162 
<< m1 >>
rect 253 161 254 162 
<< pdiffusion >>
rect 264 161 265 162 
<< pdiffusion >>
rect 265 161 266 162 
<< pdiffusion >>
rect 266 161 267 162 
<< pdiffusion >>
rect 267 161 268 162 
<< pdiffusion >>
rect 268 161 269 162 
<< pdiffusion >>
rect 269 161 270 162 
<< m1 >>
rect 271 161 272 162 
<< pdiffusion >>
rect 282 161 283 162 
<< m1 >>
rect 283 161 284 162 
<< pdiffusion >>
rect 283 161 284 162 
<< pdiffusion >>
rect 284 161 285 162 
<< pdiffusion >>
rect 285 161 286 162 
<< pdiffusion >>
rect 286 161 287 162 
<< pdiffusion >>
rect 287 161 288 162 
<< m1 >>
rect 298 161 299 162 
<< pdiffusion >>
rect 300 161 301 162 
<< pdiffusion >>
rect 301 161 302 162 
<< pdiffusion >>
rect 302 161 303 162 
<< pdiffusion >>
rect 303 161 304 162 
<< pdiffusion >>
rect 304 161 305 162 
<< pdiffusion >>
rect 305 161 306 162 
<< m1 >>
rect 307 161 308 162 
<< m1 >>
rect 311 161 312 162 
<< pdiffusion >>
rect 318 161 319 162 
<< pdiffusion >>
rect 319 161 320 162 
<< pdiffusion >>
rect 320 161 321 162 
<< pdiffusion >>
rect 321 161 322 162 
<< pdiffusion >>
rect 322 161 323 162 
<< pdiffusion >>
rect 323 161 324 162 
<< pdiffusion >>
rect 336 161 337 162 
<< pdiffusion >>
rect 337 161 338 162 
<< pdiffusion >>
rect 338 161 339 162 
<< pdiffusion >>
rect 339 161 340 162 
<< pdiffusion >>
rect 340 161 341 162 
<< pdiffusion >>
rect 341 161 342 162 
<< m1 >>
rect 343 161 344 162 
<< m1 >>
rect 347 161 348 162 
<< pdiffusion >>
rect 354 161 355 162 
<< pdiffusion >>
rect 355 161 356 162 
<< pdiffusion >>
rect 356 161 357 162 
<< pdiffusion >>
rect 357 161 358 162 
<< pdiffusion >>
rect 358 161 359 162 
<< pdiffusion >>
rect 359 161 360 162 
<< pdiffusion >>
rect 372 161 373 162 
<< pdiffusion >>
rect 373 161 374 162 
<< pdiffusion >>
rect 374 161 375 162 
<< pdiffusion >>
rect 375 161 376 162 
<< pdiffusion >>
rect 376 161 377 162 
<< pdiffusion >>
rect 377 161 378 162 
<< pdiffusion >>
rect 390 161 391 162 
<< m1 >>
rect 391 161 392 162 
<< pdiffusion >>
rect 391 161 392 162 
<< pdiffusion >>
rect 392 161 393 162 
<< pdiffusion >>
rect 393 161 394 162 
<< pdiffusion >>
rect 394 161 395 162 
<< pdiffusion >>
rect 395 161 396 162 
<< m1 >>
rect 406 161 407 162 
<< pdiffusion >>
rect 408 161 409 162 
<< pdiffusion >>
rect 409 161 410 162 
<< pdiffusion >>
rect 410 161 411 162 
<< pdiffusion >>
rect 411 161 412 162 
<< pdiffusion >>
rect 412 161 413 162 
<< pdiffusion >>
rect 413 161 414 162 
<< pdiffusion >>
rect 426 161 427 162 
<< pdiffusion >>
rect 427 161 428 162 
<< pdiffusion >>
rect 428 161 429 162 
<< pdiffusion >>
rect 429 161 430 162 
<< pdiffusion >>
rect 430 161 431 162 
<< pdiffusion >>
rect 431 161 432 162 
<< pdiffusion >>
rect 444 161 445 162 
<< pdiffusion >>
rect 445 161 446 162 
<< pdiffusion >>
rect 446 161 447 162 
<< pdiffusion >>
rect 447 161 448 162 
<< pdiffusion >>
rect 448 161 449 162 
<< pdiffusion >>
rect 449 161 450 162 
<< m1 >>
rect 49 162 50 163 
<< m2 >>
rect 63 162 64 163 
<< m1 >>
rect 64 162 65 163 
<< m1 >>
rect 91 162 92 163 
<< m1 >>
rect 93 162 94 163 
<< m1 >>
rect 106 162 107 163 
<< m1 >>
rect 118 162 119 163 
<< m1 >>
rect 121 162 122 163 
<< m1 >>
rect 160 162 161 163 
<< m1 >>
rect 170 162 171 163 
<< m1 >>
rect 172 162 173 163 
<< m1 >>
rect 181 162 182 163 
<< m1 >>
rect 193 162 194 163 
<< m1 >>
rect 208 162 209 163 
<< m1 >>
rect 226 162 227 163 
<< m2 >>
rect 226 162 227 163 
<< m1 >>
rect 232 162 233 163 
<< m1 >>
rect 235 162 236 163 
<< m1 >>
rect 244 162 245 163 
<< m1 >>
rect 247 162 248 163 
<< m1 >>
rect 253 162 254 163 
<< m1 >>
rect 271 162 272 163 
<< m1 >>
rect 283 162 284 163 
<< m1 >>
rect 298 162 299 163 
<< m1 >>
rect 307 162 308 163 
<< m1 >>
rect 311 162 312 163 
<< m1 >>
rect 343 162 344 163 
<< m1 >>
rect 347 162 348 163 
<< m1 >>
rect 391 162 392 163 
<< m1 >>
rect 406 162 407 163 
<< m1 >>
rect 49 163 50 164 
<< m2 >>
rect 63 163 64 164 
<< m1 >>
rect 64 163 65 164 
<< m1 >>
rect 91 163 92 164 
<< m1 >>
rect 93 163 94 164 
<< m1 >>
rect 106 163 107 164 
<< m1 >>
rect 118 163 119 164 
<< m1 >>
rect 121 163 122 164 
<< m1 >>
rect 160 163 161 164 
<< m1 >>
rect 162 163 163 164 
<< m1 >>
rect 163 163 164 164 
<< m1 >>
rect 164 163 165 164 
<< m1 >>
rect 165 163 166 164 
<< m1 >>
rect 166 163 167 164 
<< m1 >>
rect 167 163 168 164 
<< m1 >>
rect 168 163 169 164 
<< m2 >>
rect 168 163 169 164 
<< m2c >>
rect 168 163 169 164 
<< m1 >>
rect 168 163 169 164 
<< m2 >>
rect 168 163 169 164 
<< m2 >>
rect 169 163 170 164 
<< m1 >>
rect 170 163 171 164 
<< m2 >>
rect 170 163 171 164 
<< m2 >>
rect 171 163 172 164 
<< m1 >>
rect 172 163 173 164 
<< m2 >>
rect 172 163 173 164 
<< m2c >>
rect 172 163 173 164 
<< m1 >>
rect 172 163 173 164 
<< m2 >>
rect 172 163 173 164 
<< m1 >>
rect 181 163 182 164 
<< m1 >>
rect 193 163 194 164 
<< m1 >>
rect 208 163 209 164 
<< m1 >>
rect 226 163 227 164 
<< m2 >>
rect 226 163 227 164 
<< m1 >>
rect 232 163 233 164 
<< m1 >>
rect 235 163 236 164 
<< m1 >>
rect 244 163 245 164 
<< m1 >>
rect 247 163 248 164 
<< m1 >>
rect 253 163 254 164 
<< m1 >>
rect 271 163 272 164 
<< m1 >>
rect 283 163 284 164 
<< m1 >>
rect 298 163 299 164 
<< m1 >>
rect 307 163 308 164 
<< m1 >>
rect 311 163 312 164 
<< m1 >>
rect 343 163 344 164 
<< m1 >>
rect 347 163 348 164 
<< m1 >>
rect 391 163 392 164 
<< m1 >>
rect 406 163 407 164 
<< m1 >>
rect 49 164 50 165 
<< m1 >>
rect 50 164 51 165 
<< m1 >>
rect 51 164 52 165 
<< m1 >>
rect 52 164 53 165 
<< m1 >>
rect 53 164 54 165 
<< m1 >>
rect 54 164 55 165 
<< m1 >>
rect 55 164 56 165 
<< m1 >>
rect 56 164 57 165 
<< m1 >>
rect 57 164 58 165 
<< m1 >>
rect 58 164 59 165 
<< m1 >>
rect 59 164 60 165 
<< m1 >>
rect 60 164 61 165 
<< m1 >>
rect 61 164 62 165 
<< m1 >>
rect 62 164 63 165 
<< m2 >>
rect 62 164 63 165 
<< m2c >>
rect 62 164 63 165 
<< m1 >>
rect 62 164 63 165 
<< m2 >>
rect 62 164 63 165 
<< m2 >>
rect 63 164 64 165 
<< m1 >>
rect 64 164 65 165 
<< m1 >>
rect 91 164 92 165 
<< m1 >>
rect 93 164 94 165 
<< m1 >>
rect 106 164 107 165 
<< m1 >>
rect 118 164 119 165 
<< m1 >>
rect 121 164 122 165 
<< m1 >>
rect 160 164 161 165 
<< m1 >>
rect 162 164 163 165 
<< m1 >>
rect 170 164 171 165 
<< m1 >>
rect 181 164 182 165 
<< m1 >>
rect 193 164 194 165 
<< m1 >>
rect 194 164 195 165 
<< m1 >>
rect 195 164 196 165 
<< m1 >>
rect 196 164 197 165 
<< m1 >>
rect 197 164 198 165 
<< m1 >>
rect 198 164 199 165 
<< m1 >>
rect 199 164 200 165 
<< m1 >>
rect 200 164 201 165 
<< m1 >>
rect 201 164 202 165 
<< m1 >>
rect 202 164 203 165 
<< m1 >>
rect 203 164 204 165 
<< m1 >>
rect 204 164 205 165 
<< m1 >>
rect 205 164 206 165 
<< m1 >>
rect 206 164 207 165 
<< m1 >>
rect 207 164 208 165 
<< m1 >>
rect 208 164 209 165 
<< m1 >>
rect 226 164 227 165 
<< m2 >>
rect 226 164 227 165 
<< m1 >>
rect 232 164 233 165 
<< m1 >>
rect 235 164 236 165 
<< m1 >>
rect 244 164 245 165 
<< m1 >>
rect 247 164 248 165 
<< m1 >>
rect 248 164 249 165 
<< m1 >>
rect 249 164 250 165 
<< m1 >>
rect 250 164 251 165 
<< m1 >>
rect 251 164 252 165 
<< m1 >>
rect 252 164 253 165 
<< m1 >>
rect 253 164 254 165 
<< m1 >>
rect 271 164 272 165 
<< m1 >>
rect 283 164 284 165 
<< m1 >>
rect 298 164 299 165 
<< m1 >>
rect 307 164 308 165 
<< m1 >>
rect 311 164 312 165 
<< m1 >>
rect 343 164 344 165 
<< m1 >>
rect 347 164 348 165 
<< m1 >>
rect 391 164 392 165 
<< m1 >>
rect 392 164 393 165 
<< m1 >>
rect 393 164 394 165 
<< m1 >>
rect 394 164 395 165 
<< m1 >>
rect 395 164 396 165 
<< m1 >>
rect 396 164 397 165 
<< m1 >>
rect 397 164 398 165 
<< m1 >>
rect 398 164 399 165 
<< m1 >>
rect 399 164 400 165 
<< m1 >>
rect 400 164 401 165 
<< m1 >>
rect 401 164 402 165 
<< m1 >>
rect 402 164 403 165 
<< m1 >>
rect 403 164 404 165 
<< m1 >>
rect 404 164 405 165 
<< m1 >>
rect 405 164 406 165 
<< m1 >>
rect 406 164 407 165 
<< m1 >>
rect 64 165 65 166 
<< m1 >>
rect 91 165 92 166 
<< m1 >>
rect 93 165 94 166 
<< m1 >>
rect 106 165 107 166 
<< m1 >>
rect 118 165 119 166 
<< m1 >>
rect 121 165 122 166 
<< m2 >>
rect 159 165 160 166 
<< m1 >>
rect 160 165 161 166 
<< m2 >>
rect 160 165 161 166 
<< m2 >>
rect 161 165 162 166 
<< m1 >>
rect 162 165 163 166 
<< m2 >>
rect 162 165 163 166 
<< m2c >>
rect 162 165 163 166 
<< m1 >>
rect 162 165 163 166 
<< m2 >>
rect 162 165 163 166 
<< m1 >>
rect 170 165 171 166 
<< m2 >>
rect 170 165 171 166 
<< m2c >>
rect 170 165 171 166 
<< m1 >>
rect 170 165 171 166 
<< m2 >>
rect 170 165 171 166 
<< m1 >>
rect 181 165 182 166 
<< m1 >>
rect 226 165 227 166 
<< m2 >>
rect 226 165 227 166 
<< m1 >>
rect 232 165 233 166 
<< m1 >>
rect 235 165 236 166 
<< m1 >>
rect 244 165 245 166 
<< m1 >>
rect 271 165 272 166 
<< m1 >>
rect 283 165 284 166 
<< m1 >>
rect 298 165 299 166 
<< m1 >>
rect 307 165 308 166 
<< m1 >>
rect 311 165 312 166 
<< m1 >>
rect 343 165 344 166 
<< m1 >>
rect 347 165 348 166 
<< m1 >>
rect 64 166 65 167 
<< m1 >>
rect 91 166 92 167 
<< m1 >>
rect 93 166 94 167 
<< m1 >>
rect 106 166 107 167 
<< m1 >>
rect 118 166 119 167 
<< m1 >>
rect 121 166 122 167 
<< m2 >>
rect 159 166 160 167 
<< m1 >>
rect 160 166 161 167 
<< m2 >>
rect 170 166 171 167 
<< m1 >>
rect 181 166 182 167 
<< m1 >>
rect 226 166 227 167 
<< m2 >>
rect 226 166 227 167 
<< m1 >>
rect 232 166 233 167 
<< m1 >>
rect 235 166 236 167 
<< m1 >>
rect 244 166 245 167 
<< m1 >>
rect 271 166 272 167 
<< m1 >>
rect 283 166 284 167 
<< m1 >>
rect 298 166 299 167 
<< m1 >>
rect 307 166 308 167 
<< m1 >>
rect 311 166 312 167 
<< m1 >>
rect 343 166 344 167 
<< m1 >>
rect 347 166 348 167 
<< m1 >>
rect 64 167 65 168 
<< m2 >>
rect 64 167 65 168 
<< m2c >>
rect 64 167 65 168 
<< m1 >>
rect 64 167 65 168 
<< m2 >>
rect 64 167 65 168 
<< m1 >>
rect 91 167 92 168 
<< m2 >>
rect 91 167 92 168 
<< m2c >>
rect 91 167 92 168 
<< m1 >>
rect 91 167 92 168 
<< m2 >>
rect 91 167 92 168 
<< m1 >>
rect 93 167 94 168 
<< m2 >>
rect 93 167 94 168 
<< m2c >>
rect 93 167 94 168 
<< m1 >>
rect 93 167 94 168 
<< m2 >>
rect 93 167 94 168 
<< m1 >>
rect 100 167 101 168 
<< m2 >>
rect 100 167 101 168 
<< m2c >>
rect 100 167 101 168 
<< m1 >>
rect 100 167 101 168 
<< m2 >>
rect 100 167 101 168 
<< m1 >>
rect 101 167 102 168 
<< m1 >>
rect 102 167 103 168 
<< m1 >>
rect 103 167 104 168 
<< m1 >>
rect 104 167 105 168 
<< m1 >>
rect 105 167 106 168 
<< m1 >>
rect 106 167 107 168 
<< m1 >>
rect 118 167 119 168 
<< m2 >>
rect 118 167 119 168 
<< m2c >>
rect 118 167 119 168 
<< m1 >>
rect 118 167 119 168 
<< m2 >>
rect 118 167 119 168 
<< m1 >>
rect 121 167 122 168 
<< m1 >>
rect 122 167 123 168 
<< m1 >>
rect 123 167 124 168 
<< m1 >>
rect 124 167 125 168 
<< m2 >>
rect 124 167 125 168 
<< m2c >>
rect 124 167 125 168 
<< m1 >>
rect 124 167 125 168 
<< m2 >>
rect 124 167 125 168 
<< m2 >>
rect 159 167 160 168 
<< m1 >>
rect 160 167 161 168 
<< m1 >>
rect 161 167 162 168 
<< m1 >>
rect 162 167 163 168 
<< m1 >>
rect 163 167 164 168 
<< m1 >>
rect 164 167 165 168 
<< m1 >>
rect 165 167 166 168 
<< m1 >>
rect 166 167 167 168 
<< m1 >>
rect 167 167 168 168 
<< m1 >>
rect 168 167 169 168 
<< m1 >>
rect 169 167 170 168 
<< m1 >>
rect 170 167 171 168 
<< m2 >>
rect 170 167 171 168 
<< m1 >>
rect 171 167 172 168 
<< m1 >>
rect 172 167 173 168 
<< m2 >>
rect 172 167 173 168 
<< m2c >>
rect 172 167 173 168 
<< m1 >>
rect 172 167 173 168 
<< m2 >>
rect 172 167 173 168 
<< m1 >>
rect 181 167 182 168 
<< m2 >>
rect 181 167 182 168 
<< m2c >>
rect 181 167 182 168 
<< m1 >>
rect 181 167 182 168 
<< m2 >>
rect 181 167 182 168 
<< m1 >>
rect 226 167 227 168 
<< m2 >>
rect 226 167 227 168 
<< m1 >>
rect 227 167 228 168 
<< m1 >>
rect 228 167 229 168 
<< m1 >>
rect 229 167 230 168 
<< m2 >>
rect 229 167 230 168 
<< m2c >>
rect 229 167 230 168 
<< m1 >>
rect 229 167 230 168 
<< m2 >>
rect 229 167 230 168 
<< m1 >>
rect 232 167 233 168 
<< m1 >>
rect 235 167 236 168 
<< m1 >>
rect 244 167 245 168 
<< m1 >>
rect 271 167 272 168 
<< m2 >>
rect 271 167 272 168 
<< m2c >>
rect 271 167 272 168 
<< m1 >>
rect 271 167 272 168 
<< m2 >>
rect 271 167 272 168 
<< m1 >>
rect 283 167 284 168 
<< m2 >>
rect 283 167 284 168 
<< m2c >>
rect 283 167 284 168 
<< m1 >>
rect 283 167 284 168 
<< m2 >>
rect 283 167 284 168 
<< m1 >>
rect 298 167 299 168 
<< m2 >>
rect 298 167 299 168 
<< m2c >>
rect 298 167 299 168 
<< m1 >>
rect 298 167 299 168 
<< m2 >>
rect 298 167 299 168 
<< m1 >>
rect 307 167 308 168 
<< m2 >>
rect 307 167 308 168 
<< m2c >>
rect 307 167 308 168 
<< m1 >>
rect 307 167 308 168 
<< m2 >>
rect 307 167 308 168 
<< m1 >>
rect 311 167 312 168 
<< m2 >>
rect 311 167 312 168 
<< m2c >>
rect 311 167 312 168 
<< m1 >>
rect 311 167 312 168 
<< m2 >>
rect 311 167 312 168 
<< m1 >>
rect 343 167 344 168 
<< m1 >>
rect 347 167 348 168 
<< m2 >>
rect 347 167 348 168 
<< m2c >>
rect 347 167 348 168 
<< m1 >>
rect 347 167 348 168 
<< m2 >>
rect 347 167 348 168 
<< m2 >>
rect 64 168 65 169 
<< m2 >>
rect 84 168 85 169 
<< m2 >>
rect 85 168 86 169 
<< m2 >>
rect 86 168 87 169 
<< m2 >>
rect 87 168 88 169 
<< m2 >>
rect 88 168 89 169 
<< m2 >>
rect 89 168 90 169 
<< m2 >>
rect 90 168 91 169 
<< m2 >>
rect 91 168 92 169 
<< m2 >>
rect 93 168 94 169 
<< m2 >>
rect 100 168 101 169 
<< m2 >>
rect 118 168 119 169 
<< m2 >>
rect 124 168 125 169 
<< m2 >>
rect 159 168 160 169 
<< m2 >>
rect 170 168 171 169 
<< m2 >>
rect 172 168 173 169 
<< m2 >>
rect 181 168 182 169 
<< m2 >>
rect 226 168 227 169 
<< m2 >>
rect 229 168 230 169 
<< m1 >>
rect 232 168 233 169 
<< m1 >>
rect 235 168 236 169 
<< m1 >>
rect 244 168 245 169 
<< m2 >>
rect 271 168 272 169 
<< m2 >>
rect 283 168 284 169 
<< m2 >>
rect 284 168 285 169 
<< m2 >>
rect 298 168 299 169 
<< m2 >>
rect 307 168 308 169 
<< m2 >>
rect 311 168 312 169 
<< m1 >>
rect 343 168 344 169 
<< m2 >>
rect 347 168 348 169 
<< m1 >>
rect 19 169 20 170 
<< m1 >>
rect 20 169 21 170 
<< m1 >>
rect 21 169 22 170 
<< m1 >>
rect 22 169 23 170 
<< m1 >>
rect 23 169 24 170 
<< m1 >>
rect 24 169 25 170 
<< m1 >>
rect 25 169 26 170 
<< m1 >>
rect 26 169 27 170 
<< m1 >>
rect 27 169 28 170 
<< m1 >>
rect 28 169 29 170 
<< m1 >>
rect 29 169 30 170 
<< m1 >>
rect 30 169 31 170 
<< m1 >>
rect 31 169 32 170 
<< m1 >>
rect 32 169 33 170 
<< m1 >>
rect 33 169 34 170 
<< m1 >>
rect 34 169 35 170 
<< m1 >>
rect 35 169 36 170 
<< m1 >>
rect 36 169 37 170 
<< m1 >>
rect 37 169 38 170 
<< m1 >>
rect 38 169 39 170 
<< m1 >>
rect 39 169 40 170 
<< m1 >>
rect 40 169 41 170 
<< m1 >>
rect 41 169 42 170 
<< m1 >>
rect 42 169 43 170 
<< m1 >>
rect 43 169 44 170 
<< m1 >>
rect 44 169 45 170 
<< m1 >>
rect 45 169 46 170 
<< m1 >>
rect 46 169 47 170 
<< m1 >>
rect 47 169 48 170 
<< m1 >>
rect 48 169 49 170 
<< m1 >>
rect 49 169 50 170 
<< m1 >>
rect 50 169 51 170 
<< m1 >>
rect 51 169 52 170 
<< m1 >>
rect 52 169 53 170 
<< m1 >>
rect 53 169 54 170 
<< m1 >>
rect 54 169 55 170 
<< m1 >>
rect 55 169 56 170 
<< m1 >>
rect 56 169 57 170 
<< m1 >>
rect 57 169 58 170 
<< m1 >>
rect 58 169 59 170 
<< m1 >>
rect 59 169 60 170 
<< m1 >>
rect 60 169 61 170 
<< m1 >>
rect 61 169 62 170 
<< m1 >>
rect 62 169 63 170 
<< m1 >>
rect 63 169 64 170 
<< m1 >>
rect 64 169 65 170 
<< m2 >>
rect 64 169 65 170 
<< m1 >>
rect 65 169 66 170 
<< m1 >>
rect 66 169 67 170 
<< m1 >>
rect 67 169 68 170 
<< m1 >>
rect 68 169 69 170 
<< m1 >>
rect 69 169 70 170 
<< m1 >>
rect 70 169 71 170 
<< m1 >>
rect 71 169 72 170 
<< m1 >>
rect 72 169 73 170 
<< m1 >>
rect 73 169 74 170 
<< m1 >>
rect 74 169 75 170 
<< m1 >>
rect 75 169 76 170 
<< m1 >>
rect 76 169 77 170 
<< m1 >>
rect 77 169 78 170 
<< m1 >>
rect 78 169 79 170 
<< m1 >>
rect 79 169 80 170 
<< m1 >>
rect 80 169 81 170 
<< m1 >>
rect 81 169 82 170 
<< m1 >>
rect 82 169 83 170 
<< m1 >>
rect 83 169 84 170 
<< m1 >>
rect 84 169 85 170 
<< m2 >>
rect 84 169 85 170 
<< m1 >>
rect 85 169 86 170 
<< m1 >>
rect 86 169 87 170 
<< m1 >>
rect 87 169 88 170 
<< m1 >>
rect 88 169 89 170 
<< m1 >>
rect 89 169 90 170 
<< m1 >>
rect 90 169 91 170 
<< m1 >>
rect 91 169 92 170 
<< m1 >>
rect 92 169 93 170 
<< m1 >>
rect 93 169 94 170 
<< m2 >>
rect 93 169 94 170 
<< m1 >>
rect 94 169 95 170 
<< m1 >>
rect 95 169 96 170 
<< m1 >>
rect 96 169 97 170 
<< m1 >>
rect 97 169 98 170 
<< m1 >>
rect 98 169 99 170 
<< m1 >>
rect 99 169 100 170 
<< m1 >>
rect 100 169 101 170 
<< m2 >>
rect 100 169 101 170 
<< m1 >>
rect 101 169 102 170 
<< m1 >>
rect 102 169 103 170 
<< m1 >>
rect 103 169 104 170 
<< m1 >>
rect 104 169 105 170 
<< m1 >>
rect 105 169 106 170 
<< m1 >>
rect 106 169 107 170 
<< m1 >>
rect 107 169 108 170 
<< m1 >>
rect 108 169 109 170 
<< m1 >>
rect 109 169 110 170 
<< m1 >>
rect 110 169 111 170 
<< m1 >>
rect 111 169 112 170 
<< m1 >>
rect 112 169 113 170 
<< m1 >>
rect 113 169 114 170 
<< m1 >>
rect 114 169 115 170 
<< m1 >>
rect 115 169 116 170 
<< m1 >>
rect 116 169 117 170 
<< m1 >>
rect 117 169 118 170 
<< m1 >>
rect 118 169 119 170 
<< m2 >>
rect 118 169 119 170 
<< m1 >>
rect 119 169 120 170 
<< m1 >>
rect 120 169 121 170 
<< m1 >>
rect 121 169 122 170 
<< m1 >>
rect 122 169 123 170 
<< m1 >>
rect 123 169 124 170 
<< m1 >>
rect 124 169 125 170 
<< m2 >>
rect 124 169 125 170 
<< m1 >>
rect 125 169 126 170 
<< m1 >>
rect 126 169 127 170 
<< m1 >>
rect 127 169 128 170 
<< m2 >>
rect 127 169 128 170 
<< m1 >>
rect 128 169 129 170 
<< m2 >>
rect 128 169 129 170 
<< m1 >>
rect 129 169 130 170 
<< m2 >>
rect 129 169 130 170 
<< m1 >>
rect 130 169 131 170 
<< m2 >>
rect 130 169 131 170 
<< m1 >>
rect 131 169 132 170 
<< m2 >>
rect 131 169 132 170 
<< m1 >>
rect 132 169 133 170 
<< m2 >>
rect 132 169 133 170 
<< m1 >>
rect 133 169 134 170 
<< m2 >>
rect 133 169 134 170 
<< m1 >>
rect 134 169 135 170 
<< m2 >>
rect 134 169 135 170 
<< m1 >>
rect 135 169 136 170 
<< m2 >>
rect 135 169 136 170 
<< m1 >>
rect 136 169 137 170 
<< m2 >>
rect 136 169 137 170 
<< m1 >>
rect 137 169 138 170 
<< m2 >>
rect 137 169 138 170 
<< m1 >>
rect 138 169 139 170 
<< m2 >>
rect 138 169 139 170 
<< m1 >>
rect 139 169 140 170 
<< m2 >>
rect 139 169 140 170 
<< m1 >>
rect 140 169 141 170 
<< m2 >>
rect 140 169 141 170 
<< m1 >>
rect 141 169 142 170 
<< m2 >>
rect 141 169 142 170 
<< m1 >>
rect 142 169 143 170 
<< m2 >>
rect 142 169 143 170 
<< m1 >>
rect 143 169 144 170 
<< m2 >>
rect 143 169 144 170 
<< m1 >>
rect 144 169 145 170 
<< m2 >>
rect 144 169 145 170 
<< m1 >>
rect 145 169 146 170 
<< m2 >>
rect 145 169 146 170 
<< m1 >>
rect 146 169 147 170 
<< m2 >>
rect 146 169 147 170 
<< m1 >>
rect 147 169 148 170 
<< m2 >>
rect 147 169 148 170 
<< m1 >>
rect 148 169 149 170 
<< m2 >>
rect 148 169 149 170 
<< m1 >>
rect 149 169 150 170 
<< m2 >>
rect 149 169 150 170 
<< m1 >>
rect 150 169 151 170 
<< m2 >>
rect 150 169 151 170 
<< m1 >>
rect 151 169 152 170 
<< m2 >>
rect 151 169 152 170 
<< m1 >>
rect 152 169 153 170 
<< m2 >>
rect 152 169 153 170 
<< m1 >>
rect 153 169 154 170 
<< m2 >>
rect 153 169 154 170 
<< m1 >>
rect 154 169 155 170 
<< m2 >>
rect 154 169 155 170 
<< m1 >>
rect 155 169 156 170 
<< m2 >>
rect 155 169 156 170 
<< m1 >>
rect 156 169 157 170 
<< m2 >>
rect 156 169 157 170 
<< m1 >>
rect 157 169 158 170 
<< m2 >>
rect 157 169 158 170 
<< m1 >>
rect 158 169 159 170 
<< m2 >>
rect 158 169 159 170 
<< m1 >>
rect 159 169 160 170 
<< m2 >>
rect 159 169 160 170 
<< m1 >>
rect 160 169 161 170 
<< m1 >>
rect 161 169 162 170 
<< m1 >>
rect 162 169 163 170 
<< m1 >>
rect 163 169 164 170 
<< m1 >>
rect 164 169 165 170 
<< m1 >>
rect 165 169 166 170 
<< m1 >>
rect 166 169 167 170 
<< m1 >>
rect 167 169 168 170 
<< m1 >>
rect 168 169 169 170 
<< m1 >>
rect 169 169 170 170 
<< m1 >>
rect 170 169 171 170 
<< m2 >>
rect 170 169 171 170 
<< m1 >>
rect 171 169 172 170 
<< m1 >>
rect 172 169 173 170 
<< m2 >>
rect 172 169 173 170 
<< m1 >>
rect 173 169 174 170 
<< m1 >>
rect 174 169 175 170 
<< m1 >>
rect 175 169 176 170 
<< m1 >>
rect 176 169 177 170 
<< m1 >>
rect 177 169 178 170 
<< m1 >>
rect 178 169 179 170 
<< m1 >>
rect 179 169 180 170 
<< m1 >>
rect 180 169 181 170 
<< m1 >>
rect 181 169 182 170 
<< m2 >>
rect 181 169 182 170 
<< m1 >>
rect 182 169 183 170 
<< m1 >>
rect 183 169 184 170 
<< m1 >>
rect 184 169 185 170 
<< m1 >>
rect 185 169 186 170 
<< m1 >>
rect 186 169 187 170 
<< m1 >>
rect 187 169 188 170 
<< m1 >>
rect 188 169 189 170 
<< m1 >>
rect 189 169 190 170 
<< m1 >>
rect 190 169 191 170 
<< m1 >>
rect 191 169 192 170 
<< m1 >>
rect 192 169 193 170 
<< m1 >>
rect 193 169 194 170 
<< m1 >>
rect 194 169 195 170 
<< m1 >>
rect 195 169 196 170 
<< m1 >>
rect 196 169 197 170 
<< m1 >>
rect 197 169 198 170 
<< m1 >>
rect 198 169 199 170 
<< m1 >>
rect 199 169 200 170 
<< m1 >>
rect 200 169 201 170 
<< m1 >>
rect 201 169 202 170 
<< m1 >>
rect 202 169 203 170 
<< m1 >>
rect 203 169 204 170 
<< m1 >>
rect 204 169 205 170 
<< m1 >>
rect 205 169 206 170 
<< m1 >>
rect 206 169 207 170 
<< m1 >>
rect 207 169 208 170 
<< m1 >>
rect 208 169 209 170 
<< m1 >>
rect 209 169 210 170 
<< m1 >>
rect 210 169 211 170 
<< m1 >>
rect 211 169 212 170 
<< m1 >>
rect 212 169 213 170 
<< m1 >>
rect 213 169 214 170 
<< m1 >>
rect 214 169 215 170 
<< m1 >>
rect 215 169 216 170 
<< m1 >>
rect 216 169 217 170 
<< m1 >>
rect 217 169 218 170 
<< m1 >>
rect 218 169 219 170 
<< m1 >>
rect 219 169 220 170 
<< m1 >>
rect 220 169 221 170 
<< m1 >>
rect 221 169 222 170 
<< m1 >>
rect 222 169 223 170 
<< m1 >>
rect 223 169 224 170 
<< m1 >>
rect 224 169 225 170 
<< m1 >>
rect 225 169 226 170 
<< m1 >>
rect 226 169 227 170 
<< m2 >>
rect 226 169 227 170 
<< m1 >>
rect 227 169 228 170 
<< m1 >>
rect 228 169 229 170 
<< m1 >>
rect 229 169 230 170 
<< m2 >>
rect 229 169 230 170 
<< m1 >>
rect 230 169 231 170 
<< m1 >>
rect 231 169 232 170 
<< m1 >>
rect 232 169 233 170 
<< m1 >>
rect 235 169 236 170 
<< m1 >>
rect 244 169 245 170 
<< m1 >>
rect 245 169 246 170 
<< m1 >>
rect 246 169 247 170 
<< m1 >>
rect 247 169 248 170 
<< m1 >>
rect 248 169 249 170 
<< m1 >>
rect 249 169 250 170 
<< m1 >>
rect 250 169 251 170 
<< m1 >>
rect 251 169 252 170 
<< m1 >>
rect 252 169 253 170 
<< m1 >>
rect 253 169 254 170 
<< m1 >>
rect 254 169 255 170 
<< m1 >>
rect 255 169 256 170 
<< m1 >>
rect 256 169 257 170 
<< m1 >>
rect 257 169 258 170 
<< m1 >>
rect 258 169 259 170 
<< m1 >>
rect 259 169 260 170 
<< m1 >>
rect 260 169 261 170 
<< m1 >>
rect 261 169 262 170 
<< m1 >>
rect 262 169 263 170 
<< m1 >>
rect 263 169 264 170 
<< m1 >>
rect 264 169 265 170 
<< m1 >>
rect 265 169 266 170 
<< m1 >>
rect 266 169 267 170 
<< m1 >>
rect 267 169 268 170 
<< m1 >>
rect 268 169 269 170 
<< m1 >>
rect 269 169 270 170 
<< m1 >>
rect 270 169 271 170 
<< m1 >>
rect 271 169 272 170 
<< m2 >>
rect 271 169 272 170 
<< m1 >>
rect 272 169 273 170 
<< m1 >>
rect 273 169 274 170 
<< m1 >>
rect 274 169 275 170 
<< m1 >>
rect 275 169 276 170 
<< m1 >>
rect 276 169 277 170 
<< m1 >>
rect 277 169 278 170 
<< m1 >>
rect 278 169 279 170 
<< m1 >>
rect 279 169 280 170 
<< m1 >>
rect 280 169 281 170 
<< m1 >>
rect 281 169 282 170 
<< m1 >>
rect 282 169 283 170 
<< m1 >>
rect 283 169 284 170 
<< m1 >>
rect 284 169 285 170 
<< m2 >>
rect 284 169 285 170 
<< m1 >>
rect 285 169 286 170 
<< m1 >>
rect 286 169 287 170 
<< m1 >>
rect 287 169 288 170 
<< m1 >>
rect 288 169 289 170 
<< m1 >>
rect 289 169 290 170 
<< m1 >>
rect 290 169 291 170 
<< m1 >>
rect 291 169 292 170 
<< m1 >>
rect 292 169 293 170 
<< m1 >>
rect 293 169 294 170 
<< m1 >>
rect 294 169 295 170 
<< m1 >>
rect 295 169 296 170 
<< m1 >>
rect 296 169 297 170 
<< m1 >>
rect 297 169 298 170 
<< m1 >>
rect 298 169 299 170 
<< m2 >>
rect 298 169 299 170 
<< m1 >>
rect 299 169 300 170 
<< m1 >>
rect 300 169 301 170 
<< m1 >>
rect 301 169 302 170 
<< m1 >>
rect 302 169 303 170 
<< m1 >>
rect 303 169 304 170 
<< m1 >>
rect 304 169 305 170 
<< m1 >>
rect 305 169 306 170 
<< m1 >>
rect 306 169 307 170 
<< m1 >>
rect 307 169 308 170 
<< m2 >>
rect 307 169 308 170 
<< m1 >>
rect 308 169 309 170 
<< m1 >>
rect 309 169 310 170 
<< m1 >>
rect 310 169 311 170 
<< m1 >>
rect 311 169 312 170 
<< m2 >>
rect 311 169 312 170 
<< m1 >>
rect 312 169 313 170 
<< m1 >>
rect 313 169 314 170 
<< m1 >>
rect 314 169 315 170 
<< m1 >>
rect 315 169 316 170 
<< m1 >>
rect 316 169 317 170 
<< m1 >>
rect 317 169 318 170 
<< m1 >>
rect 318 169 319 170 
<< m1 >>
rect 319 169 320 170 
<< m1 >>
rect 320 169 321 170 
<< m1 >>
rect 321 169 322 170 
<< m1 >>
rect 322 169 323 170 
<< m1 >>
rect 323 169 324 170 
<< m1 >>
rect 324 169 325 170 
<< m1 >>
rect 325 169 326 170 
<< m1 >>
rect 326 169 327 170 
<< m1 >>
rect 327 169 328 170 
<< m1 >>
rect 328 169 329 170 
<< m1 >>
rect 329 169 330 170 
<< m1 >>
rect 330 169 331 170 
<< m1 >>
rect 331 169 332 170 
<< m1 >>
rect 332 169 333 170 
<< m1 >>
rect 333 169 334 170 
<< m1 >>
rect 334 169 335 170 
<< m1 >>
rect 335 169 336 170 
<< m1 >>
rect 336 169 337 170 
<< m1 >>
rect 337 169 338 170 
<< m1 >>
rect 338 169 339 170 
<< m1 >>
rect 339 169 340 170 
<< m1 >>
rect 340 169 341 170 
<< m1 >>
rect 341 169 342 170 
<< m2 >>
rect 341 169 342 170 
<< m2c >>
rect 341 169 342 170 
<< m1 >>
rect 341 169 342 170 
<< m2 >>
rect 341 169 342 170 
<< m2 >>
rect 342 169 343 170 
<< m1 >>
rect 343 169 344 170 
<< m2 >>
rect 343 169 344 170 
<< m2 >>
rect 344 169 345 170 
<< m1 >>
rect 345 169 346 170 
<< m2 >>
rect 345 169 346 170 
<< m2c >>
rect 345 169 346 170 
<< m1 >>
rect 345 169 346 170 
<< m2 >>
rect 345 169 346 170 
<< m1 >>
rect 346 169 347 170 
<< m1 >>
rect 347 169 348 170 
<< m2 >>
rect 347 169 348 170 
<< m1 >>
rect 348 169 349 170 
<< m1 >>
rect 349 169 350 170 
<< m1 >>
rect 350 169 351 170 
<< m1 >>
rect 351 169 352 170 
<< m1 >>
rect 352 169 353 170 
<< m1 >>
rect 353 169 354 170 
<< m1 >>
rect 354 169 355 170 
<< m1 >>
rect 355 169 356 170 
<< m1 >>
rect 356 169 357 170 
<< m1 >>
rect 357 169 358 170 
<< m1 >>
rect 358 169 359 170 
<< m1 >>
rect 359 169 360 170 
<< m1 >>
rect 360 169 361 170 
<< m1 >>
rect 361 169 362 170 
<< m1 >>
rect 362 169 363 170 
<< m1 >>
rect 363 169 364 170 
<< m1 >>
rect 364 169 365 170 
<< m1 >>
rect 365 169 366 170 
<< m1 >>
rect 366 169 367 170 
<< m1 >>
rect 367 169 368 170 
<< m1 >>
rect 368 169 369 170 
<< m1 >>
rect 369 169 370 170 
<< m1 >>
rect 370 169 371 170 
<< m1 >>
rect 371 169 372 170 
<< m1 >>
rect 372 169 373 170 
<< m1 >>
rect 373 169 374 170 
<< m1 >>
rect 374 169 375 170 
<< m1 >>
rect 375 169 376 170 
<< m1 >>
rect 376 169 377 170 
<< m1 >>
rect 377 169 378 170 
<< m1 >>
rect 378 169 379 170 
<< m1 >>
rect 379 169 380 170 
<< m1 >>
rect 380 169 381 170 
<< m1 >>
rect 381 169 382 170 
<< m1 >>
rect 382 169 383 170 
<< m1 >>
rect 383 169 384 170 
<< m1 >>
rect 384 169 385 170 
<< m1 >>
rect 385 169 386 170 
<< m1 >>
rect 386 169 387 170 
<< m1 >>
rect 387 169 388 170 
<< m1 >>
rect 388 169 389 170 
<< m1 >>
rect 389 169 390 170 
<< m1 >>
rect 390 169 391 170 
<< m1 >>
rect 391 169 392 170 
<< m1 >>
rect 392 169 393 170 
<< m1 >>
rect 393 169 394 170 
<< m1 >>
rect 394 169 395 170 
<< m1 >>
rect 19 170 20 171 
<< m2 >>
rect 64 170 65 171 
<< m2 >>
rect 84 170 85 171 
<< m2 >>
rect 93 170 94 171 
<< m2 >>
rect 100 170 101 171 
<< m2 >>
rect 118 170 119 171 
<< m2 >>
rect 124 170 125 171 
<< m2 >>
rect 127 170 128 171 
<< m2 >>
rect 170 170 171 171 
<< m2 >>
rect 172 170 173 171 
<< m2 >>
rect 181 170 182 171 
<< m2 >>
rect 226 170 227 171 
<< m2 >>
rect 229 170 230 171 
<< m1 >>
rect 235 170 236 171 
<< m2 >>
rect 271 170 272 171 
<< m2 >>
rect 284 170 285 171 
<< m2 >>
rect 298 170 299 171 
<< m2 >>
rect 307 170 308 171 
<< m2 >>
rect 311 170 312 171 
<< m1 >>
rect 343 170 344 171 
<< m2 >>
rect 347 170 348 171 
<< m1 >>
rect 394 170 395 171 
<< m1 >>
rect 19 171 20 172 
<< m1 >>
rect 64 171 65 172 
<< m2 >>
rect 64 171 65 172 
<< m2c >>
rect 64 171 65 172 
<< m1 >>
rect 64 171 65 172 
<< m2 >>
rect 64 171 65 172 
<< m1 >>
rect 82 171 83 172 
<< m1 >>
rect 83 171 84 172 
<< m1 >>
rect 84 171 85 172 
<< m2 >>
rect 84 171 85 172 
<< m2c >>
rect 84 171 85 172 
<< m1 >>
rect 84 171 85 172 
<< m2 >>
rect 84 171 85 172 
<< m1 >>
rect 93 171 94 172 
<< m2 >>
rect 93 171 94 172 
<< m2c >>
rect 93 171 94 172 
<< m1 >>
rect 93 171 94 172 
<< m2 >>
rect 93 171 94 172 
<< m1 >>
rect 100 171 101 172 
<< m2 >>
rect 100 171 101 172 
<< m2c >>
rect 100 171 101 172 
<< m1 >>
rect 100 171 101 172 
<< m2 >>
rect 100 171 101 172 
<< m1 >>
rect 118 171 119 172 
<< m2 >>
rect 118 171 119 172 
<< m2c >>
rect 118 171 119 172 
<< m1 >>
rect 118 171 119 172 
<< m2 >>
rect 118 171 119 172 
<< m1 >>
rect 124 171 125 172 
<< m2 >>
rect 124 171 125 172 
<< m2c >>
rect 124 171 125 172 
<< m1 >>
rect 124 171 125 172 
<< m2 >>
rect 124 171 125 172 
<< m1 >>
rect 127 171 128 172 
<< m2 >>
rect 127 171 128 172 
<< m2c >>
rect 127 171 128 172 
<< m1 >>
rect 127 171 128 172 
<< m2 >>
rect 127 171 128 172 
<< m1 >>
rect 170 171 171 172 
<< m2 >>
rect 170 171 171 172 
<< m2c >>
rect 170 171 171 172 
<< m1 >>
rect 170 171 171 172 
<< m2 >>
rect 170 171 171 172 
<< m1 >>
rect 172 171 173 172 
<< m2 >>
rect 172 171 173 172 
<< m2c >>
rect 172 171 173 172 
<< m1 >>
rect 172 171 173 172 
<< m2 >>
rect 172 171 173 172 
<< m1 >>
rect 181 171 182 172 
<< m2 >>
rect 181 171 182 172 
<< m2c >>
rect 181 171 182 172 
<< m1 >>
rect 181 171 182 172 
<< m2 >>
rect 181 171 182 172 
<< m1 >>
rect 226 171 227 172 
<< m2 >>
rect 226 171 227 172 
<< m2c >>
rect 226 171 227 172 
<< m1 >>
rect 226 171 227 172 
<< m2 >>
rect 226 171 227 172 
<< m1 >>
rect 229 171 230 172 
<< m2 >>
rect 229 171 230 172 
<< m2c >>
rect 229 171 230 172 
<< m1 >>
rect 229 171 230 172 
<< m2 >>
rect 229 171 230 172 
<< m1 >>
rect 235 171 236 172 
<< m1 >>
rect 271 171 272 172 
<< m2 >>
rect 271 171 272 172 
<< m2c >>
rect 271 171 272 172 
<< m1 >>
rect 271 171 272 172 
<< m2 >>
rect 271 171 272 172 
<< m1 >>
rect 284 171 285 172 
<< m2 >>
rect 284 171 285 172 
<< m2c >>
rect 284 171 285 172 
<< m1 >>
rect 284 171 285 172 
<< m2 >>
rect 284 171 285 172 
<< m1 >>
rect 285 171 286 172 
<< m1 >>
rect 286 171 287 172 
<< m1 >>
rect 287 171 288 172 
<< m1 >>
rect 288 171 289 172 
<< m1 >>
rect 289 171 290 172 
<< m1 >>
rect 298 171 299 172 
<< m2 >>
rect 298 171 299 172 
<< m2c >>
rect 298 171 299 172 
<< m1 >>
rect 298 171 299 172 
<< m2 >>
rect 298 171 299 172 
<< m1 >>
rect 307 171 308 172 
<< m2 >>
rect 307 171 308 172 
<< m2c >>
rect 307 171 308 172 
<< m1 >>
rect 307 171 308 172 
<< m2 >>
rect 307 171 308 172 
<< m1 >>
rect 311 171 312 172 
<< m2 >>
rect 311 171 312 172 
<< m2c >>
rect 311 171 312 172 
<< m1 >>
rect 311 171 312 172 
<< m2 >>
rect 311 171 312 172 
<< m1 >>
rect 343 171 344 172 
<< m1 >>
rect 347 171 348 172 
<< m2 >>
rect 347 171 348 172 
<< m2c >>
rect 347 171 348 172 
<< m1 >>
rect 347 171 348 172 
<< m2 >>
rect 347 171 348 172 
<< m1 >>
rect 394 171 395 172 
<< m1 >>
rect 19 172 20 173 
<< m1 >>
rect 64 172 65 173 
<< m1 >>
rect 82 172 83 173 
<< m1 >>
rect 93 172 94 173 
<< m1 >>
rect 100 172 101 173 
<< m1 >>
rect 118 172 119 173 
<< m1 >>
rect 124 172 125 173 
<< m1 >>
rect 127 172 128 173 
<< m1 >>
rect 170 172 171 173 
<< m1 >>
rect 172 172 173 173 
<< m1 >>
rect 181 172 182 173 
<< m1 >>
rect 226 172 227 173 
<< m1 >>
rect 229 172 230 173 
<< m1 >>
rect 235 172 236 173 
<< m1 >>
rect 271 172 272 173 
<< m1 >>
rect 289 172 290 173 
<< m1 >>
rect 298 172 299 173 
<< m1 >>
rect 307 172 308 173 
<< m1 >>
rect 311 172 312 173 
<< m1 >>
rect 343 172 344 173 
<< m1 >>
rect 347 172 348 173 
<< m1 >>
rect 394 172 395 173 
<< m1 >>
rect 19 173 20 174 
<< m1 >>
rect 64 173 65 174 
<< m1 >>
rect 82 173 83 174 
<< m1 >>
rect 93 173 94 174 
<< m1 >>
rect 100 173 101 174 
<< m1 >>
rect 118 173 119 174 
<< m1 >>
rect 124 173 125 174 
<< m1 >>
rect 127 173 128 174 
<< m1 >>
rect 170 173 171 174 
<< m1 >>
rect 172 173 173 174 
<< m1 >>
rect 181 173 182 174 
<< m1 >>
rect 226 173 227 174 
<< m1 >>
rect 229 173 230 174 
<< m1 >>
rect 235 173 236 174 
<< m1 >>
rect 271 173 272 174 
<< m1 >>
rect 289 173 290 174 
<< m1 >>
rect 290 173 291 174 
<< m1 >>
rect 291 173 292 174 
<< m1 >>
rect 292 173 293 174 
<< m1 >>
rect 293 173 294 174 
<< m1 >>
rect 294 173 295 174 
<< m1 >>
rect 295 173 296 174 
<< m1 >>
rect 296 173 297 174 
<< m2 >>
rect 296 173 297 174 
<< m2c >>
rect 296 173 297 174 
<< m1 >>
rect 296 173 297 174 
<< m2 >>
rect 296 173 297 174 
<< m2 >>
rect 297 173 298 174 
<< m1 >>
rect 298 173 299 174 
<< m1 >>
rect 307 173 308 174 
<< m1 >>
rect 311 173 312 174 
<< m1 >>
rect 343 173 344 174 
<< m1 >>
rect 347 173 348 174 
<< m1 >>
rect 394 173 395 174 
<< pdiffusion >>
rect 12 174 13 175 
<< pdiffusion >>
rect 13 174 14 175 
<< pdiffusion >>
rect 14 174 15 175 
<< pdiffusion >>
rect 15 174 16 175 
<< pdiffusion >>
rect 16 174 17 175 
<< pdiffusion >>
rect 17 174 18 175 
<< m1 >>
rect 19 174 20 175 
<< pdiffusion >>
rect 30 174 31 175 
<< pdiffusion >>
rect 31 174 32 175 
<< pdiffusion >>
rect 32 174 33 175 
<< pdiffusion >>
rect 33 174 34 175 
<< pdiffusion >>
rect 34 174 35 175 
<< pdiffusion >>
rect 35 174 36 175 
<< pdiffusion >>
rect 48 174 49 175 
<< pdiffusion >>
rect 49 174 50 175 
<< pdiffusion >>
rect 50 174 51 175 
<< pdiffusion >>
rect 51 174 52 175 
<< pdiffusion >>
rect 52 174 53 175 
<< pdiffusion >>
rect 53 174 54 175 
<< m1 >>
rect 64 174 65 175 
<< pdiffusion >>
rect 66 174 67 175 
<< pdiffusion >>
rect 67 174 68 175 
<< pdiffusion >>
rect 68 174 69 175 
<< pdiffusion >>
rect 69 174 70 175 
<< pdiffusion >>
rect 70 174 71 175 
<< pdiffusion >>
rect 71 174 72 175 
<< m1 >>
rect 82 174 83 175 
<< pdiffusion >>
rect 84 174 85 175 
<< pdiffusion >>
rect 85 174 86 175 
<< pdiffusion >>
rect 86 174 87 175 
<< pdiffusion >>
rect 87 174 88 175 
<< pdiffusion >>
rect 88 174 89 175 
<< pdiffusion >>
rect 89 174 90 175 
<< m1 >>
rect 93 174 94 175 
<< m1 >>
rect 100 174 101 175 
<< pdiffusion >>
rect 102 174 103 175 
<< pdiffusion >>
rect 103 174 104 175 
<< pdiffusion >>
rect 104 174 105 175 
<< pdiffusion >>
rect 105 174 106 175 
<< pdiffusion >>
rect 106 174 107 175 
<< pdiffusion >>
rect 107 174 108 175 
<< m1 >>
rect 118 174 119 175 
<< pdiffusion >>
rect 120 174 121 175 
<< pdiffusion >>
rect 121 174 122 175 
<< pdiffusion >>
rect 122 174 123 175 
<< pdiffusion >>
rect 123 174 124 175 
<< m1 >>
rect 124 174 125 175 
<< pdiffusion >>
rect 124 174 125 175 
<< pdiffusion >>
rect 125 174 126 175 
<< m1 >>
rect 127 174 128 175 
<< pdiffusion >>
rect 138 174 139 175 
<< pdiffusion >>
rect 139 174 140 175 
<< pdiffusion >>
rect 140 174 141 175 
<< pdiffusion >>
rect 141 174 142 175 
<< pdiffusion >>
rect 142 174 143 175 
<< pdiffusion >>
rect 143 174 144 175 
<< pdiffusion >>
rect 156 174 157 175 
<< pdiffusion >>
rect 157 174 158 175 
<< pdiffusion >>
rect 158 174 159 175 
<< pdiffusion >>
rect 159 174 160 175 
<< pdiffusion >>
rect 160 174 161 175 
<< pdiffusion >>
rect 161 174 162 175 
<< m1 >>
rect 170 174 171 175 
<< m1 >>
rect 172 174 173 175 
<< pdiffusion >>
rect 174 174 175 175 
<< pdiffusion >>
rect 175 174 176 175 
<< pdiffusion >>
rect 176 174 177 175 
<< pdiffusion >>
rect 177 174 178 175 
<< pdiffusion >>
rect 178 174 179 175 
<< pdiffusion >>
rect 179 174 180 175 
<< m1 >>
rect 181 174 182 175 
<< pdiffusion >>
rect 192 174 193 175 
<< pdiffusion >>
rect 193 174 194 175 
<< pdiffusion >>
rect 194 174 195 175 
<< pdiffusion >>
rect 195 174 196 175 
<< pdiffusion >>
rect 196 174 197 175 
<< pdiffusion >>
rect 197 174 198 175 
<< pdiffusion >>
rect 210 174 211 175 
<< pdiffusion >>
rect 211 174 212 175 
<< pdiffusion >>
rect 212 174 213 175 
<< pdiffusion >>
rect 213 174 214 175 
<< pdiffusion >>
rect 214 174 215 175 
<< pdiffusion >>
rect 215 174 216 175 
<< m1 >>
rect 226 174 227 175 
<< pdiffusion >>
rect 228 174 229 175 
<< m1 >>
rect 229 174 230 175 
<< pdiffusion >>
rect 229 174 230 175 
<< pdiffusion >>
rect 230 174 231 175 
<< pdiffusion >>
rect 231 174 232 175 
<< pdiffusion >>
rect 232 174 233 175 
<< pdiffusion >>
rect 233 174 234 175 
<< m1 >>
rect 235 174 236 175 
<< pdiffusion >>
rect 246 174 247 175 
<< pdiffusion >>
rect 247 174 248 175 
<< pdiffusion >>
rect 248 174 249 175 
<< pdiffusion >>
rect 249 174 250 175 
<< pdiffusion >>
rect 250 174 251 175 
<< pdiffusion >>
rect 251 174 252 175 
<< pdiffusion >>
rect 264 174 265 175 
<< pdiffusion >>
rect 265 174 266 175 
<< pdiffusion >>
rect 266 174 267 175 
<< pdiffusion >>
rect 267 174 268 175 
<< pdiffusion >>
rect 268 174 269 175 
<< pdiffusion >>
rect 269 174 270 175 
<< m1 >>
rect 271 174 272 175 
<< pdiffusion >>
rect 282 174 283 175 
<< pdiffusion >>
rect 283 174 284 175 
<< pdiffusion >>
rect 284 174 285 175 
<< pdiffusion >>
rect 285 174 286 175 
<< pdiffusion >>
rect 286 174 287 175 
<< pdiffusion >>
rect 287 174 288 175 
<< m2 >>
rect 297 174 298 175 
<< m1 >>
rect 298 174 299 175 
<< pdiffusion >>
rect 300 174 301 175 
<< pdiffusion >>
rect 301 174 302 175 
<< pdiffusion >>
rect 302 174 303 175 
<< pdiffusion >>
rect 303 174 304 175 
<< pdiffusion >>
rect 304 174 305 175 
<< pdiffusion >>
rect 305 174 306 175 
<< m1 >>
rect 307 174 308 175 
<< m1 >>
rect 311 174 312 175 
<< pdiffusion >>
rect 336 174 337 175 
<< pdiffusion >>
rect 337 174 338 175 
<< pdiffusion >>
rect 338 174 339 175 
<< pdiffusion >>
rect 339 174 340 175 
<< pdiffusion >>
rect 340 174 341 175 
<< pdiffusion >>
rect 341 174 342 175 
<< m1 >>
rect 343 174 344 175 
<< m1 >>
rect 347 174 348 175 
<< pdiffusion >>
rect 354 174 355 175 
<< pdiffusion >>
rect 355 174 356 175 
<< pdiffusion >>
rect 356 174 357 175 
<< pdiffusion >>
rect 357 174 358 175 
<< pdiffusion >>
rect 358 174 359 175 
<< pdiffusion >>
rect 359 174 360 175 
<< pdiffusion >>
rect 372 174 373 175 
<< pdiffusion >>
rect 373 174 374 175 
<< pdiffusion >>
rect 374 174 375 175 
<< pdiffusion >>
rect 375 174 376 175 
<< pdiffusion >>
rect 376 174 377 175 
<< pdiffusion >>
rect 377 174 378 175 
<< pdiffusion >>
rect 390 174 391 175 
<< pdiffusion >>
rect 391 174 392 175 
<< pdiffusion >>
rect 392 174 393 175 
<< pdiffusion >>
rect 393 174 394 175 
<< m1 >>
rect 394 174 395 175 
<< pdiffusion >>
rect 394 174 395 175 
<< pdiffusion >>
rect 395 174 396 175 
<< pdiffusion >>
rect 408 174 409 175 
<< pdiffusion >>
rect 409 174 410 175 
<< pdiffusion >>
rect 410 174 411 175 
<< pdiffusion >>
rect 411 174 412 175 
<< pdiffusion >>
rect 412 174 413 175 
<< pdiffusion >>
rect 413 174 414 175 
<< pdiffusion >>
rect 426 174 427 175 
<< pdiffusion >>
rect 427 174 428 175 
<< pdiffusion >>
rect 428 174 429 175 
<< pdiffusion >>
rect 429 174 430 175 
<< pdiffusion >>
rect 430 174 431 175 
<< pdiffusion >>
rect 431 174 432 175 
<< pdiffusion >>
rect 12 175 13 176 
<< pdiffusion >>
rect 13 175 14 176 
<< pdiffusion >>
rect 14 175 15 176 
<< pdiffusion >>
rect 15 175 16 176 
<< pdiffusion >>
rect 16 175 17 176 
<< pdiffusion >>
rect 17 175 18 176 
<< m1 >>
rect 19 175 20 176 
<< pdiffusion >>
rect 30 175 31 176 
<< pdiffusion >>
rect 31 175 32 176 
<< pdiffusion >>
rect 32 175 33 176 
<< pdiffusion >>
rect 33 175 34 176 
<< pdiffusion >>
rect 34 175 35 176 
<< pdiffusion >>
rect 35 175 36 176 
<< pdiffusion >>
rect 48 175 49 176 
<< pdiffusion >>
rect 49 175 50 176 
<< pdiffusion >>
rect 50 175 51 176 
<< pdiffusion >>
rect 51 175 52 176 
<< pdiffusion >>
rect 52 175 53 176 
<< pdiffusion >>
rect 53 175 54 176 
<< m1 >>
rect 64 175 65 176 
<< pdiffusion >>
rect 66 175 67 176 
<< pdiffusion >>
rect 67 175 68 176 
<< pdiffusion >>
rect 68 175 69 176 
<< pdiffusion >>
rect 69 175 70 176 
<< pdiffusion >>
rect 70 175 71 176 
<< pdiffusion >>
rect 71 175 72 176 
<< m1 >>
rect 82 175 83 176 
<< pdiffusion >>
rect 84 175 85 176 
<< pdiffusion >>
rect 85 175 86 176 
<< pdiffusion >>
rect 86 175 87 176 
<< pdiffusion >>
rect 87 175 88 176 
<< pdiffusion >>
rect 88 175 89 176 
<< pdiffusion >>
rect 89 175 90 176 
<< m1 >>
rect 93 175 94 176 
<< m1 >>
rect 100 175 101 176 
<< pdiffusion >>
rect 102 175 103 176 
<< pdiffusion >>
rect 103 175 104 176 
<< pdiffusion >>
rect 104 175 105 176 
<< pdiffusion >>
rect 105 175 106 176 
<< pdiffusion >>
rect 106 175 107 176 
<< pdiffusion >>
rect 107 175 108 176 
<< m1 >>
rect 118 175 119 176 
<< pdiffusion >>
rect 120 175 121 176 
<< pdiffusion >>
rect 121 175 122 176 
<< pdiffusion >>
rect 122 175 123 176 
<< pdiffusion >>
rect 123 175 124 176 
<< pdiffusion >>
rect 124 175 125 176 
<< pdiffusion >>
rect 125 175 126 176 
<< m1 >>
rect 127 175 128 176 
<< pdiffusion >>
rect 138 175 139 176 
<< pdiffusion >>
rect 139 175 140 176 
<< pdiffusion >>
rect 140 175 141 176 
<< pdiffusion >>
rect 141 175 142 176 
<< pdiffusion >>
rect 142 175 143 176 
<< pdiffusion >>
rect 143 175 144 176 
<< pdiffusion >>
rect 156 175 157 176 
<< pdiffusion >>
rect 157 175 158 176 
<< pdiffusion >>
rect 158 175 159 176 
<< pdiffusion >>
rect 159 175 160 176 
<< pdiffusion >>
rect 160 175 161 176 
<< pdiffusion >>
rect 161 175 162 176 
<< m1 >>
rect 170 175 171 176 
<< m1 >>
rect 172 175 173 176 
<< pdiffusion >>
rect 174 175 175 176 
<< pdiffusion >>
rect 175 175 176 176 
<< pdiffusion >>
rect 176 175 177 176 
<< pdiffusion >>
rect 177 175 178 176 
<< pdiffusion >>
rect 178 175 179 176 
<< pdiffusion >>
rect 179 175 180 176 
<< m1 >>
rect 181 175 182 176 
<< pdiffusion >>
rect 192 175 193 176 
<< pdiffusion >>
rect 193 175 194 176 
<< pdiffusion >>
rect 194 175 195 176 
<< pdiffusion >>
rect 195 175 196 176 
<< pdiffusion >>
rect 196 175 197 176 
<< pdiffusion >>
rect 197 175 198 176 
<< pdiffusion >>
rect 210 175 211 176 
<< pdiffusion >>
rect 211 175 212 176 
<< pdiffusion >>
rect 212 175 213 176 
<< pdiffusion >>
rect 213 175 214 176 
<< pdiffusion >>
rect 214 175 215 176 
<< pdiffusion >>
rect 215 175 216 176 
<< m1 >>
rect 226 175 227 176 
<< pdiffusion >>
rect 228 175 229 176 
<< pdiffusion >>
rect 229 175 230 176 
<< pdiffusion >>
rect 230 175 231 176 
<< pdiffusion >>
rect 231 175 232 176 
<< pdiffusion >>
rect 232 175 233 176 
<< pdiffusion >>
rect 233 175 234 176 
<< m1 >>
rect 235 175 236 176 
<< pdiffusion >>
rect 246 175 247 176 
<< pdiffusion >>
rect 247 175 248 176 
<< pdiffusion >>
rect 248 175 249 176 
<< pdiffusion >>
rect 249 175 250 176 
<< pdiffusion >>
rect 250 175 251 176 
<< pdiffusion >>
rect 251 175 252 176 
<< pdiffusion >>
rect 264 175 265 176 
<< pdiffusion >>
rect 265 175 266 176 
<< pdiffusion >>
rect 266 175 267 176 
<< pdiffusion >>
rect 267 175 268 176 
<< pdiffusion >>
rect 268 175 269 176 
<< pdiffusion >>
rect 269 175 270 176 
<< m1 >>
rect 271 175 272 176 
<< pdiffusion >>
rect 282 175 283 176 
<< pdiffusion >>
rect 283 175 284 176 
<< pdiffusion >>
rect 284 175 285 176 
<< pdiffusion >>
rect 285 175 286 176 
<< pdiffusion >>
rect 286 175 287 176 
<< pdiffusion >>
rect 287 175 288 176 
<< m2 >>
rect 297 175 298 176 
<< m1 >>
rect 298 175 299 176 
<< pdiffusion >>
rect 300 175 301 176 
<< pdiffusion >>
rect 301 175 302 176 
<< pdiffusion >>
rect 302 175 303 176 
<< pdiffusion >>
rect 303 175 304 176 
<< pdiffusion >>
rect 304 175 305 176 
<< pdiffusion >>
rect 305 175 306 176 
<< m1 >>
rect 307 175 308 176 
<< m1 >>
rect 311 175 312 176 
<< pdiffusion >>
rect 336 175 337 176 
<< pdiffusion >>
rect 337 175 338 176 
<< pdiffusion >>
rect 338 175 339 176 
<< pdiffusion >>
rect 339 175 340 176 
<< pdiffusion >>
rect 340 175 341 176 
<< pdiffusion >>
rect 341 175 342 176 
<< m1 >>
rect 343 175 344 176 
<< m1 >>
rect 347 175 348 176 
<< pdiffusion >>
rect 354 175 355 176 
<< pdiffusion >>
rect 355 175 356 176 
<< pdiffusion >>
rect 356 175 357 176 
<< pdiffusion >>
rect 357 175 358 176 
<< pdiffusion >>
rect 358 175 359 176 
<< pdiffusion >>
rect 359 175 360 176 
<< pdiffusion >>
rect 372 175 373 176 
<< pdiffusion >>
rect 373 175 374 176 
<< pdiffusion >>
rect 374 175 375 176 
<< pdiffusion >>
rect 375 175 376 176 
<< pdiffusion >>
rect 376 175 377 176 
<< pdiffusion >>
rect 377 175 378 176 
<< pdiffusion >>
rect 390 175 391 176 
<< pdiffusion >>
rect 391 175 392 176 
<< pdiffusion >>
rect 392 175 393 176 
<< pdiffusion >>
rect 393 175 394 176 
<< pdiffusion >>
rect 394 175 395 176 
<< pdiffusion >>
rect 395 175 396 176 
<< pdiffusion >>
rect 408 175 409 176 
<< pdiffusion >>
rect 409 175 410 176 
<< pdiffusion >>
rect 410 175 411 176 
<< pdiffusion >>
rect 411 175 412 176 
<< pdiffusion >>
rect 412 175 413 176 
<< pdiffusion >>
rect 413 175 414 176 
<< pdiffusion >>
rect 426 175 427 176 
<< pdiffusion >>
rect 427 175 428 176 
<< pdiffusion >>
rect 428 175 429 176 
<< pdiffusion >>
rect 429 175 430 176 
<< pdiffusion >>
rect 430 175 431 176 
<< pdiffusion >>
rect 431 175 432 176 
<< pdiffusion >>
rect 12 176 13 177 
<< pdiffusion >>
rect 13 176 14 177 
<< pdiffusion >>
rect 14 176 15 177 
<< pdiffusion >>
rect 15 176 16 177 
<< pdiffusion >>
rect 16 176 17 177 
<< pdiffusion >>
rect 17 176 18 177 
<< m1 >>
rect 19 176 20 177 
<< pdiffusion >>
rect 30 176 31 177 
<< pdiffusion >>
rect 31 176 32 177 
<< pdiffusion >>
rect 32 176 33 177 
<< pdiffusion >>
rect 33 176 34 177 
<< pdiffusion >>
rect 34 176 35 177 
<< pdiffusion >>
rect 35 176 36 177 
<< pdiffusion >>
rect 48 176 49 177 
<< pdiffusion >>
rect 49 176 50 177 
<< pdiffusion >>
rect 50 176 51 177 
<< pdiffusion >>
rect 51 176 52 177 
<< pdiffusion >>
rect 52 176 53 177 
<< pdiffusion >>
rect 53 176 54 177 
<< m1 >>
rect 64 176 65 177 
<< pdiffusion >>
rect 66 176 67 177 
<< pdiffusion >>
rect 67 176 68 177 
<< pdiffusion >>
rect 68 176 69 177 
<< pdiffusion >>
rect 69 176 70 177 
<< pdiffusion >>
rect 70 176 71 177 
<< pdiffusion >>
rect 71 176 72 177 
<< m1 >>
rect 82 176 83 177 
<< pdiffusion >>
rect 84 176 85 177 
<< pdiffusion >>
rect 85 176 86 177 
<< pdiffusion >>
rect 86 176 87 177 
<< pdiffusion >>
rect 87 176 88 177 
<< pdiffusion >>
rect 88 176 89 177 
<< pdiffusion >>
rect 89 176 90 177 
<< m1 >>
rect 93 176 94 177 
<< m1 >>
rect 100 176 101 177 
<< pdiffusion >>
rect 102 176 103 177 
<< pdiffusion >>
rect 103 176 104 177 
<< pdiffusion >>
rect 104 176 105 177 
<< pdiffusion >>
rect 105 176 106 177 
<< pdiffusion >>
rect 106 176 107 177 
<< pdiffusion >>
rect 107 176 108 177 
<< m1 >>
rect 118 176 119 177 
<< pdiffusion >>
rect 120 176 121 177 
<< pdiffusion >>
rect 121 176 122 177 
<< pdiffusion >>
rect 122 176 123 177 
<< pdiffusion >>
rect 123 176 124 177 
<< pdiffusion >>
rect 124 176 125 177 
<< pdiffusion >>
rect 125 176 126 177 
<< m1 >>
rect 127 176 128 177 
<< pdiffusion >>
rect 138 176 139 177 
<< pdiffusion >>
rect 139 176 140 177 
<< pdiffusion >>
rect 140 176 141 177 
<< pdiffusion >>
rect 141 176 142 177 
<< pdiffusion >>
rect 142 176 143 177 
<< pdiffusion >>
rect 143 176 144 177 
<< pdiffusion >>
rect 156 176 157 177 
<< pdiffusion >>
rect 157 176 158 177 
<< pdiffusion >>
rect 158 176 159 177 
<< pdiffusion >>
rect 159 176 160 177 
<< pdiffusion >>
rect 160 176 161 177 
<< pdiffusion >>
rect 161 176 162 177 
<< m1 >>
rect 170 176 171 177 
<< m1 >>
rect 172 176 173 177 
<< pdiffusion >>
rect 174 176 175 177 
<< pdiffusion >>
rect 175 176 176 177 
<< pdiffusion >>
rect 176 176 177 177 
<< pdiffusion >>
rect 177 176 178 177 
<< pdiffusion >>
rect 178 176 179 177 
<< pdiffusion >>
rect 179 176 180 177 
<< m1 >>
rect 181 176 182 177 
<< pdiffusion >>
rect 192 176 193 177 
<< pdiffusion >>
rect 193 176 194 177 
<< pdiffusion >>
rect 194 176 195 177 
<< pdiffusion >>
rect 195 176 196 177 
<< pdiffusion >>
rect 196 176 197 177 
<< pdiffusion >>
rect 197 176 198 177 
<< pdiffusion >>
rect 210 176 211 177 
<< pdiffusion >>
rect 211 176 212 177 
<< pdiffusion >>
rect 212 176 213 177 
<< pdiffusion >>
rect 213 176 214 177 
<< pdiffusion >>
rect 214 176 215 177 
<< pdiffusion >>
rect 215 176 216 177 
<< m1 >>
rect 226 176 227 177 
<< pdiffusion >>
rect 228 176 229 177 
<< pdiffusion >>
rect 229 176 230 177 
<< pdiffusion >>
rect 230 176 231 177 
<< pdiffusion >>
rect 231 176 232 177 
<< pdiffusion >>
rect 232 176 233 177 
<< pdiffusion >>
rect 233 176 234 177 
<< m1 >>
rect 235 176 236 177 
<< pdiffusion >>
rect 246 176 247 177 
<< pdiffusion >>
rect 247 176 248 177 
<< pdiffusion >>
rect 248 176 249 177 
<< pdiffusion >>
rect 249 176 250 177 
<< pdiffusion >>
rect 250 176 251 177 
<< pdiffusion >>
rect 251 176 252 177 
<< pdiffusion >>
rect 264 176 265 177 
<< pdiffusion >>
rect 265 176 266 177 
<< pdiffusion >>
rect 266 176 267 177 
<< pdiffusion >>
rect 267 176 268 177 
<< pdiffusion >>
rect 268 176 269 177 
<< pdiffusion >>
rect 269 176 270 177 
<< m1 >>
rect 271 176 272 177 
<< pdiffusion >>
rect 282 176 283 177 
<< pdiffusion >>
rect 283 176 284 177 
<< pdiffusion >>
rect 284 176 285 177 
<< pdiffusion >>
rect 285 176 286 177 
<< pdiffusion >>
rect 286 176 287 177 
<< pdiffusion >>
rect 287 176 288 177 
<< m2 >>
rect 297 176 298 177 
<< m1 >>
rect 298 176 299 177 
<< pdiffusion >>
rect 300 176 301 177 
<< pdiffusion >>
rect 301 176 302 177 
<< pdiffusion >>
rect 302 176 303 177 
<< pdiffusion >>
rect 303 176 304 177 
<< pdiffusion >>
rect 304 176 305 177 
<< pdiffusion >>
rect 305 176 306 177 
<< m1 >>
rect 307 176 308 177 
<< m1 >>
rect 311 176 312 177 
<< pdiffusion >>
rect 336 176 337 177 
<< pdiffusion >>
rect 337 176 338 177 
<< pdiffusion >>
rect 338 176 339 177 
<< pdiffusion >>
rect 339 176 340 177 
<< pdiffusion >>
rect 340 176 341 177 
<< pdiffusion >>
rect 341 176 342 177 
<< m1 >>
rect 343 176 344 177 
<< m1 >>
rect 347 176 348 177 
<< pdiffusion >>
rect 354 176 355 177 
<< pdiffusion >>
rect 355 176 356 177 
<< pdiffusion >>
rect 356 176 357 177 
<< pdiffusion >>
rect 357 176 358 177 
<< pdiffusion >>
rect 358 176 359 177 
<< pdiffusion >>
rect 359 176 360 177 
<< pdiffusion >>
rect 372 176 373 177 
<< pdiffusion >>
rect 373 176 374 177 
<< pdiffusion >>
rect 374 176 375 177 
<< pdiffusion >>
rect 375 176 376 177 
<< pdiffusion >>
rect 376 176 377 177 
<< pdiffusion >>
rect 377 176 378 177 
<< pdiffusion >>
rect 390 176 391 177 
<< pdiffusion >>
rect 391 176 392 177 
<< pdiffusion >>
rect 392 176 393 177 
<< pdiffusion >>
rect 393 176 394 177 
<< pdiffusion >>
rect 394 176 395 177 
<< pdiffusion >>
rect 395 176 396 177 
<< pdiffusion >>
rect 408 176 409 177 
<< pdiffusion >>
rect 409 176 410 177 
<< pdiffusion >>
rect 410 176 411 177 
<< pdiffusion >>
rect 411 176 412 177 
<< pdiffusion >>
rect 412 176 413 177 
<< pdiffusion >>
rect 413 176 414 177 
<< pdiffusion >>
rect 426 176 427 177 
<< pdiffusion >>
rect 427 176 428 177 
<< pdiffusion >>
rect 428 176 429 177 
<< pdiffusion >>
rect 429 176 430 177 
<< pdiffusion >>
rect 430 176 431 177 
<< pdiffusion >>
rect 431 176 432 177 
<< pdiffusion >>
rect 12 177 13 178 
<< pdiffusion >>
rect 13 177 14 178 
<< pdiffusion >>
rect 14 177 15 178 
<< pdiffusion >>
rect 15 177 16 178 
<< pdiffusion >>
rect 16 177 17 178 
<< pdiffusion >>
rect 17 177 18 178 
<< m1 >>
rect 19 177 20 178 
<< pdiffusion >>
rect 30 177 31 178 
<< pdiffusion >>
rect 31 177 32 178 
<< pdiffusion >>
rect 32 177 33 178 
<< pdiffusion >>
rect 33 177 34 178 
<< pdiffusion >>
rect 34 177 35 178 
<< pdiffusion >>
rect 35 177 36 178 
<< pdiffusion >>
rect 48 177 49 178 
<< pdiffusion >>
rect 49 177 50 178 
<< pdiffusion >>
rect 50 177 51 178 
<< pdiffusion >>
rect 51 177 52 178 
<< pdiffusion >>
rect 52 177 53 178 
<< pdiffusion >>
rect 53 177 54 178 
<< m1 >>
rect 64 177 65 178 
<< pdiffusion >>
rect 66 177 67 178 
<< pdiffusion >>
rect 67 177 68 178 
<< pdiffusion >>
rect 68 177 69 178 
<< pdiffusion >>
rect 69 177 70 178 
<< pdiffusion >>
rect 70 177 71 178 
<< pdiffusion >>
rect 71 177 72 178 
<< m1 >>
rect 82 177 83 178 
<< pdiffusion >>
rect 84 177 85 178 
<< pdiffusion >>
rect 85 177 86 178 
<< pdiffusion >>
rect 86 177 87 178 
<< pdiffusion >>
rect 87 177 88 178 
<< pdiffusion >>
rect 88 177 89 178 
<< pdiffusion >>
rect 89 177 90 178 
<< m1 >>
rect 93 177 94 178 
<< m1 >>
rect 100 177 101 178 
<< pdiffusion >>
rect 102 177 103 178 
<< pdiffusion >>
rect 103 177 104 178 
<< pdiffusion >>
rect 104 177 105 178 
<< pdiffusion >>
rect 105 177 106 178 
<< pdiffusion >>
rect 106 177 107 178 
<< pdiffusion >>
rect 107 177 108 178 
<< m1 >>
rect 118 177 119 178 
<< pdiffusion >>
rect 120 177 121 178 
<< pdiffusion >>
rect 121 177 122 178 
<< pdiffusion >>
rect 122 177 123 178 
<< pdiffusion >>
rect 123 177 124 178 
<< pdiffusion >>
rect 124 177 125 178 
<< pdiffusion >>
rect 125 177 126 178 
<< m1 >>
rect 127 177 128 178 
<< pdiffusion >>
rect 138 177 139 178 
<< pdiffusion >>
rect 139 177 140 178 
<< pdiffusion >>
rect 140 177 141 178 
<< pdiffusion >>
rect 141 177 142 178 
<< pdiffusion >>
rect 142 177 143 178 
<< pdiffusion >>
rect 143 177 144 178 
<< pdiffusion >>
rect 156 177 157 178 
<< pdiffusion >>
rect 157 177 158 178 
<< pdiffusion >>
rect 158 177 159 178 
<< pdiffusion >>
rect 159 177 160 178 
<< pdiffusion >>
rect 160 177 161 178 
<< pdiffusion >>
rect 161 177 162 178 
<< m1 >>
rect 170 177 171 178 
<< m1 >>
rect 172 177 173 178 
<< pdiffusion >>
rect 174 177 175 178 
<< pdiffusion >>
rect 175 177 176 178 
<< pdiffusion >>
rect 176 177 177 178 
<< pdiffusion >>
rect 177 177 178 178 
<< pdiffusion >>
rect 178 177 179 178 
<< pdiffusion >>
rect 179 177 180 178 
<< m1 >>
rect 181 177 182 178 
<< pdiffusion >>
rect 192 177 193 178 
<< pdiffusion >>
rect 193 177 194 178 
<< pdiffusion >>
rect 194 177 195 178 
<< pdiffusion >>
rect 195 177 196 178 
<< pdiffusion >>
rect 196 177 197 178 
<< pdiffusion >>
rect 197 177 198 178 
<< pdiffusion >>
rect 210 177 211 178 
<< pdiffusion >>
rect 211 177 212 178 
<< pdiffusion >>
rect 212 177 213 178 
<< pdiffusion >>
rect 213 177 214 178 
<< pdiffusion >>
rect 214 177 215 178 
<< pdiffusion >>
rect 215 177 216 178 
<< m1 >>
rect 226 177 227 178 
<< pdiffusion >>
rect 228 177 229 178 
<< pdiffusion >>
rect 229 177 230 178 
<< pdiffusion >>
rect 230 177 231 178 
<< pdiffusion >>
rect 231 177 232 178 
<< pdiffusion >>
rect 232 177 233 178 
<< pdiffusion >>
rect 233 177 234 178 
<< m1 >>
rect 235 177 236 178 
<< pdiffusion >>
rect 246 177 247 178 
<< pdiffusion >>
rect 247 177 248 178 
<< pdiffusion >>
rect 248 177 249 178 
<< pdiffusion >>
rect 249 177 250 178 
<< pdiffusion >>
rect 250 177 251 178 
<< pdiffusion >>
rect 251 177 252 178 
<< pdiffusion >>
rect 264 177 265 178 
<< pdiffusion >>
rect 265 177 266 178 
<< pdiffusion >>
rect 266 177 267 178 
<< pdiffusion >>
rect 267 177 268 178 
<< pdiffusion >>
rect 268 177 269 178 
<< pdiffusion >>
rect 269 177 270 178 
<< m1 >>
rect 271 177 272 178 
<< pdiffusion >>
rect 282 177 283 178 
<< pdiffusion >>
rect 283 177 284 178 
<< pdiffusion >>
rect 284 177 285 178 
<< pdiffusion >>
rect 285 177 286 178 
<< pdiffusion >>
rect 286 177 287 178 
<< pdiffusion >>
rect 287 177 288 178 
<< m2 >>
rect 297 177 298 178 
<< m1 >>
rect 298 177 299 178 
<< pdiffusion >>
rect 300 177 301 178 
<< pdiffusion >>
rect 301 177 302 178 
<< pdiffusion >>
rect 302 177 303 178 
<< pdiffusion >>
rect 303 177 304 178 
<< pdiffusion >>
rect 304 177 305 178 
<< pdiffusion >>
rect 305 177 306 178 
<< m1 >>
rect 307 177 308 178 
<< m1 >>
rect 311 177 312 178 
<< pdiffusion >>
rect 336 177 337 178 
<< pdiffusion >>
rect 337 177 338 178 
<< pdiffusion >>
rect 338 177 339 178 
<< pdiffusion >>
rect 339 177 340 178 
<< pdiffusion >>
rect 340 177 341 178 
<< pdiffusion >>
rect 341 177 342 178 
<< m1 >>
rect 343 177 344 178 
<< m1 >>
rect 347 177 348 178 
<< pdiffusion >>
rect 354 177 355 178 
<< pdiffusion >>
rect 355 177 356 178 
<< pdiffusion >>
rect 356 177 357 178 
<< pdiffusion >>
rect 357 177 358 178 
<< pdiffusion >>
rect 358 177 359 178 
<< pdiffusion >>
rect 359 177 360 178 
<< pdiffusion >>
rect 372 177 373 178 
<< pdiffusion >>
rect 373 177 374 178 
<< pdiffusion >>
rect 374 177 375 178 
<< pdiffusion >>
rect 375 177 376 178 
<< pdiffusion >>
rect 376 177 377 178 
<< pdiffusion >>
rect 377 177 378 178 
<< pdiffusion >>
rect 390 177 391 178 
<< pdiffusion >>
rect 391 177 392 178 
<< pdiffusion >>
rect 392 177 393 178 
<< pdiffusion >>
rect 393 177 394 178 
<< pdiffusion >>
rect 394 177 395 178 
<< pdiffusion >>
rect 395 177 396 178 
<< pdiffusion >>
rect 408 177 409 178 
<< pdiffusion >>
rect 409 177 410 178 
<< pdiffusion >>
rect 410 177 411 178 
<< pdiffusion >>
rect 411 177 412 178 
<< pdiffusion >>
rect 412 177 413 178 
<< pdiffusion >>
rect 413 177 414 178 
<< pdiffusion >>
rect 426 177 427 178 
<< pdiffusion >>
rect 427 177 428 178 
<< pdiffusion >>
rect 428 177 429 178 
<< pdiffusion >>
rect 429 177 430 178 
<< pdiffusion >>
rect 430 177 431 178 
<< pdiffusion >>
rect 431 177 432 178 
<< pdiffusion >>
rect 12 178 13 179 
<< pdiffusion >>
rect 13 178 14 179 
<< pdiffusion >>
rect 14 178 15 179 
<< pdiffusion >>
rect 15 178 16 179 
<< pdiffusion >>
rect 16 178 17 179 
<< pdiffusion >>
rect 17 178 18 179 
<< m1 >>
rect 19 178 20 179 
<< pdiffusion >>
rect 30 178 31 179 
<< pdiffusion >>
rect 31 178 32 179 
<< pdiffusion >>
rect 32 178 33 179 
<< pdiffusion >>
rect 33 178 34 179 
<< pdiffusion >>
rect 34 178 35 179 
<< pdiffusion >>
rect 35 178 36 179 
<< pdiffusion >>
rect 48 178 49 179 
<< pdiffusion >>
rect 49 178 50 179 
<< pdiffusion >>
rect 50 178 51 179 
<< pdiffusion >>
rect 51 178 52 179 
<< pdiffusion >>
rect 52 178 53 179 
<< pdiffusion >>
rect 53 178 54 179 
<< m1 >>
rect 64 178 65 179 
<< pdiffusion >>
rect 66 178 67 179 
<< pdiffusion >>
rect 67 178 68 179 
<< pdiffusion >>
rect 68 178 69 179 
<< pdiffusion >>
rect 69 178 70 179 
<< pdiffusion >>
rect 70 178 71 179 
<< pdiffusion >>
rect 71 178 72 179 
<< m1 >>
rect 82 178 83 179 
<< pdiffusion >>
rect 84 178 85 179 
<< pdiffusion >>
rect 85 178 86 179 
<< pdiffusion >>
rect 86 178 87 179 
<< pdiffusion >>
rect 87 178 88 179 
<< pdiffusion >>
rect 88 178 89 179 
<< pdiffusion >>
rect 89 178 90 179 
<< m1 >>
rect 93 178 94 179 
<< m1 >>
rect 100 178 101 179 
<< pdiffusion >>
rect 102 178 103 179 
<< pdiffusion >>
rect 103 178 104 179 
<< pdiffusion >>
rect 104 178 105 179 
<< pdiffusion >>
rect 105 178 106 179 
<< pdiffusion >>
rect 106 178 107 179 
<< pdiffusion >>
rect 107 178 108 179 
<< m1 >>
rect 118 178 119 179 
<< pdiffusion >>
rect 120 178 121 179 
<< pdiffusion >>
rect 121 178 122 179 
<< pdiffusion >>
rect 122 178 123 179 
<< pdiffusion >>
rect 123 178 124 179 
<< pdiffusion >>
rect 124 178 125 179 
<< pdiffusion >>
rect 125 178 126 179 
<< m1 >>
rect 127 178 128 179 
<< pdiffusion >>
rect 138 178 139 179 
<< pdiffusion >>
rect 139 178 140 179 
<< pdiffusion >>
rect 140 178 141 179 
<< pdiffusion >>
rect 141 178 142 179 
<< pdiffusion >>
rect 142 178 143 179 
<< pdiffusion >>
rect 143 178 144 179 
<< pdiffusion >>
rect 156 178 157 179 
<< pdiffusion >>
rect 157 178 158 179 
<< pdiffusion >>
rect 158 178 159 179 
<< pdiffusion >>
rect 159 178 160 179 
<< pdiffusion >>
rect 160 178 161 179 
<< pdiffusion >>
rect 161 178 162 179 
<< m1 >>
rect 170 178 171 179 
<< m1 >>
rect 172 178 173 179 
<< pdiffusion >>
rect 174 178 175 179 
<< pdiffusion >>
rect 175 178 176 179 
<< pdiffusion >>
rect 176 178 177 179 
<< pdiffusion >>
rect 177 178 178 179 
<< pdiffusion >>
rect 178 178 179 179 
<< pdiffusion >>
rect 179 178 180 179 
<< m1 >>
rect 181 178 182 179 
<< pdiffusion >>
rect 192 178 193 179 
<< pdiffusion >>
rect 193 178 194 179 
<< pdiffusion >>
rect 194 178 195 179 
<< pdiffusion >>
rect 195 178 196 179 
<< pdiffusion >>
rect 196 178 197 179 
<< pdiffusion >>
rect 197 178 198 179 
<< pdiffusion >>
rect 210 178 211 179 
<< pdiffusion >>
rect 211 178 212 179 
<< pdiffusion >>
rect 212 178 213 179 
<< pdiffusion >>
rect 213 178 214 179 
<< pdiffusion >>
rect 214 178 215 179 
<< pdiffusion >>
rect 215 178 216 179 
<< m1 >>
rect 226 178 227 179 
<< pdiffusion >>
rect 228 178 229 179 
<< pdiffusion >>
rect 229 178 230 179 
<< pdiffusion >>
rect 230 178 231 179 
<< pdiffusion >>
rect 231 178 232 179 
<< pdiffusion >>
rect 232 178 233 179 
<< pdiffusion >>
rect 233 178 234 179 
<< m1 >>
rect 235 178 236 179 
<< pdiffusion >>
rect 246 178 247 179 
<< pdiffusion >>
rect 247 178 248 179 
<< pdiffusion >>
rect 248 178 249 179 
<< pdiffusion >>
rect 249 178 250 179 
<< pdiffusion >>
rect 250 178 251 179 
<< pdiffusion >>
rect 251 178 252 179 
<< pdiffusion >>
rect 264 178 265 179 
<< pdiffusion >>
rect 265 178 266 179 
<< pdiffusion >>
rect 266 178 267 179 
<< pdiffusion >>
rect 267 178 268 179 
<< pdiffusion >>
rect 268 178 269 179 
<< pdiffusion >>
rect 269 178 270 179 
<< m1 >>
rect 271 178 272 179 
<< pdiffusion >>
rect 282 178 283 179 
<< pdiffusion >>
rect 283 178 284 179 
<< pdiffusion >>
rect 284 178 285 179 
<< pdiffusion >>
rect 285 178 286 179 
<< pdiffusion >>
rect 286 178 287 179 
<< pdiffusion >>
rect 287 178 288 179 
<< m2 >>
rect 297 178 298 179 
<< m1 >>
rect 298 178 299 179 
<< pdiffusion >>
rect 300 178 301 179 
<< pdiffusion >>
rect 301 178 302 179 
<< pdiffusion >>
rect 302 178 303 179 
<< pdiffusion >>
rect 303 178 304 179 
<< pdiffusion >>
rect 304 178 305 179 
<< pdiffusion >>
rect 305 178 306 179 
<< m1 >>
rect 307 178 308 179 
<< m1 >>
rect 311 178 312 179 
<< pdiffusion >>
rect 336 178 337 179 
<< pdiffusion >>
rect 337 178 338 179 
<< pdiffusion >>
rect 338 178 339 179 
<< pdiffusion >>
rect 339 178 340 179 
<< pdiffusion >>
rect 340 178 341 179 
<< pdiffusion >>
rect 341 178 342 179 
<< m1 >>
rect 343 178 344 179 
<< m1 >>
rect 347 178 348 179 
<< pdiffusion >>
rect 354 178 355 179 
<< pdiffusion >>
rect 355 178 356 179 
<< pdiffusion >>
rect 356 178 357 179 
<< pdiffusion >>
rect 357 178 358 179 
<< pdiffusion >>
rect 358 178 359 179 
<< pdiffusion >>
rect 359 178 360 179 
<< pdiffusion >>
rect 372 178 373 179 
<< pdiffusion >>
rect 373 178 374 179 
<< pdiffusion >>
rect 374 178 375 179 
<< pdiffusion >>
rect 375 178 376 179 
<< pdiffusion >>
rect 376 178 377 179 
<< pdiffusion >>
rect 377 178 378 179 
<< pdiffusion >>
rect 390 178 391 179 
<< pdiffusion >>
rect 391 178 392 179 
<< pdiffusion >>
rect 392 178 393 179 
<< pdiffusion >>
rect 393 178 394 179 
<< pdiffusion >>
rect 394 178 395 179 
<< pdiffusion >>
rect 395 178 396 179 
<< pdiffusion >>
rect 408 178 409 179 
<< pdiffusion >>
rect 409 178 410 179 
<< pdiffusion >>
rect 410 178 411 179 
<< pdiffusion >>
rect 411 178 412 179 
<< pdiffusion >>
rect 412 178 413 179 
<< pdiffusion >>
rect 413 178 414 179 
<< pdiffusion >>
rect 426 178 427 179 
<< pdiffusion >>
rect 427 178 428 179 
<< pdiffusion >>
rect 428 178 429 179 
<< pdiffusion >>
rect 429 178 430 179 
<< pdiffusion >>
rect 430 178 431 179 
<< pdiffusion >>
rect 431 178 432 179 
<< pdiffusion >>
rect 12 179 13 180 
<< pdiffusion >>
rect 13 179 14 180 
<< pdiffusion >>
rect 14 179 15 180 
<< pdiffusion >>
rect 15 179 16 180 
<< pdiffusion >>
rect 16 179 17 180 
<< pdiffusion >>
rect 17 179 18 180 
<< m1 >>
rect 19 179 20 180 
<< pdiffusion >>
rect 30 179 31 180 
<< pdiffusion >>
rect 31 179 32 180 
<< pdiffusion >>
rect 32 179 33 180 
<< pdiffusion >>
rect 33 179 34 180 
<< pdiffusion >>
rect 34 179 35 180 
<< pdiffusion >>
rect 35 179 36 180 
<< pdiffusion >>
rect 48 179 49 180 
<< pdiffusion >>
rect 49 179 50 180 
<< pdiffusion >>
rect 50 179 51 180 
<< pdiffusion >>
rect 51 179 52 180 
<< m1 >>
rect 52 179 53 180 
<< pdiffusion >>
rect 52 179 53 180 
<< pdiffusion >>
rect 53 179 54 180 
<< m1 >>
rect 64 179 65 180 
<< pdiffusion >>
rect 66 179 67 180 
<< pdiffusion >>
rect 67 179 68 180 
<< pdiffusion >>
rect 68 179 69 180 
<< pdiffusion >>
rect 69 179 70 180 
<< m1 >>
rect 70 179 71 180 
<< pdiffusion >>
rect 70 179 71 180 
<< pdiffusion >>
rect 71 179 72 180 
<< m1 >>
rect 82 179 83 180 
<< pdiffusion >>
rect 84 179 85 180 
<< pdiffusion >>
rect 85 179 86 180 
<< pdiffusion >>
rect 86 179 87 180 
<< pdiffusion >>
rect 87 179 88 180 
<< pdiffusion >>
rect 88 179 89 180 
<< pdiffusion >>
rect 89 179 90 180 
<< m1 >>
rect 93 179 94 180 
<< m1 >>
rect 100 179 101 180 
<< pdiffusion >>
rect 102 179 103 180 
<< m1 >>
rect 103 179 104 180 
<< pdiffusion >>
rect 103 179 104 180 
<< pdiffusion >>
rect 104 179 105 180 
<< pdiffusion >>
rect 105 179 106 180 
<< pdiffusion >>
rect 106 179 107 180 
<< pdiffusion >>
rect 107 179 108 180 
<< m1 >>
rect 118 179 119 180 
<< pdiffusion >>
rect 120 179 121 180 
<< pdiffusion >>
rect 121 179 122 180 
<< pdiffusion >>
rect 122 179 123 180 
<< pdiffusion >>
rect 123 179 124 180 
<< pdiffusion >>
rect 124 179 125 180 
<< pdiffusion >>
rect 125 179 126 180 
<< m1 >>
rect 127 179 128 180 
<< pdiffusion >>
rect 138 179 139 180 
<< pdiffusion >>
rect 139 179 140 180 
<< pdiffusion >>
rect 140 179 141 180 
<< pdiffusion >>
rect 141 179 142 180 
<< pdiffusion >>
rect 142 179 143 180 
<< pdiffusion >>
rect 143 179 144 180 
<< pdiffusion >>
rect 156 179 157 180 
<< pdiffusion >>
rect 157 179 158 180 
<< pdiffusion >>
rect 158 179 159 180 
<< pdiffusion >>
rect 159 179 160 180 
<< pdiffusion >>
rect 160 179 161 180 
<< pdiffusion >>
rect 161 179 162 180 
<< m1 >>
rect 170 179 171 180 
<< m1 >>
rect 172 179 173 180 
<< pdiffusion >>
rect 174 179 175 180 
<< pdiffusion >>
rect 175 179 176 180 
<< pdiffusion >>
rect 176 179 177 180 
<< pdiffusion >>
rect 177 179 178 180 
<< pdiffusion >>
rect 178 179 179 180 
<< pdiffusion >>
rect 179 179 180 180 
<< m1 >>
rect 181 179 182 180 
<< pdiffusion >>
rect 192 179 193 180 
<< pdiffusion >>
rect 193 179 194 180 
<< pdiffusion >>
rect 194 179 195 180 
<< pdiffusion >>
rect 195 179 196 180 
<< m1 >>
rect 196 179 197 180 
<< pdiffusion >>
rect 196 179 197 180 
<< pdiffusion >>
rect 197 179 198 180 
<< pdiffusion >>
rect 210 179 211 180 
<< m1 >>
rect 211 179 212 180 
<< pdiffusion >>
rect 211 179 212 180 
<< pdiffusion >>
rect 212 179 213 180 
<< pdiffusion >>
rect 213 179 214 180 
<< pdiffusion >>
rect 214 179 215 180 
<< pdiffusion >>
rect 215 179 216 180 
<< m1 >>
rect 226 179 227 180 
<< pdiffusion >>
rect 228 179 229 180 
<< m1 >>
rect 229 179 230 180 
<< pdiffusion >>
rect 229 179 230 180 
<< pdiffusion >>
rect 230 179 231 180 
<< pdiffusion >>
rect 231 179 232 180 
<< pdiffusion >>
rect 232 179 233 180 
<< pdiffusion >>
rect 233 179 234 180 
<< m1 >>
rect 235 179 236 180 
<< pdiffusion >>
rect 246 179 247 180 
<< pdiffusion >>
rect 247 179 248 180 
<< pdiffusion >>
rect 248 179 249 180 
<< pdiffusion >>
rect 249 179 250 180 
<< pdiffusion >>
rect 250 179 251 180 
<< pdiffusion >>
rect 251 179 252 180 
<< pdiffusion >>
rect 264 179 265 180 
<< pdiffusion >>
rect 265 179 266 180 
<< pdiffusion >>
rect 266 179 267 180 
<< pdiffusion >>
rect 267 179 268 180 
<< m1 >>
rect 268 179 269 180 
<< pdiffusion >>
rect 268 179 269 180 
<< pdiffusion >>
rect 269 179 270 180 
<< m1 >>
rect 271 179 272 180 
<< pdiffusion >>
rect 282 179 283 180 
<< pdiffusion >>
rect 283 179 284 180 
<< pdiffusion >>
rect 284 179 285 180 
<< pdiffusion >>
rect 285 179 286 180 
<< pdiffusion >>
rect 286 179 287 180 
<< pdiffusion >>
rect 287 179 288 180 
<< m2 >>
rect 297 179 298 180 
<< m1 >>
rect 298 179 299 180 
<< pdiffusion >>
rect 300 179 301 180 
<< m1 >>
rect 301 179 302 180 
<< pdiffusion >>
rect 301 179 302 180 
<< pdiffusion >>
rect 302 179 303 180 
<< pdiffusion >>
rect 303 179 304 180 
<< pdiffusion >>
rect 304 179 305 180 
<< pdiffusion >>
rect 305 179 306 180 
<< m1 >>
rect 307 179 308 180 
<< m1 >>
rect 311 179 312 180 
<< pdiffusion >>
rect 336 179 337 180 
<< m1 >>
rect 337 179 338 180 
<< pdiffusion >>
rect 337 179 338 180 
<< pdiffusion >>
rect 338 179 339 180 
<< pdiffusion >>
rect 339 179 340 180 
<< pdiffusion >>
rect 340 179 341 180 
<< pdiffusion >>
rect 341 179 342 180 
<< m1 >>
rect 343 179 344 180 
<< m1 >>
rect 347 179 348 180 
<< pdiffusion >>
rect 354 179 355 180 
<< pdiffusion >>
rect 355 179 356 180 
<< pdiffusion >>
rect 356 179 357 180 
<< pdiffusion >>
rect 357 179 358 180 
<< m1 >>
rect 358 179 359 180 
<< pdiffusion >>
rect 358 179 359 180 
<< pdiffusion >>
rect 359 179 360 180 
<< pdiffusion >>
rect 372 179 373 180 
<< pdiffusion >>
rect 373 179 374 180 
<< pdiffusion >>
rect 374 179 375 180 
<< pdiffusion >>
rect 375 179 376 180 
<< pdiffusion >>
rect 376 179 377 180 
<< pdiffusion >>
rect 377 179 378 180 
<< pdiffusion >>
rect 390 179 391 180 
<< pdiffusion >>
rect 391 179 392 180 
<< pdiffusion >>
rect 392 179 393 180 
<< pdiffusion >>
rect 393 179 394 180 
<< pdiffusion >>
rect 394 179 395 180 
<< pdiffusion >>
rect 395 179 396 180 
<< pdiffusion >>
rect 408 179 409 180 
<< pdiffusion >>
rect 409 179 410 180 
<< pdiffusion >>
rect 410 179 411 180 
<< pdiffusion >>
rect 411 179 412 180 
<< pdiffusion >>
rect 412 179 413 180 
<< pdiffusion >>
rect 413 179 414 180 
<< pdiffusion >>
rect 426 179 427 180 
<< pdiffusion >>
rect 427 179 428 180 
<< pdiffusion >>
rect 428 179 429 180 
<< pdiffusion >>
rect 429 179 430 180 
<< pdiffusion >>
rect 430 179 431 180 
<< pdiffusion >>
rect 431 179 432 180 
<< m1 >>
rect 19 180 20 181 
<< m1 >>
rect 52 180 53 181 
<< m1 >>
rect 64 180 65 181 
<< m1 >>
rect 70 180 71 181 
<< m1 >>
rect 82 180 83 181 
<< m1 >>
rect 93 180 94 181 
<< m1 >>
rect 100 180 101 181 
<< m1 >>
rect 103 180 104 181 
<< m1 >>
rect 118 180 119 181 
<< m1 >>
rect 127 180 128 181 
<< m1 >>
rect 170 180 171 181 
<< m1 >>
rect 172 180 173 181 
<< m1 >>
rect 181 180 182 181 
<< m1 >>
rect 196 180 197 181 
<< m1 >>
rect 211 180 212 181 
<< m1 >>
rect 226 180 227 181 
<< m1 >>
rect 229 180 230 181 
<< m1 >>
rect 235 180 236 181 
<< m1 >>
rect 268 180 269 181 
<< m1 >>
rect 271 180 272 181 
<< m2 >>
rect 297 180 298 181 
<< m1 >>
rect 298 180 299 181 
<< m1 >>
rect 301 180 302 181 
<< m1 >>
rect 307 180 308 181 
<< m1 >>
rect 311 180 312 181 
<< m1 >>
rect 337 180 338 181 
<< m1 >>
rect 343 180 344 181 
<< m1 >>
rect 347 180 348 181 
<< m1 >>
rect 358 180 359 181 
<< m1 >>
rect 19 181 20 182 
<< m1 >>
rect 52 181 53 182 
<< m1 >>
rect 53 181 54 182 
<< m1 >>
rect 54 181 55 182 
<< m1 >>
rect 55 181 56 182 
<< m1 >>
rect 56 181 57 182 
<< m1 >>
rect 57 181 58 182 
<< m1 >>
rect 58 181 59 182 
<< m1 >>
rect 59 181 60 182 
<< m1 >>
rect 60 181 61 182 
<< m1 >>
rect 61 181 62 182 
<< m1 >>
rect 62 181 63 182 
<< m1 >>
rect 63 181 64 182 
<< m1 >>
rect 64 181 65 182 
<< m1 >>
rect 70 181 71 182 
<< m1 >>
rect 71 181 72 182 
<< m1 >>
rect 72 181 73 182 
<< m1 >>
rect 73 181 74 182 
<< m1 >>
rect 74 181 75 182 
<< m1 >>
rect 75 181 76 182 
<< m1 >>
rect 76 181 77 182 
<< m1 >>
rect 77 181 78 182 
<< m1 >>
rect 78 181 79 182 
<< m1 >>
rect 79 181 80 182 
<< m1 >>
rect 80 181 81 182 
<< m1 >>
rect 81 181 82 182 
<< m1 >>
rect 82 181 83 182 
<< m1 >>
rect 93 181 94 182 
<< m1 >>
rect 100 181 101 182 
<< m1 >>
rect 101 181 102 182 
<< m1 >>
rect 102 181 103 182 
<< m1 >>
rect 103 181 104 182 
<< m1 >>
rect 118 181 119 182 
<< m1 >>
rect 127 181 128 182 
<< m1 >>
rect 170 181 171 182 
<< m1 >>
rect 172 181 173 182 
<< m1 >>
rect 181 181 182 182 
<< m1 >>
rect 196 181 197 182 
<< m1 >>
rect 197 181 198 182 
<< m1 >>
rect 198 181 199 182 
<< m1 >>
rect 199 181 200 182 
<< m1 >>
rect 200 181 201 182 
<< m1 >>
rect 201 181 202 182 
<< m1 >>
rect 202 181 203 182 
<< m1 >>
rect 203 181 204 182 
<< m1 >>
rect 204 181 205 182 
<< m1 >>
rect 205 181 206 182 
<< m1 >>
rect 206 181 207 182 
<< m1 >>
rect 207 181 208 182 
<< m1 >>
rect 208 181 209 182 
<< m1 >>
rect 209 181 210 182 
<< m1 >>
rect 210 181 211 182 
<< m1 >>
rect 211 181 212 182 
<< m1 >>
rect 226 181 227 182 
<< m1 >>
rect 229 181 230 182 
<< m1 >>
rect 235 181 236 182 
<< m1 >>
rect 268 181 269 182 
<< m1 >>
rect 269 181 270 182 
<< m1 >>
rect 270 181 271 182 
<< m1 >>
rect 271 181 272 182 
<< m2 >>
rect 297 181 298 182 
<< m1 >>
rect 298 181 299 182 
<< m2 >>
rect 298 181 299 182 
<< m2 >>
rect 299 181 300 182 
<< m1 >>
rect 300 181 301 182 
<< m2 >>
rect 300 181 301 182 
<< m2c >>
rect 300 181 301 182 
<< m1 >>
rect 300 181 301 182 
<< m2 >>
rect 300 181 301 182 
<< m1 >>
rect 301 181 302 182 
<< m1 >>
rect 307 181 308 182 
<< m1 >>
rect 311 181 312 182 
<< m1 >>
rect 337 181 338 182 
<< m1 >>
rect 343 181 344 182 
<< m1 >>
rect 347 181 348 182 
<< m1 >>
rect 358 181 359 182 
<< m1 >>
rect 19 182 20 183 
<< m1 >>
rect 93 182 94 183 
<< m1 >>
rect 118 182 119 183 
<< m1 >>
rect 127 182 128 183 
<< m2 >>
rect 127 182 128 183 
<< m2c >>
rect 127 182 128 183 
<< m1 >>
rect 127 182 128 183 
<< m2 >>
rect 127 182 128 183 
<< m1 >>
rect 170 182 171 183 
<< m1 >>
rect 172 182 173 183 
<< m1 >>
rect 181 182 182 183 
<< m1 >>
rect 226 182 227 183 
<< m1 >>
rect 229 182 230 183 
<< m1 >>
rect 235 182 236 183 
<< m2 >>
rect 235 182 236 183 
<< m2c >>
rect 235 182 236 183 
<< m1 >>
rect 235 182 236 183 
<< m2 >>
rect 235 182 236 183 
<< m1 >>
rect 298 182 299 183 
<< m1 >>
rect 307 182 308 183 
<< m1 >>
rect 311 182 312 183 
<< m1 >>
rect 337 182 338 183 
<< m1 >>
rect 338 182 339 183 
<< m1 >>
rect 339 182 340 183 
<< m1 >>
rect 340 182 341 183 
<< m1 >>
rect 341 182 342 183 
<< m2 >>
rect 341 182 342 183 
<< m2c >>
rect 341 182 342 183 
<< m1 >>
rect 341 182 342 183 
<< m2 >>
rect 341 182 342 183 
<< m2 >>
rect 342 182 343 183 
<< m1 >>
rect 343 182 344 183 
<< m2 >>
rect 343 182 344 183 
<< m2 >>
rect 344 182 345 183 
<< m1 >>
rect 345 182 346 183 
<< m2 >>
rect 345 182 346 183 
<< m2c >>
rect 345 182 346 183 
<< m1 >>
rect 345 182 346 183 
<< m2 >>
rect 345 182 346 183 
<< m1 >>
rect 347 182 348 183 
<< m1 >>
rect 358 182 359 183 
<< m1 >>
rect 19 183 20 184 
<< m1 >>
rect 93 183 94 184 
<< m1 >>
rect 118 183 119 184 
<< m2 >>
rect 127 183 128 184 
<< m1 >>
rect 170 183 171 184 
<< m1 >>
rect 172 183 173 184 
<< m1 >>
rect 181 183 182 184 
<< m1 >>
rect 226 183 227 184 
<< m1 >>
rect 229 183 230 184 
<< m2 >>
rect 235 183 236 184 
<< m1 >>
rect 298 183 299 184 
<< m1 >>
rect 307 183 308 184 
<< m1 >>
rect 311 183 312 184 
<< m1 >>
rect 343 183 344 184 
<< m1 >>
rect 345 183 346 184 
<< m1 >>
rect 347 183 348 184 
<< m1 >>
rect 358 183 359 184 
<< m1 >>
rect 19 184 20 185 
<< m1 >>
rect 93 184 94 185 
<< m1 >>
rect 118 184 119 185 
<< m1 >>
rect 121 184 122 185 
<< m1 >>
rect 122 184 123 185 
<< m1 >>
rect 123 184 124 185 
<< m1 >>
rect 124 184 125 185 
<< m1 >>
rect 125 184 126 185 
<< m1 >>
rect 126 184 127 185 
<< m1 >>
rect 127 184 128 185 
<< m2 >>
rect 127 184 128 185 
<< m1 >>
rect 128 184 129 185 
<< m1 >>
rect 129 184 130 185 
<< m1 >>
rect 130 184 131 185 
<< m1 >>
rect 131 184 132 185 
<< m1 >>
rect 132 184 133 185 
<< m1 >>
rect 133 184 134 185 
<< m1 >>
rect 134 184 135 185 
<< m1 >>
rect 135 184 136 185 
<< m1 >>
rect 136 184 137 185 
<< m1 >>
rect 137 184 138 185 
<< m1 >>
rect 138 184 139 185 
<< m1 >>
rect 139 184 140 185 
<< m1 >>
rect 140 184 141 185 
<< m1 >>
rect 141 184 142 185 
<< m1 >>
rect 142 184 143 185 
<< m1 >>
rect 143 184 144 185 
<< m1 >>
rect 144 184 145 185 
<< m1 >>
rect 145 184 146 185 
<< m1 >>
rect 146 184 147 185 
<< m1 >>
rect 147 184 148 185 
<< m1 >>
rect 148 184 149 185 
<< m1 >>
rect 149 184 150 185 
<< m1 >>
rect 150 184 151 185 
<< m1 >>
rect 151 184 152 185 
<< m1 >>
rect 152 184 153 185 
<< m1 >>
rect 153 184 154 185 
<< m1 >>
rect 154 184 155 185 
<< m1 >>
rect 155 184 156 185 
<< m1 >>
rect 156 184 157 185 
<< m1 >>
rect 157 184 158 185 
<< m1 >>
rect 158 184 159 185 
<< m1 >>
rect 159 184 160 185 
<< m1 >>
rect 160 184 161 185 
<< m1 >>
rect 161 184 162 185 
<< m1 >>
rect 162 184 163 185 
<< m1 >>
rect 163 184 164 185 
<< m1 >>
rect 164 184 165 185 
<< m1 >>
rect 165 184 166 185 
<< m1 >>
rect 166 184 167 185 
<< m1 >>
rect 167 184 168 185 
<< m1 >>
rect 168 184 169 185 
<< m1 >>
rect 169 184 170 185 
<< m1 >>
rect 170 184 171 185 
<< m1 >>
rect 172 184 173 185 
<< m1 >>
rect 181 184 182 185 
<< m1 >>
rect 226 184 227 185 
<< m1 >>
rect 229 184 230 185 
<< m1 >>
rect 230 184 231 185 
<< m1 >>
rect 231 184 232 185 
<< m1 >>
rect 232 184 233 185 
<< m1 >>
rect 233 184 234 185 
<< m1 >>
rect 234 184 235 185 
<< m1 >>
rect 235 184 236 185 
<< m2 >>
rect 235 184 236 185 
<< m1 >>
rect 236 184 237 185 
<< m1 >>
rect 237 184 238 185 
<< m1 >>
rect 238 184 239 185 
<< m1 >>
rect 239 184 240 185 
<< m1 >>
rect 240 184 241 185 
<< m1 >>
rect 241 184 242 185 
<< m1 >>
rect 242 184 243 185 
<< m1 >>
rect 243 184 244 185 
<< m1 >>
rect 244 184 245 185 
<< m1 >>
rect 245 184 246 185 
<< m1 >>
rect 246 184 247 185 
<< m1 >>
rect 247 184 248 185 
<< m1 >>
rect 298 184 299 185 
<< m1 >>
rect 307 184 308 185 
<< m1 >>
rect 311 184 312 185 
<< m1 >>
rect 343 184 344 185 
<< m1 >>
rect 345 184 346 185 
<< m1 >>
rect 347 184 348 185 
<< m1 >>
rect 348 184 349 185 
<< m1 >>
rect 349 184 350 185 
<< m1 >>
rect 350 184 351 185 
<< m1 >>
rect 351 184 352 185 
<< m1 >>
rect 352 184 353 185 
<< m1 >>
rect 353 184 354 185 
<< m1 >>
rect 354 184 355 185 
<< m1 >>
rect 355 184 356 185 
<< m1 >>
rect 356 184 357 185 
<< m1 >>
rect 357 184 358 185 
<< m1 >>
rect 358 184 359 185 
<< m1 >>
rect 19 185 20 186 
<< m1 >>
rect 93 185 94 186 
<< m1 >>
rect 118 185 119 186 
<< m1 >>
rect 121 185 122 186 
<< m2 >>
rect 127 185 128 186 
<< m1 >>
rect 172 185 173 186 
<< m1 >>
rect 181 185 182 186 
<< m1 >>
rect 226 185 227 186 
<< m2 >>
rect 235 185 236 186 
<< m1 >>
rect 247 185 248 186 
<< m1 >>
rect 298 185 299 186 
<< m1 >>
rect 307 185 308 186 
<< m1 >>
rect 311 185 312 186 
<< m1 >>
rect 343 185 344 186 
<< m1 >>
rect 345 185 346 186 
<< m1 >>
rect 19 186 20 187 
<< m1 >>
rect 93 186 94 187 
<< m1 >>
rect 118 186 119 187 
<< m1 >>
rect 121 186 122 187 
<< m2 >>
rect 127 186 128 187 
<< m1 >>
rect 172 186 173 187 
<< m1 >>
rect 181 186 182 187 
<< m1 >>
rect 226 186 227 187 
<< m1 >>
rect 235 186 236 187 
<< m2 >>
rect 235 186 236 187 
<< m2c >>
rect 235 186 236 187 
<< m1 >>
rect 235 186 236 187 
<< m2 >>
rect 235 186 236 187 
<< m1 >>
rect 247 186 248 187 
<< m1 >>
rect 298 186 299 187 
<< m1 >>
rect 307 186 308 187 
<< m1 >>
rect 311 186 312 187 
<< m1 >>
rect 343 186 344 187 
<< m1 >>
rect 345 186 346 187 
<< m1 >>
rect 346 186 347 187 
<< m1 >>
rect 347 186 348 187 
<< m1 >>
rect 348 186 349 187 
<< m1 >>
rect 349 186 350 187 
<< m1 >>
rect 350 186 351 187 
<< m1 >>
rect 351 186 352 187 
<< m1 >>
rect 352 186 353 187 
<< m1 >>
rect 353 186 354 187 
<< m1 >>
rect 354 186 355 187 
<< m1 >>
rect 355 186 356 187 
<< m1 >>
rect 19 187 20 188 
<< m1 >>
rect 93 187 94 188 
<< m1 >>
rect 118 187 119 188 
<< m1 >>
rect 121 187 122 188 
<< m1 >>
rect 127 187 128 188 
<< m2 >>
rect 127 187 128 188 
<< m1 >>
rect 128 187 129 188 
<< m1 >>
rect 129 187 130 188 
<< m1 >>
rect 130 187 131 188 
<< m1 >>
rect 131 187 132 188 
<< m1 >>
rect 132 187 133 188 
<< m1 >>
rect 133 187 134 188 
<< m1 >>
rect 134 187 135 188 
<< m1 >>
rect 135 187 136 188 
<< m1 >>
rect 136 187 137 188 
<< m1 >>
rect 137 187 138 188 
<< m1 >>
rect 138 187 139 188 
<< m1 >>
rect 139 187 140 188 
<< m1 >>
rect 140 187 141 188 
<< m1 >>
rect 141 187 142 188 
<< m1 >>
rect 142 187 143 188 
<< m1 >>
rect 154 187 155 188 
<< m1 >>
rect 155 187 156 188 
<< m1 >>
rect 156 187 157 188 
<< m1 >>
rect 157 187 158 188 
<< m1 >>
rect 158 187 159 188 
<< m1 >>
rect 159 187 160 188 
<< m1 >>
rect 160 187 161 188 
<< m1 >>
rect 172 187 173 188 
<< m1 >>
rect 181 187 182 188 
<< m2 >>
rect 181 187 182 188 
<< m2c >>
rect 181 187 182 188 
<< m1 >>
rect 181 187 182 188 
<< m2 >>
rect 181 187 182 188 
<< m1 >>
rect 226 187 227 188 
<< m1 >>
rect 235 187 236 188 
<< m1 >>
rect 247 187 248 188 
<< m1 >>
rect 254 187 255 188 
<< m1 >>
rect 255 187 256 188 
<< m1 >>
rect 256 187 257 188 
<< m1 >>
rect 257 187 258 188 
<< m1 >>
rect 258 187 259 188 
<< m1 >>
rect 259 187 260 188 
<< m1 >>
rect 260 187 261 188 
<< m1 >>
rect 261 187 262 188 
<< m1 >>
rect 262 187 263 188 
<< m1 >>
rect 263 187 264 188 
<< m1 >>
rect 264 187 265 188 
<< m1 >>
rect 265 187 266 188 
<< m1 >>
rect 266 187 267 188 
<< m1 >>
rect 267 187 268 188 
<< m1 >>
rect 268 187 269 188 
<< m1 >>
rect 269 187 270 188 
<< m1 >>
rect 270 187 271 188 
<< m1 >>
rect 271 187 272 188 
<< m1 >>
rect 272 187 273 188 
<< m1 >>
rect 273 187 274 188 
<< m1 >>
rect 274 187 275 188 
<< m1 >>
rect 275 187 276 188 
<< m1 >>
rect 276 187 277 188 
<< m1 >>
rect 277 187 278 188 
<< m1 >>
rect 278 187 279 188 
<< m1 >>
rect 279 187 280 188 
<< m1 >>
rect 280 187 281 188 
<< m1 >>
rect 281 187 282 188 
<< m1 >>
rect 282 187 283 188 
<< m1 >>
rect 283 187 284 188 
<< m1 >>
rect 284 187 285 188 
<< m1 >>
rect 285 187 286 188 
<< m1 >>
rect 286 187 287 188 
<< m1 >>
rect 287 187 288 188 
<< m1 >>
rect 288 187 289 188 
<< m1 >>
rect 289 187 290 188 
<< m1 >>
rect 290 187 291 188 
<< m1 >>
rect 291 187 292 188 
<< m1 >>
rect 292 187 293 188 
<< m1 >>
rect 293 187 294 188 
<< m1 >>
rect 294 187 295 188 
<< m1 >>
rect 295 187 296 188 
<< m1 >>
rect 296 187 297 188 
<< m2 >>
rect 296 187 297 188 
<< m2c >>
rect 296 187 297 188 
<< m1 >>
rect 296 187 297 188 
<< m2 >>
rect 296 187 297 188 
<< m2 >>
rect 297 187 298 188 
<< m1 >>
rect 298 187 299 188 
<< m2 >>
rect 298 187 299 188 
<< m2 >>
rect 299 187 300 188 
<< m1 >>
rect 300 187 301 188 
<< m2 >>
rect 300 187 301 188 
<< m2c >>
rect 300 187 301 188 
<< m1 >>
rect 300 187 301 188 
<< m2 >>
rect 300 187 301 188 
<< m1 >>
rect 301 187 302 188 
<< m1 >>
rect 302 187 303 188 
<< m1 >>
rect 303 187 304 188 
<< m1 >>
rect 304 187 305 188 
<< m1 >>
rect 305 187 306 188 
<< m2 >>
rect 305 187 306 188 
<< m2c >>
rect 305 187 306 188 
<< m1 >>
rect 305 187 306 188 
<< m2 >>
rect 305 187 306 188 
<< m2 >>
rect 306 187 307 188 
<< m1 >>
rect 307 187 308 188 
<< m2 >>
rect 307 187 308 188 
<< m2 >>
rect 308 187 309 188 
<< m1 >>
rect 309 187 310 188 
<< m2 >>
rect 309 187 310 188 
<< m2c >>
rect 309 187 310 188 
<< m1 >>
rect 309 187 310 188 
<< m2 >>
rect 309 187 310 188 
<< m2 >>
rect 310 187 311 188 
<< m1 >>
rect 311 187 312 188 
<< m2 >>
rect 311 187 312 188 
<< m2 >>
rect 312 187 313 188 
<< m1 >>
rect 313 187 314 188 
<< m2 >>
rect 313 187 314 188 
<< m2c >>
rect 313 187 314 188 
<< m1 >>
rect 313 187 314 188 
<< m2 >>
rect 313 187 314 188 
<< m1 >>
rect 343 187 344 188 
<< m1 >>
rect 355 187 356 188 
<< m1 >>
rect 19 188 20 189 
<< m1 >>
rect 93 188 94 189 
<< m1 >>
rect 118 188 119 189 
<< m1 >>
rect 121 188 122 189 
<< m1 >>
rect 127 188 128 189 
<< m2 >>
rect 127 188 128 189 
<< m1 >>
rect 142 188 143 189 
<< m1 >>
rect 154 188 155 189 
<< m1 >>
rect 160 188 161 189 
<< m1 >>
rect 172 188 173 189 
<< m2 >>
rect 181 188 182 189 
<< m1 >>
rect 226 188 227 189 
<< m1 >>
rect 235 188 236 189 
<< m1 >>
rect 247 188 248 189 
<< m1 >>
rect 254 188 255 189 
<< m1 >>
rect 298 188 299 189 
<< m1 >>
rect 307 188 308 189 
<< m1 >>
rect 311 188 312 189 
<< m1 >>
rect 313 188 314 189 
<< m1 >>
rect 343 188 344 189 
<< m1 >>
rect 355 188 356 189 
<< m1 >>
rect 19 189 20 190 
<< m1 >>
rect 93 189 94 190 
<< m1 >>
rect 118 189 119 190 
<< m1 >>
rect 121 189 122 190 
<< m1 >>
rect 127 189 128 190 
<< m2 >>
rect 127 189 128 190 
<< m1 >>
rect 142 189 143 190 
<< m1 >>
rect 154 189 155 190 
<< m1 >>
rect 160 189 161 190 
<< m1 >>
rect 172 189 173 190 
<< m1 >>
rect 175 189 176 190 
<< m1 >>
rect 176 189 177 190 
<< m1 >>
rect 177 189 178 190 
<< m1 >>
rect 178 189 179 190 
<< m1 >>
rect 179 189 180 190 
<< m1 >>
rect 180 189 181 190 
<< m1 >>
rect 181 189 182 190 
<< m2 >>
rect 181 189 182 190 
<< m1 >>
rect 211 189 212 190 
<< m1 >>
rect 212 189 213 190 
<< m1 >>
rect 213 189 214 190 
<< m1 >>
rect 214 189 215 190 
<< m1 >>
rect 215 189 216 190 
<< m1 >>
rect 216 189 217 190 
<< m1 >>
rect 217 189 218 190 
<< m1 >>
rect 226 189 227 190 
<< m1 >>
rect 235 189 236 190 
<< m1 >>
rect 247 189 248 190 
<< m1 >>
rect 254 189 255 190 
<< m1 >>
rect 298 189 299 190 
<< m1 >>
rect 301 189 302 190 
<< m1 >>
rect 302 189 303 190 
<< m1 >>
rect 303 189 304 190 
<< m1 >>
rect 304 189 305 190 
<< m1 >>
rect 305 189 306 190 
<< m1 >>
rect 307 189 308 190 
<< m1 >>
rect 311 189 312 190 
<< m1 >>
rect 313 189 314 190 
<< m1 >>
rect 343 189 344 190 
<< m1 >>
rect 355 189 356 190 
<< m1 >>
rect 19 190 20 191 
<< m1 >>
rect 93 190 94 191 
<< m1 >>
rect 118 190 119 191 
<< m1 >>
rect 121 190 122 191 
<< m1 >>
rect 127 190 128 191 
<< m2 >>
rect 127 190 128 191 
<< m1 >>
rect 142 190 143 191 
<< m1 >>
rect 154 190 155 191 
<< m1 >>
rect 160 190 161 191 
<< m1 >>
rect 172 190 173 191 
<< m1 >>
rect 175 190 176 191 
<< m1 >>
rect 181 190 182 191 
<< m2 >>
rect 181 190 182 191 
<< m1 >>
rect 211 190 212 191 
<< m1 >>
rect 217 190 218 191 
<< m1 >>
rect 226 190 227 191 
<< m1 >>
rect 235 190 236 191 
<< m1 >>
rect 247 190 248 191 
<< m1 >>
rect 254 190 255 191 
<< m1 >>
rect 298 190 299 191 
<< m1 >>
rect 301 190 302 191 
<< m1 >>
rect 305 190 306 191 
<< m2 >>
rect 305 190 306 191 
<< m2c >>
rect 305 190 306 191 
<< m1 >>
rect 305 190 306 191 
<< m2 >>
rect 305 190 306 191 
<< m2 >>
rect 306 190 307 191 
<< m1 >>
rect 307 190 308 191 
<< m2 >>
rect 307 190 308 191 
<< m2 >>
rect 308 190 309 191 
<< m1 >>
rect 311 190 312 191 
<< m1 >>
rect 313 190 314 191 
<< m1 >>
rect 343 190 344 191 
<< m1 >>
rect 355 190 356 191 
<< m1 >>
rect 19 191 20 192 
<< m1 >>
rect 93 191 94 192 
<< m1 >>
rect 118 191 119 192 
<< m1 >>
rect 121 191 122 192 
<< m1 >>
rect 127 191 128 192 
<< m2 >>
rect 127 191 128 192 
<< m1 >>
rect 142 191 143 192 
<< m1 >>
rect 154 191 155 192 
<< m1 >>
rect 160 191 161 192 
<< m1 >>
rect 172 191 173 192 
<< m1 >>
rect 175 191 176 192 
<< m1 >>
rect 181 191 182 192 
<< m2 >>
rect 181 191 182 192 
<< m1 >>
rect 211 191 212 192 
<< m1 >>
rect 217 191 218 192 
<< m1 >>
rect 226 191 227 192 
<< m1 >>
rect 235 191 236 192 
<< m1 >>
rect 247 191 248 192 
<< m1 >>
rect 254 191 255 192 
<< m1 >>
rect 298 191 299 192 
<< m1 >>
rect 301 191 302 192 
<< m1 >>
rect 307 191 308 192 
<< m2 >>
rect 308 191 309 192 
<< m1 >>
rect 311 191 312 192 
<< m1 >>
rect 313 191 314 192 
<< m1 >>
rect 343 191 344 192 
<< m1 >>
rect 355 191 356 192 
<< pdiffusion >>
rect 12 192 13 193 
<< pdiffusion >>
rect 13 192 14 193 
<< pdiffusion >>
rect 14 192 15 193 
<< pdiffusion >>
rect 15 192 16 193 
<< pdiffusion >>
rect 16 192 17 193 
<< pdiffusion >>
rect 17 192 18 193 
<< m1 >>
rect 19 192 20 193 
<< pdiffusion >>
rect 30 192 31 193 
<< pdiffusion >>
rect 31 192 32 193 
<< pdiffusion >>
rect 32 192 33 193 
<< pdiffusion >>
rect 33 192 34 193 
<< pdiffusion >>
rect 34 192 35 193 
<< pdiffusion >>
rect 35 192 36 193 
<< pdiffusion >>
rect 48 192 49 193 
<< pdiffusion >>
rect 49 192 50 193 
<< pdiffusion >>
rect 50 192 51 193 
<< pdiffusion >>
rect 51 192 52 193 
<< pdiffusion >>
rect 52 192 53 193 
<< pdiffusion >>
rect 53 192 54 193 
<< pdiffusion >>
rect 66 192 67 193 
<< pdiffusion >>
rect 67 192 68 193 
<< pdiffusion >>
rect 68 192 69 193 
<< pdiffusion >>
rect 69 192 70 193 
<< pdiffusion >>
rect 70 192 71 193 
<< pdiffusion >>
rect 71 192 72 193 
<< pdiffusion >>
rect 84 192 85 193 
<< pdiffusion >>
rect 85 192 86 193 
<< pdiffusion >>
rect 86 192 87 193 
<< pdiffusion >>
rect 87 192 88 193 
<< pdiffusion >>
rect 88 192 89 193 
<< pdiffusion >>
rect 89 192 90 193 
<< m1 >>
rect 93 192 94 193 
<< pdiffusion >>
rect 102 192 103 193 
<< pdiffusion >>
rect 103 192 104 193 
<< pdiffusion >>
rect 104 192 105 193 
<< pdiffusion >>
rect 105 192 106 193 
<< pdiffusion >>
rect 106 192 107 193 
<< pdiffusion >>
rect 107 192 108 193 
<< m1 >>
rect 118 192 119 193 
<< pdiffusion >>
rect 120 192 121 193 
<< m1 >>
rect 121 192 122 193 
<< pdiffusion >>
rect 121 192 122 193 
<< pdiffusion >>
rect 122 192 123 193 
<< pdiffusion >>
rect 123 192 124 193 
<< pdiffusion >>
rect 124 192 125 193 
<< pdiffusion >>
rect 125 192 126 193 
<< m1 >>
rect 127 192 128 193 
<< m2 >>
rect 127 192 128 193 
<< pdiffusion >>
rect 138 192 139 193 
<< pdiffusion >>
rect 139 192 140 193 
<< pdiffusion >>
rect 140 192 141 193 
<< pdiffusion >>
rect 141 192 142 193 
<< m1 >>
rect 142 192 143 193 
<< pdiffusion >>
rect 142 192 143 193 
<< pdiffusion >>
rect 143 192 144 193 
<< m1 >>
rect 154 192 155 193 
<< pdiffusion >>
rect 156 192 157 193 
<< pdiffusion >>
rect 157 192 158 193 
<< pdiffusion >>
rect 158 192 159 193 
<< pdiffusion >>
rect 159 192 160 193 
<< m1 >>
rect 160 192 161 193 
<< pdiffusion >>
rect 160 192 161 193 
<< pdiffusion >>
rect 161 192 162 193 
<< m1 >>
rect 172 192 173 193 
<< pdiffusion >>
rect 174 192 175 193 
<< m1 >>
rect 175 192 176 193 
<< pdiffusion >>
rect 175 192 176 193 
<< pdiffusion >>
rect 176 192 177 193 
<< pdiffusion >>
rect 177 192 178 193 
<< pdiffusion >>
rect 178 192 179 193 
<< pdiffusion >>
rect 179 192 180 193 
<< m1 >>
rect 181 192 182 193 
<< m2 >>
rect 181 192 182 193 
<< pdiffusion >>
rect 192 192 193 193 
<< pdiffusion >>
rect 193 192 194 193 
<< pdiffusion >>
rect 194 192 195 193 
<< pdiffusion >>
rect 195 192 196 193 
<< pdiffusion >>
rect 196 192 197 193 
<< pdiffusion >>
rect 197 192 198 193 
<< pdiffusion >>
rect 210 192 211 193 
<< m1 >>
rect 211 192 212 193 
<< pdiffusion >>
rect 211 192 212 193 
<< pdiffusion >>
rect 212 192 213 193 
<< pdiffusion >>
rect 213 192 214 193 
<< pdiffusion >>
rect 214 192 215 193 
<< pdiffusion >>
rect 215 192 216 193 
<< m1 >>
rect 217 192 218 193 
<< m1 >>
rect 226 192 227 193 
<< pdiffusion >>
rect 228 192 229 193 
<< pdiffusion >>
rect 229 192 230 193 
<< pdiffusion >>
rect 230 192 231 193 
<< pdiffusion >>
rect 231 192 232 193 
<< pdiffusion >>
rect 232 192 233 193 
<< pdiffusion >>
rect 233 192 234 193 
<< m1 >>
rect 235 192 236 193 
<< pdiffusion >>
rect 246 192 247 193 
<< m1 >>
rect 247 192 248 193 
<< pdiffusion >>
rect 247 192 248 193 
<< pdiffusion >>
rect 248 192 249 193 
<< pdiffusion >>
rect 249 192 250 193 
<< pdiffusion >>
rect 250 192 251 193 
<< pdiffusion >>
rect 251 192 252 193 
<< m1 >>
rect 254 192 255 193 
<< pdiffusion >>
rect 264 192 265 193 
<< pdiffusion >>
rect 265 192 266 193 
<< pdiffusion >>
rect 266 192 267 193 
<< pdiffusion >>
rect 267 192 268 193 
<< pdiffusion >>
rect 268 192 269 193 
<< pdiffusion >>
rect 269 192 270 193 
<< pdiffusion >>
rect 282 192 283 193 
<< pdiffusion >>
rect 283 192 284 193 
<< pdiffusion >>
rect 284 192 285 193 
<< pdiffusion >>
rect 285 192 286 193 
<< pdiffusion >>
rect 286 192 287 193 
<< pdiffusion >>
rect 287 192 288 193 
<< m1 >>
rect 298 192 299 193 
<< pdiffusion >>
rect 300 192 301 193 
<< m1 >>
rect 301 192 302 193 
<< pdiffusion >>
rect 301 192 302 193 
<< pdiffusion >>
rect 302 192 303 193 
<< pdiffusion >>
rect 303 192 304 193 
<< pdiffusion >>
rect 304 192 305 193 
<< pdiffusion >>
rect 305 192 306 193 
<< m1 >>
rect 307 192 308 193 
<< m2 >>
rect 308 192 309 193 
<< m1 >>
rect 311 192 312 193 
<< m1 >>
rect 313 192 314 193 
<< pdiffusion >>
rect 318 192 319 193 
<< pdiffusion >>
rect 319 192 320 193 
<< pdiffusion >>
rect 320 192 321 193 
<< pdiffusion >>
rect 321 192 322 193 
<< pdiffusion >>
rect 322 192 323 193 
<< pdiffusion >>
rect 323 192 324 193 
<< pdiffusion >>
rect 336 192 337 193 
<< pdiffusion >>
rect 337 192 338 193 
<< pdiffusion >>
rect 338 192 339 193 
<< pdiffusion >>
rect 339 192 340 193 
<< pdiffusion >>
rect 340 192 341 193 
<< pdiffusion >>
rect 341 192 342 193 
<< m1 >>
rect 343 192 344 193 
<< pdiffusion >>
rect 354 192 355 193 
<< m1 >>
rect 355 192 356 193 
<< pdiffusion >>
rect 355 192 356 193 
<< pdiffusion >>
rect 356 192 357 193 
<< pdiffusion >>
rect 357 192 358 193 
<< pdiffusion >>
rect 358 192 359 193 
<< pdiffusion >>
rect 359 192 360 193 
<< pdiffusion >>
rect 372 192 373 193 
<< pdiffusion >>
rect 373 192 374 193 
<< pdiffusion >>
rect 374 192 375 193 
<< pdiffusion >>
rect 375 192 376 193 
<< pdiffusion >>
rect 376 192 377 193 
<< pdiffusion >>
rect 377 192 378 193 
<< pdiffusion >>
rect 390 192 391 193 
<< pdiffusion >>
rect 391 192 392 193 
<< pdiffusion >>
rect 392 192 393 193 
<< pdiffusion >>
rect 393 192 394 193 
<< pdiffusion >>
rect 394 192 395 193 
<< pdiffusion >>
rect 395 192 396 193 
<< pdiffusion >>
rect 408 192 409 193 
<< pdiffusion >>
rect 409 192 410 193 
<< pdiffusion >>
rect 410 192 411 193 
<< pdiffusion >>
rect 411 192 412 193 
<< pdiffusion >>
rect 412 192 413 193 
<< pdiffusion >>
rect 413 192 414 193 
<< pdiffusion >>
rect 426 192 427 193 
<< pdiffusion >>
rect 427 192 428 193 
<< pdiffusion >>
rect 428 192 429 193 
<< pdiffusion >>
rect 429 192 430 193 
<< pdiffusion >>
rect 430 192 431 193 
<< pdiffusion >>
rect 431 192 432 193 
<< pdiffusion >>
rect 444 192 445 193 
<< pdiffusion >>
rect 445 192 446 193 
<< pdiffusion >>
rect 446 192 447 193 
<< pdiffusion >>
rect 447 192 448 193 
<< pdiffusion >>
rect 448 192 449 193 
<< pdiffusion >>
rect 449 192 450 193 
<< pdiffusion >>
rect 12 193 13 194 
<< pdiffusion >>
rect 13 193 14 194 
<< pdiffusion >>
rect 14 193 15 194 
<< pdiffusion >>
rect 15 193 16 194 
<< pdiffusion >>
rect 16 193 17 194 
<< pdiffusion >>
rect 17 193 18 194 
<< m1 >>
rect 19 193 20 194 
<< pdiffusion >>
rect 30 193 31 194 
<< pdiffusion >>
rect 31 193 32 194 
<< pdiffusion >>
rect 32 193 33 194 
<< pdiffusion >>
rect 33 193 34 194 
<< pdiffusion >>
rect 34 193 35 194 
<< pdiffusion >>
rect 35 193 36 194 
<< pdiffusion >>
rect 48 193 49 194 
<< pdiffusion >>
rect 49 193 50 194 
<< pdiffusion >>
rect 50 193 51 194 
<< pdiffusion >>
rect 51 193 52 194 
<< pdiffusion >>
rect 52 193 53 194 
<< pdiffusion >>
rect 53 193 54 194 
<< pdiffusion >>
rect 66 193 67 194 
<< pdiffusion >>
rect 67 193 68 194 
<< pdiffusion >>
rect 68 193 69 194 
<< pdiffusion >>
rect 69 193 70 194 
<< pdiffusion >>
rect 70 193 71 194 
<< pdiffusion >>
rect 71 193 72 194 
<< pdiffusion >>
rect 84 193 85 194 
<< pdiffusion >>
rect 85 193 86 194 
<< pdiffusion >>
rect 86 193 87 194 
<< pdiffusion >>
rect 87 193 88 194 
<< pdiffusion >>
rect 88 193 89 194 
<< pdiffusion >>
rect 89 193 90 194 
<< m1 >>
rect 93 193 94 194 
<< pdiffusion >>
rect 102 193 103 194 
<< pdiffusion >>
rect 103 193 104 194 
<< pdiffusion >>
rect 104 193 105 194 
<< pdiffusion >>
rect 105 193 106 194 
<< pdiffusion >>
rect 106 193 107 194 
<< pdiffusion >>
rect 107 193 108 194 
<< m1 >>
rect 118 193 119 194 
<< pdiffusion >>
rect 120 193 121 194 
<< pdiffusion >>
rect 121 193 122 194 
<< pdiffusion >>
rect 122 193 123 194 
<< pdiffusion >>
rect 123 193 124 194 
<< pdiffusion >>
rect 124 193 125 194 
<< pdiffusion >>
rect 125 193 126 194 
<< m1 >>
rect 127 193 128 194 
<< m2 >>
rect 127 193 128 194 
<< pdiffusion >>
rect 138 193 139 194 
<< pdiffusion >>
rect 139 193 140 194 
<< pdiffusion >>
rect 140 193 141 194 
<< pdiffusion >>
rect 141 193 142 194 
<< pdiffusion >>
rect 142 193 143 194 
<< pdiffusion >>
rect 143 193 144 194 
<< m1 >>
rect 154 193 155 194 
<< pdiffusion >>
rect 156 193 157 194 
<< pdiffusion >>
rect 157 193 158 194 
<< pdiffusion >>
rect 158 193 159 194 
<< pdiffusion >>
rect 159 193 160 194 
<< pdiffusion >>
rect 160 193 161 194 
<< pdiffusion >>
rect 161 193 162 194 
<< m1 >>
rect 172 193 173 194 
<< pdiffusion >>
rect 174 193 175 194 
<< pdiffusion >>
rect 175 193 176 194 
<< pdiffusion >>
rect 176 193 177 194 
<< pdiffusion >>
rect 177 193 178 194 
<< pdiffusion >>
rect 178 193 179 194 
<< pdiffusion >>
rect 179 193 180 194 
<< m1 >>
rect 181 193 182 194 
<< m2 >>
rect 181 193 182 194 
<< pdiffusion >>
rect 192 193 193 194 
<< pdiffusion >>
rect 193 193 194 194 
<< pdiffusion >>
rect 194 193 195 194 
<< pdiffusion >>
rect 195 193 196 194 
<< pdiffusion >>
rect 196 193 197 194 
<< pdiffusion >>
rect 197 193 198 194 
<< pdiffusion >>
rect 210 193 211 194 
<< pdiffusion >>
rect 211 193 212 194 
<< pdiffusion >>
rect 212 193 213 194 
<< pdiffusion >>
rect 213 193 214 194 
<< pdiffusion >>
rect 214 193 215 194 
<< pdiffusion >>
rect 215 193 216 194 
<< m1 >>
rect 217 193 218 194 
<< m1 >>
rect 226 193 227 194 
<< pdiffusion >>
rect 228 193 229 194 
<< pdiffusion >>
rect 229 193 230 194 
<< pdiffusion >>
rect 230 193 231 194 
<< pdiffusion >>
rect 231 193 232 194 
<< pdiffusion >>
rect 232 193 233 194 
<< pdiffusion >>
rect 233 193 234 194 
<< m1 >>
rect 235 193 236 194 
<< pdiffusion >>
rect 246 193 247 194 
<< pdiffusion >>
rect 247 193 248 194 
<< pdiffusion >>
rect 248 193 249 194 
<< pdiffusion >>
rect 249 193 250 194 
<< pdiffusion >>
rect 250 193 251 194 
<< pdiffusion >>
rect 251 193 252 194 
<< m1 >>
rect 254 193 255 194 
<< pdiffusion >>
rect 264 193 265 194 
<< pdiffusion >>
rect 265 193 266 194 
<< pdiffusion >>
rect 266 193 267 194 
<< pdiffusion >>
rect 267 193 268 194 
<< pdiffusion >>
rect 268 193 269 194 
<< pdiffusion >>
rect 269 193 270 194 
<< pdiffusion >>
rect 282 193 283 194 
<< pdiffusion >>
rect 283 193 284 194 
<< pdiffusion >>
rect 284 193 285 194 
<< pdiffusion >>
rect 285 193 286 194 
<< pdiffusion >>
rect 286 193 287 194 
<< pdiffusion >>
rect 287 193 288 194 
<< m1 >>
rect 298 193 299 194 
<< pdiffusion >>
rect 300 193 301 194 
<< pdiffusion >>
rect 301 193 302 194 
<< pdiffusion >>
rect 302 193 303 194 
<< pdiffusion >>
rect 303 193 304 194 
<< pdiffusion >>
rect 304 193 305 194 
<< pdiffusion >>
rect 305 193 306 194 
<< m1 >>
rect 307 193 308 194 
<< m2 >>
rect 308 193 309 194 
<< m1 >>
rect 311 193 312 194 
<< m1 >>
rect 313 193 314 194 
<< pdiffusion >>
rect 318 193 319 194 
<< pdiffusion >>
rect 319 193 320 194 
<< pdiffusion >>
rect 320 193 321 194 
<< pdiffusion >>
rect 321 193 322 194 
<< pdiffusion >>
rect 322 193 323 194 
<< pdiffusion >>
rect 323 193 324 194 
<< pdiffusion >>
rect 336 193 337 194 
<< pdiffusion >>
rect 337 193 338 194 
<< pdiffusion >>
rect 338 193 339 194 
<< pdiffusion >>
rect 339 193 340 194 
<< pdiffusion >>
rect 340 193 341 194 
<< pdiffusion >>
rect 341 193 342 194 
<< m1 >>
rect 343 193 344 194 
<< pdiffusion >>
rect 354 193 355 194 
<< pdiffusion >>
rect 355 193 356 194 
<< pdiffusion >>
rect 356 193 357 194 
<< pdiffusion >>
rect 357 193 358 194 
<< pdiffusion >>
rect 358 193 359 194 
<< pdiffusion >>
rect 359 193 360 194 
<< pdiffusion >>
rect 372 193 373 194 
<< pdiffusion >>
rect 373 193 374 194 
<< pdiffusion >>
rect 374 193 375 194 
<< pdiffusion >>
rect 375 193 376 194 
<< pdiffusion >>
rect 376 193 377 194 
<< pdiffusion >>
rect 377 193 378 194 
<< pdiffusion >>
rect 390 193 391 194 
<< pdiffusion >>
rect 391 193 392 194 
<< pdiffusion >>
rect 392 193 393 194 
<< pdiffusion >>
rect 393 193 394 194 
<< pdiffusion >>
rect 394 193 395 194 
<< pdiffusion >>
rect 395 193 396 194 
<< pdiffusion >>
rect 408 193 409 194 
<< pdiffusion >>
rect 409 193 410 194 
<< pdiffusion >>
rect 410 193 411 194 
<< pdiffusion >>
rect 411 193 412 194 
<< pdiffusion >>
rect 412 193 413 194 
<< pdiffusion >>
rect 413 193 414 194 
<< pdiffusion >>
rect 426 193 427 194 
<< pdiffusion >>
rect 427 193 428 194 
<< pdiffusion >>
rect 428 193 429 194 
<< pdiffusion >>
rect 429 193 430 194 
<< pdiffusion >>
rect 430 193 431 194 
<< pdiffusion >>
rect 431 193 432 194 
<< pdiffusion >>
rect 444 193 445 194 
<< pdiffusion >>
rect 445 193 446 194 
<< pdiffusion >>
rect 446 193 447 194 
<< pdiffusion >>
rect 447 193 448 194 
<< pdiffusion >>
rect 448 193 449 194 
<< pdiffusion >>
rect 449 193 450 194 
<< pdiffusion >>
rect 12 194 13 195 
<< pdiffusion >>
rect 13 194 14 195 
<< pdiffusion >>
rect 14 194 15 195 
<< pdiffusion >>
rect 15 194 16 195 
<< pdiffusion >>
rect 16 194 17 195 
<< pdiffusion >>
rect 17 194 18 195 
<< m1 >>
rect 19 194 20 195 
<< pdiffusion >>
rect 30 194 31 195 
<< pdiffusion >>
rect 31 194 32 195 
<< pdiffusion >>
rect 32 194 33 195 
<< pdiffusion >>
rect 33 194 34 195 
<< pdiffusion >>
rect 34 194 35 195 
<< pdiffusion >>
rect 35 194 36 195 
<< pdiffusion >>
rect 48 194 49 195 
<< pdiffusion >>
rect 49 194 50 195 
<< pdiffusion >>
rect 50 194 51 195 
<< pdiffusion >>
rect 51 194 52 195 
<< pdiffusion >>
rect 52 194 53 195 
<< pdiffusion >>
rect 53 194 54 195 
<< pdiffusion >>
rect 66 194 67 195 
<< pdiffusion >>
rect 67 194 68 195 
<< pdiffusion >>
rect 68 194 69 195 
<< pdiffusion >>
rect 69 194 70 195 
<< pdiffusion >>
rect 70 194 71 195 
<< pdiffusion >>
rect 71 194 72 195 
<< pdiffusion >>
rect 84 194 85 195 
<< pdiffusion >>
rect 85 194 86 195 
<< pdiffusion >>
rect 86 194 87 195 
<< pdiffusion >>
rect 87 194 88 195 
<< pdiffusion >>
rect 88 194 89 195 
<< pdiffusion >>
rect 89 194 90 195 
<< m1 >>
rect 93 194 94 195 
<< pdiffusion >>
rect 102 194 103 195 
<< pdiffusion >>
rect 103 194 104 195 
<< pdiffusion >>
rect 104 194 105 195 
<< pdiffusion >>
rect 105 194 106 195 
<< pdiffusion >>
rect 106 194 107 195 
<< pdiffusion >>
rect 107 194 108 195 
<< m1 >>
rect 118 194 119 195 
<< pdiffusion >>
rect 120 194 121 195 
<< pdiffusion >>
rect 121 194 122 195 
<< pdiffusion >>
rect 122 194 123 195 
<< pdiffusion >>
rect 123 194 124 195 
<< pdiffusion >>
rect 124 194 125 195 
<< pdiffusion >>
rect 125 194 126 195 
<< m1 >>
rect 127 194 128 195 
<< m2 >>
rect 127 194 128 195 
<< pdiffusion >>
rect 138 194 139 195 
<< pdiffusion >>
rect 139 194 140 195 
<< pdiffusion >>
rect 140 194 141 195 
<< pdiffusion >>
rect 141 194 142 195 
<< pdiffusion >>
rect 142 194 143 195 
<< pdiffusion >>
rect 143 194 144 195 
<< m1 >>
rect 154 194 155 195 
<< pdiffusion >>
rect 156 194 157 195 
<< pdiffusion >>
rect 157 194 158 195 
<< pdiffusion >>
rect 158 194 159 195 
<< pdiffusion >>
rect 159 194 160 195 
<< pdiffusion >>
rect 160 194 161 195 
<< pdiffusion >>
rect 161 194 162 195 
<< m1 >>
rect 172 194 173 195 
<< pdiffusion >>
rect 174 194 175 195 
<< pdiffusion >>
rect 175 194 176 195 
<< pdiffusion >>
rect 176 194 177 195 
<< pdiffusion >>
rect 177 194 178 195 
<< pdiffusion >>
rect 178 194 179 195 
<< pdiffusion >>
rect 179 194 180 195 
<< m1 >>
rect 181 194 182 195 
<< m2 >>
rect 181 194 182 195 
<< pdiffusion >>
rect 192 194 193 195 
<< pdiffusion >>
rect 193 194 194 195 
<< pdiffusion >>
rect 194 194 195 195 
<< pdiffusion >>
rect 195 194 196 195 
<< pdiffusion >>
rect 196 194 197 195 
<< pdiffusion >>
rect 197 194 198 195 
<< pdiffusion >>
rect 210 194 211 195 
<< pdiffusion >>
rect 211 194 212 195 
<< pdiffusion >>
rect 212 194 213 195 
<< pdiffusion >>
rect 213 194 214 195 
<< pdiffusion >>
rect 214 194 215 195 
<< pdiffusion >>
rect 215 194 216 195 
<< m1 >>
rect 217 194 218 195 
<< m1 >>
rect 226 194 227 195 
<< pdiffusion >>
rect 228 194 229 195 
<< pdiffusion >>
rect 229 194 230 195 
<< pdiffusion >>
rect 230 194 231 195 
<< pdiffusion >>
rect 231 194 232 195 
<< pdiffusion >>
rect 232 194 233 195 
<< pdiffusion >>
rect 233 194 234 195 
<< m1 >>
rect 235 194 236 195 
<< pdiffusion >>
rect 246 194 247 195 
<< pdiffusion >>
rect 247 194 248 195 
<< pdiffusion >>
rect 248 194 249 195 
<< pdiffusion >>
rect 249 194 250 195 
<< pdiffusion >>
rect 250 194 251 195 
<< pdiffusion >>
rect 251 194 252 195 
<< m1 >>
rect 254 194 255 195 
<< pdiffusion >>
rect 264 194 265 195 
<< pdiffusion >>
rect 265 194 266 195 
<< pdiffusion >>
rect 266 194 267 195 
<< pdiffusion >>
rect 267 194 268 195 
<< pdiffusion >>
rect 268 194 269 195 
<< pdiffusion >>
rect 269 194 270 195 
<< pdiffusion >>
rect 282 194 283 195 
<< pdiffusion >>
rect 283 194 284 195 
<< pdiffusion >>
rect 284 194 285 195 
<< pdiffusion >>
rect 285 194 286 195 
<< pdiffusion >>
rect 286 194 287 195 
<< pdiffusion >>
rect 287 194 288 195 
<< m1 >>
rect 298 194 299 195 
<< pdiffusion >>
rect 300 194 301 195 
<< pdiffusion >>
rect 301 194 302 195 
<< pdiffusion >>
rect 302 194 303 195 
<< pdiffusion >>
rect 303 194 304 195 
<< pdiffusion >>
rect 304 194 305 195 
<< pdiffusion >>
rect 305 194 306 195 
<< m1 >>
rect 307 194 308 195 
<< m2 >>
rect 308 194 309 195 
<< m1 >>
rect 311 194 312 195 
<< m1 >>
rect 313 194 314 195 
<< pdiffusion >>
rect 318 194 319 195 
<< pdiffusion >>
rect 319 194 320 195 
<< pdiffusion >>
rect 320 194 321 195 
<< pdiffusion >>
rect 321 194 322 195 
<< pdiffusion >>
rect 322 194 323 195 
<< pdiffusion >>
rect 323 194 324 195 
<< pdiffusion >>
rect 336 194 337 195 
<< pdiffusion >>
rect 337 194 338 195 
<< pdiffusion >>
rect 338 194 339 195 
<< pdiffusion >>
rect 339 194 340 195 
<< pdiffusion >>
rect 340 194 341 195 
<< pdiffusion >>
rect 341 194 342 195 
<< m1 >>
rect 343 194 344 195 
<< pdiffusion >>
rect 354 194 355 195 
<< pdiffusion >>
rect 355 194 356 195 
<< pdiffusion >>
rect 356 194 357 195 
<< pdiffusion >>
rect 357 194 358 195 
<< pdiffusion >>
rect 358 194 359 195 
<< pdiffusion >>
rect 359 194 360 195 
<< pdiffusion >>
rect 372 194 373 195 
<< pdiffusion >>
rect 373 194 374 195 
<< pdiffusion >>
rect 374 194 375 195 
<< pdiffusion >>
rect 375 194 376 195 
<< pdiffusion >>
rect 376 194 377 195 
<< pdiffusion >>
rect 377 194 378 195 
<< pdiffusion >>
rect 390 194 391 195 
<< pdiffusion >>
rect 391 194 392 195 
<< pdiffusion >>
rect 392 194 393 195 
<< pdiffusion >>
rect 393 194 394 195 
<< pdiffusion >>
rect 394 194 395 195 
<< pdiffusion >>
rect 395 194 396 195 
<< pdiffusion >>
rect 408 194 409 195 
<< pdiffusion >>
rect 409 194 410 195 
<< pdiffusion >>
rect 410 194 411 195 
<< pdiffusion >>
rect 411 194 412 195 
<< pdiffusion >>
rect 412 194 413 195 
<< pdiffusion >>
rect 413 194 414 195 
<< pdiffusion >>
rect 426 194 427 195 
<< pdiffusion >>
rect 427 194 428 195 
<< pdiffusion >>
rect 428 194 429 195 
<< pdiffusion >>
rect 429 194 430 195 
<< pdiffusion >>
rect 430 194 431 195 
<< pdiffusion >>
rect 431 194 432 195 
<< pdiffusion >>
rect 444 194 445 195 
<< pdiffusion >>
rect 445 194 446 195 
<< pdiffusion >>
rect 446 194 447 195 
<< pdiffusion >>
rect 447 194 448 195 
<< pdiffusion >>
rect 448 194 449 195 
<< pdiffusion >>
rect 449 194 450 195 
<< pdiffusion >>
rect 12 195 13 196 
<< pdiffusion >>
rect 13 195 14 196 
<< pdiffusion >>
rect 14 195 15 196 
<< pdiffusion >>
rect 15 195 16 196 
<< pdiffusion >>
rect 16 195 17 196 
<< pdiffusion >>
rect 17 195 18 196 
<< m1 >>
rect 19 195 20 196 
<< pdiffusion >>
rect 30 195 31 196 
<< pdiffusion >>
rect 31 195 32 196 
<< pdiffusion >>
rect 32 195 33 196 
<< pdiffusion >>
rect 33 195 34 196 
<< pdiffusion >>
rect 34 195 35 196 
<< pdiffusion >>
rect 35 195 36 196 
<< pdiffusion >>
rect 48 195 49 196 
<< pdiffusion >>
rect 49 195 50 196 
<< pdiffusion >>
rect 50 195 51 196 
<< pdiffusion >>
rect 51 195 52 196 
<< pdiffusion >>
rect 52 195 53 196 
<< pdiffusion >>
rect 53 195 54 196 
<< pdiffusion >>
rect 66 195 67 196 
<< pdiffusion >>
rect 67 195 68 196 
<< pdiffusion >>
rect 68 195 69 196 
<< pdiffusion >>
rect 69 195 70 196 
<< pdiffusion >>
rect 70 195 71 196 
<< pdiffusion >>
rect 71 195 72 196 
<< pdiffusion >>
rect 84 195 85 196 
<< pdiffusion >>
rect 85 195 86 196 
<< pdiffusion >>
rect 86 195 87 196 
<< pdiffusion >>
rect 87 195 88 196 
<< pdiffusion >>
rect 88 195 89 196 
<< pdiffusion >>
rect 89 195 90 196 
<< m1 >>
rect 93 195 94 196 
<< pdiffusion >>
rect 102 195 103 196 
<< pdiffusion >>
rect 103 195 104 196 
<< pdiffusion >>
rect 104 195 105 196 
<< pdiffusion >>
rect 105 195 106 196 
<< pdiffusion >>
rect 106 195 107 196 
<< pdiffusion >>
rect 107 195 108 196 
<< m1 >>
rect 118 195 119 196 
<< pdiffusion >>
rect 120 195 121 196 
<< pdiffusion >>
rect 121 195 122 196 
<< pdiffusion >>
rect 122 195 123 196 
<< pdiffusion >>
rect 123 195 124 196 
<< pdiffusion >>
rect 124 195 125 196 
<< pdiffusion >>
rect 125 195 126 196 
<< m1 >>
rect 127 195 128 196 
<< m2 >>
rect 127 195 128 196 
<< pdiffusion >>
rect 138 195 139 196 
<< pdiffusion >>
rect 139 195 140 196 
<< pdiffusion >>
rect 140 195 141 196 
<< pdiffusion >>
rect 141 195 142 196 
<< pdiffusion >>
rect 142 195 143 196 
<< pdiffusion >>
rect 143 195 144 196 
<< m1 >>
rect 154 195 155 196 
<< pdiffusion >>
rect 156 195 157 196 
<< pdiffusion >>
rect 157 195 158 196 
<< pdiffusion >>
rect 158 195 159 196 
<< pdiffusion >>
rect 159 195 160 196 
<< pdiffusion >>
rect 160 195 161 196 
<< pdiffusion >>
rect 161 195 162 196 
<< m1 >>
rect 172 195 173 196 
<< pdiffusion >>
rect 174 195 175 196 
<< pdiffusion >>
rect 175 195 176 196 
<< pdiffusion >>
rect 176 195 177 196 
<< pdiffusion >>
rect 177 195 178 196 
<< pdiffusion >>
rect 178 195 179 196 
<< pdiffusion >>
rect 179 195 180 196 
<< m1 >>
rect 181 195 182 196 
<< m2 >>
rect 181 195 182 196 
<< pdiffusion >>
rect 192 195 193 196 
<< pdiffusion >>
rect 193 195 194 196 
<< pdiffusion >>
rect 194 195 195 196 
<< pdiffusion >>
rect 195 195 196 196 
<< pdiffusion >>
rect 196 195 197 196 
<< pdiffusion >>
rect 197 195 198 196 
<< pdiffusion >>
rect 210 195 211 196 
<< pdiffusion >>
rect 211 195 212 196 
<< pdiffusion >>
rect 212 195 213 196 
<< pdiffusion >>
rect 213 195 214 196 
<< pdiffusion >>
rect 214 195 215 196 
<< pdiffusion >>
rect 215 195 216 196 
<< m1 >>
rect 217 195 218 196 
<< m1 >>
rect 226 195 227 196 
<< pdiffusion >>
rect 228 195 229 196 
<< pdiffusion >>
rect 229 195 230 196 
<< pdiffusion >>
rect 230 195 231 196 
<< pdiffusion >>
rect 231 195 232 196 
<< pdiffusion >>
rect 232 195 233 196 
<< pdiffusion >>
rect 233 195 234 196 
<< m1 >>
rect 235 195 236 196 
<< pdiffusion >>
rect 246 195 247 196 
<< pdiffusion >>
rect 247 195 248 196 
<< pdiffusion >>
rect 248 195 249 196 
<< pdiffusion >>
rect 249 195 250 196 
<< pdiffusion >>
rect 250 195 251 196 
<< pdiffusion >>
rect 251 195 252 196 
<< m1 >>
rect 254 195 255 196 
<< pdiffusion >>
rect 264 195 265 196 
<< pdiffusion >>
rect 265 195 266 196 
<< pdiffusion >>
rect 266 195 267 196 
<< pdiffusion >>
rect 267 195 268 196 
<< pdiffusion >>
rect 268 195 269 196 
<< pdiffusion >>
rect 269 195 270 196 
<< pdiffusion >>
rect 282 195 283 196 
<< pdiffusion >>
rect 283 195 284 196 
<< pdiffusion >>
rect 284 195 285 196 
<< pdiffusion >>
rect 285 195 286 196 
<< pdiffusion >>
rect 286 195 287 196 
<< pdiffusion >>
rect 287 195 288 196 
<< m1 >>
rect 298 195 299 196 
<< pdiffusion >>
rect 300 195 301 196 
<< pdiffusion >>
rect 301 195 302 196 
<< pdiffusion >>
rect 302 195 303 196 
<< pdiffusion >>
rect 303 195 304 196 
<< pdiffusion >>
rect 304 195 305 196 
<< pdiffusion >>
rect 305 195 306 196 
<< m1 >>
rect 307 195 308 196 
<< m2 >>
rect 308 195 309 196 
<< m1 >>
rect 311 195 312 196 
<< m1 >>
rect 313 195 314 196 
<< pdiffusion >>
rect 318 195 319 196 
<< pdiffusion >>
rect 319 195 320 196 
<< pdiffusion >>
rect 320 195 321 196 
<< pdiffusion >>
rect 321 195 322 196 
<< pdiffusion >>
rect 322 195 323 196 
<< pdiffusion >>
rect 323 195 324 196 
<< pdiffusion >>
rect 336 195 337 196 
<< pdiffusion >>
rect 337 195 338 196 
<< pdiffusion >>
rect 338 195 339 196 
<< pdiffusion >>
rect 339 195 340 196 
<< pdiffusion >>
rect 340 195 341 196 
<< pdiffusion >>
rect 341 195 342 196 
<< m1 >>
rect 343 195 344 196 
<< pdiffusion >>
rect 354 195 355 196 
<< pdiffusion >>
rect 355 195 356 196 
<< pdiffusion >>
rect 356 195 357 196 
<< pdiffusion >>
rect 357 195 358 196 
<< pdiffusion >>
rect 358 195 359 196 
<< pdiffusion >>
rect 359 195 360 196 
<< pdiffusion >>
rect 372 195 373 196 
<< pdiffusion >>
rect 373 195 374 196 
<< pdiffusion >>
rect 374 195 375 196 
<< pdiffusion >>
rect 375 195 376 196 
<< pdiffusion >>
rect 376 195 377 196 
<< pdiffusion >>
rect 377 195 378 196 
<< pdiffusion >>
rect 390 195 391 196 
<< pdiffusion >>
rect 391 195 392 196 
<< pdiffusion >>
rect 392 195 393 196 
<< pdiffusion >>
rect 393 195 394 196 
<< pdiffusion >>
rect 394 195 395 196 
<< pdiffusion >>
rect 395 195 396 196 
<< pdiffusion >>
rect 408 195 409 196 
<< pdiffusion >>
rect 409 195 410 196 
<< pdiffusion >>
rect 410 195 411 196 
<< pdiffusion >>
rect 411 195 412 196 
<< pdiffusion >>
rect 412 195 413 196 
<< pdiffusion >>
rect 413 195 414 196 
<< pdiffusion >>
rect 426 195 427 196 
<< pdiffusion >>
rect 427 195 428 196 
<< pdiffusion >>
rect 428 195 429 196 
<< pdiffusion >>
rect 429 195 430 196 
<< pdiffusion >>
rect 430 195 431 196 
<< pdiffusion >>
rect 431 195 432 196 
<< pdiffusion >>
rect 444 195 445 196 
<< pdiffusion >>
rect 445 195 446 196 
<< pdiffusion >>
rect 446 195 447 196 
<< pdiffusion >>
rect 447 195 448 196 
<< pdiffusion >>
rect 448 195 449 196 
<< pdiffusion >>
rect 449 195 450 196 
<< pdiffusion >>
rect 12 196 13 197 
<< pdiffusion >>
rect 13 196 14 197 
<< pdiffusion >>
rect 14 196 15 197 
<< pdiffusion >>
rect 15 196 16 197 
<< pdiffusion >>
rect 16 196 17 197 
<< pdiffusion >>
rect 17 196 18 197 
<< m1 >>
rect 19 196 20 197 
<< pdiffusion >>
rect 30 196 31 197 
<< pdiffusion >>
rect 31 196 32 197 
<< pdiffusion >>
rect 32 196 33 197 
<< pdiffusion >>
rect 33 196 34 197 
<< pdiffusion >>
rect 34 196 35 197 
<< pdiffusion >>
rect 35 196 36 197 
<< pdiffusion >>
rect 48 196 49 197 
<< pdiffusion >>
rect 49 196 50 197 
<< pdiffusion >>
rect 50 196 51 197 
<< pdiffusion >>
rect 51 196 52 197 
<< pdiffusion >>
rect 52 196 53 197 
<< pdiffusion >>
rect 53 196 54 197 
<< pdiffusion >>
rect 66 196 67 197 
<< pdiffusion >>
rect 67 196 68 197 
<< pdiffusion >>
rect 68 196 69 197 
<< pdiffusion >>
rect 69 196 70 197 
<< pdiffusion >>
rect 70 196 71 197 
<< pdiffusion >>
rect 71 196 72 197 
<< pdiffusion >>
rect 84 196 85 197 
<< pdiffusion >>
rect 85 196 86 197 
<< pdiffusion >>
rect 86 196 87 197 
<< pdiffusion >>
rect 87 196 88 197 
<< pdiffusion >>
rect 88 196 89 197 
<< pdiffusion >>
rect 89 196 90 197 
<< m1 >>
rect 93 196 94 197 
<< pdiffusion >>
rect 102 196 103 197 
<< pdiffusion >>
rect 103 196 104 197 
<< pdiffusion >>
rect 104 196 105 197 
<< pdiffusion >>
rect 105 196 106 197 
<< pdiffusion >>
rect 106 196 107 197 
<< pdiffusion >>
rect 107 196 108 197 
<< m1 >>
rect 118 196 119 197 
<< pdiffusion >>
rect 120 196 121 197 
<< pdiffusion >>
rect 121 196 122 197 
<< pdiffusion >>
rect 122 196 123 197 
<< pdiffusion >>
rect 123 196 124 197 
<< pdiffusion >>
rect 124 196 125 197 
<< pdiffusion >>
rect 125 196 126 197 
<< m1 >>
rect 127 196 128 197 
<< m2 >>
rect 127 196 128 197 
<< pdiffusion >>
rect 138 196 139 197 
<< pdiffusion >>
rect 139 196 140 197 
<< pdiffusion >>
rect 140 196 141 197 
<< pdiffusion >>
rect 141 196 142 197 
<< pdiffusion >>
rect 142 196 143 197 
<< pdiffusion >>
rect 143 196 144 197 
<< m1 >>
rect 154 196 155 197 
<< pdiffusion >>
rect 156 196 157 197 
<< pdiffusion >>
rect 157 196 158 197 
<< pdiffusion >>
rect 158 196 159 197 
<< pdiffusion >>
rect 159 196 160 197 
<< pdiffusion >>
rect 160 196 161 197 
<< pdiffusion >>
rect 161 196 162 197 
<< m1 >>
rect 172 196 173 197 
<< pdiffusion >>
rect 174 196 175 197 
<< pdiffusion >>
rect 175 196 176 197 
<< pdiffusion >>
rect 176 196 177 197 
<< pdiffusion >>
rect 177 196 178 197 
<< pdiffusion >>
rect 178 196 179 197 
<< pdiffusion >>
rect 179 196 180 197 
<< m1 >>
rect 181 196 182 197 
<< m2 >>
rect 181 196 182 197 
<< pdiffusion >>
rect 192 196 193 197 
<< pdiffusion >>
rect 193 196 194 197 
<< pdiffusion >>
rect 194 196 195 197 
<< pdiffusion >>
rect 195 196 196 197 
<< pdiffusion >>
rect 196 196 197 197 
<< pdiffusion >>
rect 197 196 198 197 
<< pdiffusion >>
rect 210 196 211 197 
<< pdiffusion >>
rect 211 196 212 197 
<< pdiffusion >>
rect 212 196 213 197 
<< pdiffusion >>
rect 213 196 214 197 
<< pdiffusion >>
rect 214 196 215 197 
<< pdiffusion >>
rect 215 196 216 197 
<< m1 >>
rect 217 196 218 197 
<< m1 >>
rect 226 196 227 197 
<< pdiffusion >>
rect 228 196 229 197 
<< pdiffusion >>
rect 229 196 230 197 
<< pdiffusion >>
rect 230 196 231 197 
<< pdiffusion >>
rect 231 196 232 197 
<< pdiffusion >>
rect 232 196 233 197 
<< pdiffusion >>
rect 233 196 234 197 
<< m1 >>
rect 235 196 236 197 
<< pdiffusion >>
rect 246 196 247 197 
<< pdiffusion >>
rect 247 196 248 197 
<< pdiffusion >>
rect 248 196 249 197 
<< pdiffusion >>
rect 249 196 250 197 
<< pdiffusion >>
rect 250 196 251 197 
<< pdiffusion >>
rect 251 196 252 197 
<< m1 >>
rect 254 196 255 197 
<< pdiffusion >>
rect 264 196 265 197 
<< pdiffusion >>
rect 265 196 266 197 
<< pdiffusion >>
rect 266 196 267 197 
<< pdiffusion >>
rect 267 196 268 197 
<< pdiffusion >>
rect 268 196 269 197 
<< pdiffusion >>
rect 269 196 270 197 
<< pdiffusion >>
rect 282 196 283 197 
<< pdiffusion >>
rect 283 196 284 197 
<< pdiffusion >>
rect 284 196 285 197 
<< pdiffusion >>
rect 285 196 286 197 
<< pdiffusion >>
rect 286 196 287 197 
<< pdiffusion >>
rect 287 196 288 197 
<< m1 >>
rect 298 196 299 197 
<< pdiffusion >>
rect 300 196 301 197 
<< pdiffusion >>
rect 301 196 302 197 
<< pdiffusion >>
rect 302 196 303 197 
<< pdiffusion >>
rect 303 196 304 197 
<< pdiffusion >>
rect 304 196 305 197 
<< pdiffusion >>
rect 305 196 306 197 
<< m1 >>
rect 307 196 308 197 
<< m2 >>
rect 308 196 309 197 
<< m1 >>
rect 311 196 312 197 
<< m1 >>
rect 313 196 314 197 
<< pdiffusion >>
rect 318 196 319 197 
<< pdiffusion >>
rect 319 196 320 197 
<< pdiffusion >>
rect 320 196 321 197 
<< pdiffusion >>
rect 321 196 322 197 
<< pdiffusion >>
rect 322 196 323 197 
<< pdiffusion >>
rect 323 196 324 197 
<< pdiffusion >>
rect 336 196 337 197 
<< pdiffusion >>
rect 337 196 338 197 
<< pdiffusion >>
rect 338 196 339 197 
<< pdiffusion >>
rect 339 196 340 197 
<< pdiffusion >>
rect 340 196 341 197 
<< pdiffusion >>
rect 341 196 342 197 
<< m1 >>
rect 343 196 344 197 
<< pdiffusion >>
rect 354 196 355 197 
<< pdiffusion >>
rect 355 196 356 197 
<< pdiffusion >>
rect 356 196 357 197 
<< pdiffusion >>
rect 357 196 358 197 
<< pdiffusion >>
rect 358 196 359 197 
<< pdiffusion >>
rect 359 196 360 197 
<< pdiffusion >>
rect 372 196 373 197 
<< pdiffusion >>
rect 373 196 374 197 
<< pdiffusion >>
rect 374 196 375 197 
<< pdiffusion >>
rect 375 196 376 197 
<< pdiffusion >>
rect 376 196 377 197 
<< pdiffusion >>
rect 377 196 378 197 
<< pdiffusion >>
rect 390 196 391 197 
<< pdiffusion >>
rect 391 196 392 197 
<< pdiffusion >>
rect 392 196 393 197 
<< pdiffusion >>
rect 393 196 394 197 
<< pdiffusion >>
rect 394 196 395 197 
<< pdiffusion >>
rect 395 196 396 197 
<< pdiffusion >>
rect 408 196 409 197 
<< pdiffusion >>
rect 409 196 410 197 
<< pdiffusion >>
rect 410 196 411 197 
<< pdiffusion >>
rect 411 196 412 197 
<< pdiffusion >>
rect 412 196 413 197 
<< pdiffusion >>
rect 413 196 414 197 
<< pdiffusion >>
rect 426 196 427 197 
<< pdiffusion >>
rect 427 196 428 197 
<< pdiffusion >>
rect 428 196 429 197 
<< pdiffusion >>
rect 429 196 430 197 
<< pdiffusion >>
rect 430 196 431 197 
<< pdiffusion >>
rect 431 196 432 197 
<< pdiffusion >>
rect 444 196 445 197 
<< pdiffusion >>
rect 445 196 446 197 
<< pdiffusion >>
rect 446 196 447 197 
<< pdiffusion >>
rect 447 196 448 197 
<< pdiffusion >>
rect 448 196 449 197 
<< pdiffusion >>
rect 449 196 450 197 
<< pdiffusion >>
rect 12 197 13 198 
<< pdiffusion >>
rect 13 197 14 198 
<< pdiffusion >>
rect 14 197 15 198 
<< pdiffusion >>
rect 15 197 16 198 
<< m1 >>
rect 16 197 17 198 
<< pdiffusion >>
rect 16 197 17 198 
<< pdiffusion >>
rect 17 197 18 198 
<< m1 >>
rect 19 197 20 198 
<< pdiffusion >>
rect 30 197 31 198 
<< pdiffusion >>
rect 31 197 32 198 
<< pdiffusion >>
rect 32 197 33 198 
<< pdiffusion >>
rect 33 197 34 198 
<< pdiffusion >>
rect 34 197 35 198 
<< pdiffusion >>
rect 35 197 36 198 
<< pdiffusion >>
rect 48 197 49 198 
<< m1 >>
rect 49 197 50 198 
<< pdiffusion >>
rect 49 197 50 198 
<< pdiffusion >>
rect 50 197 51 198 
<< pdiffusion >>
rect 51 197 52 198 
<< pdiffusion >>
rect 52 197 53 198 
<< pdiffusion >>
rect 53 197 54 198 
<< pdiffusion >>
rect 66 197 67 198 
<< pdiffusion >>
rect 67 197 68 198 
<< pdiffusion >>
rect 68 197 69 198 
<< pdiffusion >>
rect 69 197 70 198 
<< pdiffusion >>
rect 70 197 71 198 
<< pdiffusion >>
rect 71 197 72 198 
<< pdiffusion >>
rect 84 197 85 198 
<< pdiffusion >>
rect 85 197 86 198 
<< pdiffusion >>
rect 86 197 87 198 
<< pdiffusion >>
rect 87 197 88 198 
<< pdiffusion >>
rect 88 197 89 198 
<< pdiffusion >>
rect 89 197 90 198 
<< m1 >>
rect 93 197 94 198 
<< pdiffusion >>
rect 102 197 103 198 
<< pdiffusion >>
rect 103 197 104 198 
<< pdiffusion >>
rect 104 197 105 198 
<< pdiffusion >>
rect 105 197 106 198 
<< pdiffusion >>
rect 106 197 107 198 
<< pdiffusion >>
rect 107 197 108 198 
<< m1 >>
rect 118 197 119 198 
<< pdiffusion >>
rect 120 197 121 198 
<< pdiffusion >>
rect 121 197 122 198 
<< pdiffusion >>
rect 122 197 123 198 
<< pdiffusion >>
rect 123 197 124 198 
<< pdiffusion >>
rect 124 197 125 198 
<< pdiffusion >>
rect 125 197 126 198 
<< m1 >>
rect 127 197 128 198 
<< m2 >>
rect 127 197 128 198 
<< pdiffusion >>
rect 138 197 139 198 
<< pdiffusion >>
rect 139 197 140 198 
<< pdiffusion >>
rect 140 197 141 198 
<< pdiffusion >>
rect 141 197 142 198 
<< pdiffusion >>
rect 142 197 143 198 
<< pdiffusion >>
rect 143 197 144 198 
<< m1 >>
rect 154 197 155 198 
<< pdiffusion >>
rect 156 197 157 198 
<< pdiffusion >>
rect 157 197 158 198 
<< pdiffusion >>
rect 158 197 159 198 
<< pdiffusion >>
rect 159 197 160 198 
<< pdiffusion >>
rect 160 197 161 198 
<< pdiffusion >>
rect 161 197 162 198 
<< m1 >>
rect 172 197 173 198 
<< pdiffusion >>
rect 174 197 175 198 
<< pdiffusion >>
rect 175 197 176 198 
<< pdiffusion >>
rect 176 197 177 198 
<< pdiffusion >>
rect 177 197 178 198 
<< pdiffusion >>
rect 178 197 179 198 
<< pdiffusion >>
rect 179 197 180 198 
<< m1 >>
rect 181 197 182 198 
<< m2 >>
rect 181 197 182 198 
<< pdiffusion >>
rect 192 197 193 198 
<< pdiffusion >>
rect 193 197 194 198 
<< pdiffusion >>
rect 194 197 195 198 
<< pdiffusion >>
rect 195 197 196 198 
<< pdiffusion >>
rect 196 197 197 198 
<< pdiffusion >>
rect 197 197 198 198 
<< pdiffusion >>
rect 210 197 211 198 
<< m1 >>
rect 211 197 212 198 
<< pdiffusion >>
rect 211 197 212 198 
<< pdiffusion >>
rect 212 197 213 198 
<< pdiffusion >>
rect 213 197 214 198 
<< m1 >>
rect 214 197 215 198 
<< pdiffusion >>
rect 214 197 215 198 
<< pdiffusion >>
rect 215 197 216 198 
<< m1 >>
rect 217 197 218 198 
<< m2 >>
rect 217 197 218 198 
<< m2c >>
rect 217 197 218 198 
<< m1 >>
rect 217 197 218 198 
<< m2 >>
rect 217 197 218 198 
<< m1 >>
rect 226 197 227 198 
<< pdiffusion >>
rect 228 197 229 198 
<< pdiffusion >>
rect 229 197 230 198 
<< pdiffusion >>
rect 230 197 231 198 
<< pdiffusion >>
rect 231 197 232 198 
<< pdiffusion >>
rect 232 197 233 198 
<< pdiffusion >>
rect 233 197 234 198 
<< m1 >>
rect 235 197 236 198 
<< pdiffusion >>
rect 246 197 247 198 
<< pdiffusion >>
rect 247 197 248 198 
<< pdiffusion >>
rect 248 197 249 198 
<< pdiffusion >>
rect 249 197 250 198 
<< pdiffusion >>
rect 250 197 251 198 
<< pdiffusion >>
rect 251 197 252 198 
<< m1 >>
rect 254 197 255 198 
<< pdiffusion >>
rect 264 197 265 198 
<< m1 >>
rect 265 197 266 198 
<< pdiffusion >>
rect 265 197 266 198 
<< pdiffusion >>
rect 266 197 267 198 
<< pdiffusion >>
rect 267 197 268 198 
<< m1 >>
rect 268 197 269 198 
<< pdiffusion >>
rect 268 197 269 198 
<< pdiffusion >>
rect 269 197 270 198 
<< pdiffusion >>
rect 282 197 283 198 
<< pdiffusion >>
rect 283 197 284 198 
<< pdiffusion >>
rect 284 197 285 198 
<< pdiffusion >>
rect 285 197 286 198 
<< m1 >>
rect 286 197 287 198 
<< pdiffusion >>
rect 286 197 287 198 
<< pdiffusion >>
rect 287 197 288 198 
<< m1 >>
rect 298 197 299 198 
<< pdiffusion >>
rect 300 197 301 198 
<< pdiffusion >>
rect 301 197 302 198 
<< pdiffusion >>
rect 302 197 303 198 
<< pdiffusion >>
rect 303 197 304 198 
<< pdiffusion >>
rect 304 197 305 198 
<< pdiffusion >>
rect 305 197 306 198 
<< m1 >>
rect 307 197 308 198 
<< m2 >>
rect 308 197 309 198 
<< m1 >>
rect 311 197 312 198 
<< m1 >>
rect 313 197 314 198 
<< pdiffusion >>
rect 318 197 319 198 
<< pdiffusion >>
rect 319 197 320 198 
<< pdiffusion >>
rect 320 197 321 198 
<< pdiffusion >>
rect 321 197 322 198 
<< pdiffusion >>
rect 322 197 323 198 
<< pdiffusion >>
rect 323 197 324 198 
<< pdiffusion >>
rect 336 197 337 198 
<< pdiffusion >>
rect 337 197 338 198 
<< pdiffusion >>
rect 338 197 339 198 
<< pdiffusion >>
rect 339 197 340 198 
<< pdiffusion >>
rect 340 197 341 198 
<< pdiffusion >>
rect 341 197 342 198 
<< m1 >>
rect 343 197 344 198 
<< pdiffusion >>
rect 354 197 355 198 
<< pdiffusion >>
rect 355 197 356 198 
<< pdiffusion >>
rect 356 197 357 198 
<< pdiffusion >>
rect 357 197 358 198 
<< pdiffusion >>
rect 358 197 359 198 
<< pdiffusion >>
rect 359 197 360 198 
<< pdiffusion >>
rect 372 197 373 198 
<< pdiffusion >>
rect 373 197 374 198 
<< pdiffusion >>
rect 374 197 375 198 
<< pdiffusion >>
rect 375 197 376 198 
<< pdiffusion >>
rect 376 197 377 198 
<< pdiffusion >>
rect 377 197 378 198 
<< pdiffusion >>
rect 390 197 391 198 
<< pdiffusion >>
rect 391 197 392 198 
<< pdiffusion >>
rect 392 197 393 198 
<< pdiffusion >>
rect 393 197 394 198 
<< pdiffusion >>
rect 394 197 395 198 
<< pdiffusion >>
rect 395 197 396 198 
<< pdiffusion >>
rect 408 197 409 198 
<< pdiffusion >>
rect 409 197 410 198 
<< pdiffusion >>
rect 410 197 411 198 
<< pdiffusion >>
rect 411 197 412 198 
<< pdiffusion >>
rect 412 197 413 198 
<< pdiffusion >>
rect 413 197 414 198 
<< pdiffusion >>
rect 426 197 427 198 
<< pdiffusion >>
rect 427 197 428 198 
<< pdiffusion >>
rect 428 197 429 198 
<< pdiffusion >>
rect 429 197 430 198 
<< pdiffusion >>
rect 430 197 431 198 
<< pdiffusion >>
rect 431 197 432 198 
<< pdiffusion >>
rect 444 197 445 198 
<< pdiffusion >>
rect 445 197 446 198 
<< pdiffusion >>
rect 446 197 447 198 
<< pdiffusion >>
rect 447 197 448 198 
<< pdiffusion >>
rect 448 197 449 198 
<< pdiffusion >>
rect 449 197 450 198 
<< m1 >>
rect 16 198 17 199 
<< m1 >>
rect 19 198 20 199 
<< m1 >>
rect 49 198 50 199 
<< m1 >>
rect 93 198 94 199 
<< m1 >>
rect 118 198 119 199 
<< m1 >>
rect 127 198 128 199 
<< m2 >>
rect 127 198 128 199 
<< m1 >>
rect 154 198 155 199 
<< m1 >>
rect 172 198 173 199 
<< m1 >>
rect 181 198 182 199 
<< m2 >>
rect 181 198 182 199 
<< m1 >>
rect 211 198 212 199 
<< m1 >>
rect 214 198 215 199 
<< m2 >>
rect 217 198 218 199 
<< m1 >>
rect 226 198 227 199 
<< m1 >>
rect 235 198 236 199 
<< m1 >>
rect 254 198 255 199 
<< m1 >>
rect 265 198 266 199 
<< m1 >>
rect 268 198 269 199 
<< m1 >>
rect 286 198 287 199 
<< m1 >>
rect 298 198 299 199 
<< m1 >>
rect 307 198 308 199 
<< m2 >>
rect 308 198 309 199 
<< m1 >>
rect 311 198 312 199 
<< m1 >>
rect 313 198 314 199 
<< m1 >>
rect 343 198 344 199 
<< m1 >>
rect 16 199 17 200 
<< m1 >>
rect 19 199 20 200 
<< m1 >>
rect 49 199 50 200 
<< m1 >>
rect 93 199 94 200 
<< m1 >>
rect 118 199 119 200 
<< m1 >>
rect 127 199 128 200 
<< m2 >>
rect 127 199 128 200 
<< m1 >>
rect 154 199 155 200 
<< m1 >>
rect 172 199 173 200 
<< m1 >>
rect 181 199 182 200 
<< m2 >>
rect 181 199 182 200 
<< m1 >>
rect 211 199 212 200 
<< m1 >>
rect 214 199 215 200 
<< m1 >>
rect 215 199 216 200 
<< m1 >>
rect 216 199 217 200 
<< m1 >>
rect 217 199 218 200 
<< m2 >>
rect 217 199 218 200 
<< m1 >>
rect 218 199 219 200 
<< m1 >>
rect 219 199 220 200 
<< m1 >>
rect 220 199 221 200 
<< m1 >>
rect 221 199 222 200 
<< m1 >>
rect 222 199 223 200 
<< m1 >>
rect 223 199 224 200 
<< m1 >>
rect 224 199 225 200 
<< m1 >>
rect 225 199 226 200 
<< m1 >>
rect 226 199 227 200 
<< m1 >>
rect 235 199 236 200 
<< m1 >>
rect 254 199 255 200 
<< m1 >>
rect 265 199 266 200 
<< m1 >>
rect 266 199 267 200 
<< m2 >>
rect 266 199 267 200 
<< m2c >>
rect 266 199 267 200 
<< m1 >>
rect 266 199 267 200 
<< m2 >>
rect 266 199 267 200 
<< m2 >>
rect 267 199 268 200 
<< m1 >>
rect 268 199 269 200 
<< m1 >>
rect 286 199 287 200 
<< m1 >>
rect 298 199 299 200 
<< m1 >>
rect 307 199 308 200 
<< m2 >>
rect 308 199 309 200 
<< m1 >>
rect 311 199 312 200 
<< m1 >>
rect 313 199 314 200 
<< m1 >>
rect 343 199 344 200 
<< m1 >>
rect 16 200 17 201 
<< m1 >>
rect 19 200 20 201 
<< m1 >>
rect 49 200 50 201 
<< m1 >>
rect 93 200 94 201 
<< m1 >>
rect 118 200 119 201 
<< m1 >>
rect 127 200 128 201 
<< m2 >>
rect 127 200 128 201 
<< m1 >>
rect 154 200 155 201 
<< m1 >>
rect 172 200 173 201 
<< m1 >>
rect 181 200 182 201 
<< m2 >>
rect 181 200 182 201 
<< m1 >>
rect 200 200 201 201 
<< m2 >>
rect 200 200 201 201 
<< m2c >>
rect 200 200 201 201 
<< m1 >>
rect 200 200 201 201 
<< m2 >>
rect 200 200 201 201 
<< m1 >>
rect 201 200 202 201 
<< m1 >>
rect 202 200 203 201 
<< m1 >>
rect 203 200 204 201 
<< m1 >>
rect 204 200 205 201 
<< m1 >>
rect 205 200 206 201 
<< m1 >>
rect 206 200 207 201 
<< m1 >>
rect 207 200 208 201 
<< m1 >>
rect 208 200 209 201 
<< m1 >>
rect 209 200 210 201 
<< m1 >>
rect 210 200 211 201 
<< m1 >>
rect 211 200 212 201 
<< m2 >>
rect 217 200 218 201 
<< m1 >>
rect 235 200 236 201 
<< m2 >>
rect 235 200 236 201 
<< m2c >>
rect 235 200 236 201 
<< m1 >>
rect 235 200 236 201 
<< m2 >>
rect 235 200 236 201 
<< m1 >>
rect 254 200 255 201 
<< m2 >>
rect 254 200 255 201 
<< m2c >>
rect 254 200 255 201 
<< m1 >>
rect 254 200 255 201 
<< m2 >>
rect 254 200 255 201 
<< m2 >>
rect 267 200 268 201 
<< m1 >>
rect 268 200 269 201 
<< m2 >>
rect 268 200 269 201 
<< m2 >>
rect 269 200 270 201 
<< m1 >>
rect 270 200 271 201 
<< m2 >>
rect 270 200 271 201 
<< m2c >>
rect 270 200 271 201 
<< m1 >>
rect 270 200 271 201 
<< m2 >>
rect 270 200 271 201 
<< m1 >>
rect 286 200 287 201 
<< m1 >>
rect 298 200 299 201 
<< m1 >>
rect 307 200 308 201 
<< m2 >>
rect 308 200 309 201 
<< m1 >>
rect 311 200 312 201 
<< m1 >>
rect 313 200 314 201 
<< m1 >>
rect 343 200 344 201 
<< m1 >>
rect 16 201 17 202 
<< m1 >>
rect 19 201 20 202 
<< m1 >>
rect 49 201 50 202 
<< m1 >>
rect 93 201 94 202 
<< m1 >>
rect 118 201 119 202 
<< m1 >>
rect 127 201 128 202 
<< m2 >>
rect 127 201 128 202 
<< m1 >>
rect 154 201 155 202 
<< m1 >>
rect 172 201 173 202 
<< m1 >>
rect 181 201 182 202 
<< m2 >>
rect 181 201 182 202 
<< m2 >>
rect 200 201 201 202 
<< m2 >>
rect 217 201 218 202 
<< m2 >>
rect 235 201 236 202 
<< m2 >>
rect 254 201 255 202 
<< m1 >>
rect 268 201 269 202 
<< m1 >>
rect 270 201 271 202 
<< m1 >>
rect 286 201 287 202 
<< m1 >>
rect 298 201 299 202 
<< m1 >>
rect 307 201 308 202 
<< m2 >>
rect 308 201 309 202 
<< m1 >>
rect 311 201 312 202 
<< m1 >>
rect 313 201 314 202 
<< m1 >>
rect 343 201 344 202 
<< m1 >>
rect 16 202 17 203 
<< m1 >>
rect 19 202 20 203 
<< m1 >>
rect 49 202 50 203 
<< m1 >>
rect 93 202 94 203 
<< m2 >>
rect 93 202 94 203 
<< m2c >>
rect 93 202 94 203 
<< m1 >>
rect 93 202 94 203 
<< m2 >>
rect 93 202 94 203 
<< m1 >>
rect 118 202 119 203 
<< m2 >>
rect 118 202 119 203 
<< m2c >>
rect 118 202 119 203 
<< m1 >>
rect 118 202 119 203 
<< m2 >>
rect 118 202 119 203 
<< m1 >>
rect 121 202 122 203 
<< m2 >>
rect 121 202 122 203 
<< m2c >>
rect 121 202 122 203 
<< m1 >>
rect 121 202 122 203 
<< m2 >>
rect 121 202 122 203 
<< m1 >>
rect 122 202 123 203 
<< m1 >>
rect 123 202 124 203 
<< m1 >>
rect 124 202 125 203 
<< m1 >>
rect 125 202 126 203 
<< m1 >>
rect 126 202 127 203 
<< m1 >>
rect 127 202 128 203 
<< m2 >>
rect 127 202 128 203 
<< m1 >>
rect 154 202 155 203 
<< m2 >>
rect 154 202 155 203 
<< m2c >>
rect 154 202 155 203 
<< m1 >>
rect 154 202 155 203 
<< m2 >>
rect 154 202 155 203 
<< m1 >>
rect 172 202 173 203 
<< m1 >>
rect 173 202 174 203 
<< m1 >>
rect 174 202 175 203 
<< m1 >>
rect 175 202 176 203 
<< m1 >>
rect 176 202 177 203 
<< m1 >>
rect 177 202 178 203 
<< m1 >>
rect 178 202 179 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m2c >>
rect 179 202 180 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m1 >>
rect 181 202 182 203 
<< m2 >>
rect 181 202 182 203 
<< m1 >>
rect 182 202 183 203 
<< m1 >>
rect 183 202 184 203 
<< m1 >>
rect 184 202 185 203 
<< m1 >>
rect 185 202 186 203 
<< m1 >>
rect 186 202 187 203 
<< m1 >>
rect 187 202 188 203 
<< m1 >>
rect 188 202 189 203 
<< m1 >>
rect 189 202 190 203 
<< m1 >>
rect 190 202 191 203 
<< m1 >>
rect 191 202 192 203 
<< m1 >>
rect 192 202 193 203 
<< m1 >>
rect 193 202 194 203 
<< m1 >>
rect 194 202 195 203 
<< m1 >>
rect 195 202 196 203 
<< m1 >>
rect 196 202 197 203 
<< m1 >>
rect 197 202 198 203 
<< m1 >>
rect 198 202 199 203 
<< m1 >>
rect 199 202 200 203 
<< m1 >>
rect 200 202 201 203 
<< m2 >>
rect 200 202 201 203 
<< m1 >>
rect 201 202 202 203 
<< m1 >>
rect 202 202 203 203 
<< m1 >>
rect 203 202 204 203 
<< m1 >>
rect 204 202 205 203 
<< m1 >>
rect 205 202 206 203 
<< m1 >>
rect 206 202 207 203 
<< m1 >>
rect 207 202 208 203 
<< m1 >>
rect 208 202 209 203 
<< m1 >>
rect 209 202 210 203 
<< m1 >>
rect 210 202 211 203 
<< m1 >>
rect 211 202 212 203 
<< m1 >>
rect 212 202 213 203 
<< m1 >>
rect 213 202 214 203 
<< m1 >>
rect 214 202 215 203 
<< m1 >>
rect 215 202 216 203 
<< m1 >>
rect 216 202 217 203 
<< m1 >>
rect 217 202 218 203 
<< m2 >>
rect 217 202 218 203 
<< m1 >>
rect 218 202 219 203 
<< m1 >>
rect 219 202 220 203 
<< m1 >>
rect 220 202 221 203 
<< m1 >>
rect 221 202 222 203 
<< m1 >>
rect 222 202 223 203 
<< m1 >>
rect 223 202 224 203 
<< m1 >>
rect 224 202 225 203 
<< m1 >>
rect 225 202 226 203 
<< m1 >>
rect 226 202 227 203 
<< m1 >>
rect 227 202 228 203 
<< m1 >>
rect 228 202 229 203 
<< m1 >>
rect 229 202 230 203 
<< m1 >>
rect 230 202 231 203 
<< m1 >>
rect 231 202 232 203 
<< m1 >>
rect 232 202 233 203 
<< m1 >>
rect 233 202 234 203 
<< m1 >>
rect 234 202 235 203 
<< m1 >>
rect 235 202 236 203 
<< m2 >>
rect 235 202 236 203 
<< m1 >>
rect 236 202 237 203 
<< m1 >>
rect 237 202 238 203 
<< m1 >>
rect 238 202 239 203 
<< m1 >>
rect 239 202 240 203 
<< m1 >>
rect 240 202 241 203 
<< m1 >>
rect 241 202 242 203 
<< m1 >>
rect 242 202 243 203 
<< m1 >>
rect 243 202 244 203 
<< m1 >>
rect 244 202 245 203 
<< m1 >>
rect 245 202 246 203 
<< m1 >>
rect 246 202 247 203 
<< m1 >>
rect 247 202 248 203 
<< m1 >>
rect 248 202 249 203 
<< m1 >>
rect 249 202 250 203 
<< m1 >>
rect 250 202 251 203 
<< m2 >>
rect 251 202 252 203 
<< m1 >>
rect 252 202 253 203 
<< m2 >>
rect 252 202 253 203 
<< m2c >>
rect 252 202 253 203 
<< m1 >>
rect 252 202 253 203 
<< m2 >>
rect 252 202 253 203 
<< m1 >>
rect 253 202 254 203 
<< m1 >>
rect 254 202 255 203 
<< m2 >>
rect 254 202 255 203 
<< m1 >>
rect 255 202 256 203 
<< m1 >>
rect 256 202 257 203 
<< m1 >>
rect 257 202 258 203 
<< m1 >>
rect 258 202 259 203 
<< m1 >>
rect 259 202 260 203 
<< m1 >>
rect 260 202 261 203 
<< m1 >>
rect 261 202 262 203 
<< m1 >>
rect 262 202 263 203 
<< m1 >>
rect 263 202 264 203 
<< m1 >>
rect 264 202 265 203 
<< m1 >>
rect 265 202 266 203 
<< m1 >>
rect 266 202 267 203 
<< m1 >>
rect 267 202 268 203 
<< m1 >>
rect 268 202 269 203 
<< m1 >>
rect 270 202 271 203 
<< m1 >>
rect 271 202 272 203 
<< m1 >>
rect 272 202 273 203 
<< m1 >>
rect 273 202 274 203 
<< m1 >>
rect 274 202 275 203 
<< m1 >>
rect 275 202 276 203 
<< m1 >>
rect 276 202 277 203 
<< m1 >>
rect 277 202 278 203 
<< m1 >>
rect 278 202 279 203 
<< m1 >>
rect 279 202 280 203 
<< m1 >>
rect 280 202 281 203 
<< m1 >>
rect 281 202 282 203 
<< m1 >>
rect 282 202 283 203 
<< m1 >>
rect 283 202 284 203 
<< m1 >>
rect 284 202 285 203 
<< m2 >>
rect 284 202 285 203 
<< m2c >>
rect 284 202 285 203 
<< m1 >>
rect 284 202 285 203 
<< m2 >>
rect 284 202 285 203 
<< m2 >>
rect 285 202 286 203 
<< m1 >>
rect 286 202 287 203 
<< m1 >>
rect 298 202 299 203 
<< m1 >>
rect 307 202 308 203 
<< m2 >>
rect 308 202 309 203 
<< m1 >>
rect 311 202 312 203 
<< m1 >>
rect 313 202 314 203 
<< m1 >>
rect 314 202 315 203 
<< m1 >>
rect 315 202 316 203 
<< m1 >>
rect 316 202 317 203 
<< m1 >>
rect 317 202 318 203 
<< m1 >>
rect 318 202 319 203 
<< m1 >>
rect 319 202 320 203 
<< m1 >>
rect 320 202 321 203 
<< m1 >>
rect 321 202 322 203 
<< m1 >>
rect 322 202 323 203 
<< m1 >>
rect 323 202 324 203 
<< m1 >>
rect 324 202 325 203 
<< m1 >>
rect 325 202 326 203 
<< m1 >>
rect 326 202 327 203 
<< m1 >>
rect 327 202 328 203 
<< m1 >>
rect 328 202 329 203 
<< m1 >>
rect 329 202 330 203 
<< m1 >>
rect 330 202 331 203 
<< m1 >>
rect 331 202 332 203 
<< m1 >>
rect 332 202 333 203 
<< m1 >>
rect 333 202 334 203 
<< m1 >>
rect 334 202 335 203 
<< m1 >>
rect 335 202 336 203 
<< m1 >>
rect 336 202 337 203 
<< m1 >>
rect 337 202 338 203 
<< m1 >>
rect 343 202 344 203 
<< m1 >>
rect 16 203 17 204 
<< m1 >>
rect 19 203 20 204 
<< m1 >>
rect 49 203 50 204 
<< m2 >>
rect 93 203 94 204 
<< m2 >>
rect 118 203 119 204 
<< m2 >>
rect 121 203 122 204 
<< m2 >>
rect 127 203 128 204 
<< m2 >>
rect 154 203 155 204 
<< m2 >>
rect 179 203 180 204 
<< m2 >>
rect 181 203 182 204 
<< m2 >>
rect 200 203 201 204 
<< m2 >>
rect 217 203 218 204 
<< m2 >>
rect 235 203 236 204 
<< m1 >>
rect 250 203 251 204 
<< m2 >>
rect 251 203 252 204 
<< m2 >>
rect 254 203 255 204 
<< m2 >>
rect 285 203 286 204 
<< m1 >>
rect 286 203 287 204 
<< m1 >>
rect 298 203 299 204 
<< m1 >>
rect 307 203 308 204 
<< m2 >>
rect 308 203 309 204 
<< m1 >>
rect 311 203 312 204 
<< m1 >>
rect 337 203 338 204 
<< m1 >>
rect 343 203 344 204 
<< m1 >>
rect 16 204 17 205 
<< m1 >>
rect 19 204 20 205 
<< m1 >>
rect 49 204 50 205 
<< m1 >>
rect 50 204 51 205 
<< m1 >>
rect 51 204 52 205 
<< m1 >>
rect 52 204 53 205 
<< m1 >>
rect 53 204 54 205 
<< m1 >>
rect 54 204 55 205 
<< m1 >>
rect 55 204 56 205 
<< m1 >>
rect 56 204 57 205 
<< m1 >>
rect 57 204 58 205 
<< m1 >>
rect 58 204 59 205 
<< m1 >>
rect 59 204 60 205 
<< m1 >>
rect 60 204 61 205 
<< m1 >>
rect 61 204 62 205 
<< m1 >>
rect 62 204 63 205 
<< m1 >>
rect 63 204 64 205 
<< m1 >>
rect 64 204 65 205 
<< m1 >>
rect 65 204 66 205 
<< m1 >>
rect 66 204 67 205 
<< m1 >>
rect 67 204 68 205 
<< m1 >>
rect 68 204 69 205 
<< m1 >>
rect 69 204 70 205 
<< m1 >>
rect 70 204 71 205 
<< m1 >>
rect 71 204 72 205 
<< m1 >>
rect 72 204 73 205 
<< m1 >>
rect 73 204 74 205 
<< m1 >>
rect 74 204 75 205 
<< m1 >>
rect 75 204 76 205 
<< m1 >>
rect 76 204 77 205 
<< m1 >>
rect 77 204 78 205 
<< m1 >>
rect 78 204 79 205 
<< m1 >>
rect 79 204 80 205 
<< m1 >>
rect 80 204 81 205 
<< m1 >>
rect 81 204 82 205 
<< m1 >>
rect 82 204 83 205 
<< m1 >>
rect 83 204 84 205 
<< m1 >>
rect 84 204 85 205 
<< m1 >>
rect 85 204 86 205 
<< m1 >>
rect 86 204 87 205 
<< m1 >>
rect 87 204 88 205 
<< m1 >>
rect 88 204 89 205 
<< m1 >>
rect 89 204 90 205 
<< m1 >>
rect 90 204 91 205 
<< m1 >>
rect 91 204 92 205 
<< m1 >>
rect 92 204 93 205 
<< m1 >>
rect 93 204 94 205 
<< m2 >>
rect 93 204 94 205 
<< m1 >>
rect 94 204 95 205 
<< m1 >>
rect 95 204 96 205 
<< m1 >>
rect 96 204 97 205 
<< m1 >>
rect 97 204 98 205 
<< m1 >>
rect 98 204 99 205 
<< m1 >>
rect 99 204 100 205 
<< m1 >>
rect 100 204 101 205 
<< m1 >>
rect 101 204 102 205 
<< m1 >>
rect 102 204 103 205 
<< m1 >>
rect 103 204 104 205 
<< m1 >>
rect 104 204 105 205 
<< m1 >>
rect 105 204 106 205 
<< m1 >>
rect 106 204 107 205 
<< m1 >>
rect 107 204 108 205 
<< m1 >>
rect 108 204 109 205 
<< m1 >>
rect 109 204 110 205 
<< m1 >>
rect 110 204 111 205 
<< m1 >>
rect 111 204 112 205 
<< m1 >>
rect 112 204 113 205 
<< m1 >>
rect 113 204 114 205 
<< m1 >>
rect 114 204 115 205 
<< m1 >>
rect 115 204 116 205 
<< m1 >>
rect 116 204 117 205 
<< m1 >>
rect 117 204 118 205 
<< m1 >>
rect 118 204 119 205 
<< m2 >>
rect 118 204 119 205 
<< m1 >>
rect 119 204 120 205 
<< m1 >>
rect 120 204 121 205 
<< m1 >>
rect 121 204 122 205 
<< m2 >>
rect 121 204 122 205 
<< m1 >>
rect 122 204 123 205 
<< m1 >>
rect 123 204 124 205 
<< m1 >>
rect 124 204 125 205 
<< m1 >>
rect 125 204 126 205 
<< m1 >>
rect 126 204 127 205 
<< m1 >>
rect 127 204 128 205 
<< m2 >>
rect 127 204 128 205 
<< m1 >>
rect 128 204 129 205 
<< m1 >>
rect 129 204 130 205 
<< m1 >>
rect 130 204 131 205 
<< m1 >>
rect 131 204 132 205 
<< m1 >>
rect 132 204 133 205 
<< m1 >>
rect 133 204 134 205 
<< m1 >>
rect 134 204 135 205 
<< m1 >>
rect 135 204 136 205 
<< m1 >>
rect 136 204 137 205 
<< m1 >>
rect 137 204 138 205 
<< m1 >>
rect 138 204 139 205 
<< m1 >>
rect 139 204 140 205 
<< m1 >>
rect 140 204 141 205 
<< m1 >>
rect 141 204 142 205 
<< m1 >>
rect 142 204 143 205 
<< m1 >>
rect 143 204 144 205 
<< m1 >>
rect 144 204 145 205 
<< m1 >>
rect 145 204 146 205 
<< m1 >>
rect 146 204 147 205 
<< m1 >>
rect 147 204 148 205 
<< m1 >>
rect 148 204 149 205 
<< m1 >>
rect 149 204 150 205 
<< m1 >>
rect 150 204 151 205 
<< m1 >>
rect 151 204 152 205 
<< m1 >>
rect 152 204 153 205 
<< m1 >>
rect 153 204 154 205 
<< m1 >>
rect 154 204 155 205 
<< m2 >>
rect 154 204 155 205 
<< m1 >>
rect 155 204 156 205 
<< m1 >>
rect 156 204 157 205 
<< m1 >>
rect 157 204 158 205 
<< m1 >>
rect 158 204 159 205 
<< m1 >>
rect 159 204 160 205 
<< m1 >>
rect 160 204 161 205 
<< m1 >>
rect 161 204 162 205 
<< m1 >>
rect 162 204 163 205 
<< m1 >>
rect 163 204 164 205 
<< m1 >>
rect 164 204 165 205 
<< m1 >>
rect 165 204 166 205 
<< m1 >>
rect 166 204 167 205 
<< m1 >>
rect 167 204 168 205 
<< m1 >>
rect 168 204 169 205 
<< m1 >>
rect 169 204 170 205 
<< m1 >>
rect 170 204 171 205 
<< m1 >>
rect 171 204 172 205 
<< m1 >>
rect 172 204 173 205 
<< m1 >>
rect 173 204 174 205 
<< m1 >>
rect 174 204 175 205 
<< m1 >>
rect 175 204 176 205 
<< m1 >>
rect 176 204 177 205 
<< m1 >>
rect 177 204 178 205 
<< m1 >>
rect 178 204 179 205 
<< m1 >>
rect 179 204 180 205 
<< m2 >>
rect 179 204 180 205 
<< m1 >>
rect 180 204 181 205 
<< m1 >>
rect 181 204 182 205 
<< m2 >>
rect 181 204 182 205 
<< m1 >>
rect 182 204 183 205 
<< m2 >>
rect 182 204 183 205 
<< m1 >>
rect 183 204 184 205 
<< m2 >>
rect 183 204 184 205 
<< m1 >>
rect 184 204 185 205 
<< m2 >>
rect 184 204 185 205 
<< m1 >>
rect 185 204 186 205 
<< m2 >>
rect 185 204 186 205 
<< m1 >>
rect 186 204 187 205 
<< m2 >>
rect 186 204 187 205 
<< m1 >>
rect 187 204 188 205 
<< m2 >>
rect 187 204 188 205 
<< m1 >>
rect 188 204 189 205 
<< m2 >>
rect 188 204 189 205 
<< m1 >>
rect 189 204 190 205 
<< m2 >>
rect 189 204 190 205 
<< m1 >>
rect 190 204 191 205 
<< m2 >>
rect 190 204 191 205 
<< m1 >>
rect 191 204 192 205 
<< m2 >>
rect 191 204 192 205 
<< m1 >>
rect 192 204 193 205 
<< m2 >>
rect 192 204 193 205 
<< m1 >>
rect 193 204 194 205 
<< m2 >>
rect 193 204 194 205 
<< m1 >>
rect 194 204 195 205 
<< m2 >>
rect 194 204 195 205 
<< m1 >>
rect 195 204 196 205 
<< m2 >>
rect 195 204 196 205 
<< m1 >>
rect 196 204 197 205 
<< m2 >>
rect 196 204 197 205 
<< m2 >>
rect 197 204 198 205 
<< m1 >>
rect 198 204 199 205 
<< m2 >>
rect 198 204 199 205 
<< m2c >>
rect 198 204 199 205 
<< m1 >>
rect 198 204 199 205 
<< m2 >>
rect 198 204 199 205 
<< m1 >>
rect 199 204 200 205 
<< m1 >>
rect 200 204 201 205 
<< m2 >>
rect 200 204 201 205 
<< m1 >>
rect 201 204 202 205 
<< m1 >>
rect 202 204 203 205 
<< m1 >>
rect 203 204 204 205 
<< m1 >>
rect 204 204 205 205 
<< m1 >>
rect 205 204 206 205 
<< m1 >>
rect 206 204 207 205 
<< m1 >>
rect 207 204 208 205 
<< m1 >>
rect 217 204 218 205 
<< m2 >>
rect 217 204 218 205 
<< m2c >>
rect 217 204 218 205 
<< m1 >>
rect 217 204 218 205 
<< m2 >>
rect 217 204 218 205 
<< m1 >>
rect 235 204 236 205 
<< m2 >>
rect 235 204 236 205 
<< m2c >>
rect 235 204 236 205 
<< m1 >>
rect 235 204 236 205 
<< m2 >>
rect 235 204 236 205 
<< m1 >>
rect 244 204 245 205 
<< m1 >>
rect 245 204 246 205 
<< m1 >>
rect 246 204 247 205 
<< m1 >>
rect 247 204 248 205 
<< m1 >>
rect 248 204 249 205 
<< m2 >>
rect 248 204 249 205 
<< m2c >>
rect 248 204 249 205 
<< m1 >>
rect 248 204 249 205 
<< m2 >>
rect 248 204 249 205 
<< m2 >>
rect 249 204 250 205 
<< m1 >>
rect 250 204 251 205 
<< m2 >>
rect 250 204 251 205 
<< m2 >>
rect 251 204 252 205 
<< m1 >>
rect 254 204 255 205 
<< m2 >>
rect 254 204 255 205 
<< m2c >>
rect 254 204 255 205 
<< m1 >>
rect 254 204 255 205 
<< m2 >>
rect 254 204 255 205 
<< m2 >>
rect 285 204 286 205 
<< m1 >>
rect 286 204 287 205 
<< m1 >>
rect 298 204 299 205 
<< m1 >>
rect 307 204 308 205 
<< m2 >>
rect 308 204 309 205 
<< m1 >>
rect 311 204 312 205 
<< m1 >>
rect 337 204 338 205 
<< m1 >>
rect 343 204 344 205 
<< m1 >>
rect 16 205 17 206 
<< m1 >>
rect 19 205 20 206 
<< m2 >>
rect 93 205 94 206 
<< m2 >>
rect 118 205 119 206 
<< m2 >>
rect 121 205 122 206 
<< m2 >>
rect 127 205 128 206 
<< m2 >>
rect 154 205 155 206 
<< m2 >>
rect 179 205 180 206 
<< m1 >>
rect 196 205 197 206 
<< m2 >>
rect 200 205 201 206 
<< m1 >>
rect 207 205 208 206 
<< m1 >>
rect 217 205 218 206 
<< m1 >>
rect 235 205 236 206 
<< m1 >>
rect 244 205 245 206 
<< m1 >>
rect 250 205 251 206 
<< m1 >>
rect 254 205 255 206 
<< m2 >>
rect 285 205 286 206 
<< m1 >>
rect 286 205 287 206 
<< m1 >>
rect 298 205 299 206 
<< m2 >>
rect 298 205 299 206 
<< m2c >>
rect 298 205 299 206 
<< m1 >>
rect 298 205 299 206 
<< m2 >>
rect 298 205 299 206 
<< m1 >>
rect 307 205 308 206 
<< m2 >>
rect 308 205 309 206 
<< m1 >>
rect 311 205 312 206 
<< m1 >>
rect 337 205 338 206 
<< m1 >>
rect 343 205 344 206 
<< m1 >>
rect 16 206 17 207 
<< m1 >>
rect 19 206 20 207 
<< m1 >>
rect 93 206 94 207 
<< m2 >>
rect 93 206 94 207 
<< m2c >>
rect 93 206 94 207 
<< m1 >>
rect 93 206 94 207 
<< m2 >>
rect 93 206 94 207 
<< m1 >>
rect 118 206 119 207 
<< m2 >>
rect 118 206 119 207 
<< m2c >>
rect 118 206 119 207 
<< m1 >>
rect 118 206 119 207 
<< m2 >>
rect 118 206 119 207 
<< m1 >>
rect 121 206 122 207 
<< m2 >>
rect 121 206 122 207 
<< m2c >>
rect 121 206 122 207 
<< m1 >>
rect 121 206 122 207 
<< m2 >>
rect 121 206 122 207 
<< m1 >>
rect 127 206 128 207 
<< m2 >>
rect 127 206 128 207 
<< m2c >>
rect 127 206 128 207 
<< m1 >>
rect 127 206 128 207 
<< m2 >>
rect 127 206 128 207 
<< m1 >>
rect 154 206 155 207 
<< m2 >>
rect 154 206 155 207 
<< m2c >>
rect 154 206 155 207 
<< m1 >>
rect 154 206 155 207 
<< m2 >>
rect 154 206 155 207 
<< m1 >>
rect 179 206 180 207 
<< m2 >>
rect 179 206 180 207 
<< m2c >>
rect 179 206 180 207 
<< m1 >>
rect 179 206 180 207 
<< m2 >>
rect 179 206 180 207 
<< m1 >>
rect 196 206 197 207 
<< m1 >>
rect 200 206 201 207 
<< m2 >>
rect 200 206 201 207 
<< m2c >>
rect 200 206 201 207 
<< m1 >>
rect 200 206 201 207 
<< m2 >>
rect 200 206 201 207 
<< m1 >>
rect 207 206 208 207 
<< m1 >>
rect 217 206 218 207 
<< m1 >>
rect 218 206 219 207 
<< m1 >>
rect 219 206 220 207 
<< m1 >>
rect 220 206 221 207 
<< m1 >>
rect 221 206 222 207 
<< m1 >>
rect 222 206 223 207 
<< m1 >>
rect 223 206 224 207 
<< m1 >>
rect 224 206 225 207 
<< m1 >>
rect 225 206 226 207 
<< m1 >>
rect 226 206 227 207 
<< m1 >>
rect 227 206 228 207 
<< m1 >>
rect 228 206 229 207 
<< m1 >>
rect 229 206 230 207 
<< m1 >>
rect 230 206 231 207 
<< m1 >>
rect 231 206 232 207 
<< m1 >>
rect 232 206 233 207 
<< m1 >>
rect 233 206 234 207 
<< m2 >>
rect 233 206 234 207 
<< m2c >>
rect 233 206 234 207 
<< m1 >>
rect 233 206 234 207 
<< m2 >>
rect 233 206 234 207 
<< m2 >>
rect 234 206 235 207 
<< m1 >>
rect 235 206 236 207 
<< m2 >>
rect 235 206 236 207 
<< m2 >>
rect 236 206 237 207 
<< m1 >>
rect 237 206 238 207 
<< m2 >>
rect 237 206 238 207 
<< m2c >>
rect 237 206 238 207 
<< m1 >>
rect 237 206 238 207 
<< m2 >>
rect 237 206 238 207 
<< m1 >>
rect 244 206 245 207 
<< m1 >>
rect 250 206 251 207 
<< m1 >>
rect 254 206 255 207 
<< m2 >>
rect 285 206 286 207 
<< m1 >>
rect 286 206 287 207 
<< m2 >>
rect 286 206 287 207 
<< m2 >>
rect 287 206 288 207 
<< m2 >>
rect 288 206 289 207 
<< m2 >>
rect 289 206 290 207 
<< m2 >>
rect 298 206 299 207 
<< m1 >>
rect 307 206 308 207 
<< m2 >>
rect 308 206 309 207 
<< m1 >>
rect 311 206 312 207 
<< m1 >>
rect 337 206 338 207 
<< m1 >>
rect 343 206 344 207 
<< m1 >>
rect 16 207 17 208 
<< m1 >>
rect 19 207 20 208 
<< m1 >>
rect 93 207 94 208 
<< m1 >>
rect 118 207 119 208 
<< m1 >>
rect 121 207 122 208 
<< m1 >>
rect 127 207 128 208 
<< m1 >>
rect 154 207 155 208 
<< m1 >>
rect 179 207 180 208 
<< m1 >>
rect 196 207 197 208 
<< m1 >>
rect 200 207 201 208 
<< m1 >>
rect 207 207 208 208 
<< m1 >>
rect 235 207 236 208 
<< m1 >>
rect 237 207 238 208 
<< m1 >>
rect 244 207 245 208 
<< m2 >>
rect 249 207 250 208 
<< m1 >>
rect 250 207 251 208 
<< m2 >>
rect 250 207 251 208 
<< m2 >>
rect 251 207 252 208 
<< m1 >>
rect 252 207 253 208 
<< m2 >>
rect 252 207 253 208 
<< m2c >>
rect 252 207 253 208 
<< m1 >>
rect 252 207 253 208 
<< m2 >>
rect 252 207 253 208 
<< m1 >>
rect 253 207 254 208 
<< m1 >>
rect 254 207 255 208 
<< m1 >>
rect 286 207 287 208 
<< m1 >>
rect 287 207 288 208 
<< m1 >>
rect 288 207 289 208 
<< m1 >>
rect 289 207 290 208 
<< m2 >>
rect 289 207 290 208 
<< m1 >>
rect 290 207 291 208 
<< m1 >>
rect 291 207 292 208 
<< m1 >>
rect 292 207 293 208 
<< m1 >>
rect 293 207 294 208 
<< m1 >>
rect 294 207 295 208 
<< m1 >>
rect 295 207 296 208 
<< m1 >>
rect 296 207 297 208 
<< m1 >>
rect 297 207 298 208 
<< m1 >>
rect 298 207 299 208 
<< m2 >>
rect 298 207 299 208 
<< m1 >>
rect 307 207 308 208 
<< m2 >>
rect 308 207 309 208 
<< m1 >>
rect 311 207 312 208 
<< m1 >>
rect 337 207 338 208 
<< m1 >>
rect 343 207 344 208 
<< m1 >>
rect 16 208 17 209 
<< m1 >>
rect 19 208 20 209 
<< m1 >>
rect 93 208 94 209 
<< m1 >>
rect 94 208 95 209 
<< m1 >>
rect 95 208 96 209 
<< m1 >>
rect 96 208 97 209 
<< m1 >>
rect 97 208 98 209 
<< m1 >>
rect 98 208 99 209 
<< m1 >>
rect 99 208 100 209 
<< m1 >>
rect 100 208 101 209 
<< m1 >>
rect 101 208 102 209 
<< m1 >>
rect 102 208 103 209 
<< m1 >>
rect 103 208 104 209 
<< m1 >>
rect 104 208 105 209 
<< m1 >>
rect 105 208 106 209 
<< m1 >>
rect 106 208 107 209 
<< m1 >>
rect 107 208 108 209 
<< m1 >>
rect 108 208 109 209 
<< m1 >>
rect 109 208 110 209 
<< m1 >>
rect 110 208 111 209 
<< m1 >>
rect 111 208 112 209 
<< m1 >>
rect 112 208 113 209 
<< m1 >>
rect 113 208 114 209 
<< m1 >>
rect 114 208 115 209 
<< m1 >>
rect 115 208 116 209 
<< m1 >>
rect 116 208 117 209 
<< m2 >>
rect 116 208 117 209 
<< m2c >>
rect 116 208 117 209 
<< m1 >>
rect 116 208 117 209 
<< m2 >>
rect 116 208 117 209 
<< m2 >>
rect 117 208 118 209 
<< m1 >>
rect 118 208 119 209 
<< m1 >>
rect 121 208 122 209 
<< m1 >>
rect 127 208 128 209 
<< m1 >>
rect 154 208 155 209 
<< m2 >>
rect 178 208 179 209 
<< m1 >>
rect 179 208 180 209 
<< m2 >>
rect 179 208 180 209 
<< m1 >>
rect 180 208 181 209 
<< m2 >>
rect 180 208 181 209 
<< m1 >>
rect 181 208 182 209 
<< m2 >>
rect 181 208 182 209 
<< m1 >>
rect 182 208 183 209 
<< m1 >>
rect 183 208 184 209 
<< m1 >>
rect 184 208 185 209 
<< m1 >>
rect 185 208 186 209 
<< m1 >>
rect 186 208 187 209 
<< m1 >>
rect 187 208 188 209 
<< m1 >>
rect 188 208 189 209 
<< m1 >>
rect 189 208 190 209 
<< m1 >>
rect 190 208 191 209 
<< m1 >>
rect 196 208 197 209 
<< m1 >>
rect 200 208 201 209 
<< m1 >>
rect 207 208 208 209 
<< m1 >>
rect 235 208 236 209 
<< m1 >>
rect 237 208 238 209 
<< m1 >>
rect 244 208 245 209 
<< m1 >>
rect 247 208 248 209 
<< m1 >>
rect 248 208 249 209 
<< m2 >>
rect 248 208 249 209 
<< m2c >>
rect 248 208 249 209 
<< m1 >>
rect 248 208 249 209 
<< m2 >>
rect 248 208 249 209 
<< m2 >>
rect 249 208 250 209 
<< m1 >>
rect 250 208 251 209 
<< m2 >>
rect 289 208 290 209 
<< m1 >>
rect 298 208 299 209 
<< m2 >>
rect 298 208 299 209 
<< m1 >>
rect 307 208 308 209 
<< m2 >>
rect 308 208 309 209 
<< m1 >>
rect 311 208 312 209 
<< m1 >>
rect 337 208 338 209 
<< m1 >>
rect 340 208 341 209 
<< m1 >>
rect 341 208 342 209 
<< m1 >>
rect 342 208 343 209 
<< m1 >>
rect 343 208 344 209 
<< m1 >>
rect 448 208 449 209 
<< m1 >>
rect 449 208 450 209 
<< m1 >>
rect 450 208 451 209 
<< m1 >>
rect 451 208 452 209 
<< m1 >>
rect 16 209 17 210 
<< m1 >>
rect 19 209 20 210 
<< m2 >>
rect 117 209 118 210 
<< m1 >>
rect 118 209 119 210 
<< m1 >>
rect 121 209 122 210 
<< m1 >>
rect 127 209 128 210 
<< m1 >>
rect 154 209 155 210 
<< m1 >>
rect 178 209 179 210 
<< m2 >>
rect 178 209 179 210 
<< m2c >>
rect 178 209 179 210 
<< m1 >>
rect 178 209 179 210 
<< m2 >>
rect 178 209 179 210 
<< m2 >>
rect 181 209 182 210 
<< m1 >>
rect 190 209 191 210 
<< m1 >>
rect 196 209 197 210 
<< m1 >>
rect 200 209 201 210 
<< m1 >>
rect 207 209 208 210 
<< m1 >>
rect 235 209 236 210 
<< m1 >>
rect 237 209 238 210 
<< m1 >>
rect 244 209 245 210 
<< m1 >>
rect 247 209 248 210 
<< m1 >>
rect 250 209 251 210 
<< m1 >>
rect 289 209 290 210 
<< m2 >>
rect 289 209 290 210 
<< m2c >>
rect 289 209 290 210 
<< m1 >>
rect 289 209 290 210 
<< m2 >>
rect 289 209 290 210 
<< m1 >>
rect 298 209 299 210 
<< m2 >>
rect 298 209 299 210 
<< m1 >>
rect 307 209 308 210 
<< m2 >>
rect 308 209 309 210 
<< m1 >>
rect 311 209 312 210 
<< m1 >>
rect 337 209 338 210 
<< m1 >>
rect 340 209 341 210 
<< m1 >>
rect 448 209 449 210 
<< m1 >>
rect 451 209 452 210 
<< pdiffusion >>
rect 12 210 13 211 
<< pdiffusion >>
rect 13 210 14 211 
<< pdiffusion >>
rect 14 210 15 211 
<< pdiffusion >>
rect 15 210 16 211 
<< m1 >>
rect 16 210 17 211 
<< pdiffusion >>
rect 16 210 17 211 
<< pdiffusion >>
rect 17 210 18 211 
<< m1 >>
rect 19 210 20 211 
<< pdiffusion >>
rect 30 210 31 211 
<< pdiffusion >>
rect 31 210 32 211 
<< pdiffusion >>
rect 32 210 33 211 
<< pdiffusion >>
rect 33 210 34 211 
<< pdiffusion >>
rect 34 210 35 211 
<< pdiffusion >>
rect 35 210 36 211 
<< pdiffusion >>
rect 48 210 49 211 
<< pdiffusion >>
rect 49 210 50 211 
<< pdiffusion >>
rect 50 210 51 211 
<< pdiffusion >>
rect 51 210 52 211 
<< pdiffusion >>
rect 52 210 53 211 
<< pdiffusion >>
rect 53 210 54 211 
<< pdiffusion >>
rect 84 210 85 211 
<< pdiffusion >>
rect 85 210 86 211 
<< pdiffusion >>
rect 86 210 87 211 
<< pdiffusion >>
rect 87 210 88 211 
<< pdiffusion >>
rect 88 210 89 211 
<< pdiffusion >>
rect 89 210 90 211 
<< m2 >>
rect 117 210 118 211 
<< m1 >>
rect 118 210 119 211 
<< pdiffusion >>
rect 120 210 121 211 
<< m1 >>
rect 121 210 122 211 
<< pdiffusion >>
rect 121 210 122 211 
<< pdiffusion >>
rect 122 210 123 211 
<< pdiffusion >>
rect 123 210 124 211 
<< pdiffusion >>
rect 124 210 125 211 
<< pdiffusion >>
rect 125 210 126 211 
<< m1 >>
rect 127 210 128 211 
<< pdiffusion >>
rect 138 210 139 211 
<< pdiffusion >>
rect 139 210 140 211 
<< pdiffusion >>
rect 140 210 141 211 
<< pdiffusion >>
rect 141 210 142 211 
<< pdiffusion >>
rect 142 210 143 211 
<< pdiffusion >>
rect 143 210 144 211 
<< m1 >>
rect 154 210 155 211 
<< pdiffusion >>
rect 156 210 157 211 
<< pdiffusion >>
rect 157 210 158 211 
<< pdiffusion >>
rect 158 210 159 211 
<< pdiffusion >>
rect 159 210 160 211 
<< pdiffusion >>
rect 160 210 161 211 
<< pdiffusion >>
rect 161 210 162 211 
<< pdiffusion >>
rect 174 210 175 211 
<< pdiffusion >>
rect 175 210 176 211 
<< pdiffusion >>
rect 176 210 177 211 
<< pdiffusion >>
rect 177 210 178 211 
<< m1 >>
rect 178 210 179 211 
<< pdiffusion >>
rect 178 210 179 211 
<< pdiffusion >>
rect 179 210 180 211 
<< m1 >>
rect 181 210 182 211 
<< m2 >>
rect 181 210 182 211 
<< m2c >>
rect 181 210 182 211 
<< m1 >>
rect 181 210 182 211 
<< m2 >>
rect 181 210 182 211 
<< m1 >>
rect 190 210 191 211 
<< pdiffusion >>
rect 192 210 193 211 
<< pdiffusion >>
rect 193 210 194 211 
<< pdiffusion >>
rect 194 210 195 211 
<< pdiffusion >>
rect 195 210 196 211 
<< m1 >>
rect 196 210 197 211 
<< pdiffusion >>
rect 196 210 197 211 
<< pdiffusion >>
rect 197 210 198 211 
<< m1 >>
rect 200 210 201 211 
<< m1 >>
rect 207 210 208 211 
<< pdiffusion >>
rect 210 210 211 211 
<< pdiffusion >>
rect 211 210 212 211 
<< pdiffusion >>
rect 212 210 213 211 
<< pdiffusion >>
rect 213 210 214 211 
<< pdiffusion >>
rect 214 210 215 211 
<< pdiffusion >>
rect 215 210 216 211 
<< m1 >>
rect 235 210 236 211 
<< m1 >>
rect 237 210 238 211 
<< m1 >>
rect 244 210 245 211 
<< pdiffusion >>
rect 246 210 247 211 
<< m1 >>
rect 247 210 248 211 
<< pdiffusion >>
rect 247 210 248 211 
<< pdiffusion >>
rect 248 210 249 211 
<< pdiffusion >>
rect 249 210 250 211 
<< m1 >>
rect 250 210 251 211 
<< pdiffusion >>
rect 250 210 251 211 
<< pdiffusion >>
rect 251 210 252 211 
<< pdiffusion >>
rect 264 210 265 211 
<< pdiffusion >>
rect 265 210 266 211 
<< pdiffusion >>
rect 266 210 267 211 
<< pdiffusion >>
rect 267 210 268 211 
<< pdiffusion >>
rect 268 210 269 211 
<< pdiffusion >>
rect 269 210 270 211 
<< pdiffusion >>
rect 282 210 283 211 
<< pdiffusion >>
rect 283 210 284 211 
<< pdiffusion >>
rect 284 210 285 211 
<< pdiffusion >>
rect 285 210 286 211 
<< pdiffusion >>
rect 286 210 287 211 
<< pdiffusion >>
rect 287 210 288 211 
<< m1 >>
rect 289 210 290 211 
<< m1 >>
rect 298 210 299 211 
<< m2 >>
rect 298 210 299 211 
<< pdiffusion >>
rect 300 210 301 211 
<< pdiffusion >>
rect 301 210 302 211 
<< pdiffusion >>
rect 302 210 303 211 
<< pdiffusion >>
rect 303 210 304 211 
<< pdiffusion >>
rect 304 210 305 211 
<< pdiffusion >>
rect 305 210 306 211 
<< m1 >>
rect 307 210 308 211 
<< m2 >>
rect 308 210 309 211 
<< m1 >>
rect 311 210 312 211 
<< pdiffusion >>
rect 318 210 319 211 
<< pdiffusion >>
rect 319 210 320 211 
<< pdiffusion >>
rect 320 210 321 211 
<< pdiffusion >>
rect 321 210 322 211 
<< pdiffusion >>
rect 322 210 323 211 
<< pdiffusion >>
rect 323 210 324 211 
<< pdiffusion >>
rect 336 210 337 211 
<< m1 >>
rect 337 210 338 211 
<< pdiffusion >>
rect 337 210 338 211 
<< pdiffusion >>
rect 338 210 339 211 
<< pdiffusion >>
rect 339 210 340 211 
<< m1 >>
rect 340 210 341 211 
<< pdiffusion >>
rect 340 210 341 211 
<< pdiffusion >>
rect 341 210 342 211 
<< pdiffusion >>
rect 354 210 355 211 
<< pdiffusion >>
rect 355 210 356 211 
<< pdiffusion >>
rect 356 210 357 211 
<< pdiffusion >>
rect 357 210 358 211 
<< pdiffusion >>
rect 358 210 359 211 
<< pdiffusion >>
rect 359 210 360 211 
<< pdiffusion >>
rect 372 210 373 211 
<< pdiffusion >>
rect 373 210 374 211 
<< pdiffusion >>
rect 374 210 375 211 
<< pdiffusion >>
rect 375 210 376 211 
<< pdiffusion >>
rect 376 210 377 211 
<< pdiffusion >>
rect 377 210 378 211 
<< pdiffusion >>
rect 390 210 391 211 
<< pdiffusion >>
rect 391 210 392 211 
<< pdiffusion >>
rect 392 210 393 211 
<< pdiffusion >>
rect 393 210 394 211 
<< pdiffusion >>
rect 394 210 395 211 
<< pdiffusion >>
rect 395 210 396 211 
<< pdiffusion >>
rect 408 210 409 211 
<< pdiffusion >>
rect 409 210 410 211 
<< pdiffusion >>
rect 410 210 411 211 
<< pdiffusion >>
rect 411 210 412 211 
<< pdiffusion >>
rect 412 210 413 211 
<< pdiffusion >>
rect 413 210 414 211 
<< pdiffusion >>
rect 426 210 427 211 
<< pdiffusion >>
rect 427 210 428 211 
<< pdiffusion >>
rect 428 210 429 211 
<< pdiffusion >>
rect 429 210 430 211 
<< pdiffusion >>
rect 430 210 431 211 
<< pdiffusion >>
rect 431 210 432 211 
<< pdiffusion >>
rect 444 210 445 211 
<< pdiffusion >>
rect 445 210 446 211 
<< pdiffusion >>
rect 446 210 447 211 
<< pdiffusion >>
rect 447 210 448 211 
<< m1 >>
rect 448 210 449 211 
<< pdiffusion >>
rect 448 210 449 211 
<< pdiffusion >>
rect 449 210 450 211 
<< m1 >>
rect 451 210 452 211 
<< pdiffusion >>
rect 12 211 13 212 
<< pdiffusion >>
rect 13 211 14 212 
<< pdiffusion >>
rect 14 211 15 212 
<< pdiffusion >>
rect 15 211 16 212 
<< pdiffusion >>
rect 16 211 17 212 
<< pdiffusion >>
rect 17 211 18 212 
<< m1 >>
rect 19 211 20 212 
<< pdiffusion >>
rect 30 211 31 212 
<< pdiffusion >>
rect 31 211 32 212 
<< pdiffusion >>
rect 32 211 33 212 
<< pdiffusion >>
rect 33 211 34 212 
<< pdiffusion >>
rect 34 211 35 212 
<< pdiffusion >>
rect 35 211 36 212 
<< pdiffusion >>
rect 48 211 49 212 
<< pdiffusion >>
rect 49 211 50 212 
<< pdiffusion >>
rect 50 211 51 212 
<< pdiffusion >>
rect 51 211 52 212 
<< pdiffusion >>
rect 52 211 53 212 
<< pdiffusion >>
rect 53 211 54 212 
<< pdiffusion >>
rect 84 211 85 212 
<< pdiffusion >>
rect 85 211 86 212 
<< pdiffusion >>
rect 86 211 87 212 
<< pdiffusion >>
rect 87 211 88 212 
<< pdiffusion >>
rect 88 211 89 212 
<< pdiffusion >>
rect 89 211 90 212 
<< m2 >>
rect 117 211 118 212 
<< m1 >>
rect 118 211 119 212 
<< pdiffusion >>
rect 120 211 121 212 
<< pdiffusion >>
rect 121 211 122 212 
<< pdiffusion >>
rect 122 211 123 212 
<< pdiffusion >>
rect 123 211 124 212 
<< pdiffusion >>
rect 124 211 125 212 
<< pdiffusion >>
rect 125 211 126 212 
<< m1 >>
rect 127 211 128 212 
<< pdiffusion >>
rect 138 211 139 212 
<< pdiffusion >>
rect 139 211 140 212 
<< pdiffusion >>
rect 140 211 141 212 
<< pdiffusion >>
rect 141 211 142 212 
<< pdiffusion >>
rect 142 211 143 212 
<< pdiffusion >>
rect 143 211 144 212 
<< m1 >>
rect 154 211 155 212 
<< pdiffusion >>
rect 156 211 157 212 
<< pdiffusion >>
rect 157 211 158 212 
<< pdiffusion >>
rect 158 211 159 212 
<< pdiffusion >>
rect 159 211 160 212 
<< pdiffusion >>
rect 160 211 161 212 
<< pdiffusion >>
rect 161 211 162 212 
<< pdiffusion >>
rect 174 211 175 212 
<< pdiffusion >>
rect 175 211 176 212 
<< pdiffusion >>
rect 176 211 177 212 
<< pdiffusion >>
rect 177 211 178 212 
<< pdiffusion >>
rect 178 211 179 212 
<< pdiffusion >>
rect 179 211 180 212 
<< m1 >>
rect 181 211 182 212 
<< m1 >>
rect 190 211 191 212 
<< pdiffusion >>
rect 192 211 193 212 
<< pdiffusion >>
rect 193 211 194 212 
<< pdiffusion >>
rect 194 211 195 212 
<< pdiffusion >>
rect 195 211 196 212 
<< pdiffusion >>
rect 196 211 197 212 
<< pdiffusion >>
rect 197 211 198 212 
<< m1 >>
rect 200 211 201 212 
<< m1 >>
rect 207 211 208 212 
<< pdiffusion >>
rect 210 211 211 212 
<< pdiffusion >>
rect 211 211 212 212 
<< pdiffusion >>
rect 212 211 213 212 
<< pdiffusion >>
rect 213 211 214 212 
<< pdiffusion >>
rect 214 211 215 212 
<< pdiffusion >>
rect 215 211 216 212 
<< m1 >>
rect 235 211 236 212 
<< m1 >>
rect 237 211 238 212 
<< m1 >>
rect 244 211 245 212 
<< pdiffusion >>
rect 246 211 247 212 
<< pdiffusion >>
rect 247 211 248 212 
<< pdiffusion >>
rect 248 211 249 212 
<< pdiffusion >>
rect 249 211 250 212 
<< pdiffusion >>
rect 250 211 251 212 
<< pdiffusion >>
rect 251 211 252 212 
<< pdiffusion >>
rect 264 211 265 212 
<< pdiffusion >>
rect 265 211 266 212 
<< pdiffusion >>
rect 266 211 267 212 
<< pdiffusion >>
rect 267 211 268 212 
<< pdiffusion >>
rect 268 211 269 212 
<< pdiffusion >>
rect 269 211 270 212 
<< pdiffusion >>
rect 282 211 283 212 
<< pdiffusion >>
rect 283 211 284 212 
<< pdiffusion >>
rect 284 211 285 212 
<< pdiffusion >>
rect 285 211 286 212 
<< pdiffusion >>
rect 286 211 287 212 
<< pdiffusion >>
rect 287 211 288 212 
<< m1 >>
rect 289 211 290 212 
<< m1 >>
rect 298 211 299 212 
<< m2 >>
rect 298 211 299 212 
<< pdiffusion >>
rect 300 211 301 212 
<< pdiffusion >>
rect 301 211 302 212 
<< pdiffusion >>
rect 302 211 303 212 
<< pdiffusion >>
rect 303 211 304 212 
<< pdiffusion >>
rect 304 211 305 212 
<< pdiffusion >>
rect 305 211 306 212 
<< m1 >>
rect 307 211 308 212 
<< m2 >>
rect 308 211 309 212 
<< m1 >>
rect 311 211 312 212 
<< pdiffusion >>
rect 318 211 319 212 
<< pdiffusion >>
rect 319 211 320 212 
<< pdiffusion >>
rect 320 211 321 212 
<< pdiffusion >>
rect 321 211 322 212 
<< pdiffusion >>
rect 322 211 323 212 
<< pdiffusion >>
rect 323 211 324 212 
<< pdiffusion >>
rect 336 211 337 212 
<< pdiffusion >>
rect 337 211 338 212 
<< pdiffusion >>
rect 338 211 339 212 
<< pdiffusion >>
rect 339 211 340 212 
<< pdiffusion >>
rect 340 211 341 212 
<< pdiffusion >>
rect 341 211 342 212 
<< pdiffusion >>
rect 354 211 355 212 
<< pdiffusion >>
rect 355 211 356 212 
<< pdiffusion >>
rect 356 211 357 212 
<< pdiffusion >>
rect 357 211 358 212 
<< pdiffusion >>
rect 358 211 359 212 
<< pdiffusion >>
rect 359 211 360 212 
<< pdiffusion >>
rect 372 211 373 212 
<< pdiffusion >>
rect 373 211 374 212 
<< pdiffusion >>
rect 374 211 375 212 
<< pdiffusion >>
rect 375 211 376 212 
<< pdiffusion >>
rect 376 211 377 212 
<< pdiffusion >>
rect 377 211 378 212 
<< pdiffusion >>
rect 390 211 391 212 
<< pdiffusion >>
rect 391 211 392 212 
<< pdiffusion >>
rect 392 211 393 212 
<< pdiffusion >>
rect 393 211 394 212 
<< pdiffusion >>
rect 394 211 395 212 
<< pdiffusion >>
rect 395 211 396 212 
<< pdiffusion >>
rect 408 211 409 212 
<< pdiffusion >>
rect 409 211 410 212 
<< pdiffusion >>
rect 410 211 411 212 
<< pdiffusion >>
rect 411 211 412 212 
<< pdiffusion >>
rect 412 211 413 212 
<< pdiffusion >>
rect 413 211 414 212 
<< pdiffusion >>
rect 426 211 427 212 
<< pdiffusion >>
rect 427 211 428 212 
<< pdiffusion >>
rect 428 211 429 212 
<< pdiffusion >>
rect 429 211 430 212 
<< pdiffusion >>
rect 430 211 431 212 
<< pdiffusion >>
rect 431 211 432 212 
<< pdiffusion >>
rect 444 211 445 212 
<< pdiffusion >>
rect 445 211 446 212 
<< pdiffusion >>
rect 446 211 447 212 
<< pdiffusion >>
rect 447 211 448 212 
<< pdiffusion >>
rect 448 211 449 212 
<< pdiffusion >>
rect 449 211 450 212 
<< m1 >>
rect 451 211 452 212 
<< pdiffusion >>
rect 12 212 13 213 
<< pdiffusion >>
rect 13 212 14 213 
<< pdiffusion >>
rect 14 212 15 213 
<< pdiffusion >>
rect 15 212 16 213 
<< pdiffusion >>
rect 16 212 17 213 
<< pdiffusion >>
rect 17 212 18 213 
<< m1 >>
rect 19 212 20 213 
<< pdiffusion >>
rect 30 212 31 213 
<< pdiffusion >>
rect 31 212 32 213 
<< pdiffusion >>
rect 32 212 33 213 
<< pdiffusion >>
rect 33 212 34 213 
<< pdiffusion >>
rect 34 212 35 213 
<< pdiffusion >>
rect 35 212 36 213 
<< pdiffusion >>
rect 48 212 49 213 
<< pdiffusion >>
rect 49 212 50 213 
<< pdiffusion >>
rect 50 212 51 213 
<< pdiffusion >>
rect 51 212 52 213 
<< pdiffusion >>
rect 52 212 53 213 
<< pdiffusion >>
rect 53 212 54 213 
<< pdiffusion >>
rect 84 212 85 213 
<< pdiffusion >>
rect 85 212 86 213 
<< pdiffusion >>
rect 86 212 87 213 
<< pdiffusion >>
rect 87 212 88 213 
<< pdiffusion >>
rect 88 212 89 213 
<< pdiffusion >>
rect 89 212 90 213 
<< m2 >>
rect 117 212 118 213 
<< m1 >>
rect 118 212 119 213 
<< pdiffusion >>
rect 120 212 121 213 
<< pdiffusion >>
rect 121 212 122 213 
<< pdiffusion >>
rect 122 212 123 213 
<< pdiffusion >>
rect 123 212 124 213 
<< pdiffusion >>
rect 124 212 125 213 
<< pdiffusion >>
rect 125 212 126 213 
<< m1 >>
rect 127 212 128 213 
<< pdiffusion >>
rect 138 212 139 213 
<< pdiffusion >>
rect 139 212 140 213 
<< pdiffusion >>
rect 140 212 141 213 
<< pdiffusion >>
rect 141 212 142 213 
<< pdiffusion >>
rect 142 212 143 213 
<< pdiffusion >>
rect 143 212 144 213 
<< m1 >>
rect 154 212 155 213 
<< pdiffusion >>
rect 156 212 157 213 
<< pdiffusion >>
rect 157 212 158 213 
<< pdiffusion >>
rect 158 212 159 213 
<< pdiffusion >>
rect 159 212 160 213 
<< pdiffusion >>
rect 160 212 161 213 
<< pdiffusion >>
rect 161 212 162 213 
<< pdiffusion >>
rect 174 212 175 213 
<< pdiffusion >>
rect 175 212 176 213 
<< pdiffusion >>
rect 176 212 177 213 
<< pdiffusion >>
rect 177 212 178 213 
<< pdiffusion >>
rect 178 212 179 213 
<< pdiffusion >>
rect 179 212 180 213 
<< m1 >>
rect 181 212 182 213 
<< m1 >>
rect 190 212 191 213 
<< pdiffusion >>
rect 192 212 193 213 
<< pdiffusion >>
rect 193 212 194 213 
<< pdiffusion >>
rect 194 212 195 213 
<< pdiffusion >>
rect 195 212 196 213 
<< pdiffusion >>
rect 196 212 197 213 
<< pdiffusion >>
rect 197 212 198 213 
<< m1 >>
rect 200 212 201 213 
<< m1 >>
rect 207 212 208 213 
<< pdiffusion >>
rect 210 212 211 213 
<< pdiffusion >>
rect 211 212 212 213 
<< pdiffusion >>
rect 212 212 213 213 
<< pdiffusion >>
rect 213 212 214 213 
<< pdiffusion >>
rect 214 212 215 213 
<< pdiffusion >>
rect 215 212 216 213 
<< m1 >>
rect 235 212 236 213 
<< m1 >>
rect 237 212 238 213 
<< m1 >>
rect 244 212 245 213 
<< pdiffusion >>
rect 246 212 247 213 
<< pdiffusion >>
rect 247 212 248 213 
<< pdiffusion >>
rect 248 212 249 213 
<< pdiffusion >>
rect 249 212 250 213 
<< pdiffusion >>
rect 250 212 251 213 
<< pdiffusion >>
rect 251 212 252 213 
<< pdiffusion >>
rect 264 212 265 213 
<< pdiffusion >>
rect 265 212 266 213 
<< pdiffusion >>
rect 266 212 267 213 
<< pdiffusion >>
rect 267 212 268 213 
<< pdiffusion >>
rect 268 212 269 213 
<< pdiffusion >>
rect 269 212 270 213 
<< pdiffusion >>
rect 282 212 283 213 
<< pdiffusion >>
rect 283 212 284 213 
<< pdiffusion >>
rect 284 212 285 213 
<< pdiffusion >>
rect 285 212 286 213 
<< pdiffusion >>
rect 286 212 287 213 
<< pdiffusion >>
rect 287 212 288 213 
<< m1 >>
rect 289 212 290 213 
<< m1 >>
rect 298 212 299 213 
<< m2 >>
rect 298 212 299 213 
<< pdiffusion >>
rect 300 212 301 213 
<< pdiffusion >>
rect 301 212 302 213 
<< pdiffusion >>
rect 302 212 303 213 
<< pdiffusion >>
rect 303 212 304 213 
<< pdiffusion >>
rect 304 212 305 213 
<< pdiffusion >>
rect 305 212 306 213 
<< m1 >>
rect 307 212 308 213 
<< m2 >>
rect 308 212 309 213 
<< m1 >>
rect 311 212 312 213 
<< pdiffusion >>
rect 318 212 319 213 
<< pdiffusion >>
rect 319 212 320 213 
<< pdiffusion >>
rect 320 212 321 213 
<< pdiffusion >>
rect 321 212 322 213 
<< pdiffusion >>
rect 322 212 323 213 
<< pdiffusion >>
rect 323 212 324 213 
<< pdiffusion >>
rect 336 212 337 213 
<< pdiffusion >>
rect 337 212 338 213 
<< pdiffusion >>
rect 338 212 339 213 
<< pdiffusion >>
rect 339 212 340 213 
<< pdiffusion >>
rect 340 212 341 213 
<< pdiffusion >>
rect 341 212 342 213 
<< pdiffusion >>
rect 354 212 355 213 
<< pdiffusion >>
rect 355 212 356 213 
<< pdiffusion >>
rect 356 212 357 213 
<< pdiffusion >>
rect 357 212 358 213 
<< pdiffusion >>
rect 358 212 359 213 
<< pdiffusion >>
rect 359 212 360 213 
<< pdiffusion >>
rect 372 212 373 213 
<< pdiffusion >>
rect 373 212 374 213 
<< pdiffusion >>
rect 374 212 375 213 
<< pdiffusion >>
rect 375 212 376 213 
<< pdiffusion >>
rect 376 212 377 213 
<< pdiffusion >>
rect 377 212 378 213 
<< pdiffusion >>
rect 390 212 391 213 
<< pdiffusion >>
rect 391 212 392 213 
<< pdiffusion >>
rect 392 212 393 213 
<< pdiffusion >>
rect 393 212 394 213 
<< pdiffusion >>
rect 394 212 395 213 
<< pdiffusion >>
rect 395 212 396 213 
<< pdiffusion >>
rect 408 212 409 213 
<< pdiffusion >>
rect 409 212 410 213 
<< pdiffusion >>
rect 410 212 411 213 
<< pdiffusion >>
rect 411 212 412 213 
<< pdiffusion >>
rect 412 212 413 213 
<< pdiffusion >>
rect 413 212 414 213 
<< pdiffusion >>
rect 426 212 427 213 
<< pdiffusion >>
rect 427 212 428 213 
<< pdiffusion >>
rect 428 212 429 213 
<< pdiffusion >>
rect 429 212 430 213 
<< pdiffusion >>
rect 430 212 431 213 
<< pdiffusion >>
rect 431 212 432 213 
<< pdiffusion >>
rect 444 212 445 213 
<< pdiffusion >>
rect 445 212 446 213 
<< pdiffusion >>
rect 446 212 447 213 
<< pdiffusion >>
rect 447 212 448 213 
<< pdiffusion >>
rect 448 212 449 213 
<< pdiffusion >>
rect 449 212 450 213 
<< m1 >>
rect 451 212 452 213 
<< pdiffusion >>
rect 12 213 13 214 
<< pdiffusion >>
rect 13 213 14 214 
<< pdiffusion >>
rect 14 213 15 214 
<< pdiffusion >>
rect 15 213 16 214 
<< pdiffusion >>
rect 16 213 17 214 
<< pdiffusion >>
rect 17 213 18 214 
<< m1 >>
rect 19 213 20 214 
<< pdiffusion >>
rect 30 213 31 214 
<< pdiffusion >>
rect 31 213 32 214 
<< pdiffusion >>
rect 32 213 33 214 
<< pdiffusion >>
rect 33 213 34 214 
<< pdiffusion >>
rect 34 213 35 214 
<< pdiffusion >>
rect 35 213 36 214 
<< pdiffusion >>
rect 48 213 49 214 
<< pdiffusion >>
rect 49 213 50 214 
<< pdiffusion >>
rect 50 213 51 214 
<< pdiffusion >>
rect 51 213 52 214 
<< pdiffusion >>
rect 52 213 53 214 
<< pdiffusion >>
rect 53 213 54 214 
<< pdiffusion >>
rect 84 213 85 214 
<< pdiffusion >>
rect 85 213 86 214 
<< pdiffusion >>
rect 86 213 87 214 
<< pdiffusion >>
rect 87 213 88 214 
<< pdiffusion >>
rect 88 213 89 214 
<< pdiffusion >>
rect 89 213 90 214 
<< m2 >>
rect 117 213 118 214 
<< m1 >>
rect 118 213 119 214 
<< pdiffusion >>
rect 120 213 121 214 
<< pdiffusion >>
rect 121 213 122 214 
<< pdiffusion >>
rect 122 213 123 214 
<< pdiffusion >>
rect 123 213 124 214 
<< pdiffusion >>
rect 124 213 125 214 
<< pdiffusion >>
rect 125 213 126 214 
<< m1 >>
rect 127 213 128 214 
<< pdiffusion >>
rect 138 213 139 214 
<< pdiffusion >>
rect 139 213 140 214 
<< pdiffusion >>
rect 140 213 141 214 
<< pdiffusion >>
rect 141 213 142 214 
<< pdiffusion >>
rect 142 213 143 214 
<< pdiffusion >>
rect 143 213 144 214 
<< m1 >>
rect 154 213 155 214 
<< pdiffusion >>
rect 156 213 157 214 
<< pdiffusion >>
rect 157 213 158 214 
<< pdiffusion >>
rect 158 213 159 214 
<< pdiffusion >>
rect 159 213 160 214 
<< pdiffusion >>
rect 160 213 161 214 
<< pdiffusion >>
rect 161 213 162 214 
<< pdiffusion >>
rect 174 213 175 214 
<< pdiffusion >>
rect 175 213 176 214 
<< pdiffusion >>
rect 176 213 177 214 
<< pdiffusion >>
rect 177 213 178 214 
<< pdiffusion >>
rect 178 213 179 214 
<< pdiffusion >>
rect 179 213 180 214 
<< m1 >>
rect 181 213 182 214 
<< m1 >>
rect 190 213 191 214 
<< pdiffusion >>
rect 192 213 193 214 
<< pdiffusion >>
rect 193 213 194 214 
<< pdiffusion >>
rect 194 213 195 214 
<< pdiffusion >>
rect 195 213 196 214 
<< pdiffusion >>
rect 196 213 197 214 
<< pdiffusion >>
rect 197 213 198 214 
<< m1 >>
rect 200 213 201 214 
<< m1 >>
rect 207 213 208 214 
<< pdiffusion >>
rect 210 213 211 214 
<< pdiffusion >>
rect 211 213 212 214 
<< pdiffusion >>
rect 212 213 213 214 
<< pdiffusion >>
rect 213 213 214 214 
<< pdiffusion >>
rect 214 213 215 214 
<< pdiffusion >>
rect 215 213 216 214 
<< m1 >>
rect 235 213 236 214 
<< m1 >>
rect 237 213 238 214 
<< m1 >>
rect 244 213 245 214 
<< pdiffusion >>
rect 246 213 247 214 
<< pdiffusion >>
rect 247 213 248 214 
<< pdiffusion >>
rect 248 213 249 214 
<< pdiffusion >>
rect 249 213 250 214 
<< pdiffusion >>
rect 250 213 251 214 
<< pdiffusion >>
rect 251 213 252 214 
<< pdiffusion >>
rect 264 213 265 214 
<< pdiffusion >>
rect 265 213 266 214 
<< pdiffusion >>
rect 266 213 267 214 
<< pdiffusion >>
rect 267 213 268 214 
<< pdiffusion >>
rect 268 213 269 214 
<< pdiffusion >>
rect 269 213 270 214 
<< pdiffusion >>
rect 282 213 283 214 
<< pdiffusion >>
rect 283 213 284 214 
<< pdiffusion >>
rect 284 213 285 214 
<< pdiffusion >>
rect 285 213 286 214 
<< pdiffusion >>
rect 286 213 287 214 
<< pdiffusion >>
rect 287 213 288 214 
<< m1 >>
rect 289 213 290 214 
<< m1 >>
rect 298 213 299 214 
<< m2 >>
rect 298 213 299 214 
<< pdiffusion >>
rect 300 213 301 214 
<< pdiffusion >>
rect 301 213 302 214 
<< pdiffusion >>
rect 302 213 303 214 
<< pdiffusion >>
rect 303 213 304 214 
<< pdiffusion >>
rect 304 213 305 214 
<< pdiffusion >>
rect 305 213 306 214 
<< m1 >>
rect 307 213 308 214 
<< m2 >>
rect 308 213 309 214 
<< m1 >>
rect 311 213 312 214 
<< pdiffusion >>
rect 318 213 319 214 
<< pdiffusion >>
rect 319 213 320 214 
<< pdiffusion >>
rect 320 213 321 214 
<< pdiffusion >>
rect 321 213 322 214 
<< pdiffusion >>
rect 322 213 323 214 
<< pdiffusion >>
rect 323 213 324 214 
<< pdiffusion >>
rect 336 213 337 214 
<< pdiffusion >>
rect 337 213 338 214 
<< pdiffusion >>
rect 338 213 339 214 
<< pdiffusion >>
rect 339 213 340 214 
<< pdiffusion >>
rect 340 213 341 214 
<< pdiffusion >>
rect 341 213 342 214 
<< pdiffusion >>
rect 354 213 355 214 
<< pdiffusion >>
rect 355 213 356 214 
<< pdiffusion >>
rect 356 213 357 214 
<< pdiffusion >>
rect 357 213 358 214 
<< pdiffusion >>
rect 358 213 359 214 
<< pdiffusion >>
rect 359 213 360 214 
<< pdiffusion >>
rect 372 213 373 214 
<< pdiffusion >>
rect 373 213 374 214 
<< pdiffusion >>
rect 374 213 375 214 
<< pdiffusion >>
rect 375 213 376 214 
<< pdiffusion >>
rect 376 213 377 214 
<< pdiffusion >>
rect 377 213 378 214 
<< pdiffusion >>
rect 390 213 391 214 
<< pdiffusion >>
rect 391 213 392 214 
<< pdiffusion >>
rect 392 213 393 214 
<< pdiffusion >>
rect 393 213 394 214 
<< pdiffusion >>
rect 394 213 395 214 
<< pdiffusion >>
rect 395 213 396 214 
<< pdiffusion >>
rect 408 213 409 214 
<< pdiffusion >>
rect 409 213 410 214 
<< pdiffusion >>
rect 410 213 411 214 
<< pdiffusion >>
rect 411 213 412 214 
<< pdiffusion >>
rect 412 213 413 214 
<< pdiffusion >>
rect 413 213 414 214 
<< pdiffusion >>
rect 426 213 427 214 
<< pdiffusion >>
rect 427 213 428 214 
<< pdiffusion >>
rect 428 213 429 214 
<< pdiffusion >>
rect 429 213 430 214 
<< pdiffusion >>
rect 430 213 431 214 
<< pdiffusion >>
rect 431 213 432 214 
<< pdiffusion >>
rect 444 213 445 214 
<< pdiffusion >>
rect 445 213 446 214 
<< pdiffusion >>
rect 446 213 447 214 
<< pdiffusion >>
rect 447 213 448 214 
<< pdiffusion >>
rect 448 213 449 214 
<< pdiffusion >>
rect 449 213 450 214 
<< m1 >>
rect 451 213 452 214 
<< pdiffusion >>
rect 12 214 13 215 
<< pdiffusion >>
rect 13 214 14 215 
<< pdiffusion >>
rect 14 214 15 215 
<< pdiffusion >>
rect 15 214 16 215 
<< pdiffusion >>
rect 16 214 17 215 
<< pdiffusion >>
rect 17 214 18 215 
<< m1 >>
rect 19 214 20 215 
<< pdiffusion >>
rect 30 214 31 215 
<< pdiffusion >>
rect 31 214 32 215 
<< pdiffusion >>
rect 32 214 33 215 
<< pdiffusion >>
rect 33 214 34 215 
<< pdiffusion >>
rect 34 214 35 215 
<< pdiffusion >>
rect 35 214 36 215 
<< pdiffusion >>
rect 48 214 49 215 
<< pdiffusion >>
rect 49 214 50 215 
<< pdiffusion >>
rect 50 214 51 215 
<< pdiffusion >>
rect 51 214 52 215 
<< pdiffusion >>
rect 52 214 53 215 
<< pdiffusion >>
rect 53 214 54 215 
<< pdiffusion >>
rect 84 214 85 215 
<< pdiffusion >>
rect 85 214 86 215 
<< pdiffusion >>
rect 86 214 87 215 
<< pdiffusion >>
rect 87 214 88 215 
<< pdiffusion >>
rect 88 214 89 215 
<< pdiffusion >>
rect 89 214 90 215 
<< m2 >>
rect 117 214 118 215 
<< m1 >>
rect 118 214 119 215 
<< pdiffusion >>
rect 120 214 121 215 
<< pdiffusion >>
rect 121 214 122 215 
<< pdiffusion >>
rect 122 214 123 215 
<< pdiffusion >>
rect 123 214 124 215 
<< pdiffusion >>
rect 124 214 125 215 
<< pdiffusion >>
rect 125 214 126 215 
<< m1 >>
rect 127 214 128 215 
<< pdiffusion >>
rect 138 214 139 215 
<< pdiffusion >>
rect 139 214 140 215 
<< pdiffusion >>
rect 140 214 141 215 
<< pdiffusion >>
rect 141 214 142 215 
<< pdiffusion >>
rect 142 214 143 215 
<< pdiffusion >>
rect 143 214 144 215 
<< m1 >>
rect 154 214 155 215 
<< pdiffusion >>
rect 156 214 157 215 
<< pdiffusion >>
rect 157 214 158 215 
<< pdiffusion >>
rect 158 214 159 215 
<< pdiffusion >>
rect 159 214 160 215 
<< pdiffusion >>
rect 160 214 161 215 
<< pdiffusion >>
rect 161 214 162 215 
<< pdiffusion >>
rect 174 214 175 215 
<< pdiffusion >>
rect 175 214 176 215 
<< pdiffusion >>
rect 176 214 177 215 
<< pdiffusion >>
rect 177 214 178 215 
<< pdiffusion >>
rect 178 214 179 215 
<< pdiffusion >>
rect 179 214 180 215 
<< m1 >>
rect 181 214 182 215 
<< m1 >>
rect 190 214 191 215 
<< pdiffusion >>
rect 192 214 193 215 
<< pdiffusion >>
rect 193 214 194 215 
<< pdiffusion >>
rect 194 214 195 215 
<< pdiffusion >>
rect 195 214 196 215 
<< pdiffusion >>
rect 196 214 197 215 
<< pdiffusion >>
rect 197 214 198 215 
<< m1 >>
rect 200 214 201 215 
<< m1 >>
rect 207 214 208 215 
<< pdiffusion >>
rect 210 214 211 215 
<< pdiffusion >>
rect 211 214 212 215 
<< pdiffusion >>
rect 212 214 213 215 
<< pdiffusion >>
rect 213 214 214 215 
<< pdiffusion >>
rect 214 214 215 215 
<< pdiffusion >>
rect 215 214 216 215 
<< m1 >>
rect 235 214 236 215 
<< m1 >>
rect 237 214 238 215 
<< m1 >>
rect 244 214 245 215 
<< pdiffusion >>
rect 246 214 247 215 
<< pdiffusion >>
rect 247 214 248 215 
<< pdiffusion >>
rect 248 214 249 215 
<< pdiffusion >>
rect 249 214 250 215 
<< pdiffusion >>
rect 250 214 251 215 
<< pdiffusion >>
rect 251 214 252 215 
<< pdiffusion >>
rect 264 214 265 215 
<< pdiffusion >>
rect 265 214 266 215 
<< pdiffusion >>
rect 266 214 267 215 
<< pdiffusion >>
rect 267 214 268 215 
<< pdiffusion >>
rect 268 214 269 215 
<< pdiffusion >>
rect 269 214 270 215 
<< pdiffusion >>
rect 282 214 283 215 
<< pdiffusion >>
rect 283 214 284 215 
<< pdiffusion >>
rect 284 214 285 215 
<< pdiffusion >>
rect 285 214 286 215 
<< pdiffusion >>
rect 286 214 287 215 
<< pdiffusion >>
rect 287 214 288 215 
<< m1 >>
rect 289 214 290 215 
<< m1 >>
rect 298 214 299 215 
<< m2 >>
rect 298 214 299 215 
<< pdiffusion >>
rect 300 214 301 215 
<< pdiffusion >>
rect 301 214 302 215 
<< pdiffusion >>
rect 302 214 303 215 
<< pdiffusion >>
rect 303 214 304 215 
<< pdiffusion >>
rect 304 214 305 215 
<< pdiffusion >>
rect 305 214 306 215 
<< m1 >>
rect 307 214 308 215 
<< m2 >>
rect 308 214 309 215 
<< m1 >>
rect 311 214 312 215 
<< pdiffusion >>
rect 318 214 319 215 
<< pdiffusion >>
rect 319 214 320 215 
<< pdiffusion >>
rect 320 214 321 215 
<< pdiffusion >>
rect 321 214 322 215 
<< pdiffusion >>
rect 322 214 323 215 
<< pdiffusion >>
rect 323 214 324 215 
<< pdiffusion >>
rect 336 214 337 215 
<< pdiffusion >>
rect 337 214 338 215 
<< pdiffusion >>
rect 338 214 339 215 
<< pdiffusion >>
rect 339 214 340 215 
<< pdiffusion >>
rect 340 214 341 215 
<< pdiffusion >>
rect 341 214 342 215 
<< pdiffusion >>
rect 354 214 355 215 
<< pdiffusion >>
rect 355 214 356 215 
<< pdiffusion >>
rect 356 214 357 215 
<< pdiffusion >>
rect 357 214 358 215 
<< pdiffusion >>
rect 358 214 359 215 
<< pdiffusion >>
rect 359 214 360 215 
<< pdiffusion >>
rect 372 214 373 215 
<< pdiffusion >>
rect 373 214 374 215 
<< pdiffusion >>
rect 374 214 375 215 
<< pdiffusion >>
rect 375 214 376 215 
<< pdiffusion >>
rect 376 214 377 215 
<< pdiffusion >>
rect 377 214 378 215 
<< pdiffusion >>
rect 390 214 391 215 
<< pdiffusion >>
rect 391 214 392 215 
<< pdiffusion >>
rect 392 214 393 215 
<< pdiffusion >>
rect 393 214 394 215 
<< pdiffusion >>
rect 394 214 395 215 
<< pdiffusion >>
rect 395 214 396 215 
<< pdiffusion >>
rect 408 214 409 215 
<< pdiffusion >>
rect 409 214 410 215 
<< pdiffusion >>
rect 410 214 411 215 
<< pdiffusion >>
rect 411 214 412 215 
<< pdiffusion >>
rect 412 214 413 215 
<< pdiffusion >>
rect 413 214 414 215 
<< pdiffusion >>
rect 426 214 427 215 
<< pdiffusion >>
rect 427 214 428 215 
<< pdiffusion >>
rect 428 214 429 215 
<< pdiffusion >>
rect 429 214 430 215 
<< pdiffusion >>
rect 430 214 431 215 
<< pdiffusion >>
rect 431 214 432 215 
<< pdiffusion >>
rect 444 214 445 215 
<< pdiffusion >>
rect 445 214 446 215 
<< pdiffusion >>
rect 446 214 447 215 
<< pdiffusion >>
rect 447 214 448 215 
<< pdiffusion >>
rect 448 214 449 215 
<< pdiffusion >>
rect 449 214 450 215 
<< m1 >>
rect 451 214 452 215 
<< pdiffusion >>
rect 12 215 13 216 
<< pdiffusion >>
rect 13 215 14 216 
<< pdiffusion >>
rect 14 215 15 216 
<< pdiffusion >>
rect 15 215 16 216 
<< pdiffusion >>
rect 16 215 17 216 
<< pdiffusion >>
rect 17 215 18 216 
<< m1 >>
rect 19 215 20 216 
<< pdiffusion >>
rect 30 215 31 216 
<< pdiffusion >>
rect 31 215 32 216 
<< pdiffusion >>
rect 32 215 33 216 
<< pdiffusion >>
rect 33 215 34 216 
<< pdiffusion >>
rect 34 215 35 216 
<< pdiffusion >>
rect 35 215 36 216 
<< pdiffusion >>
rect 48 215 49 216 
<< m1 >>
rect 49 215 50 216 
<< pdiffusion >>
rect 49 215 50 216 
<< pdiffusion >>
rect 50 215 51 216 
<< pdiffusion >>
rect 51 215 52 216 
<< pdiffusion >>
rect 52 215 53 216 
<< pdiffusion >>
rect 53 215 54 216 
<< pdiffusion >>
rect 84 215 85 216 
<< pdiffusion >>
rect 85 215 86 216 
<< pdiffusion >>
rect 86 215 87 216 
<< pdiffusion >>
rect 87 215 88 216 
<< pdiffusion >>
rect 88 215 89 216 
<< pdiffusion >>
rect 89 215 90 216 
<< m2 >>
rect 117 215 118 216 
<< m1 >>
rect 118 215 119 216 
<< pdiffusion >>
rect 120 215 121 216 
<< m1 >>
rect 121 215 122 216 
<< pdiffusion >>
rect 121 215 122 216 
<< pdiffusion >>
rect 122 215 123 216 
<< pdiffusion >>
rect 123 215 124 216 
<< pdiffusion >>
rect 124 215 125 216 
<< pdiffusion >>
rect 125 215 126 216 
<< m1 >>
rect 127 215 128 216 
<< pdiffusion >>
rect 138 215 139 216 
<< pdiffusion >>
rect 139 215 140 216 
<< pdiffusion >>
rect 140 215 141 216 
<< pdiffusion >>
rect 141 215 142 216 
<< m1 >>
rect 142 215 143 216 
<< pdiffusion >>
rect 142 215 143 216 
<< pdiffusion >>
rect 143 215 144 216 
<< m1 >>
rect 154 215 155 216 
<< pdiffusion >>
rect 156 215 157 216 
<< pdiffusion >>
rect 157 215 158 216 
<< pdiffusion >>
rect 158 215 159 216 
<< pdiffusion >>
rect 159 215 160 216 
<< pdiffusion >>
rect 160 215 161 216 
<< pdiffusion >>
rect 161 215 162 216 
<< pdiffusion >>
rect 174 215 175 216 
<< pdiffusion >>
rect 175 215 176 216 
<< pdiffusion >>
rect 176 215 177 216 
<< pdiffusion >>
rect 177 215 178 216 
<< m1 >>
rect 178 215 179 216 
<< pdiffusion >>
rect 178 215 179 216 
<< pdiffusion >>
rect 179 215 180 216 
<< m1 >>
rect 181 215 182 216 
<< m2 >>
rect 181 215 182 216 
<< m2c >>
rect 181 215 182 216 
<< m1 >>
rect 181 215 182 216 
<< m2 >>
rect 181 215 182 216 
<< m1 >>
rect 190 215 191 216 
<< pdiffusion >>
rect 192 215 193 216 
<< pdiffusion >>
rect 193 215 194 216 
<< pdiffusion >>
rect 194 215 195 216 
<< pdiffusion >>
rect 195 215 196 216 
<< m1 >>
rect 196 215 197 216 
<< pdiffusion >>
rect 196 215 197 216 
<< pdiffusion >>
rect 197 215 198 216 
<< m1 >>
rect 200 215 201 216 
<< m1 >>
rect 207 215 208 216 
<< pdiffusion >>
rect 210 215 211 216 
<< pdiffusion >>
rect 211 215 212 216 
<< pdiffusion >>
rect 212 215 213 216 
<< pdiffusion >>
rect 213 215 214 216 
<< pdiffusion >>
rect 214 215 215 216 
<< pdiffusion >>
rect 215 215 216 216 
<< m1 >>
rect 235 215 236 216 
<< m1 >>
rect 237 215 238 216 
<< m1 >>
rect 244 215 245 216 
<< pdiffusion >>
rect 246 215 247 216 
<< pdiffusion >>
rect 247 215 248 216 
<< pdiffusion >>
rect 248 215 249 216 
<< pdiffusion >>
rect 249 215 250 216 
<< pdiffusion >>
rect 250 215 251 216 
<< pdiffusion >>
rect 251 215 252 216 
<< pdiffusion >>
rect 264 215 265 216 
<< pdiffusion >>
rect 265 215 266 216 
<< pdiffusion >>
rect 266 215 267 216 
<< pdiffusion >>
rect 267 215 268 216 
<< m1 >>
rect 268 215 269 216 
<< pdiffusion >>
rect 268 215 269 216 
<< pdiffusion >>
rect 269 215 270 216 
<< pdiffusion >>
rect 282 215 283 216 
<< pdiffusion >>
rect 283 215 284 216 
<< pdiffusion >>
rect 284 215 285 216 
<< pdiffusion >>
rect 285 215 286 216 
<< pdiffusion >>
rect 286 215 287 216 
<< pdiffusion >>
rect 287 215 288 216 
<< m1 >>
rect 289 215 290 216 
<< m1 >>
rect 298 215 299 216 
<< m2 >>
rect 298 215 299 216 
<< pdiffusion >>
rect 300 215 301 216 
<< m1 >>
rect 301 215 302 216 
<< pdiffusion >>
rect 301 215 302 216 
<< pdiffusion >>
rect 302 215 303 216 
<< pdiffusion >>
rect 303 215 304 216 
<< pdiffusion >>
rect 304 215 305 216 
<< pdiffusion >>
rect 305 215 306 216 
<< m1 >>
rect 307 215 308 216 
<< m2 >>
rect 308 215 309 216 
<< m1 >>
rect 311 215 312 216 
<< pdiffusion >>
rect 318 215 319 216 
<< pdiffusion >>
rect 319 215 320 216 
<< pdiffusion >>
rect 320 215 321 216 
<< pdiffusion >>
rect 321 215 322 216 
<< pdiffusion >>
rect 322 215 323 216 
<< pdiffusion >>
rect 323 215 324 216 
<< pdiffusion >>
rect 336 215 337 216 
<< pdiffusion >>
rect 337 215 338 216 
<< pdiffusion >>
rect 338 215 339 216 
<< pdiffusion >>
rect 339 215 340 216 
<< m1 >>
rect 340 215 341 216 
<< pdiffusion >>
rect 340 215 341 216 
<< pdiffusion >>
rect 341 215 342 216 
<< pdiffusion >>
rect 354 215 355 216 
<< pdiffusion >>
rect 355 215 356 216 
<< pdiffusion >>
rect 356 215 357 216 
<< pdiffusion >>
rect 357 215 358 216 
<< pdiffusion >>
rect 358 215 359 216 
<< pdiffusion >>
rect 359 215 360 216 
<< pdiffusion >>
rect 372 215 373 216 
<< pdiffusion >>
rect 373 215 374 216 
<< pdiffusion >>
rect 374 215 375 216 
<< pdiffusion >>
rect 375 215 376 216 
<< pdiffusion >>
rect 376 215 377 216 
<< pdiffusion >>
rect 377 215 378 216 
<< pdiffusion >>
rect 390 215 391 216 
<< pdiffusion >>
rect 391 215 392 216 
<< pdiffusion >>
rect 392 215 393 216 
<< pdiffusion >>
rect 393 215 394 216 
<< pdiffusion >>
rect 394 215 395 216 
<< pdiffusion >>
rect 395 215 396 216 
<< pdiffusion >>
rect 408 215 409 216 
<< pdiffusion >>
rect 409 215 410 216 
<< pdiffusion >>
rect 410 215 411 216 
<< pdiffusion >>
rect 411 215 412 216 
<< pdiffusion >>
rect 412 215 413 216 
<< pdiffusion >>
rect 413 215 414 216 
<< pdiffusion >>
rect 426 215 427 216 
<< pdiffusion >>
rect 427 215 428 216 
<< pdiffusion >>
rect 428 215 429 216 
<< pdiffusion >>
rect 429 215 430 216 
<< pdiffusion >>
rect 430 215 431 216 
<< pdiffusion >>
rect 431 215 432 216 
<< pdiffusion >>
rect 444 215 445 216 
<< pdiffusion >>
rect 445 215 446 216 
<< pdiffusion >>
rect 446 215 447 216 
<< pdiffusion >>
rect 447 215 448 216 
<< pdiffusion >>
rect 448 215 449 216 
<< pdiffusion >>
rect 449 215 450 216 
<< m1 >>
rect 451 215 452 216 
<< m1 >>
rect 19 216 20 217 
<< m1 >>
rect 49 216 50 217 
<< m2 >>
rect 117 216 118 217 
<< m1 >>
rect 118 216 119 217 
<< m1 >>
rect 121 216 122 217 
<< m1 >>
rect 127 216 128 217 
<< m1 >>
rect 142 216 143 217 
<< m1 >>
rect 154 216 155 217 
<< m1 >>
rect 178 216 179 217 
<< m2 >>
rect 181 216 182 217 
<< m1 >>
rect 190 216 191 217 
<< m1 >>
rect 196 216 197 217 
<< m1 >>
rect 200 216 201 217 
<< m1 >>
rect 207 216 208 217 
<< m1 >>
rect 235 216 236 217 
<< m1 >>
rect 237 216 238 217 
<< m1 >>
rect 244 216 245 217 
<< m1 >>
rect 268 216 269 217 
<< m1 >>
rect 289 216 290 217 
<< m1 >>
rect 298 216 299 217 
<< m2 >>
rect 298 216 299 217 
<< m1 >>
rect 301 216 302 217 
<< m1 >>
rect 307 216 308 217 
<< m2 >>
rect 308 216 309 217 
<< m1 >>
rect 311 216 312 217 
<< m1 >>
rect 340 216 341 217 
<< m1 >>
rect 451 216 452 217 
<< m1 >>
rect 19 217 20 218 
<< m1 >>
rect 49 217 50 218 
<< m2 >>
rect 117 217 118 218 
<< m1 >>
rect 118 217 119 218 
<< m2 >>
rect 118 217 119 218 
<< m2 >>
rect 119 217 120 218 
<< m1 >>
rect 120 217 121 218 
<< m2 >>
rect 120 217 121 218 
<< m2c >>
rect 120 217 121 218 
<< m1 >>
rect 120 217 121 218 
<< m2 >>
rect 120 217 121 218 
<< m1 >>
rect 121 217 122 218 
<< m1 >>
rect 127 217 128 218 
<< m1 >>
rect 142 217 143 218 
<< m1 >>
rect 154 217 155 218 
<< m1 >>
rect 178 217 179 218 
<< m1 >>
rect 179 217 180 218 
<< m1 >>
rect 180 217 181 218 
<< m1 >>
rect 181 217 182 218 
<< m2 >>
rect 181 217 182 218 
<< m1 >>
rect 182 217 183 218 
<< m1 >>
rect 183 217 184 218 
<< m1 >>
rect 184 217 185 218 
<< m1 >>
rect 185 217 186 218 
<< m1 >>
rect 186 217 187 218 
<< m1 >>
rect 187 217 188 218 
<< m1 >>
rect 188 217 189 218 
<< m2 >>
rect 188 217 189 218 
<< m2c >>
rect 188 217 189 218 
<< m1 >>
rect 188 217 189 218 
<< m2 >>
rect 188 217 189 218 
<< m2 >>
rect 189 217 190 218 
<< m1 >>
rect 190 217 191 218 
<< m2 >>
rect 190 217 191 218 
<< m2 >>
rect 191 217 192 218 
<< m1 >>
rect 192 217 193 218 
<< m2 >>
rect 192 217 193 218 
<< m2c >>
rect 192 217 193 218 
<< m1 >>
rect 192 217 193 218 
<< m2 >>
rect 192 217 193 218 
<< m1 >>
rect 196 217 197 218 
<< m1 >>
rect 200 217 201 218 
<< m1 >>
rect 207 217 208 218 
<< m1 >>
rect 235 217 236 218 
<< m1 >>
rect 237 217 238 218 
<< m1 >>
rect 244 217 245 218 
<< m1 >>
rect 268 217 269 218 
<< m1 >>
rect 289 217 290 218 
<< m1 >>
rect 298 217 299 218 
<< m2 >>
rect 298 217 299 218 
<< m1 >>
rect 299 217 300 218 
<< m1 >>
rect 300 217 301 218 
<< m1 >>
rect 301 217 302 218 
<< m1 >>
rect 307 217 308 218 
<< m2 >>
rect 308 217 309 218 
<< m1 >>
rect 311 217 312 218 
<< m1 >>
rect 340 217 341 218 
<< m1 >>
rect 451 217 452 218 
<< m1 >>
rect 19 218 20 219 
<< m1 >>
rect 49 218 50 219 
<< m1 >>
rect 118 218 119 219 
<< m1 >>
rect 127 218 128 219 
<< m1 >>
rect 142 218 143 219 
<< m1 >>
rect 154 218 155 219 
<< m2 >>
rect 154 218 155 219 
<< m2c >>
rect 154 218 155 219 
<< m1 >>
rect 154 218 155 219 
<< m2 >>
rect 154 218 155 219 
<< m2 >>
rect 181 218 182 219 
<< m1 >>
rect 190 218 191 219 
<< m1 >>
rect 192 218 193 219 
<< m1 >>
rect 196 218 197 219 
<< m1 >>
rect 200 218 201 219 
<< m1 >>
rect 207 218 208 219 
<< m1 >>
rect 235 218 236 219 
<< m1 >>
rect 237 218 238 219 
<< m1 >>
rect 244 218 245 219 
<< m1 >>
rect 268 218 269 219 
<< m1 >>
rect 289 218 290 219 
<< m2 >>
rect 298 218 299 219 
<< m1 >>
rect 307 218 308 219 
<< m2 >>
rect 308 218 309 219 
<< m1 >>
rect 311 218 312 219 
<< m1 >>
rect 340 218 341 219 
<< m1 >>
rect 448 218 449 219 
<< m1 >>
rect 449 218 450 219 
<< m1 >>
rect 450 218 451 219 
<< m1 >>
rect 451 218 452 219 
<< m1 >>
rect 19 219 20 220 
<< m1 >>
rect 49 219 50 220 
<< m1 >>
rect 118 219 119 220 
<< m1 >>
rect 127 219 128 220 
<< m1 >>
rect 142 219 143 220 
<< m2 >>
rect 154 219 155 220 
<< m2 >>
rect 181 219 182 220 
<< m1 >>
rect 190 219 191 220 
<< m1 >>
rect 192 219 193 220 
<< m2 >>
rect 195 219 196 220 
<< m1 >>
rect 196 219 197 220 
<< m2 >>
rect 196 219 197 220 
<< m2 >>
rect 197 219 198 220 
<< m1 >>
rect 198 219 199 220 
<< m2 >>
rect 198 219 199 220 
<< m2c >>
rect 198 219 199 220 
<< m1 >>
rect 198 219 199 220 
<< m2 >>
rect 198 219 199 220 
<< m1 >>
rect 199 219 200 220 
<< m1 >>
rect 200 219 201 220 
<< m1 >>
rect 207 219 208 220 
<< m1 >>
rect 235 219 236 220 
<< m1 >>
rect 237 219 238 220 
<< m1 >>
rect 244 219 245 220 
<< m1 >>
rect 268 219 269 220 
<< m1 >>
rect 289 219 290 220 
<< m1 >>
rect 298 219 299 220 
<< m2 >>
rect 298 219 299 220 
<< m2c >>
rect 298 219 299 220 
<< m1 >>
rect 298 219 299 220 
<< m2 >>
rect 298 219 299 220 
<< m1 >>
rect 307 219 308 220 
<< m2 >>
rect 308 219 309 220 
<< m1 >>
rect 311 219 312 220 
<< m1 >>
rect 340 219 341 220 
<< m1 >>
rect 448 219 449 220 
<< m1 >>
rect 19 220 20 221 
<< m1 >>
rect 49 220 50 221 
<< m1 >>
rect 118 220 119 221 
<< m1 >>
rect 127 220 128 221 
<< m1 >>
rect 142 220 143 221 
<< m1 >>
rect 143 220 144 221 
<< m1 >>
rect 144 220 145 221 
<< m1 >>
rect 145 220 146 221 
<< m1 >>
rect 146 220 147 221 
<< m1 >>
rect 147 220 148 221 
<< m1 >>
rect 148 220 149 221 
<< m1 >>
rect 149 220 150 221 
<< m1 >>
rect 150 220 151 221 
<< m1 >>
rect 151 220 152 221 
<< m1 >>
rect 152 220 153 221 
<< m1 >>
rect 153 220 154 221 
<< m1 >>
rect 154 220 155 221 
<< m2 >>
rect 154 220 155 221 
<< m1 >>
rect 155 220 156 221 
<< m1 >>
rect 156 220 157 221 
<< m1 >>
rect 157 220 158 221 
<< m1 >>
rect 158 220 159 221 
<< m1 >>
rect 159 220 160 221 
<< m1 >>
rect 160 220 161 221 
<< m1 >>
rect 161 220 162 221 
<< m1 >>
rect 162 220 163 221 
<< m1 >>
rect 163 220 164 221 
<< m1 >>
rect 164 220 165 221 
<< m1 >>
rect 165 220 166 221 
<< m1 >>
rect 166 220 167 221 
<< m1 >>
rect 167 220 168 221 
<< m1 >>
rect 168 220 169 221 
<< m1 >>
rect 169 220 170 221 
<< m1 >>
rect 170 220 171 221 
<< m1 >>
rect 171 220 172 221 
<< m1 >>
rect 172 220 173 221 
<< m1 >>
rect 173 220 174 221 
<< m1 >>
rect 174 220 175 221 
<< m1 >>
rect 175 220 176 221 
<< m1 >>
rect 176 220 177 221 
<< m1 >>
rect 177 220 178 221 
<< m1 >>
rect 178 220 179 221 
<< m1 >>
rect 179 220 180 221 
<< m1 >>
rect 180 220 181 221 
<< m1 >>
rect 181 220 182 221 
<< m2 >>
rect 181 220 182 221 
<< m1 >>
rect 182 220 183 221 
<< m1 >>
rect 183 220 184 221 
<< m1 >>
rect 184 220 185 221 
<< m1 >>
rect 185 220 186 221 
<< m1 >>
rect 186 220 187 221 
<< m1 >>
rect 187 220 188 221 
<< m1 >>
rect 188 220 189 221 
<< m2 >>
rect 188 220 189 221 
<< m2c >>
rect 188 220 189 221 
<< m1 >>
rect 188 220 189 221 
<< m2 >>
rect 188 220 189 221 
<< m2 >>
rect 189 220 190 221 
<< m1 >>
rect 190 220 191 221 
<< m2 >>
rect 190 220 191 221 
<< m2 >>
rect 191 220 192 221 
<< m1 >>
rect 192 220 193 221 
<< m2 >>
rect 192 220 193 221 
<< m2 >>
rect 193 220 194 221 
<< m1 >>
rect 194 220 195 221 
<< m2 >>
rect 194 220 195 221 
<< m2c >>
rect 194 220 195 221 
<< m1 >>
rect 194 220 195 221 
<< m2 >>
rect 194 220 195 221 
<< m2 >>
rect 195 220 196 221 
<< m1 >>
rect 196 220 197 221 
<< m1 >>
rect 207 220 208 221 
<< m1 >>
rect 235 220 236 221 
<< m1 >>
rect 237 220 238 221 
<< m1 >>
rect 244 220 245 221 
<< m1 >>
rect 268 220 269 221 
<< m1 >>
rect 269 220 270 221 
<< m1 >>
rect 270 220 271 221 
<< m1 >>
rect 271 220 272 221 
<< m1 >>
rect 272 220 273 221 
<< m1 >>
rect 273 220 274 221 
<< m1 >>
rect 274 220 275 221 
<< m1 >>
rect 275 220 276 221 
<< m1 >>
rect 276 220 277 221 
<< m1 >>
rect 277 220 278 221 
<< m1 >>
rect 278 220 279 221 
<< m1 >>
rect 279 220 280 221 
<< m1 >>
rect 280 220 281 221 
<< m1 >>
rect 281 220 282 221 
<< m1 >>
rect 282 220 283 221 
<< m1 >>
rect 283 220 284 221 
<< m2 >>
rect 283 220 284 221 
<< m2c >>
rect 283 220 284 221 
<< m1 >>
rect 283 220 284 221 
<< m2 >>
rect 283 220 284 221 
<< m1 >>
rect 289 220 290 221 
<< m2 >>
rect 289 220 290 221 
<< m2c >>
rect 289 220 290 221 
<< m1 >>
rect 289 220 290 221 
<< m2 >>
rect 289 220 290 221 
<< m1 >>
rect 298 220 299 221 
<< m1 >>
rect 307 220 308 221 
<< m2 >>
rect 308 220 309 221 
<< m1 >>
rect 311 220 312 221 
<< m1 >>
rect 340 220 341 221 
<< m1 >>
rect 448 220 449 221 
<< m1 >>
rect 19 221 20 222 
<< m1 >>
rect 49 221 50 222 
<< m1 >>
rect 118 221 119 222 
<< m1 >>
rect 127 221 128 222 
<< m2 >>
rect 154 221 155 222 
<< m2 >>
rect 181 221 182 222 
<< m1 >>
rect 190 221 191 222 
<< m1 >>
rect 192 221 193 222 
<< m1 >>
rect 196 221 197 222 
<< m1 >>
rect 197 221 198 222 
<< m1 >>
rect 198 221 199 222 
<< m1 >>
rect 199 221 200 222 
<< m1 >>
rect 200 221 201 222 
<< m1 >>
rect 201 221 202 222 
<< m1 >>
rect 202 221 203 222 
<< m1 >>
rect 203 221 204 222 
<< m2 >>
rect 203 221 204 222 
<< m2c >>
rect 203 221 204 222 
<< m1 >>
rect 203 221 204 222 
<< m2 >>
rect 203 221 204 222 
<< m1 >>
rect 207 221 208 222 
<< m2 >>
rect 207 221 208 222 
<< m2c >>
rect 207 221 208 222 
<< m1 >>
rect 207 221 208 222 
<< m2 >>
rect 207 221 208 222 
<< m1 >>
rect 235 221 236 222 
<< m2 >>
rect 235 221 236 222 
<< m2c >>
rect 235 221 236 222 
<< m1 >>
rect 235 221 236 222 
<< m2 >>
rect 235 221 236 222 
<< m1 >>
rect 237 221 238 222 
<< m2 >>
rect 237 221 238 222 
<< m2c >>
rect 237 221 238 222 
<< m1 >>
rect 237 221 238 222 
<< m2 >>
rect 237 221 238 222 
<< m1 >>
rect 244 221 245 222 
<< m2 >>
rect 283 221 284 222 
<< m2 >>
rect 289 221 290 222 
<< m2 >>
rect 290 221 291 222 
<< m2 >>
rect 291 221 292 222 
<< m2 >>
rect 292 221 293 222 
<< m2 >>
rect 293 221 294 222 
<< m2 >>
rect 294 221 295 222 
<< m2 >>
rect 295 221 296 222 
<< m2 >>
rect 296 221 297 222 
<< m2 >>
rect 297 221 298 222 
<< m1 >>
rect 298 221 299 222 
<< m2 >>
rect 298 221 299 222 
<< m2 >>
rect 299 221 300 222 
<< m1 >>
rect 300 221 301 222 
<< m2 >>
rect 300 221 301 222 
<< m2c >>
rect 300 221 301 222 
<< m1 >>
rect 300 221 301 222 
<< m2 >>
rect 300 221 301 222 
<< m1 >>
rect 301 221 302 222 
<< m1 >>
rect 302 221 303 222 
<< m1 >>
rect 303 221 304 222 
<< m1 >>
rect 304 221 305 222 
<< m1 >>
rect 305 221 306 222 
<< m2 >>
rect 305 221 306 222 
<< m2c >>
rect 305 221 306 222 
<< m1 >>
rect 305 221 306 222 
<< m2 >>
rect 305 221 306 222 
<< m2 >>
rect 306 221 307 222 
<< m1 >>
rect 307 221 308 222 
<< m2 >>
rect 308 221 309 222 
<< m1 >>
rect 311 221 312 222 
<< m2 >>
rect 311 221 312 222 
<< m2c >>
rect 311 221 312 222 
<< m1 >>
rect 311 221 312 222 
<< m2 >>
rect 311 221 312 222 
<< m1 >>
rect 340 221 341 222 
<< m1 >>
rect 448 221 449 222 
<< m1 >>
rect 19 222 20 223 
<< m1 >>
rect 49 222 50 223 
<< m1 >>
rect 118 222 119 223 
<< m1 >>
rect 127 222 128 223 
<< m1 >>
rect 154 222 155 223 
<< m2 >>
rect 154 222 155 223 
<< m2c >>
rect 154 222 155 223 
<< m1 >>
rect 154 222 155 223 
<< m2 >>
rect 154 222 155 223 
<< m1 >>
rect 174 222 175 223 
<< m1 >>
rect 175 222 176 223 
<< m1 >>
rect 176 222 177 223 
<< m1 >>
rect 177 222 178 223 
<< m1 >>
rect 178 222 179 223 
<< m1 >>
rect 179 222 180 223 
<< m1 >>
rect 180 222 181 223 
<< m1 >>
rect 181 222 182 223 
<< m2 >>
rect 181 222 182 223 
<< m2c >>
rect 181 222 182 223 
<< m1 >>
rect 181 222 182 223 
<< m2 >>
rect 181 222 182 223 
<< m1 >>
rect 190 222 191 223 
<< m1 >>
rect 192 222 193 223 
<< m2 >>
rect 203 222 204 223 
<< m2 >>
rect 207 222 208 223 
<< m2 >>
rect 208 222 209 223 
<< m2 >>
rect 209 222 210 223 
<< m2 >>
rect 210 222 211 223 
<< m2 >>
rect 211 222 212 223 
<< m2 >>
rect 212 222 213 223 
<< m2 >>
rect 213 222 214 223 
<< m2 >>
rect 214 222 215 223 
<< m2 >>
rect 215 222 216 223 
<< m2 >>
rect 216 222 217 223 
<< m2 >>
rect 217 222 218 223 
<< m2 >>
rect 218 222 219 223 
<< m2 >>
rect 219 222 220 223 
<< m2 >>
rect 220 222 221 223 
<< m2 >>
rect 221 222 222 223 
<< m2 >>
rect 222 222 223 223 
<< m2 >>
rect 223 222 224 223 
<< m2 >>
rect 224 222 225 223 
<< m2 >>
rect 225 222 226 223 
<< m2 >>
rect 226 222 227 223 
<< m2 >>
rect 227 222 228 223 
<< m2 >>
rect 228 222 229 223 
<< m2 >>
rect 229 222 230 223 
<< m2 >>
rect 230 222 231 223 
<< m2 >>
rect 235 222 236 223 
<< m2 >>
rect 237 222 238 223 
<< m1 >>
rect 244 222 245 223 
<< m2 >>
rect 269 222 270 223 
<< m1 >>
rect 270 222 271 223 
<< m2 >>
rect 270 222 271 223 
<< m2c >>
rect 270 222 271 223 
<< m1 >>
rect 270 222 271 223 
<< m2 >>
rect 270 222 271 223 
<< m1 >>
rect 271 222 272 223 
<< m1 >>
rect 272 222 273 223 
<< m1 >>
rect 273 222 274 223 
<< m1 >>
rect 274 222 275 223 
<< m1 >>
rect 275 222 276 223 
<< m1 >>
rect 276 222 277 223 
<< m1 >>
rect 277 222 278 223 
<< m1 >>
rect 278 222 279 223 
<< m1 >>
rect 279 222 280 223 
<< m1 >>
rect 280 222 281 223 
<< m1 >>
rect 281 222 282 223 
<< m1 >>
rect 282 222 283 223 
<< m1 >>
rect 283 222 284 223 
<< m2 >>
rect 283 222 284 223 
<< m1 >>
rect 284 222 285 223 
<< m1 >>
rect 285 222 286 223 
<< m1 >>
rect 286 222 287 223 
<< m1 >>
rect 287 222 288 223 
<< m1 >>
rect 288 222 289 223 
<< m1 >>
rect 289 222 290 223 
<< m1 >>
rect 290 222 291 223 
<< m1 >>
rect 291 222 292 223 
<< m1 >>
rect 292 222 293 223 
<< m1 >>
rect 293 222 294 223 
<< m1 >>
rect 294 222 295 223 
<< m1 >>
rect 295 222 296 223 
<< m1 >>
rect 296 222 297 223 
<< m1 >>
rect 297 222 298 223 
<< m1 >>
rect 298 222 299 223 
<< m2 >>
rect 306 222 307 223 
<< m1 >>
rect 307 222 308 223 
<< m2 >>
rect 308 222 309 223 
<< m2 >>
rect 311 222 312 223 
<< m1 >>
rect 340 222 341 223 
<< m1 >>
rect 448 222 449 223 
<< m1 >>
rect 19 223 20 224 
<< m1 >>
rect 49 223 50 224 
<< m1 >>
rect 50 223 51 224 
<< m1 >>
rect 51 223 52 224 
<< m1 >>
rect 52 223 53 224 
<< m1 >>
rect 53 223 54 224 
<< m1 >>
rect 54 223 55 224 
<< m1 >>
rect 55 223 56 224 
<< m1 >>
rect 56 223 57 224 
<< m1 >>
rect 57 223 58 224 
<< m1 >>
rect 58 223 59 224 
<< m1 >>
rect 59 223 60 224 
<< m1 >>
rect 60 223 61 224 
<< m1 >>
rect 61 223 62 224 
<< m1 >>
rect 62 223 63 224 
<< m1 >>
rect 63 223 64 224 
<< m1 >>
rect 64 223 65 224 
<< m1 >>
rect 118 223 119 224 
<< m1 >>
rect 127 223 128 224 
<< m1 >>
rect 154 223 155 224 
<< m1 >>
rect 174 223 175 224 
<< m1 >>
rect 190 223 191 224 
<< m1 >>
rect 192 223 193 224 
<< m1 >>
rect 193 223 194 224 
<< m1 >>
rect 194 223 195 224 
<< m1 >>
rect 195 223 196 224 
<< m1 >>
rect 196 223 197 224 
<< m1 >>
rect 197 223 198 224 
<< m1 >>
rect 198 223 199 224 
<< m1 >>
rect 199 223 200 224 
<< m1 >>
rect 200 223 201 224 
<< m1 >>
rect 201 223 202 224 
<< m1 >>
rect 202 223 203 224 
<< m1 >>
rect 203 223 204 224 
<< m2 >>
rect 203 223 204 224 
<< m1 >>
rect 204 223 205 224 
<< m1 >>
rect 205 223 206 224 
<< m2 >>
rect 205 223 206 224 
<< m2c >>
rect 205 223 206 224 
<< m1 >>
rect 205 223 206 224 
<< m2 >>
rect 205 223 206 224 
<< m2 >>
rect 206 223 207 224 
<< m2 >>
rect 207 223 208 224 
<< m1 >>
rect 208 223 209 224 
<< m1 >>
rect 209 223 210 224 
<< m1 >>
rect 210 223 211 224 
<< m1 >>
rect 211 223 212 224 
<< m1 >>
rect 212 223 213 224 
<< m1 >>
rect 213 223 214 224 
<< m1 >>
rect 214 223 215 224 
<< m1 >>
rect 215 223 216 224 
<< m1 >>
rect 216 223 217 224 
<< m1 >>
rect 217 223 218 224 
<< m1 >>
rect 218 223 219 224 
<< m1 >>
rect 219 223 220 224 
<< m1 >>
rect 220 223 221 224 
<< m1 >>
rect 221 223 222 224 
<< m1 >>
rect 222 223 223 224 
<< m1 >>
rect 223 223 224 224 
<< m1 >>
rect 224 223 225 224 
<< m1 >>
rect 225 223 226 224 
<< m1 >>
rect 226 223 227 224 
<< m1 >>
rect 227 223 228 224 
<< m1 >>
rect 228 223 229 224 
<< m1 >>
rect 229 223 230 224 
<< m1 >>
rect 230 223 231 224 
<< m2 >>
rect 230 223 231 224 
<< m1 >>
rect 231 223 232 224 
<< m1 >>
rect 232 223 233 224 
<< m1 >>
rect 233 223 234 224 
<< m1 >>
rect 234 223 235 224 
<< m1 >>
rect 235 223 236 224 
<< m2 >>
rect 235 223 236 224 
<< m1 >>
rect 236 223 237 224 
<< m1 >>
rect 237 223 238 224 
<< m2 >>
rect 237 223 238 224 
<< m1 >>
rect 238 223 239 224 
<< m1 >>
rect 239 223 240 224 
<< m1 >>
rect 240 223 241 224 
<< m1 >>
rect 241 223 242 224 
<< m1 >>
rect 242 223 243 224 
<< m2 >>
rect 242 223 243 224 
<< m2c >>
rect 242 223 243 224 
<< m1 >>
rect 242 223 243 224 
<< m2 >>
rect 242 223 243 224 
<< m2 >>
rect 243 223 244 224 
<< m1 >>
rect 244 223 245 224 
<< m2 >>
rect 244 223 245 224 
<< m2 >>
rect 245 223 246 224 
<< m1 >>
rect 246 223 247 224 
<< m2 >>
rect 246 223 247 224 
<< m2c >>
rect 246 223 247 224 
<< m1 >>
rect 246 223 247 224 
<< m2 >>
rect 246 223 247 224 
<< m1 >>
rect 247 223 248 224 
<< m1 >>
rect 248 223 249 224 
<< m1 >>
rect 249 223 250 224 
<< m1 >>
rect 250 223 251 224 
<< m1 >>
rect 251 223 252 224 
<< m1 >>
rect 252 223 253 224 
<< m1 >>
rect 253 223 254 224 
<< m1 >>
rect 254 223 255 224 
<< m1 >>
rect 255 223 256 224 
<< m1 >>
rect 256 223 257 224 
<< m1 >>
rect 257 223 258 224 
<< m1 >>
rect 258 223 259 224 
<< m1 >>
rect 259 223 260 224 
<< m1 >>
rect 260 223 261 224 
<< m1 >>
rect 261 223 262 224 
<< m1 >>
rect 262 223 263 224 
<< m1 >>
rect 263 223 264 224 
<< m1 >>
rect 264 223 265 224 
<< m1 >>
rect 265 223 266 224 
<< m1 >>
rect 266 223 267 224 
<< m1 >>
rect 267 223 268 224 
<< m1 >>
rect 268 223 269 224 
<< m2 >>
rect 269 223 270 224 
<< m2 >>
rect 283 223 284 224 
<< m2 >>
rect 306 223 307 224 
<< m1 >>
rect 307 223 308 224 
<< m2 >>
rect 308 223 309 224 
<< m1 >>
rect 309 223 310 224 
<< m2 >>
rect 309 223 310 224 
<< m2c >>
rect 309 223 310 224 
<< m1 >>
rect 309 223 310 224 
<< m2 >>
rect 309 223 310 224 
<< m1 >>
rect 310 223 311 224 
<< m1 >>
rect 311 223 312 224 
<< m2 >>
rect 311 223 312 224 
<< m1 >>
rect 312 223 313 224 
<< m1 >>
rect 313 223 314 224 
<< m2 >>
rect 313 223 314 224 
<< m1 >>
rect 314 223 315 224 
<< m2 >>
rect 314 223 315 224 
<< m1 >>
rect 315 223 316 224 
<< m2 >>
rect 315 223 316 224 
<< m1 >>
rect 316 223 317 224 
<< m2 >>
rect 316 223 317 224 
<< m1 >>
rect 317 223 318 224 
<< m2 >>
rect 317 223 318 224 
<< m1 >>
rect 318 223 319 224 
<< m2 >>
rect 318 223 319 224 
<< m1 >>
rect 319 223 320 224 
<< m2 >>
rect 319 223 320 224 
<< m1 >>
rect 320 223 321 224 
<< m2 >>
rect 320 223 321 224 
<< m1 >>
rect 321 223 322 224 
<< m2 >>
rect 321 223 322 224 
<< m1 >>
rect 322 223 323 224 
<< m2 >>
rect 322 223 323 224 
<< m1 >>
rect 323 223 324 224 
<< m2 >>
rect 323 223 324 224 
<< m1 >>
rect 324 223 325 224 
<< m2 >>
rect 324 223 325 224 
<< m1 >>
rect 325 223 326 224 
<< m2 >>
rect 325 223 326 224 
<< m1 >>
rect 326 223 327 224 
<< m2 >>
rect 326 223 327 224 
<< m1 >>
rect 327 223 328 224 
<< m2 >>
rect 327 223 328 224 
<< m1 >>
rect 328 223 329 224 
<< m2 >>
rect 328 223 329 224 
<< m1 >>
rect 329 223 330 224 
<< m2 >>
rect 329 223 330 224 
<< m1 >>
rect 330 223 331 224 
<< m2 >>
rect 330 223 331 224 
<< m1 >>
rect 331 223 332 224 
<< m2 >>
rect 331 223 332 224 
<< m1 >>
rect 332 223 333 224 
<< m2 >>
rect 332 223 333 224 
<< m1 >>
rect 333 223 334 224 
<< m2 >>
rect 333 223 334 224 
<< m1 >>
rect 334 223 335 224 
<< m2 >>
rect 334 223 335 224 
<< m1 >>
rect 335 223 336 224 
<< m2 >>
rect 335 223 336 224 
<< m1 >>
rect 336 223 337 224 
<< m2 >>
rect 336 223 337 224 
<< m1 >>
rect 337 223 338 224 
<< m2 >>
rect 337 223 338 224 
<< m2 >>
rect 338 223 339 224 
<< m2 >>
rect 339 223 340 224 
<< m1 >>
rect 340 223 341 224 
<< m2 >>
rect 340 223 341 224 
<< m2 >>
rect 341 223 342 224 
<< m1 >>
rect 342 223 343 224 
<< m2 >>
rect 342 223 343 224 
<< m2c >>
rect 342 223 343 224 
<< m1 >>
rect 342 223 343 224 
<< m2 >>
rect 342 223 343 224 
<< m1 >>
rect 343 223 344 224 
<< m1 >>
rect 344 223 345 224 
<< m1 >>
rect 345 223 346 224 
<< m1 >>
rect 346 223 347 224 
<< m1 >>
rect 347 223 348 224 
<< m1 >>
rect 348 223 349 224 
<< m1 >>
rect 349 223 350 224 
<< m1 >>
rect 350 223 351 224 
<< m1 >>
rect 351 223 352 224 
<< m1 >>
rect 352 223 353 224 
<< m1 >>
rect 353 223 354 224 
<< m1 >>
rect 354 223 355 224 
<< m1 >>
rect 355 223 356 224 
<< m1 >>
rect 356 223 357 224 
<< m1 >>
rect 357 223 358 224 
<< m1 >>
rect 358 223 359 224 
<< m1 >>
rect 359 223 360 224 
<< m1 >>
rect 360 223 361 224 
<< m1 >>
rect 361 223 362 224 
<< m1 >>
rect 362 223 363 224 
<< m1 >>
rect 363 223 364 224 
<< m1 >>
rect 364 223 365 224 
<< m1 >>
rect 365 223 366 224 
<< m1 >>
rect 366 223 367 224 
<< m1 >>
rect 367 223 368 224 
<< m1 >>
rect 368 223 369 224 
<< m1 >>
rect 369 223 370 224 
<< m1 >>
rect 370 223 371 224 
<< m1 >>
rect 371 223 372 224 
<< m1 >>
rect 372 223 373 224 
<< m1 >>
rect 373 223 374 224 
<< m1 >>
rect 374 223 375 224 
<< m1 >>
rect 375 223 376 224 
<< m1 >>
rect 376 223 377 224 
<< m1 >>
rect 448 223 449 224 
<< m1 >>
rect 19 224 20 225 
<< m1 >>
rect 64 224 65 225 
<< m1 >>
rect 118 224 119 225 
<< m1 >>
rect 127 224 128 225 
<< m1 >>
rect 154 224 155 225 
<< m2 >>
rect 164 224 165 225 
<< m1 >>
rect 165 224 166 225 
<< m2 >>
rect 165 224 166 225 
<< m2c >>
rect 165 224 166 225 
<< m1 >>
rect 165 224 166 225 
<< m2 >>
rect 165 224 166 225 
<< m1 >>
rect 166 224 167 225 
<< m1 >>
rect 167 224 168 225 
<< m1 >>
rect 168 224 169 225 
<< m1 >>
rect 169 224 170 225 
<< m1 >>
rect 170 224 171 225 
<< m1 >>
rect 171 224 172 225 
<< m1 >>
rect 172 224 173 225 
<< m1 >>
rect 173 224 174 225 
<< m1 >>
rect 174 224 175 225 
<< m1 >>
rect 190 224 191 225 
<< m2 >>
rect 203 224 204 225 
<< m2 >>
rect 207 224 208 225 
<< m1 >>
rect 208 224 209 225 
<< m2 >>
rect 230 224 231 225 
<< m2 >>
rect 235 224 236 225 
<< m2 >>
rect 237 224 238 225 
<< m1 >>
rect 244 224 245 225 
<< m1 >>
rect 268 224 269 225 
<< m2 >>
rect 269 224 270 225 
<< m1 >>
rect 283 224 284 225 
<< m2 >>
rect 283 224 284 225 
<< m2c >>
rect 283 224 284 225 
<< m1 >>
rect 283 224 284 225 
<< m2 >>
rect 283 224 284 225 
<< m2 >>
rect 306 224 307 225 
<< m1 >>
rect 307 224 308 225 
<< m2 >>
rect 311 224 312 225 
<< m2 >>
rect 313 224 314 225 
<< m1 >>
rect 337 224 338 225 
<< m1 >>
rect 340 224 341 225 
<< m1 >>
rect 376 224 377 225 
<< m1 >>
rect 448 224 449 225 
<< m1 >>
rect 19 225 20 226 
<< m1 >>
rect 64 225 65 226 
<< m1 >>
rect 118 225 119 226 
<< m1 >>
rect 127 225 128 226 
<< m1 >>
rect 154 225 155 226 
<< m1 >>
rect 157 225 158 226 
<< m1 >>
rect 158 225 159 226 
<< m1 >>
rect 159 225 160 226 
<< m1 >>
rect 160 225 161 226 
<< m1 >>
rect 161 225 162 226 
<< m1 >>
rect 162 225 163 226 
<< m1 >>
rect 163 225 164 226 
<< m2 >>
rect 164 225 165 226 
<< m1 >>
rect 190 225 191 226 
<< m1 >>
rect 203 225 204 226 
<< m2 >>
rect 203 225 204 226 
<< m2c >>
rect 203 225 204 226 
<< m1 >>
rect 203 225 204 226 
<< m2 >>
rect 203 225 204 226 
<< m2 >>
rect 207 225 208 226 
<< m1 >>
rect 208 225 209 226 
<< m1 >>
rect 230 225 231 226 
<< m2 >>
rect 230 225 231 226 
<< m2c >>
rect 230 225 231 226 
<< m1 >>
rect 230 225 231 226 
<< m2 >>
rect 230 225 231 226 
<< m1 >>
rect 231 225 232 226 
<< m1 >>
rect 232 225 233 226 
<< m1 >>
rect 233 225 234 226 
<< m1 >>
rect 234 225 235 226 
<< m1 >>
rect 235 225 236 226 
<< m2 >>
rect 235 225 236 226 
<< m1 >>
rect 236 225 237 226 
<< m1 >>
rect 237 225 238 226 
<< m2 >>
rect 237 225 238 226 
<< m1 >>
rect 238 225 239 226 
<< m1 >>
rect 239 225 240 226 
<< m1 >>
rect 240 225 241 226 
<< m1 >>
rect 241 225 242 226 
<< m1 >>
rect 242 225 243 226 
<< m2 >>
rect 242 225 243 226 
<< m2c >>
rect 242 225 243 226 
<< m1 >>
rect 242 225 243 226 
<< m2 >>
rect 242 225 243 226 
<< m2 >>
rect 243 225 244 226 
<< m1 >>
rect 244 225 245 226 
<< m1 >>
rect 265 225 266 226 
<< m1 >>
rect 266 225 267 226 
<< m2 >>
rect 266 225 267 226 
<< m2c >>
rect 266 225 267 226 
<< m1 >>
rect 266 225 267 226 
<< m2 >>
rect 266 225 267 226 
<< m2 >>
rect 267 225 268 226 
<< m1 >>
rect 268 225 269 226 
<< m2 >>
rect 268 225 269 226 
<< m2 >>
rect 269 225 270 226 
<< m1 >>
rect 283 225 284 226 
<< m2 >>
rect 306 225 307 226 
<< m1 >>
rect 307 225 308 226 
<< m2 >>
rect 307 225 308 226 
<< m2 >>
rect 308 225 309 226 
<< m1 >>
rect 309 225 310 226 
<< m2 >>
rect 309 225 310 226 
<< m2c >>
rect 309 225 310 226 
<< m1 >>
rect 309 225 310 226 
<< m2 >>
rect 309 225 310 226 
<< m1 >>
rect 311 225 312 226 
<< m2 >>
rect 311 225 312 226 
<< m2c >>
rect 311 225 312 226 
<< m1 >>
rect 311 225 312 226 
<< m2 >>
rect 311 225 312 226 
<< m1 >>
rect 313 225 314 226 
<< m2 >>
rect 313 225 314 226 
<< m2c >>
rect 313 225 314 226 
<< m1 >>
rect 313 225 314 226 
<< m2 >>
rect 313 225 314 226 
<< m1 >>
rect 337 225 338 226 
<< m1 >>
rect 340 225 341 226 
<< m1 >>
rect 341 225 342 226 
<< m1 >>
rect 342 225 343 226 
<< m1 >>
rect 343 225 344 226 
<< m1 >>
rect 344 225 345 226 
<< m1 >>
rect 345 225 346 226 
<< m1 >>
rect 346 225 347 226 
<< m1 >>
rect 347 225 348 226 
<< m1 >>
rect 348 225 349 226 
<< m1 >>
rect 349 225 350 226 
<< m1 >>
rect 350 225 351 226 
<< m1 >>
rect 351 225 352 226 
<< m1 >>
rect 352 225 353 226 
<< m1 >>
rect 376 225 377 226 
<< m1 >>
rect 448 225 449 226 
<< m1 >>
rect 16 226 17 227 
<< m1 >>
rect 17 226 18 227 
<< m1 >>
rect 18 226 19 227 
<< m1 >>
rect 19 226 20 227 
<< m1 >>
rect 64 226 65 227 
<< m1 >>
rect 118 226 119 227 
<< m1 >>
rect 127 226 128 227 
<< m1 >>
rect 154 226 155 227 
<< m1 >>
rect 157 226 158 227 
<< m1 >>
rect 163 226 164 227 
<< m2 >>
rect 164 226 165 227 
<< m1 >>
rect 190 226 191 227 
<< m1 >>
rect 203 226 204 227 
<< m2 >>
rect 207 226 208 227 
<< m1 >>
rect 208 226 209 227 
<< m2 >>
rect 235 226 236 227 
<< m2 >>
rect 237 226 238 227 
<< m2 >>
rect 243 226 244 227 
<< m1 >>
rect 244 226 245 227 
<< m1 >>
rect 265 226 266 227 
<< m1 >>
rect 268 226 269 227 
<< m1 >>
rect 283 226 284 227 
<< m1 >>
rect 307 226 308 227 
<< m1 >>
rect 309 226 310 227 
<< m1 >>
rect 311 226 312 227 
<< m1 >>
rect 313 226 314 227 
<< m1 >>
rect 337 226 338 227 
<< m1 >>
rect 352 226 353 227 
<< m1 >>
rect 376 226 377 227 
<< m1 >>
rect 448 226 449 227 
<< m1 >>
rect 16 227 17 228 
<< m1 >>
rect 64 227 65 228 
<< m1 >>
rect 118 227 119 228 
<< m1 >>
rect 127 227 128 228 
<< m1 >>
rect 154 227 155 228 
<< m1 >>
rect 157 227 158 228 
<< m1 >>
rect 163 227 164 228 
<< m2 >>
rect 164 227 165 228 
<< m1 >>
rect 190 227 191 228 
<< m1 >>
rect 203 227 204 228 
<< m2 >>
rect 207 227 208 228 
<< m1 >>
rect 208 227 209 228 
<< m1 >>
rect 235 227 236 228 
<< m2 >>
rect 235 227 236 228 
<< m2c >>
rect 235 227 236 228 
<< m1 >>
rect 235 227 236 228 
<< m2 >>
rect 235 227 236 228 
<< m1 >>
rect 237 227 238 228 
<< m2 >>
rect 237 227 238 228 
<< m2c >>
rect 237 227 238 228 
<< m1 >>
rect 237 227 238 228 
<< m2 >>
rect 237 227 238 228 
<< m2 >>
rect 243 227 244 228 
<< m1 >>
rect 244 227 245 228 
<< m1 >>
rect 265 227 266 228 
<< m1 >>
rect 268 227 269 228 
<< m1 >>
rect 283 227 284 228 
<< m1 >>
rect 307 227 308 228 
<< m1 >>
rect 309 227 310 228 
<< m2 >>
rect 309 227 310 228 
<< m2c >>
rect 309 227 310 228 
<< m1 >>
rect 309 227 310 228 
<< m2 >>
rect 309 227 310 228 
<< m2 >>
rect 310 227 311 228 
<< m1 >>
rect 311 227 312 228 
<< m2 >>
rect 311 227 312 228 
<< m2 >>
rect 312 227 313 228 
<< m1 >>
rect 313 227 314 228 
<< m2 >>
rect 313 227 314 228 
<< m2c >>
rect 313 227 314 228 
<< m1 >>
rect 313 227 314 228 
<< m2 >>
rect 313 227 314 228 
<< m1 >>
rect 337 227 338 228 
<< m1 >>
rect 352 227 353 228 
<< m1 >>
rect 376 227 377 228 
<< m1 >>
rect 448 227 449 228 
<< pdiffusion >>
rect 12 228 13 229 
<< pdiffusion >>
rect 13 228 14 229 
<< pdiffusion >>
rect 14 228 15 229 
<< pdiffusion >>
rect 15 228 16 229 
<< m1 >>
rect 16 228 17 229 
<< pdiffusion >>
rect 16 228 17 229 
<< pdiffusion >>
rect 17 228 18 229 
<< pdiffusion >>
rect 30 228 31 229 
<< pdiffusion >>
rect 31 228 32 229 
<< pdiffusion >>
rect 32 228 33 229 
<< pdiffusion >>
rect 33 228 34 229 
<< pdiffusion >>
rect 34 228 35 229 
<< pdiffusion >>
rect 35 228 36 229 
<< pdiffusion >>
rect 48 228 49 229 
<< pdiffusion >>
rect 49 228 50 229 
<< pdiffusion >>
rect 50 228 51 229 
<< pdiffusion >>
rect 51 228 52 229 
<< pdiffusion >>
rect 52 228 53 229 
<< pdiffusion >>
rect 53 228 54 229 
<< m1 >>
rect 64 228 65 229 
<< pdiffusion >>
rect 66 228 67 229 
<< pdiffusion >>
rect 67 228 68 229 
<< pdiffusion >>
rect 68 228 69 229 
<< pdiffusion >>
rect 69 228 70 229 
<< pdiffusion >>
rect 70 228 71 229 
<< pdiffusion >>
rect 71 228 72 229 
<< pdiffusion >>
rect 84 228 85 229 
<< pdiffusion >>
rect 85 228 86 229 
<< pdiffusion >>
rect 86 228 87 229 
<< pdiffusion >>
rect 87 228 88 229 
<< pdiffusion >>
rect 88 228 89 229 
<< pdiffusion >>
rect 89 228 90 229 
<< pdiffusion >>
rect 102 228 103 229 
<< pdiffusion >>
rect 103 228 104 229 
<< pdiffusion >>
rect 104 228 105 229 
<< pdiffusion >>
rect 105 228 106 229 
<< pdiffusion >>
rect 106 228 107 229 
<< pdiffusion >>
rect 107 228 108 229 
<< m1 >>
rect 118 228 119 229 
<< pdiffusion >>
rect 120 228 121 229 
<< pdiffusion >>
rect 121 228 122 229 
<< pdiffusion >>
rect 122 228 123 229 
<< pdiffusion >>
rect 123 228 124 229 
<< pdiffusion >>
rect 124 228 125 229 
<< pdiffusion >>
rect 125 228 126 229 
<< m1 >>
rect 127 228 128 229 
<< pdiffusion >>
rect 138 228 139 229 
<< pdiffusion >>
rect 139 228 140 229 
<< pdiffusion >>
rect 140 228 141 229 
<< pdiffusion >>
rect 141 228 142 229 
<< pdiffusion >>
rect 142 228 143 229 
<< pdiffusion >>
rect 143 228 144 229 
<< m1 >>
rect 154 228 155 229 
<< pdiffusion >>
rect 156 228 157 229 
<< m1 >>
rect 157 228 158 229 
<< pdiffusion >>
rect 157 228 158 229 
<< pdiffusion >>
rect 158 228 159 229 
<< pdiffusion >>
rect 159 228 160 229 
<< pdiffusion >>
rect 160 228 161 229 
<< pdiffusion >>
rect 161 228 162 229 
<< m1 >>
rect 163 228 164 229 
<< m2 >>
rect 164 228 165 229 
<< pdiffusion >>
rect 174 228 175 229 
<< pdiffusion >>
rect 175 228 176 229 
<< pdiffusion >>
rect 176 228 177 229 
<< pdiffusion >>
rect 177 228 178 229 
<< pdiffusion >>
rect 178 228 179 229 
<< pdiffusion >>
rect 179 228 180 229 
<< m1 >>
rect 190 228 191 229 
<< pdiffusion >>
rect 192 228 193 229 
<< pdiffusion >>
rect 193 228 194 229 
<< pdiffusion >>
rect 194 228 195 229 
<< pdiffusion >>
rect 195 228 196 229 
<< pdiffusion >>
rect 196 228 197 229 
<< pdiffusion >>
rect 197 228 198 229 
<< m1 >>
rect 203 228 204 229 
<< m2 >>
rect 207 228 208 229 
<< m1 >>
rect 208 228 209 229 
<< pdiffusion >>
rect 210 228 211 229 
<< pdiffusion >>
rect 211 228 212 229 
<< pdiffusion >>
rect 212 228 213 229 
<< pdiffusion >>
rect 213 228 214 229 
<< pdiffusion >>
rect 214 228 215 229 
<< pdiffusion >>
rect 215 228 216 229 
<< pdiffusion >>
rect 228 228 229 229 
<< pdiffusion >>
rect 229 228 230 229 
<< pdiffusion >>
rect 230 228 231 229 
<< pdiffusion >>
rect 231 228 232 229 
<< pdiffusion >>
rect 232 228 233 229 
<< pdiffusion >>
rect 233 228 234 229 
<< m1 >>
rect 235 228 236 229 
<< m1 >>
rect 237 228 238 229 
<< m2 >>
rect 243 228 244 229 
<< m1 >>
rect 244 228 245 229 
<< pdiffusion >>
rect 246 228 247 229 
<< pdiffusion >>
rect 247 228 248 229 
<< pdiffusion >>
rect 248 228 249 229 
<< pdiffusion >>
rect 249 228 250 229 
<< pdiffusion >>
rect 250 228 251 229 
<< pdiffusion >>
rect 251 228 252 229 
<< pdiffusion >>
rect 264 228 265 229 
<< m1 >>
rect 265 228 266 229 
<< pdiffusion >>
rect 265 228 266 229 
<< pdiffusion >>
rect 266 228 267 229 
<< pdiffusion >>
rect 267 228 268 229 
<< m1 >>
rect 268 228 269 229 
<< pdiffusion >>
rect 268 228 269 229 
<< pdiffusion >>
rect 269 228 270 229 
<< pdiffusion >>
rect 282 228 283 229 
<< m1 >>
rect 283 228 284 229 
<< pdiffusion >>
rect 283 228 284 229 
<< pdiffusion >>
rect 284 228 285 229 
<< pdiffusion >>
rect 285 228 286 229 
<< pdiffusion >>
rect 286 228 287 229 
<< pdiffusion >>
rect 287 228 288 229 
<< pdiffusion >>
rect 300 228 301 229 
<< pdiffusion >>
rect 301 228 302 229 
<< pdiffusion >>
rect 302 228 303 229 
<< pdiffusion >>
rect 303 228 304 229 
<< pdiffusion >>
rect 304 228 305 229 
<< pdiffusion >>
rect 305 228 306 229 
<< m1 >>
rect 307 228 308 229 
<< m1 >>
rect 311 228 312 229 
<< pdiffusion >>
rect 318 228 319 229 
<< pdiffusion >>
rect 319 228 320 229 
<< pdiffusion >>
rect 320 228 321 229 
<< pdiffusion >>
rect 321 228 322 229 
<< pdiffusion >>
rect 322 228 323 229 
<< pdiffusion >>
rect 323 228 324 229 
<< pdiffusion >>
rect 336 228 337 229 
<< m1 >>
rect 337 228 338 229 
<< pdiffusion >>
rect 337 228 338 229 
<< pdiffusion >>
rect 338 228 339 229 
<< pdiffusion >>
rect 339 228 340 229 
<< pdiffusion >>
rect 340 228 341 229 
<< pdiffusion >>
rect 341 228 342 229 
<< m1 >>
rect 352 228 353 229 
<< pdiffusion >>
rect 354 228 355 229 
<< pdiffusion >>
rect 355 228 356 229 
<< pdiffusion >>
rect 356 228 357 229 
<< pdiffusion >>
rect 357 228 358 229 
<< pdiffusion >>
rect 358 228 359 229 
<< pdiffusion >>
rect 359 228 360 229 
<< pdiffusion >>
rect 372 228 373 229 
<< pdiffusion >>
rect 373 228 374 229 
<< pdiffusion >>
rect 374 228 375 229 
<< pdiffusion >>
rect 375 228 376 229 
<< m1 >>
rect 376 228 377 229 
<< pdiffusion >>
rect 376 228 377 229 
<< pdiffusion >>
rect 377 228 378 229 
<< pdiffusion >>
rect 390 228 391 229 
<< pdiffusion >>
rect 391 228 392 229 
<< pdiffusion >>
rect 392 228 393 229 
<< pdiffusion >>
rect 393 228 394 229 
<< pdiffusion >>
rect 394 228 395 229 
<< pdiffusion >>
rect 395 228 396 229 
<< pdiffusion >>
rect 408 228 409 229 
<< pdiffusion >>
rect 409 228 410 229 
<< pdiffusion >>
rect 410 228 411 229 
<< pdiffusion >>
rect 411 228 412 229 
<< pdiffusion >>
rect 412 228 413 229 
<< pdiffusion >>
rect 413 228 414 229 
<< pdiffusion >>
rect 426 228 427 229 
<< pdiffusion >>
rect 427 228 428 229 
<< pdiffusion >>
rect 428 228 429 229 
<< pdiffusion >>
rect 429 228 430 229 
<< pdiffusion >>
rect 430 228 431 229 
<< pdiffusion >>
rect 431 228 432 229 
<< pdiffusion >>
rect 444 228 445 229 
<< pdiffusion >>
rect 445 228 446 229 
<< pdiffusion >>
rect 446 228 447 229 
<< pdiffusion >>
rect 447 228 448 229 
<< m1 >>
rect 448 228 449 229 
<< pdiffusion >>
rect 448 228 449 229 
<< pdiffusion >>
rect 449 228 450 229 
<< pdiffusion >>
rect 12 229 13 230 
<< pdiffusion >>
rect 13 229 14 230 
<< pdiffusion >>
rect 14 229 15 230 
<< pdiffusion >>
rect 15 229 16 230 
<< pdiffusion >>
rect 16 229 17 230 
<< pdiffusion >>
rect 17 229 18 230 
<< pdiffusion >>
rect 30 229 31 230 
<< pdiffusion >>
rect 31 229 32 230 
<< pdiffusion >>
rect 32 229 33 230 
<< pdiffusion >>
rect 33 229 34 230 
<< pdiffusion >>
rect 34 229 35 230 
<< pdiffusion >>
rect 35 229 36 230 
<< pdiffusion >>
rect 48 229 49 230 
<< pdiffusion >>
rect 49 229 50 230 
<< pdiffusion >>
rect 50 229 51 230 
<< pdiffusion >>
rect 51 229 52 230 
<< pdiffusion >>
rect 52 229 53 230 
<< pdiffusion >>
rect 53 229 54 230 
<< m1 >>
rect 64 229 65 230 
<< pdiffusion >>
rect 66 229 67 230 
<< pdiffusion >>
rect 67 229 68 230 
<< pdiffusion >>
rect 68 229 69 230 
<< pdiffusion >>
rect 69 229 70 230 
<< pdiffusion >>
rect 70 229 71 230 
<< pdiffusion >>
rect 71 229 72 230 
<< pdiffusion >>
rect 84 229 85 230 
<< pdiffusion >>
rect 85 229 86 230 
<< pdiffusion >>
rect 86 229 87 230 
<< pdiffusion >>
rect 87 229 88 230 
<< pdiffusion >>
rect 88 229 89 230 
<< pdiffusion >>
rect 89 229 90 230 
<< pdiffusion >>
rect 102 229 103 230 
<< pdiffusion >>
rect 103 229 104 230 
<< pdiffusion >>
rect 104 229 105 230 
<< pdiffusion >>
rect 105 229 106 230 
<< pdiffusion >>
rect 106 229 107 230 
<< pdiffusion >>
rect 107 229 108 230 
<< m1 >>
rect 118 229 119 230 
<< pdiffusion >>
rect 120 229 121 230 
<< pdiffusion >>
rect 121 229 122 230 
<< pdiffusion >>
rect 122 229 123 230 
<< pdiffusion >>
rect 123 229 124 230 
<< pdiffusion >>
rect 124 229 125 230 
<< pdiffusion >>
rect 125 229 126 230 
<< m1 >>
rect 127 229 128 230 
<< pdiffusion >>
rect 138 229 139 230 
<< pdiffusion >>
rect 139 229 140 230 
<< pdiffusion >>
rect 140 229 141 230 
<< pdiffusion >>
rect 141 229 142 230 
<< pdiffusion >>
rect 142 229 143 230 
<< pdiffusion >>
rect 143 229 144 230 
<< m1 >>
rect 154 229 155 230 
<< pdiffusion >>
rect 156 229 157 230 
<< pdiffusion >>
rect 157 229 158 230 
<< pdiffusion >>
rect 158 229 159 230 
<< pdiffusion >>
rect 159 229 160 230 
<< pdiffusion >>
rect 160 229 161 230 
<< pdiffusion >>
rect 161 229 162 230 
<< m1 >>
rect 163 229 164 230 
<< m2 >>
rect 164 229 165 230 
<< pdiffusion >>
rect 174 229 175 230 
<< pdiffusion >>
rect 175 229 176 230 
<< pdiffusion >>
rect 176 229 177 230 
<< pdiffusion >>
rect 177 229 178 230 
<< pdiffusion >>
rect 178 229 179 230 
<< pdiffusion >>
rect 179 229 180 230 
<< m1 >>
rect 190 229 191 230 
<< pdiffusion >>
rect 192 229 193 230 
<< pdiffusion >>
rect 193 229 194 230 
<< pdiffusion >>
rect 194 229 195 230 
<< pdiffusion >>
rect 195 229 196 230 
<< pdiffusion >>
rect 196 229 197 230 
<< pdiffusion >>
rect 197 229 198 230 
<< m1 >>
rect 203 229 204 230 
<< m2 >>
rect 207 229 208 230 
<< m1 >>
rect 208 229 209 230 
<< pdiffusion >>
rect 210 229 211 230 
<< pdiffusion >>
rect 211 229 212 230 
<< pdiffusion >>
rect 212 229 213 230 
<< pdiffusion >>
rect 213 229 214 230 
<< pdiffusion >>
rect 214 229 215 230 
<< pdiffusion >>
rect 215 229 216 230 
<< pdiffusion >>
rect 228 229 229 230 
<< pdiffusion >>
rect 229 229 230 230 
<< pdiffusion >>
rect 230 229 231 230 
<< pdiffusion >>
rect 231 229 232 230 
<< pdiffusion >>
rect 232 229 233 230 
<< pdiffusion >>
rect 233 229 234 230 
<< m1 >>
rect 235 229 236 230 
<< m1 >>
rect 237 229 238 230 
<< m2 >>
rect 243 229 244 230 
<< m1 >>
rect 244 229 245 230 
<< pdiffusion >>
rect 246 229 247 230 
<< pdiffusion >>
rect 247 229 248 230 
<< pdiffusion >>
rect 248 229 249 230 
<< pdiffusion >>
rect 249 229 250 230 
<< pdiffusion >>
rect 250 229 251 230 
<< pdiffusion >>
rect 251 229 252 230 
<< pdiffusion >>
rect 264 229 265 230 
<< pdiffusion >>
rect 265 229 266 230 
<< pdiffusion >>
rect 266 229 267 230 
<< pdiffusion >>
rect 267 229 268 230 
<< pdiffusion >>
rect 268 229 269 230 
<< pdiffusion >>
rect 269 229 270 230 
<< pdiffusion >>
rect 282 229 283 230 
<< pdiffusion >>
rect 283 229 284 230 
<< pdiffusion >>
rect 284 229 285 230 
<< pdiffusion >>
rect 285 229 286 230 
<< pdiffusion >>
rect 286 229 287 230 
<< pdiffusion >>
rect 287 229 288 230 
<< pdiffusion >>
rect 300 229 301 230 
<< pdiffusion >>
rect 301 229 302 230 
<< pdiffusion >>
rect 302 229 303 230 
<< pdiffusion >>
rect 303 229 304 230 
<< pdiffusion >>
rect 304 229 305 230 
<< pdiffusion >>
rect 305 229 306 230 
<< m1 >>
rect 307 229 308 230 
<< m1 >>
rect 311 229 312 230 
<< pdiffusion >>
rect 318 229 319 230 
<< pdiffusion >>
rect 319 229 320 230 
<< pdiffusion >>
rect 320 229 321 230 
<< pdiffusion >>
rect 321 229 322 230 
<< pdiffusion >>
rect 322 229 323 230 
<< pdiffusion >>
rect 323 229 324 230 
<< pdiffusion >>
rect 336 229 337 230 
<< pdiffusion >>
rect 337 229 338 230 
<< pdiffusion >>
rect 338 229 339 230 
<< pdiffusion >>
rect 339 229 340 230 
<< pdiffusion >>
rect 340 229 341 230 
<< pdiffusion >>
rect 341 229 342 230 
<< m1 >>
rect 352 229 353 230 
<< pdiffusion >>
rect 354 229 355 230 
<< pdiffusion >>
rect 355 229 356 230 
<< pdiffusion >>
rect 356 229 357 230 
<< pdiffusion >>
rect 357 229 358 230 
<< pdiffusion >>
rect 358 229 359 230 
<< pdiffusion >>
rect 359 229 360 230 
<< pdiffusion >>
rect 372 229 373 230 
<< pdiffusion >>
rect 373 229 374 230 
<< pdiffusion >>
rect 374 229 375 230 
<< pdiffusion >>
rect 375 229 376 230 
<< pdiffusion >>
rect 376 229 377 230 
<< pdiffusion >>
rect 377 229 378 230 
<< pdiffusion >>
rect 390 229 391 230 
<< pdiffusion >>
rect 391 229 392 230 
<< pdiffusion >>
rect 392 229 393 230 
<< pdiffusion >>
rect 393 229 394 230 
<< pdiffusion >>
rect 394 229 395 230 
<< pdiffusion >>
rect 395 229 396 230 
<< pdiffusion >>
rect 408 229 409 230 
<< pdiffusion >>
rect 409 229 410 230 
<< pdiffusion >>
rect 410 229 411 230 
<< pdiffusion >>
rect 411 229 412 230 
<< pdiffusion >>
rect 412 229 413 230 
<< pdiffusion >>
rect 413 229 414 230 
<< pdiffusion >>
rect 426 229 427 230 
<< pdiffusion >>
rect 427 229 428 230 
<< pdiffusion >>
rect 428 229 429 230 
<< pdiffusion >>
rect 429 229 430 230 
<< pdiffusion >>
rect 430 229 431 230 
<< pdiffusion >>
rect 431 229 432 230 
<< pdiffusion >>
rect 444 229 445 230 
<< pdiffusion >>
rect 445 229 446 230 
<< pdiffusion >>
rect 446 229 447 230 
<< pdiffusion >>
rect 447 229 448 230 
<< pdiffusion >>
rect 448 229 449 230 
<< pdiffusion >>
rect 449 229 450 230 
<< pdiffusion >>
rect 12 230 13 231 
<< pdiffusion >>
rect 13 230 14 231 
<< pdiffusion >>
rect 14 230 15 231 
<< pdiffusion >>
rect 15 230 16 231 
<< pdiffusion >>
rect 16 230 17 231 
<< pdiffusion >>
rect 17 230 18 231 
<< pdiffusion >>
rect 30 230 31 231 
<< pdiffusion >>
rect 31 230 32 231 
<< pdiffusion >>
rect 32 230 33 231 
<< pdiffusion >>
rect 33 230 34 231 
<< pdiffusion >>
rect 34 230 35 231 
<< pdiffusion >>
rect 35 230 36 231 
<< pdiffusion >>
rect 48 230 49 231 
<< pdiffusion >>
rect 49 230 50 231 
<< pdiffusion >>
rect 50 230 51 231 
<< pdiffusion >>
rect 51 230 52 231 
<< pdiffusion >>
rect 52 230 53 231 
<< pdiffusion >>
rect 53 230 54 231 
<< m1 >>
rect 64 230 65 231 
<< pdiffusion >>
rect 66 230 67 231 
<< pdiffusion >>
rect 67 230 68 231 
<< pdiffusion >>
rect 68 230 69 231 
<< pdiffusion >>
rect 69 230 70 231 
<< pdiffusion >>
rect 70 230 71 231 
<< pdiffusion >>
rect 71 230 72 231 
<< pdiffusion >>
rect 84 230 85 231 
<< pdiffusion >>
rect 85 230 86 231 
<< pdiffusion >>
rect 86 230 87 231 
<< pdiffusion >>
rect 87 230 88 231 
<< pdiffusion >>
rect 88 230 89 231 
<< pdiffusion >>
rect 89 230 90 231 
<< pdiffusion >>
rect 102 230 103 231 
<< pdiffusion >>
rect 103 230 104 231 
<< pdiffusion >>
rect 104 230 105 231 
<< pdiffusion >>
rect 105 230 106 231 
<< pdiffusion >>
rect 106 230 107 231 
<< pdiffusion >>
rect 107 230 108 231 
<< m1 >>
rect 118 230 119 231 
<< pdiffusion >>
rect 120 230 121 231 
<< pdiffusion >>
rect 121 230 122 231 
<< pdiffusion >>
rect 122 230 123 231 
<< pdiffusion >>
rect 123 230 124 231 
<< pdiffusion >>
rect 124 230 125 231 
<< pdiffusion >>
rect 125 230 126 231 
<< m1 >>
rect 127 230 128 231 
<< pdiffusion >>
rect 138 230 139 231 
<< pdiffusion >>
rect 139 230 140 231 
<< pdiffusion >>
rect 140 230 141 231 
<< pdiffusion >>
rect 141 230 142 231 
<< pdiffusion >>
rect 142 230 143 231 
<< pdiffusion >>
rect 143 230 144 231 
<< m1 >>
rect 154 230 155 231 
<< pdiffusion >>
rect 156 230 157 231 
<< pdiffusion >>
rect 157 230 158 231 
<< pdiffusion >>
rect 158 230 159 231 
<< pdiffusion >>
rect 159 230 160 231 
<< pdiffusion >>
rect 160 230 161 231 
<< pdiffusion >>
rect 161 230 162 231 
<< m1 >>
rect 163 230 164 231 
<< m2 >>
rect 164 230 165 231 
<< pdiffusion >>
rect 174 230 175 231 
<< pdiffusion >>
rect 175 230 176 231 
<< pdiffusion >>
rect 176 230 177 231 
<< pdiffusion >>
rect 177 230 178 231 
<< pdiffusion >>
rect 178 230 179 231 
<< pdiffusion >>
rect 179 230 180 231 
<< m1 >>
rect 190 230 191 231 
<< pdiffusion >>
rect 192 230 193 231 
<< pdiffusion >>
rect 193 230 194 231 
<< pdiffusion >>
rect 194 230 195 231 
<< pdiffusion >>
rect 195 230 196 231 
<< pdiffusion >>
rect 196 230 197 231 
<< pdiffusion >>
rect 197 230 198 231 
<< m1 >>
rect 203 230 204 231 
<< m2 >>
rect 207 230 208 231 
<< m1 >>
rect 208 230 209 231 
<< pdiffusion >>
rect 210 230 211 231 
<< pdiffusion >>
rect 211 230 212 231 
<< pdiffusion >>
rect 212 230 213 231 
<< pdiffusion >>
rect 213 230 214 231 
<< pdiffusion >>
rect 214 230 215 231 
<< pdiffusion >>
rect 215 230 216 231 
<< pdiffusion >>
rect 228 230 229 231 
<< pdiffusion >>
rect 229 230 230 231 
<< pdiffusion >>
rect 230 230 231 231 
<< pdiffusion >>
rect 231 230 232 231 
<< pdiffusion >>
rect 232 230 233 231 
<< pdiffusion >>
rect 233 230 234 231 
<< m1 >>
rect 235 230 236 231 
<< m1 >>
rect 237 230 238 231 
<< m2 >>
rect 243 230 244 231 
<< m1 >>
rect 244 230 245 231 
<< pdiffusion >>
rect 246 230 247 231 
<< pdiffusion >>
rect 247 230 248 231 
<< pdiffusion >>
rect 248 230 249 231 
<< pdiffusion >>
rect 249 230 250 231 
<< pdiffusion >>
rect 250 230 251 231 
<< pdiffusion >>
rect 251 230 252 231 
<< pdiffusion >>
rect 264 230 265 231 
<< pdiffusion >>
rect 265 230 266 231 
<< pdiffusion >>
rect 266 230 267 231 
<< pdiffusion >>
rect 267 230 268 231 
<< pdiffusion >>
rect 268 230 269 231 
<< pdiffusion >>
rect 269 230 270 231 
<< pdiffusion >>
rect 282 230 283 231 
<< pdiffusion >>
rect 283 230 284 231 
<< pdiffusion >>
rect 284 230 285 231 
<< pdiffusion >>
rect 285 230 286 231 
<< pdiffusion >>
rect 286 230 287 231 
<< pdiffusion >>
rect 287 230 288 231 
<< pdiffusion >>
rect 300 230 301 231 
<< pdiffusion >>
rect 301 230 302 231 
<< pdiffusion >>
rect 302 230 303 231 
<< pdiffusion >>
rect 303 230 304 231 
<< pdiffusion >>
rect 304 230 305 231 
<< pdiffusion >>
rect 305 230 306 231 
<< m1 >>
rect 307 230 308 231 
<< m1 >>
rect 311 230 312 231 
<< pdiffusion >>
rect 318 230 319 231 
<< pdiffusion >>
rect 319 230 320 231 
<< pdiffusion >>
rect 320 230 321 231 
<< pdiffusion >>
rect 321 230 322 231 
<< pdiffusion >>
rect 322 230 323 231 
<< pdiffusion >>
rect 323 230 324 231 
<< pdiffusion >>
rect 336 230 337 231 
<< pdiffusion >>
rect 337 230 338 231 
<< pdiffusion >>
rect 338 230 339 231 
<< pdiffusion >>
rect 339 230 340 231 
<< pdiffusion >>
rect 340 230 341 231 
<< pdiffusion >>
rect 341 230 342 231 
<< m1 >>
rect 352 230 353 231 
<< pdiffusion >>
rect 354 230 355 231 
<< pdiffusion >>
rect 355 230 356 231 
<< pdiffusion >>
rect 356 230 357 231 
<< pdiffusion >>
rect 357 230 358 231 
<< pdiffusion >>
rect 358 230 359 231 
<< pdiffusion >>
rect 359 230 360 231 
<< pdiffusion >>
rect 372 230 373 231 
<< pdiffusion >>
rect 373 230 374 231 
<< pdiffusion >>
rect 374 230 375 231 
<< pdiffusion >>
rect 375 230 376 231 
<< pdiffusion >>
rect 376 230 377 231 
<< pdiffusion >>
rect 377 230 378 231 
<< pdiffusion >>
rect 390 230 391 231 
<< pdiffusion >>
rect 391 230 392 231 
<< pdiffusion >>
rect 392 230 393 231 
<< pdiffusion >>
rect 393 230 394 231 
<< pdiffusion >>
rect 394 230 395 231 
<< pdiffusion >>
rect 395 230 396 231 
<< pdiffusion >>
rect 408 230 409 231 
<< pdiffusion >>
rect 409 230 410 231 
<< pdiffusion >>
rect 410 230 411 231 
<< pdiffusion >>
rect 411 230 412 231 
<< pdiffusion >>
rect 412 230 413 231 
<< pdiffusion >>
rect 413 230 414 231 
<< pdiffusion >>
rect 426 230 427 231 
<< pdiffusion >>
rect 427 230 428 231 
<< pdiffusion >>
rect 428 230 429 231 
<< pdiffusion >>
rect 429 230 430 231 
<< pdiffusion >>
rect 430 230 431 231 
<< pdiffusion >>
rect 431 230 432 231 
<< pdiffusion >>
rect 444 230 445 231 
<< pdiffusion >>
rect 445 230 446 231 
<< pdiffusion >>
rect 446 230 447 231 
<< pdiffusion >>
rect 447 230 448 231 
<< pdiffusion >>
rect 448 230 449 231 
<< pdiffusion >>
rect 449 230 450 231 
<< pdiffusion >>
rect 12 231 13 232 
<< pdiffusion >>
rect 13 231 14 232 
<< pdiffusion >>
rect 14 231 15 232 
<< pdiffusion >>
rect 15 231 16 232 
<< pdiffusion >>
rect 16 231 17 232 
<< pdiffusion >>
rect 17 231 18 232 
<< pdiffusion >>
rect 30 231 31 232 
<< pdiffusion >>
rect 31 231 32 232 
<< pdiffusion >>
rect 32 231 33 232 
<< pdiffusion >>
rect 33 231 34 232 
<< pdiffusion >>
rect 34 231 35 232 
<< pdiffusion >>
rect 35 231 36 232 
<< pdiffusion >>
rect 48 231 49 232 
<< pdiffusion >>
rect 49 231 50 232 
<< pdiffusion >>
rect 50 231 51 232 
<< pdiffusion >>
rect 51 231 52 232 
<< pdiffusion >>
rect 52 231 53 232 
<< pdiffusion >>
rect 53 231 54 232 
<< m1 >>
rect 64 231 65 232 
<< pdiffusion >>
rect 66 231 67 232 
<< pdiffusion >>
rect 67 231 68 232 
<< pdiffusion >>
rect 68 231 69 232 
<< pdiffusion >>
rect 69 231 70 232 
<< pdiffusion >>
rect 70 231 71 232 
<< pdiffusion >>
rect 71 231 72 232 
<< pdiffusion >>
rect 84 231 85 232 
<< pdiffusion >>
rect 85 231 86 232 
<< pdiffusion >>
rect 86 231 87 232 
<< pdiffusion >>
rect 87 231 88 232 
<< pdiffusion >>
rect 88 231 89 232 
<< pdiffusion >>
rect 89 231 90 232 
<< pdiffusion >>
rect 102 231 103 232 
<< pdiffusion >>
rect 103 231 104 232 
<< pdiffusion >>
rect 104 231 105 232 
<< pdiffusion >>
rect 105 231 106 232 
<< pdiffusion >>
rect 106 231 107 232 
<< pdiffusion >>
rect 107 231 108 232 
<< m1 >>
rect 118 231 119 232 
<< pdiffusion >>
rect 120 231 121 232 
<< pdiffusion >>
rect 121 231 122 232 
<< pdiffusion >>
rect 122 231 123 232 
<< pdiffusion >>
rect 123 231 124 232 
<< pdiffusion >>
rect 124 231 125 232 
<< pdiffusion >>
rect 125 231 126 232 
<< m1 >>
rect 127 231 128 232 
<< pdiffusion >>
rect 138 231 139 232 
<< pdiffusion >>
rect 139 231 140 232 
<< pdiffusion >>
rect 140 231 141 232 
<< pdiffusion >>
rect 141 231 142 232 
<< pdiffusion >>
rect 142 231 143 232 
<< pdiffusion >>
rect 143 231 144 232 
<< m1 >>
rect 154 231 155 232 
<< pdiffusion >>
rect 156 231 157 232 
<< pdiffusion >>
rect 157 231 158 232 
<< pdiffusion >>
rect 158 231 159 232 
<< pdiffusion >>
rect 159 231 160 232 
<< pdiffusion >>
rect 160 231 161 232 
<< pdiffusion >>
rect 161 231 162 232 
<< m1 >>
rect 163 231 164 232 
<< m2 >>
rect 164 231 165 232 
<< pdiffusion >>
rect 174 231 175 232 
<< pdiffusion >>
rect 175 231 176 232 
<< pdiffusion >>
rect 176 231 177 232 
<< pdiffusion >>
rect 177 231 178 232 
<< pdiffusion >>
rect 178 231 179 232 
<< pdiffusion >>
rect 179 231 180 232 
<< m1 >>
rect 190 231 191 232 
<< pdiffusion >>
rect 192 231 193 232 
<< pdiffusion >>
rect 193 231 194 232 
<< pdiffusion >>
rect 194 231 195 232 
<< pdiffusion >>
rect 195 231 196 232 
<< pdiffusion >>
rect 196 231 197 232 
<< pdiffusion >>
rect 197 231 198 232 
<< m1 >>
rect 203 231 204 232 
<< m2 >>
rect 207 231 208 232 
<< m1 >>
rect 208 231 209 232 
<< pdiffusion >>
rect 210 231 211 232 
<< pdiffusion >>
rect 211 231 212 232 
<< pdiffusion >>
rect 212 231 213 232 
<< pdiffusion >>
rect 213 231 214 232 
<< pdiffusion >>
rect 214 231 215 232 
<< pdiffusion >>
rect 215 231 216 232 
<< pdiffusion >>
rect 228 231 229 232 
<< pdiffusion >>
rect 229 231 230 232 
<< pdiffusion >>
rect 230 231 231 232 
<< pdiffusion >>
rect 231 231 232 232 
<< pdiffusion >>
rect 232 231 233 232 
<< pdiffusion >>
rect 233 231 234 232 
<< m1 >>
rect 235 231 236 232 
<< m1 >>
rect 237 231 238 232 
<< m2 >>
rect 243 231 244 232 
<< m1 >>
rect 244 231 245 232 
<< pdiffusion >>
rect 246 231 247 232 
<< pdiffusion >>
rect 247 231 248 232 
<< pdiffusion >>
rect 248 231 249 232 
<< pdiffusion >>
rect 249 231 250 232 
<< pdiffusion >>
rect 250 231 251 232 
<< pdiffusion >>
rect 251 231 252 232 
<< pdiffusion >>
rect 264 231 265 232 
<< pdiffusion >>
rect 265 231 266 232 
<< pdiffusion >>
rect 266 231 267 232 
<< pdiffusion >>
rect 267 231 268 232 
<< pdiffusion >>
rect 268 231 269 232 
<< pdiffusion >>
rect 269 231 270 232 
<< pdiffusion >>
rect 282 231 283 232 
<< pdiffusion >>
rect 283 231 284 232 
<< pdiffusion >>
rect 284 231 285 232 
<< pdiffusion >>
rect 285 231 286 232 
<< pdiffusion >>
rect 286 231 287 232 
<< pdiffusion >>
rect 287 231 288 232 
<< pdiffusion >>
rect 300 231 301 232 
<< pdiffusion >>
rect 301 231 302 232 
<< pdiffusion >>
rect 302 231 303 232 
<< pdiffusion >>
rect 303 231 304 232 
<< pdiffusion >>
rect 304 231 305 232 
<< pdiffusion >>
rect 305 231 306 232 
<< m1 >>
rect 307 231 308 232 
<< m1 >>
rect 311 231 312 232 
<< pdiffusion >>
rect 318 231 319 232 
<< pdiffusion >>
rect 319 231 320 232 
<< pdiffusion >>
rect 320 231 321 232 
<< pdiffusion >>
rect 321 231 322 232 
<< pdiffusion >>
rect 322 231 323 232 
<< pdiffusion >>
rect 323 231 324 232 
<< pdiffusion >>
rect 336 231 337 232 
<< pdiffusion >>
rect 337 231 338 232 
<< pdiffusion >>
rect 338 231 339 232 
<< pdiffusion >>
rect 339 231 340 232 
<< pdiffusion >>
rect 340 231 341 232 
<< pdiffusion >>
rect 341 231 342 232 
<< m1 >>
rect 352 231 353 232 
<< pdiffusion >>
rect 354 231 355 232 
<< pdiffusion >>
rect 355 231 356 232 
<< pdiffusion >>
rect 356 231 357 232 
<< pdiffusion >>
rect 357 231 358 232 
<< pdiffusion >>
rect 358 231 359 232 
<< pdiffusion >>
rect 359 231 360 232 
<< pdiffusion >>
rect 372 231 373 232 
<< pdiffusion >>
rect 373 231 374 232 
<< pdiffusion >>
rect 374 231 375 232 
<< pdiffusion >>
rect 375 231 376 232 
<< pdiffusion >>
rect 376 231 377 232 
<< pdiffusion >>
rect 377 231 378 232 
<< pdiffusion >>
rect 390 231 391 232 
<< pdiffusion >>
rect 391 231 392 232 
<< pdiffusion >>
rect 392 231 393 232 
<< pdiffusion >>
rect 393 231 394 232 
<< pdiffusion >>
rect 394 231 395 232 
<< pdiffusion >>
rect 395 231 396 232 
<< pdiffusion >>
rect 408 231 409 232 
<< pdiffusion >>
rect 409 231 410 232 
<< pdiffusion >>
rect 410 231 411 232 
<< pdiffusion >>
rect 411 231 412 232 
<< pdiffusion >>
rect 412 231 413 232 
<< pdiffusion >>
rect 413 231 414 232 
<< pdiffusion >>
rect 426 231 427 232 
<< pdiffusion >>
rect 427 231 428 232 
<< pdiffusion >>
rect 428 231 429 232 
<< pdiffusion >>
rect 429 231 430 232 
<< pdiffusion >>
rect 430 231 431 232 
<< pdiffusion >>
rect 431 231 432 232 
<< pdiffusion >>
rect 444 231 445 232 
<< pdiffusion >>
rect 445 231 446 232 
<< pdiffusion >>
rect 446 231 447 232 
<< pdiffusion >>
rect 447 231 448 232 
<< pdiffusion >>
rect 448 231 449 232 
<< pdiffusion >>
rect 449 231 450 232 
<< pdiffusion >>
rect 12 232 13 233 
<< pdiffusion >>
rect 13 232 14 233 
<< pdiffusion >>
rect 14 232 15 233 
<< pdiffusion >>
rect 15 232 16 233 
<< pdiffusion >>
rect 16 232 17 233 
<< pdiffusion >>
rect 17 232 18 233 
<< pdiffusion >>
rect 30 232 31 233 
<< pdiffusion >>
rect 31 232 32 233 
<< pdiffusion >>
rect 32 232 33 233 
<< pdiffusion >>
rect 33 232 34 233 
<< pdiffusion >>
rect 34 232 35 233 
<< pdiffusion >>
rect 35 232 36 233 
<< pdiffusion >>
rect 48 232 49 233 
<< pdiffusion >>
rect 49 232 50 233 
<< pdiffusion >>
rect 50 232 51 233 
<< pdiffusion >>
rect 51 232 52 233 
<< pdiffusion >>
rect 52 232 53 233 
<< pdiffusion >>
rect 53 232 54 233 
<< m1 >>
rect 64 232 65 233 
<< pdiffusion >>
rect 66 232 67 233 
<< pdiffusion >>
rect 67 232 68 233 
<< pdiffusion >>
rect 68 232 69 233 
<< pdiffusion >>
rect 69 232 70 233 
<< pdiffusion >>
rect 70 232 71 233 
<< pdiffusion >>
rect 71 232 72 233 
<< pdiffusion >>
rect 84 232 85 233 
<< pdiffusion >>
rect 85 232 86 233 
<< pdiffusion >>
rect 86 232 87 233 
<< pdiffusion >>
rect 87 232 88 233 
<< pdiffusion >>
rect 88 232 89 233 
<< pdiffusion >>
rect 89 232 90 233 
<< pdiffusion >>
rect 102 232 103 233 
<< pdiffusion >>
rect 103 232 104 233 
<< pdiffusion >>
rect 104 232 105 233 
<< pdiffusion >>
rect 105 232 106 233 
<< pdiffusion >>
rect 106 232 107 233 
<< pdiffusion >>
rect 107 232 108 233 
<< m1 >>
rect 118 232 119 233 
<< pdiffusion >>
rect 120 232 121 233 
<< pdiffusion >>
rect 121 232 122 233 
<< pdiffusion >>
rect 122 232 123 233 
<< pdiffusion >>
rect 123 232 124 233 
<< pdiffusion >>
rect 124 232 125 233 
<< pdiffusion >>
rect 125 232 126 233 
<< m1 >>
rect 127 232 128 233 
<< pdiffusion >>
rect 138 232 139 233 
<< pdiffusion >>
rect 139 232 140 233 
<< pdiffusion >>
rect 140 232 141 233 
<< pdiffusion >>
rect 141 232 142 233 
<< pdiffusion >>
rect 142 232 143 233 
<< pdiffusion >>
rect 143 232 144 233 
<< m1 >>
rect 154 232 155 233 
<< pdiffusion >>
rect 156 232 157 233 
<< pdiffusion >>
rect 157 232 158 233 
<< pdiffusion >>
rect 158 232 159 233 
<< pdiffusion >>
rect 159 232 160 233 
<< pdiffusion >>
rect 160 232 161 233 
<< pdiffusion >>
rect 161 232 162 233 
<< m1 >>
rect 163 232 164 233 
<< m2 >>
rect 164 232 165 233 
<< pdiffusion >>
rect 174 232 175 233 
<< pdiffusion >>
rect 175 232 176 233 
<< pdiffusion >>
rect 176 232 177 233 
<< pdiffusion >>
rect 177 232 178 233 
<< pdiffusion >>
rect 178 232 179 233 
<< pdiffusion >>
rect 179 232 180 233 
<< m1 >>
rect 190 232 191 233 
<< pdiffusion >>
rect 192 232 193 233 
<< pdiffusion >>
rect 193 232 194 233 
<< pdiffusion >>
rect 194 232 195 233 
<< pdiffusion >>
rect 195 232 196 233 
<< pdiffusion >>
rect 196 232 197 233 
<< pdiffusion >>
rect 197 232 198 233 
<< m1 >>
rect 203 232 204 233 
<< m2 >>
rect 207 232 208 233 
<< m1 >>
rect 208 232 209 233 
<< pdiffusion >>
rect 210 232 211 233 
<< pdiffusion >>
rect 211 232 212 233 
<< pdiffusion >>
rect 212 232 213 233 
<< pdiffusion >>
rect 213 232 214 233 
<< pdiffusion >>
rect 214 232 215 233 
<< pdiffusion >>
rect 215 232 216 233 
<< pdiffusion >>
rect 228 232 229 233 
<< pdiffusion >>
rect 229 232 230 233 
<< pdiffusion >>
rect 230 232 231 233 
<< pdiffusion >>
rect 231 232 232 233 
<< pdiffusion >>
rect 232 232 233 233 
<< pdiffusion >>
rect 233 232 234 233 
<< m1 >>
rect 235 232 236 233 
<< m1 >>
rect 237 232 238 233 
<< m2 >>
rect 243 232 244 233 
<< m1 >>
rect 244 232 245 233 
<< pdiffusion >>
rect 246 232 247 233 
<< pdiffusion >>
rect 247 232 248 233 
<< pdiffusion >>
rect 248 232 249 233 
<< pdiffusion >>
rect 249 232 250 233 
<< pdiffusion >>
rect 250 232 251 233 
<< pdiffusion >>
rect 251 232 252 233 
<< pdiffusion >>
rect 264 232 265 233 
<< pdiffusion >>
rect 265 232 266 233 
<< pdiffusion >>
rect 266 232 267 233 
<< pdiffusion >>
rect 267 232 268 233 
<< pdiffusion >>
rect 268 232 269 233 
<< pdiffusion >>
rect 269 232 270 233 
<< pdiffusion >>
rect 282 232 283 233 
<< pdiffusion >>
rect 283 232 284 233 
<< pdiffusion >>
rect 284 232 285 233 
<< pdiffusion >>
rect 285 232 286 233 
<< pdiffusion >>
rect 286 232 287 233 
<< pdiffusion >>
rect 287 232 288 233 
<< pdiffusion >>
rect 300 232 301 233 
<< pdiffusion >>
rect 301 232 302 233 
<< pdiffusion >>
rect 302 232 303 233 
<< pdiffusion >>
rect 303 232 304 233 
<< pdiffusion >>
rect 304 232 305 233 
<< pdiffusion >>
rect 305 232 306 233 
<< m1 >>
rect 307 232 308 233 
<< m1 >>
rect 311 232 312 233 
<< pdiffusion >>
rect 318 232 319 233 
<< pdiffusion >>
rect 319 232 320 233 
<< pdiffusion >>
rect 320 232 321 233 
<< pdiffusion >>
rect 321 232 322 233 
<< pdiffusion >>
rect 322 232 323 233 
<< pdiffusion >>
rect 323 232 324 233 
<< pdiffusion >>
rect 336 232 337 233 
<< pdiffusion >>
rect 337 232 338 233 
<< pdiffusion >>
rect 338 232 339 233 
<< pdiffusion >>
rect 339 232 340 233 
<< pdiffusion >>
rect 340 232 341 233 
<< pdiffusion >>
rect 341 232 342 233 
<< m1 >>
rect 352 232 353 233 
<< pdiffusion >>
rect 354 232 355 233 
<< pdiffusion >>
rect 355 232 356 233 
<< pdiffusion >>
rect 356 232 357 233 
<< pdiffusion >>
rect 357 232 358 233 
<< pdiffusion >>
rect 358 232 359 233 
<< pdiffusion >>
rect 359 232 360 233 
<< pdiffusion >>
rect 372 232 373 233 
<< pdiffusion >>
rect 373 232 374 233 
<< pdiffusion >>
rect 374 232 375 233 
<< pdiffusion >>
rect 375 232 376 233 
<< pdiffusion >>
rect 376 232 377 233 
<< pdiffusion >>
rect 377 232 378 233 
<< pdiffusion >>
rect 390 232 391 233 
<< pdiffusion >>
rect 391 232 392 233 
<< pdiffusion >>
rect 392 232 393 233 
<< pdiffusion >>
rect 393 232 394 233 
<< pdiffusion >>
rect 394 232 395 233 
<< pdiffusion >>
rect 395 232 396 233 
<< pdiffusion >>
rect 408 232 409 233 
<< pdiffusion >>
rect 409 232 410 233 
<< pdiffusion >>
rect 410 232 411 233 
<< pdiffusion >>
rect 411 232 412 233 
<< pdiffusion >>
rect 412 232 413 233 
<< pdiffusion >>
rect 413 232 414 233 
<< pdiffusion >>
rect 426 232 427 233 
<< pdiffusion >>
rect 427 232 428 233 
<< pdiffusion >>
rect 428 232 429 233 
<< pdiffusion >>
rect 429 232 430 233 
<< pdiffusion >>
rect 430 232 431 233 
<< pdiffusion >>
rect 431 232 432 233 
<< pdiffusion >>
rect 444 232 445 233 
<< pdiffusion >>
rect 445 232 446 233 
<< pdiffusion >>
rect 446 232 447 233 
<< pdiffusion >>
rect 447 232 448 233 
<< pdiffusion >>
rect 448 232 449 233 
<< pdiffusion >>
rect 449 232 450 233 
<< pdiffusion >>
rect 12 233 13 234 
<< pdiffusion >>
rect 13 233 14 234 
<< pdiffusion >>
rect 14 233 15 234 
<< pdiffusion >>
rect 15 233 16 234 
<< pdiffusion >>
rect 16 233 17 234 
<< pdiffusion >>
rect 17 233 18 234 
<< pdiffusion >>
rect 30 233 31 234 
<< pdiffusion >>
rect 31 233 32 234 
<< pdiffusion >>
rect 32 233 33 234 
<< pdiffusion >>
rect 33 233 34 234 
<< pdiffusion >>
rect 34 233 35 234 
<< pdiffusion >>
rect 35 233 36 234 
<< pdiffusion >>
rect 48 233 49 234 
<< pdiffusion >>
rect 49 233 50 234 
<< pdiffusion >>
rect 50 233 51 234 
<< pdiffusion >>
rect 51 233 52 234 
<< pdiffusion >>
rect 52 233 53 234 
<< pdiffusion >>
rect 53 233 54 234 
<< m1 >>
rect 64 233 65 234 
<< pdiffusion >>
rect 66 233 67 234 
<< pdiffusion >>
rect 67 233 68 234 
<< pdiffusion >>
rect 68 233 69 234 
<< pdiffusion >>
rect 69 233 70 234 
<< pdiffusion >>
rect 70 233 71 234 
<< pdiffusion >>
rect 71 233 72 234 
<< pdiffusion >>
rect 84 233 85 234 
<< m1 >>
rect 85 233 86 234 
<< pdiffusion >>
rect 85 233 86 234 
<< pdiffusion >>
rect 86 233 87 234 
<< pdiffusion >>
rect 87 233 88 234 
<< pdiffusion >>
rect 88 233 89 234 
<< pdiffusion >>
rect 89 233 90 234 
<< pdiffusion >>
rect 102 233 103 234 
<< pdiffusion >>
rect 103 233 104 234 
<< pdiffusion >>
rect 104 233 105 234 
<< pdiffusion >>
rect 105 233 106 234 
<< pdiffusion >>
rect 106 233 107 234 
<< pdiffusion >>
rect 107 233 108 234 
<< m1 >>
rect 118 233 119 234 
<< pdiffusion >>
rect 120 233 121 234 
<< pdiffusion >>
rect 121 233 122 234 
<< pdiffusion >>
rect 122 233 123 234 
<< pdiffusion >>
rect 123 233 124 234 
<< pdiffusion >>
rect 124 233 125 234 
<< pdiffusion >>
rect 125 233 126 234 
<< m1 >>
rect 127 233 128 234 
<< pdiffusion >>
rect 138 233 139 234 
<< pdiffusion >>
rect 139 233 140 234 
<< pdiffusion >>
rect 140 233 141 234 
<< pdiffusion >>
rect 141 233 142 234 
<< pdiffusion >>
rect 142 233 143 234 
<< pdiffusion >>
rect 143 233 144 234 
<< m1 >>
rect 154 233 155 234 
<< pdiffusion >>
rect 156 233 157 234 
<< m1 >>
rect 157 233 158 234 
<< pdiffusion >>
rect 157 233 158 234 
<< pdiffusion >>
rect 158 233 159 234 
<< pdiffusion >>
rect 159 233 160 234 
<< pdiffusion >>
rect 160 233 161 234 
<< pdiffusion >>
rect 161 233 162 234 
<< m1 >>
rect 163 233 164 234 
<< m2 >>
rect 164 233 165 234 
<< pdiffusion >>
rect 174 233 175 234 
<< pdiffusion >>
rect 175 233 176 234 
<< pdiffusion >>
rect 176 233 177 234 
<< pdiffusion >>
rect 177 233 178 234 
<< pdiffusion >>
rect 178 233 179 234 
<< pdiffusion >>
rect 179 233 180 234 
<< m1 >>
rect 190 233 191 234 
<< pdiffusion >>
rect 192 233 193 234 
<< pdiffusion >>
rect 193 233 194 234 
<< pdiffusion >>
rect 194 233 195 234 
<< pdiffusion >>
rect 195 233 196 234 
<< pdiffusion >>
rect 196 233 197 234 
<< pdiffusion >>
rect 197 233 198 234 
<< m1 >>
rect 203 233 204 234 
<< m2 >>
rect 207 233 208 234 
<< m1 >>
rect 208 233 209 234 
<< pdiffusion >>
rect 210 233 211 234 
<< pdiffusion >>
rect 211 233 212 234 
<< pdiffusion >>
rect 212 233 213 234 
<< pdiffusion >>
rect 213 233 214 234 
<< m1 >>
rect 214 233 215 234 
<< pdiffusion >>
rect 214 233 215 234 
<< pdiffusion >>
rect 215 233 216 234 
<< pdiffusion >>
rect 228 233 229 234 
<< pdiffusion >>
rect 229 233 230 234 
<< pdiffusion >>
rect 230 233 231 234 
<< pdiffusion >>
rect 231 233 232 234 
<< m1 >>
rect 232 233 233 234 
<< pdiffusion >>
rect 232 233 233 234 
<< pdiffusion >>
rect 233 233 234 234 
<< m1 >>
rect 235 233 236 234 
<< m1 >>
rect 237 233 238 234 
<< m2 >>
rect 243 233 244 234 
<< m1 >>
rect 244 233 245 234 
<< pdiffusion >>
rect 246 233 247 234 
<< m1 >>
rect 247 233 248 234 
<< pdiffusion >>
rect 247 233 248 234 
<< pdiffusion >>
rect 248 233 249 234 
<< pdiffusion >>
rect 249 233 250 234 
<< pdiffusion >>
rect 250 233 251 234 
<< pdiffusion >>
rect 251 233 252 234 
<< pdiffusion >>
rect 264 233 265 234 
<< pdiffusion >>
rect 265 233 266 234 
<< pdiffusion >>
rect 266 233 267 234 
<< pdiffusion >>
rect 267 233 268 234 
<< pdiffusion >>
rect 268 233 269 234 
<< pdiffusion >>
rect 269 233 270 234 
<< pdiffusion >>
rect 282 233 283 234 
<< pdiffusion >>
rect 283 233 284 234 
<< pdiffusion >>
rect 284 233 285 234 
<< pdiffusion >>
rect 285 233 286 234 
<< pdiffusion >>
rect 286 233 287 234 
<< pdiffusion >>
rect 287 233 288 234 
<< pdiffusion >>
rect 300 233 301 234 
<< pdiffusion >>
rect 301 233 302 234 
<< pdiffusion >>
rect 302 233 303 234 
<< pdiffusion >>
rect 303 233 304 234 
<< pdiffusion >>
rect 304 233 305 234 
<< pdiffusion >>
rect 305 233 306 234 
<< m1 >>
rect 307 233 308 234 
<< m1 >>
rect 311 233 312 234 
<< pdiffusion >>
rect 318 233 319 234 
<< pdiffusion >>
rect 319 233 320 234 
<< pdiffusion >>
rect 320 233 321 234 
<< pdiffusion >>
rect 321 233 322 234 
<< m1 >>
rect 322 233 323 234 
<< pdiffusion >>
rect 322 233 323 234 
<< pdiffusion >>
rect 323 233 324 234 
<< pdiffusion >>
rect 336 233 337 234 
<< pdiffusion >>
rect 337 233 338 234 
<< pdiffusion >>
rect 338 233 339 234 
<< pdiffusion >>
rect 339 233 340 234 
<< pdiffusion >>
rect 340 233 341 234 
<< pdiffusion >>
rect 341 233 342 234 
<< m1 >>
rect 352 233 353 234 
<< pdiffusion >>
rect 354 233 355 234 
<< pdiffusion >>
rect 355 233 356 234 
<< pdiffusion >>
rect 356 233 357 234 
<< pdiffusion >>
rect 357 233 358 234 
<< pdiffusion >>
rect 358 233 359 234 
<< pdiffusion >>
rect 359 233 360 234 
<< pdiffusion >>
rect 372 233 373 234 
<< pdiffusion >>
rect 373 233 374 234 
<< pdiffusion >>
rect 374 233 375 234 
<< pdiffusion >>
rect 375 233 376 234 
<< pdiffusion >>
rect 376 233 377 234 
<< pdiffusion >>
rect 377 233 378 234 
<< pdiffusion >>
rect 390 233 391 234 
<< m1 >>
rect 391 233 392 234 
<< pdiffusion >>
rect 391 233 392 234 
<< pdiffusion >>
rect 392 233 393 234 
<< pdiffusion >>
rect 393 233 394 234 
<< pdiffusion >>
rect 394 233 395 234 
<< pdiffusion >>
rect 395 233 396 234 
<< pdiffusion >>
rect 408 233 409 234 
<< pdiffusion >>
rect 409 233 410 234 
<< pdiffusion >>
rect 410 233 411 234 
<< pdiffusion >>
rect 411 233 412 234 
<< pdiffusion >>
rect 412 233 413 234 
<< pdiffusion >>
rect 413 233 414 234 
<< pdiffusion >>
rect 426 233 427 234 
<< pdiffusion >>
rect 427 233 428 234 
<< pdiffusion >>
rect 428 233 429 234 
<< pdiffusion >>
rect 429 233 430 234 
<< pdiffusion >>
rect 430 233 431 234 
<< pdiffusion >>
rect 431 233 432 234 
<< pdiffusion >>
rect 444 233 445 234 
<< pdiffusion >>
rect 445 233 446 234 
<< pdiffusion >>
rect 446 233 447 234 
<< pdiffusion >>
rect 447 233 448 234 
<< pdiffusion >>
rect 448 233 449 234 
<< pdiffusion >>
rect 449 233 450 234 
<< m1 >>
rect 64 234 65 235 
<< m1 >>
rect 85 234 86 235 
<< m1 >>
rect 118 234 119 235 
<< m1 >>
rect 127 234 128 235 
<< m1 >>
rect 154 234 155 235 
<< m1 >>
rect 157 234 158 235 
<< m1 >>
rect 163 234 164 235 
<< m2 >>
rect 164 234 165 235 
<< m1 >>
rect 190 234 191 235 
<< m1 >>
rect 203 234 204 235 
<< m2 >>
rect 207 234 208 235 
<< m1 >>
rect 208 234 209 235 
<< m1 >>
rect 214 234 215 235 
<< m1 >>
rect 232 234 233 235 
<< m1 >>
rect 235 234 236 235 
<< m1 >>
rect 237 234 238 235 
<< m2 >>
rect 243 234 244 235 
<< m1 >>
rect 244 234 245 235 
<< m1 >>
rect 247 234 248 235 
<< m1 >>
rect 307 234 308 235 
<< m1 >>
rect 311 234 312 235 
<< m1 >>
rect 322 234 323 235 
<< m1 >>
rect 352 234 353 235 
<< m1 >>
rect 391 234 392 235 
<< m1 >>
rect 64 235 65 236 
<< m1 >>
rect 85 235 86 236 
<< m1 >>
rect 118 235 119 236 
<< m1 >>
rect 127 235 128 236 
<< m1 >>
rect 154 235 155 236 
<< m1 >>
rect 155 235 156 236 
<< m1 >>
rect 156 235 157 236 
<< m1 >>
rect 157 235 158 236 
<< m1 >>
rect 161 235 162 236 
<< m2 >>
rect 161 235 162 236 
<< m2c >>
rect 161 235 162 236 
<< m1 >>
rect 161 235 162 236 
<< m2 >>
rect 161 235 162 236 
<< m2 >>
rect 162 235 163 236 
<< m1 >>
rect 163 235 164 236 
<< m2 >>
rect 163 235 164 236 
<< m2 >>
rect 164 235 165 236 
<< m1 >>
rect 190 235 191 236 
<< m1 >>
rect 203 235 204 236 
<< m2 >>
rect 207 235 208 236 
<< m1 >>
rect 208 235 209 236 
<< m2 >>
rect 208 235 209 236 
<< m2 >>
rect 209 235 210 236 
<< m1 >>
rect 210 235 211 236 
<< m2 >>
rect 210 235 211 236 
<< m2c >>
rect 210 235 211 236 
<< m1 >>
rect 210 235 211 236 
<< m2 >>
rect 210 235 211 236 
<< m1 >>
rect 214 235 215 236 
<< m1 >>
rect 232 235 233 236 
<< m1 >>
rect 233 235 234 236 
<< m1 >>
rect 234 235 235 236 
<< m1 >>
rect 235 235 236 236 
<< m1 >>
rect 237 235 238 236 
<< m2 >>
rect 243 235 244 236 
<< m1 >>
rect 244 235 245 236 
<< m2 >>
rect 244 235 245 236 
<< m2 >>
rect 245 235 246 236 
<< m1 >>
rect 246 235 247 236 
<< m2 >>
rect 246 235 247 236 
<< m2c >>
rect 246 235 247 236 
<< m1 >>
rect 246 235 247 236 
<< m2 >>
rect 246 235 247 236 
<< m1 >>
rect 247 235 248 236 
<< m1 >>
rect 307 235 308 236 
<< m1 >>
rect 311 235 312 236 
<< m1 >>
rect 322 235 323 236 
<< m1 >>
rect 352 235 353 236 
<< m1 >>
rect 391 235 392 236 
<< m1 >>
rect 64 236 65 237 
<< m1 >>
rect 85 236 86 237 
<< m1 >>
rect 118 236 119 237 
<< m1 >>
rect 127 236 128 237 
<< m1 >>
rect 161 236 162 237 
<< m1 >>
rect 163 236 164 237 
<< m1 >>
rect 190 236 191 237 
<< m1 >>
rect 203 236 204 237 
<< m1 >>
rect 208 236 209 237 
<< m1 >>
rect 210 236 211 237 
<< m1 >>
rect 214 236 215 237 
<< m1 >>
rect 237 236 238 237 
<< m1 >>
rect 244 236 245 237 
<< m1 >>
rect 307 236 308 237 
<< m1 >>
rect 311 236 312 237 
<< m1 >>
rect 322 236 323 237 
<< m1 >>
rect 352 236 353 237 
<< m1 >>
rect 391 236 392 237 
<< m1 >>
rect 64 237 65 238 
<< m1 >>
rect 85 237 86 238 
<< m1 >>
rect 118 237 119 238 
<< m1 >>
rect 127 237 128 238 
<< m1 >>
rect 161 237 162 238 
<< m1 >>
rect 163 237 164 238 
<< m1 >>
rect 190 237 191 238 
<< m1 >>
rect 203 237 204 238 
<< m1 >>
rect 208 237 209 238 
<< m1 >>
rect 210 237 211 238 
<< m1 >>
rect 214 237 215 238 
<< m1 >>
rect 237 237 238 238 
<< m1 >>
rect 238 237 239 238 
<< m1 >>
rect 239 237 240 238 
<< m1 >>
rect 240 237 241 238 
<< m1 >>
rect 241 237 242 238 
<< m1 >>
rect 242 237 243 238 
<< m2 >>
rect 242 237 243 238 
<< m2c >>
rect 242 237 243 238 
<< m1 >>
rect 242 237 243 238 
<< m2 >>
rect 242 237 243 238 
<< m2 >>
rect 243 237 244 238 
<< m1 >>
rect 244 237 245 238 
<< m1 >>
rect 307 237 308 238 
<< m1 >>
rect 311 237 312 238 
<< m1 >>
rect 322 237 323 238 
<< m1 >>
rect 352 237 353 238 
<< m1 >>
rect 391 237 392 238 
<< m1 >>
rect 64 238 65 239 
<< m1 >>
rect 85 238 86 239 
<< m1 >>
rect 86 238 87 239 
<< m1 >>
rect 87 238 88 239 
<< m1 >>
rect 88 238 89 239 
<< m1 >>
rect 89 238 90 239 
<< m1 >>
rect 90 238 91 239 
<< m1 >>
rect 91 238 92 239 
<< m1 >>
rect 92 238 93 239 
<< m1 >>
rect 93 238 94 239 
<< m1 >>
rect 94 238 95 239 
<< m1 >>
rect 95 238 96 239 
<< m1 >>
rect 96 238 97 239 
<< m1 >>
rect 97 238 98 239 
<< m1 >>
rect 98 238 99 239 
<< m1 >>
rect 99 238 100 239 
<< m1 >>
rect 100 238 101 239 
<< m1 >>
rect 101 238 102 239 
<< m1 >>
rect 102 238 103 239 
<< m1 >>
rect 103 238 104 239 
<< m1 >>
rect 104 238 105 239 
<< m1 >>
rect 105 238 106 239 
<< m1 >>
rect 106 238 107 239 
<< m1 >>
rect 118 238 119 239 
<< m1 >>
rect 127 238 128 239 
<< m1 >>
rect 138 238 139 239 
<< m1 >>
rect 139 238 140 239 
<< m1 >>
rect 140 238 141 239 
<< m1 >>
rect 141 238 142 239 
<< m1 >>
rect 142 238 143 239 
<< m1 >>
rect 143 238 144 239 
<< m1 >>
rect 144 238 145 239 
<< m1 >>
rect 145 238 146 239 
<< m1 >>
rect 146 238 147 239 
<< m1 >>
rect 147 238 148 239 
<< m1 >>
rect 148 238 149 239 
<< m1 >>
rect 149 238 150 239 
<< m1 >>
rect 150 238 151 239 
<< m1 >>
rect 151 238 152 239 
<< m1 >>
rect 152 238 153 239 
<< m1 >>
rect 153 238 154 239 
<< m1 >>
rect 154 238 155 239 
<< m1 >>
rect 155 238 156 239 
<< m1 >>
rect 156 238 157 239 
<< m1 >>
rect 157 238 158 239 
<< m1 >>
rect 158 238 159 239 
<< m1 >>
rect 159 238 160 239 
<< m1 >>
rect 160 238 161 239 
<< m1 >>
rect 161 238 162 239 
<< m1 >>
rect 163 238 164 239 
<< m1 >>
rect 190 238 191 239 
<< m1 >>
rect 203 238 204 239 
<< m1 >>
rect 208 238 209 239 
<< m1 >>
rect 210 238 211 239 
<< m1 >>
rect 211 238 212 239 
<< m1 >>
rect 212 238 213 239 
<< m1 >>
rect 213 238 214 239 
<< m1 >>
rect 214 238 215 239 
<< m2 >>
rect 243 238 244 239 
<< m1 >>
rect 244 238 245 239 
<< m1 >>
rect 247 238 248 239 
<< m1 >>
rect 248 238 249 239 
<< m1 >>
rect 249 238 250 239 
<< m1 >>
rect 250 238 251 239 
<< m1 >>
rect 251 238 252 239 
<< m1 >>
rect 252 238 253 239 
<< m1 >>
rect 253 238 254 239 
<< m1 >>
rect 254 238 255 239 
<< m1 >>
rect 255 238 256 239 
<< m1 >>
rect 256 238 257 239 
<< m1 >>
rect 257 238 258 239 
<< m1 >>
rect 258 238 259 239 
<< m1 >>
rect 259 238 260 239 
<< m1 >>
rect 260 238 261 239 
<< m1 >>
rect 261 238 262 239 
<< m1 >>
rect 262 238 263 239 
<< m1 >>
rect 263 238 264 239 
<< m1 >>
rect 264 238 265 239 
<< m1 >>
rect 265 238 266 239 
<< m1 >>
rect 266 238 267 239 
<< m1 >>
rect 267 238 268 239 
<< m1 >>
rect 268 238 269 239 
<< m1 >>
rect 269 238 270 239 
<< m1 >>
rect 270 238 271 239 
<< m1 >>
rect 271 238 272 239 
<< m1 >>
rect 272 238 273 239 
<< m1 >>
rect 273 238 274 239 
<< m1 >>
rect 274 238 275 239 
<< m1 >>
rect 275 238 276 239 
<< m1 >>
rect 276 238 277 239 
<< m1 >>
rect 277 238 278 239 
<< m1 >>
rect 278 238 279 239 
<< m1 >>
rect 279 238 280 239 
<< m1 >>
rect 280 238 281 239 
<< m1 >>
rect 281 238 282 239 
<< m1 >>
rect 282 238 283 239 
<< m1 >>
rect 283 238 284 239 
<< m1 >>
rect 284 238 285 239 
<< m1 >>
rect 285 238 286 239 
<< m1 >>
rect 286 238 287 239 
<< m1 >>
rect 287 238 288 239 
<< m1 >>
rect 288 238 289 239 
<< m1 >>
rect 289 238 290 239 
<< m1 >>
rect 290 238 291 239 
<< m1 >>
rect 291 238 292 239 
<< m1 >>
rect 292 238 293 239 
<< m1 >>
rect 293 238 294 239 
<< m1 >>
rect 294 238 295 239 
<< m1 >>
rect 295 238 296 239 
<< m1 >>
rect 296 238 297 239 
<< m1 >>
rect 297 238 298 239 
<< m1 >>
rect 298 238 299 239 
<< m1 >>
rect 299 238 300 239 
<< m1 >>
rect 300 238 301 239 
<< m1 >>
rect 301 238 302 239 
<< m1 >>
rect 302 238 303 239 
<< m1 >>
rect 303 238 304 239 
<< m1 >>
rect 304 238 305 239 
<< m1 >>
rect 305 238 306 239 
<< m1 >>
rect 306 238 307 239 
<< m1 >>
rect 307 238 308 239 
<< m1 >>
rect 311 238 312 239 
<< m1 >>
rect 322 238 323 239 
<< m1 >>
rect 352 238 353 239 
<< m1 >>
rect 391 238 392 239 
<< m1 >>
rect 64 239 65 240 
<< m1 >>
rect 106 239 107 240 
<< m1 >>
rect 118 239 119 240 
<< m1 >>
rect 127 239 128 240 
<< m1 >>
rect 138 239 139 240 
<< m1 >>
rect 163 239 164 240 
<< m1 >>
rect 190 239 191 240 
<< m1 >>
rect 203 239 204 240 
<< m1 >>
rect 208 239 209 240 
<< m2 >>
rect 243 239 244 240 
<< m1 >>
rect 244 239 245 240 
<< m1 >>
rect 247 239 248 240 
<< m2 >>
rect 304 239 305 240 
<< m2 >>
rect 305 239 306 240 
<< m2 >>
rect 306 239 307 240 
<< m2 >>
rect 307 239 308 240 
<< m2 >>
rect 308 239 309 240 
<< m1 >>
rect 309 239 310 240 
<< m2 >>
rect 309 239 310 240 
<< m2c >>
rect 309 239 310 240 
<< m1 >>
rect 309 239 310 240 
<< m2 >>
rect 309 239 310 240 
<< m1 >>
rect 310 239 311 240 
<< m1 >>
rect 311 239 312 240 
<< m1 >>
rect 322 239 323 240 
<< m1 >>
rect 352 239 353 240 
<< m1 >>
rect 391 239 392 240 
<< m1 >>
rect 64 240 65 241 
<< m1 >>
rect 106 240 107 241 
<< m1 >>
rect 118 240 119 241 
<< m1 >>
rect 127 240 128 241 
<< m1 >>
rect 138 240 139 241 
<< m1 >>
rect 163 240 164 241 
<< m1 >>
rect 190 240 191 241 
<< m1 >>
rect 203 240 204 241 
<< m1 >>
rect 208 240 209 241 
<< m2 >>
rect 243 240 244 241 
<< m1 >>
rect 244 240 245 241 
<< m2 >>
rect 244 240 245 241 
<< m2 >>
rect 245 240 246 241 
<< m2 >>
rect 246 240 247 241 
<< m1 >>
rect 247 240 248 241 
<< m2 >>
rect 247 240 248 241 
<< m2 >>
rect 248 240 249 241 
<< m1 >>
rect 249 240 250 241 
<< m2 >>
rect 249 240 250 241 
<< m2c >>
rect 249 240 250 241 
<< m1 >>
rect 249 240 250 241 
<< m2 >>
rect 249 240 250 241 
<< m1 >>
rect 250 240 251 241 
<< m1 >>
rect 251 240 252 241 
<< m1 >>
rect 252 240 253 241 
<< m1 >>
rect 253 240 254 241 
<< m1 >>
rect 254 240 255 241 
<< m1 >>
rect 304 240 305 241 
<< m2 >>
rect 304 240 305 241 
<< m2c >>
rect 304 240 305 241 
<< m1 >>
rect 304 240 305 241 
<< m2 >>
rect 304 240 305 241 
<< m1 >>
rect 322 240 323 241 
<< m1 >>
rect 352 240 353 241 
<< m1 >>
rect 391 240 392 241 
<< m1 >>
rect 16 241 17 242 
<< m1 >>
rect 17 241 18 242 
<< m1 >>
rect 18 241 19 242 
<< m1 >>
rect 19 241 20 242 
<< m1 >>
rect 20 241 21 242 
<< m1 >>
rect 21 241 22 242 
<< m1 >>
rect 22 241 23 242 
<< m1 >>
rect 23 241 24 242 
<< m1 >>
rect 24 241 25 242 
<< m1 >>
rect 25 241 26 242 
<< m1 >>
rect 26 241 27 242 
<< m1 >>
rect 27 241 28 242 
<< m1 >>
rect 28 241 29 242 
<< m1 >>
rect 29 241 30 242 
<< m1 >>
rect 30 241 31 242 
<< m1 >>
rect 31 241 32 242 
<< m1 >>
rect 32 241 33 242 
<< m1 >>
rect 33 241 34 242 
<< m1 >>
rect 34 241 35 242 
<< m1 >>
rect 64 241 65 242 
<< m1 >>
rect 106 241 107 242 
<< m1 >>
rect 118 241 119 242 
<< m1 >>
rect 119 241 120 242 
<< m1 >>
rect 120 241 121 242 
<< m1 >>
rect 121 241 122 242 
<< m1 >>
rect 122 241 123 242 
<< m1 >>
rect 123 241 124 242 
<< m1 >>
rect 124 241 125 242 
<< m1 >>
rect 125 241 126 242 
<< m1 >>
rect 127 241 128 242 
<< m1 >>
rect 138 241 139 242 
<< m1 >>
rect 163 241 164 242 
<< m1 >>
rect 190 241 191 242 
<< m1 >>
rect 203 241 204 242 
<< m1 >>
rect 208 241 209 242 
<< m1 >>
rect 244 241 245 242 
<< m1 >>
rect 247 241 248 242 
<< m1 >>
rect 254 241 255 242 
<< m1 >>
rect 304 241 305 242 
<< m1 >>
rect 307 241 308 242 
<< m1 >>
rect 308 241 309 242 
<< m1 >>
rect 309 241 310 242 
<< m1 >>
rect 310 241 311 242 
<< m1 >>
rect 311 241 312 242 
<< m1 >>
rect 312 241 313 242 
<< m1 >>
rect 313 241 314 242 
<< m1 >>
rect 314 241 315 242 
<< m1 >>
rect 315 241 316 242 
<< m1 >>
rect 316 241 317 242 
<< m1 >>
rect 317 241 318 242 
<< m1 >>
rect 318 241 319 242 
<< m1 >>
rect 319 241 320 242 
<< m1 >>
rect 320 241 321 242 
<< m1 >>
rect 321 241 322 242 
<< m1 >>
rect 322 241 323 242 
<< m1 >>
rect 350 241 351 242 
<< m2 >>
rect 350 241 351 242 
<< m2c >>
rect 350 241 351 242 
<< m1 >>
rect 350 241 351 242 
<< m2 >>
rect 350 241 351 242 
<< m2 >>
rect 351 241 352 242 
<< m1 >>
rect 352 241 353 242 
<< m2 >>
rect 352 241 353 242 
<< m2 >>
rect 353 241 354 242 
<< m1 >>
rect 354 241 355 242 
<< m2 >>
rect 354 241 355 242 
<< m2c >>
rect 354 241 355 242 
<< m1 >>
rect 354 241 355 242 
<< m2 >>
rect 354 241 355 242 
<< m1 >>
rect 355 241 356 242 
<< m1 >>
rect 356 241 357 242 
<< m1 >>
rect 357 241 358 242 
<< m1 >>
rect 358 241 359 242 
<< m1 >>
rect 359 241 360 242 
<< m1 >>
rect 360 241 361 242 
<< m1 >>
rect 361 241 362 242 
<< m1 >>
rect 362 241 363 242 
<< m1 >>
rect 363 241 364 242 
<< m1 >>
rect 364 241 365 242 
<< m1 >>
rect 365 241 366 242 
<< m1 >>
rect 366 241 367 242 
<< m1 >>
rect 367 241 368 242 
<< m1 >>
rect 368 241 369 242 
<< m1 >>
rect 369 241 370 242 
<< m1 >>
rect 370 241 371 242 
<< m1 >>
rect 371 241 372 242 
<< m1 >>
rect 372 241 373 242 
<< m1 >>
rect 373 241 374 242 
<< m1 >>
rect 374 241 375 242 
<< m1 >>
rect 375 241 376 242 
<< m1 >>
rect 376 241 377 242 
<< m1 >>
rect 377 241 378 242 
<< m1 >>
rect 378 241 379 242 
<< m1 >>
rect 379 241 380 242 
<< m1 >>
rect 380 241 381 242 
<< m1 >>
rect 381 241 382 242 
<< m1 >>
rect 382 241 383 242 
<< m1 >>
rect 383 241 384 242 
<< m1 >>
rect 384 241 385 242 
<< m1 >>
rect 385 241 386 242 
<< m1 >>
rect 386 241 387 242 
<< m1 >>
rect 387 241 388 242 
<< m1 >>
rect 388 241 389 242 
<< m1 >>
rect 389 241 390 242 
<< m2 >>
rect 389 241 390 242 
<< m2c >>
rect 389 241 390 242 
<< m1 >>
rect 389 241 390 242 
<< m2 >>
rect 389 241 390 242 
<< m2 >>
rect 390 241 391 242 
<< m1 >>
rect 391 241 392 242 
<< m2 >>
rect 391 241 392 242 
<< m2 >>
rect 392 241 393 242 
<< m1 >>
rect 393 241 394 242 
<< m2 >>
rect 393 241 394 242 
<< m2c >>
rect 393 241 394 242 
<< m1 >>
rect 393 241 394 242 
<< m2 >>
rect 393 241 394 242 
<< m1 >>
rect 394 241 395 242 
<< m1 >>
rect 395 241 396 242 
<< m1 >>
rect 396 241 397 242 
<< m1 >>
rect 397 241 398 242 
<< m1 >>
rect 398 241 399 242 
<< m1 >>
rect 399 241 400 242 
<< m1 >>
rect 400 241 401 242 
<< m1 >>
rect 401 241 402 242 
<< m1 >>
rect 402 241 403 242 
<< m1 >>
rect 403 241 404 242 
<< m1 >>
rect 404 241 405 242 
<< m1 >>
rect 405 241 406 242 
<< m1 >>
rect 406 241 407 242 
<< m1 >>
rect 407 241 408 242 
<< m1 >>
rect 408 241 409 242 
<< m1 >>
rect 409 241 410 242 
<< m1 >>
rect 410 241 411 242 
<< m1 >>
rect 411 241 412 242 
<< m1 >>
rect 412 241 413 242 
<< m1 >>
rect 16 242 17 243 
<< m1 >>
rect 34 242 35 243 
<< m1 >>
rect 64 242 65 243 
<< m1 >>
rect 106 242 107 243 
<< m1 >>
rect 125 242 126 243 
<< m1 >>
rect 127 242 128 243 
<< m1 >>
rect 138 242 139 243 
<< m2 >>
rect 138 242 139 243 
<< m2c >>
rect 138 242 139 243 
<< m1 >>
rect 138 242 139 243 
<< m2 >>
rect 138 242 139 243 
<< m1 >>
rect 163 242 164 243 
<< m1 >>
rect 190 242 191 243 
<< m1 >>
rect 203 242 204 243 
<< m1 >>
rect 208 242 209 243 
<< m1 >>
rect 244 242 245 243 
<< m1 >>
rect 247 242 248 243 
<< m1 >>
rect 254 242 255 243 
<< m1 >>
rect 304 242 305 243 
<< m1 >>
rect 307 242 308 243 
<< m1 >>
rect 350 242 351 243 
<< m1 >>
rect 352 242 353 243 
<< m1 >>
rect 391 242 392 243 
<< m1 >>
rect 412 242 413 243 
<< m1 >>
rect 16 243 17 244 
<< m1 >>
rect 34 243 35 244 
<< m1 >>
rect 64 243 65 244 
<< m1 >>
rect 106 243 107 244 
<< m1 >>
rect 125 243 126 244 
<< m1 >>
rect 127 243 128 244 
<< m2 >>
rect 136 243 137 244 
<< m2 >>
rect 137 243 138 244 
<< m2 >>
rect 138 243 139 244 
<< m1 >>
rect 163 243 164 244 
<< m1 >>
rect 190 243 191 244 
<< m1 >>
rect 203 243 204 244 
<< m1 >>
rect 208 243 209 244 
<< m1 >>
rect 244 243 245 244 
<< m1 >>
rect 247 243 248 244 
<< m1 >>
rect 254 243 255 244 
<< m1 >>
rect 304 243 305 244 
<< m1 >>
rect 307 243 308 244 
<< m1 >>
rect 350 243 351 244 
<< m1 >>
rect 352 243 353 244 
<< m1 >>
rect 391 243 392 244 
<< m1 >>
rect 412 243 413 244 
<< m1 >>
rect 16 244 17 245 
<< m1 >>
rect 34 244 35 245 
<< m1 >>
rect 64 244 65 245 
<< m1 >>
rect 106 244 107 245 
<< m1 >>
rect 125 244 126 245 
<< m2 >>
rect 125 244 126 245 
<< m2c >>
rect 125 244 126 245 
<< m1 >>
rect 125 244 126 245 
<< m2 >>
rect 125 244 126 245 
<< m2 >>
rect 126 244 127 245 
<< m1 >>
rect 127 244 128 245 
<< m2 >>
rect 127 244 128 245 
<< m2 >>
rect 128 244 129 245 
<< m1 >>
rect 129 244 130 245 
<< m2 >>
rect 129 244 130 245 
<< m2c >>
rect 129 244 130 245 
<< m1 >>
rect 129 244 130 245 
<< m2 >>
rect 129 244 130 245 
<< m1 >>
rect 130 244 131 245 
<< m1 >>
rect 131 244 132 245 
<< m1 >>
rect 132 244 133 245 
<< m1 >>
rect 133 244 134 245 
<< m1 >>
rect 134 244 135 245 
<< m1 >>
rect 135 244 136 245 
<< m1 >>
rect 136 244 137 245 
<< m2 >>
rect 136 244 137 245 
<< m1 >>
rect 137 244 138 245 
<< m1 >>
rect 138 244 139 245 
<< m1 >>
rect 139 244 140 245 
<< m1 >>
rect 163 244 164 245 
<< m1 >>
rect 190 244 191 245 
<< m1 >>
rect 191 244 192 245 
<< m1 >>
rect 192 244 193 245 
<< m1 >>
rect 193 244 194 245 
<< m1 >>
rect 203 244 204 245 
<< m1 >>
rect 208 244 209 245 
<< m1 >>
rect 226 244 227 245 
<< m1 >>
rect 227 244 228 245 
<< m1 >>
rect 228 244 229 245 
<< m1 >>
rect 229 244 230 245 
<< m1 >>
rect 244 244 245 245 
<< m1 >>
rect 247 244 248 245 
<< m1 >>
rect 254 244 255 245 
<< m1 >>
rect 286 244 287 245 
<< m1 >>
rect 287 244 288 245 
<< m1 >>
rect 288 244 289 245 
<< m1 >>
rect 289 244 290 245 
<< m1 >>
rect 304 244 305 245 
<< m1 >>
rect 307 244 308 245 
<< m1 >>
rect 350 244 351 245 
<< m1 >>
rect 352 244 353 245 
<< m1 >>
rect 376 244 377 245 
<< m1 >>
rect 377 244 378 245 
<< m1 >>
rect 378 244 379 245 
<< m1 >>
rect 379 244 380 245 
<< m1 >>
rect 391 244 392 245 
<< m1 >>
rect 412 244 413 245 
<< m1 >>
rect 16 245 17 246 
<< m1 >>
rect 34 245 35 246 
<< m1 >>
rect 64 245 65 246 
<< m1 >>
rect 106 245 107 246 
<< m1 >>
rect 127 245 128 246 
<< m2 >>
rect 136 245 137 246 
<< m1 >>
rect 139 245 140 246 
<< m1 >>
rect 163 245 164 246 
<< m1 >>
rect 193 245 194 246 
<< m1 >>
rect 203 245 204 246 
<< m1 >>
rect 208 245 209 246 
<< m1 >>
rect 226 245 227 246 
<< m1 >>
rect 229 245 230 246 
<< m1 >>
rect 244 245 245 246 
<< m1 >>
rect 247 245 248 246 
<< m1 >>
rect 254 245 255 246 
<< m1 >>
rect 286 245 287 246 
<< m1 >>
rect 289 245 290 246 
<< m1 >>
rect 304 245 305 246 
<< m1 >>
rect 307 245 308 246 
<< m1 >>
rect 350 245 351 246 
<< m1 >>
rect 352 245 353 246 
<< m1 >>
rect 376 245 377 246 
<< m1 >>
rect 379 245 380 246 
<< m1 >>
rect 391 245 392 246 
<< m1 >>
rect 412 245 413 246 
<< pdiffusion >>
rect 12 246 13 247 
<< pdiffusion >>
rect 13 246 14 247 
<< pdiffusion >>
rect 14 246 15 247 
<< pdiffusion >>
rect 15 246 16 247 
<< m1 >>
rect 16 246 17 247 
<< pdiffusion >>
rect 16 246 17 247 
<< pdiffusion >>
rect 17 246 18 247 
<< pdiffusion >>
rect 30 246 31 247 
<< pdiffusion >>
rect 31 246 32 247 
<< pdiffusion >>
rect 32 246 33 247 
<< pdiffusion >>
rect 33 246 34 247 
<< m1 >>
rect 34 246 35 247 
<< pdiffusion >>
rect 34 246 35 247 
<< pdiffusion >>
rect 35 246 36 247 
<< pdiffusion >>
rect 48 246 49 247 
<< pdiffusion >>
rect 49 246 50 247 
<< pdiffusion >>
rect 50 246 51 247 
<< pdiffusion >>
rect 51 246 52 247 
<< pdiffusion >>
rect 52 246 53 247 
<< pdiffusion >>
rect 53 246 54 247 
<< m1 >>
rect 64 246 65 247 
<< pdiffusion >>
rect 84 246 85 247 
<< pdiffusion >>
rect 85 246 86 247 
<< pdiffusion >>
rect 86 246 87 247 
<< pdiffusion >>
rect 87 246 88 247 
<< pdiffusion >>
rect 88 246 89 247 
<< pdiffusion >>
rect 89 246 90 247 
<< pdiffusion >>
rect 102 246 103 247 
<< pdiffusion >>
rect 103 246 104 247 
<< pdiffusion >>
rect 104 246 105 247 
<< pdiffusion >>
rect 105 246 106 247 
<< m1 >>
rect 106 246 107 247 
<< pdiffusion >>
rect 106 246 107 247 
<< pdiffusion >>
rect 107 246 108 247 
<< pdiffusion >>
rect 120 246 121 247 
<< pdiffusion >>
rect 121 246 122 247 
<< pdiffusion >>
rect 122 246 123 247 
<< pdiffusion >>
rect 123 246 124 247 
<< pdiffusion >>
rect 124 246 125 247 
<< pdiffusion >>
rect 125 246 126 247 
<< m1 >>
rect 127 246 128 247 
<< m2 >>
rect 128 246 129 247 
<< m1 >>
rect 129 246 130 247 
<< m2 >>
rect 129 246 130 247 
<< m2c >>
rect 129 246 130 247 
<< m1 >>
rect 129 246 130 247 
<< m2 >>
rect 129 246 130 247 
<< m1 >>
rect 130 246 131 247 
<< m1 >>
rect 131 246 132 247 
<< m1 >>
rect 132 246 133 247 
<< m1 >>
rect 133 246 134 247 
<< m1 >>
rect 134 246 135 247 
<< m1 >>
rect 135 246 136 247 
<< m1 >>
rect 136 246 137 247 
<< m2 >>
rect 136 246 137 247 
<< m2c >>
rect 136 246 137 247 
<< m1 >>
rect 136 246 137 247 
<< m2 >>
rect 136 246 137 247 
<< pdiffusion >>
rect 138 246 139 247 
<< m1 >>
rect 139 246 140 247 
<< pdiffusion >>
rect 139 246 140 247 
<< pdiffusion >>
rect 140 246 141 247 
<< pdiffusion >>
rect 141 246 142 247 
<< pdiffusion >>
rect 142 246 143 247 
<< pdiffusion >>
rect 143 246 144 247 
<< pdiffusion >>
rect 156 246 157 247 
<< pdiffusion >>
rect 157 246 158 247 
<< pdiffusion >>
rect 158 246 159 247 
<< pdiffusion >>
rect 159 246 160 247 
<< pdiffusion >>
rect 160 246 161 247 
<< pdiffusion >>
rect 161 246 162 247 
<< m1 >>
rect 163 246 164 247 
<< pdiffusion >>
rect 174 246 175 247 
<< pdiffusion >>
rect 175 246 176 247 
<< pdiffusion >>
rect 176 246 177 247 
<< pdiffusion >>
rect 177 246 178 247 
<< pdiffusion >>
rect 178 246 179 247 
<< pdiffusion >>
rect 179 246 180 247 
<< pdiffusion >>
rect 192 246 193 247 
<< m1 >>
rect 193 246 194 247 
<< pdiffusion >>
rect 193 246 194 247 
<< pdiffusion >>
rect 194 246 195 247 
<< pdiffusion >>
rect 195 246 196 247 
<< pdiffusion >>
rect 196 246 197 247 
<< pdiffusion >>
rect 197 246 198 247 
<< m1 >>
rect 203 246 204 247 
<< m1 >>
rect 208 246 209 247 
<< pdiffusion >>
rect 210 246 211 247 
<< pdiffusion >>
rect 211 246 212 247 
<< pdiffusion >>
rect 212 246 213 247 
<< pdiffusion >>
rect 213 246 214 247 
<< pdiffusion >>
rect 214 246 215 247 
<< pdiffusion >>
rect 215 246 216 247 
<< m1 >>
rect 226 246 227 247 
<< pdiffusion >>
rect 228 246 229 247 
<< m1 >>
rect 229 246 230 247 
<< pdiffusion >>
rect 229 246 230 247 
<< pdiffusion >>
rect 230 246 231 247 
<< pdiffusion >>
rect 231 246 232 247 
<< pdiffusion >>
rect 232 246 233 247 
<< pdiffusion >>
rect 233 246 234 247 
<< m1 >>
rect 244 246 245 247 
<< pdiffusion >>
rect 246 246 247 247 
<< m1 >>
rect 247 246 248 247 
<< pdiffusion >>
rect 247 246 248 247 
<< pdiffusion >>
rect 248 246 249 247 
<< pdiffusion >>
rect 249 246 250 247 
<< pdiffusion >>
rect 250 246 251 247 
<< pdiffusion >>
rect 251 246 252 247 
<< m1 >>
rect 254 246 255 247 
<< pdiffusion >>
rect 264 246 265 247 
<< pdiffusion >>
rect 265 246 266 247 
<< pdiffusion >>
rect 266 246 267 247 
<< pdiffusion >>
rect 267 246 268 247 
<< pdiffusion >>
rect 268 246 269 247 
<< pdiffusion >>
rect 269 246 270 247 
<< pdiffusion >>
rect 282 246 283 247 
<< pdiffusion >>
rect 283 246 284 247 
<< pdiffusion >>
rect 284 246 285 247 
<< pdiffusion >>
rect 285 246 286 247 
<< m1 >>
rect 286 246 287 247 
<< pdiffusion >>
rect 286 246 287 247 
<< pdiffusion >>
rect 287 246 288 247 
<< m1 >>
rect 289 246 290 247 
<< pdiffusion >>
rect 300 246 301 247 
<< pdiffusion >>
rect 301 246 302 247 
<< pdiffusion >>
rect 302 246 303 247 
<< pdiffusion >>
rect 303 246 304 247 
<< m1 >>
rect 304 246 305 247 
<< pdiffusion >>
rect 304 246 305 247 
<< pdiffusion >>
rect 305 246 306 247 
<< m1 >>
rect 307 246 308 247 
<< pdiffusion >>
rect 318 246 319 247 
<< pdiffusion >>
rect 319 246 320 247 
<< pdiffusion >>
rect 320 246 321 247 
<< pdiffusion >>
rect 321 246 322 247 
<< pdiffusion >>
rect 322 246 323 247 
<< pdiffusion >>
rect 323 246 324 247 
<< pdiffusion >>
rect 336 246 337 247 
<< pdiffusion >>
rect 337 246 338 247 
<< pdiffusion >>
rect 338 246 339 247 
<< pdiffusion >>
rect 339 246 340 247 
<< pdiffusion >>
rect 340 246 341 247 
<< pdiffusion >>
rect 341 246 342 247 
<< m1 >>
rect 350 246 351 247 
<< m1 >>
rect 352 246 353 247 
<< pdiffusion >>
rect 354 246 355 247 
<< pdiffusion >>
rect 355 246 356 247 
<< pdiffusion >>
rect 356 246 357 247 
<< pdiffusion >>
rect 357 246 358 247 
<< pdiffusion >>
rect 358 246 359 247 
<< pdiffusion >>
rect 359 246 360 247 
<< pdiffusion >>
rect 372 246 373 247 
<< pdiffusion >>
rect 373 246 374 247 
<< pdiffusion >>
rect 374 246 375 247 
<< pdiffusion >>
rect 375 246 376 247 
<< m1 >>
rect 376 246 377 247 
<< pdiffusion >>
rect 376 246 377 247 
<< pdiffusion >>
rect 377 246 378 247 
<< m1 >>
rect 379 246 380 247 
<< pdiffusion >>
rect 390 246 391 247 
<< m1 >>
rect 391 246 392 247 
<< pdiffusion >>
rect 391 246 392 247 
<< pdiffusion >>
rect 392 246 393 247 
<< pdiffusion >>
rect 393 246 394 247 
<< pdiffusion >>
rect 394 246 395 247 
<< pdiffusion >>
rect 395 246 396 247 
<< pdiffusion >>
rect 408 246 409 247 
<< pdiffusion >>
rect 409 246 410 247 
<< pdiffusion >>
rect 410 246 411 247 
<< pdiffusion >>
rect 411 246 412 247 
<< m1 >>
rect 412 246 413 247 
<< pdiffusion >>
rect 412 246 413 247 
<< pdiffusion >>
rect 413 246 414 247 
<< pdiffusion >>
rect 426 246 427 247 
<< pdiffusion >>
rect 427 246 428 247 
<< pdiffusion >>
rect 428 246 429 247 
<< pdiffusion >>
rect 429 246 430 247 
<< pdiffusion >>
rect 430 246 431 247 
<< pdiffusion >>
rect 431 246 432 247 
<< pdiffusion >>
rect 444 246 445 247 
<< pdiffusion >>
rect 445 246 446 247 
<< pdiffusion >>
rect 446 246 447 247 
<< pdiffusion >>
rect 447 246 448 247 
<< pdiffusion >>
rect 448 246 449 247 
<< pdiffusion >>
rect 449 246 450 247 
<< pdiffusion >>
rect 12 247 13 248 
<< pdiffusion >>
rect 13 247 14 248 
<< pdiffusion >>
rect 14 247 15 248 
<< pdiffusion >>
rect 15 247 16 248 
<< pdiffusion >>
rect 16 247 17 248 
<< pdiffusion >>
rect 17 247 18 248 
<< pdiffusion >>
rect 30 247 31 248 
<< pdiffusion >>
rect 31 247 32 248 
<< pdiffusion >>
rect 32 247 33 248 
<< pdiffusion >>
rect 33 247 34 248 
<< pdiffusion >>
rect 34 247 35 248 
<< pdiffusion >>
rect 35 247 36 248 
<< pdiffusion >>
rect 48 247 49 248 
<< pdiffusion >>
rect 49 247 50 248 
<< pdiffusion >>
rect 50 247 51 248 
<< pdiffusion >>
rect 51 247 52 248 
<< pdiffusion >>
rect 52 247 53 248 
<< pdiffusion >>
rect 53 247 54 248 
<< m1 >>
rect 64 247 65 248 
<< pdiffusion >>
rect 84 247 85 248 
<< pdiffusion >>
rect 85 247 86 248 
<< pdiffusion >>
rect 86 247 87 248 
<< pdiffusion >>
rect 87 247 88 248 
<< pdiffusion >>
rect 88 247 89 248 
<< pdiffusion >>
rect 89 247 90 248 
<< pdiffusion >>
rect 102 247 103 248 
<< pdiffusion >>
rect 103 247 104 248 
<< pdiffusion >>
rect 104 247 105 248 
<< pdiffusion >>
rect 105 247 106 248 
<< pdiffusion >>
rect 106 247 107 248 
<< pdiffusion >>
rect 107 247 108 248 
<< pdiffusion >>
rect 120 247 121 248 
<< pdiffusion >>
rect 121 247 122 248 
<< pdiffusion >>
rect 122 247 123 248 
<< pdiffusion >>
rect 123 247 124 248 
<< pdiffusion >>
rect 124 247 125 248 
<< pdiffusion >>
rect 125 247 126 248 
<< m1 >>
rect 127 247 128 248 
<< m2 >>
rect 128 247 129 248 
<< pdiffusion >>
rect 138 247 139 248 
<< pdiffusion >>
rect 139 247 140 248 
<< pdiffusion >>
rect 140 247 141 248 
<< pdiffusion >>
rect 141 247 142 248 
<< pdiffusion >>
rect 142 247 143 248 
<< pdiffusion >>
rect 143 247 144 248 
<< pdiffusion >>
rect 156 247 157 248 
<< pdiffusion >>
rect 157 247 158 248 
<< pdiffusion >>
rect 158 247 159 248 
<< pdiffusion >>
rect 159 247 160 248 
<< pdiffusion >>
rect 160 247 161 248 
<< pdiffusion >>
rect 161 247 162 248 
<< m1 >>
rect 163 247 164 248 
<< pdiffusion >>
rect 174 247 175 248 
<< pdiffusion >>
rect 175 247 176 248 
<< pdiffusion >>
rect 176 247 177 248 
<< pdiffusion >>
rect 177 247 178 248 
<< pdiffusion >>
rect 178 247 179 248 
<< pdiffusion >>
rect 179 247 180 248 
<< pdiffusion >>
rect 192 247 193 248 
<< pdiffusion >>
rect 193 247 194 248 
<< pdiffusion >>
rect 194 247 195 248 
<< pdiffusion >>
rect 195 247 196 248 
<< pdiffusion >>
rect 196 247 197 248 
<< pdiffusion >>
rect 197 247 198 248 
<< m1 >>
rect 203 247 204 248 
<< m1 >>
rect 208 247 209 248 
<< pdiffusion >>
rect 210 247 211 248 
<< pdiffusion >>
rect 211 247 212 248 
<< pdiffusion >>
rect 212 247 213 248 
<< pdiffusion >>
rect 213 247 214 248 
<< pdiffusion >>
rect 214 247 215 248 
<< pdiffusion >>
rect 215 247 216 248 
<< m1 >>
rect 226 247 227 248 
<< pdiffusion >>
rect 228 247 229 248 
<< pdiffusion >>
rect 229 247 230 248 
<< pdiffusion >>
rect 230 247 231 248 
<< pdiffusion >>
rect 231 247 232 248 
<< pdiffusion >>
rect 232 247 233 248 
<< pdiffusion >>
rect 233 247 234 248 
<< m1 >>
rect 244 247 245 248 
<< pdiffusion >>
rect 246 247 247 248 
<< pdiffusion >>
rect 247 247 248 248 
<< pdiffusion >>
rect 248 247 249 248 
<< pdiffusion >>
rect 249 247 250 248 
<< pdiffusion >>
rect 250 247 251 248 
<< pdiffusion >>
rect 251 247 252 248 
<< m1 >>
rect 254 247 255 248 
<< pdiffusion >>
rect 264 247 265 248 
<< pdiffusion >>
rect 265 247 266 248 
<< pdiffusion >>
rect 266 247 267 248 
<< pdiffusion >>
rect 267 247 268 248 
<< pdiffusion >>
rect 268 247 269 248 
<< pdiffusion >>
rect 269 247 270 248 
<< pdiffusion >>
rect 282 247 283 248 
<< pdiffusion >>
rect 283 247 284 248 
<< pdiffusion >>
rect 284 247 285 248 
<< pdiffusion >>
rect 285 247 286 248 
<< pdiffusion >>
rect 286 247 287 248 
<< pdiffusion >>
rect 287 247 288 248 
<< m1 >>
rect 289 247 290 248 
<< pdiffusion >>
rect 300 247 301 248 
<< pdiffusion >>
rect 301 247 302 248 
<< pdiffusion >>
rect 302 247 303 248 
<< pdiffusion >>
rect 303 247 304 248 
<< pdiffusion >>
rect 304 247 305 248 
<< pdiffusion >>
rect 305 247 306 248 
<< m1 >>
rect 307 247 308 248 
<< pdiffusion >>
rect 318 247 319 248 
<< pdiffusion >>
rect 319 247 320 248 
<< pdiffusion >>
rect 320 247 321 248 
<< pdiffusion >>
rect 321 247 322 248 
<< pdiffusion >>
rect 322 247 323 248 
<< pdiffusion >>
rect 323 247 324 248 
<< pdiffusion >>
rect 336 247 337 248 
<< pdiffusion >>
rect 337 247 338 248 
<< pdiffusion >>
rect 338 247 339 248 
<< pdiffusion >>
rect 339 247 340 248 
<< pdiffusion >>
rect 340 247 341 248 
<< pdiffusion >>
rect 341 247 342 248 
<< m1 >>
rect 350 247 351 248 
<< m1 >>
rect 352 247 353 248 
<< pdiffusion >>
rect 354 247 355 248 
<< pdiffusion >>
rect 355 247 356 248 
<< pdiffusion >>
rect 356 247 357 248 
<< pdiffusion >>
rect 357 247 358 248 
<< pdiffusion >>
rect 358 247 359 248 
<< pdiffusion >>
rect 359 247 360 248 
<< pdiffusion >>
rect 372 247 373 248 
<< pdiffusion >>
rect 373 247 374 248 
<< pdiffusion >>
rect 374 247 375 248 
<< pdiffusion >>
rect 375 247 376 248 
<< pdiffusion >>
rect 376 247 377 248 
<< pdiffusion >>
rect 377 247 378 248 
<< m1 >>
rect 379 247 380 248 
<< pdiffusion >>
rect 390 247 391 248 
<< pdiffusion >>
rect 391 247 392 248 
<< pdiffusion >>
rect 392 247 393 248 
<< pdiffusion >>
rect 393 247 394 248 
<< pdiffusion >>
rect 394 247 395 248 
<< pdiffusion >>
rect 395 247 396 248 
<< pdiffusion >>
rect 408 247 409 248 
<< pdiffusion >>
rect 409 247 410 248 
<< pdiffusion >>
rect 410 247 411 248 
<< pdiffusion >>
rect 411 247 412 248 
<< pdiffusion >>
rect 412 247 413 248 
<< pdiffusion >>
rect 413 247 414 248 
<< pdiffusion >>
rect 426 247 427 248 
<< pdiffusion >>
rect 427 247 428 248 
<< pdiffusion >>
rect 428 247 429 248 
<< pdiffusion >>
rect 429 247 430 248 
<< pdiffusion >>
rect 430 247 431 248 
<< pdiffusion >>
rect 431 247 432 248 
<< pdiffusion >>
rect 444 247 445 248 
<< pdiffusion >>
rect 445 247 446 248 
<< pdiffusion >>
rect 446 247 447 248 
<< pdiffusion >>
rect 447 247 448 248 
<< pdiffusion >>
rect 448 247 449 248 
<< pdiffusion >>
rect 449 247 450 248 
<< pdiffusion >>
rect 12 248 13 249 
<< pdiffusion >>
rect 13 248 14 249 
<< pdiffusion >>
rect 14 248 15 249 
<< pdiffusion >>
rect 15 248 16 249 
<< pdiffusion >>
rect 16 248 17 249 
<< pdiffusion >>
rect 17 248 18 249 
<< pdiffusion >>
rect 30 248 31 249 
<< pdiffusion >>
rect 31 248 32 249 
<< pdiffusion >>
rect 32 248 33 249 
<< pdiffusion >>
rect 33 248 34 249 
<< pdiffusion >>
rect 34 248 35 249 
<< pdiffusion >>
rect 35 248 36 249 
<< pdiffusion >>
rect 48 248 49 249 
<< pdiffusion >>
rect 49 248 50 249 
<< pdiffusion >>
rect 50 248 51 249 
<< pdiffusion >>
rect 51 248 52 249 
<< pdiffusion >>
rect 52 248 53 249 
<< pdiffusion >>
rect 53 248 54 249 
<< m1 >>
rect 64 248 65 249 
<< pdiffusion >>
rect 84 248 85 249 
<< pdiffusion >>
rect 85 248 86 249 
<< pdiffusion >>
rect 86 248 87 249 
<< pdiffusion >>
rect 87 248 88 249 
<< pdiffusion >>
rect 88 248 89 249 
<< pdiffusion >>
rect 89 248 90 249 
<< pdiffusion >>
rect 102 248 103 249 
<< pdiffusion >>
rect 103 248 104 249 
<< pdiffusion >>
rect 104 248 105 249 
<< pdiffusion >>
rect 105 248 106 249 
<< pdiffusion >>
rect 106 248 107 249 
<< pdiffusion >>
rect 107 248 108 249 
<< pdiffusion >>
rect 120 248 121 249 
<< pdiffusion >>
rect 121 248 122 249 
<< pdiffusion >>
rect 122 248 123 249 
<< pdiffusion >>
rect 123 248 124 249 
<< pdiffusion >>
rect 124 248 125 249 
<< pdiffusion >>
rect 125 248 126 249 
<< m1 >>
rect 127 248 128 249 
<< m2 >>
rect 128 248 129 249 
<< pdiffusion >>
rect 138 248 139 249 
<< pdiffusion >>
rect 139 248 140 249 
<< pdiffusion >>
rect 140 248 141 249 
<< pdiffusion >>
rect 141 248 142 249 
<< pdiffusion >>
rect 142 248 143 249 
<< pdiffusion >>
rect 143 248 144 249 
<< pdiffusion >>
rect 156 248 157 249 
<< pdiffusion >>
rect 157 248 158 249 
<< pdiffusion >>
rect 158 248 159 249 
<< pdiffusion >>
rect 159 248 160 249 
<< pdiffusion >>
rect 160 248 161 249 
<< pdiffusion >>
rect 161 248 162 249 
<< m1 >>
rect 163 248 164 249 
<< pdiffusion >>
rect 174 248 175 249 
<< pdiffusion >>
rect 175 248 176 249 
<< pdiffusion >>
rect 176 248 177 249 
<< pdiffusion >>
rect 177 248 178 249 
<< pdiffusion >>
rect 178 248 179 249 
<< pdiffusion >>
rect 179 248 180 249 
<< pdiffusion >>
rect 192 248 193 249 
<< pdiffusion >>
rect 193 248 194 249 
<< pdiffusion >>
rect 194 248 195 249 
<< pdiffusion >>
rect 195 248 196 249 
<< pdiffusion >>
rect 196 248 197 249 
<< pdiffusion >>
rect 197 248 198 249 
<< m1 >>
rect 203 248 204 249 
<< m1 >>
rect 208 248 209 249 
<< pdiffusion >>
rect 210 248 211 249 
<< pdiffusion >>
rect 211 248 212 249 
<< pdiffusion >>
rect 212 248 213 249 
<< pdiffusion >>
rect 213 248 214 249 
<< pdiffusion >>
rect 214 248 215 249 
<< pdiffusion >>
rect 215 248 216 249 
<< m1 >>
rect 226 248 227 249 
<< pdiffusion >>
rect 228 248 229 249 
<< pdiffusion >>
rect 229 248 230 249 
<< pdiffusion >>
rect 230 248 231 249 
<< pdiffusion >>
rect 231 248 232 249 
<< pdiffusion >>
rect 232 248 233 249 
<< pdiffusion >>
rect 233 248 234 249 
<< m1 >>
rect 244 248 245 249 
<< pdiffusion >>
rect 246 248 247 249 
<< pdiffusion >>
rect 247 248 248 249 
<< pdiffusion >>
rect 248 248 249 249 
<< pdiffusion >>
rect 249 248 250 249 
<< pdiffusion >>
rect 250 248 251 249 
<< pdiffusion >>
rect 251 248 252 249 
<< m1 >>
rect 254 248 255 249 
<< pdiffusion >>
rect 264 248 265 249 
<< pdiffusion >>
rect 265 248 266 249 
<< pdiffusion >>
rect 266 248 267 249 
<< pdiffusion >>
rect 267 248 268 249 
<< pdiffusion >>
rect 268 248 269 249 
<< pdiffusion >>
rect 269 248 270 249 
<< pdiffusion >>
rect 282 248 283 249 
<< pdiffusion >>
rect 283 248 284 249 
<< pdiffusion >>
rect 284 248 285 249 
<< pdiffusion >>
rect 285 248 286 249 
<< pdiffusion >>
rect 286 248 287 249 
<< pdiffusion >>
rect 287 248 288 249 
<< m1 >>
rect 289 248 290 249 
<< pdiffusion >>
rect 300 248 301 249 
<< pdiffusion >>
rect 301 248 302 249 
<< pdiffusion >>
rect 302 248 303 249 
<< pdiffusion >>
rect 303 248 304 249 
<< pdiffusion >>
rect 304 248 305 249 
<< pdiffusion >>
rect 305 248 306 249 
<< m1 >>
rect 307 248 308 249 
<< pdiffusion >>
rect 318 248 319 249 
<< pdiffusion >>
rect 319 248 320 249 
<< pdiffusion >>
rect 320 248 321 249 
<< pdiffusion >>
rect 321 248 322 249 
<< pdiffusion >>
rect 322 248 323 249 
<< pdiffusion >>
rect 323 248 324 249 
<< pdiffusion >>
rect 336 248 337 249 
<< pdiffusion >>
rect 337 248 338 249 
<< pdiffusion >>
rect 338 248 339 249 
<< pdiffusion >>
rect 339 248 340 249 
<< pdiffusion >>
rect 340 248 341 249 
<< pdiffusion >>
rect 341 248 342 249 
<< m1 >>
rect 350 248 351 249 
<< m1 >>
rect 352 248 353 249 
<< pdiffusion >>
rect 354 248 355 249 
<< pdiffusion >>
rect 355 248 356 249 
<< pdiffusion >>
rect 356 248 357 249 
<< pdiffusion >>
rect 357 248 358 249 
<< pdiffusion >>
rect 358 248 359 249 
<< pdiffusion >>
rect 359 248 360 249 
<< pdiffusion >>
rect 372 248 373 249 
<< pdiffusion >>
rect 373 248 374 249 
<< pdiffusion >>
rect 374 248 375 249 
<< pdiffusion >>
rect 375 248 376 249 
<< pdiffusion >>
rect 376 248 377 249 
<< pdiffusion >>
rect 377 248 378 249 
<< m1 >>
rect 379 248 380 249 
<< pdiffusion >>
rect 390 248 391 249 
<< pdiffusion >>
rect 391 248 392 249 
<< pdiffusion >>
rect 392 248 393 249 
<< pdiffusion >>
rect 393 248 394 249 
<< pdiffusion >>
rect 394 248 395 249 
<< pdiffusion >>
rect 395 248 396 249 
<< pdiffusion >>
rect 408 248 409 249 
<< pdiffusion >>
rect 409 248 410 249 
<< pdiffusion >>
rect 410 248 411 249 
<< pdiffusion >>
rect 411 248 412 249 
<< pdiffusion >>
rect 412 248 413 249 
<< pdiffusion >>
rect 413 248 414 249 
<< pdiffusion >>
rect 426 248 427 249 
<< pdiffusion >>
rect 427 248 428 249 
<< pdiffusion >>
rect 428 248 429 249 
<< pdiffusion >>
rect 429 248 430 249 
<< pdiffusion >>
rect 430 248 431 249 
<< pdiffusion >>
rect 431 248 432 249 
<< pdiffusion >>
rect 444 248 445 249 
<< pdiffusion >>
rect 445 248 446 249 
<< pdiffusion >>
rect 446 248 447 249 
<< pdiffusion >>
rect 447 248 448 249 
<< pdiffusion >>
rect 448 248 449 249 
<< pdiffusion >>
rect 449 248 450 249 
<< pdiffusion >>
rect 12 249 13 250 
<< pdiffusion >>
rect 13 249 14 250 
<< pdiffusion >>
rect 14 249 15 250 
<< pdiffusion >>
rect 15 249 16 250 
<< pdiffusion >>
rect 16 249 17 250 
<< pdiffusion >>
rect 17 249 18 250 
<< pdiffusion >>
rect 30 249 31 250 
<< pdiffusion >>
rect 31 249 32 250 
<< pdiffusion >>
rect 32 249 33 250 
<< pdiffusion >>
rect 33 249 34 250 
<< pdiffusion >>
rect 34 249 35 250 
<< pdiffusion >>
rect 35 249 36 250 
<< pdiffusion >>
rect 48 249 49 250 
<< pdiffusion >>
rect 49 249 50 250 
<< pdiffusion >>
rect 50 249 51 250 
<< pdiffusion >>
rect 51 249 52 250 
<< pdiffusion >>
rect 52 249 53 250 
<< pdiffusion >>
rect 53 249 54 250 
<< m1 >>
rect 64 249 65 250 
<< pdiffusion >>
rect 84 249 85 250 
<< pdiffusion >>
rect 85 249 86 250 
<< pdiffusion >>
rect 86 249 87 250 
<< pdiffusion >>
rect 87 249 88 250 
<< pdiffusion >>
rect 88 249 89 250 
<< pdiffusion >>
rect 89 249 90 250 
<< pdiffusion >>
rect 102 249 103 250 
<< pdiffusion >>
rect 103 249 104 250 
<< pdiffusion >>
rect 104 249 105 250 
<< pdiffusion >>
rect 105 249 106 250 
<< pdiffusion >>
rect 106 249 107 250 
<< pdiffusion >>
rect 107 249 108 250 
<< pdiffusion >>
rect 120 249 121 250 
<< pdiffusion >>
rect 121 249 122 250 
<< pdiffusion >>
rect 122 249 123 250 
<< pdiffusion >>
rect 123 249 124 250 
<< pdiffusion >>
rect 124 249 125 250 
<< pdiffusion >>
rect 125 249 126 250 
<< m1 >>
rect 127 249 128 250 
<< m2 >>
rect 128 249 129 250 
<< pdiffusion >>
rect 138 249 139 250 
<< pdiffusion >>
rect 139 249 140 250 
<< pdiffusion >>
rect 140 249 141 250 
<< pdiffusion >>
rect 141 249 142 250 
<< pdiffusion >>
rect 142 249 143 250 
<< pdiffusion >>
rect 143 249 144 250 
<< pdiffusion >>
rect 156 249 157 250 
<< pdiffusion >>
rect 157 249 158 250 
<< pdiffusion >>
rect 158 249 159 250 
<< pdiffusion >>
rect 159 249 160 250 
<< pdiffusion >>
rect 160 249 161 250 
<< pdiffusion >>
rect 161 249 162 250 
<< m1 >>
rect 163 249 164 250 
<< pdiffusion >>
rect 174 249 175 250 
<< pdiffusion >>
rect 175 249 176 250 
<< pdiffusion >>
rect 176 249 177 250 
<< pdiffusion >>
rect 177 249 178 250 
<< pdiffusion >>
rect 178 249 179 250 
<< pdiffusion >>
rect 179 249 180 250 
<< pdiffusion >>
rect 192 249 193 250 
<< pdiffusion >>
rect 193 249 194 250 
<< pdiffusion >>
rect 194 249 195 250 
<< pdiffusion >>
rect 195 249 196 250 
<< pdiffusion >>
rect 196 249 197 250 
<< pdiffusion >>
rect 197 249 198 250 
<< m1 >>
rect 203 249 204 250 
<< m1 >>
rect 208 249 209 250 
<< pdiffusion >>
rect 210 249 211 250 
<< pdiffusion >>
rect 211 249 212 250 
<< pdiffusion >>
rect 212 249 213 250 
<< pdiffusion >>
rect 213 249 214 250 
<< pdiffusion >>
rect 214 249 215 250 
<< pdiffusion >>
rect 215 249 216 250 
<< m1 >>
rect 226 249 227 250 
<< pdiffusion >>
rect 228 249 229 250 
<< pdiffusion >>
rect 229 249 230 250 
<< pdiffusion >>
rect 230 249 231 250 
<< pdiffusion >>
rect 231 249 232 250 
<< pdiffusion >>
rect 232 249 233 250 
<< pdiffusion >>
rect 233 249 234 250 
<< m1 >>
rect 244 249 245 250 
<< pdiffusion >>
rect 246 249 247 250 
<< pdiffusion >>
rect 247 249 248 250 
<< pdiffusion >>
rect 248 249 249 250 
<< pdiffusion >>
rect 249 249 250 250 
<< pdiffusion >>
rect 250 249 251 250 
<< pdiffusion >>
rect 251 249 252 250 
<< m1 >>
rect 254 249 255 250 
<< pdiffusion >>
rect 264 249 265 250 
<< pdiffusion >>
rect 265 249 266 250 
<< pdiffusion >>
rect 266 249 267 250 
<< pdiffusion >>
rect 267 249 268 250 
<< pdiffusion >>
rect 268 249 269 250 
<< pdiffusion >>
rect 269 249 270 250 
<< pdiffusion >>
rect 282 249 283 250 
<< pdiffusion >>
rect 283 249 284 250 
<< pdiffusion >>
rect 284 249 285 250 
<< pdiffusion >>
rect 285 249 286 250 
<< pdiffusion >>
rect 286 249 287 250 
<< pdiffusion >>
rect 287 249 288 250 
<< m1 >>
rect 289 249 290 250 
<< pdiffusion >>
rect 300 249 301 250 
<< pdiffusion >>
rect 301 249 302 250 
<< pdiffusion >>
rect 302 249 303 250 
<< pdiffusion >>
rect 303 249 304 250 
<< pdiffusion >>
rect 304 249 305 250 
<< pdiffusion >>
rect 305 249 306 250 
<< m1 >>
rect 307 249 308 250 
<< pdiffusion >>
rect 318 249 319 250 
<< pdiffusion >>
rect 319 249 320 250 
<< pdiffusion >>
rect 320 249 321 250 
<< pdiffusion >>
rect 321 249 322 250 
<< pdiffusion >>
rect 322 249 323 250 
<< pdiffusion >>
rect 323 249 324 250 
<< pdiffusion >>
rect 336 249 337 250 
<< pdiffusion >>
rect 337 249 338 250 
<< pdiffusion >>
rect 338 249 339 250 
<< pdiffusion >>
rect 339 249 340 250 
<< pdiffusion >>
rect 340 249 341 250 
<< pdiffusion >>
rect 341 249 342 250 
<< m1 >>
rect 350 249 351 250 
<< m1 >>
rect 352 249 353 250 
<< pdiffusion >>
rect 354 249 355 250 
<< pdiffusion >>
rect 355 249 356 250 
<< pdiffusion >>
rect 356 249 357 250 
<< pdiffusion >>
rect 357 249 358 250 
<< pdiffusion >>
rect 358 249 359 250 
<< pdiffusion >>
rect 359 249 360 250 
<< pdiffusion >>
rect 372 249 373 250 
<< pdiffusion >>
rect 373 249 374 250 
<< pdiffusion >>
rect 374 249 375 250 
<< pdiffusion >>
rect 375 249 376 250 
<< pdiffusion >>
rect 376 249 377 250 
<< pdiffusion >>
rect 377 249 378 250 
<< m1 >>
rect 379 249 380 250 
<< pdiffusion >>
rect 390 249 391 250 
<< pdiffusion >>
rect 391 249 392 250 
<< pdiffusion >>
rect 392 249 393 250 
<< pdiffusion >>
rect 393 249 394 250 
<< pdiffusion >>
rect 394 249 395 250 
<< pdiffusion >>
rect 395 249 396 250 
<< pdiffusion >>
rect 408 249 409 250 
<< pdiffusion >>
rect 409 249 410 250 
<< pdiffusion >>
rect 410 249 411 250 
<< pdiffusion >>
rect 411 249 412 250 
<< pdiffusion >>
rect 412 249 413 250 
<< pdiffusion >>
rect 413 249 414 250 
<< pdiffusion >>
rect 426 249 427 250 
<< pdiffusion >>
rect 427 249 428 250 
<< pdiffusion >>
rect 428 249 429 250 
<< pdiffusion >>
rect 429 249 430 250 
<< pdiffusion >>
rect 430 249 431 250 
<< pdiffusion >>
rect 431 249 432 250 
<< pdiffusion >>
rect 444 249 445 250 
<< pdiffusion >>
rect 445 249 446 250 
<< pdiffusion >>
rect 446 249 447 250 
<< pdiffusion >>
rect 447 249 448 250 
<< pdiffusion >>
rect 448 249 449 250 
<< pdiffusion >>
rect 449 249 450 250 
<< pdiffusion >>
rect 12 250 13 251 
<< pdiffusion >>
rect 13 250 14 251 
<< pdiffusion >>
rect 14 250 15 251 
<< pdiffusion >>
rect 15 250 16 251 
<< pdiffusion >>
rect 16 250 17 251 
<< pdiffusion >>
rect 17 250 18 251 
<< pdiffusion >>
rect 30 250 31 251 
<< pdiffusion >>
rect 31 250 32 251 
<< pdiffusion >>
rect 32 250 33 251 
<< pdiffusion >>
rect 33 250 34 251 
<< pdiffusion >>
rect 34 250 35 251 
<< pdiffusion >>
rect 35 250 36 251 
<< pdiffusion >>
rect 48 250 49 251 
<< pdiffusion >>
rect 49 250 50 251 
<< pdiffusion >>
rect 50 250 51 251 
<< pdiffusion >>
rect 51 250 52 251 
<< pdiffusion >>
rect 52 250 53 251 
<< pdiffusion >>
rect 53 250 54 251 
<< m1 >>
rect 64 250 65 251 
<< pdiffusion >>
rect 84 250 85 251 
<< pdiffusion >>
rect 85 250 86 251 
<< pdiffusion >>
rect 86 250 87 251 
<< pdiffusion >>
rect 87 250 88 251 
<< pdiffusion >>
rect 88 250 89 251 
<< pdiffusion >>
rect 89 250 90 251 
<< pdiffusion >>
rect 102 250 103 251 
<< pdiffusion >>
rect 103 250 104 251 
<< pdiffusion >>
rect 104 250 105 251 
<< pdiffusion >>
rect 105 250 106 251 
<< pdiffusion >>
rect 106 250 107 251 
<< pdiffusion >>
rect 107 250 108 251 
<< pdiffusion >>
rect 120 250 121 251 
<< pdiffusion >>
rect 121 250 122 251 
<< pdiffusion >>
rect 122 250 123 251 
<< pdiffusion >>
rect 123 250 124 251 
<< pdiffusion >>
rect 124 250 125 251 
<< pdiffusion >>
rect 125 250 126 251 
<< m1 >>
rect 127 250 128 251 
<< m2 >>
rect 128 250 129 251 
<< pdiffusion >>
rect 138 250 139 251 
<< pdiffusion >>
rect 139 250 140 251 
<< pdiffusion >>
rect 140 250 141 251 
<< pdiffusion >>
rect 141 250 142 251 
<< pdiffusion >>
rect 142 250 143 251 
<< pdiffusion >>
rect 143 250 144 251 
<< pdiffusion >>
rect 156 250 157 251 
<< pdiffusion >>
rect 157 250 158 251 
<< pdiffusion >>
rect 158 250 159 251 
<< pdiffusion >>
rect 159 250 160 251 
<< pdiffusion >>
rect 160 250 161 251 
<< pdiffusion >>
rect 161 250 162 251 
<< m1 >>
rect 163 250 164 251 
<< pdiffusion >>
rect 174 250 175 251 
<< pdiffusion >>
rect 175 250 176 251 
<< pdiffusion >>
rect 176 250 177 251 
<< pdiffusion >>
rect 177 250 178 251 
<< pdiffusion >>
rect 178 250 179 251 
<< pdiffusion >>
rect 179 250 180 251 
<< pdiffusion >>
rect 192 250 193 251 
<< pdiffusion >>
rect 193 250 194 251 
<< pdiffusion >>
rect 194 250 195 251 
<< pdiffusion >>
rect 195 250 196 251 
<< pdiffusion >>
rect 196 250 197 251 
<< pdiffusion >>
rect 197 250 198 251 
<< m1 >>
rect 203 250 204 251 
<< m1 >>
rect 208 250 209 251 
<< pdiffusion >>
rect 210 250 211 251 
<< pdiffusion >>
rect 211 250 212 251 
<< pdiffusion >>
rect 212 250 213 251 
<< pdiffusion >>
rect 213 250 214 251 
<< pdiffusion >>
rect 214 250 215 251 
<< pdiffusion >>
rect 215 250 216 251 
<< m1 >>
rect 226 250 227 251 
<< pdiffusion >>
rect 228 250 229 251 
<< pdiffusion >>
rect 229 250 230 251 
<< pdiffusion >>
rect 230 250 231 251 
<< pdiffusion >>
rect 231 250 232 251 
<< pdiffusion >>
rect 232 250 233 251 
<< pdiffusion >>
rect 233 250 234 251 
<< m1 >>
rect 244 250 245 251 
<< pdiffusion >>
rect 246 250 247 251 
<< pdiffusion >>
rect 247 250 248 251 
<< pdiffusion >>
rect 248 250 249 251 
<< pdiffusion >>
rect 249 250 250 251 
<< pdiffusion >>
rect 250 250 251 251 
<< pdiffusion >>
rect 251 250 252 251 
<< m1 >>
rect 254 250 255 251 
<< pdiffusion >>
rect 264 250 265 251 
<< pdiffusion >>
rect 265 250 266 251 
<< pdiffusion >>
rect 266 250 267 251 
<< pdiffusion >>
rect 267 250 268 251 
<< pdiffusion >>
rect 268 250 269 251 
<< pdiffusion >>
rect 269 250 270 251 
<< pdiffusion >>
rect 282 250 283 251 
<< pdiffusion >>
rect 283 250 284 251 
<< pdiffusion >>
rect 284 250 285 251 
<< pdiffusion >>
rect 285 250 286 251 
<< pdiffusion >>
rect 286 250 287 251 
<< pdiffusion >>
rect 287 250 288 251 
<< m1 >>
rect 289 250 290 251 
<< pdiffusion >>
rect 300 250 301 251 
<< pdiffusion >>
rect 301 250 302 251 
<< pdiffusion >>
rect 302 250 303 251 
<< pdiffusion >>
rect 303 250 304 251 
<< pdiffusion >>
rect 304 250 305 251 
<< pdiffusion >>
rect 305 250 306 251 
<< m1 >>
rect 307 250 308 251 
<< pdiffusion >>
rect 318 250 319 251 
<< pdiffusion >>
rect 319 250 320 251 
<< pdiffusion >>
rect 320 250 321 251 
<< pdiffusion >>
rect 321 250 322 251 
<< pdiffusion >>
rect 322 250 323 251 
<< pdiffusion >>
rect 323 250 324 251 
<< pdiffusion >>
rect 336 250 337 251 
<< pdiffusion >>
rect 337 250 338 251 
<< pdiffusion >>
rect 338 250 339 251 
<< pdiffusion >>
rect 339 250 340 251 
<< pdiffusion >>
rect 340 250 341 251 
<< pdiffusion >>
rect 341 250 342 251 
<< m1 >>
rect 350 250 351 251 
<< m1 >>
rect 352 250 353 251 
<< pdiffusion >>
rect 354 250 355 251 
<< pdiffusion >>
rect 355 250 356 251 
<< pdiffusion >>
rect 356 250 357 251 
<< pdiffusion >>
rect 357 250 358 251 
<< pdiffusion >>
rect 358 250 359 251 
<< pdiffusion >>
rect 359 250 360 251 
<< pdiffusion >>
rect 372 250 373 251 
<< pdiffusion >>
rect 373 250 374 251 
<< pdiffusion >>
rect 374 250 375 251 
<< pdiffusion >>
rect 375 250 376 251 
<< pdiffusion >>
rect 376 250 377 251 
<< pdiffusion >>
rect 377 250 378 251 
<< m1 >>
rect 379 250 380 251 
<< pdiffusion >>
rect 390 250 391 251 
<< pdiffusion >>
rect 391 250 392 251 
<< pdiffusion >>
rect 392 250 393 251 
<< pdiffusion >>
rect 393 250 394 251 
<< pdiffusion >>
rect 394 250 395 251 
<< pdiffusion >>
rect 395 250 396 251 
<< pdiffusion >>
rect 408 250 409 251 
<< pdiffusion >>
rect 409 250 410 251 
<< pdiffusion >>
rect 410 250 411 251 
<< pdiffusion >>
rect 411 250 412 251 
<< pdiffusion >>
rect 412 250 413 251 
<< pdiffusion >>
rect 413 250 414 251 
<< pdiffusion >>
rect 426 250 427 251 
<< pdiffusion >>
rect 427 250 428 251 
<< pdiffusion >>
rect 428 250 429 251 
<< pdiffusion >>
rect 429 250 430 251 
<< pdiffusion >>
rect 430 250 431 251 
<< pdiffusion >>
rect 431 250 432 251 
<< pdiffusion >>
rect 444 250 445 251 
<< pdiffusion >>
rect 445 250 446 251 
<< pdiffusion >>
rect 446 250 447 251 
<< pdiffusion >>
rect 447 250 448 251 
<< pdiffusion >>
rect 448 250 449 251 
<< pdiffusion >>
rect 449 250 450 251 
<< pdiffusion >>
rect 12 251 13 252 
<< pdiffusion >>
rect 13 251 14 252 
<< pdiffusion >>
rect 14 251 15 252 
<< pdiffusion >>
rect 15 251 16 252 
<< pdiffusion >>
rect 16 251 17 252 
<< pdiffusion >>
rect 17 251 18 252 
<< pdiffusion >>
rect 30 251 31 252 
<< pdiffusion >>
rect 31 251 32 252 
<< pdiffusion >>
rect 32 251 33 252 
<< pdiffusion >>
rect 33 251 34 252 
<< pdiffusion >>
rect 34 251 35 252 
<< pdiffusion >>
rect 35 251 36 252 
<< pdiffusion >>
rect 48 251 49 252 
<< pdiffusion >>
rect 49 251 50 252 
<< pdiffusion >>
rect 50 251 51 252 
<< pdiffusion >>
rect 51 251 52 252 
<< pdiffusion >>
rect 52 251 53 252 
<< pdiffusion >>
rect 53 251 54 252 
<< m1 >>
rect 64 251 65 252 
<< pdiffusion >>
rect 84 251 85 252 
<< pdiffusion >>
rect 85 251 86 252 
<< pdiffusion >>
rect 86 251 87 252 
<< pdiffusion >>
rect 87 251 88 252 
<< pdiffusion >>
rect 88 251 89 252 
<< pdiffusion >>
rect 89 251 90 252 
<< pdiffusion >>
rect 102 251 103 252 
<< pdiffusion >>
rect 103 251 104 252 
<< pdiffusion >>
rect 104 251 105 252 
<< pdiffusion >>
rect 105 251 106 252 
<< pdiffusion >>
rect 106 251 107 252 
<< pdiffusion >>
rect 107 251 108 252 
<< pdiffusion >>
rect 120 251 121 252 
<< m1 >>
rect 121 251 122 252 
<< pdiffusion >>
rect 121 251 122 252 
<< pdiffusion >>
rect 122 251 123 252 
<< pdiffusion >>
rect 123 251 124 252 
<< pdiffusion >>
rect 124 251 125 252 
<< pdiffusion >>
rect 125 251 126 252 
<< m1 >>
rect 127 251 128 252 
<< m2 >>
rect 128 251 129 252 
<< pdiffusion >>
rect 138 251 139 252 
<< pdiffusion >>
rect 139 251 140 252 
<< pdiffusion >>
rect 140 251 141 252 
<< pdiffusion >>
rect 141 251 142 252 
<< pdiffusion >>
rect 142 251 143 252 
<< pdiffusion >>
rect 143 251 144 252 
<< pdiffusion >>
rect 156 251 157 252 
<< pdiffusion >>
rect 157 251 158 252 
<< pdiffusion >>
rect 158 251 159 252 
<< pdiffusion >>
rect 159 251 160 252 
<< pdiffusion >>
rect 160 251 161 252 
<< pdiffusion >>
rect 161 251 162 252 
<< m1 >>
rect 163 251 164 252 
<< pdiffusion >>
rect 174 251 175 252 
<< pdiffusion >>
rect 175 251 176 252 
<< pdiffusion >>
rect 176 251 177 252 
<< pdiffusion >>
rect 177 251 178 252 
<< pdiffusion >>
rect 178 251 179 252 
<< pdiffusion >>
rect 179 251 180 252 
<< pdiffusion >>
rect 192 251 193 252 
<< pdiffusion >>
rect 193 251 194 252 
<< pdiffusion >>
rect 194 251 195 252 
<< pdiffusion >>
rect 195 251 196 252 
<< pdiffusion >>
rect 196 251 197 252 
<< pdiffusion >>
rect 197 251 198 252 
<< m1 >>
rect 203 251 204 252 
<< m1 >>
rect 208 251 209 252 
<< pdiffusion >>
rect 210 251 211 252 
<< m1 >>
rect 211 251 212 252 
<< pdiffusion >>
rect 211 251 212 252 
<< pdiffusion >>
rect 212 251 213 252 
<< pdiffusion >>
rect 213 251 214 252 
<< pdiffusion >>
rect 214 251 215 252 
<< pdiffusion >>
rect 215 251 216 252 
<< m1 >>
rect 226 251 227 252 
<< pdiffusion >>
rect 228 251 229 252 
<< pdiffusion >>
rect 229 251 230 252 
<< pdiffusion >>
rect 230 251 231 252 
<< pdiffusion >>
rect 231 251 232 252 
<< pdiffusion >>
rect 232 251 233 252 
<< pdiffusion >>
rect 233 251 234 252 
<< m1 >>
rect 244 251 245 252 
<< pdiffusion >>
rect 246 251 247 252 
<< pdiffusion >>
rect 247 251 248 252 
<< pdiffusion >>
rect 248 251 249 252 
<< pdiffusion >>
rect 249 251 250 252 
<< m1 >>
rect 250 251 251 252 
<< pdiffusion >>
rect 250 251 251 252 
<< pdiffusion >>
rect 251 251 252 252 
<< m1 >>
rect 254 251 255 252 
<< pdiffusion >>
rect 264 251 265 252 
<< pdiffusion >>
rect 265 251 266 252 
<< pdiffusion >>
rect 266 251 267 252 
<< pdiffusion >>
rect 267 251 268 252 
<< pdiffusion >>
rect 268 251 269 252 
<< pdiffusion >>
rect 269 251 270 252 
<< pdiffusion >>
rect 282 251 283 252 
<< pdiffusion >>
rect 283 251 284 252 
<< pdiffusion >>
rect 284 251 285 252 
<< pdiffusion >>
rect 285 251 286 252 
<< pdiffusion >>
rect 286 251 287 252 
<< pdiffusion >>
rect 287 251 288 252 
<< m1 >>
rect 289 251 290 252 
<< pdiffusion >>
rect 300 251 301 252 
<< m1 >>
rect 301 251 302 252 
<< pdiffusion >>
rect 301 251 302 252 
<< pdiffusion >>
rect 302 251 303 252 
<< pdiffusion >>
rect 303 251 304 252 
<< pdiffusion >>
rect 304 251 305 252 
<< pdiffusion >>
rect 305 251 306 252 
<< m1 >>
rect 307 251 308 252 
<< pdiffusion >>
rect 318 251 319 252 
<< pdiffusion >>
rect 319 251 320 252 
<< pdiffusion >>
rect 320 251 321 252 
<< pdiffusion >>
rect 321 251 322 252 
<< pdiffusion >>
rect 322 251 323 252 
<< pdiffusion >>
rect 323 251 324 252 
<< pdiffusion >>
rect 336 251 337 252 
<< m1 >>
rect 337 251 338 252 
<< pdiffusion >>
rect 337 251 338 252 
<< pdiffusion >>
rect 338 251 339 252 
<< pdiffusion >>
rect 339 251 340 252 
<< pdiffusion >>
rect 340 251 341 252 
<< pdiffusion >>
rect 341 251 342 252 
<< m1 >>
rect 350 251 351 252 
<< m1 >>
rect 352 251 353 252 
<< pdiffusion >>
rect 354 251 355 252 
<< pdiffusion >>
rect 355 251 356 252 
<< pdiffusion >>
rect 356 251 357 252 
<< pdiffusion >>
rect 357 251 358 252 
<< pdiffusion >>
rect 358 251 359 252 
<< pdiffusion >>
rect 359 251 360 252 
<< pdiffusion >>
rect 372 251 373 252 
<< m1 >>
rect 373 251 374 252 
<< pdiffusion >>
rect 373 251 374 252 
<< pdiffusion >>
rect 374 251 375 252 
<< pdiffusion >>
rect 375 251 376 252 
<< pdiffusion >>
rect 376 251 377 252 
<< pdiffusion >>
rect 377 251 378 252 
<< m1 >>
rect 379 251 380 252 
<< pdiffusion >>
rect 390 251 391 252 
<< pdiffusion >>
rect 391 251 392 252 
<< pdiffusion >>
rect 392 251 393 252 
<< pdiffusion >>
rect 393 251 394 252 
<< pdiffusion >>
rect 394 251 395 252 
<< pdiffusion >>
rect 395 251 396 252 
<< pdiffusion >>
rect 408 251 409 252 
<< pdiffusion >>
rect 409 251 410 252 
<< pdiffusion >>
rect 410 251 411 252 
<< pdiffusion >>
rect 411 251 412 252 
<< pdiffusion >>
rect 412 251 413 252 
<< pdiffusion >>
rect 413 251 414 252 
<< pdiffusion >>
rect 426 251 427 252 
<< pdiffusion >>
rect 427 251 428 252 
<< pdiffusion >>
rect 428 251 429 252 
<< pdiffusion >>
rect 429 251 430 252 
<< pdiffusion >>
rect 430 251 431 252 
<< pdiffusion >>
rect 431 251 432 252 
<< pdiffusion >>
rect 444 251 445 252 
<< pdiffusion >>
rect 445 251 446 252 
<< pdiffusion >>
rect 446 251 447 252 
<< pdiffusion >>
rect 447 251 448 252 
<< pdiffusion >>
rect 448 251 449 252 
<< pdiffusion >>
rect 449 251 450 252 
<< m1 >>
rect 64 252 65 253 
<< m1 >>
rect 121 252 122 253 
<< m1 >>
rect 127 252 128 253 
<< m2 >>
rect 128 252 129 253 
<< m1 >>
rect 163 252 164 253 
<< m1 >>
rect 203 252 204 253 
<< m1 >>
rect 208 252 209 253 
<< m1 >>
rect 211 252 212 253 
<< m1 >>
rect 226 252 227 253 
<< m1 >>
rect 244 252 245 253 
<< m1 >>
rect 250 252 251 253 
<< m1 >>
rect 254 252 255 253 
<< m1 >>
rect 289 252 290 253 
<< m1 >>
rect 301 252 302 253 
<< m1 >>
rect 307 252 308 253 
<< m2 >>
rect 307 252 308 253 
<< m2c >>
rect 307 252 308 253 
<< m1 >>
rect 307 252 308 253 
<< m2 >>
rect 307 252 308 253 
<< m1 >>
rect 337 252 338 253 
<< m1 >>
rect 350 252 351 253 
<< m1 >>
rect 352 252 353 253 
<< m1 >>
rect 373 252 374 253 
<< m1 >>
rect 379 252 380 253 
<< m1 >>
rect 64 253 65 254 
<< m1 >>
rect 121 253 122 254 
<< m1 >>
rect 125 253 126 254 
<< m2 >>
rect 125 253 126 254 
<< m2c >>
rect 125 253 126 254 
<< m1 >>
rect 125 253 126 254 
<< m2 >>
rect 125 253 126 254 
<< m2 >>
rect 126 253 127 254 
<< m1 >>
rect 127 253 128 254 
<< m2 >>
rect 127 253 128 254 
<< m2 >>
rect 128 253 129 254 
<< m1 >>
rect 163 253 164 254 
<< m1 >>
rect 203 253 204 254 
<< m1 >>
rect 208 253 209 254 
<< m1 >>
rect 211 253 212 254 
<< m1 >>
rect 226 253 227 254 
<< m1 >>
rect 244 253 245 254 
<< m1 >>
rect 250 253 251 254 
<< m1 >>
rect 254 253 255 254 
<< m1 >>
rect 289 253 290 254 
<< m1 >>
rect 301 253 302 254 
<< m2 >>
rect 307 253 308 254 
<< m1 >>
rect 337 253 338 254 
<< m1 >>
rect 350 253 351 254 
<< m1 >>
rect 352 253 353 254 
<< m1 >>
rect 373 253 374 254 
<< m1 >>
rect 379 253 380 254 
<< m1 >>
rect 64 254 65 255 
<< m1 >>
rect 121 254 122 255 
<< m1 >>
rect 122 254 123 255 
<< m1 >>
rect 123 254 124 255 
<< m1 >>
rect 124 254 125 255 
<< m1 >>
rect 125 254 126 255 
<< m1 >>
rect 127 254 128 255 
<< m1 >>
rect 163 254 164 255 
<< m1 >>
rect 203 254 204 255 
<< m1 >>
rect 208 254 209 255 
<< m1 >>
rect 211 254 212 255 
<< m1 >>
rect 212 254 213 255 
<< m1 >>
rect 213 254 214 255 
<< m1 >>
rect 214 254 215 255 
<< m1 >>
rect 215 254 216 255 
<< m1 >>
rect 216 254 217 255 
<< m1 >>
rect 217 254 218 255 
<< m1 >>
rect 218 254 219 255 
<< m1 >>
rect 219 254 220 255 
<< m1 >>
rect 220 254 221 255 
<< m1 >>
rect 221 254 222 255 
<< m1 >>
rect 222 254 223 255 
<< m1 >>
rect 223 254 224 255 
<< m1 >>
rect 224 254 225 255 
<< m1 >>
rect 225 254 226 255 
<< m1 >>
rect 226 254 227 255 
<< m1 >>
rect 244 254 245 255 
<< m1 >>
rect 250 254 251 255 
<< m1 >>
rect 254 254 255 255 
<< m1 >>
rect 289 254 290 255 
<< m1 >>
rect 301 254 302 255 
<< m1 >>
rect 302 254 303 255 
<< m1 >>
rect 303 254 304 255 
<< m1 >>
rect 304 254 305 255 
<< m1 >>
rect 305 254 306 255 
<< m1 >>
rect 306 254 307 255 
<< m1 >>
rect 307 254 308 255 
<< m2 >>
rect 307 254 308 255 
<< m1 >>
rect 337 254 338 255 
<< m1 >>
rect 350 254 351 255 
<< m1 >>
rect 352 254 353 255 
<< m1 >>
rect 373 254 374 255 
<< m1 >>
rect 379 254 380 255 
<< m1 >>
rect 64 255 65 256 
<< m1 >>
rect 127 255 128 256 
<< m1 >>
rect 163 255 164 256 
<< m1 >>
rect 203 255 204 256 
<< m1 >>
rect 208 255 209 256 
<< m1 >>
rect 244 255 245 256 
<< m1 >>
rect 250 255 251 256 
<< m1 >>
rect 254 255 255 256 
<< m1 >>
rect 289 255 290 256 
<< m1 >>
rect 307 255 308 256 
<< m2 >>
rect 307 255 308 256 
<< m1 >>
rect 337 255 338 256 
<< m1 >>
rect 350 255 351 256 
<< m1 >>
rect 352 255 353 256 
<< m1 >>
rect 373 255 374 256 
<< m1 >>
rect 379 255 380 256 
<< m1 >>
rect 64 256 65 257 
<< m1 >>
rect 127 256 128 257 
<< m1 >>
rect 163 256 164 257 
<< m1 >>
rect 203 256 204 257 
<< m1 >>
rect 208 256 209 257 
<< m1 >>
rect 244 256 245 257 
<< m1 >>
rect 250 256 251 257 
<< m1 >>
rect 254 256 255 257 
<< m1 >>
rect 282 256 283 257 
<< m1 >>
rect 283 256 284 257 
<< m1 >>
rect 284 256 285 257 
<< m1 >>
rect 285 256 286 257 
<< m1 >>
rect 286 256 287 257 
<< m1 >>
rect 287 256 288 257 
<< m1 >>
rect 288 256 289 257 
<< m1 >>
rect 289 256 290 257 
<< m1 >>
rect 307 256 308 257 
<< m2 >>
rect 307 256 308 257 
<< m1 >>
rect 337 256 338 257 
<< m1 >>
rect 350 256 351 257 
<< m1 >>
rect 352 256 353 257 
<< m1 >>
rect 373 256 374 257 
<< m1 >>
rect 379 256 380 257 
<< m1 >>
rect 64 257 65 258 
<< m1 >>
rect 127 257 128 258 
<< m1 >>
rect 163 257 164 258 
<< m1 >>
rect 203 257 204 258 
<< m1 >>
rect 208 257 209 258 
<< m1 >>
rect 244 257 245 258 
<< m1 >>
rect 250 257 251 258 
<< m1 >>
rect 254 257 255 258 
<< m1 >>
rect 282 257 283 258 
<< m1 >>
rect 307 257 308 258 
<< m2 >>
rect 307 257 308 258 
<< m1 >>
rect 337 257 338 258 
<< m1 >>
rect 350 257 351 258 
<< m2 >>
rect 350 257 351 258 
<< m2c >>
rect 350 257 351 258 
<< m1 >>
rect 350 257 351 258 
<< m2 >>
rect 350 257 351 258 
<< m1 >>
rect 352 257 353 258 
<< m2 >>
rect 352 257 353 258 
<< m2c >>
rect 352 257 353 258 
<< m1 >>
rect 352 257 353 258 
<< m2 >>
rect 352 257 353 258 
<< m1 >>
rect 373 257 374 258 
<< m1 >>
rect 379 257 380 258 
<< m1 >>
rect 64 258 65 259 
<< m1 >>
rect 127 258 128 259 
<< m1 >>
rect 163 258 164 259 
<< m1 >>
rect 203 258 204 259 
<< m1 >>
rect 208 258 209 259 
<< m1 >>
rect 244 258 245 259 
<< m1 >>
rect 250 258 251 259 
<< m1 >>
rect 254 258 255 259 
<< m2 >>
rect 254 258 255 259 
<< m2c >>
rect 254 258 255 259 
<< m1 >>
rect 254 258 255 259 
<< m2 >>
rect 254 258 255 259 
<< m1 >>
rect 282 258 283 259 
<< m1 >>
rect 307 258 308 259 
<< m2 >>
rect 307 258 308 259 
<< m1 >>
rect 337 258 338 259 
<< m2 >>
rect 350 258 351 259 
<< m2 >>
rect 352 258 353 259 
<< m2 >>
rect 354 258 355 259 
<< m2 >>
rect 355 258 356 259 
<< m2 >>
rect 356 258 357 259 
<< m2 >>
rect 357 258 358 259 
<< m2 >>
rect 358 258 359 259 
<< m2 >>
rect 359 258 360 259 
<< m1 >>
rect 360 258 361 259 
<< m2 >>
rect 360 258 361 259 
<< m2c >>
rect 360 258 361 259 
<< m1 >>
rect 360 258 361 259 
<< m2 >>
rect 360 258 361 259 
<< m1 >>
rect 361 258 362 259 
<< m1 >>
rect 362 258 363 259 
<< m1 >>
rect 363 258 364 259 
<< m1 >>
rect 364 258 365 259 
<< m1 >>
rect 365 258 366 259 
<< m1 >>
rect 366 258 367 259 
<< m1 >>
rect 367 258 368 259 
<< m1 >>
rect 368 258 369 259 
<< m1 >>
rect 369 258 370 259 
<< m1 >>
rect 370 258 371 259 
<< m1 >>
rect 371 258 372 259 
<< m1 >>
rect 372 258 373 259 
<< m1 >>
rect 373 258 374 259 
<< m1 >>
rect 379 258 380 259 
<< m1 >>
rect 64 259 65 260 
<< m1 >>
rect 127 259 128 260 
<< m1 >>
rect 163 259 164 260 
<< m1 >>
rect 203 259 204 260 
<< m1 >>
rect 204 259 205 260 
<< m1 >>
rect 205 259 206 260 
<< m1 >>
rect 206 259 207 260 
<< m2 >>
rect 206 259 207 260 
<< m2c >>
rect 206 259 207 260 
<< m1 >>
rect 206 259 207 260 
<< m2 >>
rect 206 259 207 260 
<< m2 >>
rect 207 259 208 260 
<< m1 >>
rect 208 259 209 260 
<< m2 >>
rect 208 259 209 260 
<< m2 >>
rect 209 259 210 260 
<< m1 >>
rect 210 259 211 260 
<< m2 >>
rect 210 259 211 260 
<< m2c >>
rect 210 259 211 260 
<< m1 >>
rect 210 259 211 260 
<< m2 >>
rect 210 259 211 260 
<< m1 >>
rect 211 259 212 260 
<< m1 >>
rect 212 259 213 260 
<< m1 >>
rect 213 259 214 260 
<< m1 >>
rect 214 259 215 260 
<< m1 >>
rect 215 259 216 260 
<< m1 >>
rect 216 259 217 260 
<< m1 >>
rect 217 259 218 260 
<< m1 >>
rect 218 259 219 260 
<< m1 >>
rect 219 259 220 260 
<< m1 >>
rect 220 259 221 260 
<< m1 >>
rect 221 259 222 260 
<< m1 >>
rect 222 259 223 260 
<< m1 >>
rect 223 259 224 260 
<< m1 >>
rect 224 259 225 260 
<< m1 >>
rect 225 259 226 260 
<< m1 >>
rect 226 259 227 260 
<< m1 >>
rect 227 259 228 260 
<< m1 >>
rect 228 259 229 260 
<< m1 >>
rect 229 259 230 260 
<< m1 >>
rect 230 259 231 260 
<< m1 >>
rect 231 259 232 260 
<< m1 >>
rect 232 259 233 260 
<< m1 >>
rect 233 259 234 260 
<< m1 >>
rect 234 259 235 260 
<< m1 >>
rect 235 259 236 260 
<< m1 >>
rect 236 259 237 260 
<< m1 >>
rect 237 259 238 260 
<< m1 >>
rect 238 259 239 260 
<< m1 >>
rect 239 259 240 260 
<< m1 >>
rect 240 259 241 260 
<< m1 >>
rect 241 259 242 260 
<< m1 >>
rect 242 259 243 260 
<< m2 >>
rect 242 259 243 260 
<< m2c >>
rect 242 259 243 260 
<< m1 >>
rect 242 259 243 260 
<< m2 >>
rect 242 259 243 260 
<< m2 >>
rect 243 259 244 260 
<< m1 >>
rect 244 259 245 260 
<< m2 >>
rect 244 259 245 260 
<< m2 >>
rect 245 259 246 260 
<< m1 >>
rect 246 259 247 260 
<< m2 >>
rect 246 259 247 260 
<< m1 >>
rect 247 259 248 260 
<< m2 >>
rect 247 259 248 260 
<< m1 >>
rect 248 259 249 260 
<< m2 >>
rect 248 259 249 260 
<< m1 >>
rect 249 259 250 260 
<< m2 >>
rect 249 259 250 260 
<< m1 >>
rect 250 259 251 260 
<< m2 >>
rect 250 259 251 260 
<< m2 >>
rect 251 259 252 260 
<< m2 >>
rect 254 259 255 260 
<< m1 >>
rect 282 259 283 260 
<< m1 >>
rect 300 259 301 260 
<< m1 >>
rect 301 259 302 260 
<< m1 >>
rect 302 259 303 260 
<< m1 >>
rect 303 259 304 260 
<< m1 >>
rect 304 259 305 260 
<< m1 >>
rect 307 259 308 260 
<< m2 >>
rect 307 259 308 260 
<< m1 >>
rect 337 259 338 260 
<< m1 >>
rect 338 259 339 260 
<< m1 >>
rect 339 259 340 260 
<< m1 >>
rect 340 259 341 260 
<< m1 >>
rect 341 259 342 260 
<< m1 >>
rect 342 259 343 260 
<< m1 >>
rect 343 259 344 260 
<< m1 >>
rect 344 259 345 260 
<< m1 >>
rect 345 259 346 260 
<< m1 >>
rect 346 259 347 260 
<< m1 >>
rect 347 259 348 260 
<< m1 >>
rect 348 259 349 260 
<< m1 >>
rect 349 259 350 260 
<< m1 >>
rect 350 259 351 260 
<< m2 >>
rect 350 259 351 260 
<< m1 >>
rect 351 259 352 260 
<< m1 >>
rect 352 259 353 260 
<< m2 >>
rect 352 259 353 260 
<< m1 >>
rect 353 259 354 260 
<< m1 >>
rect 354 259 355 260 
<< m2 >>
rect 354 259 355 260 
<< m1 >>
rect 355 259 356 260 
<< m1 >>
rect 356 259 357 260 
<< m1 >>
rect 357 259 358 260 
<< m1 >>
rect 358 259 359 260 
<< m1 >>
rect 379 259 380 260 
<< m1 >>
rect 64 260 65 261 
<< m1 >>
rect 127 260 128 261 
<< m1 >>
rect 163 260 164 261 
<< m1 >>
rect 208 260 209 261 
<< m1 >>
rect 244 260 245 261 
<< m1 >>
rect 246 260 247 261 
<< m2 >>
rect 251 260 252 261 
<< m1 >>
rect 252 260 253 261 
<< m2 >>
rect 252 260 253 261 
<< m2c >>
rect 252 260 253 261 
<< m1 >>
rect 252 260 253 261 
<< m2 >>
rect 252 260 253 261 
<< m1 >>
rect 253 260 254 261 
<< m1 >>
rect 254 260 255 261 
<< m2 >>
rect 254 260 255 261 
<< m1 >>
rect 255 260 256 261 
<< m1 >>
rect 256 260 257 261 
<< m1 >>
rect 257 260 258 261 
<< m1 >>
rect 258 260 259 261 
<< m1 >>
rect 259 260 260 261 
<< m1 >>
rect 260 260 261 261 
<< m1 >>
rect 261 260 262 261 
<< m1 >>
rect 262 260 263 261 
<< m1 >>
rect 282 260 283 261 
<< m1 >>
rect 300 260 301 261 
<< m2 >>
rect 300 260 301 261 
<< m2c >>
rect 300 260 301 261 
<< m1 >>
rect 300 260 301 261 
<< m2 >>
rect 300 260 301 261 
<< m1 >>
rect 304 260 305 261 
<< m1 >>
rect 307 260 308 261 
<< m2 >>
rect 307 260 308 261 
<< m2 >>
rect 350 260 351 261 
<< m2 >>
rect 352 260 353 261 
<< m2 >>
rect 354 260 355 261 
<< m1 >>
rect 358 260 359 261 
<< m1 >>
rect 379 260 380 261 
<< m2 >>
rect 379 260 380 261 
<< m2c >>
rect 379 260 380 261 
<< m1 >>
rect 379 260 380 261 
<< m2 >>
rect 379 260 380 261 
<< m1 >>
rect 64 261 65 262 
<< m1 >>
rect 121 261 122 262 
<< m1 >>
rect 122 261 123 262 
<< m1 >>
rect 123 261 124 262 
<< m1 >>
rect 124 261 125 262 
<< m1 >>
rect 125 261 126 262 
<< m1 >>
rect 126 261 127 262 
<< m1 >>
rect 127 261 128 262 
<< m1 >>
rect 163 261 164 262 
<< m1 >>
rect 175 261 176 262 
<< m1 >>
rect 176 261 177 262 
<< m2 >>
rect 176 261 177 262 
<< m2c >>
rect 176 261 177 262 
<< m1 >>
rect 176 261 177 262 
<< m2 >>
rect 176 261 177 262 
<< m2 >>
rect 177 261 178 262 
<< m2 >>
rect 178 261 179 262 
<< m2 >>
rect 179 261 180 262 
<< m2 >>
rect 180 261 181 262 
<< m2 >>
rect 181 261 182 262 
<< m2 >>
rect 182 261 183 262 
<< m1 >>
rect 208 261 209 262 
<< m1 >>
rect 244 261 245 262 
<< m1 >>
rect 246 261 247 262 
<< m2 >>
rect 254 261 255 262 
<< m1 >>
rect 262 261 263 262 
<< m2 >>
rect 272 261 273 262 
<< m1 >>
rect 273 261 274 262 
<< m2 >>
rect 273 261 274 262 
<< m2c >>
rect 273 261 274 262 
<< m1 >>
rect 273 261 274 262 
<< m2 >>
rect 273 261 274 262 
<< m1 >>
rect 274 261 275 262 
<< m1 >>
rect 275 261 276 262 
<< m1 >>
rect 276 261 277 262 
<< m1 >>
rect 277 261 278 262 
<< m1 >>
rect 278 261 279 262 
<< m1 >>
rect 279 261 280 262 
<< m1 >>
rect 280 261 281 262 
<< m1 >>
rect 281 261 282 262 
<< m1 >>
rect 282 261 283 262 
<< m2 >>
rect 298 261 299 262 
<< m2 >>
rect 299 261 300 262 
<< m2 >>
rect 300 261 301 262 
<< m1 >>
rect 304 261 305 262 
<< m1 >>
rect 307 261 308 262 
<< m2 >>
rect 307 261 308 262 
<< m1 >>
rect 350 261 351 262 
<< m2 >>
rect 350 261 351 262 
<< m2c >>
rect 350 261 351 262 
<< m1 >>
rect 350 261 351 262 
<< m2 >>
rect 350 261 351 262 
<< m1 >>
rect 352 261 353 262 
<< m2 >>
rect 352 261 353 262 
<< m1 >>
rect 353 261 354 262 
<< m1 >>
rect 354 261 355 262 
<< m2 >>
rect 354 261 355 262 
<< m2c >>
rect 354 261 355 262 
<< m1 >>
rect 354 261 355 262 
<< m2 >>
rect 354 261 355 262 
<< m1 >>
rect 358 261 359 262 
<< m2 >>
rect 379 261 380 262 
<< m1 >>
rect 52 262 53 263 
<< m1 >>
rect 53 262 54 263 
<< m1 >>
rect 54 262 55 263 
<< m1 >>
rect 55 262 56 263 
<< m1 >>
rect 64 262 65 263 
<< m1 >>
rect 121 262 122 263 
<< m1 >>
rect 163 262 164 263 
<< m1 >>
rect 175 262 176 263 
<< m1 >>
rect 178 262 179 263 
<< m1 >>
rect 179 262 180 263 
<< m1 >>
rect 180 262 181 263 
<< m1 >>
rect 181 262 182 263 
<< m2 >>
rect 182 262 183 263 
<< m1 >>
rect 196 262 197 263 
<< m1 >>
rect 197 262 198 263 
<< m1 >>
rect 198 262 199 263 
<< m1 >>
rect 199 262 200 263 
<< m1 >>
rect 200 262 201 263 
<< m1 >>
rect 201 262 202 263 
<< m1 >>
rect 202 262 203 263 
<< m1 >>
rect 203 262 204 263 
<< m1 >>
rect 204 262 205 263 
<< m1 >>
rect 205 262 206 263 
<< m1 >>
rect 206 262 207 263 
<< m1 >>
rect 208 262 209 263 
<< m2 >>
rect 243 262 244 263 
<< m1 >>
rect 244 262 245 263 
<< m2 >>
rect 244 262 245 263 
<< m2 >>
rect 245 262 246 263 
<< m1 >>
rect 246 262 247 263 
<< m2 >>
rect 246 262 247 263 
<< m2c >>
rect 246 262 247 263 
<< m1 >>
rect 246 262 247 263 
<< m2 >>
rect 246 262 247 263 
<< m1 >>
rect 254 262 255 263 
<< m2 >>
rect 254 262 255 263 
<< m2c >>
rect 254 262 255 263 
<< m1 >>
rect 254 262 255 263 
<< m2 >>
rect 254 262 255 263 
<< m1 >>
rect 262 262 263 263 
<< m1 >>
rect 268 262 269 263 
<< m1 >>
rect 269 262 270 263 
<< m1 >>
rect 270 262 271 263 
<< m1 >>
rect 271 262 272 263 
<< m2 >>
rect 272 262 273 263 
<< m1 >>
rect 286 262 287 263 
<< m1 >>
rect 287 262 288 263 
<< m1 >>
rect 288 262 289 263 
<< m1 >>
rect 289 262 290 263 
<< m1 >>
rect 290 262 291 263 
<< m1 >>
rect 291 262 292 263 
<< m1 >>
rect 292 262 293 263 
<< m1 >>
rect 293 262 294 263 
<< m1 >>
rect 294 262 295 263 
<< m1 >>
rect 295 262 296 263 
<< m1 >>
rect 296 262 297 263 
<< m1 >>
rect 297 262 298 263 
<< m1 >>
rect 298 262 299 263 
<< m2 >>
rect 298 262 299 263 
<< m1 >>
rect 299 262 300 263 
<< m1 >>
rect 300 262 301 263 
<< m1 >>
rect 301 262 302 263 
<< m1 >>
rect 304 262 305 263 
<< m1 >>
rect 307 262 308 263 
<< m2 >>
rect 307 262 308 263 
<< m1 >>
rect 325 262 326 263 
<< m1 >>
rect 326 262 327 263 
<< m1 >>
rect 327 262 328 263 
<< m1 >>
rect 328 262 329 263 
<< m1 >>
rect 329 262 330 263 
<< m1 >>
rect 330 262 331 263 
<< m1 >>
rect 331 262 332 263 
<< m1 >>
rect 332 262 333 263 
<< m1 >>
rect 333 262 334 263 
<< m1 >>
rect 334 262 335 263 
<< m1 >>
rect 335 262 336 263 
<< m1 >>
rect 336 262 337 263 
<< m1 >>
rect 337 262 338 263 
<< m1 >>
rect 350 262 351 263 
<< m1 >>
rect 352 262 353 263 
<< m2 >>
rect 352 262 353 263 
<< m1 >>
rect 358 262 359 263 
<< m1 >>
rect 376 262 377 263 
<< m1 >>
rect 377 262 378 263 
<< m1 >>
rect 378 262 379 263 
<< m1 >>
rect 379 262 380 263 
<< m2 >>
rect 379 262 380 263 
<< m1 >>
rect 380 262 381 263 
<< m1 >>
rect 381 262 382 263 
<< m1 >>
rect 382 262 383 263 
<< m1 >>
rect 383 262 384 263 
<< m1 >>
rect 384 262 385 263 
<< m1 >>
rect 385 262 386 263 
<< m1 >>
rect 386 262 387 263 
<< m1 >>
rect 387 262 388 263 
<< m1 >>
rect 388 262 389 263 
<< m1 >>
rect 52 263 53 264 
<< m1 >>
rect 55 263 56 264 
<< m1 >>
rect 64 263 65 264 
<< m1 >>
rect 121 263 122 264 
<< m1 >>
rect 163 263 164 264 
<< m1 >>
rect 175 263 176 264 
<< m1 >>
rect 178 263 179 264 
<< m1 >>
rect 181 263 182 264 
<< m2 >>
rect 182 263 183 264 
<< m1 >>
rect 196 263 197 264 
<< m1 >>
rect 206 263 207 264 
<< m1 >>
rect 208 263 209 264 
<< m2 >>
rect 243 263 244 264 
<< m1 >>
rect 244 263 245 264 
<< m1 >>
rect 254 263 255 264 
<< m1 >>
rect 262 263 263 264 
<< m1 >>
rect 268 263 269 264 
<< m1 >>
rect 271 263 272 264 
<< m2 >>
rect 272 263 273 264 
<< m1 >>
rect 286 263 287 264 
<< m2 >>
rect 298 263 299 264 
<< m1 >>
rect 301 263 302 264 
<< m1 >>
rect 304 263 305 264 
<< m1 >>
rect 307 263 308 264 
<< m2 >>
rect 307 263 308 264 
<< m1 >>
rect 325 263 326 264 
<< m1 >>
rect 337 263 338 264 
<< m1 >>
rect 350 263 351 264 
<< m1 >>
rect 352 263 353 264 
<< m2 >>
rect 352 263 353 264 
<< m1 >>
rect 358 263 359 264 
<< m1 >>
rect 376 263 377 264 
<< m2 >>
rect 379 263 380 264 
<< m1 >>
rect 388 263 389 264 
<< pdiffusion >>
rect 12 264 13 265 
<< pdiffusion >>
rect 13 264 14 265 
<< pdiffusion >>
rect 14 264 15 265 
<< pdiffusion >>
rect 15 264 16 265 
<< pdiffusion >>
rect 16 264 17 265 
<< pdiffusion >>
rect 17 264 18 265 
<< pdiffusion >>
rect 48 264 49 265 
<< pdiffusion >>
rect 49 264 50 265 
<< pdiffusion >>
rect 50 264 51 265 
<< pdiffusion >>
rect 51 264 52 265 
<< m1 >>
rect 52 264 53 265 
<< pdiffusion >>
rect 52 264 53 265 
<< pdiffusion >>
rect 53 264 54 265 
<< m1 >>
rect 55 264 56 265 
<< m1 >>
rect 64 264 65 265 
<< pdiffusion >>
rect 66 264 67 265 
<< pdiffusion >>
rect 67 264 68 265 
<< pdiffusion >>
rect 68 264 69 265 
<< pdiffusion >>
rect 69 264 70 265 
<< pdiffusion >>
rect 70 264 71 265 
<< pdiffusion >>
rect 71 264 72 265 
<< pdiffusion >>
rect 84 264 85 265 
<< pdiffusion >>
rect 85 264 86 265 
<< pdiffusion >>
rect 86 264 87 265 
<< pdiffusion >>
rect 87 264 88 265 
<< pdiffusion >>
rect 88 264 89 265 
<< pdiffusion >>
rect 89 264 90 265 
<< pdiffusion >>
rect 102 264 103 265 
<< pdiffusion >>
rect 103 264 104 265 
<< pdiffusion >>
rect 104 264 105 265 
<< pdiffusion >>
rect 105 264 106 265 
<< pdiffusion >>
rect 106 264 107 265 
<< pdiffusion >>
rect 107 264 108 265 
<< pdiffusion >>
rect 120 264 121 265 
<< m1 >>
rect 121 264 122 265 
<< pdiffusion >>
rect 121 264 122 265 
<< pdiffusion >>
rect 122 264 123 265 
<< pdiffusion >>
rect 123 264 124 265 
<< pdiffusion >>
rect 124 264 125 265 
<< pdiffusion >>
rect 125 264 126 265 
<< pdiffusion >>
rect 156 264 157 265 
<< pdiffusion >>
rect 157 264 158 265 
<< pdiffusion >>
rect 158 264 159 265 
<< pdiffusion >>
rect 159 264 160 265 
<< pdiffusion >>
rect 160 264 161 265 
<< pdiffusion >>
rect 161 264 162 265 
<< m1 >>
rect 163 264 164 265 
<< pdiffusion >>
rect 174 264 175 265 
<< m1 >>
rect 175 264 176 265 
<< pdiffusion >>
rect 175 264 176 265 
<< pdiffusion >>
rect 176 264 177 265 
<< pdiffusion >>
rect 177 264 178 265 
<< m1 >>
rect 178 264 179 265 
<< pdiffusion >>
rect 178 264 179 265 
<< pdiffusion >>
rect 179 264 180 265 
<< m1 >>
rect 181 264 182 265 
<< m2 >>
rect 182 264 183 265 
<< pdiffusion >>
rect 192 264 193 265 
<< pdiffusion >>
rect 193 264 194 265 
<< pdiffusion >>
rect 194 264 195 265 
<< pdiffusion >>
rect 195 264 196 265 
<< m1 >>
rect 196 264 197 265 
<< pdiffusion >>
rect 196 264 197 265 
<< pdiffusion >>
rect 197 264 198 265 
<< m1 >>
rect 206 264 207 265 
<< m1 >>
rect 208 264 209 265 
<< pdiffusion >>
rect 210 264 211 265 
<< pdiffusion >>
rect 211 264 212 265 
<< pdiffusion >>
rect 212 264 213 265 
<< pdiffusion >>
rect 213 264 214 265 
<< pdiffusion >>
rect 214 264 215 265 
<< pdiffusion >>
rect 215 264 216 265 
<< pdiffusion >>
rect 228 264 229 265 
<< pdiffusion >>
rect 229 264 230 265 
<< pdiffusion >>
rect 230 264 231 265 
<< pdiffusion >>
rect 231 264 232 265 
<< pdiffusion >>
rect 232 264 233 265 
<< pdiffusion >>
rect 233 264 234 265 
<< m2 >>
rect 243 264 244 265 
<< m1 >>
rect 244 264 245 265 
<< pdiffusion >>
rect 246 264 247 265 
<< pdiffusion >>
rect 247 264 248 265 
<< pdiffusion >>
rect 248 264 249 265 
<< pdiffusion >>
rect 249 264 250 265 
<< pdiffusion >>
rect 250 264 251 265 
<< pdiffusion >>
rect 251 264 252 265 
<< m1 >>
rect 254 264 255 265 
<< m1 >>
rect 262 264 263 265 
<< pdiffusion >>
rect 264 264 265 265 
<< pdiffusion >>
rect 265 264 266 265 
<< pdiffusion >>
rect 266 264 267 265 
<< pdiffusion >>
rect 267 264 268 265 
<< m1 >>
rect 268 264 269 265 
<< pdiffusion >>
rect 268 264 269 265 
<< pdiffusion >>
rect 269 264 270 265 
<< m1 >>
rect 271 264 272 265 
<< m2 >>
rect 272 264 273 265 
<< pdiffusion >>
rect 282 264 283 265 
<< pdiffusion >>
rect 283 264 284 265 
<< pdiffusion >>
rect 284 264 285 265 
<< pdiffusion >>
rect 285 264 286 265 
<< m1 >>
rect 286 264 287 265 
<< pdiffusion >>
rect 286 264 287 265 
<< pdiffusion >>
rect 287 264 288 265 
<< m1 >>
rect 298 264 299 265 
<< m2 >>
rect 298 264 299 265 
<< m2c >>
rect 298 264 299 265 
<< m1 >>
rect 298 264 299 265 
<< m2 >>
rect 298 264 299 265 
<< pdiffusion >>
rect 300 264 301 265 
<< m1 >>
rect 301 264 302 265 
<< pdiffusion >>
rect 301 264 302 265 
<< pdiffusion >>
rect 302 264 303 265 
<< pdiffusion >>
rect 303 264 304 265 
<< m1 >>
rect 304 264 305 265 
<< pdiffusion >>
rect 304 264 305 265 
<< pdiffusion >>
rect 305 264 306 265 
<< m1 >>
rect 307 264 308 265 
<< m2 >>
rect 307 264 308 265 
<< pdiffusion >>
rect 318 264 319 265 
<< pdiffusion >>
rect 319 264 320 265 
<< pdiffusion >>
rect 320 264 321 265 
<< pdiffusion >>
rect 321 264 322 265 
<< pdiffusion >>
rect 322 264 323 265 
<< pdiffusion >>
rect 323 264 324 265 
<< m1 >>
rect 325 264 326 265 
<< pdiffusion >>
rect 336 264 337 265 
<< m1 >>
rect 337 264 338 265 
<< pdiffusion >>
rect 337 264 338 265 
<< pdiffusion >>
rect 338 264 339 265 
<< pdiffusion >>
rect 339 264 340 265 
<< pdiffusion >>
rect 340 264 341 265 
<< pdiffusion >>
rect 341 264 342 265 
<< m1 >>
rect 350 264 351 265 
<< m1 >>
rect 352 264 353 265 
<< m2 >>
rect 352 264 353 265 
<< pdiffusion >>
rect 354 264 355 265 
<< pdiffusion >>
rect 355 264 356 265 
<< pdiffusion >>
rect 356 264 357 265 
<< pdiffusion >>
rect 357 264 358 265 
<< m1 >>
rect 358 264 359 265 
<< pdiffusion >>
rect 358 264 359 265 
<< pdiffusion >>
rect 359 264 360 265 
<< pdiffusion >>
rect 372 264 373 265 
<< pdiffusion >>
rect 373 264 374 265 
<< pdiffusion >>
rect 374 264 375 265 
<< pdiffusion >>
rect 375 264 376 265 
<< m1 >>
rect 376 264 377 265 
<< pdiffusion >>
rect 376 264 377 265 
<< pdiffusion >>
rect 377 264 378 265 
<< m1 >>
rect 379 264 380 265 
<< m2 >>
rect 379 264 380 265 
<< m2c >>
rect 379 264 380 265 
<< m1 >>
rect 379 264 380 265 
<< m2 >>
rect 379 264 380 265 
<< m1 >>
rect 388 264 389 265 
<< pdiffusion >>
rect 390 264 391 265 
<< pdiffusion >>
rect 391 264 392 265 
<< pdiffusion >>
rect 392 264 393 265 
<< pdiffusion >>
rect 393 264 394 265 
<< pdiffusion >>
rect 394 264 395 265 
<< pdiffusion >>
rect 395 264 396 265 
<< pdiffusion >>
rect 408 264 409 265 
<< pdiffusion >>
rect 409 264 410 265 
<< pdiffusion >>
rect 410 264 411 265 
<< pdiffusion >>
rect 411 264 412 265 
<< pdiffusion >>
rect 412 264 413 265 
<< pdiffusion >>
rect 413 264 414 265 
<< pdiffusion >>
rect 426 264 427 265 
<< pdiffusion >>
rect 427 264 428 265 
<< pdiffusion >>
rect 428 264 429 265 
<< pdiffusion >>
rect 429 264 430 265 
<< pdiffusion >>
rect 430 264 431 265 
<< pdiffusion >>
rect 431 264 432 265 
<< pdiffusion >>
rect 444 264 445 265 
<< pdiffusion >>
rect 445 264 446 265 
<< pdiffusion >>
rect 446 264 447 265 
<< pdiffusion >>
rect 447 264 448 265 
<< pdiffusion >>
rect 448 264 449 265 
<< pdiffusion >>
rect 449 264 450 265 
<< pdiffusion >>
rect 12 265 13 266 
<< pdiffusion >>
rect 13 265 14 266 
<< pdiffusion >>
rect 14 265 15 266 
<< pdiffusion >>
rect 15 265 16 266 
<< pdiffusion >>
rect 16 265 17 266 
<< pdiffusion >>
rect 17 265 18 266 
<< pdiffusion >>
rect 48 265 49 266 
<< pdiffusion >>
rect 49 265 50 266 
<< pdiffusion >>
rect 50 265 51 266 
<< pdiffusion >>
rect 51 265 52 266 
<< pdiffusion >>
rect 52 265 53 266 
<< pdiffusion >>
rect 53 265 54 266 
<< m1 >>
rect 55 265 56 266 
<< m1 >>
rect 64 265 65 266 
<< pdiffusion >>
rect 66 265 67 266 
<< pdiffusion >>
rect 67 265 68 266 
<< pdiffusion >>
rect 68 265 69 266 
<< pdiffusion >>
rect 69 265 70 266 
<< pdiffusion >>
rect 70 265 71 266 
<< pdiffusion >>
rect 71 265 72 266 
<< pdiffusion >>
rect 84 265 85 266 
<< pdiffusion >>
rect 85 265 86 266 
<< pdiffusion >>
rect 86 265 87 266 
<< pdiffusion >>
rect 87 265 88 266 
<< pdiffusion >>
rect 88 265 89 266 
<< pdiffusion >>
rect 89 265 90 266 
<< pdiffusion >>
rect 102 265 103 266 
<< pdiffusion >>
rect 103 265 104 266 
<< pdiffusion >>
rect 104 265 105 266 
<< pdiffusion >>
rect 105 265 106 266 
<< pdiffusion >>
rect 106 265 107 266 
<< pdiffusion >>
rect 107 265 108 266 
<< pdiffusion >>
rect 120 265 121 266 
<< pdiffusion >>
rect 121 265 122 266 
<< pdiffusion >>
rect 122 265 123 266 
<< pdiffusion >>
rect 123 265 124 266 
<< pdiffusion >>
rect 124 265 125 266 
<< pdiffusion >>
rect 125 265 126 266 
<< pdiffusion >>
rect 156 265 157 266 
<< pdiffusion >>
rect 157 265 158 266 
<< pdiffusion >>
rect 158 265 159 266 
<< pdiffusion >>
rect 159 265 160 266 
<< pdiffusion >>
rect 160 265 161 266 
<< pdiffusion >>
rect 161 265 162 266 
<< m1 >>
rect 163 265 164 266 
<< pdiffusion >>
rect 174 265 175 266 
<< pdiffusion >>
rect 175 265 176 266 
<< pdiffusion >>
rect 176 265 177 266 
<< pdiffusion >>
rect 177 265 178 266 
<< pdiffusion >>
rect 178 265 179 266 
<< pdiffusion >>
rect 179 265 180 266 
<< m1 >>
rect 181 265 182 266 
<< m2 >>
rect 182 265 183 266 
<< pdiffusion >>
rect 192 265 193 266 
<< pdiffusion >>
rect 193 265 194 266 
<< pdiffusion >>
rect 194 265 195 266 
<< pdiffusion >>
rect 195 265 196 266 
<< pdiffusion >>
rect 196 265 197 266 
<< pdiffusion >>
rect 197 265 198 266 
<< m1 >>
rect 206 265 207 266 
<< m1 >>
rect 208 265 209 266 
<< pdiffusion >>
rect 210 265 211 266 
<< pdiffusion >>
rect 211 265 212 266 
<< pdiffusion >>
rect 212 265 213 266 
<< pdiffusion >>
rect 213 265 214 266 
<< pdiffusion >>
rect 214 265 215 266 
<< pdiffusion >>
rect 215 265 216 266 
<< pdiffusion >>
rect 228 265 229 266 
<< pdiffusion >>
rect 229 265 230 266 
<< pdiffusion >>
rect 230 265 231 266 
<< pdiffusion >>
rect 231 265 232 266 
<< pdiffusion >>
rect 232 265 233 266 
<< pdiffusion >>
rect 233 265 234 266 
<< m2 >>
rect 243 265 244 266 
<< m1 >>
rect 244 265 245 266 
<< pdiffusion >>
rect 246 265 247 266 
<< pdiffusion >>
rect 247 265 248 266 
<< pdiffusion >>
rect 248 265 249 266 
<< pdiffusion >>
rect 249 265 250 266 
<< pdiffusion >>
rect 250 265 251 266 
<< pdiffusion >>
rect 251 265 252 266 
<< m1 >>
rect 254 265 255 266 
<< m1 >>
rect 262 265 263 266 
<< pdiffusion >>
rect 264 265 265 266 
<< pdiffusion >>
rect 265 265 266 266 
<< pdiffusion >>
rect 266 265 267 266 
<< pdiffusion >>
rect 267 265 268 266 
<< pdiffusion >>
rect 268 265 269 266 
<< pdiffusion >>
rect 269 265 270 266 
<< m1 >>
rect 271 265 272 266 
<< m2 >>
rect 272 265 273 266 
<< pdiffusion >>
rect 282 265 283 266 
<< pdiffusion >>
rect 283 265 284 266 
<< pdiffusion >>
rect 284 265 285 266 
<< pdiffusion >>
rect 285 265 286 266 
<< pdiffusion >>
rect 286 265 287 266 
<< pdiffusion >>
rect 287 265 288 266 
<< m1 >>
rect 298 265 299 266 
<< pdiffusion >>
rect 300 265 301 266 
<< pdiffusion >>
rect 301 265 302 266 
<< pdiffusion >>
rect 302 265 303 266 
<< pdiffusion >>
rect 303 265 304 266 
<< pdiffusion >>
rect 304 265 305 266 
<< pdiffusion >>
rect 305 265 306 266 
<< m1 >>
rect 307 265 308 266 
<< m2 >>
rect 307 265 308 266 
<< pdiffusion >>
rect 318 265 319 266 
<< pdiffusion >>
rect 319 265 320 266 
<< pdiffusion >>
rect 320 265 321 266 
<< pdiffusion >>
rect 321 265 322 266 
<< pdiffusion >>
rect 322 265 323 266 
<< pdiffusion >>
rect 323 265 324 266 
<< m1 >>
rect 325 265 326 266 
<< pdiffusion >>
rect 336 265 337 266 
<< pdiffusion >>
rect 337 265 338 266 
<< pdiffusion >>
rect 338 265 339 266 
<< pdiffusion >>
rect 339 265 340 266 
<< pdiffusion >>
rect 340 265 341 266 
<< pdiffusion >>
rect 341 265 342 266 
<< m1 >>
rect 350 265 351 266 
<< m1 >>
rect 352 265 353 266 
<< m2 >>
rect 352 265 353 266 
<< pdiffusion >>
rect 354 265 355 266 
<< pdiffusion >>
rect 355 265 356 266 
<< pdiffusion >>
rect 356 265 357 266 
<< pdiffusion >>
rect 357 265 358 266 
<< pdiffusion >>
rect 358 265 359 266 
<< pdiffusion >>
rect 359 265 360 266 
<< pdiffusion >>
rect 372 265 373 266 
<< pdiffusion >>
rect 373 265 374 266 
<< pdiffusion >>
rect 374 265 375 266 
<< pdiffusion >>
rect 375 265 376 266 
<< pdiffusion >>
rect 376 265 377 266 
<< pdiffusion >>
rect 377 265 378 266 
<< m1 >>
rect 379 265 380 266 
<< m1 >>
rect 388 265 389 266 
<< pdiffusion >>
rect 390 265 391 266 
<< pdiffusion >>
rect 391 265 392 266 
<< pdiffusion >>
rect 392 265 393 266 
<< pdiffusion >>
rect 393 265 394 266 
<< pdiffusion >>
rect 394 265 395 266 
<< pdiffusion >>
rect 395 265 396 266 
<< pdiffusion >>
rect 408 265 409 266 
<< pdiffusion >>
rect 409 265 410 266 
<< pdiffusion >>
rect 410 265 411 266 
<< pdiffusion >>
rect 411 265 412 266 
<< pdiffusion >>
rect 412 265 413 266 
<< pdiffusion >>
rect 413 265 414 266 
<< pdiffusion >>
rect 426 265 427 266 
<< pdiffusion >>
rect 427 265 428 266 
<< pdiffusion >>
rect 428 265 429 266 
<< pdiffusion >>
rect 429 265 430 266 
<< pdiffusion >>
rect 430 265 431 266 
<< pdiffusion >>
rect 431 265 432 266 
<< pdiffusion >>
rect 444 265 445 266 
<< pdiffusion >>
rect 445 265 446 266 
<< pdiffusion >>
rect 446 265 447 266 
<< pdiffusion >>
rect 447 265 448 266 
<< pdiffusion >>
rect 448 265 449 266 
<< pdiffusion >>
rect 449 265 450 266 
<< pdiffusion >>
rect 12 266 13 267 
<< pdiffusion >>
rect 13 266 14 267 
<< pdiffusion >>
rect 14 266 15 267 
<< pdiffusion >>
rect 15 266 16 267 
<< pdiffusion >>
rect 16 266 17 267 
<< pdiffusion >>
rect 17 266 18 267 
<< pdiffusion >>
rect 48 266 49 267 
<< pdiffusion >>
rect 49 266 50 267 
<< pdiffusion >>
rect 50 266 51 267 
<< pdiffusion >>
rect 51 266 52 267 
<< pdiffusion >>
rect 52 266 53 267 
<< pdiffusion >>
rect 53 266 54 267 
<< m1 >>
rect 55 266 56 267 
<< m1 >>
rect 64 266 65 267 
<< pdiffusion >>
rect 66 266 67 267 
<< pdiffusion >>
rect 67 266 68 267 
<< pdiffusion >>
rect 68 266 69 267 
<< pdiffusion >>
rect 69 266 70 267 
<< pdiffusion >>
rect 70 266 71 267 
<< pdiffusion >>
rect 71 266 72 267 
<< pdiffusion >>
rect 84 266 85 267 
<< pdiffusion >>
rect 85 266 86 267 
<< pdiffusion >>
rect 86 266 87 267 
<< pdiffusion >>
rect 87 266 88 267 
<< pdiffusion >>
rect 88 266 89 267 
<< pdiffusion >>
rect 89 266 90 267 
<< pdiffusion >>
rect 102 266 103 267 
<< pdiffusion >>
rect 103 266 104 267 
<< pdiffusion >>
rect 104 266 105 267 
<< pdiffusion >>
rect 105 266 106 267 
<< pdiffusion >>
rect 106 266 107 267 
<< pdiffusion >>
rect 107 266 108 267 
<< pdiffusion >>
rect 120 266 121 267 
<< pdiffusion >>
rect 121 266 122 267 
<< pdiffusion >>
rect 122 266 123 267 
<< pdiffusion >>
rect 123 266 124 267 
<< pdiffusion >>
rect 124 266 125 267 
<< pdiffusion >>
rect 125 266 126 267 
<< pdiffusion >>
rect 156 266 157 267 
<< pdiffusion >>
rect 157 266 158 267 
<< pdiffusion >>
rect 158 266 159 267 
<< pdiffusion >>
rect 159 266 160 267 
<< pdiffusion >>
rect 160 266 161 267 
<< pdiffusion >>
rect 161 266 162 267 
<< m1 >>
rect 163 266 164 267 
<< pdiffusion >>
rect 174 266 175 267 
<< pdiffusion >>
rect 175 266 176 267 
<< pdiffusion >>
rect 176 266 177 267 
<< pdiffusion >>
rect 177 266 178 267 
<< pdiffusion >>
rect 178 266 179 267 
<< pdiffusion >>
rect 179 266 180 267 
<< m1 >>
rect 181 266 182 267 
<< m2 >>
rect 182 266 183 267 
<< pdiffusion >>
rect 192 266 193 267 
<< pdiffusion >>
rect 193 266 194 267 
<< pdiffusion >>
rect 194 266 195 267 
<< pdiffusion >>
rect 195 266 196 267 
<< pdiffusion >>
rect 196 266 197 267 
<< pdiffusion >>
rect 197 266 198 267 
<< m1 >>
rect 206 266 207 267 
<< m1 >>
rect 208 266 209 267 
<< pdiffusion >>
rect 210 266 211 267 
<< pdiffusion >>
rect 211 266 212 267 
<< pdiffusion >>
rect 212 266 213 267 
<< pdiffusion >>
rect 213 266 214 267 
<< pdiffusion >>
rect 214 266 215 267 
<< pdiffusion >>
rect 215 266 216 267 
<< pdiffusion >>
rect 228 266 229 267 
<< pdiffusion >>
rect 229 266 230 267 
<< pdiffusion >>
rect 230 266 231 267 
<< pdiffusion >>
rect 231 266 232 267 
<< pdiffusion >>
rect 232 266 233 267 
<< pdiffusion >>
rect 233 266 234 267 
<< m2 >>
rect 243 266 244 267 
<< m1 >>
rect 244 266 245 267 
<< pdiffusion >>
rect 246 266 247 267 
<< pdiffusion >>
rect 247 266 248 267 
<< pdiffusion >>
rect 248 266 249 267 
<< pdiffusion >>
rect 249 266 250 267 
<< pdiffusion >>
rect 250 266 251 267 
<< pdiffusion >>
rect 251 266 252 267 
<< m1 >>
rect 254 266 255 267 
<< m1 >>
rect 262 266 263 267 
<< pdiffusion >>
rect 264 266 265 267 
<< pdiffusion >>
rect 265 266 266 267 
<< pdiffusion >>
rect 266 266 267 267 
<< pdiffusion >>
rect 267 266 268 267 
<< pdiffusion >>
rect 268 266 269 267 
<< pdiffusion >>
rect 269 266 270 267 
<< m1 >>
rect 271 266 272 267 
<< m2 >>
rect 272 266 273 267 
<< pdiffusion >>
rect 282 266 283 267 
<< pdiffusion >>
rect 283 266 284 267 
<< pdiffusion >>
rect 284 266 285 267 
<< pdiffusion >>
rect 285 266 286 267 
<< pdiffusion >>
rect 286 266 287 267 
<< pdiffusion >>
rect 287 266 288 267 
<< m1 >>
rect 298 266 299 267 
<< pdiffusion >>
rect 300 266 301 267 
<< pdiffusion >>
rect 301 266 302 267 
<< pdiffusion >>
rect 302 266 303 267 
<< pdiffusion >>
rect 303 266 304 267 
<< pdiffusion >>
rect 304 266 305 267 
<< pdiffusion >>
rect 305 266 306 267 
<< m1 >>
rect 307 266 308 267 
<< m2 >>
rect 307 266 308 267 
<< pdiffusion >>
rect 318 266 319 267 
<< pdiffusion >>
rect 319 266 320 267 
<< pdiffusion >>
rect 320 266 321 267 
<< pdiffusion >>
rect 321 266 322 267 
<< pdiffusion >>
rect 322 266 323 267 
<< pdiffusion >>
rect 323 266 324 267 
<< m1 >>
rect 325 266 326 267 
<< pdiffusion >>
rect 336 266 337 267 
<< pdiffusion >>
rect 337 266 338 267 
<< pdiffusion >>
rect 338 266 339 267 
<< pdiffusion >>
rect 339 266 340 267 
<< pdiffusion >>
rect 340 266 341 267 
<< pdiffusion >>
rect 341 266 342 267 
<< m1 >>
rect 350 266 351 267 
<< m1 >>
rect 352 266 353 267 
<< m2 >>
rect 352 266 353 267 
<< pdiffusion >>
rect 354 266 355 267 
<< pdiffusion >>
rect 355 266 356 267 
<< pdiffusion >>
rect 356 266 357 267 
<< pdiffusion >>
rect 357 266 358 267 
<< pdiffusion >>
rect 358 266 359 267 
<< pdiffusion >>
rect 359 266 360 267 
<< pdiffusion >>
rect 372 266 373 267 
<< pdiffusion >>
rect 373 266 374 267 
<< pdiffusion >>
rect 374 266 375 267 
<< pdiffusion >>
rect 375 266 376 267 
<< pdiffusion >>
rect 376 266 377 267 
<< pdiffusion >>
rect 377 266 378 267 
<< m1 >>
rect 379 266 380 267 
<< m1 >>
rect 388 266 389 267 
<< pdiffusion >>
rect 390 266 391 267 
<< pdiffusion >>
rect 391 266 392 267 
<< pdiffusion >>
rect 392 266 393 267 
<< pdiffusion >>
rect 393 266 394 267 
<< pdiffusion >>
rect 394 266 395 267 
<< pdiffusion >>
rect 395 266 396 267 
<< pdiffusion >>
rect 408 266 409 267 
<< pdiffusion >>
rect 409 266 410 267 
<< pdiffusion >>
rect 410 266 411 267 
<< pdiffusion >>
rect 411 266 412 267 
<< pdiffusion >>
rect 412 266 413 267 
<< pdiffusion >>
rect 413 266 414 267 
<< pdiffusion >>
rect 426 266 427 267 
<< pdiffusion >>
rect 427 266 428 267 
<< pdiffusion >>
rect 428 266 429 267 
<< pdiffusion >>
rect 429 266 430 267 
<< pdiffusion >>
rect 430 266 431 267 
<< pdiffusion >>
rect 431 266 432 267 
<< pdiffusion >>
rect 444 266 445 267 
<< pdiffusion >>
rect 445 266 446 267 
<< pdiffusion >>
rect 446 266 447 267 
<< pdiffusion >>
rect 447 266 448 267 
<< pdiffusion >>
rect 448 266 449 267 
<< pdiffusion >>
rect 449 266 450 267 
<< pdiffusion >>
rect 12 267 13 268 
<< pdiffusion >>
rect 13 267 14 268 
<< pdiffusion >>
rect 14 267 15 268 
<< pdiffusion >>
rect 15 267 16 268 
<< pdiffusion >>
rect 16 267 17 268 
<< pdiffusion >>
rect 17 267 18 268 
<< pdiffusion >>
rect 48 267 49 268 
<< pdiffusion >>
rect 49 267 50 268 
<< pdiffusion >>
rect 50 267 51 268 
<< pdiffusion >>
rect 51 267 52 268 
<< pdiffusion >>
rect 52 267 53 268 
<< pdiffusion >>
rect 53 267 54 268 
<< m1 >>
rect 55 267 56 268 
<< m1 >>
rect 64 267 65 268 
<< pdiffusion >>
rect 66 267 67 268 
<< pdiffusion >>
rect 67 267 68 268 
<< pdiffusion >>
rect 68 267 69 268 
<< pdiffusion >>
rect 69 267 70 268 
<< pdiffusion >>
rect 70 267 71 268 
<< pdiffusion >>
rect 71 267 72 268 
<< pdiffusion >>
rect 84 267 85 268 
<< pdiffusion >>
rect 85 267 86 268 
<< pdiffusion >>
rect 86 267 87 268 
<< pdiffusion >>
rect 87 267 88 268 
<< pdiffusion >>
rect 88 267 89 268 
<< pdiffusion >>
rect 89 267 90 268 
<< pdiffusion >>
rect 102 267 103 268 
<< pdiffusion >>
rect 103 267 104 268 
<< pdiffusion >>
rect 104 267 105 268 
<< pdiffusion >>
rect 105 267 106 268 
<< pdiffusion >>
rect 106 267 107 268 
<< pdiffusion >>
rect 107 267 108 268 
<< pdiffusion >>
rect 120 267 121 268 
<< pdiffusion >>
rect 121 267 122 268 
<< pdiffusion >>
rect 122 267 123 268 
<< pdiffusion >>
rect 123 267 124 268 
<< pdiffusion >>
rect 124 267 125 268 
<< pdiffusion >>
rect 125 267 126 268 
<< pdiffusion >>
rect 156 267 157 268 
<< pdiffusion >>
rect 157 267 158 268 
<< pdiffusion >>
rect 158 267 159 268 
<< pdiffusion >>
rect 159 267 160 268 
<< pdiffusion >>
rect 160 267 161 268 
<< pdiffusion >>
rect 161 267 162 268 
<< m1 >>
rect 163 267 164 268 
<< pdiffusion >>
rect 174 267 175 268 
<< pdiffusion >>
rect 175 267 176 268 
<< pdiffusion >>
rect 176 267 177 268 
<< pdiffusion >>
rect 177 267 178 268 
<< pdiffusion >>
rect 178 267 179 268 
<< pdiffusion >>
rect 179 267 180 268 
<< m1 >>
rect 181 267 182 268 
<< m2 >>
rect 182 267 183 268 
<< pdiffusion >>
rect 192 267 193 268 
<< pdiffusion >>
rect 193 267 194 268 
<< pdiffusion >>
rect 194 267 195 268 
<< pdiffusion >>
rect 195 267 196 268 
<< pdiffusion >>
rect 196 267 197 268 
<< pdiffusion >>
rect 197 267 198 268 
<< m1 >>
rect 206 267 207 268 
<< m1 >>
rect 208 267 209 268 
<< pdiffusion >>
rect 210 267 211 268 
<< pdiffusion >>
rect 211 267 212 268 
<< pdiffusion >>
rect 212 267 213 268 
<< pdiffusion >>
rect 213 267 214 268 
<< pdiffusion >>
rect 214 267 215 268 
<< pdiffusion >>
rect 215 267 216 268 
<< pdiffusion >>
rect 228 267 229 268 
<< pdiffusion >>
rect 229 267 230 268 
<< pdiffusion >>
rect 230 267 231 268 
<< pdiffusion >>
rect 231 267 232 268 
<< pdiffusion >>
rect 232 267 233 268 
<< pdiffusion >>
rect 233 267 234 268 
<< m2 >>
rect 243 267 244 268 
<< m1 >>
rect 244 267 245 268 
<< pdiffusion >>
rect 246 267 247 268 
<< pdiffusion >>
rect 247 267 248 268 
<< pdiffusion >>
rect 248 267 249 268 
<< pdiffusion >>
rect 249 267 250 268 
<< pdiffusion >>
rect 250 267 251 268 
<< pdiffusion >>
rect 251 267 252 268 
<< m1 >>
rect 254 267 255 268 
<< m1 >>
rect 262 267 263 268 
<< pdiffusion >>
rect 264 267 265 268 
<< pdiffusion >>
rect 265 267 266 268 
<< pdiffusion >>
rect 266 267 267 268 
<< pdiffusion >>
rect 267 267 268 268 
<< pdiffusion >>
rect 268 267 269 268 
<< pdiffusion >>
rect 269 267 270 268 
<< m1 >>
rect 271 267 272 268 
<< m2 >>
rect 272 267 273 268 
<< pdiffusion >>
rect 282 267 283 268 
<< pdiffusion >>
rect 283 267 284 268 
<< pdiffusion >>
rect 284 267 285 268 
<< pdiffusion >>
rect 285 267 286 268 
<< pdiffusion >>
rect 286 267 287 268 
<< pdiffusion >>
rect 287 267 288 268 
<< m1 >>
rect 298 267 299 268 
<< pdiffusion >>
rect 300 267 301 268 
<< pdiffusion >>
rect 301 267 302 268 
<< pdiffusion >>
rect 302 267 303 268 
<< pdiffusion >>
rect 303 267 304 268 
<< pdiffusion >>
rect 304 267 305 268 
<< pdiffusion >>
rect 305 267 306 268 
<< m1 >>
rect 307 267 308 268 
<< m2 >>
rect 307 267 308 268 
<< pdiffusion >>
rect 318 267 319 268 
<< pdiffusion >>
rect 319 267 320 268 
<< pdiffusion >>
rect 320 267 321 268 
<< pdiffusion >>
rect 321 267 322 268 
<< pdiffusion >>
rect 322 267 323 268 
<< pdiffusion >>
rect 323 267 324 268 
<< m1 >>
rect 325 267 326 268 
<< pdiffusion >>
rect 336 267 337 268 
<< pdiffusion >>
rect 337 267 338 268 
<< pdiffusion >>
rect 338 267 339 268 
<< pdiffusion >>
rect 339 267 340 268 
<< pdiffusion >>
rect 340 267 341 268 
<< pdiffusion >>
rect 341 267 342 268 
<< m1 >>
rect 350 267 351 268 
<< m1 >>
rect 352 267 353 268 
<< m2 >>
rect 352 267 353 268 
<< pdiffusion >>
rect 354 267 355 268 
<< pdiffusion >>
rect 355 267 356 268 
<< pdiffusion >>
rect 356 267 357 268 
<< pdiffusion >>
rect 357 267 358 268 
<< pdiffusion >>
rect 358 267 359 268 
<< pdiffusion >>
rect 359 267 360 268 
<< pdiffusion >>
rect 372 267 373 268 
<< pdiffusion >>
rect 373 267 374 268 
<< pdiffusion >>
rect 374 267 375 268 
<< pdiffusion >>
rect 375 267 376 268 
<< pdiffusion >>
rect 376 267 377 268 
<< pdiffusion >>
rect 377 267 378 268 
<< m1 >>
rect 379 267 380 268 
<< m1 >>
rect 388 267 389 268 
<< pdiffusion >>
rect 390 267 391 268 
<< pdiffusion >>
rect 391 267 392 268 
<< pdiffusion >>
rect 392 267 393 268 
<< pdiffusion >>
rect 393 267 394 268 
<< pdiffusion >>
rect 394 267 395 268 
<< pdiffusion >>
rect 395 267 396 268 
<< pdiffusion >>
rect 408 267 409 268 
<< pdiffusion >>
rect 409 267 410 268 
<< pdiffusion >>
rect 410 267 411 268 
<< pdiffusion >>
rect 411 267 412 268 
<< pdiffusion >>
rect 412 267 413 268 
<< pdiffusion >>
rect 413 267 414 268 
<< pdiffusion >>
rect 426 267 427 268 
<< pdiffusion >>
rect 427 267 428 268 
<< pdiffusion >>
rect 428 267 429 268 
<< pdiffusion >>
rect 429 267 430 268 
<< pdiffusion >>
rect 430 267 431 268 
<< pdiffusion >>
rect 431 267 432 268 
<< pdiffusion >>
rect 444 267 445 268 
<< pdiffusion >>
rect 445 267 446 268 
<< pdiffusion >>
rect 446 267 447 268 
<< pdiffusion >>
rect 447 267 448 268 
<< pdiffusion >>
rect 448 267 449 268 
<< pdiffusion >>
rect 449 267 450 268 
<< pdiffusion >>
rect 12 268 13 269 
<< pdiffusion >>
rect 13 268 14 269 
<< pdiffusion >>
rect 14 268 15 269 
<< pdiffusion >>
rect 15 268 16 269 
<< pdiffusion >>
rect 16 268 17 269 
<< pdiffusion >>
rect 17 268 18 269 
<< pdiffusion >>
rect 48 268 49 269 
<< pdiffusion >>
rect 49 268 50 269 
<< pdiffusion >>
rect 50 268 51 269 
<< pdiffusion >>
rect 51 268 52 269 
<< pdiffusion >>
rect 52 268 53 269 
<< pdiffusion >>
rect 53 268 54 269 
<< m1 >>
rect 55 268 56 269 
<< m1 >>
rect 64 268 65 269 
<< pdiffusion >>
rect 66 268 67 269 
<< pdiffusion >>
rect 67 268 68 269 
<< pdiffusion >>
rect 68 268 69 269 
<< pdiffusion >>
rect 69 268 70 269 
<< pdiffusion >>
rect 70 268 71 269 
<< pdiffusion >>
rect 71 268 72 269 
<< pdiffusion >>
rect 84 268 85 269 
<< pdiffusion >>
rect 85 268 86 269 
<< pdiffusion >>
rect 86 268 87 269 
<< pdiffusion >>
rect 87 268 88 269 
<< pdiffusion >>
rect 88 268 89 269 
<< pdiffusion >>
rect 89 268 90 269 
<< pdiffusion >>
rect 102 268 103 269 
<< pdiffusion >>
rect 103 268 104 269 
<< pdiffusion >>
rect 104 268 105 269 
<< pdiffusion >>
rect 105 268 106 269 
<< pdiffusion >>
rect 106 268 107 269 
<< pdiffusion >>
rect 107 268 108 269 
<< pdiffusion >>
rect 120 268 121 269 
<< pdiffusion >>
rect 121 268 122 269 
<< pdiffusion >>
rect 122 268 123 269 
<< pdiffusion >>
rect 123 268 124 269 
<< pdiffusion >>
rect 124 268 125 269 
<< pdiffusion >>
rect 125 268 126 269 
<< pdiffusion >>
rect 156 268 157 269 
<< pdiffusion >>
rect 157 268 158 269 
<< pdiffusion >>
rect 158 268 159 269 
<< pdiffusion >>
rect 159 268 160 269 
<< pdiffusion >>
rect 160 268 161 269 
<< pdiffusion >>
rect 161 268 162 269 
<< m1 >>
rect 163 268 164 269 
<< pdiffusion >>
rect 174 268 175 269 
<< pdiffusion >>
rect 175 268 176 269 
<< pdiffusion >>
rect 176 268 177 269 
<< pdiffusion >>
rect 177 268 178 269 
<< pdiffusion >>
rect 178 268 179 269 
<< pdiffusion >>
rect 179 268 180 269 
<< m1 >>
rect 181 268 182 269 
<< m2 >>
rect 182 268 183 269 
<< pdiffusion >>
rect 192 268 193 269 
<< pdiffusion >>
rect 193 268 194 269 
<< pdiffusion >>
rect 194 268 195 269 
<< pdiffusion >>
rect 195 268 196 269 
<< pdiffusion >>
rect 196 268 197 269 
<< pdiffusion >>
rect 197 268 198 269 
<< m1 >>
rect 206 268 207 269 
<< m1 >>
rect 208 268 209 269 
<< pdiffusion >>
rect 210 268 211 269 
<< pdiffusion >>
rect 211 268 212 269 
<< pdiffusion >>
rect 212 268 213 269 
<< pdiffusion >>
rect 213 268 214 269 
<< pdiffusion >>
rect 214 268 215 269 
<< pdiffusion >>
rect 215 268 216 269 
<< pdiffusion >>
rect 228 268 229 269 
<< pdiffusion >>
rect 229 268 230 269 
<< pdiffusion >>
rect 230 268 231 269 
<< pdiffusion >>
rect 231 268 232 269 
<< pdiffusion >>
rect 232 268 233 269 
<< pdiffusion >>
rect 233 268 234 269 
<< m2 >>
rect 243 268 244 269 
<< m1 >>
rect 244 268 245 269 
<< pdiffusion >>
rect 246 268 247 269 
<< pdiffusion >>
rect 247 268 248 269 
<< pdiffusion >>
rect 248 268 249 269 
<< pdiffusion >>
rect 249 268 250 269 
<< pdiffusion >>
rect 250 268 251 269 
<< pdiffusion >>
rect 251 268 252 269 
<< m1 >>
rect 254 268 255 269 
<< m1 >>
rect 262 268 263 269 
<< pdiffusion >>
rect 264 268 265 269 
<< pdiffusion >>
rect 265 268 266 269 
<< pdiffusion >>
rect 266 268 267 269 
<< pdiffusion >>
rect 267 268 268 269 
<< pdiffusion >>
rect 268 268 269 269 
<< pdiffusion >>
rect 269 268 270 269 
<< m1 >>
rect 271 268 272 269 
<< m2 >>
rect 272 268 273 269 
<< pdiffusion >>
rect 282 268 283 269 
<< pdiffusion >>
rect 283 268 284 269 
<< pdiffusion >>
rect 284 268 285 269 
<< pdiffusion >>
rect 285 268 286 269 
<< pdiffusion >>
rect 286 268 287 269 
<< pdiffusion >>
rect 287 268 288 269 
<< m1 >>
rect 298 268 299 269 
<< pdiffusion >>
rect 300 268 301 269 
<< pdiffusion >>
rect 301 268 302 269 
<< pdiffusion >>
rect 302 268 303 269 
<< pdiffusion >>
rect 303 268 304 269 
<< pdiffusion >>
rect 304 268 305 269 
<< pdiffusion >>
rect 305 268 306 269 
<< m1 >>
rect 307 268 308 269 
<< m2 >>
rect 307 268 308 269 
<< pdiffusion >>
rect 318 268 319 269 
<< pdiffusion >>
rect 319 268 320 269 
<< pdiffusion >>
rect 320 268 321 269 
<< pdiffusion >>
rect 321 268 322 269 
<< pdiffusion >>
rect 322 268 323 269 
<< pdiffusion >>
rect 323 268 324 269 
<< m1 >>
rect 325 268 326 269 
<< pdiffusion >>
rect 336 268 337 269 
<< pdiffusion >>
rect 337 268 338 269 
<< pdiffusion >>
rect 338 268 339 269 
<< pdiffusion >>
rect 339 268 340 269 
<< pdiffusion >>
rect 340 268 341 269 
<< pdiffusion >>
rect 341 268 342 269 
<< m1 >>
rect 350 268 351 269 
<< m1 >>
rect 352 268 353 269 
<< m2 >>
rect 352 268 353 269 
<< pdiffusion >>
rect 354 268 355 269 
<< pdiffusion >>
rect 355 268 356 269 
<< pdiffusion >>
rect 356 268 357 269 
<< pdiffusion >>
rect 357 268 358 269 
<< pdiffusion >>
rect 358 268 359 269 
<< pdiffusion >>
rect 359 268 360 269 
<< pdiffusion >>
rect 372 268 373 269 
<< pdiffusion >>
rect 373 268 374 269 
<< pdiffusion >>
rect 374 268 375 269 
<< pdiffusion >>
rect 375 268 376 269 
<< pdiffusion >>
rect 376 268 377 269 
<< pdiffusion >>
rect 377 268 378 269 
<< m1 >>
rect 379 268 380 269 
<< m1 >>
rect 388 268 389 269 
<< pdiffusion >>
rect 390 268 391 269 
<< pdiffusion >>
rect 391 268 392 269 
<< pdiffusion >>
rect 392 268 393 269 
<< pdiffusion >>
rect 393 268 394 269 
<< pdiffusion >>
rect 394 268 395 269 
<< pdiffusion >>
rect 395 268 396 269 
<< pdiffusion >>
rect 408 268 409 269 
<< pdiffusion >>
rect 409 268 410 269 
<< pdiffusion >>
rect 410 268 411 269 
<< pdiffusion >>
rect 411 268 412 269 
<< pdiffusion >>
rect 412 268 413 269 
<< pdiffusion >>
rect 413 268 414 269 
<< pdiffusion >>
rect 426 268 427 269 
<< pdiffusion >>
rect 427 268 428 269 
<< pdiffusion >>
rect 428 268 429 269 
<< pdiffusion >>
rect 429 268 430 269 
<< pdiffusion >>
rect 430 268 431 269 
<< pdiffusion >>
rect 431 268 432 269 
<< pdiffusion >>
rect 444 268 445 269 
<< pdiffusion >>
rect 445 268 446 269 
<< pdiffusion >>
rect 446 268 447 269 
<< pdiffusion >>
rect 447 268 448 269 
<< pdiffusion >>
rect 448 268 449 269 
<< pdiffusion >>
rect 449 268 450 269 
<< pdiffusion >>
rect 12 269 13 270 
<< pdiffusion >>
rect 13 269 14 270 
<< pdiffusion >>
rect 14 269 15 270 
<< pdiffusion >>
rect 15 269 16 270 
<< pdiffusion >>
rect 16 269 17 270 
<< pdiffusion >>
rect 17 269 18 270 
<< pdiffusion >>
rect 48 269 49 270 
<< pdiffusion >>
rect 49 269 50 270 
<< pdiffusion >>
rect 50 269 51 270 
<< pdiffusion >>
rect 51 269 52 270 
<< pdiffusion >>
rect 52 269 53 270 
<< pdiffusion >>
rect 53 269 54 270 
<< m1 >>
rect 55 269 56 270 
<< m1 >>
rect 64 269 65 270 
<< pdiffusion >>
rect 66 269 67 270 
<< pdiffusion >>
rect 67 269 68 270 
<< pdiffusion >>
rect 68 269 69 270 
<< pdiffusion >>
rect 69 269 70 270 
<< m1 >>
rect 70 269 71 270 
<< pdiffusion >>
rect 70 269 71 270 
<< pdiffusion >>
rect 71 269 72 270 
<< pdiffusion >>
rect 84 269 85 270 
<< pdiffusion >>
rect 85 269 86 270 
<< pdiffusion >>
rect 86 269 87 270 
<< pdiffusion >>
rect 87 269 88 270 
<< m1 >>
rect 88 269 89 270 
<< pdiffusion >>
rect 88 269 89 270 
<< pdiffusion >>
rect 89 269 90 270 
<< pdiffusion >>
rect 102 269 103 270 
<< pdiffusion >>
rect 103 269 104 270 
<< pdiffusion >>
rect 104 269 105 270 
<< pdiffusion >>
rect 105 269 106 270 
<< pdiffusion >>
rect 106 269 107 270 
<< pdiffusion >>
rect 107 269 108 270 
<< pdiffusion >>
rect 120 269 121 270 
<< pdiffusion >>
rect 121 269 122 270 
<< pdiffusion >>
rect 122 269 123 270 
<< pdiffusion >>
rect 123 269 124 270 
<< m1 >>
rect 124 269 125 270 
<< pdiffusion >>
rect 124 269 125 270 
<< pdiffusion >>
rect 125 269 126 270 
<< pdiffusion >>
rect 156 269 157 270 
<< m1 >>
rect 157 269 158 270 
<< pdiffusion >>
rect 157 269 158 270 
<< pdiffusion >>
rect 158 269 159 270 
<< pdiffusion >>
rect 159 269 160 270 
<< m1 >>
rect 160 269 161 270 
<< pdiffusion >>
rect 160 269 161 270 
<< pdiffusion >>
rect 161 269 162 270 
<< m1 >>
rect 163 269 164 270 
<< pdiffusion >>
rect 174 269 175 270 
<< pdiffusion >>
rect 175 269 176 270 
<< pdiffusion >>
rect 176 269 177 270 
<< pdiffusion >>
rect 177 269 178 270 
<< pdiffusion >>
rect 178 269 179 270 
<< pdiffusion >>
rect 179 269 180 270 
<< m1 >>
rect 181 269 182 270 
<< m2 >>
rect 182 269 183 270 
<< pdiffusion >>
rect 192 269 193 270 
<< m1 >>
rect 193 269 194 270 
<< pdiffusion >>
rect 193 269 194 270 
<< pdiffusion >>
rect 194 269 195 270 
<< pdiffusion >>
rect 195 269 196 270 
<< pdiffusion >>
rect 196 269 197 270 
<< pdiffusion >>
rect 197 269 198 270 
<< m1 >>
rect 206 269 207 270 
<< m1 >>
rect 208 269 209 270 
<< pdiffusion >>
rect 210 269 211 270 
<< pdiffusion >>
rect 211 269 212 270 
<< pdiffusion >>
rect 212 269 213 270 
<< pdiffusion >>
rect 213 269 214 270 
<< pdiffusion >>
rect 214 269 215 270 
<< pdiffusion >>
rect 215 269 216 270 
<< pdiffusion >>
rect 228 269 229 270 
<< pdiffusion >>
rect 229 269 230 270 
<< pdiffusion >>
rect 230 269 231 270 
<< pdiffusion >>
rect 231 269 232 270 
<< pdiffusion >>
rect 232 269 233 270 
<< pdiffusion >>
rect 233 269 234 270 
<< m2 >>
rect 243 269 244 270 
<< m1 >>
rect 244 269 245 270 
<< pdiffusion >>
rect 246 269 247 270 
<< m1 >>
rect 247 269 248 270 
<< pdiffusion >>
rect 247 269 248 270 
<< pdiffusion >>
rect 248 269 249 270 
<< pdiffusion >>
rect 249 269 250 270 
<< pdiffusion >>
rect 250 269 251 270 
<< pdiffusion >>
rect 251 269 252 270 
<< m1 >>
rect 254 269 255 270 
<< m1 >>
rect 262 269 263 270 
<< pdiffusion >>
rect 264 269 265 270 
<< m1 >>
rect 265 269 266 270 
<< pdiffusion >>
rect 265 269 266 270 
<< pdiffusion >>
rect 266 269 267 270 
<< pdiffusion >>
rect 267 269 268 270 
<< pdiffusion >>
rect 268 269 269 270 
<< pdiffusion >>
rect 269 269 270 270 
<< m1 >>
rect 271 269 272 270 
<< m2 >>
rect 272 269 273 270 
<< pdiffusion >>
rect 282 269 283 270 
<< pdiffusion >>
rect 283 269 284 270 
<< pdiffusion >>
rect 284 269 285 270 
<< pdiffusion >>
rect 285 269 286 270 
<< pdiffusion >>
rect 286 269 287 270 
<< pdiffusion >>
rect 287 269 288 270 
<< m1 >>
rect 298 269 299 270 
<< pdiffusion >>
rect 300 269 301 270 
<< m1 >>
rect 301 269 302 270 
<< pdiffusion >>
rect 301 269 302 270 
<< pdiffusion >>
rect 302 269 303 270 
<< pdiffusion >>
rect 303 269 304 270 
<< pdiffusion >>
rect 304 269 305 270 
<< pdiffusion >>
rect 305 269 306 270 
<< m1 >>
rect 307 269 308 270 
<< m2 >>
rect 307 269 308 270 
<< pdiffusion >>
rect 318 269 319 270 
<< pdiffusion >>
rect 319 269 320 270 
<< pdiffusion >>
rect 320 269 321 270 
<< pdiffusion >>
rect 321 269 322 270 
<< pdiffusion >>
rect 322 269 323 270 
<< pdiffusion >>
rect 323 269 324 270 
<< m1 >>
rect 325 269 326 270 
<< pdiffusion >>
rect 336 269 337 270 
<< pdiffusion >>
rect 337 269 338 270 
<< pdiffusion >>
rect 338 269 339 270 
<< pdiffusion >>
rect 339 269 340 270 
<< m1 >>
rect 340 269 341 270 
<< pdiffusion >>
rect 340 269 341 270 
<< pdiffusion >>
rect 341 269 342 270 
<< m1 >>
rect 350 269 351 270 
<< m2 >>
rect 350 269 351 270 
<< m2c >>
rect 350 269 351 270 
<< m1 >>
rect 350 269 351 270 
<< m2 >>
rect 350 269 351 270 
<< m1 >>
rect 352 269 353 270 
<< m2 >>
rect 352 269 353 270 
<< pdiffusion >>
rect 354 269 355 270 
<< pdiffusion >>
rect 355 269 356 270 
<< pdiffusion >>
rect 356 269 357 270 
<< pdiffusion >>
rect 357 269 358 270 
<< pdiffusion >>
rect 358 269 359 270 
<< pdiffusion >>
rect 359 269 360 270 
<< pdiffusion >>
rect 372 269 373 270 
<< pdiffusion >>
rect 373 269 374 270 
<< pdiffusion >>
rect 374 269 375 270 
<< pdiffusion >>
rect 375 269 376 270 
<< pdiffusion >>
rect 376 269 377 270 
<< pdiffusion >>
rect 377 269 378 270 
<< m1 >>
rect 379 269 380 270 
<< m1 >>
rect 388 269 389 270 
<< pdiffusion >>
rect 390 269 391 270 
<< m1 >>
rect 391 269 392 270 
<< pdiffusion >>
rect 391 269 392 270 
<< pdiffusion >>
rect 392 269 393 270 
<< pdiffusion >>
rect 393 269 394 270 
<< pdiffusion >>
rect 394 269 395 270 
<< pdiffusion >>
rect 395 269 396 270 
<< pdiffusion >>
rect 408 269 409 270 
<< pdiffusion >>
rect 409 269 410 270 
<< pdiffusion >>
rect 410 269 411 270 
<< pdiffusion >>
rect 411 269 412 270 
<< m1 >>
rect 412 269 413 270 
<< pdiffusion >>
rect 412 269 413 270 
<< pdiffusion >>
rect 413 269 414 270 
<< pdiffusion >>
rect 426 269 427 270 
<< pdiffusion >>
rect 427 269 428 270 
<< pdiffusion >>
rect 428 269 429 270 
<< pdiffusion >>
rect 429 269 430 270 
<< pdiffusion >>
rect 430 269 431 270 
<< pdiffusion >>
rect 431 269 432 270 
<< pdiffusion >>
rect 444 269 445 270 
<< pdiffusion >>
rect 445 269 446 270 
<< pdiffusion >>
rect 446 269 447 270 
<< pdiffusion >>
rect 447 269 448 270 
<< pdiffusion >>
rect 448 269 449 270 
<< pdiffusion >>
rect 449 269 450 270 
<< m1 >>
rect 55 270 56 271 
<< m1 >>
rect 64 270 65 271 
<< m1 >>
rect 70 270 71 271 
<< m1 >>
rect 88 270 89 271 
<< m1 >>
rect 124 270 125 271 
<< m1 >>
rect 157 270 158 271 
<< m1 >>
rect 160 270 161 271 
<< m1 >>
rect 163 270 164 271 
<< m1 >>
rect 181 270 182 271 
<< m2 >>
rect 182 270 183 271 
<< m1 >>
rect 193 270 194 271 
<< m1 >>
rect 206 270 207 271 
<< m2 >>
rect 206 270 207 271 
<< m2c >>
rect 206 270 207 271 
<< m1 >>
rect 206 270 207 271 
<< m2 >>
rect 206 270 207 271 
<< m2 >>
rect 207 270 208 271 
<< m1 >>
rect 208 270 209 271 
<< m2 >>
rect 208 270 209 271 
<< m2 >>
rect 243 270 244 271 
<< m1 >>
rect 244 270 245 271 
<< m1 >>
rect 247 270 248 271 
<< m1 >>
rect 254 270 255 271 
<< m1 >>
rect 262 270 263 271 
<< m1 >>
rect 265 270 266 271 
<< m1 >>
rect 271 270 272 271 
<< m2 >>
rect 272 270 273 271 
<< m1 >>
rect 298 270 299 271 
<< m1 >>
rect 301 270 302 271 
<< m1 >>
rect 307 270 308 271 
<< m2 >>
rect 307 270 308 271 
<< m1 >>
rect 325 270 326 271 
<< m1 >>
rect 340 270 341 271 
<< m2 >>
rect 350 270 351 271 
<< m1 >>
rect 352 270 353 271 
<< m2 >>
rect 352 270 353 271 
<< m1 >>
rect 379 270 380 271 
<< m1 >>
rect 388 270 389 271 
<< m1 >>
rect 391 270 392 271 
<< m1 >>
rect 412 270 413 271 
<< m1 >>
rect 55 271 56 272 
<< m1 >>
rect 64 271 65 272 
<< m1 >>
rect 70 271 71 272 
<< m1 >>
rect 88 271 89 272 
<< m1 >>
rect 124 271 125 272 
<< m1 >>
rect 157 271 158 272 
<< m1 >>
rect 160 271 161 272 
<< m1 >>
rect 161 271 162 272 
<< m1 >>
rect 162 271 163 272 
<< m1 >>
rect 163 271 164 272 
<< m1 >>
rect 181 271 182 272 
<< m2 >>
rect 182 271 183 272 
<< m1 >>
rect 193 271 194 272 
<< m1 >>
rect 208 271 209 272 
<< m2 >>
rect 208 271 209 272 
<< m2 >>
rect 243 271 244 272 
<< m1 >>
rect 244 271 245 272 
<< m1 >>
rect 247 271 248 272 
<< m1 >>
rect 254 271 255 272 
<< m1 >>
rect 262 271 263 272 
<< m1 >>
rect 265 271 266 272 
<< m1 >>
rect 269 271 270 272 
<< m2 >>
rect 269 271 270 272 
<< m2c >>
rect 269 271 270 272 
<< m1 >>
rect 269 271 270 272 
<< m2 >>
rect 269 271 270 272 
<< m2 >>
rect 270 271 271 272 
<< m1 >>
rect 271 271 272 272 
<< m2 >>
rect 271 271 272 272 
<< m2 >>
rect 272 271 273 272 
<< m1 >>
rect 298 271 299 272 
<< m1 >>
rect 301 271 302 272 
<< m1 >>
rect 307 271 308 272 
<< m2 >>
rect 307 271 308 272 
<< m1 >>
rect 325 271 326 272 
<< m1 >>
rect 340 271 341 272 
<< m1 >>
rect 341 271 342 272 
<< m1 >>
rect 342 271 343 272 
<< m1 >>
rect 343 271 344 272 
<< m1 >>
rect 344 271 345 272 
<< m1 >>
rect 345 271 346 272 
<< m1 >>
rect 346 271 347 272 
<< m1 >>
rect 347 271 348 272 
<< m1 >>
rect 348 271 349 272 
<< m1 >>
rect 349 271 350 272 
<< m1 >>
rect 350 271 351 272 
<< m2 >>
rect 350 271 351 272 
<< m1 >>
rect 351 271 352 272 
<< m1 >>
rect 352 271 353 272 
<< m2 >>
rect 352 271 353 272 
<< m1 >>
rect 379 271 380 272 
<< m1 >>
rect 388 271 389 272 
<< m1 >>
rect 389 271 390 272 
<< m1 >>
rect 390 271 391 272 
<< m1 >>
rect 391 271 392 272 
<< m1 >>
rect 412 271 413 272 
<< m1 >>
rect 55 272 56 273 
<< m1 >>
rect 64 272 65 273 
<< m1 >>
rect 70 272 71 273 
<< m1 >>
rect 88 272 89 273 
<< m1 >>
rect 124 272 125 273 
<< m1 >>
rect 157 272 158 273 
<< m1 >>
rect 181 272 182 273 
<< m2 >>
rect 182 272 183 273 
<< m1 >>
rect 193 272 194 273 
<< m1 >>
rect 194 272 195 273 
<< m1 >>
rect 195 272 196 273 
<< m1 >>
rect 196 272 197 273 
<< m1 >>
rect 197 272 198 273 
<< m1 >>
rect 198 272 199 273 
<< m1 >>
rect 199 272 200 273 
<< m1 >>
rect 200 272 201 273 
<< m1 >>
rect 201 272 202 273 
<< m1 >>
rect 202 272 203 273 
<< m1 >>
rect 203 272 204 273 
<< m1 >>
rect 204 272 205 273 
<< m1 >>
rect 205 272 206 273 
<< m1 >>
rect 206 272 207 273 
<< m1 >>
rect 207 272 208 273 
<< m1 >>
rect 208 272 209 273 
<< m2 >>
rect 208 272 209 273 
<< m2 >>
rect 243 272 244 273 
<< m1 >>
rect 244 272 245 273 
<< m1 >>
rect 247 272 248 273 
<< m1 >>
rect 254 272 255 273 
<< m1 >>
rect 262 272 263 273 
<< m1 >>
rect 265 272 266 273 
<< m1 >>
rect 266 272 267 273 
<< m1 >>
rect 267 272 268 273 
<< m1 >>
rect 268 272 269 273 
<< m1 >>
rect 269 272 270 273 
<< m1 >>
rect 271 272 272 273 
<< m1 >>
rect 298 272 299 273 
<< m1 >>
rect 301 272 302 273 
<< m1 >>
rect 302 272 303 273 
<< m1 >>
rect 303 272 304 273 
<< m1 >>
rect 304 272 305 273 
<< m1 >>
rect 305 272 306 273 
<< m2 >>
rect 305 272 306 273 
<< m2c >>
rect 305 272 306 273 
<< m1 >>
rect 305 272 306 273 
<< m2 >>
rect 305 272 306 273 
<< m2 >>
rect 306 272 307 273 
<< m1 >>
rect 307 272 308 273 
<< m2 >>
rect 307 272 308 273 
<< m1 >>
rect 325 272 326 273 
<< m2 >>
rect 350 272 351 273 
<< m2 >>
rect 352 272 353 273 
<< m1 >>
rect 379 272 380 273 
<< m1 >>
rect 412 272 413 273 
<< m1 >>
rect 55 273 56 274 
<< m1 >>
rect 64 273 65 274 
<< m1 >>
rect 70 273 71 274 
<< m1 >>
rect 88 273 89 274 
<< m1 >>
rect 124 273 125 274 
<< m1 >>
rect 157 273 158 274 
<< m1 >>
rect 158 273 159 274 
<< m1 >>
rect 159 273 160 274 
<< m1 >>
rect 160 273 161 274 
<< m1 >>
rect 161 273 162 274 
<< m1 >>
rect 162 273 163 274 
<< m1 >>
rect 163 273 164 274 
<< m1 >>
rect 181 273 182 274 
<< m2 >>
rect 182 273 183 274 
<< m2 >>
rect 208 273 209 274 
<< m2 >>
rect 209 273 210 274 
<< m1 >>
rect 210 273 211 274 
<< m2 >>
rect 210 273 211 274 
<< m2c >>
rect 210 273 211 274 
<< m1 >>
rect 210 273 211 274 
<< m2 >>
rect 210 273 211 274 
<< m2 >>
rect 243 273 244 274 
<< m1 >>
rect 244 273 245 274 
<< m1 >>
rect 247 273 248 274 
<< m1 >>
rect 254 273 255 274 
<< m1 >>
rect 262 273 263 274 
<< m1 >>
rect 271 273 272 274 
<< m1 >>
rect 298 273 299 274 
<< m1 >>
rect 307 273 308 274 
<< m1 >>
rect 325 273 326 274 
<< m1 >>
rect 350 273 351 274 
<< m2 >>
rect 350 273 351 274 
<< m2c >>
rect 350 273 351 274 
<< m1 >>
rect 350 273 351 274 
<< m2 >>
rect 350 273 351 274 
<< m1 >>
rect 352 273 353 274 
<< m2 >>
rect 352 273 353 274 
<< m2c >>
rect 352 273 353 274 
<< m1 >>
rect 352 273 353 274 
<< m2 >>
rect 352 273 353 274 
<< m1 >>
rect 379 273 380 274 
<< m1 >>
rect 412 273 413 274 
<< m1 >>
rect 55 274 56 275 
<< m1 >>
rect 64 274 65 275 
<< m1 >>
rect 70 274 71 275 
<< m1 >>
rect 71 274 72 275 
<< m1 >>
rect 72 274 73 275 
<< m1 >>
rect 73 274 74 275 
<< m1 >>
rect 74 274 75 275 
<< m1 >>
rect 75 274 76 275 
<< m1 >>
rect 76 274 77 275 
<< m1 >>
rect 77 274 78 275 
<< m1 >>
rect 78 274 79 275 
<< m1 >>
rect 79 274 80 275 
<< m1 >>
rect 80 274 81 275 
<< m1 >>
rect 81 274 82 275 
<< m1 >>
rect 82 274 83 275 
<< m1 >>
rect 83 274 84 275 
<< m1 >>
rect 84 274 85 275 
<< m1 >>
rect 85 274 86 275 
<< m1 >>
rect 86 274 87 275 
<< m1 >>
rect 87 274 88 275 
<< m1 >>
rect 88 274 89 275 
<< m1 >>
rect 124 274 125 275 
<< m1 >>
rect 163 274 164 275 
<< m1 >>
rect 181 274 182 275 
<< m2 >>
rect 182 274 183 275 
<< m1 >>
rect 210 274 211 275 
<< m2 >>
rect 243 274 244 275 
<< m1 >>
rect 244 274 245 275 
<< m1 >>
rect 247 274 248 275 
<< m1 >>
rect 254 274 255 275 
<< m1 >>
rect 262 274 263 275 
<< m1 >>
rect 271 274 272 275 
<< m1 >>
rect 298 274 299 275 
<< m1 >>
rect 299 274 300 275 
<< m1 >>
rect 300 274 301 275 
<< m1 >>
rect 301 274 302 275 
<< m1 >>
rect 302 274 303 275 
<< m1 >>
rect 303 274 304 275 
<< m1 >>
rect 304 274 305 275 
<< m1 >>
rect 305 274 306 275 
<< m2 >>
rect 305 274 306 275 
<< m2c >>
rect 305 274 306 275 
<< m1 >>
rect 305 274 306 275 
<< m2 >>
rect 305 274 306 275 
<< m2 >>
rect 306 274 307 275 
<< m1 >>
rect 307 274 308 275 
<< m2 >>
rect 307 274 308 275 
<< m2 >>
rect 308 274 309 275 
<< m1 >>
rect 309 274 310 275 
<< m2 >>
rect 309 274 310 275 
<< m2c >>
rect 309 274 310 275 
<< m1 >>
rect 309 274 310 275 
<< m2 >>
rect 309 274 310 275 
<< m1 >>
rect 310 274 311 275 
<< m1 >>
rect 311 274 312 275 
<< m1 >>
rect 312 274 313 275 
<< m1 >>
rect 313 274 314 275 
<< m1 >>
rect 314 274 315 275 
<< m1 >>
rect 315 274 316 275 
<< m1 >>
rect 316 274 317 275 
<< m1 >>
rect 317 274 318 275 
<< m1 >>
rect 318 274 319 275 
<< m1 >>
rect 319 274 320 275 
<< m1 >>
rect 320 274 321 275 
<< m1 >>
rect 321 274 322 275 
<< m1 >>
rect 322 274 323 275 
<< m1 >>
rect 323 274 324 275 
<< m1 >>
rect 324 274 325 275 
<< m1 >>
rect 325 274 326 275 
<< m1 >>
rect 350 274 351 275 
<< m1 >>
rect 352 274 353 275 
<< m1 >>
rect 379 274 380 275 
<< m1 >>
rect 380 274 381 275 
<< m1 >>
rect 381 274 382 275 
<< m1 >>
rect 382 274 383 275 
<< m1 >>
rect 383 274 384 275 
<< m1 >>
rect 384 274 385 275 
<< m1 >>
rect 385 274 386 275 
<< m1 >>
rect 386 274 387 275 
<< m1 >>
rect 387 274 388 275 
<< m1 >>
rect 388 274 389 275 
<< m1 >>
rect 389 274 390 275 
<< m1 >>
rect 390 274 391 275 
<< m1 >>
rect 391 274 392 275 
<< m1 >>
rect 392 274 393 275 
<< m1 >>
rect 393 274 394 275 
<< m1 >>
rect 394 274 395 275 
<< m1 >>
rect 395 274 396 275 
<< m1 >>
rect 396 274 397 275 
<< m1 >>
rect 397 274 398 275 
<< m1 >>
rect 398 274 399 275 
<< m1 >>
rect 399 274 400 275 
<< m1 >>
rect 400 274 401 275 
<< m1 >>
rect 401 274 402 275 
<< m1 >>
rect 402 274 403 275 
<< m1 >>
rect 403 274 404 275 
<< m1 >>
rect 404 274 405 275 
<< m1 >>
rect 405 274 406 275 
<< m1 >>
rect 406 274 407 275 
<< m1 >>
rect 407 274 408 275 
<< m1 >>
rect 408 274 409 275 
<< m1 >>
rect 409 274 410 275 
<< m1 >>
rect 410 274 411 275 
<< m2 >>
rect 410 274 411 275 
<< m2c >>
rect 410 274 411 275 
<< m1 >>
rect 410 274 411 275 
<< m2 >>
rect 410 274 411 275 
<< m2 >>
rect 411 274 412 275 
<< m1 >>
rect 412 274 413 275 
<< m2 >>
rect 412 274 413 275 
<< m2 >>
rect 413 274 414 275 
<< m1 >>
rect 414 274 415 275 
<< m2 >>
rect 414 274 415 275 
<< m2c >>
rect 414 274 415 275 
<< m1 >>
rect 414 274 415 275 
<< m2 >>
rect 414 274 415 275 
<< m1 >>
rect 415 274 416 275 
<< m1 >>
rect 416 274 417 275 
<< m1 >>
rect 417 274 418 275 
<< m1 >>
rect 418 274 419 275 
<< m1 >>
rect 419 274 420 275 
<< m1 >>
rect 420 274 421 275 
<< m1 >>
rect 421 274 422 275 
<< m1 >>
rect 422 274 423 275 
<< m1 >>
rect 423 274 424 275 
<< m1 >>
rect 424 274 425 275 
<< m1 >>
rect 425 274 426 275 
<< m1 >>
rect 426 274 427 275 
<< m1 >>
rect 427 274 428 275 
<< m1 >>
rect 428 274 429 275 
<< m1 >>
rect 429 274 430 275 
<< m1 >>
rect 430 274 431 275 
<< m1 >>
rect 431 274 432 275 
<< m1 >>
rect 432 274 433 275 
<< m1 >>
rect 433 274 434 275 
<< m1 >>
rect 434 274 435 275 
<< m1 >>
rect 435 274 436 275 
<< m1 >>
rect 436 274 437 275 
<< m1 >>
rect 437 274 438 275 
<< m1 >>
rect 438 274 439 275 
<< m1 >>
rect 439 274 440 275 
<< m1 >>
rect 440 274 441 275 
<< m1 >>
rect 441 274 442 275 
<< m1 >>
rect 442 274 443 275 
<< m1 >>
rect 443 274 444 275 
<< m1 >>
rect 444 274 445 275 
<< m1 >>
rect 445 274 446 275 
<< m1 >>
rect 55 275 56 276 
<< m1 >>
rect 64 275 65 276 
<< m1 >>
rect 124 275 125 276 
<< m1 >>
rect 163 275 164 276 
<< m1 >>
rect 181 275 182 276 
<< m2 >>
rect 182 275 183 276 
<< m1 >>
rect 210 275 211 276 
<< m2 >>
rect 243 275 244 276 
<< m1 >>
rect 244 275 245 276 
<< m1 >>
rect 247 275 248 276 
<< m1 >>
rect 254 275 255 276 
<< m2 >>
rect 254 275 255 276 
<< m2c >>
rect 254 275 255 276 
<< m1 >>
rect 254 275 255 276 
<< m2 >>
rect 254 275 255 276 
<< m1 >>
rect 262 275 263 276 
<< m1 >>
rect 271 275 272 276 
<< m1 >>
rect 307 275 308 276 
<< m1 >>
rect 350 275 351 276 
<< m2 >>
rect 350 275 351 276 
<< m2c >>
rect 350 275 351 276 
<< m1 >>
rect 350 275 351 276 
<< m2 >>
rect 350 275 351 276 
<< m1 >>
rect 352 275 353 276 
<< m2 >>
rect 352 275 353 276 
<< m2c >>
rect 352 275 353 276 
<< m1 >>
rect 352 275 353 276 
<< m2 >>
rect 352 275 353 276 
<< m1 >>
rect 412 275 413 276 
<< m1 >>
rect 445 275 446 276 
<< m1 >>
rect 55 276 56 277 
<< m1 >>
rect 64 276 65 277 
<< m1 >>
rect 124 276 125 277 
<< m1 >>
rect 163 276 164 277 
<< m1 >>
rect 181 276 182 277 
<< m2 >>
rect 182 276 183 277 
<< m1 >>
rect 210 276 211 277 
<< m2 >>
rect 243 276 244 277 
<< m1 >>
rect 244 276 245 277 
<< m1 >>
rect 247 276 248 277 
<< m2 >>
rect 254 276 255 277 
<< m1 >>
rect 262 276 263 277 
<< m1 >>
rect 271 276 272 277 
<< m1 >>
rect 307 276 308 277 
<< m2 >>
rect 318 276 319 277 
<< m2 >>
rect 319 276 320 277 
<< m2 >>
rect 320 276 321 277 
<< m2 >>
rect 321 276 322 277 
<< m2 >>
rect 322 276 323 277 
<< m2 >>
rect 323 276 324 277 
<< m2 >>
rect 324 276 325 277 
<< m2 >>
rect 325 276 326 277 
<< m2 >>
rect 326 276 327 277 
<< m2 >>
rect 327 276 328 277 
<< m2 >>
rect 328 276 329 277 
<< m2 >>
rect 329 276 330 277 
<< m2 >>
rect 330 276 331 277 
<< m2 >>
rect 331 276 332 277 
<< m2 >>
rect 332 276 333 277 
<< m2 >>
rect 333 276 334 277 
<< m2 >>
rect 334 276 335 277 
<< m2 >>
rect 335 276 336 277 
<< m2 >>
rect 336 276 337 277 
<< m2 >>
rect 337 276 338 277 
<< m2 >>
rect 338 276 339 277 
<< m2 >>
rect 339 276 340 277 
<< m2 >>
rect 340 276 341 277 
<< m2 >>
rect 341 276 342 277 
<< m2 >>
rect 342 276 343 277 
<< m2 >>
rect 343 276 344 277 
<< m2 >>
rect 344 276 345 277 
<< m2 >>
rect 345 276 346 277 
<< m2 >>
rect 346 276 347 277 
<< m2 >>
rect 347 276 348 277 
<< m2 >>
rect 348 276 349 277 
<< m2 >>
rect 349 276 350 277 
<< m2 >>
rect 350 276 351 277 
<< m2 >>
rect 352 276 353 277 
<< m1 >>
rect 412 276 413 277 
<< m1 >>
rect 445 276 446 277 
<< m1 >>
rect 55 277 56 278 
<< m1 >>
rect 64 277 65 278 
<< m1 >>
rect 91 277 92 278 
<< m1 >>
rect 92 277 93 278 
<< m1 >>
rect 93 277 94 278 
<< m1 >>
rect 94 277 95 278 
<< m1 >>
rect 95 277 96 278 
<< m1 >>
rect 96 277 97 278 
<< m1 >>
rect 97 277 98 278 
<< m1 >>
rect 98 277 99 278 
<< m1 >>
rect 99 277 100 278 
<< m1 >>
rect 100 277 101 278 
<< m1 >>
rect 101 277 102 278 
<< m1 >>
rect 102 277 103 278 
<< m1 >>
rect 103 277 104 278 
<< m1 >>
rect 104 277 105 278 
<< m1 >>
rect 105 277 106 278 
<< m1 >>
rect 106 277 107 278 
<< m1 >>
rect 107 277 108 278 
<< m1 >>
rect 108 277 109 278 
<< m1 >>
rect 109 277 110 278 
<< m1 >>
rect 110 277 111 278 
<< m1 >>
rect 111 277 112 278 
<< m1 >>
rect 112 277 113 278 
<< m1 >>
rect 113 277 114 278 
<< m1 >>
rect 114 277 115 278 
<< m1 >>
rect 115 277 116 278 
<< m1 >>
rect 116 277 117 278 
<< m1 >>
rect 117 277 118 278 
<< m1 >>
rect 118 277 119 278 
<< m1 >>
rect 119 277 120 278 
<< m1 >>
rect 120 277 121 278 
<< m1 >>
rect 121 277 122 278 
<< m1 >>
rect 122 277 123 278 
<< m1 >>
rect 123 277 124 278 
<< m1 >>
rect 124 277 125 278 
<< m1 >>
rect 127 277 128 278 
<< m1 >>
rect 128 277 129 278 
<< m1 >>
rect 129 277 130 278 
<< m1 >>
rect 130 277 131 278 
<< m1 >>
rect 131 277 132 278 
<< m1 >>
rect 132 277 133 278 
<< m1 >>
rect 133 277 134 278 
<< m1 >>
rect 134 277 135 278 
<< m1 >>
rect 135 277 136 278 
<< m1 >>
rect 136 277 137 278 
<< m1 >>
rect 137 277 138 278 
<< m1 >>
rect 138 277 139 278 
<< m1 >>
rect 139 277 140 278 
<< m1 >>
rect 140 277 141 278 
<< m2 >>
rect 140 277 141 278 
<< m2c >>
rect 140 277 141 278 
<< m1 >>
rect 140 277 141 278 
<< m2 >>
rect 140 277 141 278 
<< m1 >>
rect 163 277 164 278 
<< m1 >>
rect 181 277 182 278 
<< m2 >>
rect 182 277 183 278 
<< m1 >>
rect 210 277 211 278 
<< m1 >>
rect 211 277 212 278 
<< m1 >>
rect 212 277 213 278 
<< m1 >>
rect 213 277 214 278 
<< m1 >>
rect 214 277 215 278 
<< m1 >>
rect 215 277 216 278 
<< m1 >>
rect 216 277 217 278 
<< m1 >>
rect 217 277 218 278 
<< m1 >>
rect 218 277 219 278 
<< m1 >>
rect 219 277 220 278 
<< m1 >>
rect 220 277 221 278 
<< m1 >>
rect 221 277 222 278 
<< m1 >>
rect 222 277 223 278 
<< m1 >>
rect 223 277 224 278 
<< m1 >>
rect 224 277 225 278 
<< m1 >>
rect 225 277 226 278 
<< m1 >>
rect 226 277 227 278 
<< m2 >>
rect 243 277 244 278 
<< m1 >>
rect 244 277 245 278 
<< m1 >>
rect 247 277 248 278 
<< m1 >>
rect 248 277 249 278 
<< m1 >>
rect 249 277 250 278 
<< m1 >>
rect 250 277 251 278 
<< m1 >>
rect 251 277 252 278 
<< m1 >>
rect 252 277 253 278 
<< m1 >>
rect 253 277 254 278 
<< m1 >>
rect 254 277 255 278 
<< m2 >>
rect 254 277 255 278 
<< m1 >>
rect 255 277 256 278 
<< m1 >>
rect 256 277 257 278 
<< m1 >>
rect 257 277 258 278 
<< m1 >>
rect 258 277 259 278 
<< m1 >>
rect 259 277 260 278 
<< m1 >>
rect 260 277 261 278 
<< m1 >>
rect 262 277 263 278 
<< m1 >>
rect 263 277 264 278 
<< m1 >>
rect 264 277 265 278 
<< m1 >>
rect 265 277 266 278 
<< m1 >>
rect 266 277 267 278 
<< m1 >>
rect 267 277 268 278 
<< m1 >>
rect 268 277 269 278 
<< m1 >>
rect 269 277 270 278 
<< m2 >>
rect 269 277 270 278 
<< m2c >>
rect 269 277 270 278 
<< m1 >>
rect 269 277 270 278 
<< m2 >>
rect 269 277 270 278 
<< m2 >>
rect 270 277 271 278 
<< m1 >>
rect 271 277 272 278 
<< m2 >>
rect 271 277 272 278 
<< m2 >>
rect 272 277 273 278 
<< m1 >>
rect 273 277 274 278 
<< m2 >>
rect 273 277 274 278 
<< m2c >>
rect 273 277 274 278 
<< m1 >>
rect 273 277 274 278 
<< m2 >>
rect 273 277 274 278 
<< m1 >>
rect 274 277 275 278 
<< m1 >>
rect 275 277 276 278 
<< m1 >>
rect 276 277 277 278 
<< m1 >>
rect 277 277 278 278 
<< m1 >>
rect 278 277 279 278 
<< m1 >>
rect 279 277 280 278 
<< m1 >>
rect 280 277 281 278 
<< m1 >>
rect 281 277 282 278 
<< m1 >>
rect 282 277 283 278 
<< m1 >>
rect 283 277 284 278 
<< m1 >>
rect 284 277 285 278 
<< m1 >>
rect 285 277 286 278 
<< m1 >>
rect 286 277 287 278 
<< m1 >>
rect 287 277 288 278 
<< m1 >>
rect 288 277 289 278 
<< m1 >>
rect 289 277 290 278 
<< m1 >>
rect 290 277 291 278 
<< m1 >>
rect 291 277 292 278 
<< m1 >>
rect 292 277 293 278 
<< m1 >>
rect 293 277 294 278 
<< m1 >>
rect 294 277 295 278 
<< m1 >>
rect 295 277 296 278 
<< m1 >>
rect 296 277 297 278 
<< m1 >>
rect 297 277 298 278 
<< m1 >>
rect 298 277 299 278 
<< m1 >>
rect 299 277 300 278 
<< m1 >>
rect 300 277 301 278 
<< m1 >>
rect 301 277 302 278 
<< m1 >>
rect 302 277 303 278 
<< m1 >>
rect 303 277 304 278 
<< m1 >>
rect 304 277 305 278 
<< m1 >>
rect 305 277 306 278 
<< m2 >>
rect 305 277 306 278 
<< m2c >>
rect 305 277 306 278 
<< m1 >>
rect 305 277 306 278 
<< m2 >>
rect 305 277 306 278 
<< m2 >>
rect 306 277 307 278 
<< m1 >>
rect 307 277 308 278 
<< m2 >>
rect 307 277 308 278 
<< m2 >>
rect 308 277 309 278 
<< m1 >>
rect 309 277 310 278 
<< m2 >>
rect 309 277 310 278 
<< m2c >>
rect 309 277 310 278 
<< m1 >>
rect 309 277 310 278 
<< m2 >>
rect 309 277 310 278 
<< m1 >>
rect 310 277 311 278 
<< m1 >>
rect 311 277 312 278 
<< m1 >>
rect 312 277 313 278 
<< m1 >>
rect 313 277 314 278 
<< m1 >>
rect 314 277 315 278 
<< m1 >>
rect 315 277 316 278 
<< m1 >>
rect 316 277 317 278 
<< m1 >>
rect 317 277 318 278 
<< m1 >>
rect 318 277 319 278 
<< m2 >>
rect 318 277 319 278 
<< m1 >>
rect 319 277 320 278 
<< m1 >>
rect 320 277 321 278 
<< m1 >>
rect 321 277 322 278 
<< m1 >>
rect 322 277 323 278 
<< m1 >>
rect 323 277 324 278 
<< m1 >>
rect 324 277 325 278 
<< m1 >>
rect 325 277 326 278 
<< m1 >>
rect 326 277 327 278 
<< m1 >>
rect 327 277 328 278 
<< m1 >>
rect 328 277 329 278 
<< m1 >>
rect 329 277 330 278 
<< m1 >>
rect 330 277 331 278 
<< m1 >>
rect 331 277 332 278 
<< m1 >>
rect 332 277 333 278 
<< m1 >>
rect 333 277 334 278 
<< m1 >>
rect 334 277 335 278 
<< m1 >>
rect 335 277 336 278 
<< m1 >>
rect 336 277 337 278 
<< m1 >>
rect 337 277 338 278 
<< m1 >>
rect 338 277 339 278 
<< m1 >>
rect 339 277 340 278 
<< m1 >>
rect 340 277 341 278 
<< m1 >>
rect 341 277 342 278 
<< m1 >>
rect 342 277 343 278 
<< m1 >>
rect 343 277 344 278 
<< m1 >>
rect 344 277 345 278 
<< m1 >>
rect 345 277 346 278 
<< m1 >>
rect 346 277 347 278 
<< m1 >>
rect 347 277 348 278 
<< m1 >>
rect 348 277 349 278 
<< m1 >>
rect 349 277 350 278 
<< m1 >>
rect 350 277 351 278 
<< m1 >>
rect 351 277 352 278 
<< m1 >>
rect 352 277 353 278 
<< m2 >>
rect 352 277 353 278 
<< m1 >>
rect 353 277 354 278 
<< m1 >>
rect 354 277 355 278 
<< m1 >>
rect 355 277 356 278 
<< m1 >>
rect 356 277 357 278 
<< m1 >>
rect 357 277 358 278 
<< m1 >>
rect 358 277 359 278 
<< m1 >>
rect 359 277 360 278 
<< m1 >>
rect 360 277 361 278 
<< m1 >>
rect 361 277 362 278 
<< m1 >>
rect 362 277 363 278 
<< m1 >>
rect 363 277 364 278 
<< m1 >>
rect 364 277 365 278 
<< m1 >>
rect 365 277 366 278 
<< m1 >>
rect 366 277 367 278 
<< m1 >>
rect 367 277 368 278 
<< m1 >>
rect 368 277 369 278 
<< m1 >>
rect 369 277 370 278 
<< m1 >>
rect 370 277 371 278 
<< m1 >>
rect 371 277 372 278 
<< m1 >>
rect 372 277 373 278 
<< m1 >>
rect 373 277 374 278 
<< m1 >>
rect 374 277 375 278 
<< m1 >>
rect 375 277 376 278 
<< m1 >>
rect 376 277 377 278 
<< m1 >>
rect 377 277 378 278 
<< m1 >>
rect 378 277 379 278 
<< m1 >>
rect 379 277 380 278 
<< m1 >>
rect 380 277 381 278 
<< m1 >>
rect 381 277 382 278 
<< m1 >>
rect 382 277 383 278 
<< m1 >>
rect 383 277 384 278 
<< m1 >>
rect 384 277 385 278 
<< m1 >>
rect 385 277 386 278 
<< m1 >>
rect 386 277 387 278 
<< m1 >>
rect 387 277 388 278 
<< m1 >>
rect 388 277 389 278 
<< m1 >>
rect 389 277 390 278 
<< m1 >>
rect 390 277 391 278 
<< m1 >>
rect 391 277 392 278 
<< m1 >>
rect 392 277 393 278 
<< m1 >>
rect 393 277 394 278 
<< m1 >>
rect 394 277 395 278 
<< m1 >>
rect 395 277 396 278 
<< m1 >>
rect 396 277 397 278 
<< m1 >>
rect 397 277 398 278 
<< m1 >>
rect 398 277 399 278 
<< m1 >>
rect 399 277 400 278 
<< m1 >>
rect 400 277 401 278 
<< m1 >>
rect 401 277 402 278 
<< m1 >>
rect 402 277 403 278 
<< m1 >>
rect 403 277 404 278 
<< m1 >>
rect 404 277 405 278 
<< m2 >>
rect 404 277 405 278 
<< m2c >>
rect 404 277 405 278 
<< m1 >>
rect 404 277 405 278 
<< m2 >>
rect 404 277 405 278 
<< m2 >>
rect 405 277 406 278 
<< m1 >>
rect 406 277 407 278 
<< m2 >>
rect 406 277 407 278 
<< m1 >>
rect 407 277 408 278 
<< m2 >>
rect 407 277 408 278 
<< m1 >>
rect 408 277 409 278 
<< m2 >>
rect 408 277 409 278 
<< m1 >>
rect 409 277 410 278 
<< m2 >>
rect 409 277 410 278 
<< m1 >>
rect 410 277 411 278 
<< m2 >>
rect 410 277 411 278 
<< m1 >>
rect 411 277 412 278 
<< m2 >>
rect 411 277 412 278 
<< m1 >>
rect 412 277 413 278 
<< m2 >>
rect 412 277 413 278 
<< m2 >>
rect 413 277 414 278 
<< m1 >>
rect 445 277 446 278 
<< m1 >>
rect 55 278 56 279 
<< m1 >>
rect 64 278 65 279 
<< m1 >>
rect 91 278 92 279 
<< m1 >>
rect 127 278 128 279 
<< m2 >>
rect 140 278 141 279 
<< m2 >>
rect 141 278 142 279 
<< m2 >>
rect 142 278 143 279 
<< m1 >>
rect 163 278 164 279 
<< m1 >>
rect 181 278 182 279 
<< m2 >>
rect 182 278 183 279 
<< m1 >>
rect 226 278 227 279 
<< m2 >>
rect 243 278 244 279 
<< m1 >>
rect 244 278 245 279 
<< m2 >>
rect 254 278 255 279 
<< m1 >>
rect 260 278 261 279 
<< m1 >>
rect 271 278 272 279 
<< m1 >>
rect 307 278 308 279 
<< m2 >>
rect 318 278 319 279 
<< m2 >>
rect 352 278 353 279 
<< m1 >>
rect 406 278 407 279 
<< m2 >>
rect 413 278 414 279 
<< m1 >>
rect 414 278 415 279 
<< m2 >>
rect 414 278 415 279 
<< m2c >>
rect 414 278 415 279 
<< m1 >>
rect 414 278 415 279 
<< m2 >>
rect 414 278 415 279 
<< m1 >>
rect 415 278 416 279 
<< m1 >>
rect 416 278 417 279 
<< m1 >>
rect 417 278 418 279 
<< m1 >>
rect 418 278 419 279 
<< m1 >>
rect 419 278 420 279 
<< m1 >>
rect 420 278 421 279 
<< m1 >>
rect 421 278 422 279 
<< m1 >>
rect 422 278 423 279 
<< m1 >>
rect 423 278 424 279 
<< m1 >>
rect 424 278 425 279 
<< m1 >>
rect 425 278 426 279 
<< m1 >>
rect 426 278 427 279 
<< m1 >>
rect 427 278 428 279 
<< m1 >>
rect 445 278 446 279 
<< m1 >>
rect 55 279 56 280 
<< m1 >>
rect 64 279 65 280 
<< m1 >>
rect 91 279 92 280 
<< m1 >>
rect 127 279 128 280 
<< m1 >>
rect 139 279 140 280 
<< m1 >>
rect 140 279 141 280 
<< m1 >>
rect 141 279 142 280 
<< m1 >>
rect 142 279 143 280 
<< m2 >>
rect 142 279 143 280 
<< m1 >>
rect 143 279 144 280 
<< m1 >>
rect 144 279 145 280 
<< m1 >>
rect 145 279 146 280 
<< m1 >>
rect 163 279 164 280 
<< m1 >>
rect 181 279 182 280 
<< m2 >>
rect 182 279 183 280 
<< m1 >>
rect 226 279 227 280 
<< m2 >>
rect 243 279 244 280 
<< m1 >>
rect 244 279 245 280 
<< m1 >>
rect 254 279 255 280 
<< m2 >>
rect 254 279 255 280 
<< m2c >>
rect 254 279 255 280 
<< m1 >>
rect 254 279 255 280 
<< m2 >>
rect 254 279 255 280 
<< m1 >>
rect 260 279 261 280 
<< m1 >>
rect 271 279 272 280 
<< m1 >>
rect 307 279 308 280 
<< m2 >>
rect 308 279 309 280 
<< m1 >>
rect 309 279 310 280 
<< m2 >>
rect 309 279 310 280 
<< m2c >>
rect 309 279 310 280 
<< m1 >>
rect 309 279 310 280 
<< m2 >>
rect 309 279 310 280 
<< m1 >>
rect 310 279 311 280 
<< m1 >>
rect 311 279 312 280 
<< m1 >>
rect 312 279 313 280 
<< m1 >>
rect 313 279 314 280 
<< m1 >>
rect 314 279 315 280 
<< m1 >>
rect 315 279 316 280 
<< m1 >>
rect 316 279 317 280 
<< m1 >>
rect 317 279 318 280 
<< m1 >>
rect 318 279 319 280 
<< m2 >>
rect 318 279 319 280 
<< m2c >>
rect 318 279 319 280 
<< m1 >>
rect 318 279 319 280 
<< m2 >>
rect 318 279 319 280 
<< m1 >>
rect 352 279 353 280 
<< m2 >>
rect 352 279 353 280 
<< m2c >>
rect 352 279 353 280 
<< m1 >>
rect 352 279 353 280 
<< m2 >>
rect 352 279 353 280 
<< m1 >>
rect 406 279 407 280 
<< m1 >>
rect 427 279 428 280 
<< m1 >>
rect 445 279 446 280 
<< m1 >>
rect 55 280 56 281 
<< m1 >>
rect 64 280 65 281 
<< m1 >>
rect 91 280 92 281 
<< m1 >>
rect 127 280 128 281 
<< m1 >>
rect 139 280 140 281 
<< m2 >>
rect 142 280 143 281 
<< m1 >>
rect 145 280 146 281 
<< m1 >>
rect 163 280 164 281 
<< m1 >>
rect 181 280 182 281 
<< m2 >>
rect 182 280 183 281 
<< m1 >>
rect 224 280 225 281 
<< m2 >>
rect 224 280 225 281 
<< m2c >>
rect 224 280 225 281 
<< m1 >>
rect 224 280 225 281 
<< m2 >>
rect 224 280 225 281 
<< m2 >>
rect 225 280 226 281 
<< m1 >>
rect 226 280 227 281 
<< m2 >>
rect 226 280 227 281 
<< m2 >>
rect 227 280 228 281 
<< m1 >>
rect 228 280 229 281 
<< m2 >>
rect 228 280 229 281 
<< m2c >>
rect 228 280 229 281 
<< m1 >>
rect 228 280 229 281 
<< m2 >>
rect 228 280 229 281 
<< m1 >>
rect 229 280 230 281 
<< m2 >>
rect 243 280 244 281 
<< m1 >>
rect 244 280 245 281 
<< m1 >>
rect 254 280 255 281 
<< m1 >>
rect 260 280 261 281 
<< m1 >>
rect 268 280 269 281 
<< m1 >>
rect 269 280 270 281 
<< m1 >>
rect 270 280 271 281 
<< m1 >>
rect 271 280 272 281 
<< m1 >>
rect 307 280 308 281 
<< m2 >>
rect 308 280 309 281 
<< m1 >>
rect 352 280 353 281 
<< m1 >>
rect 406 280 407 281 
<< m1 >>
rect 427 280 428 281 
<< m1 >>
rect 445 280 446 281 
<< m1 >>
rect 55 281 56 282 
<< m1 >>
rect 64 281 65 282 
<< m1 >>
rect 91 281 92 282 
<< m1 >>
rect 127 281 128 282 
<< m1 >>
rect 139 281 140 282 
<< m1 >>
rect 142 281 143 282 
<< m2 >>
rect 142 281 143 282 
<< m2c >>
rect 142 281 143 282 
<< m1 >>
rect 142 281 143 282 
<< m2 >>
rect 142 281 143 282 
<< m1 >>
rect 145 281 146 282 
<< m1 >>
rect 163 281 164 282 
<< m1 >>
rect 181 281 182 282 
<< m2 >>
rect 182 281 183 282 
<< m1 >>
rect 224 281 225 282 
<< m1 >>
rect 226 281 227 282 
<< m1 >>
rect 229 281 230 282 
<< m2 >>
rect 243 281 244 282 
<< m1 >>
rect 244 281 245 282 
<< m1 >>
rect 254 281 255 282 
<< m1 >>
rect 260 281 261 282 
<< m1 >>
rect 268 281 269 282 
<< m1 >>
rect 307 281 308 282 
<< m2 >>
rect 308 281 309 282 
<< m1 >>
rect 352 281 353 282 
<< m1 >>
rect 406 281 407 282 
<< m1 >>
rect 427 281 428 282 
<< m1 >>
rect 445 281 446 282 
<< pdiffusion >>
rect 12 282 13 283 
<< pdiffusion >>
rect 13 282 14 283 
<< pdiffusion >>
rect 14 282 15 283 
<< pdiffusion >>
rect 15 282 16 283 
<< pdiffusion >>
rect 16 282 17 283 
<< pdiffusion >>
rect 17 282 18 283 
<< pdiffusion >>
rect 30 282 31 283 
<< pdiffusion >>
rect 31 282 32 283 
<< pdiffusion >>
rect 32 282 33 283 
<< pdiffusion >>
rect 33 282 34 283 
<< pdiffusion >>
rect 34 282 35 283 
<< pdiffusion >>
rect 35 282 36 283 
<< pdiffusion >>
rect 48 282 49 283 
<< pdiffusion >>
rect 49 282 50 283 
<< pdiffusion >>
rect 50 282 51 283 
<< pdiffusion >>
rect 51 282 52 283 
<< pdiffusion >>
rect 52 282 53 283 
<< pdiffusion >>
rect 53 282 54 283 
<< m1 >>
rect 55 282 56 283 
<< m1 >>
rect 64 282 65 283 
<< pdiffusion >>
rect 66 282 67 283 
<< pdiffusion >>
rect 67 282 68 283 
<< pdiffusion >>
rect 68 282 69 283 
<< pdiffusion >>
rect 69 282 70 283 
<< pdiffusion >>
rect 70 282 71 283 
<< pdiffusion >>
rect 71 282 72 283 
<< pdiffusion >>
rect 84 282 85 283 
<< pdiffusion >>
rect 85 282 86 283 
<< pdiffusion >>
rect 86 282 87 283 
<< pdiffusion >>
rect 87 282 88 283 
<< pdiffusion >>
rect 88 282 89 283 
<< pdiffusion >>
rect 89 282 90 283 
<< m1 >>
rect 91 282 92 283 
<< pdiffusion >>
rect 102 282 103 283 
<< pdiffusion >>
rect 103 282 104 283 
<< pdiffusion >>
rect 104 282 105 283 
<< pdiffusion >>
rect 105 282 106 283 
<< pdiffusion >>
rect 106 282 107 283 
<< pdiffusion >>
rect 107 282 108 283 
<< pdiffusion >>
rect 120 282 121 283 
<< pdiffusion >>
rect 121 282 122 283 
<< pdiffusion >>
rect 122 282 123 283 
<< pdiffusion >>
rect 123 282 124 283 
<< pdiffusion >>
rect 124 282 125 283 
<< pdiffusion >>
rect 125 282 126 283 
<< m1 >>
rect 127 282 128 283 
<< pdiffusion >>
rect 138 282 139 283 
<< m1 >>
rect 139 282 140 283 
<< pdiffusion >>
rect 139 282 140 283 
<< pdiffusion >>
rect 140 282 141 283 
<< pdiffusion >>
rect 141 282 142 283 
<< m1 >>
rect 142 282 143 283 
<< pdiffusion >>
rect 142 282 143 283 
<< pdiffusion >>
rect 143 282 144 283 
<< m1 >>
rect 145 282 146 283 
<< pdiffusion >>
rect 156 282 157 283 
<< pdiffusion >>
rect 157 282 158 283 
<< pdiffusion >>
rect 158 282 159 283 
<< pdiffusion >>
rect 159 282 160 283 
<< pdiffusion >>
rect 160 282 161 283 
<< pdiffusion >>
rect 161 282 162 283 
<< m1 >>
rect 163 282 164 283 
<< pdiffusion >>
rect 174 282 175 283 
<< pdiffusion >>
rect 175 282 176 283 
<< pdiffusion >>
rect 176 282 177 283 
<< pdiffusion >>
rect 177 282 178 283 
<< pdiffusion >>
rect 178 282 179 283 
<< pdiffusion >>
rect 179 282 180 283 
<< m1 >>
rect 181 282 182 283 
<< m2 >>
rect 182 282 183 283 
<< pdiffusion >>
rect 192 282 193 283 
<< pdiffusion >>
rect 193 282 194 283 
<< pdiffusion >>
rect 194 282 195 283 
<< pdiffusion >>
rect 195 282 196 283 
<< pdiffusion >>
rect 196 282 197 283 
<< pdiffusion >>
rect 197 282 198 283 
<< pdiffusion >>
rect 210 282 211 283 
<< pdiffusion >>
rect 211 282 212 283 
<< pdiffusion >>
rect 212 282 213 283 
<< pdiffusion >>
rect 213 282 214 283 
<< pdiffusion >>
rect 214 282 215 283 
<< pdiffusion >>
rect 215 282 216 283 
<< m1 >>
rect 224 282 225 283 
<< m1 >>
rect 226 282 227 283 
<< pdiffusion >>
rect 228 282 229 283 
<< m1 >>
rect 229 282 230 283 
<< pdiffusion >>
rect 229 282 230 283 
<< pdiffusion >>
rect 230 282 231 283 
<< pdiffusion >>
rect 231 282 232 283 
<< pdiffusion >>
rect 232 282 233 283 
<< pdiffusion >>
rect 233 282 234 283 
<< m2 >>
rect 243 282 244 283 
<< m1 >>
rect 244 282 245 283 
<< pdiffusion >>
rect 246 282 247 283 
<< pdiffusion >>
rect 247 282 248 283 
<< pdiffusion >>
rect 248 282 249 283 
<< pdiffusion >>
rect 249 282 250 283 
<< pdiffusion >>
rect 250 282 251 283 
<< pdiffusion >>
rect 251 282 252 283 
<< m1 >>
rect 254 282 255 283 
<< m1 >>
rect 260 282 261 283 
<< pdiffusion >>
rect 264 282 265 283 
<< pdiffusion >>
rect 265 282 266 283 
<< pdiffusion >>
rect 266 282 267 283 
<< pdiffusion >>
rect 267 282 268 283 
<< m1 >>
rect 268 282 269 283 
<< pdiffusion >>
rect 268 282 269 283 
<< pdiffusion >>
rect 269 282 270 283 
<< pdiffusion >>
rect 300 282 301 283 
<< pdiffusion >>
rect 301 282 302 283 
<< pdiffusion >>
rect 302 282 303 283 
<< pdiffusion >>
rect 303 282 304 283 
<< pdiffusion >>
rect 304 282 305 283 
<< pdiffusion >>
rect 305 282 306 283 
<< m1 >>
rect 307 282 308 283 
<< m2 >>
rect 308 282 309 283 
<< pdiffusion >>
rect 318 282 319 283 
<< pdiffusion >>
rect 319 282 320 283 
<< pdiffusion >>
rect 320 282 321 283 
<< pdiffusion >>
rect 321 282 322 283 
<< pdiffusion >>
rect 322 282 323 283 
<< pdiffusion >>
rect 323 282 324 283 
<< pdiffusion >>
rect 336 282 337 283 
<< pdiffusion >>
rect 337 282 338 283 
<< pdiffusion >>
rect 338 282 339 283 
<< pdiffusion >>
rect 339 282 340 283 
<< pdiffusion >>
rect 340 282 341 283 
<< pdiffusion >>
rect 341 282 342 283 
<< m1 >>
rect 352 282 353 283 
<< pdiffusion >>
rect 354 282 355 283 
<< pdiffusion >>
rect 355 282 356 283 
<< pdiffusion >>
rect 356 282 357 283 
<< pdiffusion >>
rect 357 282 358 283 
<< pdiffusion >>
rect 358 282 359 283 
<< pdiffusion >>
rect 359 282 360 283 
<< pdiffusion >>
rect 372 282 373 283 
<< pdiffusion >>
rect 373 282 374 283 
<< pdiffusion >>
rect 374 282 375 283 
<< pdiffusion >>
rect 375 282 376 283 
<< pdiffusion >>
rect 376 282 377 283 
<< pdiffusion >>
rect 377 282 378 283 
<< pdiffusion >>
rect 390 282 391 283 
<< pdiffusion >>
rect 391 282 392 283 
<< pdiffusion >>
rect 392 282 393 283 
<< pdiffusion >>
rect 393 282 394 283 
<< pdiffusion >>
rect 394 282 395 283 
<< pdiffusion >>
rect 395 282 396 283 
<< m1 >>
rect 406 282 407 283 
<< pdiffusion >>
rect 408 282 409 283 
<< pdiffusion >>
rect 409 282 410 283 
<< pdiffusion >>
rect 410 282 411 283 
<< pdiffusion >>
rect 411 282 412 283 
<< pdiffusion >>
rect 412 282 413 283 
<< pdiffusion >>
rect 413 282 414 283 
<< pdiffusion >>
rect 426 282 427 283 
<< m1 >>
rect 427 282 428 283 
<< pdiffusion >>
rect 427 282 428 283 
<< pdiffusion >>
rect 428 282 429 283 
<< pdiffusion >>
rect 429 282 430 283 
<< pdiffusion >>
rect 430 282 431 283 
<< pdiffusion >>
rect 431 282 432 283 
<< pdiffusion >>
rect 444 282 445 283 
<< m1 >>
rect 445 282 446 283 
<< pdiffusion >>
rect 445 282 446 283 
<< pdiffusion >>
rect 446 282 447 283 
<< pdiffusion >>
rect 447 282 448 283 
<< pdiffusion >>
rect 448 282 449 283 
<< pdiffusion >>
rect 449 282 450 283 
<< pdiffusion >>
rect 12 283 13 284 
<< pdiffusion >>
rect 13 283 14 284 
<< pdiffusion >>
rect 14 283 15 284 
<< pdiffusion >>
rect 15 283 16 284 
<< pdiffusion >>
rect 16 283 17 284 
<< pdiffusion >>
rect 17 283 18 284 
<< pdiffusion >>
rect 30 283 31 284 
<< pdiffusion >>
rect 31 283 32 284 
<< pdiffusion >>
rect 32 283 33 284 
<< pdiffusion >>
rect 33 283 34 284 
<< pdiffusion >>
rect 34 283 35 284 
<< pdiffusion >>
rect 35 283 36 284 
<< pdiffusion >>
rect 48 283 49 284 
<< pdiffusion >>
rect 49 283 50 284 
<< pdiffusion >>
rect 50 283 51 284 
<< pdiffusion >>
rect 51 283 52 284 
<< pdiffusion >>
rect 52 283 53 284 
<< pdiffusion >>
rect 53 283 54 284 
<< m1 >>
rect 55 283 56 284 
<< m1 >>
rect 64 283 65 284 
<< pdiffusion >>
rect 66 283 67 284 
<< pdiffusion >>
rect 67 283 68 284 
<< pdiffusion >>
rect 68 283 69 284 
<< pdiffusion >>
rect 69 283 70 284 
<< pdiffusion >>
rect 70 283 71 284 
<< pdiffusion >>
rect 71 283 72 284 
<< pdiffusion >>
rect 84 283 85 284 
<< pdiffusion >>
rect 85 283 86 284 
<< pdiffusion >>
rect 86 283 87 284 
<< pdiffusion >>
rect 87 283 88 284 
<< pdiffusion >>
rect 88 283 89 284 
<< pdiffusion >>
rect 89 283 90 284 
<< m1 >>
rect 91 283 92 284 
<< pdiffusion >>
rect 102 283 103 284 
<< pdiffusion >>
rect 103 283 104 284 
<< pdiffusion >>
rect 104 283 105 284 
<< pdiffusion >>
rect 105 283 106 284 
<< pdiffusion >>
rect 106 283 107 284 
<< pdiffusion >>
rect 107 283 108 284 
<< pdiffusion >>
rect 120 283 121 284 
<< pdiffusion >>
rect 121 283 122 284 
<< pdiffusion >>
rect 122 283 123 284 
<< pdiffusion >>
rect 123 283 124 284 
<< pdiffusion >>
rect 124 283 125 284 
<< pdiffusion >>
rect 125 283 126 284 
<< m1 >>
rect 127 283 128 284 
<< pdiffusion >>
rect 138 283 139 284 
<< pdiffusion >>
rect 139 283 140 284 
<< pdiffusion >>
rect 140 283 141 284 
<< pdiffusion >>
rect 141 283 142 284 
<< pdiffusion >>
rect 142 283 143 284 
<< pdiffusion >>
rect 143 283 144 284 
<< m1 >>
rect 145 283 146 284 
<< pdiffusion >>
rect 156 283 157 284 
<< pdiffusion >>
rect 157 283 158 284 
<< pdiffusion >>
rect 158 283 159 284 
<< pdiffusion >>
rect 159 283 160 284 
<< pdiffusion >>
rect 160 283 161 284 
<< pdiffusion >>
rect 161 283 162 284 
<< m1 >>
rect 163 283 164 284 
<< pdiffusion >>
rect 174 283 175 284 
<< pdiffusion >>
rect 175 283 176 284 
<< pdiffusion >>
rect 176 283 177 284 
<< pdiffusion >>
rect 177 283 178 284 
<< pdiffusion >>
rect 178 283 179 284 
<< pdiffusion >>
rect 179 283 180 284 
<< m1 >>
rect 181 283 182 284 
<< m2 >>
rect 182 283 183 284 
<< pdiffusion >>
rect 192 283 193 284 
<< pdiffusion >>
rect 193 283 194 284 
<< pdiffusion >>
rect 194 283 195 284 
<< pdiffusion >>
rect 195 283 196 284 
<< pdiffusion >>
rect 196 283 197 284 
<< pdiffusion >>
rect 197 283 198 284 
<< pdiffusion >>
rect 210 283 211 284 
<< pdiffusion >>
rect 211 283 212 284 
<< pdiffusion >>
rect 212 283 213 284 
<< pdiffusion >>
rect 213 283 214 284 
<< pdiffusion >>
rect 214 283 215 284 
<< pdiffusion >>
rect 215 283 216 284 
<< m1 >>
rect 224 283 225 284 
<< m1 >>
rect 226 283 227 284 
<< pdiffusion >>
rect 228 283 229 284 
<< pdiffusion >>
rect 229 283 230 284 
<< pdiffusion >>
rect 230 283 231 284 
<< pdiffusion >>
rect 231 283 232 284 
<< pdiffusion >>
rect 232 283 233 284 
<< pdiffusion >>
rect 233 283 234 284 
<< m2 >>
rect 243 283 244 284 
<< m1 >>
rect 244 283 245 284 
<< pdiffusion >>
rect 246 283 247 284 
<< pdiffusion >>
rect 247 283 248 284 
<< pdiffusion >>
rect 248 283 249 284 
<< pdiffusion >>
rect 249 283 250 284 
<< pdiffusion >>
rect 250 283 251 284 
<< pdiffusion >>
rect 251 283 252 284 
<< m1 >>
rect 254 283 255 284 
<< m1 >>
rect 260 283 261 284 
<< pdiffusion >>
rect 264 283 265 284 
<< pdiffusion >>
rect 265 283 266 284 
<< pdiffusion >>
rect 266 283 267 284 
<< pdiffusion >>
rect 267 283 268 284 
<< pdiffusion >>
rect 268 283 269 284 
<< pdiffusion >>
rect 269 283 270 284 
<< pdiffusion >>
rect 300 283 301 284 
<< pdiffusion >>
rect 301 283 302 284 
<< pdiffusion >>
rect 302 283 303 284 
<< pdiffusion >>
rect 303 283 304 284 
<< pdiffusion >>
rect 304 283 305 284 
<< pdiffusion >>
rect 305 283 306 284 
<< m1 >>
rect 307 283 308 284 
<< m2 >>
rect 308 283 309 284 
<< pdiffusion >>
rect 318 283 319 284 
<< pdiffusion >>
rect 319 283 320 284 
<< pdiffusion >>
rect 320 283 321 284 
<< pdiffusion >>
rect 321 283 322 284 
<< pdiffusion >>
rect 322 283 323 284 
<< pdiffusion >>
rect 323 283 324 284 
<< pdiffusion >>
rect 336 283 337 284 
<< pdiffusion >>
rect 337 283 338 284 
<< pdiffusion >>
rect 338 283 339 284 
<< pdiffusion >>
rect 339 283 340 284 
<< pdiffusion >>
rect 340 283 341 284 
<< pdiffusion >>
rect 341 283 342 284 
<< m1 >>
rect 352 283 353 284 
<< pdiffusion >>
rect 354 283 355 284 
<< pdiffusion >>
rect 355 283 356 284 
<< pdiffusion >>
rect 356 283 357 284 
<< pdiffusion >>
rect 357 283 358 284 
<< pdiffusion >>
rect 358 283 359 284 
<< pdiffusion >>
rect 359 283 360 284 
<< pdiffusion >>
rect 372 283 373 284 
<< pdiffusion >>
rect 373 283 374 284 
<< pdiffusion >>
rect 374 283 375 284 
<< pdiffusion >>
rect 375 283 376 284 
<< pdiffusion >>
rect 376 283 377 284 
<< pdiffusion >>
rect 377 283 378 284 
<< pdiffusion >>
rect 390 283 391 284 
<< pdiffusion >>
rect 391 283 392 284 
<< pdiffusion >>
rect 392 283 393 284 
<< pdiffusion >>
rect 393 283 394 284 
<< pdiffusion >>
rect 394 283 395 284 
<< pdiffusion >>
rect 395 283 396 284 
<< m1 >>
rect 406 283 407 284 
<< pdiffusion >>
rect 408 283 409 284 
<< pdiffusion >>
rect 409 283 410 284 
<< pdiffusion >>
rect 410 283 411 284 
<< pdiffusion >>
rect 411 283 412 284 
<< pdiffusion >>
rect 412 283 413 284 
<< pdiffusion >>
rect 413 283 414 284 
<< pdiffusion >>
rect 426 283 427 284 
<< pdiffusion >>
rect 427 283 428 284 
<< pdiffusion >>
rect 428 283 429 284 
<< pdiffusion >>
rect 429 283 430 284 
<< pdiffusion >>
rect 430 283 431 284 
<< pdiffusion >>
rect 431 283 432 284 
<< pdiffusion >>
rect 444 283 445 284 
<< pdiffusion >>
rect 445 283 446 284 
<< pdiffusion >>
rect 446 283 447 284 
<< pdiffusion >>
rect 447 283 448 284 
<< pdiffusion >>
rect 448 283 449 284 
<< pdiffusion >>
rect 449 283 450 284 
<< pdiffusion >>
rect 12 284 13 285 
<< pdiffusion >>
rect 13 284 14 285 
<< pdiffusion >>
rect 14 284 15 285 
<< pdiffusion >>
rect 15 284 16 285 
<< pdiffusion >>
rect 16 284 17 285 
<< pdiffusion >>
rect 17 284 18 285 
<< pdiffusion >>
rect 30 284 31 285 
<< pdiffusion >>
rect 31 284 32 285 
<< pdiffusion >>
rect 32 284 33 285 
<< pdiffusion >>
rect 33 284 34 285 
<< pdiffusion >>
rect 34 284 35 285 
<< pdiffusion >>
rect 35 284 36 285 
<< pdiffusion >>
rect 48 284 49 285 
<< pdiffusion >>
rect 49 284 50 285 
<< pdiffusion >>
rect 50 284 51 285 
<< pdiffusion >>
rect 51 284 52 285 
<< pdiffusion >>
rect 52 284 53 285 
<< pdiffusion >>
rect 53 284 54 285 
<< m1 >>
rect 55 284 56 285 
<< m1 >>
rect 64 284 65 285 
<< pdiffusion >>
rect 66 284 67 285 
<< pdiffusion >>
rect 67 284 68 285 
<< pdiffusion >>
rect 68 284 69 285 
<< pdiffusion >>
rect 69 284 70 285 
<< pdiffusion >>
rect 70 284 71 285 
<< pdiffusion >>
rect 71 284 72 285 
<< pdiffusion >>
rect 84 284 85 285 
<< pdiffusion >>
rect 85 284 86 285 
<< pdiffusion >>
rect 86 284 87 285 
<< pdiffusion >>
rect 87 284 88 285 
<< pdiffusion >>
rect 88 284 89 285 
<< pdiffusion >>
rect 89 284 90 285 
<< m1 >>
rect 91 284 92 285 
<< pdiffusion >>
rect 102 284 103 285 
<< pdiffusion >>
rect 103 284 104 285 
<< pdiffusion >>
rect 104 284 105 285 
<< pdiffusion >>
rect 105 284 106 285 
<< pdiffusion >>
rect 106 284 107 285 
<< pdiffusion >>
rect 107 284 108 285 
<< pdiffusion >>
rect 120 284 121 285 
<< pdiffusion >>
rect 121 284 122 285 
<< pdiffusion >>
rect 122 284 123 285 
<< pdiffusion >>
rect 123 284 124 285 
<< pdiffusion >>
rect 124 284 125 285 
<< pdiffusion >>
rect 125 284 126 285 
<< m1 >>
rect 127 284 128 285 
<< pdiffusion >>
rect 138 284 139 285 
<< pdiffusion >>
rect 139 284 140 285 
<< pdiffusion >>
rect 140 284 141 285 
<< pdiffusion >>
rect 141 284 142 285 
<< pdiffusion >>
rect 142 284 143 285 
<< pdiffusion >>
rect 143 284 144 285 
<< m1 >>
rect 145 284 146 285 
<< pdiffusion >>
rect 156 284 157 285 
<< pdiffusion >>
rect 157 284 158 285 
<< pdiffusion >>
rect 158 284 159 285 
<< pdiffusion >>
rect 159 284 160 285 
<< pdiffusion >>
rect 160 284 161 285 
<< pdiffusion >>
rect 161 284 162 285 
<< m1 >>
rect 163 284 164 285 
<< pdiffusion >>
rect 174 284 175 285 
<< pdiffusion >>
rect 175 284 176 285 
<< pdiffusion >>
rect 176 284 177 285 
<< pdiffusion >>
rect 177 284 178 285 
<< pdiffusion >>
rect 178 284 179 285 
<< pdiffusion >>
rect 179 284 180 285 
<< m1 >>
rect 181 284 182 285 
<< m2 >>
rect 182 284 183 285 
<< pdiffusion >>
rect 192 284 193 285 
<< pdiffusion >>
rect 193 284 194 285 
<< pdiffusion >>
rect 194 284 195 285 
<< pdiffusion >>
rect 195 284 196 285 
<< pdiffusion >>
rect 196 284 197 285 
<< pdiffusion >>
rect 197 284 198 285 
<< pdiffusion >>
rect 210 284 211 285 
<< pdiffusion >>
rect 211 284 212 285 
<< pdiffusion >>
rect 212 284 213 285 
<< pdiffusion >>
rect 213 284 214 285 
<< pdiffusion >>
rect 214 284 215 285 
<< pdiffusion >>
rect 215 284 216 285 
<< m1 >>
rect 224 284 225 285 
<< m1 >>
rect 226 284 227 285 
<< pdiffusion >>
rect 228 284 229 285 
<< pdiffusion >>
rect 229 284 230 285 
<< pdiffusion >>
rect 230 284 231 285 
<< pdiffusion >>
rect 231 284 232 285 
<< pdiffusion >>
rect 232 284 233 285 
<< pdiffusion >>
rect 233 284 234 285 
<< m2 >>
rect 243 284 244 285 
<< m1 >>
rect 244 284 245 285 
<< pdiffusion >>
rect 246 284 247 285 
<< pdiffusion >>
rect 247 284 248 285 
<< pdiffusion >>
rect 248 284 249 285 
<< pdiffusion >>
rect 249 284 250 285 
<< pdiffusion >>
rect 250 284 251 285 
<< pdiffusion >>
rect 251 284 252 285 
<< m1 >>
rect 254 284 255 285 
<< m1 >>
rect 260 284 261 285 
<< pdiffusion >>
rect 264 284 265 285 
<< pdiffusion >>
rect 265 284 266 285 
<< pdiffusion >>
rect 266 284 267 285 
<< pdiffusion >>
rect 267 284 268 285 
<< pdiffusion >>
rect 268 284 269 285 
<< pdiffusion >>
rect 269 284 270 285 
<< pdiffusion >>
rect 300 284 301 285 
<< pdiffusion >>
rect 301 284 302 285 
<< pdiffusion >>
rect 302 284 303 285 
<< pdiffusion >>
rect 303 284 304 285 
<< pdiffusion >>
rect 304 284 305 285 
<< pdiffusion >>
rect 305 284 306 285 
<< m1 >>
rect 307 284 308 285 
<< m2 >>
rect 308 284 309 285 
<< pdiffusion >>
rect 318 284 319 285 
<< pdiffusion >>
rect 319 284 320 285 
<< pdiffusion >>
rect 320 284 321 285 
<< pdiffusion >>
rect 321 284 322 285 
<< pdiffusion >>
rect 322 284 323 285 
<< pdiffusion >>
rect 323 284 324 285 
<< pdiffusion >>
rect 336 284 337 285 
<< pdiffusion >>
rect 337 284 338 285 
<< pdiffusion >>
rect 338 284 339 285 
<< pdiffusion >>
rect 339 284 340 285 
<< pdiffusion >>
rect 340 284 341 285 
<< pdiffusion >>
rect 341 284 342 285 
<< m1 >>
rect 352 284 353 285 
<< pdiffusion >>
rect 354 284 355 285 
<< pdiffusion >>
rect 355 284 356 285 
<< pdiffusion >>
rect 356 284 357 285 
<< pdiffusion >>
rect 357 284 358 285 
<< pdiffusion >>
rect 358 284 359 285 
<< pdiffusion >>
rect 359 284 360 285 
<< pdiffusion >>
rect 372 284 373 285 
<< pdiffusion >>
rect 373 284 374 285 
<< pdiffusion >>
rect 374 284 375 285 
<< pdiffusion >>
rect 375 284 376 285 
<< pdiffusion >>
rect 376 284 377 285 
<< pdiffusion >>
rect 377 284 378 285 
<< pdiffusion >>
rect 390 284 391 285 
<< pdiffusion >>
rect 391 284 392 285 
<< pdiffusion >>
rect 392 284 393 285 
<< pdiffusion >>
rect 393 284 394 285 
<< pdiffusion >>
rect 394 284 395 285 
<< pdiffusion >>
rect 395 284 396 285 
<< m1 >>
rect 406 284 407 285 
<< pdiffusion >>
rect 408 284 409 285 
<< pdiffusion >>
rect 409 284 410 285 
<< pdiffusion >>
rect 410 284 411 285 
<< pdiffusion >>
rect 411 284 412 285 
<< pdiffusion >>
rect 412 284 413 285 
<< pdiffusion >>
rect 413 284 414 285 
<< pdiffusion >>
rect 426 284 427 285 
<< pdiffusion >>
rect 427 284 428 285 
<< pdiffusion >>
rect 428 284 429 285 
<< pdiffusion >>
rect 429 284 430 285 
<< pdiffusion >>
rect 430 284 431 285 
<< pdiffusion >>
rect 431 284 432 285 
<< pdiffusion >>
rect 444 284 445 285 
<< pdiffusion >>
rect 445 284 446 285 
<< pdiffusion >>
rect 446 284 447 285 
<< pdiffusion >>
rect 447 284 448 285 
<< pdiffusion >>
rect 448 284 449 285 
<< pdiffusion >>
rect 449 284 450 285 
<< pdiffusion >>
rect 12 285 13 286 
<< pdiffusion >>
rect 13 285 14 286 
<< pdiffusion >>
rect 14 285 15 286 
<< pdiffusion >>
rect 15 285 16 286 
<< pdiffusion >>
rect 16 285 17 286 
<< pdiffusion >>
rect 17 285 18 286 
<< pdiffusion >>
rect 30 285 31 286 
<< pdiffusion >>
rect 31 285 32 286 
<< pdiffusion >>
rect 32 285 33 286 
<< pdiffusion >>
rect 33 285 34 286 
<< pdiffusion >>
rect 34 285 35 286 
<< pdiffusion >>
rect 35 285 36 286 
<< pdiffusion >>
rect 48 285 49 286 
<< pdiffusion >>
rect 49 285 50 286 
<< pdiffusion >>
rect 50 285 51 286 
<< pdiffusion >>
rect 51 285 52 286 
<< pdiffusion >>
rect 52 285 53 286 
<< pdiffusion >>
rect 53 285 54 286 
<< m1 >>
rect 55 285 56 286 
<< m1 >>
rect 64 285 65 286 
<< pdiffusion >>
rect 66 285 67 286 
<< pdiffusion >>
rect 67 285 68 286 
<< pdiffusion >>
rect 68 285 69 286 
<< pdiffusion >>
rect 69 285 70 286 
<< pdiffusion >>
rect 70 285 71 286 
<< pdiffusion >>
rect 71 285 72 286 
<< pdiffusion >>
rect 84 285 85 286 
<< pdiffusion >>
rect 85 285 86 286 
<< pdiffusion >>
rect 86 285 87 286 
<< pdiffusion >>
rect 87 285 88 286 
<< pdiffusion >>
rect 88 285 89 286 
<< pdiffusion >>
rect 89 285 90 286 
<< m1 >>
rect 91 285 92 286 
<< pdiffusion >>
rect 102 285 103 286 
<< pdiffusion >>
rect 103 285 104 286 
<< pdiffusion >>
rect 104 285 105 286 
<< pdiffusion >>
rect 105 285 106 286 
<< pdiffusion >>
rect 106 285 107 286 
<< pdiffusion >>
rect 107 285 108 286 
<< pdiffusion >>
rect 120 285 121 286 
<< pdiffusion >>
rect 121 285 122 286 
<< pdiffusion >>
rect 122 285 123 286 
<< pdiffusion >>
rect 123 285 124 286 
<< pdiffusion >>
rect 124 285 125 286 
<< pdiffusion >>
rect 125 285 126 286 
<< m1 >>
rect 127 285 128 286 
<< pdiffusion >>
rect 138 285 139 286 
<< pdiffusion >>
rect 139 285 140 286 
<< pdiffusion >>
rect 140 285 141 286 
<< pdiffusion >>
rect 141 285 142 286 
<< pdiffusion >>
rect 142 285 143 286 
<< pdiffusion >>
rect 143 285 144 286 
<< m1 >>
rect 145 285 146 286 
<< pdiffusion >>
rect 156 285 157 286 
<< pdiffusion >>
rect 157 285 158 286 
<< pdiffusion >>
rect 158 285 159 286 
<< pdiffusion >>
rect 159 285 160 286 
<< pdiffusion >>
rect 160 285 161 286 
<< pdiffusion >>
rect 161 285 162 286 
<< m1 >>
rect 163 285 164 286 
<< pdiffusion >>
rect 174 285 175 286 
<< pdiffusion >>
rect 175 285 176 286 
<< pdiffusion >>
rect 176 285 177 286 
<< pdiffusion >>
rect 177 285 178 286 
<< pdiffusion >>
rect 178 285 179 286 
<< pdiffusion >>
rect 179 285 180 286 
<< m1 >>
rect 181 285 182 286 
<< m2 >>
rect 182 285 183 286 
<< pdiffusion >>
rect 192 285 193 286 
<< pdiffusion >>
rect 193 285 194 286 
<< pdiffusion >>
rect 194 285 195 286 
<< pdiffusion >>
rect 195 285 196 286 
<< pdiffusion >>
rect 196 285 197 286 
<< pdiffusion >>
rect 197 285 198 286 
<< pdiffusion >>
rect 210 285 211 286 
<< pdiffusion >>
rect 211 285 212 286 
<< pdiffusion >>
rect 212 285 213 286 
<< pdiffusion >>
rect 213 285 214 286 
<< pdiffusion >>
rect 214 285 215 286 
<< pdiffusion >>
rect 215 285 216 286 
<< m1 >>
rect 224 285 225 286 
<< m1 >>
rect 226 285 227 286 
<< pdiffusion >>
rect 228 285 229 286 
<< pdiffusion >>
rect 229 285 230 286 
<< pdiffusion >>
rect 230 285 231 286 
<< pdiffusion >>
rect 231 285 232 286 
<< pdiffusion >>
rect 232 285 233 286 
<< pdiffusion >>
rect 233 285 234 286 
<< m2 >>
rect 243 285 244 286 
<< m1 >>
rect 244 285 245 286 
<< pdiffusion >>
rect 246 285 247 286 
<< pdiffusion >>
rect 247 285 248 286 
<< pdiffusion >>
rect 248 285 249 286 
<< pdiffusion >>
rect 249 285 250 286 
<< pdiffusion >>
rect 250 285 251 286 
<< pdiffusion >>
rect 251 285 252 286 
<< m1 >>
rect 254 285 255 286 
<< m1 >>
rect 260 285 261 286 
<< pdiffusion >>
rect 264 285 265 286 
<< pdiffusion >>
rect 265 285 266 286 
<< pdiffusion >>
rect 266 285 267 286 
<< pdiffusion >>
rect 267 285 268 286 
<< pdiffusion >>
rect 268 285 269 286 
<< pdiffusion >>
rect 269 285 270 286 
<< pdiffusion >>
rect 300 285 301 286 
<< pdiffusion >>
rect 301 285 302 286 
<< pdiffusion >>
rect 302 285 303 286 
<< pdiffusion >>
rect 303 285 304 286 
<< pdiffusion >>
rect 304 285 305 286 
<< pdiffusion >>
rect 305 285 306 286 
<< m1 >>
rect 307 285 308 286 
<< m2 >>
rect 308 285 309 286 
<< pdiffusion >>
rect 318 285 319 286 
<< pdiffusion >>
rect 319 285 320 286 
<< pdiffusion >>
rect 320 285 321 286 
<< pdiffusion >>
rect 321 285 322 286 
<< pdiffusion >>
rect 322 285 323 286 
<< pdiffusion >>
rect 323 285 324 286 
<< pdiffusion >>
rect 336 285 337 286 
<< pdiffusion >>
rect 337 285 338 286 
<< pdiffusion >>
rect 338 285 339 286 
<< pdiffusion >>
rect 339 285 340 286 
<< pdiffusion >>
rect 340 285 341 286 
<< pdiffusion >>
rect 341 285 342 286 
<< m1 >>
rect 352 285 353 286 
<< pdiffusion >>
rect 354 285 355 286 
<< pdiffusion >>
rect 355 285 356 286 
<< pdiffusion >>
rect 356 285 357 286 
<< pdiffusion >>
rect 357 285 358 286 
<< pdiffusion >>
rect 358 285 359 286 
<< pdiffusion >>
rect 359 285 360 286 
<< pdiffusion >>
rect 372 285 373 286 
<< pdiffusion >>
rect 373 285 374 286 
<< pdiffusion >>
rect 374 285 375 286 
<< pdiffusion >>
rect 375 285 376 286 
<< pdiffusion >>
rect 376 285 377 286 
<< pdiffusion >>
rect 377 285 378 286 
<< pdiffusion >>
rect 390 285 391 286 
<< pdiffusion >>
rect 391 285 392 286 
<< pdiffusion >>
rect 392 285 393 286 
<< pdiffusion >>
rect 393 285 394 286 
<< pdiffusion >>
rect 394 285 395 286 
<< pdiffusion >>
rect 395 285 396 286 
<< m1 >>
rect 406 285 407 286 
<< pdiffusion >>
rect 408 285 409 286 
<< pdiffusion >>
rect 409 285 410 286 
<< pdiffusion >>
rect 410 285 411 286 
<< pdiffusion >>
rect 411 285 412 286 
<< pdiffusion >>
rect 412 285 413 286 
<< pdiffusion >>
rect 413 285 414 286 
<< pdiffusion >>
rect 426 285 427 286 
<< pdiffusion >>
rect 427 285 428 286 
<< pdiffusion >>
rect 428 285 429 286 
<< pdiffusion >>
rect 429 285 430 286 
<< pdiffusion >>
rect 430 285 431 286 
<< pdiffusion >>
rect 431 285 432 286 
<< pdiffusion >>
rect 444 285 445 286 
<< pdiffusion >>
rect 445 285 446 286 
<< pdiffusion >>
rect 446 285 447 286 
<< pdiffusion >>
rect 447 285 448 286 
<< pdiffusion >>
rect 448 285 449 286 
<< pdiffusion >>
rect 449 285 450 286 
<< pdiffusion >>
rect 12 286 13 287 
<< pdiffusion >>
rect 13 286 14 287 
<< pdiffusion >>
rect 14 286 15 287 
<< pdiffusion >>
rect 15 286 16 287 
<< pdiffusion >>
rect 16 286 17 287 
<< pdiffusion >>
rect 17 286 18 287 
<< pdiffusion >>
rect 30 286 31 287 
<< pdiffusion >>
rect 31 286 32 287 
<< pdiffusion >>
rect 32 286 33 287 
<< pdiffusion >>
rect 33 286 34 287 
<< pdiffusion >>
rect 34 286 35 287 
<< pdiffusion >>
rect 35 286 36 287 
<< pdiffusion >>
rect 48 286 49 287 
<< pdiffusion >>
rect 49 286 50 287 
<< pdiffusion >>
rect 50 286 51 287 
<< pdiffusion >>
rect 51 286 52 287 
<< pdiffusion >>
rect 52 286 53 287 
<< pdiffusion >>
rect 53 286 54 287 
<< m1 >>
rect 55 286 56 287 
<< m1 >>
rect 64 286 65 287 
<< pdiffusion >>
rect 66 286 67 287 
<< pdiffusion >>
rect 67 286 68 287 
<< pdiffusion >>
rect 68 286 69 287 
<< pdiffusion >>
rect 69 286 70 287 
<< pdiffusion >>
rect 70 286 71 287 
<< pdiffusion >>
rect 71 286 72 287 
<< pdiffusion >>
rect 84 286 85 287 
<< pdiffusion >>
rect 85 286 86 287 
<< pdiffusion >>
rect 86 286 87 287 
<< pdiffusion >>
rect 87 286 88 287 
<< pdiffusion >>
rect 88 286 89 287 
<< pdiffusion >>
rect 89 286 90 287 
<< m1 >>
rect 91 286 92 287 
<< pdiffusion >>
rect 102 286 103 287 
<< pdiffusion >>
rect 103 286 104 287 
<< pdiffusion >>
rect 104 286 105 287 
<< pdiffusion >>
rect 105 286 106 287 
<< pdiffusion >>
rect 106 286 107 287 
<< pdiffusion >>
rect 107 286 108 287 
<< pdiffusion >>
rect 120 286 121 287 
<< pdiffusion >>
rect 121 286 122 287 
<< pdiffusion >>
rect 122 286 123 287 
<< pdiffusion >>
rect 123 286 124 287 
<< pdiffusion >>
rect 124 286 125 287 
<< pdiffusion >>
rect 125 286 126 287 
<< m1 >>
rect 127 286 128 287 
<< pdiffusion >>
rect 138 286 139 287 
<< pdiffusion >>
rect 139 286 140 287 
<< pdiffusion >>
rect 140 286 141 287 
<< pdiffusion >>
rect 141 286 142 287 
<< pdiffusion >>
rect 142 286 143 287 
<< pdiffusion >>
rect 143 286 144 287 
<< m1 >>
rect 145 286 146 287 
<< pdiffusion >>
rect 156 286 157 287 
<< pdiffusion >>
rect 157 286 158 287 
<< pdiffusion >>
rect 158 286 159 287 
<< pdiffusion >>
rect 159 286 160 287 
<< pdiffusion >>
rect 160 286 161 287 
<< pdiffusion >>
rect 161 286 162 287 
<< m1 >>
rect 163 286 164 287 
<< pdiffusion >>
rect 174 286 175 287 
<< pdiffusion >>
rect 175 286 176 287 
<< pdiffusion >>
rect 176 286 177 287 
<< pdiffusion >>
rect 177 286 178 287 
<< pdiffusion >>
rect 178 286 179 287 
<< pdiffusion >>
rect 179 286 180 287 
<< m1 >>
rect 181 286 182 287 
<< m2 >>
rect 182 286 183 287 
<< pdiffusion >>
rect 192 286 193 287 
<< pdiffusion >>
rect 193 286 194 287 
<< pdiffusion >>
rect 194 286 195 287 
<< pdiffusion >>
rect 195 286 196 287 
<< pdiffusion >>
rect 196 286 197 287 
<< pdiffusion >>
rect 197 286 198 287 
<< pdiffusion >>
rect 210 286 211 287 
<< pdiffusion >>
rect 211 286 212 287 
<< pdiffusion >>
rect 212 286 213 287 
<< pdiffusion >>
rect 213 286 214 287 
<< pdiffusion >>
rect 214 286 215 287 
<< pdiffusion >>
rect 215 286 216 287 
<< m1 >>
rect 224 286 225 287 
<< m1 >>
rect 226 286 227 287 
<< pdiffusion >>
rect 228 286 229 287 
<< pdiffusion >>
rect 229 286 230 287 
<< pdiffusion >>
rect 230 286 231 287 
<< pdiffusion >>
rect 231 286 232 287 
<< pdiffusion >>
rect 232 286 233 287 
<< pdiffusion >>
rect 233 286 234 287 
<< m2 >>
rect 243 286 244 287 
<< m1 >>
rect 244 286 245 287 
<< pdiffusion >>
rect 246 286 247 287 
<< pdiffusion >>
rect 247 286 248 287 
<< pdiffusion >>
rect 248 286 249 287 
<< pdiffusion >>
rect 249 286 250 287 
<< pdiffusion >>
rect 250 286 251 287 
<< pdiffusion >>
rect 251 286 252 287 
<< m1 >>
rect 254 286 255 287 
<< m1 >>
rect 260 286 261 287 
<< pdiffusion >>
rect 264 286 265 287 
<< pdiffusion >>
rect 265 286 266 287 
<< pdiffusion >>
rect 266 286 267 287 
<< pdiffusion >>
rect 267 286 268 287 
<< pdiffusion >>
rect 268 286 269 287 
<< pdiffusion >>
rect 269 286 270 287 
<< pdiffusion >>
rect 300 286 301 287 
<< pdiffusion >>
rect 301 286 302 287 
<< pdiffusion >>
rect 302 286 303 287 
<< pdiffusion >>
rect 303 286 304 287 
<< pdiffusion >>
rect 304 286 305 287 
<< pdiffusion >>
rect 305 286 306 287 
<< m1 >>
rect 307 286 308 287 
<< m2 >>
rect 308 286 309 287 
<< pdiffusion >>
rect 318 286 319 287 
<< pdiffusion >>
rect 319 286 320 287 
<< pdiffusion >>
rect 320 286 321 287 
<< pdiffusion >>
rect 321 286 322 287 
<< pdiffusion >>
rect 322 286 323 287 
<< pdiffusion >>
rect 323 286 324 287 
<< pdiffusion >>
rect 336 286 337 287 
<< pdiffusion >>
rect 337 286 338 287 
<< pdiffusion >>
rect 338 286 339 287 
<< pdiffusion >>
rect 339 286 340 287 
<< pdiffusion >>
rect 340 286 341 287 
<< pdiffusion >>
rect 341 286 342 287 
<< m1 >>
rect 352 286 353 287 
<< pdiffusion >>
rect 354 286 355 287 
<< pdiffusion >>
rect 355 286 356 287 
<< pdiffusion >>
rect 356 286 357 287 
<< pdiffusion >>
rect 357 286 358 287 
<< pdiffusion >>
rect 358 286 359 287 
<< pdiffusion >>
rect 359 286 360 287 
<< pdiffusion >>
rect 372 286 373 287 
<< pdiffusion >>
rect 373 286 374 287 
<< pdiffusion >>
rect 374 286 375 287 
<< pdiffusion >>
rect 375 286 376 287 
<< pdiffusion >>
rect 376 286 377 287 
<< pdiffusion >>
rect 377 286 378 287 
<< pdiffusion >>
rect 390 286 391 287 
<< pdiffusion >>
rect 391 286 392 287 
<< pdiffusion >>
rect 392 286 393 287 
<< pdiffusion >>
rect 393 286 394 287 
<< pdiffusion >>
rect 394 286 395 287 
<< pdiffusion >>
rect 395 286 396 287 
<< m1 >>
rect 406 286 407 287 
<< pdiffusion >>
rect 408 286 409 287 
<< pdiffusion >>
rect 409 286 410 287 
<< pdiffusion >>
rect 410 286 411 287 
<< pdiffusion >>
rect 411 286 412 287 
<< pdiffusion >>
rect 412 286 413 287 
<< pdiffusion >>
rect 413 286 414 287 
<< pdiffusion >>
rect 426 286 427 287 
<< pdiffusion >>
rect 427 286 428 287 
<< pdiffusion >>
rect 428 286 429 287 
<< pdiffusion >>
rect 429 286 430 287 
<< pdiffusion >>
rect 430 286 431 287 
<< pdiffusion >>
rect 431 286 432 287 
<< pdiffusion >>
rect 444 286 445 287 
<< pdiffusion >>
rect 445 286 446 287 
<< pdiffusion >>
rect 446 286 447 287 
<< pdiffusion >>
rect 447 286 448 287 
<< pdiffusion >>
rect 448 286 449 287 
<< pdiffusion >>
rect 449 286 450 287 
<< pdiffusion >>
rect 12 287 13 288 
<< pdiffusion >>
rect 13 287 14 288 
<< pdiffusion >>
rect 14 287 15 288 
<< pdiffusion >>
rect 15 287 16 288 
<< pdiffusion >>
rect 16 287 17 288 
<< pdiffusion >>
rect 17 287 18 288 
<< pdiffusion >>
rect 30 287 31 288 
<< pdiffusion >>
rect 31 287 32 288 
<< pdiffusion >>
rect 32 287 33 288 
<< pdiffusion >>
rect 33 287 34 288 
<< pdiffusion >>
rect 34 287 35 288 
<< pdiffusion >>
rect 35 287 36 288 
<< pdiffusion >>
rect 48 287 49 288 
<< pdiffusion >>
rect 49 287 50 288 
<< pdiffusion >>
rect 50 287 51 288 
<< pdiffusion >>
rect 51 287 52 288 
<< pdiffusion >>
rect 52 287 53 288 
<< pdiffusion >>
rect 53 287 54 288 
<< m1 >>
rect 55 287 56 288 
<< m1 >>
rect 64 287 65 288 
<< pdiffusion >>
rect 66 287 67 288 
<< pdiffusion >>
rect 67 287 68 288 
<< pdiffusion >>
rect 68 287 69 288 
<< pdiffusion >>
rect 69 287 70 288 
<< pdiffusion >>
rect 70 287 71 288 
<< pdiffusion >>
rect 71 287 72 288 
<< pdiffusion >>
rect 84 287 85 288 
<< pdiffusion >>
rect 85 287 86 288 
<< pdiffusion >>
rect 86 287 87 288 
<< pdiffusion >>
rect 87 287 88 288 
<< m1 >>
rect 88 287 89 288 
<< pdiffusion >>
rect 88 287 89 288 
<< pdiffusion >>
rect 89 287 90 288 
<< m1 >>
rect 91 287 92 288 
<< pdiffusion >>
rect 102 287 103 288 
<< m1 >>
rect 103 287 104 288 
<< pdiffusion >>
rect 103 287 104 288 
<< pdiffusion >>
rect 104 287 105 288 
<< pdiffusion >>
rect 105 287 106 288 
<< pdiffusion >>
rect 106 287 107 288 
<< pdiffusion >>
rect 107 287 108 288 
<< pdiffusion >>
rect 120 287 121 288 
<< pdiffusion >>
rect 121 287 122 288 
<< pdiffusion >>
rect 122 287 123 288 
<< pdiffusion >>
rect 123 287 124 288 
<< pdiffusion >>
rect 124 287 125 288 
<< pdiffusion >>
rect 125 287 126 288 
<< m1 >>
rect 127 287 128 288 
<< pdiffusion >>
rect 138 287 139 288 
<< pdiffusion >>
rect 139 287 140 288 
<< pdiffusion >>
rect 140 287 141 288 
<< pdiffusion >>
rect 141 287 142 288 
<< pdiffusion >>
rect 142 287 143 288 
<< pdiffusion >>
rect 143 287 144 288 
<< m1 >>
rect 145 287 146 288 
<< pdiffusion >>
rect 156 287 157 288 
<< pdiffusion >>
rect 157 287 158 288 
<< pdiffusion >>
rect 158 287 159 288 
<< pdiffusion >>
rect 159 287 160 288 
<< pdiffusion >>
rect 160 287 161 288 
<< pdiffusion >>
rect 161 287 162 288 
<< m1 >>
rect 163 287 164 288 
<< pdiffusion >>
rect 174 287 175 288 
<< pdiffusion >>
rect 175 287 176 288 
<< pdiffusion >>
rect 176 287 177 288 
<< pdiffusion >>
rect 177 287 178 288 
<< pdiffusion >>
rect 178 287 179 288 
<< pdiffusion >>
rect 179 287 180 288 
<< m1 >>
rect 181 287 182 288 
<< m2 >>
rect 182 287 183 288 
<< pdiffusion >>
rect 192 287 193 288 
<< pdiffusion >>
rect 193 287 194 288 
<< pdiffusion >>
rect 194 287 195 288 
<< pdiffusion >>
rect 195 287 196 288 
<< m1 >>
rect 196 287 197 288 
<< pdiffusion >>
rect 196 287 197 288 
<< pdiffusion >>
rect 197 287 198 288 
<< pdiffusion >>
rect 210 287 211 288 
<< pdiffusion >>
rect 211 287 212 288 
<< pdiffusion >>
rect 212 287 213 288 
<< pdiffusion >>
rect 213 287 214 288 
<< pdiffusion >>
rect 214 287 215 288 
<< pdiffusion >>
rect 215 287 216 288 
<< m1 >>
rect 224 287 225 288 
<< m1 >>
rect 226 287 227 288 
<< pdiffusion >>
rect 228 287 229 288 
<< m1 >>
rect 229 287 230 288 
<< pdiffusion >>
rect 229 287 230 288 
<< pdiffusion >>
rect 230 287 231 288 
<< pdiffusion >>
rect 231 287 232 288 
<< m1 >>
rect 232 287 233 288 
<< pdiffusion >>
rect 232 287 233 288 
<< pdiffusion >>
rect 233 287 234 288 
<< m2 >>
rect 243 287 244 288 
<< m1 >>
rect 244 287 245 288 
<< pdiffusion >>
rect 246 287 247 288 
<< pdiffusion >>
rect 247 287 248 288 
<< pdiffusion >>
rect 248 287 249 288 
<< pdiffusion >>
rect 249 287 250 288 
<< pdiffusion >>
rect 250 287 251 288 
<< pdiffusion >>
rect 251 287 252 288 
<< m1 >>
rect 254 287 255 288 
<< m1 >>
rect 260 287 261 288 
<< pdiffusion >>
rect 264 287 265 288 
<< m1 >>
rect 265 287 266 288 
<< pdiffusion >>
rect 265 287 266 288 
<< pdiffusion >>
rect 266 287 267 288 
<< pdiffusion >>
rect 267 287 268 288 
<< pdiffusion >>
rect 268 287 269 288 
<< pdiffusion >>
rect 269 287 270 288 
<< pdiffusion >>
rect 300 287 301 288 
<< m1 >>
rect 301 287 302 288 
<< pdiffusion >>
rect 301 287 302 288 
<< pdiffusion >>
rect 302 287 303 288 
<< pdiffusion >>
rect 303 287 304 288 
<< m1 >>
rect 304 287 305 288 
<< pdiffusion >>
rect 304 287 305 288 
<< pdiffusion >>
rect 305 287 306 288 
<< m1 >>
rect 307 287 308 288 
<< m2 >>
rect 308 287 309 288 
<< pdiffusion >>
rect 318 287 319 288 
<< pdiffusion >>
rect 319 287 320 288 
<< pdiffusion >>
rect 320 287 321 288 
<< pdiffusion >>
rect 321 287 322 288 
<< pdiffusion >>
rect 322 287 323 288 
<< pdiffusion >>
rect 323 287 324 288 
<< pdiffusion >>
rect 336 287 337 288 
<< pdiffusion >>
rect 337 287 338 288 
<< pdiffusion >>
rect 338 287 339 288 
<< pdiffusion >>
rect 339 287 340 288 
<< pdiffusion >>
rect 340 287 341 288 
<< pdiffusion >>
rect 341 287 342 288 
<< m1 >>
rect 352 287 353 288 
<< pdiffusion >>
rect 354 287 355 288 
<< pdiffusion >>
rect 355 287 356 288 
<< pdiffusion >>
rect 356 287 357 288 
<< pdiffusion >>
rect 357 287 358 288 
<< pdiffusion >>
rect 358 287 359 288 
<< pdiffusion >>
rect 359 287 360 288 
<< pdiffusion >>
rect 372 287 373 288 
<< pdiffusion >>
rect 373 287 374 288 
<< pdiffusion >>
rect 374 287 375 288 
<< pdiffusion >>
rect 375 287 376 288 
<< pdiffusion >>
rect 376 287 377 288 
<< pdiffusion >>
rect 377 287 378 288 
<< pdiffusion >>
rect 390 287 391 288 
<< pdiffusion >>
rect 391 287 392 288 
<< pdiffusion >>
rect 392 287 393 288 
<< pdiffusion >>
rect 393 287 394 288 
<< pdiffusion >>
rect 394 287 395 288 
<< pdiffusion >>
rect 395 287 396 288 
<< m1 >>
rect 406 287 407 288 
<< pdiffusion >>
rect 408 287 409 288 
<< m1 >>
rect 409 287 410 288 
<< pdiffusion >>
rect 409 287 410 288 
<< pdiffusion >>
rect 410 287 411 288 
<< pdiffusion >>
rect 411 287 412 288 
<< pdiffusion >>
rect 412 287 413 288 
<< pdiffusion >>
rect 413 287 414 288 
<< pdiffusion >>
rect 426 287 427 288 
<< pdiffusion >>
rect 427 287 428 288 
<< pdiffusion >>
rect 428 287 429 288 
<< pdiffusion >>
rect 429 287 430 288 
<< pdiffusion >>
rect 430 287 431 288 
<< pdiffusion >>
rect 431 287 432 288 
<< pdiffusion >>
rect 444 287 445 288 
<< pdiffusion >>
rect 445 287 446 288 
<< pdiffusion >>
rect 446 287 447 288 
<< pdiffusion >>
rect 447 287 448 288 
<< pdiffusion >>
rect 448 287 449 288 
<< pdiffusion >>
rect 449 287 450 288 
<< m1 >>
rect 55 288 56 289 
<< m1 >>
rect 64 288 65 289 
<< m1 >>
rect 88 288 89 289 
<< m1 >>
rect 91 288 92 289 
<< m1 >>
rect 103 288 104 289 
<< m1 >>
rect 127 288 128 289 
<< m1 >>
rect 145 288 146 289 
<< m1 >>
rect 163 288 164 289 
<< m1 >>
rect 181 288 182 289 
<< m2 >>
rect 182 288 183 289 
<< m1 >>
rect 196 288 197 289 
<< m1 >>
rect 224 288 225 289 
<< m1 >>
rect 226 288 227 289 
<< m1 >>
rect 229 288 230 289 
<< m1 >>
rect 232 288 233 289 
<< m2 >>
rect 243 288 244 289 
<< m1 >>
rect 244 288 245 289 
<< m1 >>
rect 254 288 255 289 
<< m1 >>
rect 260 288 261 289 
<< m1 >>
rect 265 288 266 289 
<< m1 >>
rect 301 288 302 289 
<< m1 >>
rect 304 288 305 289 
<< m1 >>
rect 307 288 308 289 
<< m2 >>
rect 308 288 309 289 
<< m1 >>
rect 352 288 353 289 
<< m1 >>
rect 406 288 407 289 
<< m1 >>
rect 409 288 410 289 
<< m1 >>
rect 55 289 56 290 
<< m1 >>
rect 64 289 65 290 
<< m1 >>
rect 88 289 89 290 
<< m1 >>
rect 89 289 90 290 
<< m2 >>
rect 89 289 90 290 
<< m2c >>
rect 89 289 90 290 
<< m1 >>
rect 89 289 90 290 
<< m2 >>
rect 89 289 90 290 
<< m2 >>
rect 90 289 91 290 
<< m1 >>
rect 91 289 92 290 
<< m2 >>
rect 91 289 92 290 
<< m2 >>
rect 92 289 93 290 
<< m1 >>
rect 93 289 94 290 
<< m2 >>
rect 93 289 94 290 
<< m2c >>
rect 93 289 94 290 
<< m1 >>
rect 93 289 94 290 
<< m2 >>
rect 93 289 94 290 
<< m1 >>
rect 94 289 95 290 
<< m1 >>
rect 95 289 96 290 
<< m1 >>
rect 96 289 97 290 
<< m1 >>
rect 97 289 98 290 
<< m1 >>
rect 98 289 99 290 
<< m1 >>
rect 99 289 100 290 
<< m1 >>
rect 100 289 101 290 
<< m1 >>
rect 101 289 102 290 
<< m1 >>
rect 102 289 103 290 
<< m1 >>
rect 103 289 104 290 
<< m1 >>
rect 127 289 128 290 
<< m1 >>
rect 145 289 146 290 
<< m1 >>
rect 163 289 164 290 
<< m1 >>
rect 181 289 182 290 
<< m2 >>
rect 182 289 183 290 
<< m1 >>
rect 196 289 197 290 
<< m1 >>
rect 224 289 225 290 
<< m1 >>
rect 226 289 227 290 
<< m1 >>
rect 229 289 230 290 
<< m1 >>
rect 232 289 233 290 
<< m1 >>
rect 233 289 234 290 
<< m1 >>
rect 234 289 235 290 
<< m1 >>
rect 235 289 236 290 
<< m1 >>
rect 236 289 237 290 
<< m1 >>
rect 237 289 238 290 
<< m1 >>
rect 238 289 239 290 
<< m1 >>
rect 239 289 240 290 
<< m1 >>
rect 240 289 241 290 
<< m1 >>
rect 241 289 242 290 
<< m1 >>
rect 242 289 243 290 
<< m1 >>
rect 243 289 244 290 
<< m2 >>
rect 243 289 244 290 
<< m1 >>
rect 244 289 245 290 
<< m1 >>
rect 254 289 255 290 
<< m1 >>
rect 260 289 261 290 
<< m1 >>
rect 265 289 266 290 
<< m1 >>
rect 301 289 302 290 
<< m1 >>
rect 304 289 305 290 
<< m1 >>
rect 307 289 308 290 
<< m2 >>
rect 308 289 309 290 
<< m1 >>
rect 352 289 353 290 
<< m1 >>
rect 406 289 407 290 
<< m1 >>
rect 407 289 408 290 
<< m1 >>
rect 408 289 409 290 
<< m1 >>
rect 409 289 410 290 
<< m1 >>
rect 55 290 56 291 
<< m1 >>
rect 64 290 65 291 
<< m1 >>
rect 91 290 92 291 
<< m1 >>
rect 127 290 128 291 
<< m1 >>
rect 145 290 146 291 
<< m1 >>
rect 163 290 164 291 
<< m1 >>
rect 181 290 182 291 
<< m2 >>
rect 182 290 183 291 
<< m1 >>
rect 196 290 197 291 
<< m1 >>
rect 224 290 225 291 
<< m1 >>
rect 226 290 227 291 
<< m1 >>
rect 229 290 230 291 
<< m2 >>
rect 230 290 231 291 
<< m2 >>
rect 231 290 232 291 
<< m2 >>
rect 232 290 233 291 
<< m2 >>
rect 233 290 234 291 
<< m2 >>
rect 234 290 235 291 
<< m2 >>
rect 235 290 236 291 
<< m2 >>
rect 236 290 237 291 
<< m2 >>
rect 237 290 238 291 
<< m2 >>
rect 238 290 239 291 
<< m2 >>
rect 239 290 240 291 
<< m2 >>
rect 240 290 241 291 
<< m2 >>
rect 241 290 242 291 
<< m2 >>
rect 242 290 243 291 
<< m2 >>
rect 243 290 244 291 
<< m1 >>
rect 254 290 255 291 
<< m1 >>
rect 260 290 261 291 
<< m1 >>
rect 265 290 266 291 
<< m1 >>
rect 301 290 302 291 
<< m1 >>
rect 302 290 303 291 
<< m2 >>
rect 302 290 303 291 
<< m2c >>
rect 302 290 303 291 
<< m1 >>
rect 302 290 303 291 
<< m2 >>
rect 302 290 303 291 
<< m2 >>
rect 303 290 304 291 
<< m1 >>
rect 304 290 305 291 
<< m2 >>
rect 304 290 305 291 
<< m2 >>
rect 305 290 306 291 
<< m2 >>
rect 306 290 307 291 
<< m1 >>
rect 307 290 308 291 
<< m2 >>
rect 307 290 308 291 
<< m2 >>
rect 308 290 309 291 
<< m1 >>
rect 352 290 353 291 
<< m1 >>
rect 55 291 56 292 
<< m1 >>
rect 64 291 65 292 
<< m1 >>
rect 91 291 92 292 
<< m1 >>
rect 127 291 128 292 
<< m1 >>
rect 145 291 146 292 
<< m1 >>
rect 163 291 164 292 
<< m1 >>
rect 181 291 182 292 
<< m2 >>
rect 182 291 183 292 
<< m1 >>
rect 196 291 197 292 
<< m1 >>
rect 224 291 225 292 
<< m1 >>
rect 226 291 227 292 
<< m1 >>
rect 229 291 230 292 
<< m1 >>
rect 230 291 231 292 
<< m2 >>
rect 230 291 231 292 
<< m1 >>
rect 231 291 232 292 
<< m1 >>
rect 232 291 233 292 
<< m1 >>
rect 233 291 234 292 
<< m1 >>
rect 234 291 235 292 
<< m1 >>
rect 235 291 236 292 
<< m1 >>
rect 254 291 255 292 
<< m1 >>
rect 260 291 261 292 
<< m1 >>
rect 265 291 266 292 
<< m2 >>
rect 265 291 266 292 
<< m2c >>
rect 265 291 266 292 
<< m1 >>
rect 265 291 266 292 
<< m2 >>
rect 265 291 266 292 
<< m1 >>
rect 304 291 305 292 
<< m1 >>
rect 307 291 308 292 
<< m1 >>
rect 352 291 353 292 
<< m1 >>
rect 55 292 56 293 
<< m1 >>
rect 64 292 65 293 
<< m1 >>
rect 91 292 92 293 
<< m1 >>
rect 127 292 128 293 
<< m1 >>
rect 145 292 146 293 
<< m1 >>
rect 146 292 147 293 
<< m1 >>
rect 147 292 148 293 
<< m1 >>
rect 148 292 149 293 
<< m1 >>
rect 149 292 150 293 
<< m1 >>
rect 150 292 151 293 
<< m1 >>
rect 151 292 152 293 
<< m1 >>
rect 152 292 153 293 
<< m1 >>
rect 153 292 154 293 
<< m1 >>
rect 154 292 155 293 
<< m1 >>
rect 155 292 156 293 
<< m1 >>
rect 156 292 157 293 
<< m1 >>
rect 157 292 158 293 
<< m1 >>
rect 158 292 159 293 
<< m1 >>
rect 159 292 160 293 
<< m1 >>
rect 160 292 161 293 
<< m1 >>
rect 161 292 162 293 
<< m2 >>
rect 161 292 162 293 
<< m2c >>
rect 161 292 162 293 
<< m1 >>
rect 161 292 162 293 
<< m2 >>
rect 161 292 162 293 
<< m2 >>
rect 162 292 163 293 
<< m1 >>
rect 163 292 164 293 
<< m2 >>
rect 163 292 164 293 
<< m2 >>
rect 164 292 165 293 
<< m1 >>
rect 165 292 166 293 
<< m2 >>
rect 165 292 166 293 
<< m2c >>
rect 165 292 166 293 
<< m1 >>
rect 165 292 166 293 
<< m2 >>
rect 165 292 166 293 
<< m1 >>
rect 166 292 167 293 
<< m1 >>
rect 167 292 168 293 
<< m1 >>
rect 168 292 169 293 
<< m1 >>
rect 169 292 170 293 
<< m1 >>
rect 170 292 171 293 
<< m1 >>
rect 171 292 172 293 
<< m1 >>
rect 172 292 173 293 
<< m1 >>
rect 173 292 174 293 
<< m1 >>
rect 174 292 175 293 
<< m1 >>
rect 175 292 176 293 
<< m1 >>
rect 181 292 182 293 
<< m1 >>
rect 182 292 183 293 
<< m2 >>
rect 182 292 183 293 
<< m1 >>
rect 183 292 184 293 
<< m1 >>
rect 184 292 185 293 
<< m1 >>
rect 185 292 186 293 
<< m1 >>
rect 186 292 187 293 
<< m1 >>
rect 187 292 188 293 
<< m1 >>
rect 188 292 189 293 
<< m1 >>
rect 189 292 190 293 
<< m1 >>
rect 190 292 191 293 
<< m1 >>
rect 191 292 192 293 
<< m1 >>
rect 192 292 193 293 
<< m1 >>
rect 193 292 194 293 
<< m1 >>
rect 194 292 195 293 
<< m1 >>
rect 195 292 196 293 
<< m1 >>
rect 196 292 197 293 
<< m2 >>
rect 206 292 207 293 
<< m2 >>
rect 207 292 208 293 
<< m2 >>
rect 208 292 209 293 
<< m2 >>
rect 209 292 210 293 
<< m1 >>
rect 210 292 211 293 
<< m2 >>
rect 210 292 211 293 
<< m2c >>
rect 210 292 211 293 
<< m1 >>
rect 210 292 211 293 
<< m2 >>
rect 210 292 211 293 
<< m1 >>
rect 211 292 212 293 
<< m1 >>
rect 212 292 213 293 
<< m1 >>
rect 213 292 214 293 
<< m1 >>
rect 214 292 215 293 
<< m1 >>
rect 215 292 216 293 
<< m1 >>
rect 216 292 217 293 
<< m1 >>
rect 217 292 218 293 
<< m1 >>
rect 218 292 219 293 
<< m1 >>
rect 219 292 220 293 
<< m1 >>
rect 220 292 221 293 
<< m1 >>
rect 221 292 222 293 
<< m1 >>
rect 222 292 223 293 
<< m1 >>
rect 223 292 224 293 
<< m1 >>
rect 224 292 225 293 
<< m1 >>
rect 226 292 227 293 
<< m2 >>
rect 228 292 229 293 
<< m2 >>
rect 229 292 230 293 
<< m2 >>
rect 230 292 231 293 
<< m1 >>
rect 235 292 236 293 
<< m1 >>
rect 254 292 255 293 
<< m1 >>
rect 260 292 261 293 
<< m2 >>
rect 265 292 266 293 
<< m2 >>
rect 266 292 267 293 
<< m1 >>
rect 304 292 305 293 
<< m1 >>
rect 307 292 308 293 
<< m1 >>
rect 352 292 353 293 
<< m1 >>
rect 55 293 56 294 
<< m1 >>
rect 64 293 65 294 
<< m1 >>
rect 91 293 92 294 
<< m1 >>
rect 127 293 128 294 
<< m1 >>
rect 163 293 164 294 
<< m1 >>
rect 175 293 176 294 
<< m2 >>
rect 182 293 183 294 
<< m2 >>
rect 183 293 184 294 
<< m2 >>
rect 184 293 185 294 
<< m2 >>
rect 185 293 186 294 
<< m2 >>
rect 186 293 187 294 
<< m2 >>
rect 187 293 188 294 
<< m2 >>
rect 188 293 189 294 
<< m2 >>
rect 189 293 190 294 
<< m2 >>
rect 190 293 191 294 
<< m2 >>
rect 191 293 192 294 
<< m2 >>
rect 192 293 193 294 
<< m2 >>
rect 193 293 194 294 
<< m2 >>
rect 194 293 195 294 
<< m2 >>
rect 195 293 196 294 
<< m2 >>
rect 196 293 197 294 
<< m2 >>
rect 197 293 198 294 
<< m1 >>
rect 198 293 199 294 
<< m2 >>
rect 198 293 199 294 
<< m2c >>
rect 198 293 199 294 
<< m1 >>
rect 198 293 199 294 
<< m2 >>
rect 198 293 199 294 
<< m1 >>
rect 199 293 200 294 
<< m1 >>
rect 200 293 201 294 
<< m1 >>
rect 201 293 202 294 
<< m1 >>
rect 202 293 203 294 
<< m1 >>
rect 203 293 204 294 
<< m1 >>
rect 204 293 205 294 
<< m1 >>
rect 205 293 206 294 
<< m1 >>
rect 206 293 207 294 
<< m2 >>
rect 206 293 207 294 
<< m1 >>
rect 207 293 208 294 
<< m1 >>
rect 208 293 209 294 
<< m1 >>
rect 226 293 227 294 
<< m1 >>
rect 228 293 229 294 
<< m2 >>
rect 228 293 229 294 
<< m2c >>
rect 228 293 229 294 
<< m1 >>
rect 228 293 229 294 
<< m2 >>
rect 228 293 229 294 
<< m1 >>
rect 235 293 236 294 
<< m1 >>
rect 254 293 255 294 
<< m2 >>
rect 254 293 255 294 
<< m2c >>
rect 254 293 255 294 
<< m1 >>
rect 254 293 255 294 
<< m2 >>
rect 254 293 255 294 
<< m1 >>
rect 260 293 261 294 
<< m1 >>
rect 261 293 262 294 
<< m1 >>
rect 262 293 263 294 
<< m1 >>
rect 263 293 264 294 
<< m1 >>
rect 264 293 265 294 
<< m1 >>
rect 265 293 266 294 
<< m1 >>
rect 266 293 267 294 
<< m2 >>
rect 266 293 267 294 
<< m1 >>
rect 267 293 268 294 
<< m1 >>
rect 268 293 269 294 
<< m1 >>
rect 269 293 270 294 
<< m1 >>
rect 270 293 271 294 
<< m1 >>
rect 271 293 272 294 
<< m1 >>
rect 272 293 273 294 
<< m1 >>
rect 273 293 274 294 
<< m1 >>
rect 274 293 275 294 
<< m1 >>
rect 275 293 276 294 
<< m1 >>
rect 276 293 277 294 
<< m1 >>
rect 277 293 278 294 
<< m1 >>
rect 278 293 279 294 
<< m1 >>
rect 279 293 280 294 
<< m1 >>
rect 280 293 281 294 
<< m2 >>
rect 280 293 281 294 
<< m2c >>
rect 280 293 281 294 
<< m1 >>
rect 280 293 281 294 
<< m2 >>
rect 280 293 281 294 
<< m1 >>
rect 304 293 305 294 
<< m1 >>
rect 307 293 308 294 
<< m1 >>
rect 352 293 353 294 
<< m1 >>
rect 55 294 56 295 
<< m1 >>
rect 64 294 65 295 
<< m1 >>
rect 91 294 92 295 
<< m1 >>
rect 127 294 128 295 
<< m1 >>
rect 163 294 164 295 
<< m1 >>
rect 175 294 176 295 
<< m2 >>
rect 206 294 207 295 
<< m1 >>
rect 208 294 209 295 
<< m1 >>
rect 226 294 227 295 
<< m1 >>
rect 228 294 229 295 
<< m1 >>
rect 235 294 236 295 
<< m2 >>
rect 254 294 255 295 
<< m2 >>
rect 266 294 267 295 
<< m2 >>
rect 280 294 281 295 
<< m1 >>
rect 304 294 305 295 
<< m1 >>
rect 307 294 308 295 
<< m1 >>
rect 352 294 353 295 
<< m1 >>
rect 55 295 56 296 
<< m1 >>
rect 64 295 65 296 
<< m1 >>
rect 91 295 92 296 
<< m1 >>
rect 127 295 128 296 
<< m1 >>
rect 163 295 164 296 
<< m1 >>
rect 175 295 176 296 
<< m1 >>
rect 206 295 207 296 
<< m2 >>
rect 206 295 207 296 
<< m2c >>
rect 206 295 207 296 
<< m1 >>
rect 206 295 207 296 
<< m2 >>
rect 206 295 207 296 
<< m1 >>
rect 208 295 209 296 
<< m1 >>
rect 226 295 227 296 
<< m1 >>
rect 228 295 229 296 
<< m1 >>
rect 235 295 236 296 
<< m1 >>
rect 237 295 238 296 
<< m1 >>
rect 238 295 239 296 
<< m1 >>
rect 239 295 240 296 
<< m1 >>
rect 240 295 241 296 
<< m1 >>
rect 241 295 242 296 
<< m1 >>
rect 242 295 243 296 
<< m1 >>
rect 243 295 244 296 
<< m1 >>
rect 244 295 245 296 
<< m1 >>
rect 245 295 246 296 
<< m1 >>
rect 246 295 247 296 
<< m1 >>
rect 247 295 248 296 
<< m1 >>
rect 248 295 249 296 
<< m1 >>
rect 249 295 250 296 
<< m1 >>
rect 250 295 251 296 
<< m1 >>
rect 251 295 252 296 
<< m1 >>
rect 252 295 253 296 
<< m1 >>
rect 253 295 254 296 
<< m1 >>
rect 254 295 255 296 
<< m2 >>
rect 254 295 255 296 
<< m1 >>
rect 255 295 256 296 
<< m1 >>
rect 256 295 257 296 
<< m1 >>
rect 257 295 258 296 
<< m1 >>
rect 258 295 259 296 
<< m1 >>
rect 259 295 260 296 
<< m1 >>
rect 260 295 261 296 
<< m1 >>
rect 261 295 262 296 
<< m1 >>
rect 262 295 263 296 
<< m1 >>
rect 263 295 264 296 
<< m1 >>
rect 264 295 265 296 
<< m1 >>
rect 265 295 266 296 
<< m1 >>
rect 266 295 267 296 
<< m2 >>
rect 266 295 267 296 
<< m1 >>
rect 267 295 268 296 
<< m1 >>
rect 268 295 269 296 
<< m1 >>
rect 269 295 270 296 
<< m1 >>
rect 270 295 271 296 
<< m1 >>
rect 271 295 272 296 
<< m1 >>
rect 272 295 273 296 
<< m1 >>
rect 273 295 274 296 
<< m1 >>
rect 274 295 275 296 
<< m1 >>
rect 275 295 276 296 
<< m1 >>
rect 276 295 277 296 
<< m1 >>
rect 277 295 278 296 
<< m1 >>
rect 278 295 279 296 
<< m1 >>
rect 279 295 280 296 
<< m1 >>
rect 280 295 281 296 
<< m2 >>
rect 280 295 281 296 
<< m1 >>
rect 281 295 282 296 
<< m1 >>
rect 282 295 283 296 
<< m1 >>
rect 283 295 284 296 
<< m1 >>
rect 284 295 285 296 
<< m1 >>
rect 285 295 286 296 
<< m1 >>
rect 286 295 287 296 
<< m1 >>
rect 287 295 288 296 
<< m1 >>
rect 288 295 289 296 
<< m1 >>
rect 289 295 290 296 
<< m1 >>
rect 290 295 291 296 
<< m1 >>
rect 291 295 292 296 
<< m1 >>
rect 292 295 293 296 
<< m1 >>
rect 293 295 294 296 
<< m1 >>
rect 294 295 295 296 
<< m1 >>
rect 295 295 296 296 
<< m1 >>
rect 296 295 297 296 
<< m1 >>
rect 297 295 298 296 
<< m1 >>
rect 298 295 299 296 
<< m1 >>
rect 299 295 300 296 
<< m1 >>
rect 300 295 301 296 
<< m1 >>
rect 301 295 302 296 
<< m1 >>
rect 302 295 303 296 
<< m1 >>
rect 303 295 304 296 
<< m1 >>
rect 304 295 305 296 
<< m1 >>
rect 307 295 308 296 
<< m1 >>
rect 352 295 353 296 
<< m1 >>
rect 55 296 56 297 
<< m1 >>
rect 64 296 65 297 
<< m1 >>
rect 91 296 92 297 
<< m1 >>
rect 127 296 128 297 
<< m1 >>
rect 163 296 164 297 
<< m1 >>
rect 175 296 176 297 
<< m1 >>
rect 206 296 207 297 
<< m2 >>
rect 206 296 207 297 
<< m1 >>
rect 208 296 209 297 
<< m2 >>
rect 208 296 209 297 
<< m2c >>
rect 208 296 209 297 
<< m1 >>
rect 208 296 209 297 
<< m2 >>
rect 208 296 209 297 
<< m1 >>
rect 226 296 227 297 
<< m2 >>
rect 226 296 227 297 
<< m2c >>
rect 226 296 227 297 
<< m1 >>
rect 226 296 227 297 
<< m2 >>
rect 226 296 227 297 
<< m1 >>
rect 228 296 229 297 
<< m1 >>
rect 235 296 236 297 
<< m1 >>
rect 237 296 238 297 
<< m2 >>
rect 254 296 255 297 
<< m2 >>
rect 266 296 267 297 
<< m2 >>
rect 280 296 281 297 
<< m1 >>
rect 307 296 308 297 
<< m1 >>
rect 352 296 353 297 
<< m1 >>
rect 55 297 56 298 
<< m1 >>
rect 64 297 65 298 
<< m1 >>
rect 91 297 92 298 
<< m1 >>
rect 127 297 128 298 
<< m1 >>
rect 163 297 164 298 
<< m1 >>
rect 175 297 176 298 
<< m2 >>
rect 206 297 207 298 
<< m2 >>
rect 208 297 209 298 
<< m2 >>
rect 226 297 227 298 
<< m1 >>
rect 228 297 229 298 
<< m1 >>
rect 235 297 236 298 
<< m1 >>
rect 237 297 238 298 
<< m1 >>
rect 254 297 255 298 
<< m2 >>
rect 254 297 255 298 
<< m2c >>
rect 254 297 255 298 
<< m1 >>
rect 254 297 255 298 
<< m2 >>
rect 254 297 255 298 
<< m1 >>
rect 255 297 256 298 
<< m1 >>
rect 256 297 257 298 
<< m1 >>
rect 257 297 258 298 
<< m1 >>
rect 266 297 267 298 
<< m2 >>
rect 266 297 267 298 
<< m2c >>
rect 266 297 267 298 
<< m1 >>
rect 266 297 267 298 
<< m2 >>
rect 266 297 267 298 
<< m1 >>
rect 267 297 268 298 
<< m1 >>
rect 268 297 269 298 
<< m1 >>
rect 269 297 270 298 
<< m1 >>
rect 270 297 271 298 
<< m1 >>
rect 271 297 272 298 
<< m1 >>
rect 280 297 281 298 
<< m2 >>
rect 280 297 281 298 
<< m2c >>
rect 280 297 281 298 
<< m1 >>
rect 280 297 281 298 
<< m2 >>
rect 280 297 281 298 
<< m1 >>
rect 283 297 284 298 
<< m1 >>
rect 284 297 285 298 
<< m1 >>
rect 285 297 286 298 
<< m1 >>
rect 286 297 287 298 
<< m1 >>
rect 287 297 288 298 
<< m1 >>
rect 288 297 289 298 
<< m1 >>
rect 289 297 290 298 
<< m1 >>
rect 307 297 308 298 
<< m1 >>
rect 352 297 353 298 
<< m1 >>
rect 55 298 56 299 
<< m1 >>
rect 64 298 65 299 
<< m1 >>
rect 91 298 92 299 
<< m1 >>
rect 124 298 125 299 
<< m1 >>
rect 125 298 126 299 
<< m1 >>
rect 126 298 127 299 
<< m1 >>
rect 127 298 128 299 
<< m1 >>
rect 163 298 164 299 
<< m1 >>
rect 175 298 176 299 
<< m1 >>
rect 196 298 197 299 
<< m1 >>
rect 197 298 198 299 
<< m1 >>
rect 198 298 199 299 
<< m1 >>
rect 199 298 200 299 
<< m1 >>
rect 200 298 201 299 
<< m1 >>
rect 201 298 202 299 
<< m1 >>
rect 202 298 203 299 
<< m1 >>
rect 203 298 204 299 
<< m1 >>
rect 204 298 205 299 
<< m1 >>
rect 205 298 206 299 
<< m1 >>
rect 206 298 207 299 
<< m2 >>
rect 206 298 207 299 
<< m1 >>
rect 207 298 208 299 
<< m1 >>
rect 208 298 209 299 
<< m2 >>
rect 208 298 209 299 
<< m1 >>
rect 217 298 218 299 
<< m1 >>
rect 218 298 219 299 
<< m1 >>
rect 219 298 220 299 
<< m1 >>
rect 220 298 221 299 
<< m1 >>
rect 221 298 222 299 
<< m1 >>
rect 222 298 223 299 
<< m1 >>
rect 223 298 224 299 
<< m1 >>
rect 224 298 225 299 
<< m1 >>
rect 225 298 226 299 
<< m1 >>
rect 226 298 227 299 
<< m2 >>
rect 226 298 227 299 
<< m1 >>
rect 227 298 228 299 
<< m1 >>
rect 228 298 229 299 
<< m1 >>
rect 235 298 236 299 
<< m1 >>
rect 237 298 238 299 
<< m1 >>
rect 257 298 258 299 
<< m1 >>
rect 271 298 272 299 
<< m1 >>
rect 280 298 281 299 
<< m1 >>
rect 283 298 284 299 
<< m1 >>
rect 289 298 290 299 
<< m1 >>
rect 307 298 308 299 
<< m1 >>
rect 352 298 353 299 
<< m1 >>
rect 55 299 56 300 
<< m1 >>
rect 64 299 65 300 
<< m1 >>
rect 91 299 92 300 
<< m1 >>
rect 124 299 125 300 
<< m1 >>
rect 163 299 164 300 
<< m1 >>
rect 175 299 176 300 
<< m1 >>
rect 196 299 197 300 
<< m2 >>
rect 206 299 207 300 
<< m1 >>
rect 208 299 209 300 
<< m2 >>
rect 208 299 209 300 
<< m1 >>
rect 217 299 218 300 
<< m2 >>
rect 226 299 227 300 
<< m1 >>
rect 235 299 236 300 
<< m1 >>
rect 237 299 238 300 
<< m1 >>
rect 257 299 258 300 
<< m1 >>
rect 271 299 272 300 
<< m1 >>
rect 280 299 281 300 
<< m1 >>
rect 283 299 284 300 
<< m1 >>
rect 289 299 290 300 
<< m1 >>
rect 307 299 308 300 
<< m1 >>
rect 352 299 353 300 
<< pdiffusion >>
rect 12 300 13 301 
<< pdiffusion >>
rect 13 300 14 301 
<< pdiffusion >>
rect 14 300 15 301 
<< pdiffusion >>
rect 15 300 16 301 
<< pdiffusion >>
rect 16 300 17 301 
<< pdiffusion >>
rect 17 300 18 301 
<< pdiffusion >>
rect 30 300 31 301 
<< pdiffusion >>
rect 31 300 32 301 
<< pdiffusion >>
rect 32 300 33 301 
<< pdiffusion >>
rect 33 300 34 301 
<< pdiffusion >>
rect 34 300 35 301 
<< pdiffusion >>
rect 35 300 36 301 
<< pdiffusion >>
rect 48 300 49 301 
<< pdiffusion >>
rect 49 300 50 301 
<< pdiffusion >>
rect 50 300 51 301 
<< pdiffusion >>
rect 51 300 52 301 
<< pdiffusion >>
rect 52 300 53 301 
<< pdiffusion >>
rect 53 300 54 301 
<< m1 >>
rect 55 300 56 301 
<< m1 >>
rect 64 300 65 301 
<< pdiffusion >>
rect 66 300 67 301 
<< pdiffusion >>
rect 67 300 68 301 
<< pdiffusion >>
rect 68 300 69 301 
<< pdiffusion >>
rect 69 300 70 301 
<< pdiffusion >>
rect 70 300 71 301 
<< pdiffusion >>
rect 71 300 72 301 
<< pdiffusion >>
rect 84 300 85 301 
<< pdiffusion >>
rect 85 300 86 301 
<< pdiffusion >>
rect 86 300 87 301 
<< pdiffusion >>
rect 87 300 88 301 
<< pdiffusion >>
rect 88 300 89 301 
<< pdiffusion >>
rect 89 300 90 301 
<< m1 >>
rect 91 300 92 301 
<< pdiffusion >>
rect 102 300 103 301 
<< pdiffusion >>
rect 103 300 104 301 
<< pdiffusion >>
rect 104 300 105 301 
<< pdiffusion >>
rect 105 300 106 301 
<< pdiffusion >>
rect 106 300 107 301 
<< pdiffusion >>
rect 107 300 108 301 
<< pdiffusion >>
rect 120 300 121 301 
<< pdiffusion >>
rect 121 300 122 301 
<< pdiffusion >>
rect 122 300 123 301 
<< pdiffusion >>
rect 123 300 124 301 
<< m1 >>
rect 124 300 125 301 
<< pdiffusion >>
rect 124 300 125 301 
<< pdiffusion >>
rect 125 300 126 301 
<< pdiffusion >>
rect 138 300 139 301 
<< pdiffusion >>
rect 139 300 140 301 
<< pdiffusion >>
rect 140 300 141 301 
<< pdiffusion >>
rect 141 300 142 301 
<< pdiffusion >>
rect 142 300 143 301 
<< pdiffusion >>
rect 143 300 144 301 
<< pdiffusion >>
rect 156 300 157 301 
<< pdiffusion >>
rect 157 300 158 301 
<< pdiffusion >>
rect 158 300 159 301 
<< pdiffusion >>
rect 159 300 160 301 
<< pdiffusion >>
rect 160 300 161 301 
<< pdiffusion >>
rect 161 300 162 301 
<< m1 >>
rect 163 300 164 301 
<< pdiffusion >>
rect 174 300 175 301 
<< m1 >>
rect 175 300 176 301 
<< pdiffusion >>
rect 175 300 176 301 
<< pdiffusion >>
rect 176 300 177 301 
<< pdiffusion >>
rect 177 300 178 301 
<< pdiffusion >>
rect 178 300 179 301 
<< pdiffusion >>
rect 179 300 180 301 
<< pdiffusion >>
rect 192 300 193 301 
<< pdiffusion >>
rect 193 300 194 301 
<< pdiffusion >>
rect 194 300 195 301 
<< pdiffusion >>
rect 195 300 196 301 
<< m1 >>
rect 196 300 197 301 
<< pdiffusion >>
rect 196 300 197 301 
<< pdiffusion >>
rect 197 300 198 301 
<< m1 >>
rect 206 300 207 301 
<< m2 >>
rect 206 300 207 301 
<< m2c >>
rect 206 300 207 301 
<< m1 >>
rect 206 300 207 301 
<< m2 >>
rect 206 300 207 301 
<< m1 >>
rect 208 300 209 301 
<< m2 >>
rect 208 300 209 301 
<< pdiffusion >>
rect 210 300 211 301 
<< pdiffusion >>
rect 211 300 212 301 
<< pdiffusion >>
rect 212 300 213 301 
<< pdiffusion >>
rect 213 300 214 301 
<< pdiffusion >>
rect 214 300 215 301 
<< pdiffusion >>
rect 215 300 216 301 
<< m1 >>
rect 217 300 218 301 
<< m1 >>
rect 226 300 227 301 
<< m2 >>
rect 226 300 227 301 
<< m2c >>
rect 226 300 227 301 
<< m1 >>
rect 226 300 227 301 
<< m2 >>
rect 226 300 227 301 
<< pdiffusion >>
rect 228 300 229 301 
<< pdiffusion >>
rect 229 300 230 301 
<< pdiffusion >>
rect 230 300 231 301 
<< pdiffusion >>
rect 231 300 232 301 
<< pdiffusion >>
rect 232 300 233 301 
<< pdiffusion >>
rect 233 300 234 301 
<< m1 >>
rect 235 300 236 301 
<< m1 >>
rect 237 300 238 301 
<< pdiffusion >>
rect 246 300 247 301 
<< pdiffusion >>
rect 247 300 248 301 
<< pdiffusion >>
rect 248 300 249 301 
<< pdiffusion >>
rect 249 300 250 301 
<< pdiffusion >>
rect 250 300 251 301 
<< pdiffusion >>
rect 251 300 252 301 
<< m1 >>
rect 257 300 258 301 
<< pdiffusion >>
rect 264 300 265 301 
<< pdiffusion >>
rect 265 300 266 301 
<< pdiffusion >>
rect 266 300 267 301 
<< pdiffusion >>
rect 267 300 268 301 
<< pdiffusion >>
rect 268 300 269 301 
<< pdiffusion >>
rect 269 300 270 301 
<< m1 >>
rect 271 300 272 301 
<< m1 >>
rect 280 300 281 301 
<< pdiffusion >>
rect 282 300 283 301 
<< m1 >>
rect 283 300 284 301 
<< pdiffusion >>
rect 283 300 284 301 
<< pdiffusion >>
rect 284 300 285 301 
<< pdiffusion >>
rect 285 300 286 301 
<< pdiffusion >>
rect 286 300 287 301 
<< pdiffusion >>
rect 287 300 288 301 
<< m1 >>
rect 289 300 290 301 
<< pdiffusion >>
rect 300 300 301 301 
<< pdiffusion >>
rect 301 300 302 301 
<< pdiffusion >>
rect 302 300 303 301 
<< pdiffusion >>
rect 303 300 304 301 
<< pdiffusion >>
rect 304 300 305 301 
<< pdiffusion >>
rect 305 300 306 301 
<< m1 >>
rect 307 300 308 301 
<< pdiffusion >>
rect 318 300 319 301 
<< pdiffusion >>
rect 319 300 320 301 
<< pdiffusion >>
rect 320 300 321 301 
<< pdiffusion >>
rect 321 300 322 301 
<< pdiffusion >>
rect 322 300 323 301 
<< pdiffusion >>
rect 323 300 324 301 
<< pdiffusion >>
rect 336 300 337 301 
<< pdiffusion >>
rect 337 300 338 301 
<< pdiffusion >>
rect 338 300 339 301 
<< pdiffusion >>
rect 339 300 340 301 
<< pdiffusion >>
rect 340 300 341 301 
<< pdiffusion >>
rect 341 300 342 301 
<< m1 >>
rect 352 300 353 301 
<< pdiffusion >>
rect 354 300 355 301 
<< pdiffusion >>
rect 355 300 356 301 
<< pdiffusion >>
rect 356 300 357 301 
<< pdiffusion >>
rect 357 300 358 301 
<< pdiffusion >>
rect 358 300 359 301 
<< pdiffusion >>
rect 359 300 360 301 
<< pdiffusion >>
rect 372 300 373 301 
<< pdiffusion >>
rect 373 300 374 301 
<< pdiffusion >>
rect 374 300 375 301 
<< pdiffusion >>
rect 375 300 376 301 
<< pdiffusion >>
rect 376 300 377 301 
<< pdiffusion >>
rect 377 300 378 301 
<< pdiffusion >>
rect 390 300 391 301 
<< pdiffusion >>
rect 391 300 392 301 
<< pdiffusion >>
rect 392 300 393 301 
<< pdiffusion >>
rect 393 300 394 301 
<< pdiffusion >>
rect 394 300 395 301 
<< pdiffusion >>
rect 395 300 396 301 
<< pdiffusion >>
rect 408 300 409 301 
<< pdiffusion >>
rect 409 300 410 301 
<< pdiffusion >>
rect 410 300 411 301 
<< pdiffusion >>
rect 411 300 412 301 
<< pdiffusion >>
rect 412 300 413 301 
<< pdiffusion >>
rect 413 300 414 301 
<< pdiffusion >>
rect 426 300 427 301 
<< pdiffusion >>
rect 427 300 428 301 
<< pdiffusion >>
rect 428 300 429 301 
<< pdiffusion >>
rect 429 300 430 301 
<< pdiffusion >>
rect 430 300 431 301 
<< pdiffusion >>
rect 431 300 432 301 
<< pdiffusion >>
rect 444 300 445 301 
<< pdiffusion >>
rect 445 300 446 301 
<< pdiffusion >>
rect 446 300 447 301 
<< pdiffusion >>
rect 447 300 448 301 
<< pdiffusion >>
rect 448 300 449 301 
<< pdiffusion >>
rect 449 300 450 301 
<< pdiffusion >>
rect 12 301 13 302 
<< pdiffusion >>
rect 13 301 14 302 
<< pdiffusion >>
rect 14 301 15 302 
<< pdiffusion >>
rect 15 301 16 302 
<< pdiffusion >>
rect 16 301 17 302 
<< pdiffusion >>
rect 17 301 18 302 
<< pdiffusion >>
rect 30 301 31 302 
<< pdiffusion >>
rect 31 301 32 302 
<< pdiffusion >>
rect 32 301 33 302 
<< pdiffusion >>
rect 33 301 34 302 
<< pdiffusion >>
rect 34 301 35 302 
<< pdiffusion >>
rect 35 301 36 302 
<< pdiffusion >>
rect 48 301 49 302 
<< pdiffusion >>
rect 49 301 50 302 
<< pdiffusion >>
rect 50 301 51 302 
<< pdiffusion >>
rect 51 301 52 302 
<< pdiffusion >>
rect 52 301 53 302 
<< pdiffusion >>
rect 53 301 54 302 
<< m1 >>
rect 55 301 56 302 
<< m1 >>
rect 64 301 65 302 
<< pdiffusion >>
rect 66 301 67 302 
<< pdiffusion >>
rect 67 301 68 302 
<< pdiffusion >>
rect 68 301 69 302 
<< pdiffusion >>
rect 69 301 70 302 
<< pdiffusion >>
rect 70 301 71 302 
<< pdiffusion >>
rect 71 301 72 302 
<< pdiffusion >>
rect 84 301 85 302 
<< pdiffusion >>
rect 85 301 86 302 
<< pdiffusion >>
rect 86 301 87 302 
<< pdiffusion >>
rect 87 301 88 302 
<< pdiffusion >>
rect 88 301 89 302 
<< pdiffusion >>
rect 89 301 90 302 
<< m1 >>
rect 91 301 92 302 
<< pdiffusion >>
rect 102 301 103 302 
<< pdiffusion >>
rect 103 301 104 302 
<< pdiffusion >>
rect 104 301 105 302 
<< pdiffusion >>
rect 105 301 106 302 
<< pdiffusion >>
rect 106 301 107 302 
<< pdiffusion >>
rect 107 301 108 302 
<< pdiffusion >>
rect 120 301 121 302 
<< pdiffusion >>
rect 121 301 122 302 
<< pdiffusion >>
rect 122 301 123 302 
<< pdiffusion >>
rect 123 301 124 302 
<< pdiffusion >>
rect 124 301 125 302 
<< pdiffusion >>
rect 125 301 126 302 
<< pdiffusion >>
rect 138 301 139 302 
<< pdiffusion >>
rect 139 301 140 302 
<< pdiffusion >>
rect 140 301 141 302 
<< pdiffusion >>
rect 141 301 142 302 
<< pdiffusion >>
rect 142 301 143 302 
<< pdiffusion >>
rect 143 301 144 302 
<< pdiffusion >>
rect 156 301 157 302 
<< pdiffusion >>
rect 157 301 158 302 
<< pdiffusion >>
rect 158 301 159 302 
<< pdiffusion >>
rect 159 301 160 302 
<< pdiffusion >>
rect 160 301 161 302 
<< pdiffusion >>
rect 161 301 162 302 
<< m1 >>
rect 163 301 164 302 
<< pdiffusion >>
rect 174 301 175 302 
<< pdiffusion >>
rect 175 301 176 302 
<< pdiffusion >>
rect 176 301 177 302 
<< pdiffusion >>
rect 177 301 178 302 
<< pdiffusion >>
rect 178 301 179 302 
<< pdiffusion >>
rect 179 301 180 302 
<< pdiffusion >>
rect 192 301 193 302 
<< pdiffusion >>
rect 193 301 194 302 
<< pdiffusion >>
rect 194 301 195 302 
<< pdiffusion >>
rect 195 301 196 302 
<< pdiffusion >>
rect 196 301 197 302 
<< pdiffusion >>
rect 197 301 198 302 
<< m1 >>
rect 206 301 207 302 
<< m1 >>
rect 208 301 209 302 
<< m2 >>
rect 208 301 209 302 
<< pdiffusion >>
rect 210 301 211 302 
<< pdiffusion >>
rect 211 301 212 302 
<< pdiffusion >>
rect 212 301 213 302 
<< pdiffusion >>
rect 213 301 214 302 
<< pdiffusion >>
rect 214 301 215 302 
<< pdiffusion >>
rect 215 301 216 302 
<< m1 >>
rect 217 301 218 302 
<< m1 >>
rect 226 301 227 302 
<< pdiffusion >>
rect 228 301 229 302 
<< pdiffusion >>
rect 229 301 230 302 
<< pdiffusion >>
rect 230 301 231 302 
<< pdiffusion >>
rect 231 301 232 302 
<< pdiffusion >>
rect 232 301 233 302 
<< pdiffusion >>
rect 233 301 234 302 
<< m1 >>
rect 235 301 236 302 
<< m1 >>
rect 237 301 238 302 
<< pdiffusion >>
rect 246 301 247 302 
<< pdiffusion >>
rect 247 301 248 302 
<< pdiffusion >>
rect 248 301 249 302 
<< pdiffusion >>
rect 249 301 250 302 
<< pdiffusion >>
rect 250 301 251 302 
<< pdiffusion >>
rect 251 301 252 302 
<< m1 >>
rect 257 301 258 302 
<< pdiffusion >>
rect 264 301 265 302 
<< pdiffusion >>
rect 265 301 266 302 
<< pdiffusion >>
rect 266 301 267 302 
<< pdiffusion >>
rect 267 301 268 302 
<< pdiffusion >>
rect 268 301 269 302 
<< pdiffusion >>
rect 269 301 270 302 
<< m1 >>
rect 271 301 272 302 
<< m1 >>
rect 280 301 281 302 
<< pdiffusion >>
rect 282 301 283 302 
<< pdiffusion >>
rect 283 301 284 302 
<< pdiffusion >>
rect 284 301 285 302 
<< pdiffusion >>
rect 285 301 286 302 
<< pdiffusion >>
rect 286 301 287 302 
<< pdiffusion >>
rect 287 301 288 302 
<< m1 >>
rect 289 301 290 302 
<< pdiffusion >>
rect 300 301 301 302 
<< pdiffusion >>
rect 301 301 302 302 
<< pdiffusion >>
rect 302 301 303 302 
<< pdiffusion >>
rect 303 301 304 302 
<< pdiffusion >>
rect 304 301 305 302 
<< pdiffusion >>
rect 305 301 306 302 
<< m1 >>
rect 307 301 308 302 
<< pdiffusion >>
rect 318 301 319 302 
<< pdiffusion >>
rect 319 301 320 302 
<< pdiffusion >>
rect 320 301 321 302 
<< pdiffusion >>
rect 321 301 322 302 
<< pdiffusion >>
rect 322 301 323 302 
<< pdiffusion >>
rect 323 301 324 302 
<< pdiffusion >>
rect 336 301 337 302 
<< pdiffusion >>
rect 337 301 338 302 
<< pdiffusion >>
rect 338 301 339 302 
<< pdiffusion >>
rect 339 301 340 302 
<< pdiffusion >>
rect 340 301 341 302 
<< pdiffusion >>
rect 341 301 342 302 
<< m1 >>
rect 352 301 353 302 
<< pdiffusion >>
rect 354 301 355 302 
<< pdiffusion >>
rect 355 301 356 302 
<< pdiffusion >>
rect 356 301 357 302 
<< pdiffusion >>
rect 357 301 358 302 
<< pdiffusion >>
rect 358 301 359 302 
<< pdiffusion >>
rect 359 301 360 302 
<< pdiffusion >>
rect 372 301 373 302 
<< pdiffusion >>
rect 373 301 374 302 
<< pdiffusion >>
rect 374 301 375 302 
<< pdiffusion >>
rect 375 301 376 302 
<< pdiffusion >>
rect 376 301 377 302 
<< pdiffusion >>
rect 377 301 378 302 
<< pdiffusion >>
rect 390 301 391 302 
<< pdiffusion >>
rect 391 301 392 302 
<< pdiffusion >>
rect 392 301 393 302 
<< pdiffusion >>
rect 393 301 394 302 
<< pdiffusion >>
rect 394 301 395 302 
<< pdiffusion >>
rect 395 301 396 302 
<< pdiffusion >>
rect 408 301 409 302 
<< pdiffusion >>
rect 409 301 410 302 
<< pdiffusion >>
rect 410 301 411 302 
<< pdiffusion >>
rect 411 301 412 302 
<< pdiffusion >>
rect 412 301 413 302 
<< pdiffusion >>
rect 413 301 414 302 
<< pdiffusion >>
rect 426 301 427 302 
<< pdiffusion >>
rect 427 301 428 302 
<< pdiffusion >>
rect 428 301 429 302 
<< pdiffusion >>
rect 429 301 430 302 
<< pdiffusion >>
rect 430 301 431 302 
<< pdiffusion >>
rect 431 301 432 302 
<< pdiffusion >>
rect 444 301 445 302 
<< pdiffusion >>
rect 445 301 446 302 
<< pdiffusion >>
rect 446 301 447 302 
<< pdiffusion >>
rect 447 301 448 302 
<< pdiffusion >>
rect 448 301 449 302 
<< pdiffusion >>
rect 449 301 450 302 
<< pdiffusion >>
rect 12 302 13 303 
<< pdiffusion >>
rect 13 302 14 303 
<< pdiffusion >>
rect 14 302 15 303 
<< pdiffusion >>
rect 15 302 16 303 
<< pdiffusion >>
rect 16 302 17 303 
<< pdiffusion >>
rect 17 302 18 303 
<< pdiffusion >>
rect 30 302 31 303 
<< pdiffusion >>
rect 31 302 32 303 
<< pdiffusion >>
rect 32 302 33 303 
<< pdiffusion >>
rect 33 302 34 303 
<< pdiffusion >>
rect 34 302 35 303 
<< pdiffusion >>
rect 35 302 36 303 
<< pdiffusion >>
rect 48 302 49 303 
<< pdiffusion >>
rect 49 302 50 303 
<< pdiffusion >>
rect 50 302 51 303 
<< pdiffusion >>
rect 51 302 52 303 
<< pdiffusion >>
rect 52 302 53 303 
<< pdiffusion >>
rect 53 302 54 303 
<< m1 >>
rect 55 302 56 303 
<< m1 >>
rect 64 302 65 303 
<< pdiffusion >>
rect 66 302 67 303 
<< pdiffusion >>
rect 67 302 68 303 
<< pdiffusion >>
rect 68 302 69 303 
<< pdiffusion >>
rect 69 302 70 303 
<< pdiffusion >>
rect 70 302 71 303 
<< pdiffusion >>
rect 71 302 72 303 
<< pdiffusion >>
rect 84 302 85 303 
<< pdiffusion >>
rect 85 302 86 303 
<< pdiffusion >>
rect 86 302 87 303 
<< pdiffusion >>
rect 87 302 88 303 
<< pdiffusion >>
rect 88 302 89 303 
<< pdiffusion >>
rect 89 302 90 303 
<< m1 >>
rect 91 302 92 303 
<< pdiffusion >>
rect 102 302 103 303 
<< pdiffusion >>
rect 103 302 104 303 
<< pdiffusion >>
rect 104 302 105 303 
<< pdiffusion >>
rect 105 302 106 303 
<< pdiffusion >>
rect 106 302 107 303 
<< pdiffusion >>
rect 107 302 108 303 
<< pdiffusion >>
rect 120 302 121 303 
<< pdiffusion >>
rect 121 302 122 303 
<< pdiffusion >>
rect 122 302 123 303 
<< pdiffusion >>
rect 123 302 124 303 
<< pdiffusion >>
rect 124 302 125 303 
<< pdiffusion >>
rect 125 302 126 303 
<< pdiffusion >>
rect 138 302 139 303 
<< pdiffusion >>
rect 139 302 140 303 
<< pdiffusion >>
rect 140 302 141 303 
<< pdiffusion >>
rect 141 302 142 303 
<< pdiffusion >>
rect 142 302 143 303 
<< pdiffusion >>
rect 143 302 144 303 
<< pdiffusion >>
rect 156 302 157 303 
<< pdiffusion >>
rect 157 302 158 303 
<< pdiffusion >>
rect 158 302 159 303 
<< pdiffusion >>
rect 159 302 160 303 
<< pdiffusion >>
rect 160 302 161 303 
<< pdiffusion >>
rect 161 302 162 303 
<< m1 >>
rect 163 302 164 303 
<< pdiffusion >>
rect 174 302 175 303 
<< pdiffusion >>
rect 175 302 176 303 
<< pdiffusion >>
rect 176 302 177 303 
<< pdiffusion >>
rect 177 302 178 303 
<< pdiffusion >>
rect 178 302 179 303 
<< pdiffusion >>
rect 179 302 180 303 
<< pdiffusion >>
rect 192 302 193 303 
<< pdiffusion >>
rect 193 302 194 303 
<< pdiffusion >>
rect 194 302 195 303 
<< pdiffusion >>
rect 195 302 196 303 
<< pdiffusion >>
rect 196 302 197 303 
<< pdiffusion >>
rect 197 302 198 303 
<< m1 >>
rect 206 302 207 303 
<< m1 >>
rect 208 302 209 303 
<< m2 >>
rect 208 302 209 303 
<< pdiffusion >>
rect 210 302 211 303 
<< pdiffusion >>
rect 211 302 212 303 
<< pdiffusion >>
rect 212 302 213 303 
<< pdiffusion >>
rect 213 302 214 303 
<< pdiffusion >>
rect 214 302 215 303 
<< pdiffusion >>
rect 215 302 216 303 
<< m1 >>
rect 217 302 218 303 
<< m1 >>
rect 226 302 227 303 
<< pdiffusion >>
rect 228 302 229 303 
<< pdiffusion >>
rect 229 302 230 303 
<< pdiffusion >>
rect 230 302 231 303 
<< pdiffusion >>
rect 231 302 232 303 
<< pdiffusion >>
rect 232 302 233 303 
<< pdiffusion >>
rect 233 302 234 303 
<< m1 >>
rect 235 302 236 303 
<< m1 >>
rect 237 302 238 303 
<< pdiffusion >>
rect 246 302 247 303 
<< pdiffusion >>
rect 247 302 248 303 
<< pdiffusion >>
rect 248 302 249 303 
<< pdiffusion >>
rect 249 302 250 303 
<< pdiffusion >>
rect 250 302 251 303 
<< pdiffusion >>
rect 251 302 252 303 
<< m1 >>
rect 257 302 258 303 
<< pdiffusion >>
rect 264 302 265 303 
<< pdiffusion >>
rect 265 302 266 303 
<< pdiffusion >>
rect 266 302 267 303 
<< pdiffusion >>
rect 267 302 268 303 
<< pdiffusion >>
rect 268 302 269 303 
<< pdiffusion >>
rect 269 302 270 303 
<< m1 >>
rect 271 302 272 303 
<< m1 >>
rect 280 302 281 303 
<< pdiffusion >>
rect 282 302 283 303 
<< pdiffusion >>
rect 283 302 284 303 
<< pdiffusion >>
rect 284 302 285 303 
<< pdiffusion >>
rect 285 302 286 303 
<< pdiffusion >>
rect 286 302 287 303 
<< pdiffusion >>
rect 287 302 288 303 
<< m1 >>
rect 289 302 290 303 
<< pdiffusion >>
rect 300 302 301 303 
<< pdiffusion >>
rect 301 302 302 303 
<< pdiffusion >>
rect 302 302 303 303 
<< pdiffusion >>
rect 303 302 304 303 
<< pdiffusion >>
rect 304 302 305 303 
<< pdiffusion >>
rect 305 302 306 303 
<< m1 >>
rect 307 302 308 303 
<< pdiffusion >>
rect 318 302 319 303 
<< pdiffusion >>
rect 319 302 320 303 
<< pdiffusion >>
rect 320 302 321 303 
<< pdiffusion >>
rect 321 302 322 303 
<< pdiffusion >>
rect 322 302 323 303 
<< pdiffusion >>
rect 323 302 324 303 
<< pdiffusion >>
rect 336 302 337 303 
<< pdiffusion >>
rect 337 302 338 303 
<< pdiffusion >>
rect 338 302 339 303 
<< pdiffusion >>
rect 339 302 340 303 
<< pdiffusion >>
rect 340 302 341 303 
<< pdiffusion >>
rect 341 302 342 303 
<< m1 >>
rect 352 302 353 303 
<< pdiffusion >>
rect 354 302 355 303 
<< pdiffusion >>
rect 355 302 356 303 
<< pdiffusion >>
rect 356 302 357 303 
<< pdiffusion >>
rect 357 302 358 303 
<< pdiffusion >>
rect 358 302 359 303 
<< pdiffusion >>
rect 359 302 360 303 
<< pdiffusion >>
rect 372 302 373 303 
<< pdiffusion >>
rect 373 302 374 303 
<< pdiffusion >>
rect 374 302 375 303 
<< pdiffusion >>
rect 375 302 376 303 
<< pdiffusion >>
rect 376 302 377 303 
<< pdiffusion >>
rect 377 302 378 303 
<< pdiffusion >>
rect 390 302 391 303 
<< pdiffusion >>
rect 391 302 392 303 
<< pdiffusion >>
rect 392 302 393 303 
<< pdiffusion >>
rect 393 302 394 303 
<< pdiffusion >>
rect 394 302 395 303 
<< pdiffusion >>
rect 395 302 396 303 
<< pdiffusion >>
rect 408 302 409 303 
<< pdiffusion >>
rect 409 302 410 303 
<< pdiffusion >>
rect 410 302 411 303 
<< pdiffusion >>
rect 411 302 412 303 
<< pdiffusion >>
rect 412 302 413 303 
<< pdiffusion >>
rect 413 302 414 303 
<< pdiffusion >>
rect 426 302 427 303 
<< pdiffusion >>
rect 427 302 428 303 
<< pdiffusion >>
rect 428 302 429 303 
<< pdiffusion >>
rect 429 302 430 303 
<< pdiffusion >>
rect 430 302 431 303 
<< pdiffusion >>
rect 431 302 432 303 
<< pdiffusion >>
rect 444 302 445 303 
<< pdiffusion >>
rect 445 302 446 303 
<< pdiffusion >>
rect 446 302 447 303 
<< pdiffusion >>
rect 447 302 448 303 
<< pdiffusion >>
rect 448 302 449 303 
<< pdiffusion >>
rect 449 302 450 303 
<< pdiffusion >>
rect 12 303 13 304 
<< pdiffusion >>
rect 13 303 14 304 
<< pdiffusion >>
rect 14 303 15 304 
<< pdiffusion >>
rect 15 303 16 304 
<< pdiffusion >>
rect 16 303 17 304 
<< pdiffusion >>
rect 17 303 18 304 
<< pdiffusion >>
rect 30 303 31 304 
<< pdiffusion >>
rect 31 303 32 304 
<< pdiffusion >>
rect 32 303 33 304 
<< pdiffusion >>
rect 33 303 34 304 
<< pdiffusion >>
rect 34 303 35 304 
<< pdiffusion >>
rect 35 303 36 304 
<< pdiffusion >>
rect 48 303 49 304 
<< pdiffusion >>
rect 49 303 50 304 
<< pdiffusion >>
rect 50 303 51 304 
<< pdiffusion >>
rect 51 303 52 304 
<< pdiffusion >>
rect 52 303 53 304 
<< pdiffusion >>
rect 53 303 54 304 
<< m1 >>
rect 55 303 56 304 
<< m1 >>
rect 64 303 65 304 
<< pdiffusion >>
rect 66 303 67 304 
<< pdiffusion >>
rect 67 303 68 304 
<< pdiffusion >>
rect 68 303 69 304 
<< pdiffusion >>
rect 69 303 70 304 
<< pdiffusion >>
rect 70 303 71 304 
<< pdiffusion >>
rect 71 303 72 304 
<< pdiffusion >>
rect 84 303 85 304 
<< pdiffusion >>
rect 85 303 86 304 
<< pdiffusion >>
rect 86 303 87 304 
<< pdiffusion >>
rect 87 303 88 304 
<< pdiffusion >>
rect 88 303 89 304 
<< pdiffusion >>
rect 89 303 90 304 
<< m1 >>
rect 91 303 92 304 
<< pdiffusion >>
rect 102 303 103 304 
<< pdiffusion >>
rect 103 303 104 304 
<< pdiffusion >>
rect 104 303 105 304 
<< pdiffusion >>
rect 105 303 106 304 
<< pdiffusion >>
rect 106 303 107 304 
<< pdiffusion >>
rect 107 303 108 304 
<< pdiffusion >>
rect 120 303 121 304 
<< pdiffusion >>
rect 121 303 122 304 
<< pdiffusion >>
rect 122 303 123 304 
<< pdiffusion >>
rect 123 303 124 304 
<< pdiffusion >>
rect 124 303 125 304 
<< pdiffusion >>
rect 125 303 126 304 
<< pdiffusion >>
rect 138 303 139 304 
<< pdiffusion >>
rect 139 303 140 304 
<< pdiffusion >>
rect 140 303 141 304 
<< pdiffusion >>
rect 141 303 142 304 
<< pdiffusion >>
rect 142 303 143 304 
<< pdiffusion >>
rect 143 303 144 304 
<< pdiffusion >>
rect 156 303 157 304 
<< pdiffusion >>
rect 157 303 158 304 
<< pdiffusion >>
rect 158 303 159 304 
<< pdiffusion >>
rect 159 303 160 304 
<< pdiffusion >>
rect 160 303 161 304 
<< pdiffusion >>
rect 161 303 162 304 
<< m1 >>
rect 163 303 164 304 
<< pdiffusion >>
rect 174 303 175 304 
<< pdiffusion >>
rect 175 303 176 304 
<< pdiffusion >>
rect 176 303 177 304 
<< pdiffusion >>
rect 177 303 178 304 
<< pdiffusion >>
rect 178 303 179 304 
<< pdiffusion >>
rect 179 303 180 304 
<< pdiffusion >>
rect 192 303 193 304 
<< pdiffusion >>
rect 193 303 194 304 
<< pdiffusion >>
rect 194 303 195 304 
<< pdiffusion >>
rect 195 303 196 304 
<< pdiffusion >>
rect 196 303 197 304 
<< pdiffusion >>
rect 197 303 198 304 
<< m1 >>
rect 206 303 207 304 
<< m1 >>
rect 208 303 209 304 
<< m2 >>
rect 208 303 209 304 
<< pdiffusion >>
rect 210 303 211 304 
<< pdiffusion >>
rect 211 303 212 304 
<< pdiffusion >>
rect 212 303 213 304 
<< pdiffusion >>
rect 213 303 214 304 
<< pdiffusion >>
rect 214 303 215 304 
<< pdiffusion >>
rect 215 303 216 304 
<< m1 >>
rect 217 303 218 304 
<< m1 >>
rect 226 303 227 304 
<< pdiffusion >>
rect 228 303 229 304 
<< pdiffusion >>
rect 229 303 230 304 
<< pdiffusion >>
rect 230 303 231 304 
<< pdiffusion >>
rect 231 303 232 304 
<< pdiffusion >>
rect 232 303 233 304 
<< pdiffusion >>
rect 233 303 234 304 
<< m1 >>
rect 235 303 236 304 
<< m1 >>
rect 237 303 238 304 
<< pdiffusion >>
rect 246 303 247 304 
<< pdiffusion >>
rect 247 303 248 304 
<< pdiffusion >>
rect 248 303 249 304 
<< pdiffusion >>
rect 249 303 250 304 
<< pdiffusion >>
rect 250 303 251 304 
<< pdiffusion >>
rect 251 303 252 304 
<< m1 >>
rect 257 303 258 304 
<< pdiffusion >>
rect 264 303 265 304 
<< pdiffusion >>
rect 265 303 266 304 
<< pdiffusion >>
rect 266 303 267 304 
<< pdiffusion >>
rect 267 303 268 304 
<< pdiffusion >>
rect 268 303 269 304 
<< pdiffusion >>
rect 269 303 270 304 
<< m1 >>
rect 271 303 272 304 
<< m1 >>
rect 280 303 281 304 
<< pdiffusion >>
rect 282 303 283 304 
<< pdiffusion >>
rect 283 303 284 304 
<< pdiffusion >>
rect 284 303 285 304 
<< pdiffusion >>
rect 285 303 286 304 
<< pdiffusion >>
rect 286 303 287 304 
<< pdiffusion >>
rect 287 303 288 304 
<< m1 >>
rect 289 303 290 304 
<< pdiffusion >>
rect 300 303 301 304 
<< pdiffusion >>
rect 301 303 302 304 
<< pdiffusion >>
rect 302 303 303 304 
<< pdiffusion >>
rect 303 303 304 304 
<< pdiffusion >>
rect 304 303 305 304 
<< pdiffusion >>
rect 305 303 306 304 
<< m1 >>
rect 307 303 308 304 
<< pdiffusion >>
rect 318 303 319 304 
<< pdiffusion >>
rect 319 303 320 304 
<< pdiffusion >>
rect 320 303 321 304 
<< pdiffusion >>
rect 321 303 322 304 
<< pdiffusion >>
rect 322 303 323 304 
<< pdiffusion >>
rect 323 303 324 304 
<< pdiffusion >>
rect 336 303 337 304 
<< pdiffusion >>
rect 337 303 338 304 
<< pdiffusion >>
rect 338 303 339 304 
<< pdiffusion >>
rect 339 303 340 304 
<< pdiffusion >>
rect 340 303 341 304 
<< pdiffusion >>
rect 341 303 342 304 
<< m1 >>
rect 352 303 353 304 
<< pdiffusion >>
rect 354 303 355 304 
<< pdiffusion >>
rect 355 303 356 304 
<< pdiffusion >>
rect 356 303 357 304 
<< pdiffusion >>
rect 357 303 358 304 
<< pdiffusion >>
rect 358 303 359 304 
<< pdiffusion >>
rect 359 303 360 304 
<< pdiffusion >>
rect 372 303 373 304 
<< pdiffusion >>
rect 373 303 374 304 
<< pdiffusion >>
rect 374 303 375 304 
<< pdiffusion >>
rect 375 303 376 304 
<< pdiffusion >>
rect 376 303 377 304 
<< pdiffusion >>
rect 377 303 378 304 
<< pdiffusion >>
rect 390 303 391 304 
<< pdiffusion >>
rect 391 303 392 304 
<< pdiffusion >>
rect 392 303 393 304 
<< pdiffusion >>
rect 393 303 394 304 
<< pdiffusion >>
rect 394 303 395 304 
<< pdiffusion >>
rect 395 303 396 304 
<< pdiffusion >>
rect 408 303 409 304 
<< pdiffusion >>
rect 409 303 410 304 
<< pdiffusion >>
rect 410 303 411 304 
<< pdiffusion >>
rect 411 303 412 304 
<< pdiffusion >>
rect 412 303 413 304 
<< pdiffusion >>
rect 413 303 414 304 
<< pdiffusion >>
rect 426 303 427 304 
<< pdiffusion >>
rect 427 303 428 304 
<< pdiffusion >>
rect 428 303 429 304 
<< pdiffusion >>
rect 429 303 430 304 
<< pdiffusion >>
rect 430 303 431 304 
<< pdiffusion >>
rect 431 303 432 304 
<< pdiffusion >>
rect 444 303 445 304 
<< pdiffusion >>
rect 445 303 446 304 
<< pdiffusion >>
rect 446 303 447 304 
<< pdiffusion >>
rect 447 303 448 304 
<< pdiffusion >>
rect 448 303 449 304 
<< pdiffusion >>
rect 449 303 450 304 
<< pdiffusion >>
rect 12 304 13 305 
<< pdiffusion >>
rect 13 304 14 305 
<< pdiffusion >>
rect 14 304 15 305 
<< pdiffusion >>
rect 15 304 16 305 
<< pdiffusion >>
rect 16 304 17 305 
<< pdiffusion >>
rect 17 304 18 305 
<< pdiffusion >>
rect 30 304 31 305 
<< pdiffusion >>
rect 31 304 32 305 
<< pdiffusion >>
rect 32 304 33 305 
<< pdiffusion >>
rect 33 304 34 305 
<< pdiffusion >>
rect 34 304 35 305 
<< pdiffusion >>
rect 35 304 36 305 
<< pdiffusion >>
rect 48 304 49 305 
<< pdiffusion >>
rect 49 304 50 305 
<< pdiffusion >>
rect 50 304 51 305 
<< pdiffusion >>
rect 51 304 52 305 
<< pdiffusion >>
rect 52 304 53 305 
<< pdiffusion >>
rect 53 304 54 305 
<< m1 >>
rect 55 304 56 305 
<< m1 >>
rect 64 304 65 305 
<< pdiffusion >>
rect 66 304 67 305 
<< pdiffusion >>
rect 67 304 68 305 
<< pdiffusion >>
rect 68 304 69 305 
<< pdiffusion >>
rect 69 304 70 305 
<< pdiffusion >>
rect 70 304 71 305 
<< pdiffusion >>
rect 71 304 72 305 
<< pdiffusion >>
rect 84 304 85 305 
<< pdiffusion >>
rect 85 304 86 305 
<< pdiffusion >>
rect 86 304 87 305 
<< pdiffusion >>
rect 87 304 88 305 
<< pdiffusion >>
rect 88 304 89 305 
<< pdiffusion >>
rect 89 304 90 305 
<< m1 >>
rect 91 304 92 305 
<< pdiffusion >>
rect 102 304 103 305 
<< pdiffusion >>
rect 103 304 104 305 
<< pdiffusion >>
rect 104 304 105 305 
<< pdiffusion >>
rect 105 304 106 305 
<< pdiffusion >>
rect 106 304 107 305 
<< pdiffusion >>
rect 107 304 108 305 
<< pdiffusion >>
rect 120 304 121 305 
<< pdiffusion >>
rect 121 304 122 305 
<< pdiffusion >>
rect 122 304 123 305 
<< pdiffusion >>
rect 123 304 124 305 
<< pdiffusion >>
rect 124 304 125 305 
<< pdiffusion >>
rect 125 304 126 305 
<< pdiffusion >>
rect 138 304 139 305 
<< pdiffusion >>
rect 139 304 140 305 
<< pdiffusion >>
rect 140 304 141 305 
<< pdiffusion >>
rect 141 304 142 305 
<< pdiffusion >>
rect 142 304 143 305 
<< pdiffusion >>
rect 143 304 144 305 
<< pdiffusion >>
rect 156 304 157 305 
<< pdiffusion >>
rect 157 304 158 305 
<< pdiffusion >>
rect 158 304 159 305 
<< pdiffusion >>
rect 159 304 160 305 
<< pdiffusion >>
rect 160 304 161 305 
<< pdiffusion >>
rect 161 304 162 305 
<< m1 >>
rect 163 304 164 305 
<< pdiffusion >>
rect 174 304 175 305 
<< pdiffusion >>
rect 175 304 176 305 
<< pdiffusion >>
rect 176 304 177 305 
<< pdiffusion >>
rect 177 304 178 305 
<< pdiffusion >>
rect 178 304 179 305 
<< pdiffusion >>
rect 179 304 180 305 
<< pdiffusion >>
rect 192 304 193 305 
<< pdiffusion >>
rect 193 304 194 305 
<< pdiffusion >>
rect 194 304 195 305 
<< pdiffusion >>
rect 195 304 196 305 
<< pdiffusion >>
rect 196 304 197 305 
<< pdiffusion >>
rect 197 304 198 305 
<< m1 >>
rect 206 304 207 305 
<< m1 >>
rect 208 304 209 305 
<< m2 >>
rect 208 304 209 305 
<< pdiffusion >>
rect 210 304 211 305 
<< pdiffusion >>
rect 211 304 212 305 
<< pdiffusion >>
rect 212 304 213 305 
<< pdiffusion >>
rect 213 304 214 305 
<< pdiffusion >>
rect 214 304 215 305 
<< pdiffusion >>
rect 215 304 216 305 
<< m1 >>
rect 217 304 218 305 
<< m1 >>
rect 226 304 227 305 
<< pdiffusion >>
rect 228 304 229 305 
<< pdiffusion >>
rect 229 304 230 305 
<< pdiffusion >>
rect 230 304 231 305 
<< pdiffusion >>
rect 231 304 232 305 
<< pdiffusion >>
rect 232 304 233 305 
<< pdiffusion >>
rect 233 304 234 305 
<< m1 >>
rect 235 304 236 305 
<< m1 >>
rect 237 304 238 305 
<< pdiffusion >>
rect 246 304 247 305 
<< pdiffusion >>
rect 247 304 248 305 
<< pdiffusion >>
rect 248 304 249 305 
<< pdiffusion >>
rect 249 304 250 305 
<< pdiffusion >>
rect 250 304 251 305 
<< pdiffusion >>
rect 251 304 252 305 
<< m1 >>
rect 257 304 258 305 
<< pdiffusion >>
rect 264 304 265 305 
<< pdiffusion >>
rect 265 304 266 305 
<< pdiffusion >>
rect 266 304 267 305 
<< pdiffusion >>
rect 267 304 268 305 
<< pdiffusion >>
rect 268 304 269 305 
<< pdiffusion >>
rect 269 304 270 305 
<< m1 >>
rect 271 304 272 305 
<< m1 >>
rect 280 304 281 305 
<< pdiffusion >>
rect 282 304 283 305 
<< pdiffusion >>
rect 283 304 284 305 
<< pdiffusion >>
rect 284 304 285 305 
<< pdiffusion >>
rect 285 304 286 305 
<< pdiffusion >>
rect 286 304 287 305 
<< pdiffusion >>
rect 287 304 288 305 
<< m1 >>
rect 289 304 290 305 
<< pdiffusion >>
rect 300 304 301 305 
<< pdiffusion >>
rect 301 304 302 305 
<< pdiffusion >>
rect 302 304 303 305 
<< pdiffusion >>
rect 303 304 304 305 
<< pdiffusion >>
rect 304 304 305 305 
<< pdiffusion >>
rect 305 304 306 305 
<< m1 >>
rect 307 304 308 305 
<< pdiffusion >>
rect 318 304 319 305 
<< pdiffusion >>
rect 319 304 320 305 
<< pdiffusion >>
rect 320 304 321 305 
<< pdiffusion >>
rect 321 304 322 305 
<< pdiffusion >>
rect 322 304 323 305 
<< pdiffusion >>
rect 323 304 324 305 
<< pdiffusion >>
rect 336 304 337 305 
<< pdiffusion >>
rect 337 304 338 305 
<< pdiffusion >>
rect 338 304 339 305 
<< pdiffusion >>
rect 339 304 340 305 
<< pdiffusion >>
rect 340 304 341 305 
<< pdiffusion >>
rect 341 304 342 305 
<< m1 >>
rect 352 304 353 305 
<< pdiffusion >>
rect 354 304 355 305 
<< pdiffusion >>
rect 355 304 356 305 
<< pdiffusion >>
rect 356 304 357 305 
<< pdiffusion >>
rect 357 304 358 305 
<< pdiffusion >>
rect 358 304 359 305 
<< pdiffusion >>
rect 359 304 360 305 
<< pdiffusion >>
rect 372 304 373 305 
<< pdiffusion >>
rect 373 304 374 305 
<< pdiffusion >>
rect 374 304 375 305 
<< pdiffusion >>
rect 375 304 376 305 
<< pdiffusion >>
rect 376 304 377 305 
<< pdiffusion >>
rect 377 304 378 305 
<< pdiffusion >>
rect 390 304 391 305 
<< pdiffusion >>
rect 391 304 392 305 
<< pdiffusion >>
rect 392 304 393 305 
<< pdiffusion >>
rect 393 304 394 305 
<< pdiffusion >>
rect 394 304 395 305 
<< pdiffusion >>
rect 395 304 396 305 
<< pdiffusion >>
rect 408 304 409 305 
<< pdiffusion >>
rect 409 304 410 305 
<< pdiffusion >>
rect 410 304 411 305 
<< pdiffusion >>
rect 411 304 412 305 
<< pdiffusion >>
rect 412 304 413 305 
<< pdiffusion >>
rect 413 304 414 305 
<< pdiffusion >>
rect 426 304 427 305 
<< pdiffusion >>
rect 427 304 428 305 
<< pdiffusion >>
rect 428 304 429 305 
<< pdiffusion >>
rect 429 304 430 305 
<< pdiffusion >>
rect 430 304 431 305 
<< pdiffusion >>
rect 431 304 432 305 
<< pdiffusion >>
rect 444 304 445 305 
<< pdiffusion >>
rect 445 304 446 305 
<< pdiffusion >>
rect 446 304 447 305 
<< pdiffusion >>
rect 447 304 448 305 
<< pdiffusion >>
rect 448 304 449 305 
<< pdiffusion >>
rect 449 304 450 305 
<< pdiffusion >>
rect 12 305 13 306 
<< pdiffusion >>
rect 13 305 14 306 
<< pdiffusion >>
rect 14 305 15 306 
<< pdiffusion >>
rect 15 305 16 306 
<< pdiffusion >>
rect 16 305 17 306 
<< pdiffusion >>
rect 17 305 18 306 
<< pdiffusion >>
rect 30 305 31 306 
<< pdiffusion >>
rect 31 305 32 306 
<< pdiffusion >>
rect 32 305 33 306 
<< pdiffusion >>
rect 33 305 34 306 
<< pdiffusion >>
rect 34 305 35 306 
<< pdiffusion >>
rect 35 305 36 306 
<< pdiffusion >>
rect 48 305 49 306 
<< pdiffusion >>
rect 49 305 50 306 
<< pdiffusion >>
rect 50 305 51 306 
<< pdiffusion >>
rect 51 305 52 306 
<< pdiffusion >>
rect 52 305 53 306 
<< pdiffusion >>
rect 53 305 54 306 
<< m1 >>
rect 55 305 56 306 
<< m1 >>
rect 64 305 65 306 
<< pdiffusion >>
rect 66 305 67 306 
<< pdiffusion >>
rect 67 305 68 306 
<< pdiffusion >>
rect 68 305 69 306 
<< pdiffusion >>
rect 69 305 70 306 
<< pdiffusion >>
rect 70 305 71 306 
<< pdiffusion >>
rect 71 305 72 306 
<< pdiffusion >>
rect 84 305 85 306 
<< pdiffusion >>
rect 85 305 86 306 
<< pdiffusion >>
rect 86 305 87 306 
<< pdiffusion >>
rect 87 305 88 306 
<< pdiffusion >>
rect 88 305 89 306 
<< pdiffusion >>
rect 89 305 90 306 
<< m1 >>
rect 91 305 92 306 
<< pdiffusion >>
rect 102 305 103 306 
<< pdiffusion >>
rect 103 305 104 306 
<< pdiffusion >>
rect 104 305 105 306 
<< pdiffusion >>
rect 105 305 106 306 
<< pdiffusion >>
rect 106 305 107 306 
<< pdiffusion >>
rect 107 305 108 306 
<< pdiffusion >>
rect 120 305 121 306 
<< pdiffusion >>
rect 121 305 122 306 
<< pdiffusion >>
rect 122 305 123 306 
<< pdiffusion >>
rect 123 305 124 306 
<< m1 >>
rect 124 305 125 306 
<< pdiffusion >>
rect 124 305 125 306 
<< pdiffusion >>
rect 125 305 126 306 
<< pdiffusion >>
rect 138 305 139 306 
<< pdiffusion >>
rect 139 305 140 306 
<< pdiffusion >>
rect 140 305 141 306 
<< pdiffusion >>
rect 141 305 142 306 
<< pdiffusion >>
rect 142 305 143 306 
<< pdiffusion >>
rect 143 305 144 306 
<< pdiffusion >>
rect 156 305 157 306 
<< pdiffusion >>
rect 157 305 158 306 
<< pdiffusion >>
rect 158 305 159 306 
<< pdiffusion >>
rect 159 305 160 306 
<< pdiffusion >>
rect 160 305 161 306 
<< pdiffusion >>
rect 161 305 162 306 
<< m1 >>
rect 163 305 164 306 
<< pdiffusion >>
rect 174 305 175 306 
<< pdiffusion >>
rect 175 305 176 306 
<< pdiffusion >>
rect 176 305 177 306 
<< pdiffusion >>
rect 177 305 178 306 
<< pdiffusion >>
rect 178 305 179 306 
<< pdiffusion >>
rect 179 305 180 306 
<< pdiffusion >>
rect 192 305 193 306 
<< pdiffusion >>
rect 193 305 194 306 
<< pdiffusion >>
rect 194 305 195 306 
<< pdiffusion >>
rect 195 305 196 306 
<< pdiffusion >>
rect 196 305 197 306 
<< pdiffusion >>
rect 197 305 198 306 
<< m1 >>
rect 206 305 207 306 
<< m1 >>
rect 208 305 209 306 
<< m2 >>
rect 208 305 209 306 
<< pdiffusion >>
rect 210 305 211 306 
<< pdiffusion >>
rect 211 305 212 306 
<< pdiffusion >>
rect 212 305 213 306 
<< pdiffusion >>
rect 213 305 214 306 
<< pdiffusion >>
rect 214 305 215 306 
<< pdiffusion >>
rect 215 305 216 306 
<< m1 >>
rect 217 305 218 306 
<< m1 >>
rect 226 305 227 306 
<< pdiffusion >>
rect 228 305 229 306 
<< pdiffusion >>
rect 229 305 230 306 
<< pdiffusion >>
rect 230 305 231 306 
<< pdiffusion >>
rect 231 305 232 306 
<< pdiffusion >>
rect 232 305 233 306 
<< pdiffusion >>
rect 233 305 234 306 
<< m1 >>
rect 235 305 236 306 
<< m1 >>
rect 237 305 238 306 
<< pdiffusion >>
rect 246 305 247 306 
<< pdiffusion >>
rect 247 305 248 306 
<< pdiffusion >>
rect 248 305 249 306 
<< pdiffusion >>
rect 249 305 250 306 
<< pdiffusion >>
rect 250 305 251 306 
<< pdiffusion >>
rect 251 305 252 306 
<< m1 >>
rect 257 305 258 306 
<< pdiffusion >>
rect 264 305 265 306 
<< pdiffusion >>
rect 265 305 266 306 
<< pdiffusion >>
rect 266 305 267 306 
<< pdiffusion >>
rect 267 305 268 306 
<< pdiffusion >>
rect 268 305 269 306 
<< pdiffusion >>
rect 269 305 270 306 
<< m1 >>
rect 271 305 272 306 
<< m1 >>
rect 280 305 281 306 
<< pdiffusion >>
rect 282 305 283 306 
<< pdiffusion >>
rect 283 305 284 306 
<< pdiffusion >>
rect 284 305 285 306 
<< pdiffusion >>
rect 285 305 286 306 
<< pdiffusion >>
rect 286 305 287 306 
<< pdiffusion >>
rect 287 305 288 306 
<< m1 >>
rect 289 305 290 306 
<< pdiffusion >>
rect 300 305 301 306 
<< pdiffusion >>
rect 301 305 302 306 
<< pdiffusion >>
rect 302 305 303 306 
<< pdiffusion >>
rect 303 305 304 306 
<< pdiffusion >>
rect 304 305 305 306 
<< pdiffusion >>
rect 305 305 306 306 
<< m1 >>
rect 307 305 308 306 
<< pdiffusion >>
rect 318 305 319 306 
<< pdiffusion >>
rect 319 305 320 306 
<< pdiffusion >>
rect 320 305 321 306 
<< pdiffusion >>
rect 321 305 322 306 
<< pdiffusion >>
rect 322 305 323 306 
<< pdiffusion >>
rect 323 305 324 306 
<< pdiffusion >>
rect 336 305 337 306 
<< m1 >>
rect 337 305 338 306 
<< pdiffusion >>
rect 337 305 338 306 
<< pdiffusion >>
rect 338 305 339 306 
<< pdiffusion >>
rect 339 305 340 306 
<< pdiffusion >>
rect 340 305 341 306 
<< pdiffusion >>
rect 341 305 342 306 
<< m1 >>
rect 352 305 353 306 
<< pdiffusion >>
rect 354 305 355 306 
<< pdiffusion >>
rect 355 305 356 306 
<< pdiffusion >>
rect 356 305 357 306 
<< pdiffusion >>
rect 357 305 358 306 
<< pdiffusion >>
rect 358 305 359 306 
<< pdiffusion >>
rect 359 305 360 306 
<< pdiffusion >>
rect 372 305 373 306 
<< m1 >>
rect 373 305 374 306 
<< pdiffusion >>
rect 373 305 374 306 
<< pdiffusion >>
rect 374 305 375 306 
<< pdiffusion >>
rect 375 305 376 306 
<< pdiffusion >>
rect 376 305 377 306 
<< pdiffusion >>
rect 377 305 378 306 
<< pdiffusion >>
rect 390 305 391 306 
<< pdiffusion >>
rect 391 305 392 306 
<< pdiffusion >>
rect 392 305 393 306 
<< pdiffusion >>
rect 393 305 394 306 
<< pdiffusion >>
rect 394 305 395 306 
<< pdiffusion >>
rect 395 305 396 306 
<< pdiffusion >>
rect 408 305 409 306 
<< pdiffusion >>
rect 409 305 410 306 
<< pdiffusion >>
rect 410 305 411 306 
<< pdiffusion >>
rect 411 305 412 306 
<< pdiffusion >>
rect 412 305 413 306 
<< pdiffusion >>
rect 413 305 414 306 
<< pdiffusion >>
rect 426 305 427 306 
<< pdiffusion >>
rect 427 305 428 306 
<< pdiffusion >>
rect 428 305 429 306 
<< pdiffusion >>
rect 429 305 430 306 
<< pdiffusion >>
rect 430 305 431 306 
<< pdiffusion >>
rect 431 305 432 306 
<< pdiffusion >>
rect 444 305 445 306 
<< pdiffusion >>
rect 445 305 446 306 
<< pdiffusion >>
rect 446 305 447 306 
<< pdiffusion >>
rect 447 305 448 306 
<< pdiffusion >>
rect 448 305 449 306 
<< pdiffusion >>
rect 449 305 450 306 
<< m1 >>
rect 55 306 56 307 
<< m1 >>
rect 64 306 65 307 
<< m1 >>
rect 91 306 92 307 
<< m1 >>
rect 124 306 125 307 
<< m1 >>
rect 163 306 164 307 
<< m1 >>
rect 206 306 207 307 
<< m1 >>
rect 208 306 209 307 
<< m2 >>
rect 208 306 209 307 
<< m1 >>
rect 217 306 218 307 
<< m1 >>
rect 226 306 227 307 
<< m1 >>
rect 235 306 236 307 
<< m1 >>
rect 237 306 238 307 
<< m1 >>
rect 257 306 258 307 
<< m1 >>
rect 271 306 272 307 
<< m1 >>
rect 280 306 281 307 
<< m1 >>
rect 289 306 290 307 
<< m1 >>
rect 307 306 308 307 
<< m1 >>
rect 337 306 338 307 
<< m1 >>
rect 352 306 353 307 
<< m1 >>
rect 373 306 374 307 
<< m1 >>
rect 55 307 56 308 
<< m1 >>
rect 64 307 65 308 
<< m1 >>
rect 91 307 92 308 
<< m1 >>
rect 124 307 125 308 
<< m1 >>
rect 163 307 164 308 
<< m1 >>
rect 206 307 207 308 
<< m1 >>
rect 208 307 209 308 
<< m2 >>
rect 208 307 209 308 
<< m1 >>
rect 217 307 218 308 
<< m1 >>
rect 226 307 227 308 
<< m1 >>
rect 235 307 236 308 
<< m1 >>
rect 237 307 238 308 
<< m1 >>
rect 257 307 258 308 
<< m1 >>
rect 271 307 272 308 
<< m1 >>
rect 280 307 281 308 
<< m1 >>
rect 289 307 290 308 
<< m1 >>
rect 307 307 308 308 
<< m1 >>
rect 337 307 338 308 
<< m1 >>
rect 352 307 353 308 
<< m1 >>
rect 373 307 374 308 
<< m1 >>
rect 55 308 56 309 
<< m1 >>
rect 64 308 65 309 
<< m1 >>
rect 91 308 92 309 
<< m1 >>
rect 124 308 125 309 
<< m1 >>
rect 163 308 164 309 
<< m1 >>
rect 206 308 207 309 
<< m1 >>
rect 208 308 209 309 
<< m2 >>
rect 208 308 209 309 
<< m1 >>
rect 217 308 218 309 
<< m1 >>
rect 226 308 227 309 
<< m2 >>
rect 234 308 235 309 
<< m1 >>
rect 235 308 236 309 
<< m2 >>
rect 235 308 236 309 
<< m2 >>
rect 236 308 237 309 
<< m1 >>
rect 237 308 238 309 
<< m2 >>
rect 237 308 238 309 
<< m2c >>
rect 237 308 238 309 
<< m1 >>
rect 237 308 238 309 
<< m2 >>
rect 237 308 238 309 
<< m1 >>
rect 257 308 258 309 
<< m1 >>
rect 271 308 272 309 
<< m1 >>
rect 280 308 281 309 
<< m1 >>
rect 289 308 290 309 
<< m1 >>
rect 307 308 308 309 
<< m1 >>
rect 337 308 338 309 
<< m1 >>
rect 352 308 353 309 
<< m1 >>
rect 373 308 374 309 
<< m1 >>
rect 55 309 56 310 
<< m1 >>
rect 64 309 65 310 
<< m1 >>
rect 91 309 92 310 
<< m1 >>
rect 124 309 125 310 
<< m1 >>
rect 163 309 164 310 
<< m1 >>
rect 206 309 207 310 
<< m1 >>
rect 208 309 209 310 
<< m2 >>
rect 208 309 209 310 
<< m2 >>
rect 209 309 210 310 
<< m1 >>
rect 210 309 211 310 
<< m2 >>
rect 210 309 211 310 
<< m2c >>
rect 210 309 211 310 
<< m1 >>
rect 210 309 211 310 
<< m2 >>
rect 210 309 211 310 
<< m1 >>
rect 217 309 218 310 
<< m1 >>
rect 226 309 227 310 
<< m2 >>
rect 234 309 235 310 
<< m1 >>
rect 235 309 236 310 
<< m1 >>
rect 257 309 258 310 
<< m1 >>
rect 271 309 272 310 
<< m1 >>
rect 280 309 281 310 
<< m1 >>
rect 289 309 290 310 
<< m1 >>
rect 307 309 308 310 
<< m1 >>
rect 337 309 338 310 
<< m1 >>
rect 352 309 353 310 
<< m1 >>
rect 373 309 374 310 
<< m1 >>
rect 55 310 56 311 
<< m1 >>
rect 64 310 65 311 
<< m1 >>
rect 91 310 92 311 
<< m1 >>
rect 118 310 119 311 
<< m1 >>
rect 119 310 120 311 
<< m1 >>
rect 120 310 121 311 
<< m1 >>
rect 121 310 122 311 
<< m1 >>
rect 122 310 123 311 
<< m1 >>
rect 123 310 124 311 
<< m1 >>
rect 124 310 125 311 
<< m1 >>
rect 163 310 164 311 
<< m1 >>
rect 206 310 207 311 
<< m1 >>
rect 208 310 209 311 
<< m1 >>
rect 210 310 211 311 
<< m1 >>
rect 217 310 218 311 
<< m1 >>
rect 226 310 227 311 
<< m2 >>
rect 234 310 235 311 
<< m1 >>
rect 235 310 236 311 
<< m1 >>
rect 236 310 237 311 
<< m1 >>
rect 237 310 238 311 
<< m1 >>
rect 238 310 239 311 
<< m1 >>
rect 239 310 240 311 
<< m1 >>
rect 240 310 241 311 
<< m1 >>
rect 241 310 242 311 
<< m1 >>
rect 242 310 243 311 
<< m1 >>
rect 243 310 244 311 
<< m1 >>
rect 244 310 245 311 
<< m1 >>
rect 245 310 246 311 
<< m1 >>
rect 246 310 247 311 
<< m1 >>
rect 247 310 248 311 
<< m1 >>
rect 257 310 258 311 
<< m1 >>
rect 271 310 272 311 
<< m1 >>
rect 280 310 281 311 
<< m1 >>
rect 289 310 290 311 
<< m1 >>
rect 290 310 291 311 
<< m1 >>
rect 291 310 292 311 
<< m1 >>
rect 292 310 293 311 
<< m1 >>
rect 293 310 294 311 
<< m1 >>
rect 294 310 295 311 
<< m1 >>
rect 295 310 296 311 
<< m1 >>
rect 296 310 297 311 
<< m1 >>
rect 297 310 298 311 
<< m1 >>
rect 298 310 299 311 
<< m1 >>
rect 299 310 300 311 
<< m1 >>
rect 300 310 301 311 
<< m1 >>
rect 301 310 302 311 
<< m1 >>
rect 307 310 308 311 
<< m1 >>
rect 337 310 338 311 
<< m1 >>
rect 338 310 339 311 
<< m1 >>
rect 339 310 340 311 
<< m1 >>
rect 340 310 341 311 
<< m1 >>
rect 341 310 342 311 
<< m1 >>
rect 342 310 343 311 
<< m1 >>
rect 343 310 344 311 
<< m1 >>
rect 344 310 345 311 
<< m1 >>
rect 345 310 346 311 
<< m1 >>
rect 346 310 347 311 
<< m1 >>
rect 347 310 348 311 
<< m1 >>
rect 348 310 349 311 
<< m1 >>
rect 349 310 350 311 
<< m1 >>
rect 350 310 351 311 
<< m2 >>
rect 350 310 351 311 
<< m2c >>
rect 350 310 351 311 
<< m1 >>
rect 350 310 351 311 
<< m2 >>
rect 350 310 351 311 
<< m2 >>
rect 351 310 352 311 
<< m1 >>
rect 352 310 353 311 
<< m2 >>
rect 352 310 353 311 
<< m2 >>
rect 353 310 354 311 
<< m1 >>
rect 354 310 355 311 
<< m2 >>
rect 354 310 355 311 
<< m2c >>
rect 354 310 355 311 
<< m1 >>
rect 354 310 355 311 
<< m2 >>
rect 354 310 355 311 
<< m1 >>
rect 355 310 356 311 
<< m1 >>
rect 356 310 357 311 
<< m1 >>
rect 357 310 358 311 
<< m1 >>
rect 358 310 359 311 
<< m1 >>
rect 359 310 360 311 
<< m1 >>
rect 360 310 361 311 
<< m1 >>
rect 361 310 362 311 
<< m1 >>
rect 362 310 363 311 
<< m1 >>
rect 363 310 364 311 
<< m1 >>
rect 364 310 365 311 
<< m1 >>
rect 365 310 366 311 
<< m1 >>
rect 366 310 367 311 
<< m1 >>
rect 367 310 368 311 
<< m1 >>
rect 368 310 369 311 
<< m1 >>
rect 369 310 370 311 
<< m1 >>
rect 370 310 371 311 
<< m1 >>
rect 371 310 372 311 
<< m1 >>
rect 372 310 373 311 
<< m1 >>
rect 373 310 374 311 
<< m1 >>
rect 55 311 56 312 
<< m1 >>
rect 64 311 65 312 
<< m1 >>
rect 91 311 92 312 
<< m1 >>
rect 118 311 119 312 
<< m1 >>
rect 163 311 164 312 
<< m1 >>
rect 206 311 207 312 
<< m2 >>
rect 206 311 207 312 
<< m2c >>
rect 206 311 207 312 
<< m1 >>
rect 206 311 207 312 
<< m2 >>
rect 206 311 207 312 
<< m1 >>
rect 208 311 209 312 
<< m2 >>
rect 208 311 209 312 
<< m2c >>
rect 208 311 209 312 
<< m1 >>
rect 208 311 209 312 
<< m2 >>
rect 208 311 209 312 
<< m1 >>
rect 210 311 211 312 
<< m1 >>
rect 211 311 212 312 
<< m1 >>
rect 212 311 213 312 
<< m1 >>
rect 213 311 214 312 
<< m2 >>
rect 213 311 214 312 
<< m2c >>
rect 213 311 214 312 
<< m1 >>
rect 213 311 214 312 
<< m2 >>
rect 213 311 214 312 
<< m1 >>
rect 217 311 218 312 
<< m1 >>
rect 226 311 227 312 
<< m1 >>
rect 227 311 228 312 
<< m1 >>
rect 228 311 229 312 
<< m1 >>
rect 229 311 230 312 
<< m1 >>
rect 230 311 231 312 
<< m1 >>
rect 231 311 232 312 
<< m1 >>
rect 232 311 233 312 
<< m2 >>
rect 232 311 233 312 
<< m2c >>
rect 232 311 233 312 
<< m1 >>
rect 232 311 233 312 
<< m2 >>
rect 232 311 233 312 
<< m2 >>
rect 234 311 235 312 
<< m1 >>
rect 247 311 248 312 
<< m1 >>
rect 257 311 258 312 
<< m1 >>
rect 271 311 272 312 
<< m1 >>
rect 280 311 281 312 
<< m1 >>
rect 301 311 302 312 
<< m1 >>
rect 307 311 308 312 
<< m1 >>
rect 352 311 353 312 
<< m1 >>
rect 55 312 56 313 
<< m1 >>
rect 64 312 65 313 
<< m1 >>
rect 91 312 92 313 
<< m1 >>
rect 118 312 119 313 
<< m1 >>
rect 163 312 164 313 
<< m2 >>
rect 206 312 207 313 
<< m2 >>
rect 208 312 209 313 
<< m2 >>
rect 213 312 214 313 
<< m1 >>
rect 217 312 218 313 
<< m2 >>
rect 232 312 233 313 
<< m1 >>
rect 234 312 235 313 
<< m2 >>
rect 234 312 235 313 
<< m2c >>
rect 234 312 235 313 
<< m1 >>
rect 234 312 235 313 
<< m2 >>
rect 234 312 235 313 
<< m1 >>
rect 247 312 248 313 
<< m1 >>
rect 257 312 258 313 
<< m1 >>
rect 271 312 272 313 
<< m1 >>
rect 280 312 281 313 
<< m1 >>
rect 301 312 302 313 
<< m1 >>
rect 307 312 308 313 
<< m1 >>
rect 352 312 353 313 
<< m1 >>
rect 55 313 56 314 
<< m1 >>
rect 64 313 65 314 
<< m1 >>
rect 65 313 66 314 
<< m1 >>
rect 66 313 67 314 
<< m1 >>
rect 67 313 68 314 
<< m1 >>
rect 68 313 69 314 
<< m1 >>
rect 69 313 70 314 
<< m1 >>
rect 70 313 71 314 
<< m1 >>
rect 91 313 92 314 
<< m1 >>
rect 118 313 119 314 
<< m1 >>
rect 163 313 164 314 
<< m1 >>
rect 181 313 182 314 
<< m1 >>
rect 182 313 183 314 
<< m1 >>
rect 183 313 184 314 
<< m1 >>
rect 184 313 185 314 
<< m1 >>
rect 185 313 186 314 
<< m1 >>
rect 186 313 187 314 
<< m1 >>
rect 187 313 188 314 
<< m1 >>
rect 188 313 189 314 
<< m1 >>
rect 189 313 190 314 
<< m1 >>
rect 190 313 191 314 
<< m1 >>
rect 191 313 192 314 
<< m1 >>
rect 192 313 193 314 
<< m1 >>
rect 193 313 194 314 
<< m1 >>
rect 194 313 195 314 
<< m1 >>
rect 195 313 196 314 
<< m1 >>
rect 196 313 197 314 
<< m1 >>
rect 197 313 198 314 
<< m1 >>
rect 198 313 199 314 
<< m1 >>
rect 199 313 200 314 
<< m1 >>
rect 200 313 201 314 
<< m1 >>
rect 201 313 202 314 
<< m1 >>
rect 202 313 203 314 
<< m1 >>
rect 203 313 204 314 
<< m1 >>
rect 204 313 205 314 
<< m1 >>
rect 205 313 206 314 
<< m1 >>
rect 206 313 207 314 
<< m2 >>
rect 206 313 207 314 
<< m1 >>
rect 207 313 208 314 
<< m1 >>
rect 208 313 209 314 
<< m2 >>
rect 208 313 209 314 
<< m1 >>
rect 209 313 210 314 
<< m1 >>
rect 210 313 211 314 
<< m1 >>
rect 211 313 212 314 
<< m1 >>
rect 212 313 213 314 
<< m1 >>
rect 213 313 214 314 
<< m2 >>
rect 213 313 214 314 
<< m1 >>
rect 214 313 215 314 
<< m1 >>
rect 215 313 216 314 
<< m2 >>
rect 215 313 216 314 
<< m2c >>
rect 215 313 216 314 
<< m1 >>
rect 215 313 216 314 
<< m2 >>
rect 215 313 216 314 
<< m2 >>
rect 216 313 217 314 
<< m1 >>
rect 217 313 218 314 
<< m2 >>
rect 217 313 218 314 
<< m2 >>
rect 218 313 219 314 
<< m1 >>
rect 219 313 220 314 
<< m2 >>
rect 219 313 220 314 
<< m2c >>
rect 219 313 220 314 
<< m1 >>
rect 219 313 220 314 
<< m2 >>
rect 219 313 220 314 
<< m1 >>
rect 220 313 221 314 
<< m1 >>
rect 221 313 222 314 
<< m1 >>
rect 222 313 223 314 
<< m1 >>
rect 223 313 224 314 
<< m1 >>
rect 224 313 225 314 
<< m1 >>
rect 225 313 226 314 
<< m1 >>
rect 226 313 227 314 
<< m1 >>
rect 227 313 228 314 
<< m1 >>
rect 228 313 229 314 
<< m1 >>
rect 229 313 230 314 
<< m1 >>
rect 230 313 231 314 
<< m1 >>
rect 231 313 232 314 
<< m1 >>
rect 232 313 233 314 
<< m2 >>
rect 232 313 233 314 
<< m1 >>
rect 233 313 234 314 
<< m1 >>
rect 234 313 235 314 
<< m1 >>
rect 247 313 248 314 
<< m1 >>
rect 257 313 258 314 
<< m1 >>
rect 271 313 272 314 
<< m1 >>
rect 280 313 281 314 
<< m1 >>
rect 301 313 302 314 
<< m1 >>
rect 307 313 308 314 
<< m2 >>
rect 308 313 309 314 
<< m1 >>
rect 309 313 310 314 
<< m2 >>
rect 309 313 310 314 
<< m2c >>
rect 309 313 310 314 
<< m1 >>
rect 309 313 310 314 
<< m2 >>
rect 309 313 310 314 
<< m1 >>
rect 310 313 311 314 
<< m1 >>
rect 311 313 312 314 
<< m1 >>
rect 312 313 313 314 
<< m1 >>
rect 313 313 314 314 
<< m1 >>
rect 314 313 315 314 
<< m1 >>
rect 315 313 316 314 
<< m1 >>
rect 316 313 317 314 
<< m1 >>
rect 317 313 318 314 
<< m1 >>
rect 318 313 319 314 
<< m1 >>
rect 319 313 320 314 
<< m1 >>
rect 320 313 321 314 
<< m1 >>
rect 321 313 322 314 
<< m1 >>
rect 322 313 323 314 
<< m1 >>
rect 323 313 324 314 
<< m1 >>
rect 324 313 325 314 
<< m1 >>
rect 325 313 326 314 
<< m1 >>
rect 352 313 353 314 
<< m1 >>
rect 55 314 56 315 
<< m2 >>
rect 55 314 56 315 
<< m2c >>
rect 55 314 56 315 
<< m1 >>
rect 55 314 56 315 
<< m2 >>
rect 55 314 56 315 
<< m1 >>
rect 70 314 71 315 
<< m1 >>
rect 91 314 92 315 
<< m1 >>
rect 118 314 119 315 
<< m1 >>
rect 163 314 164 315 
<< m1 >>
rect 181 314 182 315 
<< m2 >>
rect 206 314 207 315 
<< m2 >>
rect 208 314 209 315 
<< m2 >>
rect 213 314 214 315 
<< m1 >>
rect 217 314 218 315 
<< m2 >>
rect 232 314 233 315 
<< m2 >>
rect 233 314 234 315 
<< m2 >>
rect 234 314 235 315 
<< m2 >>
rect 235 314 236 315 
<< m1 >>
rect 236 314 237 315 
<< m2 >>
rect 236 314 237 315 
<< m2c >>
rect 236 314 237 315 
<< m1 >>
rect 236 314 237 315 
<< m2 >>
rect 236 314 237 315 
<< m1 >>
rect 237 314 238 315 
<< m1 >>
rect 238 314 239 315 
<< m1 >>
rect 239 314 240 315 
<< m1 >>
rect 240 314 241 315 
<< m1 >>
rect 241 314 242 315 
<< m1 >>
rect 242 314 243 315 
<< m1 >>
rect 243 314 244 315 
<< m1 >>
rect 244 314 245 315 
<< m1 >>
rect 247 314 248 315 
<< m1 >>
rect 257 314 258 315 
<< m1 >>
rect 271 314 272 315 
<< m1 >>
rect 280 314 281 315 
<< m1 >>
rect 301 314 302 315 
<< m1 >>
rect 307 314 308 315 
<< m2 >>
rect 308 314 309 315 
<< m1 >>
rect 325 314 326 315 
<< m2 >>
rect 325 314 326 315 
<< m2c >>
rect 325 314 326 315 
<< m1 >>
rect 325 314 326 315 
<< m2 >>
rect 325 314 326 315 
<< m1 >>
rect 352 314 353 315 
<< m2 >>
rect 55 315 56 316 
<< m1 >>
rect 70 315 71 316 
<< m1 >>
rect 91 315 92 316 
<< m1 >>
rect 118 315 119 316 
<< m1 >>
rect 121 315 122 316 
<< m1 >>
rect 122 315 123 316 
<< m1 >>
rect 123 315 124 316 
<< m1 >>
rect 124 315 125 316 
<< m1 >>
rect 125 315 126 316 
<< m1 >>
rect 126 315 127 316 
<< m1 >>
rect 127 315 128 316 
<< m1 >>
rect 163 315 164 316 
<< m1 >>
rect 181 315 182 316 
<< m1 >>
rect 190 315 191 316 
<< m1 >>
rect 191 315 192 316 
<< m1 >>
rect 192 315 193 316 
<< m1 >>
rect 193 315 194 316 
<< m1 >>
rect 194 315 195 316 
<< m1 >>
rect 195 315 196 316 
<< m1 >>
rect 196 315 197 316 
<< m1 >>
rect 197 315 198 316 
<< m1 >>
rect 198 315 199 316 
<< m1 >>
rect 199 315 200 316 
<< m1 >>
rect 200 315 201 316 
<< m1 >>
rect 201 315 202 316 
<< m1 >>
rect 202 315 203 316 
<< m1 >>
rect 203 315 204 316 
<< m1 >>
rect 204 315 205 316 
<< m1 >>
rect 205 315 206 316 
<< m1 >>
rect 206 315 207 316 
<< m2 >>
rect 206 315 207 316 
<< m2c >>
rect 206 315 207 316 
<< m1 >>
rect 206 315 207 316 
<< m2 >>
rect 206 315 207 316 
<< m1 >>
rect 208 315 209 316 
<< m2 >>
rect 208 315 209 316 
<< m2c >>
rect 208 315 209 316 
<< m1 >>
rect 208 315 209 316 
<< m2 >>
rect 208 315 209 316 
<< m1 >>
rect 213 315 214 316 
<< m2 >>
rect 213 315 214 316 
<< m2c >>
rect 213 315 214 316 
<< m1 >>
rect 213 315 214 316 
<< m2 >>
rect 213 315 214 316 
<< m1 >>
rect 214 315 215 316 
<< m1 >>
rect 215 315 216 316 
<< m1 >>
rect 217 315 218 316 
<< m1 >>
rect 244 315 245 316 
<< m1 >>
rect 247 315 248 316 
<< m1 >>
rect 257 315 258 316 
<< m1 >>
rect 271 315 272 316 
<< m1 >>
rect 280 315 281 316 
<< m1 >>
rect 283 315 284 316 
<< m1 >>
rect 284 315 285 316 
<< m1 >>
rect 285 315 286 316 
<< m1 >>
rect 286 315 287 316 
<< m1 >>
rect 287 315 288 316 
<< m1 >>
rect 288 315 289 316 
<< m1 >>
rect 289 315 290 316 
<< m1 >>
rect 301 315 302 316 
<< m1 >>
rect 307 315 308 316 
<< m2 >>
rect 308 315 309 316 
<< m2 >>
rect 325 315 326 316 
<< m1 >>
rect 352 315 353 316 
<< m1 >>
rect 373 315 374 316 
<< m1 >>
rect 374 315 375 316 
<< m1 >>
rect 375 315 376 316 
<< m1 >>
rect 376 315 377 316 
<< m1 >>
rect 377 315 378 316 
<< m1 >>
rect 378 315 379 316 
<< m1 >>
rect 379 315 380 316 
<< m1 >>
rect 52 316 53 317 
<< m1 >>
rect 53 316 54 317 
<< m1 >>
rect 54 316 55 317 
<< m1 >>
rect 55 316 56 317 
<< m2 >>
rect 55 316 56 317 
<< m1 >>
rect 56 316 57 317 
<< m1 >>
rect 57 316 58 317 
<< m1 >>
rect 58 316 59 317 
<< m1 >>
rect 59 316 60 317 
<< m1 >>
rect 60 316 61 317 
<< m1 >>
rect 61 316 62 317 
<< m1 >>
rect 62 316 63 317 
<< m1 >>
rect 63 316 64 317 
<< m1 >>
rect 64 316 65 317 
<< m1 >>
rect 70 316 71 317 
<< m1 >>
rect 91 316 92 317 
<< m1 >>
rect 118 316 119 317 
<< m1 >>
rect 121 316 122 317 
<< m1 >>
rect 127 316 128 317 
<< m1 >>
rect 163 316 164 317 
<< m1 >>
rect 181 316 182 317 
<< m1 >>
rect 190 316 191 317 
<< m1 >>
rect 208 316 209 317 
<< m1 >>
rect 215 316 216 317 
<< m2 >>
rect 215 316 216 317 
<< m2c >>
rect 215 316 216 317 
<< m1 >>
rect 215 316 216 317 
<< m2 >>
rect 215 316 216 317 
<< m2 >>
rect 216 316 217 317 
<< m1 >>
rect 217 316 218 317 
<< m2 >>
rect 217 316 218 317 
<< m1 >>
rect 244 316 245 317 
<< m1 >>
rect 247 316 248 317 
<< m1 >>
rect 257 316 258 317 
<< m1 >>
rect 271 316 272 317 
<< m1 >>
rect 280 316 281 317 
<< m1 >>
rect 283 316 284 317 
<< m1 >>
rect 289 316 290 317 
<< m1 >>
rect 301 316 302 317 
<< m1 >>
rect 307 316 308 317 
<< m2 >>
rect 308 316 309 317 
<< m1 >>
rect 322 316 323 317 
<< m1 >>
rect 323 316 324 317 
<< m1 >>
rect 324 316 325 317 
<< m1 >>
rect 325 316 326 317 
<< m2 >>
rect 325 316 326 317 
<< m1 >>
rect 352 316 353 317 
<< m1 >>
rect 373 316 374 317 
<< m1 >>
rect 379 316 380 317 
<< m1 >>
rect 52 317 53 318 
<< m2 >>
rect 55 317 56 318 
<< m1 >>
rect 64 317 65 318 
<< m1 >>
rect 70 317 71 318 
<< m1 >>
rect 91 317 92 318 
<< m1 >>
rect 118 317 119 318 
<< m1 >>
rect 121 317 122 318 
<< m1 >>
rect 127 317 128 318 
<< m1 >>
rect 163 317 164 318 
<< m1 >>
rect 181 317 182 318 
<< m1 >>
rect 190 317 191 318 
<< m1 >>
rect 208 317 209 318 
<< m1 >>
rect 217 317 218 318 
<< m2 >>
rect 217 317 218 318 
<< m1 >>
rect 244 317 245 318 
<< m1 >>
rect 247 317 248 318 
<< m1 >>
rect 257 317 258 318 
<< m1 >>
rect 271 317 272 318 
<< m1 >>
rect 280 317 281 318 
<< m1 >>
rect 283 317 284 318 
<< m1 >>
rect 289 317 290 318 
<< m1 >>
rect 301 317 302 318 
<< m1 >>
rect 307 317 308 318 
<< m2 >>
rect 308 317 309 318 
<< m1 >>
rect 322 317 323 318 
<< m1 >>
rect 325 317 326 318 
<< m2 >>
rect 325 317 326 318 
<< m1 >>
rect 352 317 353 318 
<< m1 >>
rect 373 317 374 318 
<< m1 >>
rect 379 317 380 318 
<< pdiffusion >>
rect 12 318 13 319 
<< pdiffusion >>
rect 13 318 14 319 
<< pdiffusion >>
rect 14 318 15 319 
<< pdiffusion >>
rect 15 318 16 319 
<< pdiffusion >>
rect 16 318 17 319 
<< pdiffusion >>
rect 17 318 18 319 
<< pdiffusion >>
rect 30 318 31 319 
<< pdiffusion >>
rect 31 318 32 319 
<< pdiffusion >>
rect 32 318 33 319 
<< pdiffusion >>
rect 33 318 34 319 
<< pdiffusion >>
rect 34 318 35 319 
<< pdiffusion >>
rect 35 318 36 319 
<< pdiffusion >>
rect 48 318 49 319 
<< pdiffusion >>
rect 49 318 50 319 
<< pdiffusion >>
rect 50 318 51 319 
<< pdiffusion >>
rect 51 318 52 319 
<< m1 >>
rect 52 318 53 319 
<< pdiffusion >>
rect 52 318 53 319 
<< pdiffusion >>
rect 53 318 54 319 
<< m1 >>
rect 55 318 56 319 
<< m2 >>
rect 55 318 56 319 
<< m2c >>
rect 55 318 56 319 
<< m1 >>
rect 55 318 56 319 
<< m2 >>
rect 55 318 56 319 
<< m1 >>
rect 64 318 65 319 
<< pdiffusion >>
rect 66 318 67 319 
<< pdiffusion >>
rect 67 318 68 319 
<< pdiffusion >>
rect 68 318 69 319 
<< pdiffusion >>
rect 69 318 70 319 
<< m1 >>
rect 70 318 71 319 
<< pdiffusion >>
rect 70 318 71 319 
<< pdiffusion >>
rect 71 318 72 319 
<< pdiffusion >>
rect 84 318 85 319 
<< pdiffusion >>
rect 85 318 86 319 
<< pdiffusion >>
rect 86 318 87 319 
<< pdiffusion >>
rect 87 318 88 319 
<< pdiffusion >>
rect 88 318 89 319 
<< pdiffusion >>
rect 89 318 90 319 
<< m1 >>
rect 91 318 92 319 
<< m1 >>
rect 118 318 119 319 
<< pdiffusion >>
rect 120 318 121 319 
<< m1 >>
rect 121 318 122 319 
<< pdiffusion >>
rect 121 318 122 319 
<< pdiffusion >>
rect 122 318 123 319 
<< pdiffusion >>
rect 123 318 124 319 
<< pdiffusion >>
rect 124 318 125 319 
<< pdiffusion >>
rect 125 318 126 319 
<< m1 >>
rect 127 318 128 319 
<< pdiffusion >>
rect 138 318 139 319 
<< pdiffusion >>
rect 139 318 140 319 
<< pdiffusion >>
rect 140 318 141 319 
<< pdiffusion >>
rect 141 318 142 319 
<< pdiffusion >>
rect 142 318 143 319 
<< pdiffusion >>
rect 143 318 144 319 
<< pdiffusion >>
rect 156 318 157 319 
<< pdiffusion >>
rect 157 318 158 319 
<< pdiffusion >>
rect 158 318 159 319 
<< pdiffusion >>
rect 159 318 160 319 
<< pdiffusion >>
rect 160 318 161 319 
<< pdiffusion >>
rect 161 318 162 319 
<< m1 >>
rect 163 318 164 319 
<< pdiffusion >>
rect 174 318 175 319 
<< pdiffusion >>
rect 175 318 176 319 
<< pdiffusion >>
rect 176 318 177 319 
<< pdiffusion >>
rect 177 318 178 319 
<< pdiffusion >>
rect 178 318 179 319 
<< pdiffusion >>
rect 179 318 180 319 
<< m1 >>
rect 181 318 182 319 
<< m1 >>
rect 190 318 191 319 
<< m1 >>
rect 208 318 209 319 
<< pdiffusion >>
rect 210 318 211 319 
<< pdiffusion >>
rect 211 318 212 319 
<< pdiffusion >>
rect 212 318 213 319 
<< pdiffusion >>
rect 213 318 214 319 
<< pdiffusion >>
rect 214 318 215 319 
<< pdiffusion >>
rect 215 318 216 319 
<< m1 >>
rect 217 318 218 319 
<< m2 >>
rect 217 318 218 319 
<< pdiffusion >>
rect 228 318 229 319 
<< pdiffusion >>
rect 229 318 230 319 
<< pdiffusion >>
rect 230 318 231 319 
<< pdiffusion >>
rect 231 318 232 319 
<< pdiffusion >>
rect 232 318 233 319 
<< pdiffusion >>
rect 233 318 234 319 
<< m1 >>
rect 244 318 245 319 
<< pdiffusion >>
rect 246 318 247 319 
<< m1 >>
rect 247 318 248 319 
<< pdiffusion >>
rect 247 318 248 319 
<< pdiffusion >>
rect 248 318 249 319 
<< pdiffusion >>
rect 249 318 250 319 
<< pdiffusion >>
rect 250 318 251 319 
<< pdiffusion >>
rect 251 318 252 319 
<< m1 >>
rect 257 318 258 319 
<< pdiffusion >>
rect 264 318 265 319 
<< pdiffusion >>
rect 265 318 266 319 
<< pdiffusion >>
rect 266 318 267 319 
<< pdiffusion >>
rect 267 318 268 319 
<< pdiffusion >>
rect 268 318 269 319 
<< pdiffusion >>
rect 269 318 270 319 
<< m1 >>
rect 271 318 272 319 
<< m1 >>
rect 280 318 281 319 
<< pdiffusion >>
rect 282 318 283 319 
<< m1 >>
rect 283 318 284 319 
<< pdiffusion >>
rect 283 318 284 319 
<< pdiffusion >>
rect 284 318 285 319 
<< pdiffusion >>
rect 285 318 286 319 
<< pdiffusion >>
rect 286 318 287 319 
<< pdiffusion >>
rect 287 318 288 319 
<< m1 >>
rect 289 318 290 319 
<< pdiffusion >>
rect 300 318 301 319 
<< m1 >>
rect 301 318 302 319 
<< pdiffusion >>
rect 301 318 302 319 
<< pdiffusion >>
rect 302 318 303 319 
<< pdiffusion >>
rect 303 318 304 319 
<< pdiffusion >>
rect 304 318 305 319 
<< pdiffusion >>
rect 305 318 306 319 
<< m1 >>
rect 307 318 308 319 
<< m2 >>
rect 308 318 309 319 
<< pdiffusion >>
rect 318 318 319 319 
<< pdiffusion >>
rect 319 318 320 319 
<< pdiffusion >>
rect 320 318 321 319 
<< pdiffusion >>
rect 321 318 322 319 
<< m1 >>
rect 322 318 323 319 
<< pdiffusion >>
rect 322 318 323 319 
<< pdiffusion >>
rect 323 318 324 319 
<< m1 >>
rect 325 318 326 319 
<< m2 >>
rect 325 318 326 319 
<< pdiffusion >>
rect 336 318 337 319 
<< pdiffusion >>
rect 337 318 338 319 
<< pdiffusion >>
rect 338 318 339 319 
<< pdiffusion >>
rect 339 318 340 319 
<< pdiffusion >>
rect 340 318 341 319 
<< pdiffusion >>
rect 341 318 342 319 
<< m1 >>
rect 352 318 353 319 
<< pdiffusion >>
rect 354 318 355 319 
<< pdiffusion >>
rect 355 318 356 319 
<< pdiffusion >>
rect 356 318 357 319 
<< pdiffusion >>
rect 357 318 358 319 
<< pdiffusion >>
rect 358 318 359 319 
<< pdiffusion >>
rect 359 318 360 319 
<< pdiffusion >>
rect 372 318 373 319 
<< m1 >>
rect 373 318 374 319 
<< pdiffusion >>
rect 373 318 374 319 
<< pdiffusion >>
rect 374 318 375 319 
<< pdiffusion >>
rect 375 318 376 319 
<< pdiffusion >>
rect 376 318 377 319 
<< pdiffusion >>
rect 377 318 378 319 
<< m1 >>
rect 379 318 380 319 
<< pdiffusion >>
rect 390 318 391 319 
<< pdiffusion >>
rect 391 318 392 319 
<< pdiffusion >>
rect 392 318 393 319 
<< pdiffusion >>
rect 393 318 394 319 
<< pdiffusion >>
rect 394 318 395 319 
<< pdiffusion >>
rect 395 318 396 319 
<< pdiffusion >>
rect 408 318 409 319 
<< pdiffusion >>
rect 409 318 410 319 
<< pdiffusion >>
rect 410 318 411 319 
<< pdiffusion >>
rect 411 318 412 319 
<< pdiffusion >>
rect 412 318 413 319 
<< pdiffusion >>
rect 413 318 414 319 
<< pdiffusion >>
rect 426 318 427 319 
<< pdiffusion >>
rect 427 318 428 319 
<< pdiffusion >>
rect 428 318 429 319 
<< pdiffusion >>
rect 429 318 430 319 
<< pdiffusion >>
rect 430 318 431 319 
<< pdiffusion >>
rect 431 318 432 319 
<< pdiffusion >>
rect 444 318 445 319 
<< pdiffusion >>
rect 445 318 446 319 
<< pdiffusion >>
rect 446 318 447 319 
<< pdiffusion >>
rect 447 318 448 319 
<< pdiffusion >>
rect 448 318 449 319 
<< pdiffusion >>
rect 449 318 450 319 
<< pdiffusion >>
rect 12 319 13 320 
<< pdiffusion >>
rect 13 319 14 320 
<< pdiffusion >>
rect 14 319 15 320 
<< pdiffusion >>
rect 15 319 16 320 
<< pdiffusion >>
rect 16 319 17 320 
<< pdiffusion >>
rect 17 319 18 320 
<< pdiffusion >>
rect 30 319 31 320 
<< pdiffusion >>
rect 31 319 32 320 
<< pdiffusion >>
rect 32 319 33 320 
<< pdiffusion >>
rect 33 319 34 320 
<< pdiffusion >>
rect 34 319 35 320 
<< pdiffusion >>
rect 35 319 36 320 
<< pdiffusion >>
rect 48 319 49 320 
<< pdiffusion >>
rect 49 319 50 320 
<< pdiffusion >>
rect 50 319 51 320 
<< pdiffusion >>
rect 51 319 52 320 
<< pdiffusion >>
rect 52 319 53 320 
<< pdiffusion >>
rect 53 319 54 320 
<< m1 >>
rect 55 319 56 320 
<< m1 >>
rect 64 319 65 320 
<< pdiffusion >>
rect 66 319 67 320 
<< pdiffusion >>
rect 67 319 68 320 
<< pdiffusion >>
rect 68 319 69 320 
<< pdiffusion >>
rect 69 319 70 320 
<< pdiffusion >>
rect 70 319 71 320 
<< pdiffusion >>
rect 71 319 72 320 
<< pdiffusion >>
rect 84 319 85 320 
<< pdiffusion >>
rect 85 319 86 320 
<< pdiffusion >>
rect 86 319 87 320 
<< pdiffusion >>
rect 87 319 88 320 
<< pdiffusion >>
rect 88 319 89 320 
<< pdiffusion >>
rect 89 319 90 320 
<< m1 >>
rect 91 319 92 320 
<< m1 >>
rect 118 319 119 320 
<< pdiffusion >>
rect 120 319 121 320 
<< pdiffusion >>
rect 121 319 122 320 
<< pdiffusion >>
rect 122 319 123 320 
<< pdiffusion >>
rect 123 319 124 320 
<< pdiffusion >>
rect 124 319 125 320 
<< pdiffusion >>
rect 125 319 126 320 
<< m1 >>
rect 127 319 128 320 
<< pdiffusion >>
rect 138 319 139 320 
<< pdiffusion >>
rect 139 319 140 320 
<< pdiffusion >>
rect 140 319 141 320 
<< pdiffusion >>
rect 141 319 142 320 
<< pdiffusion >>
rect 142 319 143 320 
<< pdiffusion >>
rect 143 319 144 320 
<< pdiffusion >>
rect 156 319 157 320 
<< pdiffusion >>
rect 157 319 158 320 
<< pdiffusion >>
rect 158 319 159 320 
<< pdiffusion >>
rect 159 319 160 320 
<< pdiffusion >>
rect 160 319 161 320 
<< pdiffusion >>
rect 161 319 162 320 
<< m1 >>
rect 163 319 164 320 
<< pdiffusion >>
rect 174 319 175 320 
<< pdiffusion >>
rect 175 319 176 320 
<< pdiffusion >>
rect 176 319 177 320 
<< pdiffusion >>
rect 177 319 178 320 
<< pdiffusion >>
rect 178 319 179 320 
<< pdiffusion >>
rect 179 319 180 320 
<< m1 >>
rect 181 319 182 320 
<< m1 >>
rect 190 319 191 320 
<< m1 >>
rect 208 319 209 320 
<< pdiffusion >>
rect 210 319 211 320 
<< pdiffusion >>
rect 211 319 212 320 
<< pdiffusion >>
rect 212 319 213 320 
<< pdiffusion >>
rect 213 319 214 320 
<< pdiffusion >>
rect 214 319 215 320 
<< pdiffusion >>
rect 215 319 216 320 
<< m1 >>
rect 217 319 218 320 
<< m2 >>
rect 217 319 218 320 
<< pdiffusion >>
rect 228 319 229 320 
<< pdiffusion >>
rect 229 319 230 320 
<< pdiffusion >>
rect 230 319 231 320 
<< pdiffusion >>
rect 231 319 232 320 
<< pdiffusion >>
rect 232 319 233 320 
<< pdiffusion >>
rect 233 319 234 320 
<< m1 >>
rect 244 319 245 320 
<< pdiffusion >>
rect 246 319 247 320 
<< pdiffusion >>
rect 247 319 248 320 
<< pdiffusion >>
rect 248 319 249 320 
<< pdiffusion >>
rect 249 319 250 320 
<< pdiffusion >>
rect 250 319 251 320 
<< pdiffusion >>
rect 251 319 252 320 
<< m1 >>
rect 257 319 258 320 
<< pdiffusion >>
rect 264 319 265 320 
<< pdiffusion >>
rect 265 319 266 320 
<< pdiffusion >>
rect 266 319 267 320 
<< pdiffusion >>
rect 267 319 268 320 
<< pdiffusion >>
rect 268 319 269 320 
<< pdiffusion >>
rect 269 319 270 320 
<< m1 >>
rect 271 319 272 320 
<< m1 >>
rect 280 319 281 320 
<< pdiffusion >>
rect 282 319 283 320 
<< pdiffusion >>
rect 283 319 284 320 
<< pdiffusion >>
rect 284 319 285 320 
<< pdiffusion >>
rect 285 319 286 320 
<< pdiffusion >>
rect 286 319 287 320 
<< pdiffusion >>
rect 287 319 288 320 
<< m1 >>
rect 289 319 290 320 
<< pdiffusion >>
rect 300 319 301 320 
<< pdiffusion >>
rect 301 319 302 320 
<< pdiffusion >>
rect 302 319 303 320 
<< pdiffusion >>
rect 303 319 304 320 
<< pdiffusion >>
rect 304 319 305 320 
<< pdiffusion >>
rect 305 319 306 320 
<< m1 >>
rect 307 319 308 320 
<< m2 >>
rect 308 319 309 320 
<< pdiffusion >>
rect 318 319 319 320 
<< pdiffusion >>
rect 319 319 320 320 
<< pdiffusion >>
rect 320 319 321 320 
<< pdiffusion >>
rect 321 319 322 320 
<< pdiffusion >>
rect 322 319 323 320 
<< pdiffusion >>
rect 323 319 324 320 
<< m1 >>
rect 325 319 326 320 
<< m2 >>
rect 325 319 326 320 
<< pdiffusion >>
rect 336 319 337 320 
<< pdiffusion >>
rect 337 319 338 320 
<< pdiffusion >>
rect 338 319 339 320 
<< pdiffusion >>
rect 339 319 340 320 
<< pdiffusion >>
rect 340 319 341 320 
<< pdiffusion >>
rect 341 319 342 320 
<< m1 >>
rect 352 319 353 320 
<< pdiffusion >>
rect 354 319 355 320 
<< pdiffusion >>
rect 355 319 356 320 
<< pdiffusion >>
rect 356 319 357 320 
<< pdiffusion >>
rect 357 319 358 320 
<< pdiffusion >>
rect 358 319 359 320 
<< pdiffusion >>
rect 359 319 360 320 
<< pdiffusion >>
rect 372 319 373 320 
<< pdiffusion >>
rect 373 319 374 320 
<< pdiffusion >>
rect 374 319 375 320 
<< pdiffusion >>
rect 375 319 376 320 
<< pdiffusion >>
rect 376 319 377 320 
<< pdiffusion >>
rect 377 319 378 320 
<< m1 >>
rect 379 319 380 320 
<< pdiffusion >>
rect 390 319 391 320 
<< pdiffusion >>
rect 391 319 392 320 
<< pdiffusion >>
rect 392 319 393 320 
<< pdiffusion >>
rect 393 319 394 320 
<< pdiffusion >>
rect 394 319 395 320 
<< pdiffusion >>
rect 395 319 396 320 
<< pdiffusion >>
rect 408 319 409 320 
<< pdiffusion >>
rect 409 319 410 320 
<< pdiffusion >>
rect 410 319 411 320 
<< pdiffusion >>
rect 411 319 412 320 
<< pdiffusion >>
rect 412 319 413 320 
<< pdiffusion >>
rect 413 319 414 320 
<< pdiffusion >>
rect 426 319 427 320 
<< pdiffusion >>
rect 427 319 428 320 
<< pdiffusion >>
rect 428 319 429 320 
<< pdiffusion >>
rect 429 319 430 320 
<< pdiffusion >>
rect 430 319 431 320 
<< pdiffusion >>
rect 431 319 432 320 
<< pdiffusion >>
rect 444 319 445 320 
<< pdiffusion >>
rect 445 319 446 320 
<< pdiffusion >>
rect 446 319 447 320 
<< pdiffusion >>
rect 447 319 448 320 
<< pdiffusion >>
rect 448 319 449 320 
<< pdiffusion >>
rect 449 319 450 320 
<< pdiffusion >>
rect 12 320 13 321 
<< pdiffusion >>
rect 13 320 14 321 
<< pdiffusion >>
rect 14 320 15 321 
<< pdiffusion >>
rect 15 320 16 321 
<< pdiffusion >>
rect 16 320 17 321 
<< pdiffusion >>
rect 17 320 18 321 
<< pdiffusion >>
rect 30 320 31 321 
<< pdiffusion >>
rect 31 320 32 321 
<< pdiffusion >>
rect 32 320 33 321 
<< pdiffusion >>
rect 33 320 34 321 
<< pdiffusion >>
rect 34 320 35 321 
<< pdiffusion >>
rect 35 320 36 321 
<< pdiffusion >>
rect 48 320 49 321 
<< pdiffusion >>
rect 49 320 50 321 
<< pdiffusion >>
rect 50 320 51 321 
<< pdiffusion >>
rect 51 320 52 321 
<< pdiffusion >>
rect 52 320 53 321 
<< pdiffusion >>
rect 53 320 54 321 
<< m1 >>
rect 55 320 56 321 
<< m1 >>
rect 64 320 65 321 
<< pdiffusion >>
rect 66 320 67 321 
<< pdiffusion >>
rect 67 320 68 321 
<< pdiffusion >>
rect 68 320 69 321 
<< pdiffusion >>
rect 69 320 70 321 
<< pdiffusion >>
rect 70 320 71 321 
<< pdiffusion >>
rect 71 320 72 321 
<< pdiffusion >>
rect 84 320 85 321 
<< pdiffusion >>
rect 85 320 86 321 
<< pdiffusion >>
rect 86 320 87 321 
<< pdiffusion >>
rect 87 320 88 321 
<< pdiffusion >>
rect 88 320 89 321 
<< pdiffusion >>
rect 89 320 90 321 
<< m1 >>
rect 91 320 92 321 
<< m1 >>
rect 118 320 119 321 
<< pdiffusion >>
rect 120 320 121 321 
<< pdiffusion >>
rect 121 320 122 321 
<< pdiffusion >>
rect 122 320 123 321 
<< pdiffusion >>
rect 123 320 124 321 
<< pdiffusion >>
rect 124 320 125 321 
<< pdiffusion >>
rect 125 320 126 321 
<< m1 >>
rect 127 320 128 321 
<< pdiffusion >>
rect 138 320 139 321 
<< pdiffusion >>
rect 139 320 140 321 
<< pdiffusion >>
rect 140 320 141 321 
<< pdiffusion >>
rect 141 320 142 321 
<< pdiffusion >>
rect 142 320 143 321 
<< pdiffusion >>
rect 143 320 144 321 
<< pdiffusion >>
rect 156 320 157 321 
<< pdiffusion >>
rect 157 320 158 321 
<< pdiffusion >>
rect 158 320 159 321 
<< pdiffusion >>
rect 159 320 160 321 
<< pdiffusion >>
rect 160 320 161 321 
<< pdiffusion >>
rect 161 320 162 321 
<< m1 >>
rect 163 320 164 321 
<< pdiffusion >>
rect 174 320 175 321 
<< pdiffusion >>
rect 175 320 176 321 
<< pdiffusion >>
rect 176 320 177 321 
<< pdiffusion >>
rect 177 320 178 321 
<< pdiffusion >>
rect 178 320 179 321 
<< pdiffusion >>
rect 179 320 180 321 
<< m1 >>
rect 181 320 182 321 
<< m1 >>
rect 190 320 191 321 
<< m1 >>
rect 208 320 209 321 
<< pdiffusion >>
rect 210 320 211 321 
<< pdiffusion >>
rect 211 320 212 321 
<< pdiffusion >>
rect 212 320 213 321 
<< pdiffusion >>
rect 213 320 214 321 
<< pdiffusion >>
rect 214 320 215 321 
<< pdiffusion >>
rect 215 320 216 321 
<< m1 >>
rect 217 320 218 321 
<< m2 >>
rect 217 320 218 321 
<< pdiffusion >>
rect 228 320 229 321 
<< pdiffusion >>
rect 229 320 230 321 
<< pdiffusion >>
rect 230 320 231 321 
<< pdiffusion >>
rect 231 320 232 321 
<< pdiffusion >>
rect 232 320 233 321 
<< pdiffusion >>
rect 233 320 234 321 
<< m1 >>
rect 244 320 245 321 
<< pdiffusion >>
rect 246 320 247 321 
<< pdiffusion >>
rect 247 320 248 321 
<< pdiffusion >>
rect 248 320 249 321 
<< pdiffusion >>
rect 249 320 250 321 
<< pdiffusion >>
rect 250 320 251 321 
<< pdiffusion >>
rect 251 320 252 321 
<< m1 >>
rect 257 320 258 321 
<< pdiffusion >>
rect 264 320 265 321 
<< pdiffusion >>
rect 265 320 266 321 
<< pdiffusion >>
rect 266 320 267 321 
<< pdiffusion >>
rect 267 320 268 321 
<< pdiffusion >>
rect 268 320 269 321 
<< pdiffusion >>
rect 269 320 270 321 
<< m1 >>
rect 271 320 272 321 
<< m1 >>
rect 280 320 281 321 
<< pdiffusion >>
rect 282 320 283 321 
<< pdiffusion >>
rect 283 320 284 321 
<< pdiffusion >>
rect 284 320 285 321 
<< pdiffusion >>
rect 285 320 286 321 
<< pdiffusion >>
rect 286 320 287 321 
<< pdiffusion >>
rect 287 320 288 321 
<< m1 >>
rect 289 320 290 321 
<< pdiffusion >>
rect 300 320 301 321 
<< pdiffusion >>
rect 301 320 302 321 
<< pdiffusion >>
rect 302 320 303 321 
<< pdiffusion >>
rect 303 320 304 321 
<< pdiffusion >>
rect 304 320 305 321 
<< pdiffusion >>
rect 305 320 306 321 
<< m1 >>
rect 307 320 308 321 
<< m2 >>
rect 308 320 309 321 
<< pdiffusion >>
rect 318 320 319 321 
<< pdiffusion >>
rect 319 320 320 321 
<< pdiffusion >>
rect 320 320 321 321 
<< pdiffusion >>
rect 321 320 322 321 
<< pdiffusion >>
rect 322 320 323 321 
<< pdiffusion >>
rect 323 320 324 321 
<< m1 >>
rect 325 320 326 321 
<< m2 >>
rect 325 320 326 321 
<< pdiffusion >>
rect 336 320 337 321 
<< pdiffusion >>
rect 337 320 338 321 
<< pdiffusion >>
rect 338 320 339 321 
<< pdiffusion >>
rect 339 320 340 321 
<< pdiffusion >>
rect 340 320 341 321 
<< pdiffusion >>
rect 341 320 342 321 
<< m1 >>
rect 352 320 353 321 
<< pdiffusion >>
rect 354 320 355 321 
<< pdiffusion >>
rect 355 320 356 321 
<< pdiffusion >>
rect 356 320 357 321 
<< pdiffusion >>
rect 357 320 358 321 
<< pdiffusion >>
rect 358 320 359 321 
<< pdiffusion >>
rect 359 320 360 321 
<< pdiffusion >>
rect 372 320 373 321 
<< pdiffusion >>
rect 373 320 374 321 
<< pdiffusion >>
rect 374 320 375 321 
<< pdiffusion >>
rect 375 320 376 321 
<< pdiffusion >>
rect 376 320 377 321 
<< pdiffusion >>
rect 377 320 378 321 
<< m1 >>
rect 379 320 380 321 
<< pdiffusion >>
rect 390 320 391 321 
<< pdiffusion >>
rect 391 320 392 321 
<< pdiffusion >>
rect 392 320 393 321 
<< pdiffusion >>
rect 393 320 394 321 
<< pdiffusion >>
rect 394 320 395 321 
<< pdiffusion >>
rect 395 320 396 321 
<< pdiffusion >>
rect 408 320 409 321 
<< pdiffusion >>
rect 409 320 410 321 
<< pdiffusion >>
rect 410 320 411 321 
<< pdiffusion >>
rect 411 320 412 321 
<< pdiffusion >>
rect 412 320 413 321 
<< pdiffusion >>
rect 413 320 414 321 
<< pdiffusion >>
rect 426 320 427 321 
<< pdiffusion >>
rect 427 320 428 321 
<< pdiffusion >>
rect 428 320 429 321 
<< pdiffusion >>
rect 429 320 430 321 
<< pdiffusion >>
rect 430 320 431 321 
<< pdiffusion >>
rect 431 320 432 321 
<< pdiffusion >>
rect 444 320 445 321 
<< pdiffusion >>
rect 445 320 446 321 
<< pdiffusion >>
rect 446 320 447 321 
<< pdiffusion >>
rect 447 320 448 321 
<< pdiffusion >>
rect 448 320 449 321 
<< pdiffusion >>
rect 449 320 450 321 
<< pdiffusion >>
rect 12 321 13 322 
<< pdiffusion >>
rect 13 321 14 322 
<< pdiffusion >>
rect 14 321 15 322 
<< pdiffusion >>
rect 15 321 16 322 
<< pdiffusion >>
rect 16 321 17 322 
<< pdiffusion >>
rect 17 321 18 322 
<< pdiffusion >>
rect 30 321 31 322 
<< pdiffusion >>
rect 31 321 32 322 
<< pdiffusion >>
rect 32 321 33 322 
<< pdiffusion >>
rect 33 321 34 322 
<< pdiffusion >>
rect 34 321 35 322 
<< pdiffusion >>
rect 35 321 36 322 
<< pdiffusion >>
rect 48 321 49 322 
<< pdiffusion >>
rect 49 321 50 322 
<< pdiffusion >>
rect 50 321 51 322 
<< pdiffusion >>
rect 51 321 52 322 
<< pdiffusion >>
rect 52 321 53 322 
<< pdiffusion >>
rect 53 321 54 322 
<< m1 >>
rect 55 321 56 322 
<< m1 >>
rect 64 321 65 322 
<< pdiffusion >>
rect 66 321 67 322 
<< pdiffusion >>
rect 67 321 68 322 
<< pdiffusion >>
rect 68 321 69 322 
<< pdiffusion >>
rect 69 321 70 322 
<< pdiffusion >>
rect 70 321 71 322 
<< pdiffusion >>
rect 71 321 72 322 
<< pdiffusion >>
rect 84 321 85 322 
<< pdiffusion >>
rect 85 321 86 322 
<< pdiffusion >>
rect 86 321 87 322 
<< pdiffusion >>
rect 87 321 88 322 
<< pdiffusion >>
rect 88 321 89 322 
<< pdiffusion >>
rect 89 321 90 322 
<< m1 >>
rect 91 321 92 322 
<< m1 >>
rect 118 321 119 322 
<< pdiffusion >>
rect 120 321 121 322 
<< pdiffusion >>
rect 121 321 122 322 
<< pdiffusion >>
rect 122 321 123 322 
<< pdiffusion >>
rect 123 321 124 322 
<< pdiffusion >>
rect 124 321 125 322 
<< pdiffusion >>
rect 125 321 126 322 
<< m1 >>
rect 127 321 128 322 
<< pdiffusion >>
rect 138 321 139 322 
<< pdiffusion >>
rect 139 321 140 322 
<< pdiffusion >>
rect 140 321 141 322 
<< pdiffusion >>
rect 141 321 142 322 
<< pdiffusion >>
rect 142 321 143 322 
<< pdiffusion >>
rect 143 321 144 322 
<< pdiffusion >>
rect 156 321 157 322 
<< pdiffusion >>
rect 157 321 158 322 
<< pdiffusion >>
rect 158 321 159 322 
<< pdiffusion >>
rect 159 321 160 322 
<< pdiffusion >>
rect 160 321 161 322 
<< pdiffusion >>
rect 161 321 162 322 
<< m1 >>
rect 163 321 164 322 
<< pdiffusion >>
rect 174 321 175 322 
<< pdiffusion >>
rect 175 321 176 322 
<< pdiffusion >>
rect 176 321 177 322 
<< pdiffusion >>
rect 177 321 178 322 
<< pdiffusion >>
rect 178 321 179 322 
<< pdiffusion >>
rect 179 321 180 322 
<< m1 >>
rect 181 321 182 322 
<< m1 >>
rect 190 321 191 322 
<< m1 >>
rect 208 321 209 322 
<< pdiffusion >>
rect 210 321 211 322 
<< pdiffusion >>
rect 211 321 212 322 
<< pdiffusion >>
rect 212 321 213 322 
<< pdiffusion >>
rect 213 321 214 322 
<< pdiffusion >>
rect 214 321 215 322 
<< pdiffusion >>
rect 215 321 216 322 
<< m1 >>
rect 217 321 218 322 
<< m2 >>
rect 217 321 218 322 
<< pdiffusion >>
rect 228 321 229 322 
<< pdiffusion >>
rect 229 321 230 322 
<< pdiffusion >>
rect 230 321 231 322 
<< pdiffusion >>
rect 231 321 232 322 
<< pdiffusion >>
rect 232 321 233 322 
<< pdiffusion >>
rect 233 321 234 322 
<< m1 >>
rect 244 321 245 322 
<< pdiffusion >>
rect 246 321 247 322 
<< pdiffusion >>
rect 247 321 248 322 
<< pdiffusion >>
rect 248 321 249 322 
<< pdiffusion >>
rect 249 321 250 322 
<< pdiffusion >>
rect 250 321 251 322 
<< pdiffusion >>
rect 251 321 252 322 
<< m1 >>
rect 257 321 258 322 
<< pdiffusion >>
rect 264 321 265 322 
<< pdiffusion >>
rect 265 321 266 322 
<< pdiffusion >>
rect 266 321 267 322 
<< pdiffusion >>
rect 267 321 268 322 
<< pdiffusion >>
rect 268 321 269 322 
<< pdiffusion >>
rect 269 321 270 322 
<< m1 >>
rect 271 321 272 322 
<< m1 >>
rect 280 321 281 322 
<< pdiffusion >>
rect 282 321 283 322 
<< pdiffusion >>
rect 283 321 284 322 
<< pdiffusion >>
rect 284 321 285 322 
<< pdiffusion >>
rect 285 321 286 322 
<< pdiffusion >>
rect 286 321 287 322 
<< pdiffusion >>
rect 287 321 288 322 
<< m1 >>
rect 289 321 290 322 
<< pdiffusion >>
rect 300 321 301 322 
<< pdiffusion >>
rect 301 321 302 322 
<< pdiffusion >>
rect 302 321 303 322 
<< pdiffusion >>
rect 303 321 304 322 
<< pdiffusion >>
rect 304 321 305 322 
<< pdiffusion >>
rect 305 321 306 322 
<< m1 >>
rect 307 321 308 322 
<< m2 >>
rect 308 321 309 322 
<< pdiffusion >>
rect 318 321 319 322 
<< pdiffusion >>
rect 319 321 320 322 
<< pdiffusion >>
rect 320 321 321 322 
<< pdiffusion >>
rect 321 321 322 322 
<< pdiffusion >>
rect 322 321 323 322 
<< pdiffusion >>
rect 323 321 324 322 
<< m1 >>
rect 325 321 326 322 
<< m2 >>
rect 325 321 326 322 
<< pdiffusion >>
rect 336 321 337 322 
<< pdiffusion >>
rect 337 321 338 322 
<< pdiffusion >>
rect 338 321 339 322 
<< pdiffusion >>
rect 339 321 340 322 
<< pdiffusion >>
rect 340 321 341 322 
<< pdiffusion >>
rect 341 321 342 322 
<< m1 >>
rect 352 321 353 322 
<< pdiffusion >>
rect 354 321 355 322 
<< pdiffusion >>
rect 355 321 356 322 
<< pdiffusion >>
rect 356 321 357 322 
<< pdiffusion >>
rect 357 321 358 322 
<< pdiffusion >>
rect 358 321 359 322 
<< pdiffusion >>
rect 359 321 360 322 
<< pdiffusion >>
rect 372 321 373 322 
<< pdiffusion >>
rect 373 321 374 322 
<< pdiffusion >>
rect 374 321 375 322 
<< pdiffusion >>
rect 375 321 376 322 
<< pdiffusion >>
rect 376 321 377 322 
<< pdiffusion >>
rect 377 321 378 322 
<< m1 >>
rect 379 321 380 322 
<< pdiffusion >>
rect 390 321 391 322 
<< pdiffusion >>
rect 391 321 392 322 
<< pdiffusion >>
rect 392 321 393 322 
<< pdiffusion >>
rect 393 321 394 322 
<< pdiffusion >>
rect 394 321 395 322 
<< pdiffusion >>
rect 395 321 396 322 
<< pdiffusion >>
rect 408 321 409 322 
<< pdiffusion >>
rect 409 321 410 322 
<< pdiffusion >>
rect 410 321 411 322 
<< pdiffusion >>
rect 411 321 412 322 
<< pdiffusion >>
rect 412 321 413 322 
<< pdiffusion >>
rect 413 321 414 322 
<< pdiffusion >>
rect 426 321 427 322 
<< pdiffusion >>
rect 427 321 428 322 
<< pdiffusion >>
rect 428 321 429 322 
<< pdiffusion >>
rect 429 321 430 322 
<< pdiffusion >>
rect 430 321 431 322 
<< pdiffusion >>
rect 431 321 432 322 
<< pdiffusion >>
rect 444 321 445 322 
<< pdiffusion >>
rect 445 321 446 322 
<< pdiffusion >>
rect 446 321 447 322 
<< pdiffusion >>
rect 447 321 448 322 
<< pdiffusion >>
rect 448 321 449 322 
<< pdiffusion >>
rect 449 321 450 322 
<< pdiffusion >>
rect 12 322 13 323 
<< pdiffusion >>
rect 13 322 14 323 
<< pdiffusion >>
rect 14 322 15 323 
<< pdiffusion >>
rect 15 322 16 323 
<< pdiffusion >>
rect 16 322 17 323 
<< pdiffusion >>
rect 17 322 18 323 
<< pdiffusion >>
rect 30 322 31 323 
<< pdiffusion >>
rect 31 322 32 323 
<< pdiffusion >>
rect 32 322 33 323 
<< pdiffusion >>
rect 33 322 34 323 
<< pdiffusion >>
rect 34 322 35 323 
<< pdiffusion >>
rect 35 322 36 323 
<< pdiffusion >>
rect 48 322 49 323 
<< pdiffusion >>
rect 49 322 50 323 
<< pdiffusion >>
rect 50 322 51 323 
<< pdiffusion >>
rect 51 322 52 323 
<< pdiffusion >>
rect 52 322 53 323 
<< pdiffusion >>
rect 53 322 54 323 
<< m1 >>
rect 55 322 56 323 
<< m1 >>
rect 64 322 65 323 
<< pdiffusion >>
rect 66 322 67 323 
<< pdiffusion >>
rect 67 322 68 323 
<< pdiffusion >>
rect 68 322 69 323 
<< pdiffusion >>
rect 69 322 70 323 
<< pdiffusion >>
rect 70 322 71 323 
<< pdiffusion >>
rect 71 322 72 323 
<< pdiffusion >>
rect 84 322 85 323 
<< pdiffusion >>
rect 85 322 86 323 
<< pdiffusion >>
rect 86 322 87 323 
<< pdiffusion >>
rect 87 322 88 323 
<< pdiffusion >>
rect 88 322 89 323 
<< pdiffusion >>
rect 89 322 90 323 
<< m1 >>
rect 91 322 92 323 
<< m1 >>
rect 118 322 119 323 
<< pdiffusion >>
rect 120 322 121 323 
<< pdiffusion >>
rect 121 322 122 323 
<< pdiffusion >>
rect 122 322 123 323 
<< pdiffusion >>
rect 123 322 124 323 
<< pdiffusion >>
rect 124 322 125 323 
<< pdiffusion >>
rect 125 322 126 323 
<< m1 >>
rect 127 322 128 323 
<< pdiffusion >>
rect 138 322 139 323 
<< pdiffusion >>
rect 139 322 140 323 
<< pdiffusion >>
rect 140 322 141 323 
<< pdiffusion >>
rect 141 322 142 323 
<< pdiffusion >>
rect 142 322 143 323 
<< pdiffusion >>
rect 143 322 144 323 
<< pdiffusion >>
rect 156 322 157 323 
<< pdiffusion >>
rect 157 322 158 323 
<< pdiffusion >>
rect 158 322 159 323 
<< pdiffusion >>
rect 159 322 160 323 
<< pdiffusion >>
rect 160 322 161 323 
<< pdiffusion >>
rect 161 322 162 323 
<< m1 >>
rect 163 322 164 323 
<< pdiffusion >>
rect 174 322 175 323 
<< pdiffusion >>
rect 175 322 176 323 
<< pdiffusion >>
rect 176 322 177 323 
<< pdiffusion >>
rect 177 322 178 323 
<< pdiffusion >>
rect 178 322 179 323 
<< pdiffusion >>
rect 179 322 180 323 
<< m1 >>
rect 181 322 182 323 
<< m1 >>
rect 190 322 191 323 
<< m1 >>
rect 208 322 209 323 
<< pdiffusion >>
rect 210 322 211 323 
<< pdiffusion >>
rect 211 322 212 323 
<< pdiffusion >>
rect 212 322 213 323 
<< pdiffusion >>
rect 213 322 214 323 
<< pdiffusion >>
rect 214 322 215 323 
<< pdiffusion >>
rect 215 322 216 323 
<< m1 >>
rect 217 322 218 323 
<< m2 >>
rect 217 322 218 323 
<< pdiffusion >>
rect 228 322 229 323 
<< pdiffusion >>
rect 229 322 230 323 
<< pdiffusion >>
rect 230 322 231 323 
<< pdiffusion >>
rect 231 322 232 323 
<< pdiffusion >>
rect 232 322 233 323 
<< pdiffusion >>
rect 233 322 234 323 
<< m1 >>
rect 244 322 245 323 
<< pdiffusion >>
rect 246 322 247 323 
<< pdiffusion >>
rect 247 322 248 323 
<< pdiffusion >>
rect 248 322 249 323 
<< pdiffusion >>
rect 249 322 250 323 
<< pdiffusion >>
rect 250 322 251 323 
<< pdiffusion >>
rect 251 322 252 323 
<< m1 >>
rect 257 322 258 323 
<< pdiffusion >>
rect 264 322 265 323 
<< pdiffusion >>
rect 265 322 266 323 
<< pdiffusion >>
rect 266 322 267 323 
<< pdiffusion >>
rect 267 322 268 323 
<< pdiffusion >>
rect 268 322 269 323 
<< pdiffusion >>
rect 269 322 270 323 
<< m1 >>
rect 271 322 272 323 
<< m1 >>
rect 280 322 281 323 
<< pdiffusion >>
rect 282 322 283 323 
<< pdiffusion >>
rect 283 322 284 323 
<< pdiffusion >>
rect 284 322 285 323 
<< pdiffusion >>
rect 285 322 286 323 
<< pdiffusion >>
rect 286 322 287 323 
<< pdiffusion >>
rect 287 322 288 323 
<< m1 >>
rect 289 322 290 323 
<< pdiffusion >>
rect 300 322 301 323 
<< pdiffusion >>
rect 301 322 302 323 
<< pdiffusion >>
rect 302 322 303 323 
<< pdiffusion >>
rect 303 322 304 323 
<< pdiffusion >>
rect 304 322 305 323 
<< pdiffusion >>
rect 305 322 306 323 
<< m1 >>
rect 307 322 308 323 
<< m2 >>
rect 308 322 309 323 
<< pdiffusion >>
rect 318 322 319 323 
<< pdiffusion >>
rect 319 322 320 323 
<< pdiffusion >>
rect 320 322 321 323 
<< pdiffusion >>
rect 321 322 322 323 
<< pdiffusion >>
rect 322 322 323 323 
<< pdiffusion >>
rect 323 322 324 323 
<< m1 >>
rect 325 322 326 323 
<< m2 >>
rect 325 322 326 323 
<< pdiffusion >>
rect 336 322 337 323 
<< pdiffusion >>
rect 337 322 338 323 
<< pdiffusion >>
rect 338 322 339 323 
<< pdiffusion >>
rect 339 322 340 323 
<< pdiffusion >>
rect 340 322 341 323 
<< pdiffusion >>
rect 341 322 342 323 
<< m1 >>
rect 352 322 353 323 
<< pdiffusion >>
rect 354 322 355 323 
<< pdiffusion >>
rect 355 322 356 323 
<< pdiffusion >>
rect 356 322 357 323 
<< pdiffusion >>
rect 357 322 358 323 
<< pdiffusion >>
rect 358 322 359 323 
<< pdiffusion >>
rect 359 322 360 323 
<< pdiffusion >>
rect 372 322 373 323 
<< pdiffusion >>
rect 373 322 374 323 
<< pdiffusion >>
rect 374 322 375 323 
<< pdiffusion >>
rect 375 322 376 323 
<< pdiffusion >>
rect 376 322 377 323 
<< pdiffusion >>
rect 377 322 378 323 
<< m1 >>
rect 379 322 380 323 
<< pdiffusion >>
rect 390 322 391 323 
<< pdiffusion >>
rect 391 322 392 323 
<< pdiffusion >>
rect 392 322 393 323 
<< pdiffusion >>
rect 393 322 394 323 
<< pdiffusion >>
rect 394 322 395 323 
<< pdiffusion >>
rect 395 322 396 323 
<< pdiffusion >>
rect 408 322 409 323 
<< pdiffusion >>
rect 409 322 410 323 
<< pdiffusion >>
rect 410 322 411 323 
<< pdiffusion >>
rect 411 322 412 323 
<< pdiffusion >>
rect 412 322 413 323 
<< pdiffusion >>
rect 413 322 414 323 
<< pdiffusion >>
rect 426 322 427 323 
<< pdiffusion >>
rect 427 322 428 323 
<< pdiffusion >>
rect 428 322 429 323 
<< pdiffusion >>
rect 429 322 430 323 
<< pdiffusion >>
rect 430 322 431 323 
<< pdiffusion >>
rect 431 322 432 323 
<< pdiffusion >>
rect 444 322 445 323 
<< pdiffusion >>
rect 445 322 446 323 
<< pdiffusion >>
rect 446 322 447 323 
<< pdiffusion >>
rect 447 322 448 323 
<< pdiffusion >>
rect 448 322 449 323 
<< pdiffusion >>
rect 449 322 450 323 
<< pdiffusion >>
rect 12 323 13 324 
<< pdiffusion >>
rect 13 323 14 324 
<< pdiffusion >>
rect 14 323 15 324 
<< pdiffusion >>
rect 15 323 16 324 
<< pdiffusion >>
rect 16 323 17 324 
<< pdiffusion >>
rect 17 323 18 324 
<< pdiffusion >>
rect 30 323 31 324 
<< pdiffusion >>
rect 31 323 32 324 
<< pdiffusion >>
rect 32 323 33 324 
<< pdiffusion >>
rect 33 323 34 324 
<< pdiffusion >>
rect 34 323 35 324 
<< pdiffusion >>
rect 35 323 36 324 
<< pdiffusion >>
rect 48 323 49 324 
<< m1 >>
rect 49 323 50 324 
<< pdiffusion >>
rect 49 323 50 324 
<< pdiffusion >>
rect 50 323 51 324 
<< pdiffusion >>
rect 51 323 52 324 
<< pdiffusion >>
rect 52 323 53 324 
<< pdiffusion >>
rect 53 323 54 324 
<< m1 >>
rect 55 323 56 324 
<< m1 >>
rect 64 323 65 324 
<< pdiffusion >>
rect 66 323 67 324 
<< m1 >>
rect 67 323 68 324 
<< pdiffusion >>
rect 67 323 68 324 
<< pdiffusion >>
rect 68 323 69 324 
<< pdiffusion >>
rect 69 323 70 324 
<< pdiffusion >>
rect 70 323 71 324 
<< pdiffusion >>
rect 71 323 72 324 
<< pdiffusion >>
rect 84 323 85 324 
<< pdiffusion >>
rect 85 323 86 324 
<< pdiffusion >>
rect 86 323 87 324 
<< pdiffusion >>
rect 87 323 88 324 
<< m1 >>
rect 88 323 89 324 
<< pdiffusion >>
rect 88 323 89 324 
<< pdiffusion >>
rect 89 323 90 324 
<< m1 >>
rect 91 323 92 324 
<< m1 >>
rect 118 323 119 324 
<< pdiffusion >>
rect 120 323 121 324 
<< pdiffusion >>
rect 121 323 122 324 
<< pdiffusion >>
rect 122 323 123 324 
<< pdiffusion >>
rect 123 323 124 324 
<< m1 >>
rect 124 323 125 324 
<< pdiffusion >>
rect 124 323 125 324 
<< pdiffusion >>
rect 125 323 126 324 
<< m1 >>
rect 127 323 128 324 
<< pdiffusion >>
rect 138 323 139 324 
<< pdiffusion >>
rect 139 323 140 324 
<< pdiffusion >>
rect 140 323 141 324 
<< pdiffusion >>
rect 141 323 142 324 
<< pdiffusion >>
rect 142 323 143 324 
<< pdiffusion >>
rect 143 323 144 324 
<< pdiffusion >>
rect 156 323 157 324 
<< m1 >>
rect 157 323 158 324 
<< pdiffusion >>
rect 157 323 158 324 
<< pdiffusion >>
rect 158 323 159 324 
<< pdiffusion >>
rect 159 323 160 324 
<< pdiffusion >>
rect 160 323 161 324 
<< pdiffusion >>
rect 161 323 162 324 
<< m1 >>
rect 163 323 164 324 
<< pdiffusion >>
rect 174 323 175 324 
<< m1 >>
rect 175 323 176 324 
<< pdiffusion >>
rect 175 323 176 324 
<< pdiffusion >>
rect 176 323 177 324 
<< m1 >>
rect 177 323 178 324 
<< m2 >>
rect 177 323 178 324 
<< m2c >>
rect 177 323 178 324 
<< m1 >>
rect 177 323 178 324 
<< m2 >>
rect 177 323 178 324 
<< pdiffusion >>
rect 177 323 178 324 
<< m1 >>
rect 178 323 179 324 
<< pdiffusion >>
rect 178 323 179 324 
<< pdiffusion >>
rect 179 323 180 324 
<< m1 >>
rect 181 323 182 324 
<< m1 >>
rect 190 323 191 324 
<< m1 >>
rect 208 323 209 324 
<< pdiffusion >>
rect 210 323 211 324 
<< pdiffusion >>
rect 211 323 212 324 
<< pdiffusion >>
rect 212 323 213 324 
<< pdiffusion >>
rect 213 323 214 324 
<< m1 >>
rect 214 323 215 324 
<< pdiffusion >>
rect 214 323 215 324 
<< pdiffusion >>
rect 215 323 216 324 
<< m1 >>
rect 217 323 218 324 
<< m2 >>
rect 217 323 218 324 
<< pdiffusion >>
rect 228 323 229 324 
<< pdiffusion >>
rect 229 323 230 324 
<< pdiffusion >>
rect 230 323 231 324 
<< pdiffusion >>
rect 231 323 232 324 
<< pdiffusion >>
rect 232 323 233 324 
<< pdiffusion >>
rect 233 323 234 324 
<< m1 >>
rect 244 323 245 324 
<< pdiffusion >>
rect 246 323 247 324 
<< pdiffusion >>
rect 247 323 248 324 
<< pdiffusion >>
rect 248 323 249 324 
<< pdiffusion >>
rect 249 323 250 324 
<< m1 >>
rect 250 323 251 324 
<< pdiffusion >>
rect 250 323 251 324 
<< pdiffusion >>
rect 251 323 252 324 
<< m1 >>
rect 257 323 258 324 
<< pdiffusion >>
rect 264 323 265 324 
<< pdiffusion >>
rect 265 323 266 324 
<< pdiffusion >>
rect 266 323 267 324 
<< pdiffusion >>
rect 267 323 268 324 
<< pdiffusion >>
rect 268 323 269 324 
<< pdiffusion >>
rect 269 323 270 324 
<< m1 >>
rect 271 323 272 324 
<< m1 >>
rect 280 323 281 324 
<< pdiffusion >>
rect 282 323 283 324 
<< m1 >>
rect 283 323 284 324 
<< pdiffusion >>
rect 283 323 284 324 
<< pdiffusion >>
rect 284 323 285 324 
<< pdiffusion >>
rect 285 323 286 324 
<< m1 >>
rect 286 323 287 324 
<< pdiffusion >>
rect 286 323 287 324 
<< pdiffusion >>
rect 287 323 288 324 
<< m1 >>
rect 289 323 290 324 
<< pdiffusion >>
rect 300 323 301 324 
<< m1 >>
rect 301 323 302 324 
<< pdiffusion >>
rect 301 323 302 324 
<< pdiffusion >>
rect 302 323 303 324 
<< pdiffusion >>
rect 303 323 304 324 
<< pdiffusion >>
rect 304 323 305 324 
<< pdiffusion >>
rect 305 323 306 324 
<< m1 >>
rect 307 323 308 324 
<< m2 >>
rect 308 323 309 324 
<< pdiffusion >>
rect 318 323 319 324 
<< pdiffusion >>
rect 319 323 320 324 
<< pdiffusion >>
rect 320 323 321 324 
<< m1 >>
rect 321 323 322 324 
<< m2 >>
rect 321 323 322 324 
<< m2c >>
rect 321 323 322 324 
<< m1 >>
rect 321 323 322 324 
<< m2 >>
rect 321 323 322 324 
<< pdiffusion >>
rect 321 323 322 324 
<< m1 >>
rect 322 323 323 324 
<< pdiffusion >>
rect 322 323 323 324 
<< pdiffusion >>
rect 323 323 324 324 
<< m1 >>
rect 325 323 326 324 
<< m2 >>
rect 325 323 326 324 
<< pdiffusion >>
rect 336 323 337 324 
<< pdiffusion >>
rect 337 323 338 324 
<< pdiffusion >>
rect 338 323 339 324 
<< pdiffusion >>
rect 339 323 340 324 
<< pdiffusion >>
rect 340 323 341 324 
<< pdiffusion >>
rect 341 323 342 324 
<< m1 >>
rect 352 323 353 324 
<< pdiffusion >>
rect 354 323 355 324 
<< pdiffusion >>
rect 355 323 356 324 
<< pdiffusion >>
rect 356 323 357 324 
<< pdiffusion >>
rect 357 323 358 324 
<< pdiffusion >>
rect 358 323 359 324 
<< pdiffusion >>
rect 359 323 360 324 
<< pdiffusion >>
rect 372 323 373 324 
<< pdiffusion >>
rect 373 323 374 324 
<< pdiffusion >>
rect 374 323 375 324 
<< pdiffusion >>
rect 375 323 376 324 
<< pdiffusion >>
rect 376 323 377 324 
<< pdiffusion >>
rect 377 323 378 324 
<< m1 >>
rect 379 323 380 324 
<< pdiffusion >>
rect 390 323 391 324 
<< pdiffusion >>
rect 391 323 392 324 
<< pdiffusion >>
rect 392 323 393 324 
<< pdiffusion >>
rect 393 323 394 324 
<< pdiffusion >>
rect 394 323 395 324 
<< pdiffusion >>
rect 395 323 396 324 
<< pdiffusion >>
rect 408 323 409 324 
<< pdiffusion >>
rect 409 323 410 324 
<< pdiffusion >>
rect 410 323 411 324 
<< pdiffusion >>
rect 411 323 412 324 
<< pdiffusion >>
rect 412 323 413 324 
<< pdiffusion >>
rect 413 323 414 324 
<< pdiffusion >>
rect 426 323 427 324 
<< pdiffusion >>
rect 427 323 428 324 
<< pdiffusion >>
rect 428 323 429 324 
<< pdiffusion >>
rect 429 323 430 324 
<< pdiffusion >>
rect 430 323 431 324 
<< pdiffusion >>
rect 431 323 432 324 
<< pdiffusion >>
rect 444 323 445 324 
<< pdiffusion >>
rect 445 323 446 324 
<< pdiffusion >>
rect 446 323 447 324 
<< pdiffusion >>
rect 447 323 448 324 
<< pdiffusion >>
rect 448 323 449 324 
<< pdiffusion >>
rect 449 323 450 324 
<< m1 >>
rect 49 324 50 325 
<< m1 >>
rect 55 324 56 325 
<< m1 >>
rect 64 324 65 325 
<< m1 >>
rect 67 324 68 325 
<< m1 >>
rect 88 324 89 325 
<< m1 >>
rect 91 324 92 325 
<< m1 >>
rect 118 324 119 325 
<< m1 >>
rect 124 324 125 325 
<< m1 >>
rect 127 324 128 325 
<< m1 >>
rect 157 324 158 325 
<< m1 >>
rect 163 324 164 325 
<< m1 >>
rect 175 324 176 325 
<< m1 >>
rect 178 324 179 325 
<< m2 >>
rect 178 324 179 325 
<< m1 >>
rect 181 324 182 325 
<< m1 >>
rect 190 324 191 325 
<< m1 >>
rect 208 324 209 325 
<< m1 >>
rect 214 324 215 325 
<< m1 >>
rect 217 324 218 325 
<< m2 >>
rect 217 324 218 325 
<< m1 >>
rect 244 324 245 325 
<< m1 >>
rect 250 324 251 325 
<< m1 >>
rect 257 324 258 325 
<< m1 >>
rect 271 324 272 325 
<< m1 >>
rect 280 324 281 325 
<< m1 >>
rect 283 324 284 325 
<< m1 >>
rect 286 324 287 325 
<< m1 >>
rect 289 324 290 325 
<< m1 >>
rect 301 324 302 325 
<< m1 >>
rect 307 324 308 325 
<< m2 >>
rect 308 324 309 325 
<< m1 >>
rect 322 324 323 325 
<< m2 >>
rect 322 324 323 325 
<< m1 >>
rect 325 324 326 325 
<< m2 >>
rect 325 324 326 325 
<< m1 >>
rect 352 324 353 325 
<< m1 >>
rect 379 324 380 325 
<< m1 >>
rect 49 325 50 326 
<< m1 >>
rect 55 325 56 326 
<< m1 >>
rect 64 325 65 326 
<< m1 >>
rect 65 325 66 326 
<< m1 >>
rect 66 325 67 326 
<< m1 >>
rect 67 325 68 326 
<< m1 >>
rect 88 325 89 326 
<< m1 >>
rect 91 325 92 326 
<< m1 >>
rect 118 325 119 326 
<< m1 >>
rect 124 325 125 326 
<< m1 >>
rect 125 325 126 326 
<< m2 >>
rect 125 325 126 326 
<< m2c >>
rect 125 325 126 326 
<< m1 >>
rect 125 325 126 326 
<< m2 >>
rect 125 325 126 326 
<< m2 >>
rect 126 325 127 326 
<< m1 >>
rect 127 325 128 326 
<< m2 >>
rect 127 325 128 326 
<< m2 >>
rect 128 325 129 326 
<< m1 >>
rect 129 325 130 326 
<< m2 >>
rect 129 325 130 326 
<< m2c >>
rect 129 325 130 326 
<< m1 >>
rect 129 325 130 326 
<< m2 >>
rect 129 325 130 326 
<< m1 >>
rect 157 325 158 326 
<< m1 >>
rect 163 325 164 326 
<< m1 >>
rect 175 325 176 326 
<< m2 >>
rect 178 325 179 326 
<< m1 >>
rect 181 325 182 326 
<< m1 >>
rect 190 325 191 326 
<< m1 >>
rect 208 325 209 326 
<< m1 >>
rect 214 325 215 326 
<< m1 >>
rect 215 325 216 326 
<< m2 >>
rect 215 325 216 326 
<< m2c >>
rect 215 325 216 326 
<< m1 >>
rect 215 325 216 326 
<< m2 >>
rect 215 325 216 326 
<< m2 >>
rect 216 325 217 326 
<< m1 >>
rect 217 325 218 326 
<< m2 >>
rect 217 325 218 326 
<< m1 >>
rect 244 325 245 326 
<< m1 >>
rect 250 325 251 326 
<< m1 >>
rect 251 325 252 326 
<< m1 >>
rect 252 325 253 326 
<< m1 >>
rect 253 325 254 326 
<< m1 >>
rect 257 325 258 326 
<< m1 >>
rect 271 325 272 326 
<< m1 >>
rect 280 325 281 326 
<< m1 >>
rect 281 325 282 326 
<< m1 >>
rect 282 325 283 326 
<< m1 >>
rect 283 325 284 326 
<< m1 >>
rect 286 325 287 326 
<< m1 >>
rect 289 325 290 326 
<< m1 >>
rect 301 325 302 326 
<< m1 >>
rect 305 325 306 326 
<< m2 >>
rect 305 325 306 326 
<< m2c >>
rect 305 325 306 326 
<< m1 >>
rect 305 325 306 326 
<< m2 >>
rect 305 325 306 326 
<< m2 >>
rect 306 325 307 326 
<< m1 >>
rect 307 325 308 326 
<< m2 >>
rect 307 325 308 326 
<< m2 >>
rect 308 325 309 326 
<< m2 >>
rect 322 325 323 326 
<< m2 >>
rect 323 325 324 326 
<< m2 >>
rect 324 325 325 326 
<< m1 >>
rect 325 325 326 326 
<< m2 >>
rect 325 325 326 326 
<< m1 >>
rect 352 325 353 326 
<< m1 >>
rect 379 325 380 326 
<< m1 >>
rect 49 326 50 327 
<< m1 >>
rect 50 326 51 327 
<< m1 >>
rect 51 326 52 327 
<< m1 >>
rect 52 326 53 327 
<< m1 >>
rect 53 326 54 327 
<< m1 >>
rect 54 326 55 327 
<< m1 >>
rect 55 326 56 327 
<< m1 >>
rect 88 326 89 327 
<< m1 >>
rect 91 326 92 327 
<< m1 >>
rect 118 326 119 327 
<< m1 >>
rect 127 326 128 327 
<< m1 >>
rect 129 326 130 327 
<< m1 >>
rect 157 326 158 327 
<< m1 >>
rect 163 326 164 327 
<< m1 >>
rect 175 326 176 327 
<< m1 >>
rect 176 326 177 327 
<< m1 >>
rect 177 326 178 327 
<< m1 >>
rect 178 326 179 327 
<< m2 >>
rect 178 326 179 327 
<< m1 >>
rect 179 326 180 327 
<< m1 >>
rect 180 326 181 327 
<< m1 >>
rect 181 326 182 327 
<< m1 >>
rect 190 326 191 327 
<< m1 >>
rect 208 326 209 327 
<< m1 >>
rect 217 326 218 327 
<< m1 >>
rect 244 326 245 327 
<< m1 >>
rect 253 326 254 327 
<< m1 >>
rect 257 326 258 327 
<< m1 >>
rect 271 326 272 327 
<< m1 >>
rect 286 326 287 327 
<< m1 >>
rect 289 326 290 327 
<< m1 >>
rect 301 326 302 327 
<< m1 >>
rect 302 326 303 327 
<< m1 >>
rect 303 326 304 327 
<< m1 >>
rect 304 326 305 327 
<< m1 >>
rect 305 326 306 327 
<< m1 >>
rect 307 326 308 327 
<< m1 >>
rect 322 326 323 327 
<< m1 >>
rect 323 326 324 327 
<< m1 >>
rect 324 326 325 327 
<< m1 >>
rect 325 326 326 327 
<< m1 >>
rect 352 326 353 327 
<< m1 >>
rect 353 326 354 327 
<< m1 >>
rect 354 326 355 327 
<< m2 >>
rect 354 326 355 327 
<< m2c >>
rect 354 326 355 327 
<< m1 >>
rect 354 326 355 327 
<< m2 >>
rect 354 326 355 327 
<< m1 >>
rect 379 326 380 327 
<< m1 >>
rect 88 327 89 328 
<< m1 >>
rect 91 327 92 328 
<< m1 >>
rect 118 327 119 328 
<< m1 >>
rect 127 327 128 328 
<< m1 >>
rect 129 327 130 328 
<< m1 >>
rect 157 327 158 328 
<< m1 >>
rect 163 327 164 328 
<< m2 >>
rect 178 327 179 328 
<< m1 >>
rect 190 327 191 328 
<< m1 >>
rect 208 327 209 328 
<< m1 >>
rect 217 327 218 328 
<< m1 >>
rect 244 327 245 328 
<< m1 >>
rect 253 327 254 328 
<< m1 >>
rect 257 327 258 328 
<< m1 >>
rect 271 327 272 328 
<< m1 >>
rect 286 327 287 328 
<< m1 >>
rect 289 327 290 328 
<< m1 >>
rect 307 327 308 328 
<< m1 >>
rect 322 327 323 328 
<< m2 >>
rect 354 327 355 328 
<< m1 >>
rect 379 327 380 328 
<< m1 >>
rect 88 328 89 329 
<< m1 >>
rect 91 328 92 329 
<< m1 >>
rect 118 328 119 329 
<< m1 >>
rect 127 328 128 329 
<< m1 >>
rect 129 328 130 329 
<< m1 >>
rect 130 328 131 329 
<< m1 >>
rect 131 328 132 329 
<< m1 >>
rect 132 328 133 329 
<< m1 >>
rect 133 328 134 329 
<< m1 >>
rect 134 328 135 329 
<< m1 >>
rect 135 328 136 329 
<< m1 >>
rect 136 328 137 329 
<< m1 >>
rect 137 328 138 329 
<< m1 >>
rect 138 328 139 329 
<< m1 >>
rect 139 328 140 329 
<< m1 >>
rect 140 328 141 329 
<< m1 >>
rect 141 328 142 329 
<< m1 >>
rect 142 328 143 329 
<< m1 >>
rect 143 328 144 329 
<< m1 >>
rect 144 328 145 329 
<< m1 >>
rect 145 328 146 329 
<< m1 >>
rect 146 328 147 329 
<< m1 >>
rect 147 328 148 329 
<< m1 >>
rect 148 328 149 329 
<< m1 >>
rect 149 328 150 329 
<< m1 >>
rect 150 328 151 329 
<< m1 >>
rect 151 328 152 329 
<< m1 >>
rect 152 328 153 329 
<< m1 >>
rect 153 328 154 329 
<< m1 >>
rect 154 328 155 329 
<< m1 >>
rect 155 328 156 329 
<< m1 >>
rect 156 328 157 329 
<< m1 >>
rect 157 328 158 329 
<< m1 >>
rect 163 328 164 329 
<< m1 >>
rect 172 328 173 329 
<< m1 >>
rect 173 328 174 329 
<< m1 >>
rect 174 328 175 329 
<< m1 >>
rect 175 328 176 329 
<< m1 >>
rect 176 328 177 329 
<< m1 >>
rect 177 328 178 329 
<< m1 >>
rect 178 328 179 329 
<< m2 >>
rect 178 328 179 329 
<< m2c >>
rect 178 328 179 329 
<< m1 >>
rect 178 328 179 329 
<< m2 >>
rect 178 328 179 329 
<< m1 >>
rect 190 328 191 329 
<< m1 >>
rect 208 328 209 329 
<< m1 >>
rect 217 328 218 329 
<< m1 >>
rect 244 328 245 329 
<< m1 >>
rect 253 328 254 329 
<< m1 >>
rect 257 328 258 329 
<< m1 >>
rect 271 328 272 329 
<< m1 >>
rect 272 328 273 329 
<< m1 >>
rect 273 328 274 329 
<< m1 >>
rect 274 328 275 329 
<< m1 >>
rect 275 328 276 329 
<< m1 >>
rect 276 328 277 329 
<< m1 >>
rect 277 328 278 329 
<< m1 >>
rect 278 328 279 329 
<< m1 >>
rect 279 328 280 329 
<< m1 >>
rect 280 328 281 329 
<< m1 >>
rect 281 328 282 329 
<< m1 >>
rect 282 328 283 329 
<< m1 >>
rect 283 328 284 329 
<< m1 >>
rect 284 328 285 329 
<< m1 >>
rect 285 328 286 329 
<< m1 >>
rect 286 328 287 329 
<< m1 >>
rect 289 328 290 329 
<< m1 >>
rect 307 328 308 329 
<< m1 >>
rect 308 328 309 329 
<< m1 >>
rect 309 328 310 329 
<< m1 >>
rect 310 328 311 329 
<< m1 >>
rect 311 328 312 329 
<< m1 >>
rect 312 328 313 329 
<< m1 >>
rect 313 328 314 329 
<< m1 >>
rect 314 328 315 329 
<< m1 >>
rect 315 328 316 329 
<< m1 >>
rect 316 328 317 329 
<< m1 >>
rect 317 328 318 329 
<< m1 >>
rect 318 328 319 329 
<< m1 >>
rect 319 328 320 329 
<< m1 >>
rect 320 328 321 329 
<< m2 >>
rect 320 328 321 329 
<< m2c >>
rect 320 328 321 329 
<< m1 >>
rect 320 328 321 329 
<< m2 >>
rect 320 328 321 329 
<< m2 >>
rect 321 328 322 329 
<< m1 >>
rect 322 328 323 329 
<< m2 >>
rect 322 328 323 329 
<< m2 >>
rect 323 328 324 329 
<< m1 >>
rect 324 328 325 329 
<< m2 >>
rect 324 328 325 329 
<< m2c >>
rect 324 328 325 329 
<< m1 >>
rect 324 328 325 329 
<< m2 >>
rect 324 328 325 329 
<< m1 >>
rect 325 328 326 329 
<< m1 >>
rect 326 328 327 329 
<< m1 >>
rect 327 328 328 329 
<< m1 >>
rect 328 328 329 329 
<< m1 >>
rect 329 328 330 329 
<< m1 >>
rect 330 328 331 329 
<< m1 >>
rect 331 328 332 329 
<< m1 >>
rect 332 328 333 329 
<< m1 >>
rect 333 328 334 329 
<< m1 >>
rect 334 328 335 329 
<< m1 >>
rect 335 328 336 329 
<< m1 >>
rect 336 328 337 329 
<< m1 >>
rect 337 328 338 329 
<< m1 >>
rect 338 328 339 329 
<< m1 >>
rect 339 328 340 329 
<< m1 >>
rect 340 328 341 329 
<< m1 >>
rect 341 328 342 329 
<< m1 >>
rect 342 328 343 329 
<< m1 >>
rect 343 328 344 329 
<< m1 >>
rect 344 328 345 329 
<< m1 >>
rect 345 328 346 329 
<< m1 >>
rect 346 328 347 329 
<< m1 >>
rect 347 328 348 329 
<< m1 >>
rect 348 328 349 329 
<< m1 >>
rect 349 328 350 329 
<< m1 >>
rect 350 328 351 329 
<< m1 >>
rect 351 328 352 329 
<< m1 >>
rect 352 328 353 329 
<< m1 >>
rect 353 328 354 329 
<< m1 >>
rect 354 328 355 329 
<< m2 >>
rect 354 328 355 329 
<< m1 >>
rect 355 328 356 329 
<< m1 >>
rect 356 328 357 329 
<< m1 >>
rect 357 328 358 329 
<< m1 >>
rect 358 328 359 329 
<< m1 >>
rect 359 328 360 329 
<< m1 >>
rect 360 328 361 329 
<< m1 >>
rect 361 328 362 329 
<< m1 >>
rect 362 328 363 329 
<< m1 >>
rect 363 328 364 329 
<< m1 >>
rect 364 328 365 329 
<< m1 >>
rect 365 328 366 329 
<< m1 >>
rect 366 328 367 329 
<< m1 >>
rect 367 328 368 329 
<< m1 >>
rect 368 328 369 329 
<< m1 >>
rect 369 328 370 329 
<< m1 >>
rect 370 328 371 329 
<< m1 >>
rect 371 328 372 329 
<< m1 >>
rect 372 328 373 329 
<< m1 >>
rect 373 328 374 329 
<< m1 >>
rect 374 328 375 329 
<< m1 >>
rect 375 328 376 329 
<< m1 >>
rect 376 328 377 329 
<< m1 >>
rect 379 328 380 329 
<< m1 >>
rect 380 328 381 329 
<< m1 >>
rect 381 328 382 329 
<< m1 >>
rect 382 328 383 329 
<< m1 >>
rect 383 328 384 329 
<< m1 >>
rect 384 328 385 329 
<< m1 >>
rect 385 328 386 329 
<< m1 >>
rect 386 328 387 329 
<< m1 >>
rect 387 328 388 329 
<< m1 >>
rect 388 328 389 329 
<< m1 >>
rect 389 328 390 329 
<< m1 >>
rect 390 328 391 329 
<< m1 >>
rect 391 328 392 329 
<< m1 >>
rect 88 329 89 330 
<< m1 >>
rect 91 329 92 330 
<< m1 >>
rect 118 329 119 330 
<< m1 >>
rect 127 329 128 330 
<< m1 >>
rect 163 329 164 330 
<< m1 >>
rect 172 329 173 330 
<< m1 >>
rect 190 329 191 330 
<< m1 >>
rect 208 329 209 330 
<< m1 >>
rect 217 329 218 330 
<< m1 >>
rect 244 329 245 330 
<< m1 >>
rect 253 329 254 330 
<< m1 >>
rect 257 329 258 330 
<< m1 >>
rect 289 329 290 330 
<< m1 >>
rect 322 329 323 330 
<< m2 >>
rect 354 329 355 330 
<< m2 >>
rect 355 329 356 330 
<< m1 >>
rect 376 329 377 330 
<< m1 >>
rect 391 329 392 330 
<< m1 >>
rect 88 330 89 331 
<< m1 >>
rect 91 330 92 331 
<< m1 >>
rect 118 330 119 331 
<< m1 >>
rect 127 330 128 331 
<< m1 >>
rect 163 330 164 331 
<< m1 >>
rect 172 330 173 331 
<< m1 >>
rect 190 330 191 331 
<< m1 >>
rect 208 330 209 331 
<< m1 >>
rect 217 330 218 331 
<< m1 >>
rect 244 330 245 331 
<< m1 >>
rect 253 330 254 331 
<< m1 >>
rect 257 330 258 331 
<< m1 >>
rect 289 330 290 331 
<< m1 >>
rect 322 330 323 331 
<< m1 >>
rect 355 330 356 331 
<< m2 >>
rect 355 330 356 331 
<< m2c >>
rect 355 330 356 331 
<< m1 >>
rect 355 330 356 331 
<< m2 >>
rect 355 330 356 331 
<< m1 >>
rect 376 330 377 331 
<< m1 >>
rect 391 330 392 331 
<< m1 >>
rect 73 331 74 332 
<< m1 >>
rect 74 331 75 332 
<< m1 >>
rect 75 331 76 332 
<< m1 >>
rect 76 331 77 332 
<< m1 >>
rect 77 331 78 332 
<< m1 >>
rect 78 331 79 332 
<< m1 >>
rect 79 331 80 332 
<< m1 >>
rect 80 331 81 332 
<< m1 >>
rect 81 331 82 332 
<< m1 >>
rect 82 331 83 332 
<< m1 >>
rect 83 331 84 332 
<< m1 >>
rect 84 331 85 332 
<< m1 >>
rect 85 331 86 332 
<< m1 >>
rect 86 331 87 332 
<< m1 >>
rect 87 331 88 332 
<< m1 >>
rect 88 331 89 332 
<< m1 >>
rect 91 331 92 332 
<< m1 >>
rect 118 331 119 332 
<< m1 >>
rect 127 331 128 332 
<< m1 >>
rect 145 331 146 332 
<< m1 >>
rect 146 331 147 332 
<< m1 >>
rect 147 331 148 332 
<< m1 >>
rect 148 331 149 332 
<< m1 >>
rect 149 331 150 332 
<< m1 >>
rect 150 331 151 332 
<< m1 >>
rect 151 331 152 332 
<< m1 >>
rect 152 331 153 332 
<< m1 >>
rect 153 331 154 332 
<< m1 >>
rect 154 331 155 332 
<< m1 >>
rect 155 331 156 332 
<< m1 >>
rect 156 331 157 332 
<< m1 >>
rect 157 331 158 332 
<< m1 >>
rect 158 331 159 332 
<< m1 >>
rect 159 331 160 332 
<< m1 >>
rect 160 331 161 332 
<< m1 >>
rect 163 331 164 332 
<< m1 >>
rect 172 331 173 332 
<< m1 >>
rect 190 331 191 332 
<< m1 >>
rect 208 331 209 332 
<< m1 >>
rect 217 331 218 332 
<< m1 >>
rect 244 331 245 332 
<< m1 >>
rect 253 331 254 332 
<< m1 >>
rect 257 331 258 332 
<< m1 >>
rect 259 331 260 332 
<< m1 >>
rect 260 331 261 332 
<< m1 >>
rect 261 331 262 332 
<< m1 >>
rect 262 331 263 332 
<< m1 >>
rect 263 331 264 332 
<< m1 >>
rect 264 331 265 332 
<< m1 >>
rect 265 331 266 332 
<< m1 >>
rect 266 331 267 332 
<< m1 >>
rect 267 331 268 332 
<< m1 >>
rect 268 331 269 332 
<< m1 >>
rect 269 331 270 332 
<< m1 >>
rect 270 331 271 332 
<< m1 >>
rect 271 331 272 332 
<< m1 >>
rect 272 331 273 332 
<< m1 >>
rect 273 331 274 332 
<< m1 >>
rect 274 331 275 332 
<< m1 >>
rect 275 331 276 332 
<< m1 >>
rect 276 331 277 332 
<< m1 >>
rect 277 331 278 332 
<< m1 >>
rect 278 331 279 332 
<< m1 >>
rect 279 331 280 332 
<< m1 >>
rect 280 331 281 332 
<< m1 >>
rect 281 331 282 332 
<< m1 >>
rect 282 331 283 332 
<< m1 >>
rect 283 331 284 332 
<< m1 >>
rect 284 331 285 332 
<< m1 >>
rect 285 331 286 332 
<< m1 >>
rect 286 331 287 332 
<< m1 >>
rect 289 331 290 332 
<< m1 >>
rect 291 331 292 332 
<< m1 >>
rect 292 331 293 332 
<< m1 >>
rect 293 331 294 332 
<< m1 >>
rect 294 331 295 332 
<< m1 >>
rect 295 331 296 332 
<< m1 >>
rect 296 331 297 332 
<< m1 >>
rect 297 331 298 332 
<< m1 >>
rect 298 331 299 332 
<< m1 >>
rect 299 331 300 332 
<< m1 >>
rect 300 331 301 332 
<< m1 >>
rect 301 331 302 332 
<< m1 >>
rect 302 331 303 332 
<< m1 >>
rect 303 331 304 332 
<< m1 >>
rect 304 331 305 332 
<< m1 >>
rect 305 331 306 332 
<< m1 >>
rect 306 331 307 332 
<< m1 >>
rect 307 331 308 332 
<< m1 >>
rect 308 331 309 332 
<< m1 >>
rect 309 331 310 332 
<< m1 >>
rect 310 331 311 332 
<< m1 >>
rect 311 331 312 332 
<< m1 >>
rect 312 331 313 332 
<< m1 >>
rect 313 331 314 332 
<< m1 >>
rect 314 331 315 332 
<< m1 >>
rect 315 331 316 332 
<< m1 >>
rect 316 331 317 332 
<< m1 >>
rect 317 331 318 332 
<< m1 >>
rect 318 331 319 332 
<< m1 >>
rect 319 331 320 332 
<< m1 >>
rect 320 331 321 332 
<< m2 >>
rect 320 331 321 332 
<< m2c >>
rect 320 331 321 332 
<< m1 >>
rect 320 331 321 332 
<< m2 >>
rect 320 331 321 332 
<< m2 >>
rect 321 331 322 332 
<< m1 >>
rect 322 331 323 332 
<< m2 >>
rect 322 331 323 332 
<< m2 >>
rect 323 331 324 332 
<< m1 >>
rect 324 331 325 332 
<< m2 >>
rect 324 331 325 332 
<< m2c >>
rect 324 331 325 332 
<< m1 >>
rect 324 331 325 332 
<< m2 >>
rect 324 331 325 332 
<< m1 >>
rect 325 331 326 332 
<< m1 >>
rect 326 331 327 332 
<< m1 >>
rect 327 331 328 332 
<< m1 >>
rect 328 331 329 332 
<< m1 >>
rect 329 331 330 332 
<< m1 >>
rect 330 331 331 332 
<< m1 >>
rect 331 331 332 332 
<< m1 >>
rect 332 331 333 332 
<< m1 >>
rect 333 331 334 332 
<< m1 >>
rect 334 331 335 332 
<< m1 >>
rect 335 331 336 332 
<< m1 >>
rect 336 331 337 332 
<< m1 >>
rect 337 331 338 332 
<< m1 >>
rect 338 331 339 332 
<< m1 >>
rect 339 331 340 332 
<< m1 >>
rect 340 331 341 332 
<< m1 >>
rect 355 331 356 332 
<< m1 >>
rect 376 331 377 332 
<< m1 >>
rect 391 331 392 332 
<< m1 >>
rect 73 332 74 333 
<< m1 >>
rect 91 332 92 333 
<< m1 >>
rect 118 332 119 333 
<< m1 >>
rect 127 332 128 333 
<< m1 >>
rect 145 332 146 333 
<< m1 >>
rect 160 332 161 333 
<< m1 >>
rect 163 332 164 333 
<< m1 >>
rect 172 332 173 333 
<< m1 >>
rect 190 332 191 333 
<< m1 >>
rect 208 332 209 333 
<< m1 >>
rect 217 332 218 333 
<< m1 >>
rect 244 332 245 333 
<< m1 >>
rect 253 332 254 333 
<< m1 >>
rect 257 332 258 333 
<< m1 >>
rect 259 332 260 333 
<< m1 >>
rect 286 332 287 333 
<< m1 >>
rect 289 332 290 333 
<< m1 >>
rect 291 332 292 333 
<< m1 >>
rect 322 332 323 333 
<< m1 >>
rect 340 332 341 333 
<< m1 >>
rect 355 332 356 333 
<< m1 >>
rect 376 332 377 333 
<< m1 >>
rect 391 332 392 333 
<< m1 >>
rect 73 333 74 334 
<< m1 >>
rect 91 333 92 334 
<< m1 >>
rect 118 333 119 334 
<< m1 >>
rect 127 333 128 334 
<< m1 >>
rect 145 333 146 334 
<< m1 >>
rect 160 333 161 334 
<< m1 >>
rect 163 333 164 334 
<< m1 >>
rect 172 333 173 334 
<< m1 >>
rect 190 333 191 334 
<< m1 >>
rect 208 333 209 334 
<< m1 >>
rect 217 333 218 334 
<< m1 >>
rect 244 333 245 334 
<< m1 >>
rect 253 333 254 334 
<< m1 >>
rect 257 333 258 334 
<< m1 >>
rect 259 333 260 334 
<< m1 >>
rect 286 333 287 334 
<< m1 >>
rect 289 333 290 334 
<< m1 >>
rect 291 333 292 334 
<< m1 >>
rect 322 333 323 334 
<< m1 >>
rect 340 333 341 334 
<< m1 >>
rect 355 333 356 334 
<< m1 >>
rect 376 333 377 334 
<< m1 >>
rect 391 333 392 334 
<< m1 >>
rect 34 334 35 335 
<< m1 >>
rect 35 334 36 335 
<< m1 >>
rect 36 334 37 335 
<< m1 >>
rect 37 334 38 335 
<< m1 >>
rect 73 334 74 335 
<< m1 >>
rect 91 334 92 335 
<< m1 >>
rect 118 334 119 335 
<< m1 >>
rect 127 334 128 335 
<< m1 >>
rect 145 334 146 335 
<< m1 >>
rect 160 334 161 335 
<< m1 >>
rect 163 334 164 335 
<< m1 >>
rect 172 334 173 335 
<< m1 >>
rect 190 334 191 335 
<< m1 >>
rect 208 334 209 335 
<< m1 >>
rect 217 334 218 335 
<< m1 >>
rect 244 334 245 335 
<< m1 >>
rect 253 334 254 335 
<< m1 >>
rect 257 334 258 335 
<< m1 >>
rect 259 334 260 335 
<< m1 >>
rect 286 334 287 335 
<< m1 >>
rect 289 334 290 335 
<< m1 >>
rect 291 334 292 335 
<< m1 >>
rect 322 334 323 335 
<< m1 >>
rect 340 334 341 335 
<< m1 >>
rect 355 334 356 335 
<< m1 >>
rect 376 334 377 335 
<< m1 >>
rect 391 334 392 335 
<< m1 >>
rect 34 335 35 336 
<< m1 >>
rect 37 335 38 336 
<< m1 >>
rect 73 335 74 336 
<< m1 >>
rect 91 335 92 336 
<< m1 >>
rect 118 335 119 336 
<< m1 >>
rect 127 335 128 336 
<< m1 >>
rect 145 335 146 336 
<< m1 >>
rect 160 335 161 336 
<< m1 >>
rect 163 335 164 336 
<< m1 >>
rect 172 335 173 336 
<< m1 >>
rect 190 335 191 336 
<< m1 >>
rect 208 335 209 336 
<< m1 >>
rect 217 335 218 336 
<< m1 >>
rect 244 335 245 336 
<< m1 >>
rect 253 335 254 336 
<< m1 >>
rect 257 335 258 336 
<< m1 >>
rect 259 335 260 336 
<< m1 >>
rect 286 335 287 336 
<< m1 >>
rect 289 335 290 336 
<< m1 >>
rect 291 335 292 336 
<< m1 >>
rect 322 335 323 336 
<< m1 >>
rect 340 335 341 336 
<< m1 >>
rect 355 335 356 336 
<< m1 >>
rect 376 335 377 336 
<< m1 >>
rect 391 335 392 336 
<< pdiffusion >>
rect 12 336 13 337 
<< pdiffusion >>
rect 13 336 14 337 
<< pdiffusion >>
rect 14 336 15 337 
<< pdiffusion >>
rect 15 336 16 337 
<< pdiffusion >>
rect 16 336 17 337 
<< pdiffusion >>
rect 17 336 18 337 
<< pdiffusion >>
rect 30 336 31 337 
<< pdiffusion >>
rect 31 336 32 337 
<< pdiffusion >>
rect 32 336 33 337 
<< pdiffusion >>
rect 33 336 34 337 
<< m1 >>
rect 34 336 35 337 
<< pdiffusion >>
rect 34 336 35 337 
<< pdiffusion >>
rect 35 336 36 337 
<< m1 >>
rect 37 336 38 337 
<< pdiffusion >>
rect 48 336 49 337 
<< pdiffusion >>
rect 49 336 50 337 
<< pdiffusion >>
rect 50 336 51 337 
<< pdiffusion >>
rect 51 336 52 337 
<< pdiffusion >>
rect 52 336 53 337 
<< pdiffusion >>
rect 53 336 54 337 
<< pdiffusion >>
rect 66 336 67 337 
<< pdiffusion >>
rect 67 336 68 337 
<< pdiffusion >>
rect 68 336 69 337 
<< pdiffusion >>
rect 69 336 70 337 
<< pdiffusion >>
rect 70 336 71 337 
<< pdiffusion >>
rect 71 336 72 337 
<< m1 >>
rect 73 336 74 337 
<< pdiffusion >>
rect 84 336 85 337 
<< pdiffusion >>
rect 85 336 86 337 
<< pdiffusion >>
rect 86 336 87 337 
<< pdiffusion >>
rect 87 336 88 337 
<< pdiffusion >>
rect 88 336 89 337 
<< pdiffusion >>
rect 89 336 90 337 
<< m1 >>
rect 91 336 92 337 
<< pdiffusion >>
rect 102 336 103 337 
<< pdiffusion >>
rect 103 336 104 337 
<< pdiffusion >>
rect 104 336 105 337 
<< pdiffusion >>
rect 105 336 106 337 
<< pdiffusion >>
rect 106 336 107 337 
<< pdiffusion >>
rect 107 336 108 337 
<< m1 >>
rect 118 336 119 337 
<< pdiffusion >>
rect 120 336 121 337 
<< pdiffusion >>
rect 121 336 122 337 
<< pdiffusion >>
rect 122 336 123 337 
<< pdiffusion >>
rect 123 336 124 337 
<< pdiffusion >>
rect 124 336 125 337 
<< pdiffusion >>
rect 125 336 126 337 
<< m1 >>
rect 127 336 128 337 
<< pdiffusion >>
rect 138 336 139 337 
<< pdiffusion >>
rect 139 336 140 337 
<< pdiffusion >>
rect 140 336 141 337 
<< pdiffusion >>
rect 141 336 142 337 
<< pdiffusion >>
rect 142 336 143 337 
<< pdiffusion >>
rect 143 336 144 337 
<< m1 >>
rect 145 336 146 337 
<< pdiffusion >>
rect 156 336 157 337 
<< pdiffusion >>
rect 157 336 158 337 
<< pdiffusion >>
rect 158 336 159 337 
<< pdiffusion >>
rect 159 336 160 337 
<< m1 >>
rect 160 336 161 337 
<< pdiffusion >>
rect 160 336 161 337 
<< pdiffusion >>
rect 161 336 162 337 
<< m1 >>
rect 163 336 164 337 
<< m1 >>
rect 172 336 173 337 
<< pdiffusion >>
rect 174 336 175 337 
<< pdiffusion >>
rect 175 336 176 337 
<< pdiffusion >>
rect 176 336 177 337 
<< pdiffusion >>
rect 177 336 178 337 
<< pdiffusion >>
rect 178 336 179 337 
<< pdiffusion >>
rect 179 336 180 337 
<< m1 >>
rect 190 336 191 337 
<< pdiffusion >>
rect 192 336 193 337 
<< pdiffusion >>
rect 193 336 194 337 
<< pdiffusion >>
rect 194 336 195 337 
<< pdiffusion >>
rect 195 336 196 337 
<< pdiffusion >>
rect 196 336 197 337 
<< pdiffusion >>
rect 197 336 198 337 
<< m1 >>
rect 208 336 209 337 
<< pdiffusion >>
rect 210 336 211 337 
<< pdiffusion >>
rect 211 336 212 337 
<< pdiffusion >>
rect 212 336 213 337 
<< pdiffusion >>
rect 213 336 214 337 
<< pdiffusion >>
rect 214 336 215 337 
<< pdiffusion >>
rect 215 336 216 337 
<< m1 >>
rect 217 336 218 337 
<< pdiffusion >>
rect 228 336 229 337 
<< pdiffusion >>
rect 229 336 230 337 
<< pdiffusion >>
rect 230 336 231 337 
<< pdiffusion >>
rect 231 336 232 337 
<< pdiffusion >>
rect 232 336 233 337 
<< pdiffusion >>
rect 233 336 234 337 
<< m1 >>
rect 244 336 245 337 
<< pdiffusion >>
rect 246 336 247 337 
<< pdiffusion >>
rect 247 336 248 337 
<< pdiffusion >>
rect 248 336 249 337 
<< pdiffusion >>
rect 249 336 250 337 
<< pdiffusion >>
rect 250 336 251 337 
<< pdiffusion >>
rect 251 336 252 337 
<< m1 >>
rect 253 336 254 337 
<< m1 >>
rect 257 336 258 337 
<< m1 >>
rect 259 336 260 337 
<< pdiffusion >>
rect 264 336 265 337 
<< pdiffusion >>
rect 265 336 266 337 
<< pdiffusion >>
rect 266 336 267 337 
<< pdiffusion >>
rect 267 336 268 337 
<< pdiffusion >>
rect 268 336 269 337 
<< pdiffusion >>
rect 269 336 270 337 
<< pdiffusion >>
rect 282 336 283 337 
<< pdiffusion >>
rect 283 336 284 337 
<< pdiffusion >>
rect 284 336 285 337 
<< pdiffusion >>
rect 285 336 286 337 
<< m1 >>
rect 286 336 287 337 
<< pdiffusion >>
rect 286 336 287 337 
<< pdiffusion >>
rect 287 336 288 337 
<< m1 >>
rect 289 336 290 337 
<< m1 >>
rect 291 336 292 337 
<< pdiffusion >>
rect 300 336 301 337 
<< pdiffusion >>
rect 301 336 302 337 
<< pdiffusion >>
rect 302 336 303 337 
<< pdiffusion >>
rect 303 336 304 337 
<< pdiffusion >>
rect 304 336 305 337 
<< pdiffusion >>
rect 305 336 306 337 
<< pdiffusion >>
rect 318 336 319 337 
<< pdiffusion >>
rect 319 336 320 337 
<< pdiffusion >>
rect 320 336 321 337 
<< pdiffusion >>
rect 321 336 322 337 
<< m1 >>
rect 322 336 323 337 
<< pdiffusion >>
rect 322 336 323 337 
<< pdiffusion >>
rect 323 336 324 337 
<< pdiffusion >>
rect 336 336 337 337 
<< pdiffusion >>
rect 337 336 338 337 
<< pdiffusion >>
rect 338 336 339 337 
<< pdiffusion >>
rect 339 336 340 337 
<< m1 >>
rect 340 336 341 337 
<< pdiffusion >>
rect 340 336 341 337 
<< pdiffusion >>
rect 341 336 342 337 
<< pdiffusion >>
rect 354 336 355 337 
<< m1 >>
rect 355 336 356 337 
<< pdiffusion >>
rect 355 336 356 337 
<< pdiffusion >>
rect 356 336 357 337 
<< pdiffusion >>
rect 357 336 358 337 
<< pdiffusion >>
rect 358 336 359 337 
<< pdiffusion >>
rect 359 336 360 337 
<< pdiffusion >>
rect 372 336 373 337 
<< pdiffusion >>
rect 373 336 374 337 
<< pdiffusion >>
rect 374 336 375 337 
<< pdiffusion >>
rect 375 336 376 337 
<< m1 >>
rect 376 336 377 337 
<< pdiffusion >>
rect 376 336 377 337 
<< pdiffusion >>
rect 377 336 378 337 
<< pdiffusion >>
rect 390 336 391 337 
<< m1 >>
rect 391 336 392 337 
<< pdiffusion >>
rect 391 336 392 337 
<< pdiffusion >>
rect 392 336 393 337 
<< pdiffusion >>
rect 393 336 394 337 
<< pdiffusion >>
rect 394 336 395 337 
<< pdiffusion >>
rect 395 336 396 337 
<< pdiffusion >>
rect 408 336 409 337 
<< pdiffusion >>
rect 409 336 410 337 
<< pdiffusion >>
rect 410 336 411 337 
<< pdiffusion >>
rect 411 336 412 337 
<< pdiffusion >>
rect 412 336 413 337 
<< pdiffusion >>
rect 413 336 414 337 
<< pdiffusion >>
rect 426 336 427 337 
<< pdiffusion >>
rect 427 336 428 337 
<< pdiffusion >>
rect 428 336 429 337 
<< pdiffusion >>
rect 429 336 430 337 
<< pdiffusion >>
rect 430 336 431 337 
<< pdiffusion >>
rect 431 336 432 337 
<< pdiffusion >>
rect 444 336 445 337 
<< pdiffusion >>
rect 445 336 446 337 
<< pdiffusion >>
rect 446 336 447 337 
<< pdiffusion >>
rect 447 336 448 337 
<< pdiffusion >>
rect 448 336 449 337 
<< pdiffusion >>
rect 449 336 450 337 
<< pdiffusion >>
rect 12 337 13 338 
<< pdiffusion >>
rect 13 337 14 338 
<< pdiffusion >>
rect 14 337 15 338 
<< pdiffusion >>
rect 15 337 16 338 
<< pdiffusion >>
rect 16 337 17 338 
<< pdiffusion >>
rect 17 337 18 338 
<< pdiffusion >>
rect 30 337 31 338 
<< pdiffusion >>
rect 31 337 32 338 
<< pdiffusion >>
rect 32 337 33 338 
<< pdiffusion >>
rect 33 337 34 338 
<< pdiffusion >>
rect 34 337 35 338 
<< pdiffusion >>
rect 35 337 36 338 
<< m1 >>
rect 37 337 38 338 
<< pdiffusion >>
rect 48 337 49 338 
<< pdiffusion >>
rect 49 337 50 338 
<< pdiffusion >>
rect 50 337 51 338 
<< pdiffusion >>
rect 51 337 52 338 
<< pdiffusion >>
rect 52 337 53 338 
<< pdiffusion >>
rect 53 337 54 338 
<< pdiffusion >>
rect 66 337 67 338 
<< pdiffusion >>
rect 67 337 68 338 
<< pdiffusion >>
rect 68 337 69 338 
<< pdiffusion >>
rect 69 337 70 338 
<< pdiffusion >>
rect 70 337 71 338 
<< pdiffusion >>
rect 71 337 72 338 
<< m1 >>
rect 73 337 74 338 
<< pdiffusion >>
rect 84 337 85 338 
<< pdiffusion >>
rect 85 337 86 338 
<< pdiffusion >>
rect 86 337 87 338 
<< pdiffusion >>
rect 87 337 88 338 
<< pdiffusion >>
rect 88 337 89 338 
<< pdiffusion >>
rect 89 337 90 338 
<< m1 >>
rect 91 337 92 338 
<< pdiffusion >>
rect 102 337 103 338 
<< pdiffusion >>
rect 103 337 104 338 
<< pdiffusion >>
rect 104 337 105 338 
<< pdiffusion >>
rect 105 337 106 338 
<< pdiffusion >>
rect 106 337 107 338 
<< pdiffusion >>
rect 107 337 108 338 
<< m1 >>
rect 118 337 119 338 
<< pdiffusion >>
rect 120 337 121 338 
<< pdiffusion >>
rect 121 337 122 338 
<< pdiffusion >>
rect 122 337 123 338 
<< pdiffusion >>
rect 123 337 124 338 
<< pdiffusion >>
rect 124 337 125 338 
<< pdiffusion >>
rect 125 337 126 338 
<< m1 >>
rect 127 337 128 338 
<< pdiffusion >>
rect 138 337 139 338 
<< pdiffusion >>
rect 139 337 140 338 
<< pdiffusion >>
rect 140 337 141 338 
<< pdiffusion >>
rect 141 337 142 338 
<< pdiffusion >>
rect 142 337 143 338 
<< pdiffusion >>
rect 143 337 144 338 
<< m1 >>
rect 145 337 146 338 
<< pdiffusion >>
rect 156 337 157 338 
<< pdiffusion >>
rect 157 337 158 338 
<< pdiffusion >>
rect 158 337 159 338 
<< pdiffusion >>
rect 159 337 160 338 
<< pdiffusion >>
rect 160 337 161 338 
<< pdiffusion >>
rect 161 337 162 338 
<< m1 >>
rect 163 337 164 338 
<< m1 >>
rect 172 337 173 338 
<< pdiffusion >>
rect 174 337 175 338 
<< pdiffusion >>
rect 175 337 176 338 
<< pdiffusion >>
rect 176 337 177 338 
<< pdiffusion >>
rect 177 337 178 338 
<< pdiffusion >>
rect 178 337 179 338 
<< pdiffusion >>
rect 179 337 180 338 
<< m1 >>
rect 190 337 191 338 
<< pdiffusion >>
rect 192 337 193 338 
<< pdiffusion >>
rect 193 337 194 338 
<< pdiffusion >>
rect 194 337 195 338 
<< pdiffusion >>
rect 195 337 196 338 
<< pdiffusion >>
rect 196 337 197 338 
<< pdiffusion >>
rect 197 337 198 338 
<< m1 >>
rect 208 337 209 338 
<< pdiffusion >>
rect 210 337 211 338 
<< pdiffusion >>
rect 211 337 212 338 
<< pdiffusion >>
rect 212 337 213 338 
<< pdiffusion >>
rect 213 337 214 338 
<< pdiffusion >>
rect 214 337 215 338 
<< pdiffusion >>
rect 215 337 216 338 
<< m1 >>
rect 217 337 218 338 
<< pdiffusion >>
rect 228 337 229 338 
<< pdiffusion >>
rect 229 337 230 338 
<< pdiffusion >>
rect 230 337 231 338 
<< pdiffusion >>
rect 231 337 232 338 
<< pdiffusion >>
rect 232 337 233 338 
<< pdiffusion >>
rect 233 337 234 338 
<< m1 >>
rect 244 337 245 338 
<< pdiffusion >>
rect 246 337 247 338 
<< pdiffusion >>
rect 247 337 248 338 
<< pdiffusion >>
rect 248 337 249 338 
<< pdiffusion >>
rect 249 337 250 338 
<< pdiffusion >>
rect 250 337 251 338 
<< pdiffusion >>
rect 251 337 252 338 
<< m1 >>
rect 253 337 254 338 
<< m1 >>
rect 257 337 258 338 
<< m1 >>
rect 259 337 260 338 
<< pdiffusion >>
rect 264 337 265 338 
<< pdiffusion >>
rect 265 337 266 338 
<< pdiffusion >>
rect 266 337 267 338 
<< pdiffusion >>
rect 267 337 268 338 
<< pdiffusion >>
rect 268 337 269 338 
<< pdiffusion >>
rect 269 337 270 338 
<< pdiffusion >>
rect 282 337 283 338 
<< pdiffusion >>
rect 283 337 284 338 
<< pdiffusion >>
rect 284 337 285 338 
<< pdiffusion >>
rect 285 337 286 338 
<< pdiffusion >>
rect 286 337 287 338 
<< pdiffusion >>
rect 287 337 288 338 
<< m1 >>
rect 289 337 290 338 
<< m1 >>
rect 291 337 292 338 
<< pdiffusion >>
rect 300 337 301 338 
<< pdiffusion >>
rect 301 337 302 338 
<< pdiffusion >>
rect 302 337 303 338 
<< pdiffusion >>
rect 303 337 304 338 
<< pdiffusion >>
rect 304 337 305 338 
<< pdiffusion >>
rect 305 337 306 338 
<< pdiffusion >>
rect 318 337 319 338 
<< pdiffusion >>
rect 319 337 320 338 
<< pdiffusion >>
rect 320 337 321 338 
<< pdiffusion >>
rect 321 337 322 338 
<< pdiffusion >>
rect 322 337 323 338 
<< pdiffusion >>
rect 323 337 324 338 
<< pdiffusion >>
rect 336 337 337 338 
<< pdiffusion >>
rect 337 337 338 338 
<< pdiffusion >>
rect 338 337 339 338 
<< pdiffusion >>
rect 339 337 340 338 
<< pdiffusion >>
rect 340 337 341 338 
<< pdiffusion >>
rect 341 337 342 338 
<< pdiffusion >>
rect 354 337 355 338 
<< pdiffusion >>
rect 355 337 356 338 
<< pdiffusion >>
rect 356 337 357 338 
<< pdiffusion >>
rect 357 337 358 338 
<< pdiffusion >>
rect 358 337 359 338 
<< pdiffusion >>
rect 359 337 360 338 
<< pdiffusion >>
rect 372 337 373 338 
<< pdiffusion >>
rect 373 337 374 338 
<< pdiffusion >>
rect 374 337 375 338 
<< pdiffusion >>
rect 375 337 376 338 
<< pdiffusion >>
rect 376 337 377 338 
<< pdiffusion >>
rect 377 337 378 338 
<< pdiffusion >>
rect 390 337 391 338 
<< pdiffusion >>
rect 391 337 392 338 
<< pdiffusion >>
rect 392 337 393 338 
<< pdiffusion >>
rect 393 337 394 338 
<< pdiffusion >>
rect 394 337 395 338 
<< pdiffusion >>
rect 395 337 396 338 
<< pdiffusion >>
rect 408 337 409 338 
<< pdiffusion >>
rect 409 337 410 338 
<< pdiffusion >>
rect 410 337 411 338 
<< pdiffusion >>
rect 411 337 412 338 
<< pdiffusion >>
rect 412 337 413 338 
<< pdiffusion >>
rect 413 337 414 338 
<< pdiffusion >>
rect 426 337 427 338 
<< pdiffusion >>
rect 427 337 428 338 
<< pdiffusion >>
rect 428 337 429 338 
<< pdiffusion >>
rect 429 337 430 338 
<< pdiffusion >>
rect 430 337 431 338 
<< pdiffusion >>
rect 431 337 432 338 
<< pdiffusion >>
rect 444 337 445 338 
<< pdiffusion >>
rect 445 337 446 338 
<< pdiffusion >>
rect 446 337 447 338 
<< pdiffusion >>
rect 447 337 448 338 
<< pdiffusion >>
rect 448 337 449 338 
<< pdiffusion >>
rect 449 337 450 338 
<< pdiffusion >>
rect 12 338 13 339 
<< pdiffusion >>
rect 13 338 14 339 
<< pdiffusion >>
rect 14 338 15 339 
<< pdiffusion >>
rect 15 338 16 339 
<< pdiffusion >>
rect 16 338 17 339 
<< pdiffusion >>
rect 17 338 18 339 
<< pdiffusion >>
rect 30 338 31 339 
<< pdiffusion >>
rect 31 338 32 339 
<< pdiffusion >>
rect 32 338 33 339 
<< pdiffusion >>
rect 33 338 34 339 
<< pdiffusion >>
rect 34 338 35 339 
<< pdiffusion >>
rect 35 338 36 339 
<< m1 >>
rect 37 338 38 339 
<< pdiffusion >>
rect 48 338 49 339 
<< pdiffusion >>
rect 49 338 50 339 
<< pdiffusion >>
rect 50 338 51 339 
<< pdiffusion >>
rect 51 338 52 339 
<< pdiffusion >>
rect 52 338 53 339 
<< pdiffusion >>
rect 53 338 54 339 
<< pdiffusion >>
rect 66 338 67 339 
<< pdiffusion >>
rect 67 338 68 339 
<< pdiffusion >>
rect 68 338 69 339 
<< pdiffusion >>
rect 69 338 70 339 
<< pdiffusion >>
rect 70 338 71 339 
<< pdiffusion >>
rect 71 338 72 339 
<< m1 >>
rect 73 338 74 339 
<< pdiffusion >>
rect 84 338 85 339 
<< pdiffusion >>
rect 85 338 86 339 
<< pdiffusion >>
rect 86 338 87 339 
<< pdiffusion >>
rect 87 338 88 339 
<< pdiffusion >>
rect 88 338 89 339 
<< pdiffusion >>
rect 89 338 90 339 
<< m1 >>
rect 91 338 92 339 
<< pdiffusion >>
rect 102 338 103 339 
<< pdiffusion >>
rect 103 338 104 339 
<< pdiffusion >>
rect 104 338 105 339 
<< pdiffusion >>
rect 105 338 106 339 
<< pdiffusion >>
rect 106 338 107 339 
<< pdiffusion >>
rect 107 338 108 339 
<< m1 >>
rect 118 338 119 339 
<< pdiffusion >>
rect 120 338 121 339 
<< pdiffusion >>
rect 121 338 122 339 
<< pdiffusion >>
rect 122 338 123 339 
<< pdiffusion >>
rect 123 338 124 339 
<< pdiffusion >>
rect 124 338 125 339 
<< pdiffusion >>
rect 125 338 126 339 
<< m1 >>
rect 127 338 128 339 
<< pdiffusion >>
rect 138 338 139 339 
<< pdiffusion >>
rect 139 338 140 339 
<< pdiffusion >>
rect 140 338 141 339 
<< pdiffusion >>
rect 141 338 142 339 
<< pdiffusion >>
rect 142 338 143 339 
<< pdiffusion >>
rect 143 338 144 339 
<< m1 >>
rect 145 338 146 339 
<< pdiffusion >>
rect 156 338 157 339 
<< pdiffusion >>
rect 157 338 158 339 
<< pdiffusion >>
rect 158 338 159 339 
<< pdiffusion >>
rect 159 338 160 339 
<< pdiffusion >>
rect 160 338 161 339 
<< pdiffusion >>
rect 161 338 162 339 
<< m1 >>
rect 163 338 164 339 
<< m1 >>
rect 172 338 173 339 
<< pdiffusion >>
rect 174 338 175 339 
<< pdiffusion >>
rect 175 338 176 339 
<< pdiffusion >>
rect 176 338 177 339 
<< pdiffusion >>
rect 177 338 178 339 
<< pdiffusion >>
rect 178 338 179 339 
<< pdiffusion >>
rect 179 338 180 339 
<< m1 >>
rect 190 338 191 339 
<< pdiffusion >>
rect 192 338 193 339 
<< pdiffusion >>
rect 193 338 194 339 
<< pdiffusion >>
rect 194 338 195 339 
<< pdiffusion >>
rect 195 338 196 339 
<< pdiffusion >>
rect 196 338 197 339 
<< pdiffusion >>
rect 197 338 198 339 
<< m1 >>
rect 208 338 209 339 
<< pdiffusion >>
rect 210 338 211 339 
<< pdiffusion >>
rect 211 338 212 339 
<< pdiffusion >>
rect 212 338 213 339 
<< pdiffusion >>
rect 213 338 214 339 
<< pdiffusion >>
rect 214 338 215 339 
<< pdiffusion >>
rect 215 338 216 339 
<< m1 >>
rect 217 338 218 339 
<< pdiffusion >>
rect 228 338 229 339 
<< pdiffusion >>
rect 229 338 230 339 
<< pdiffusion >>
rect 230 338 231 339 
<< pdiffusion >>
rect 231 338 232 339 
<< pdiffusion >>
rect 232 338 233 339 
<< pdiffusion >>
rect 233 338 234 339 
<< m1 >>
rect 244 338 245 339 
<< pdiffusion >>
rect 246 338 247 339 
<< pdiffusion >>
rect 247 338 248 339 
<< pdiffusion >>
rect 248 338 249 339 
<< pdiffusion >>
rect 249 338 250 339 
<< pdiffusion >>
rect 250 338 251 339 
<< pdiffusion >>
rect 251 338 252 339 
<< m1 >>
rect 253 338 254 339 
<< m1 >>
rect 257 338 258 339 
<< m1 >>
rect 259 338 260 339 
<< pdiffusion >>
rect 264 338 265 339 
<< pdiffusion >>
rect 265 338 266 339 
<< pdiffusion >>
rect 266 338 267 339 
<< pdiffusion >>
rect 267 338 268 339 
<< pdiffusion >>
rect 268 338 269 339 
<< pdiffusion >>
rect 269 338 270 339 
<< pdiffusion >>
rect 282 338 283 339 
<< pdiffusion >>
rect 283 338 284 339 
<< pdiffusion >>
rect 284 338 285 339 
<< pdiffusion >>
rect 285 338 286 339 
<< pdiffusion >>
rect 286 338 287 339 
<< pdiffusion >>
rect 287 338 288 339 
<< m1 >>
rect 289 338 290 339 
<< m1 >>
rect 291 338 292 339 
<< pdiffusion >>
rect 300 338 301 339 
<< pdiffusion >>
rect 301 338 302 339 
<< pdiffusion >>
rect 302 338 303 339 
<< pdiffusion >>
rect 303 338 304 339 
<< pdiffusion >>
rect 304 338 305 339 
<< pdiffusion >>
rect 305 338 306 339 
<< pdiffusion >>
rect 318 338 319 339 
<< pdiffusion >>
rect 319 338 320 339 
<< pdiffusion >>
rect 320 338 321 339 
<< pdiffusion >>
rect 321 338 322 339 
<< pdiffusion >>
rect 322 338 323 339 
<< pdiffusion >>
rect 323 338 324 339 
<< pdiffusion >>
rect 336 338 337 339 
<< pdiffusion >>
rect 337 338 338 339 
<< pdiffusion >>
rect 338 338 339 339 
<< pdiffusion >>
rect 339 338 340 339 
<< pdiffusion >>
rect 340 338 341 339 
<< pdiffusion >>
rect 341 338 342 339 
<< pdiffusion >>
rect 354 338 355 339 
<< pdiffusion >>
rect 355 338 356 339 
<< pdiffusion >>
rect 356 338 357 339 
<< pdiffusion >>
rect 357 338 358 339 
<< pdiffusion >>
rect 358 338 359 339 
<< pdiffusion >>
rect 359 338 360 339 
<< pdiffusion >>
rect 372 338 373 339 
<< pdiffusion >>
rect 373 338 374 339 
<< pdiffusion >>
rect 374 338 375 339 
<< pdiffusion >>
rect 375 338 376 339 
<< pdiffusion >>
rect 376 338 377 339 
<< pdiffusion >>
rect 377 338 378 339 
<< pdiffusion >>
rect 390 338 391 339 
<< pdiffusion >>
rect 391 338 392 339 
<< pdiffusion >>
rect 392 338 393 339 
<< pdiffusion >>
rect 393 338 394 339 
<< pdiffusion >>
rect 394 338 395 339 
<< pdiffusion >>
rect 395 338 396 339 
<< pdiffusion >>
rect 408 338 409 339 
<< pdiffusion >>
rect 409 338 410 339 
<< pdiffusion >>
rect 410 338 411 339 
<< pdiffusion >>
rect 411 338 412 339 
<< pdiffusion >>
rect 412 338 413 339 
<< pdiffusion >>
rect 413 338 414 339 
<< pdiffusion >>
rect 426 338 427 339 
<< pdiffusion >>
rect 427 338 428 339 
<< pdiffusion >>
rect 428 338 429 339 
<< pdiffusion >>
rect 429 338 430 339 
<< pdiffusion >>
rect 430 338 431 339 
<< pdiffusion >>
rect 431 338 432 339 
<< pdiffusion >>
rect 444 338 445 339 
<< pdiffusion >>
rect 445 338 446 339 
<< pdiffusion >>
rect 446 338 447 339 
<< pdiffusion >>
rect 447 338 448 339 
<< pdiffusion >>
rect 448 338 449 339 
<< pdiffusion >>
rect 449 338 450 339 
<< pdiffusion >>
rect 12 339 13 340 
<< pdiffusion >>
rect 13 339 14 340 
<< pdiffusion >>
rect 14 339 15 340 
<< pdiffusion >>
rect 15 339 16 340 
<< pdiffusion >>
rect 16 339 17 340 
<< pdiffusion >>
rect 17 339 18 340 
<< pdiffusion >>
rect 30 339 31 340 
<< pdiffusion >>
rect 31 339 32 340 
<< pdiffusion >>
rect 32 339 33 340 
<< pdiffusion >>
rect 33 339 34 340 
<< pdiffusion >>
rect 34 339 35 340 
<< pdiffusion >>
rect 35 339 36 340 
<< m1 >>
rect 37 339 38 340 
<< pdiffusion >>
rect 48 339 49 340 
<< pdiffusion >>
rect 49 339 50 340 
<< pdiffusion >>
rect 50 339 51 340 
<< pdiffusion >>
rect 51 339 52 340 
<< pdiffusion >>
rect 52 339 53 340 
<< pdiffusion >>
rect 53 339 54 340 
<< pdiffusion >>
rect 66 339 67 340 
<< pdiffusion >>
rect 67 339 68 340 
<< pdiffusion >>
rect 68 339 69 340 
<< pdiffusion >>
rect 69 339 70 340 
<< pdiffusion >>
rect 70 339 71 340 
<< pdiffusion >>
rect 71 339 72 340 
<< m1 >>
rect 73 339 74 340 
<< pdiffusion >>
rect 84 339 85 340 
<< pdiffusion >>
rect 85 339 86 340 
<< pdiffusion >>
rect 86 339 87 340 
<< pdiffusion >>
rect 87 339 88 340 
<< pdiffusion >>
rect 88 339 89 340 
<< pdiffusion >>
rect 89 339 90 340 
<< m1 >>
rect 91 339 92 340 
<< pdiffusion >>
rect 102 339 103 340 
<< pdiffusion >>
rect 103 339 104 340 
<< pdiffusion >>
rect 104 339 105 340 
<< pdiffusion >>
rect 105 339 106 340 
<< pdiffusion >>
rect 106 339 107 340 
<< pdiffusion >>
rect 107 339 108 340 
<< m1 >>
rect 118 339 119 340 
<< pdiffusion >>
rect 120 339 121 340 
<< pdiffusion >>
rect 121 339 122 340 
<< pdiffusion >>
rect 122 339 123 340 
<< pdiffusion >>
rect 123 339 124 340 
<< pdiffusion >>
rect 124 339 125 340 
<< pdiffusion >>
rect 125 339 126 340 
<< m1 >>
rect 127 339 128 340 
<< pdiffusion >>
rect 138 339 139 340 
<< pdiffusion >>
rect 139 339 140 340 
<< pdiffusion >>
rect 140 339 141 340 
<< pdiffusion >>
rect 141 339 142 340 
<< pdiffusion >>
rect 142 339 143 340 
<< pdiffusion >>
rect 143 339 144 340 
<< m1 >>
rect 145 339 146 340 
<< pdiffusion >>
rect 156 339 157 340 
<< pdiffusion >>
rect 157 339 158 340 
<< pdiffusion >>
rect 158 339 159 340 
<< pdiffusion >>
rect 159 339 160 340 
<< pdiffusion >>
rect 160 339 161 340 
<< pdiffusion >>
rect 161 339 162 340 
<< m1 >>
rect 163 339 164 340 
<< m1 >>
rect 172 339 173 340 
<< pdiffusion >>
rect 174 339 175 340 
<< pdiffusion >>
rect 175 339 176 340 
<< pdiffusion >>
rect 176 339 177 340 
<< pdiffusion >>
rect 177 339 178 340 
<< pdiffusion >>
rect 178 339 179 340 
<< pdiffusion >>
rect 179 339 180 340 
<< m1 >>
rect 190 339 191 340 
<< pdiffusion >>
rect 192 339 193 340 
<< pdiffusion >>
rect 193 339 194 340 
<< pdiffusion >>
rect 194 339 195 340 
<< pdiffusion >>
rect 195 339 196 340 
<< pdiffusion >>
rect 196 339 197 340 
<< pdiffusion >>
rect 197 339 198 340 
<< m1 >>
rect 208 339 209 340 
<< pdiffusion >>
rect 210 339 211 340 
<< pdiffusion >>
rect 211 339 212 340 
<< pdiffusion >>
rect 212 339 213 340 
<< pdiffusion >>
rect 213 339 214 340 
<< pdiffusion >>
rect 214 339 215 340 
<< pdiffusion >>
rect 215 339 216 340 
<< m1 >>
rect 217 339 218 340 
<< pdiffusion >>
rect 228 339 229 340 
<< pdiffusion >>
rect 229 339 230 340 
<< pdiffusion >>
rect 230 339 231 340 
<< pdiffusion >>
rect 231 339 232 340 
<< pdiffusion >>
rect 232 339 233 340 
<< pdiffusion >>
rect 233 339 234 340 
<< m1 >>
rect 244 339 245 340 
<< pdiffusion >>
rect 246 339 247 340 
<< pdiffusion >>
rect 247 339 248 340 
<< pdiffusion >>
rect 248 339 249 340 
<< pdiffusion >>
rect 249 339 250 340 
<< pdiffusion >>
rect 250 339 251 340 
<< pdiffusion >>
rect 251 339 252 340 
<< m1 >>
rect 253 339 254 340 
<< m1 >>
rect 257 339 258 340 
<< m1 >>
rect 259 339 260 340 
<< pdiffusion >>
rect 264 339 265 340 
<< pdiffusion >>
rect 265 339 266 340 
<< pdiffusion >>
rect 266 339 267 340 
<< pdiffusion >>
rect 267 339 268 340 
<< pdiffusion >>
rect 268 339 269 340 
<< pdiffusion >>
rect 269 339 270 340 
<< pdiffusion >>
rect 282 339 283 340 
<< pdiffusion >>
rect 283 339 284 340 
<< pdiffusion >>
rect 284 339 285 340 
<< pdiffusion >>
rect 285 339 286 340 
<< pdiffusion >>
rect 286 339 287 340 
<< pdiffusion >>
rect 287 339 288 340 
<< m1 >>
rect 289 339 290 340 
<< m1 >>
rect 291 339 292 340 
<< pdiffusion >>
rect 300 339 301 340 
<< pdiffusion >>
rect 301 339 302 340 
<< pdiffusion >>
rect 302 339 303 340 
<< pdiffusion >>
rect 303 339 304 340 
<< pdiffusion >>
rect 304 339 305 340 
<< pdiffusion >>
rect 305 339 306 340 
<< pdiffusion >>
rect 318 339 319 340 
<< pdiffusion >>
rect 319 339 320 340 
<< pdiffusion >>
rect 320 339 321 340 
<< pdiffusion >>
rect 321 339 322 340 
<< pdiffusion >>
rect 322 339 323 340 
<< pdiffusion >>
rect 323 339 324 340 
<< pdiffusion >>
rect 336 339 337 340 
<< pdiffusion >>
rect 337 339 338 340 
<< pdiffusion >>
rect 338 339 339 340 
<< pdiffusion >>
rect 339 339 340 340 
<< pdiffusion >>
rect 340 339 341 340 
<< pdiffusion >>
rect 341 339 342 340 
<< pdiffusion >>
rect 354 339 355 340 
<< pdiffusion >>
rect 355 339 356 340 
<< pdiffusion >>
rect 356 339 357 340 
<< pdiffusion >>
rect 357 339 358 340 
<< pdiffusion >>
rect 358 339 359 340 
<< pdiffusion >>
rect 359 339 360 340 
<< pdiffusion >>
rect 372 339 373 340 
<< pdiffusion >>
rect 373 339 374 340 
<< pdiffusion >>
rect 374 339 375 340 
<< pdiffusion >>
rect 375 339 376 340 
<< pdiffusion >>
rect 376 339 377 340 
<< pdiffusion >>
rect 377 339 378 340 
<< pdiffusion >>
rect 390 339 391 340 
<< pdiffusion >>
rect 391 339 392 340 
<< pdiffusion >>
rect 392 339 393 340 
<< pdiffusion >>
rect 393 339 394 340 
<< pdiffusion >>
rect 394 339 395 340 
<< pdiffusion >>
rect 395 339 396 340 
<< pdiffusion >>
rect 408 339 409 340 
<< pdiffusion >>
rect 409 339 410 340 
<< pdiffusion >>
rect 410 339 411 340 
<< pdiffusion >>
rect 411 339 412 340 
<< pdiffusion >>
rect 412 339 413 340 
<< pdiffusion >>
rect 413 339 414 340 
<< pdiffusion >>
rect 426 339 427 340 
<< pdiffusion >>
rect 427 339 428 340 
<< pdiffusion >>
rect 428 339 429 340 
<< pdiffusion >>
rect 429 339 430 340 
<< pdiffusion >>
rect 430 339 431 340 
<< pdiffusion >>
rect 431 339 432 340 
<< pdiffusion >>
rect 444 339 445 340 
<< pdiffusion >>
rect 445 339 446 340 
<< pdiffusion >>
rect 446 339 447 340 
<< pdiffusion >>
rect 447 339 448 340 
<< pdiffusion >>
rect 448 339 449 340 
<< pdiffusion >>
rect 449 339 450 340 
<< pdiffusion >>
rect 12 340 13 341 
<< pdiffusion >>
rect 13 340 14 341 
<< pdiffusion >>
rect 14 340 15 341 
<< pdiffusion >>
rect 15 340 16 341 
<< pdiffusion >>
rect 16 340 17 341 
<< pdiffusion >>
rect 17 340 18 341 
<< pdiffusion >>
rect 30 340 31 341 
<< pdiffusion >>
rect 31 340 32 341 
<< pdiffusion >>
rect 32 340 33 341 
<< pdiffusion >>
rect 33 340 34 341 
<< pdiffusion >>
rect 34 340 35 341 
<< pdiffusion >>
rect 35 340 36 341 
<< m1 >>
rect 37 340 38 341 
<< pdiffusion >>
rect 48 340 49 341 
<< pdiffusion >>
rect 49 340 50 341 
<< pdiffusion >>
rect 50 340 51 341 
<< pdiffusion >>
rect 51 340 52 341 
<< pdiffusion >>
rect 52 340 53 341 
<< pdiffusion >>
rect 53 340 54 341 
<< pdiffusion >>
rect 66 340 67 341 
<< pdiffusion >>
rect 67 340 68 341 
<< pdiffusion >>
rect 68 340 69 341 
<< pdiffusion >>
rect 69 340 70 341 
<< pdiffusion >>
rect 70 340 71 341 
<< pdiffusion >>
rect 71 340 72 341 
<< m1 >>
rect 73 340 74 341 
<< pdiffusion >>
rect 84 340 85 341 
<< pdiffusion >>
rect 85 340 86 341 
<< pdiffusion >>
rect 86 340 87 341 
<< pdiffusion >>
rect 87 340 88 341 
<< pdiffusion >>
rect 88 340 89 341 
<< pdiffusion >>
rect 89 340 90 341 
<< m1 >>
rect 91 340 92 341 
<< pdiffusion >>
rect 102 340 103 341 
<< pdiffusion >>
rect 103 340 104 341 
<< pdiffusion >>
rect 104 340 105 341 
<< pdiffusion >>
rect 105 340 106 341 
<< pdiffusion >>
rect 106 340 107 341 
<< pdiffusion >>
rect 107 340 108 341 
<< m1 >>
rect 118 340 119 341 
<< pdiffusion >>
rect 120 340 121 341 
<< pdiffusion >>
rect 121 340 122 341 
<< pdiffusion >>
rect 122 340 123 341 
<< pdiffusion >>
rect 123 340 124 341 
<< pdiffusion >>
rect 124 340 125 341 
<< pdiffusion >>
rect 125 340 126 341 
<< m1 >>
rect 127 340 128 341 
<< pdiffusion >>
rect 138 340 139 341 
<< pdiffusion >>
rect 139 340 140 341 
<< pdiffusion >>
rect 140 340 141 341 
<< pdiffusion >>
rect 141 340 142 341 
<< pdiffusion >>
rect 142 340 143 341 
<< pdiffusion >>
rect 143 340 144 341 
<< m1 >>
rect 145 340 146 341 
<< pdiffusion >>
rect 156 340 157 341 
<< pdiffusion >>
rect 157 340 158 341 
<< pdiffusion >>
rect 158 340 159 341 
<< pdiffusion >>
rect 159 340 160 341 
<< pdiffusion >>
rect 160 340 161 341 
<< pdiffusion >>
rect 161 340 162 341 
<< m1 >>
rect 163 340 164 341 
<< m1 >>
rect 172 340 173 341 
<< pdiffusion >>
rect 174 340 175 341 
<< pdiffusion >>
rect 175 340 176 341 
<< pdiffusion >>
rect 176 340 177 341 
<< pdiffusion >>
rect 177 340 178 341 
<< pdiffusion >>
rect 178 340 179 341 
<< pdiffusion >>
rect 179 340 180 341 
<< m1 >>
rect 190 340 191 341 
<< pdiffusion >>
rect 192 340 193 341 
<< pdiffusion >>
rect 193 340 194 341 
<< pdiffusion >>
rect 194 340 195 341 
<< pdiffusion >>
rect 195 340 196 341 
<< pdiffusion >>
rect 196 340 197 341 
<< pdiffusion >>
rect 197 340 198 341 
<< m1 >>
rect 208 340 209 341 
<< pdiffusion >>
rect 210 340 211 341 
<< pdiffusion >>
rect 211 340 212 341 
<< pdiffusion >>
rect 212 340 213 341 
<< pdiffusion >>
rect 213 340 214 341 
<< pdiffusion >>
rect 214 340 215 341 
<< pdiffusion >>
rect 215 340 216 341 
<< m1 >>
rect 217 340 218 341 
<< pdiffusion >>
rect 228 340 229 341 
<< pdiffusion >>
rect 229 340 230 341 
<< pdiffusion >>
rect 230 340 231 341 
<< pdiffusion >>
rect 231 340 232 341 
<< pdiffusion >>
rect 232 340 233 341 
<< pdiffusion >>
rect 233 340 234 341 
<< m1 >>
rect 244 340 245 341 
<< pdiffusion >>
rect 246 340 247 341 
<< pdiffusion >>
rect 247 340 248 341 
<< pdiffusion >>
rect 248 340 249 341 
<< pdiffusion >>
rect 249 340 250 341 
<< pdiffusion >>
rect 250 340 251 341 
<< pdiffusion >>
rect 251 340 252 341 
<< m1 >>
rect 253 340 254 341 
<< m1 >>
rect 257 340 258 341 
<< m1 >>
rect 259 340 260 341 
<< pdiffusion >>
rect 264 340 265 341 
<< pdiffusion >>
rect 265 340 266 341 
<< pdiffusion >>
rect 266 340 267 341 
<< pdiffusion >>
rect 267 340 268 341 
<< pdiffusion >>
rect 268 340 269 341 
<< pdiffusion >>
rect 269 340 270 341 
<< pdiffusion >>
rect 282 340 283 341 
<< pdiffusion >>
rect 283 340 284 341 
<< pdiffusion >>
rect 284 340 285 341 
<< pdiffusion >>
rect 285 340 286 341 
<< pdiffusion >>
rect 286 340 287 341 
<< pdiffusion >>
rect 287 340 288 341 
<< m1 >>
rect 289 340 290 341 
<< m1 >>
rect 291 340 292 341 
<< pdiffusion >>
rect 300 340 301 341 
<< pdiffusion >>
rect 301 340 302 341 
<< pdiffusion >>
rect 302 340 303 341 
<< pdiffusion >>
rect 303 340 304 341 
<< pdiffusion >>
rect 304 340 305 341 
<< pdiffusion >>
rect 305 340 306 341 
<< pdiffusion >>
rect 318 340 319 341 
<< pdiffusion >>
rect 319 340 320 341 
<< pdiffusion >>
rect 320 340 321 341 
<< pdiffusion >>
rect 321 340 322 341 
<< pdiffusion >>
rect 322 340 323 341 
<< pdiffusion >>
rect 323 340 324 341 
<< pdiffusion >>
rect 336 340 337 341 
<< pdiffusion >>
rect 337 340 338 341 
<< pdiffusion >>
rect 338 340 339 341 
<< pdiffusion >>
rect 339 340 340 341 
<< pdiffusion >>
rect 340 340 341 341 
<< pdiffusion >>
rect 341 340 342 341 
<< pdiffusion >>
rect 354 340 355 341 
<< pdiffusion >>
rect 355 340 356 341 
<< pdiffusion >>
rect 356 340 357 341 
<< pdiffusion >>
rect 357 340 358 341 
<< pdiffusion >>
rect 358 340 359 341 
<< pdiffusion >>
rect 359 340 360 341 
<< pdiffusion >>
rect 372 340 373 341 
<< pdiffusion >>
rect 373 340 374 341 
<< pdiffusion >>
rect 374 340 375 341 
<< pdiffusion >>
rect 375 340 376 341 
<< pdiffusion >>
rect 376 340 377 341 
<< pdiffusion >>
rect 377 340 378 341 
<< pdiffusion >>
rect 390 340 391 341 
<< pdiffusion >>
rect 391 340 392 341 
<< pdiffusion >>
rect 392 340 393 341 
<< pdiffusion >>
rect 393 340 394 341 
<< pdiffusion >>
rect 394 340 395 341 
<< pdiffusion >>
rect 395 340 396 341 
<< pdiffusion >>
rect 408 340 409 341 
<< pdiffusion >>
rect 409 340 410 341 
<< pdiffusion >>
rect 410 340 411 341 
<< pdiffusion >>
rect 411 340 412 341 
<< pdiffusion >>
rect 412 340 413 341 
<< pdiffusion >>
rect 413 340 414 341 
<< pdiffusion >>
rect 426 340 427 341 
<< pdiffusion >>
rect 427 340 428 341 
<< pdiffusion >>
rect 428 340 429 341 
<< pdiffusion >>
rect 429 340 430 341 
<< pdiffusion >>
rect 430 340 431 341 
<< pdiffusion >>
rect 431 340 432 341 
<< pdiffusion >>
rect 444 340 445 341 
<< pdiffusion >>
rect 445 340 446 341 
<< pdiffusion >>
rect 446 340 447 341 
<< pdiffusion >>
rect 447 340 448 341 
<< pdiffusion >>
rect 448 340 449 341 
<< pdiffusion >>
rect 449 340 450 341 
<< pdiffusion >>
rect 12 341 13 342 
<< pdiffusion >>
rect 13 341 14 342 
<< pdiffusion >>
rect 14 341 15 342 
<< pdiffusion >>
rect 15 341 16 342 
<< pdiffusion >>
rect 16 341 17 342 
<< pdiffusion >>
rect 17 341 18 342 
<< pdiffusion >>
rect 30 341 31 342 
<< pdiffusion >>
rect 31 341 32 342 
<< pdiffusion >>
rect 32 341 33 342 
<< pdiffusion >>
rect 33 341 34 342 
<< pdiffusion >>
rect 34 341 35 342 
<< pdiffusion >>
rect 35 341 36 342 
<< m1 >>
rect 37 341 38 342 
<< pdiffusion >>
rect 48 341 49 342 
<< pdiffusion >>
rect 49 341 50 342 
<< pdiffusion >>
rect 50 341 51 342 
<< pdiffusion >>
rect 51 341 52 342 
<< pdiffusion >>
rect 52 341 53 342 
<< pdiffusion >>
rect 53 341 54 342 
<< pdiffusion >>
rect 66 341 67 342 
<< m1 >>
rect 67 341 68 342 
<< pdiffusion >>
rect 67 341 68 342 
<< pdiffusion >>
rect 68 341 69 342 
<< pdiffusion >>
rect 69 341 70 342 
<< pdiffusion >>
rect 70 341 71 342 
<< pdiffusion >>
rect 71 341 72 342 
<< m1 >>
rect 73 341 74 342 
<< pdiffusion >>
rect 84 341 85 342 
<< pdiffusion >>
rect 85 341 86 342 
<< pdiffusion >>
rect 86 341 87 342 
<< pdiffusion >>
rect 87 341 88 342 
<< pdiffusion >>
rect 88 341 89 342 
<< pdiffusion >>
rect 89 341 90 342 
<< m1 >>
rect 91 341 92 342 
<< pdiffusion >>
rect 102 341 103 342 
<< pdiffusion >>
rect 103 341 104 342 
<< pdiffusion >>
rect 104 341 105 342 
<< pdiffusion >>
rect 105 341 106 342 
<< pdiffusion >>
rect 106 341 107 342 
<< pdiffusion >>
rect 107 341 108 342 
<< m1 >>
rect 118 341 119 342 
<< pdiffusion >>
rect 120 341 121 342 
<< m1 >>
rect 121 341 122 342 
<< pdiffusion >>
rect 121 341 122 342 
<< pdiffusion >>
rect 122 341 123 342 
<< pdiffusion >>
rect 123 341 124 342 
<< m1 >>
rect 124 341 125 342 
<< pdiffusion >>
rect 124 341 125 342 
<< pdiffusion >>
rect 125 341 126 342 
<< m1 >>
rect 127 341 128 342 
<< pdiffusion >>
rect 138 341 139 342 
<< pdiffusion >>
rect 139 341 140 342 
<< pdiffusion >>
rect 140 341 141 342 
<< pdiffusion >>
rect 141 341 142 342 
<< m1 >>
rect 142 341 143 342 
<< pdiffusion >>
rect 142 341 143 342 
<< pdiffusion >>
rect 143 341 144 342 
<< m1 >>
rect 145 341 146 342 
<< pdiffusion >>
rect 156 341 157 342 
<< pdiffusion >>
rect 157 341 158 342 
<< pdiffusion >>
rect 158 341 159 342 
<< pdiffusion >>
rect 159 341 160 342 
<< pdiffusion >>
rect 160 341 161 342 
<< pdiffusion >>
rect 161 341 162 342 
<< m1 >>
rect 163 341 164 342 
<< m1 >>
rect 172 341 173 342 
<< pdiffusion >>
rect 174 341 175 342 
<< m1 >>
rect 175 341 176 342 
<< pdiffusion >>
rect 175 341 176 342 
<< pdiffusion >>
rect 176 341 177 342 
<< pdiffusion >>
rect 177 341 178 342 
<< pdiffusion >>
rect 178 341 179 342 
<< pdiffusion >>
rect 179 341 180 342 
<< m1 >>
rect 190 341 191 342 
<< pdiffusion >>
rect 192 341 193 342 
<< pdiffusion >>
rect 193 341 194 342 
<< pdiffusion >>
rect 194 341 195 342 
<< pdiffusion >>
rect 195 341 196 342 
<< pdiffusion >>
rect 196 341 197 342 
<< pdiffusion >>
rect 197 341 198 342 
<< m1 >>
rect 208 341 209 342 
<< pdiffusion >>
rect 210 341 211 342 
<< m1 >>
rect 211 341 212 342 
<< pdiffusion >>
rect 211 341 212 342 
<< pdiffusion >>
rect 212 341 213 342 
<< pdiffusion >>
rect 213 341 214 342 
<< pdiffusion >>
rect 214 341 215 342 
<< pdiffusion >>
rect 215 341 216 342 
<< m1 >>
rect 217 341 218 342 
<< pdiffusion >>
rect 228 341 229 342 
<< pdiffusion >>
rect 229 341 230 342 
<< pdiffusion >>
rect 230 341 231 342 
<< pdiffusion >>
rect 231 341 232 342 
<< pdiffusion >>
rect 232 341 233 342 
<< pdiffusion >>
rect 233 341 234 342 
<< m1 >>
rect 244 341 245 342 
<< pdiffusion >>
rect 246 341 247 342 
<< pdiffusion >>
rect 247 341 248 342 
<< pdiffusion >>
rect 248 341 249 342 
<< pdiffusion >>
rect 249 341 250 342 
<< pdiffusion >>
rect 250 341 251 342 
<< pdiffusion >>
rect 251 341 252 342 
<< m1 >>
rect 253 341 254 342 
<< m1 >>
rect 257 341 258 342 
<< m1 >>
rect 259 341 260 342 
<< pdiffusion >>
rect 264 341 265 342 
<< pdiffusion >>
rect 265 341 266 342 
<< pdiffusion >>
rect 266 341 267 342 
<< pdiffusion >>
rect 267 341 268 342 
<< pdiffusion >>
rect 268 341 269 342 
<< pdiffusion >>
rect 269 341 270 342 
<< pdiffusion >>
rect 282 341 283 342 
<< m1 >>
rect 283 341 284 342 
<< pdiffusion >>
rect 283 341 284 342 
<< pdiffusion >>
rect 284 341 285 342 
<< pdiffusion >>
rect 285 341 286 342 
<< pdiffusion >>
rect 286 341 287 342 
<< pdiffusion >>
rect 287 341 288 342 
<< m1 >>
rect 289 341 290 342 
<< m1 >>
rect 291 341 292 342 
<< pdiffusion >>
rect 300 341 301 342 
<< pdiffusion >>
rect 301 341 302 342 
<< pdiffusion >>
rect 302 341 303 342 
<< pdiffusion >>
rect 303 341 304 342 
<< pdiffusion >>
rect 304 341 305 342 
<< pdiffusion >>
rect 305 341 306 342 
<< pdiffusion >>
rect 318 341 319 342 
<< m1 >>
rect 319 341 320 342 
<< pdiffusion >>
rect 319 341 320 342 
<< pdiffusion >>
rect 320 341 321 342 
<< pdiffusion >>
rect 321 341 322 342 
<< pdiffusion >>
rect 322 341 323 342 
<< pdiffusion >>
rect 323 341 324 342 
<< pdiffusion >>
rect 336 341 337 342 
<< m1 >>
rect 337 341 338 342 
<< pdiffusion >>
rect 337 341 338 342 
<< pdiffusion >>
rect 338 341 339 342 
<< pdiffusion >>
rect 339 341 340 342 
<< pdiffusion >>
rect 340 341 341 342 
<< pdiffusion >>
rect 341 341 342 342 
<< pdiffusion >>
rect 354 341 355 342 
<< pdiffusion >>
rect 355 341 356 342 
<< pdiffusion >>
rect 356 341 357 342 
<< pdiffusion >>
rect 357 341 358 342 
<< pdiffusion >>
rect 358 341 359 342 
<< pdiffusion >>
rect 359 341 360 342 
<< pdiffusion >>
rect 372 341 373 342 
<< m1 >>
rect 373 341 374 342 
<< pdiffusion >>
rect 373 341 374 342 
<< pdiffusion >>
rect 374 341 375 342 
<< pdiffusion >>
rect 375 341 376 342 
<< pdiffusion >>
rect 376 341 377 342 
<< pdiffusion >>
rect 377 341 378 342 
<< pdiffusion >>
rect 390 341 391 342 
<< pdiffusion >>
rect 391 341 392 342 
<< pdiffusion >>
rect 392 341 393 342 
<< pdiffusion >>
rect 393 341 394 342 
<< pdiffusion >>
rect 394 341 395 342 
<< pdiffusion >>
rect 395 341 396 342 
<< pdiffusion >>
rect 408 341 409 342 
<< pdiffusion >>
rect 409 341 410 342 
<< pdiffusion >>
rect 410 341 411 342 
<< pdiffusion >>
rect 411 341 412 342 
<< pdiffusion >>
rect 412 341 413 342 
<< pdiffusion >>
rect 413 341 414 342 
<< pdiffusion >>
rect 426 341 427 342 
<< pdiffusion >>
rect 427 341 428 342 
<< pdiffusion >>
rect 428 341 429 342 
<< pdiffusion >>
rect 429 341 430 342 
<< pdiffusion >>
rect 430 341 431 342 
<< pdiffusion >>
rect 431 341 432 342 
<< pdiffusion >>
rect 444 341 445 342 
<< pdiffusion >>
rect 445 341 446 342 
<< pdiffusion >>
rect 446 341 447 342 
<< pdiffusion >>
rect 447 341 448 342 
<< pdiffusion >>
rect 448 341 449 342 
<< pdiffusion >>
rect 449 341 450 342 
<< m1 >>
rect 37 342 38 343 
<< m1 >>
rect 67 342 68 343 
<< m1 >>
rect 73 342 74 343 
<< m1 >>
rect 91 342 92 343 
<< m1 >>
rect 118 342 119 343 
<< m1 >>
rect 121 342 122 343 
<< m1 >>
rect 124 342 125 343 
<< m1 >>
rect 127 342 128 343 
<< m1 >>
rect 142 342 143 343 
<< m1 >>
rect 145 342 146 343 
<< m1 >>
rect 163 342 164 343 
<< m1 >>
rect 172 342 173 343 
<< m1 >>
rect 175 342 176 343 
<< m1 >>
rect 190 342 191 343 
<< m2 >>
rect 190 342 191 343 
<< m2c >>
rect 190 342 191 343 
<< m1 >>
rect 190 342 191 343 
<< m2 >>
rect 190 342 191 343 
<< m1 >>
rect 208 342 209 343 
<< m1 >>
rect 211 342 212 343 
<< m1 >>
rect 217 342 218 343 
<< m1 >>
rect 244 342 245 343 
<< m1 >>
rect 253 342 254 343 
<< m1 >>
rect 255 342 256 343 
<< m2 >>
rect 255 342 256 343 
<< m2c >>
rect 255 342 256 343 
<< m1 >>
rect 255 342 256 343 
<< m2 >>
rect 255 342 256 343 
<< m2 >>
rect 256 342 257 343 
<< m1 >>
rect 257 342 258 343 
<< m2 >>
rect 257 342 258 343 
<< m2 >>
rect 258 342 259 343 
<< m1 >>
rect 259 342 260 343 
<< m2 >>
rect 259 342 260 343 
<< m2c >>
rect 259 342 260 343 
<< m1 >>
rect 259 342 260 343 
<< m2 >>
rect 259 342 260 343 
<< m1 >>
rect 283 342 284 343 
<< m1 >>
rect 289 342 290 343 
<< m1 >>
rect 291 342 292 343 
<< m1 >>
rect 319 342 320 343 
<< m1 >>
rect 337 342 338 343 
<< m1 >>
rect 373 342 374 343 
<< m1 >>
rect 37 343 38 344 
<< m1 >>
rect 67 343 68 344 
<< m1 >>
rect 73 343 74 344 
<< m1 >>
rect 91 343 92 344 
<< m1 >>
rect 118 343 119 344 
<< m1 >>
rect 119 343 120 344 
<< m1 >>
rect 120 343 121 344 
<< m1 >>
rect 121 343 122 344 
<< m1 >>
rect 124 343 125 344 
<< m1 >>
rect 125 343 126 344 
<< m2 >>
rect 125 343 126 344 
<< m2c >>
rect 125 343 126 344 
<< m1 >>
rect 125 343 126 344 
<< m2 >>
rect 125 343 126 344 
<< m2 >>
rect 126 343 127 344 
<< m1 >>
rect 127 343 128 344 
<< m2 >>
rect 127 343 128 344 
<< m1 >>
rect 142 343 143 344 
<< m1 >>
rect 143 343 144 344 
<< m1 >>
rect 144 343 145 344 
<< m1 >>
rect 145 343 146 344 
<< m1 >>
rect 163 343 164 344 
<< m1 >>
rect 172 343 173 344 
<< m1 >>
rect 175 343 176 344 
<< m2 >>
rect 179 343 180 344 
<< m2 >>
rect 180 343 181 344 
<< m2 >>
rect 181 343 182 344 
<< m2 >>
rect 182 343 183 344 
<< m2 >>
rect 183 343 184 344 
<< m2 >>
rect 184 343 185 344 
<< m2 >>
rect 185 343 186 344 
<< m2 >>
rect 186 343 187 344 
<< m2 >>
rect 187 343 188 344 
<< m2 >>
rect 188 343 189 344 
<< m2 >>
rect 189 343 190 344 
<< m2 >>
rect 190 343 191 344 
<< m1 >>
rect 208 343 209 344 
<< m1 >>
rect 209 343 210 344 
<< m1 >>
rect 210 343 211 344 
<< m1 >>
rect 211 343 212 344 
<< m1 >>
rect 217 343 218 344 
<< m1 >>
rect 244 343 245 344 
<< m1 >>
rect 253 343 254 344 
<< m1 >>
rect 255 343 256 344 
<< m1 >>
rect 257 343 258 344 
<< m1 >>
rect 283 343 284 344 
<< m1 >>
rect 289 343 290 344 
<< m1 >>
rect 291 343 292 344 
<< m1 >>
rect 319 343 320 344 
<< m2 >>
rect 326 343 327 344 
<< m1 >>
rect 327 343 328 344 
<< m2 >>
rect 327 343 328 344 
<< m2c >>
rect 327 343 328 344 
<< m1 >>
rect 327 343 328 344 
<< m2 >>
rect 327 343 328 344 
<< m1 >>
rect 328 343 329 344 
<< m1 >>
rect 329 343 330 344 
<< m1 >>
rect 330 343 331 344 
<< m1 >>
rect 331 343 332 344 
<< m1 >>
rect 332 343 333 344 
<< m1 >>
rect 333 343 334 344 
<< m1 >>
rect 334 343 335 344 
<< m1 >>
rect 335 343 336 344 
<< m1 >>
rect 336 343 337 344 
<< m1 >>
rect 337 343 338 344 
<< m1 >>
rect 373 343 374 344 
<< m1 >>
rect 37 344 38 345 
<< m1 >>
rect 67 344 68 345 
<< m1 >>
rect 68 344 69 345 
<< m1 >>
rect 69 344 70 345 
<< m1 >>
rect 70 344 71 345 
<< m1 >>
rect 71 344 72 345 
<< m1 >>
rect 72 344 73 345 
<< m1 >>
rect 73 344 74 345 
<< m1 >>
rect 91 344 92 345 
<< m1 >>
rect 127 344 128 345 
<< m2 >>
rect 127 344 128 345 
<< m1 >>
rect 163 344 164 345 
<< m1 >>
rect 172 344 173 345 
<< m2 >>
rect 172 344 173 345 
<< m2c >>
rect 172 344 173 345 
<< m1 >>
rect 172 344 173 345 
<< m2 >>
rect 172 344 173 345 
<< m1 >>
rect 175 344 176 345 
<< m1 >>
rect 176 344 177 345 
<< m1 >>
rect 177 344 178 345 
<< m1 >>
rect 178 344 179 345 
<< m1 >>
rect 179 344 180 345 
<< m2 >>
rect 179 344 180 345 
<< m1 >>
rect 180 344 181 345 
<< m1 >>
rect 181 344 182 345 
<< m1 >>
rect 182 344 183 345 
<< m1 >>
rect 183 344 184 345 
<< m1 >>
rect 184 344 185 345 
<< m1 >>
rect 185 344 186 345 
<< m1 >>
rect 186 344 187 345 
<< m1 >>
rect 187 344 188 345 
<< m1 >>
rect 188 344 189 345 
<< m1 >>
rect 189 344 190 345 
<< m1 >>
rect 190 344 191 345 
<< m1 >>
rect 191 344 192 345 
<< m1 >>
rect 192 344 193 345 
<< m1 >>
rect 217 344 218 345 
<< m1 >>
rect 244 344 245 345 
<< m2 >>
rect 244 344 245 345 
<< m2c >>
rect 244 344 245 345 
<< m1 >>
rect 244 344 245 345 
<< m2 >>
rect 244 344 245 345 
<< m1 >>
rect 248 344 249 345 
<< m2 >>
rect 248 344 249 345 
<< m2c >>
rect 248 344 249 345 
<< m1 >>
rect 248 344 249 345 
<< m2 >>
rect 248 344 249 345 
<< m1 >>
rect 249 344 250 345 
<< m1 >>
rect 250 344 251 345 
<< m1 >>
rect 251 344 252 345 
<< m2 >>
rect 251 344 252 345 
<< m2c >>
rect 251 344 252 345 
<< m1 >>
rect 251 344 252 345 
<< m2 >>
rect 251 344 252 345 
<< m2 >>
rect 252 344 253 345 
<< m1 >>
rect 253 344 254 345 
<< m2 >>
rect 253 344 254 345 
<< m2 >>
rect 254 344 255 345 
<< m1 >>
rect 255 344 256 345 
<< m2 >>
rect 255 344 256 345 
<< m2c >>
rect 255 344 256 345 
<< m1 >>
rect 255 344 256 345 
<< m2 >>
rect 255 344 256 345 
<< m1 >>
rect 257 344 258 345 
<< m2 >>
rect 257 344 258 345 
<< m2c >>
rect 257 344 258 345 
<< m1 >>
rect 257 344 258 345 
<< m2 >>
rect 257 344 258 345 
<< m1 >>
rect 283 344 284 345 
<< m2 >>
rect 283 344 284 345 
<< m2c >>
rect 283 344 284 345 
<< m1 >>
rect 283 344 284 345 
<< m2 >>
rect 283 344 284 345 
<< m1 >>
rect 289 344 290 345 
<< m1 >>
rect 291 344 292 345 
<< m1 >>
rect 319 344 320 345 
<< m1 >>
rect 320 344 321 345 
<< m1 >>
rect 321 344 322 345 
<< m1 >>
rect 322 344 323 345 
<< m1 >>
rect 323 344 324 345 
<< m1 >>
rect 324 344 325 345 
<< m1 >>
rect 325 344 326 345 
<< m2 >>
rect 326 344 327 345 
<< m1 >>
rect 373 344 374 345 
<< m1 >>
rect 374 344 375 345 
<< m1 >>
rect 375 344 376 345 
<< m1 >>
rect 376 344 377 345 
<< m1 >>
rect 377 344 378 345 
<< m1 >>
rect 378 344 379 345 
<< m1 >>
rect 379 344 380 345 
<< m1 >>
rect 37 345 38 346 
<< m1 >>
rect 91 345 92 346 
<< m1 >>
rect 127 345 128 346 
<< m2 >>
rect 127 345 128 346 
<< m1 >>
rect 163 345 164 346 
<< m2 >>
rect 172 345 173 346 
<< m2 >>
rect 179 345 180 346 
<< m1 >>
rect 192 345 193 346 
<< m1 >>
rect 217 345 218 346 
<< m2 >>
rect 244 345 245 346 
<< m2 >>
rect 248 345 249 346 
<< m1 >>
rect 253 345 254 346 
<< m2 >>
rect 257 345 258 346 
<< m2 >>
rect 283 345 284 346 
<< m1 >>
rect 289 345 290 346 
<< m1 >>
rect 291 345 292 346 
<< m1 >>
rect 325 345 326 346 
<< m2 >>
rect 326 345 327 346 
<< m1 >>
rect 379 345 380 346 
<< m1 >>
rect 37 346 38 347 
<< m1 >>
rect 91 346 92 347 
<< m1 >>
rect 127 346 128 347 
<< m2 >>
rect 127 346 128 347 
<< m1 >>
rect 163 346 164 347 
<< m1 >>
rect 164 346 165 347 
<< m1 >>
rect 165 346 166 347 
<< m1 >>
rect 166 346 167 347 
<< m1 >>
rect 167 346 168 347 
<< m1 >>
rect 168 346 169 347 
<< m1 >>
rect 169 346 170 347 
<< m1 >>
rect 170 346 171 347 
<< m1 >>
rect 171 346 172 347 
<< m1 >>
rect 172 346 173 347 
<< m2 >>
rect 172 346 173 347 
<< m1 >>
rect 173 346 174 347 
<< m1 >>
rect 174 346 175 347 
<< m1 >>
rect 175 346 176 347 
<< m1 >>
rect 176 346 177 347 
<< m1 >>
rect 177 346 178 347 
<< m1 >>
rect 178 346 179 347 
<< m2 >>
rect 179 346 180 347 
<< m1 >>
rect 192 346 193 347 
<< m1 >>
rect 214 346 215 347 
<< m1 >>
rect 215 346 216 347 
<< m2 >>
rect 215 346 216 347 
<< m2c >>
rect 215 346 216 347 
<< m1 >>
rect 215 346 216 347 
<< m2 >>
rect 215 346 216 347 
<< m2 >>
rect 216 346 217 347 
<< m1 >>
rect 217 346 218 347 
<< m2 >>
rect 217 346 218 347 
<< m2 >>
rect 218 346 219 347 
<< m1 >>
rect 219 346 220 347 
<< m2 >>
rect 219 346 220 347 
<< m2c >>
rect 219 346 220 347 
<< m1 >>
rect 219 346 220 347 
<< m2 >>
rect 219 346 220 347 
<< m1 >>
rect 220 346 221 347 
<< m1 >>
rect 221 346 222 347 
<< m1 >>
rect 222 346 223 347 
<< m1 >>
rect 223 346 224 347 
<< m1 >>
rect 224 346 225 347 
<< m1 >>
rect 225 346 226 347 
<< m1 >>
rect 226 346 227 347 
<< m1 >>
rect 227 346 228 347 
<< m1 >>
rect 228 346 229 347 
<< m1 >>
rect 229 346 230 347 
<< m1 >>
rect 230 346 231 347 
<< m1 >>
rect 231 346 232 347 
<< m1 >>
rect 232 346 233 347 
<< m1 >>
rect 233 346 234 347 
<< m1 >>
rect 234 346 235 347 
<< m1 >>
rect 235 346 236 347 
<< m1 >>
rect 236 346 237 347 
<< m1 >>
rect 237 346 238 347 
<< m1 >>
rect 238 346 239 347 
<< m1 >>
rect 239 346 240 347 
<< m1 >>
rect 240 346 241 347 
<< m1 >>
rect 241 346 242 347 
<< m1 >>
rect 242 346 243 347 
<< m1 >>
rect 243 346 244 347 
<< m1 >>
rect 244 346 245 347 
<< m2 >>
rect 244 346 245 347 
<< m1 >>
rect 245 346 246 347 
<< m1 >>
rect 246 346 247 347 
<< m1 >>
rect 247 346 248 347 
<< m1 >>
rect 248 346 249 347 
<< m2 >>
rect 248 346 249 347 
<< m1 >>
rect 249 346 250 347 
<< m1 >>
rect 250 346 251 347 
<< m1 >>
rect 251 346 252 347 
<< m2 >>
rect 251 346 252 347 
<< m2c >>
rect 251 346 252 347 
<< m1 >>
rect 251 346 252 347 
<< m2 >>
rect 251 346 252 347 
<< m2 >>
rect 252 346 253 347 
<< m1 >>
rect 253 346 254 347 
<< m2 >>
rect 253 346 254 347 
<< m2 >>
rect 254 346 255 347 
<< m1 >>
rect 255 346 256 347 
<< m2 >>
rect 255 346 256 347 
<< m2c >>
rect 255 346 256 347 
<< m1 >>
rect 255 346 256 347 
<< m2 >>
rect 255 346 256 347 
<< m1 >>
rect 256 346 257 347 
<< m1 >>
rect 257 346 258 347 
<< m2 >>
rect 257 346 258 347 
<< m1 >>
rect 258 346 259 347 
<< m1 >>
rect 259 346 260 347 
<< m1 >>
rect 260 346 261 347 
<< m1 >>
rect 261 346 262 347 
<< m1 >>
rect 262 346 263 347 
<< m1 >>
rect 263 346 264 347 
<< m1 >>
rect 264 346 265 347 
<< m1 >>
rect 265 346 266 347 
<< m1 >>
rect 266 346 267 347 
<< m1 >>
rect 267 346 268 347 
<< m1 >>
rect 268 346 269 347 
<< m1 >>
rect 269 346 270 347 
<< m1 >>
rect 270 346 271 347 
<< m1 >>
rect 271 346 272 347 
<< m1 >>
rect 272 346 273 347 
<< m1 >>
rect 273 346 274 347 
<< m1 >>
rect 274 346 275 347 
<< m1 >>
rect 275 346 276 347 
<< m1 >>
rect 276 346 277 347 
<< m1 >>
rect 277 346 278 347 
<< m1 >>
rect 278 346 279 347 
<< m1 >>
rect 279 346 280 347 
<< m1 >>
rect 280 346 281 347 
<< m1 >>
rect 281 346 282 347 
<< m1 >>
rect 282 346 283 347 
<< m1 >>
rect 283 346 284 347 
<< m2 >>
rect 283 346 284 347 
<< m1 >>
rect 284 346 285 347 
<< m1 >>
rect 285 346 286 347 
<< m1 >>
rect 286 346 287 347 
<< m1 >>
rect 287 346 288 347 
<< m2 >>
rect 287 346 288 347 
<< m2c >>
rect 287 346 288 347 
<< m1 >>
rect 287 346 288 347 
<< m2 >>
rect 287 346 288 347 
<< m2 >>
rect 288 346 289 347 
<< m1 >>
rect 289 346 290 347 
<< m2 >>
rect 289 346 290 347 
<< m2 >>
rect 290 346 291 347 
<< m1 >>
rect 291 346 292 347 
<< m2 >>
rect 291 346 292 347 
<< m2 >>
rect 292 346 293 347 
<< m1 >>
rect 293 346 294 347 
<< m2 >>
rect 293 346 294 347 
<< m2c >>
rect 293 346 294 347 
<< m1 >>
rect 293 346 294 347 
<< m2 >>
rect 293 346 294 347 
<< m1 >>
rect 294 346 295 347 
<< m1 >>
rect 295 346 296 347 
<< m1 >>
rect 296 346 297 347 
<< m1 >>
rect 297 346 298 347 
<< m1 >>
rect 298 346 299 347 
<< m1 >>
rect 299 346 300 347 
<< m1 >>
rect 300 346 301 347 
<< m1 >>
rect 301 346 302 347 
<< m1 >>
rect 302 346 303 347 
<< m1 >>
rect 303 346 304 347 
<< m1 >>
rect 304 346 305 347 
<< m1 >>
rect 305 346 306 347 
<< m1 >>
rect 306 346 307 347 
<< m1 >>
rect 307 346 308 347 
<< m1 >>
rect 308 346 309 347 
<< m1 >>
rect 309 346 310 347 
<< m1 >>
rect 310 346 311 347 
<< m1 >>
rect 311 346 312 347 
<< m1 >>
rect 312 346 313 347 
<< m1 >>
rect 313 346 314 347 
<< m1 >>
rect 314 346 315 347 
<< m1 >>
rect 315 346 316 347 
<< m1 >>
rect 316 346 317 347 
<< m1 >>
rect 317 346 318 347 
<< m1 >>
rect 318 346 319 347 
<< m1 >>
rect 319 346 320 347 
<< m1 >>
rect 320 346 321 347 
<< m1 >>
rect 321 346 322 347 
<< m1 >>
rect 322 346 323 347 
<< m1 >>
rect 323 346 324 347 
<< m2 >>
rect 323 346 324 347 
<< m2c >>
rect 323 346 324 347 
<< m1 >>
rect 323 346 324 347 
<< m2 >>
rect 323 346 324 347 
<< m2 >>
rect 324 346 325 347 
<< m1 >>
rect 325 346 326 347 
<< m2 >>
rect 325 346 326 347 
<< m2 >>
rect 326 346 327 347 
<< m1 >>
rect 379 346 380 347 
<< m1 >>
rect 37 347 38 348 
<< m1 >>
rect 91 347 92 348 
<< m1 >>
rect 127 347 128 348 
<< m2 >>
rect 127 347 128 348 
<< m2 >>
rect 172 347 173 348 
<< m1 >>
rect 178 347 179 348 
<< m2 >>
rect 179 347 180 348 
<< m1 >>
rect 192 347 193 348 
<< m1 >>
rect 214 347 215 348 
<< m1 >>
rect 217 347 218 348 
<< m2 >>
rect 244 347 245 348 
<< m2 >>
rect 246 347 247 348 
<< m2 >>
rect 247 347 248 348 
<< m2 >>
rect 248 347 249 348 
<< m1 >>
rect 253 347 254 348 
<< m2 >>
rect 257 347 258 348 
<< m2 >>
rect 283 347 284 348 
<< m1 >>
rect 289 347 290 348 
<< m1 >>
rect 291 347 292 348 
<< m1 >>
rect 325 347 326 348 
<< m1 >>
rect 379 347 380 348 
<< m1 >>
rect 37 348 38 349 
<< m1 >>
rect 91 348 92 349 
<< m1 >>
rect 127 348 128 349 
<< m2 >>
rect 127 348 128 349 
<< m1 >>
rect 172 348 173 349 
<< m2 >>
rect 172 348 173 349 
<< m2c >>
rect 172 348 173 349 
<< m1 >>
rect 172 348 173 349 
<< m2 >>
rect 172 348 173 349 
<< m1 >>
rect 175 348 176 349 
<< m1 >>
rect 176 348 177 349 
<< m2 >>
rect 176 348 177 349 
<< m2c >>
rect 176 348 177 349 
<< m1 >>
rect 176 348 177 349 
<< m2 >>
rect 176 348 177 349 
<< m2 >>
rect 177 348 178 349 
<< m1 >>
rect 178 348 179 349 
<< m2 >>
rect 178 348 179 349 
<< m2 >>
rect 179 348 180 349 
<< m1 >>
rect 192 348 193 349 
<< m1 >>
rect 214 348 215 349 
<< m1 >>
rect 217 348 218 349 
<< m1 >>
rect 244 348 245 349 
<< m2 >>
rect 244 348 245 349 
<< m2c >>
rect 244 348 245 349 
<< m1 >>
rect 244 348 245 349 
<< m2 >>
rect 244 348 245 349 
<< m1 >>
rect 246 348 247 349 
<< m2 >>
rect 246 348 247 349 
<< m2c >>
rect 246 348 247 349 
<< m1 >>
rect 246 348 247 349 
<< m2 >>
rect 246 348 247 349 
<< m1 >>
rect 253 348 254 349 
<< m2 >>
rect 254 348 255 349 
<< m1 >>
rect 255 348 256 349 
<< m2 >>
rect 255 348 256 349 
<< m2c >>
rect 255 348 256 349 
<< m1 >>
rect 255 348 256 349 
<< m2 >>
rect 255 348 256 349 
<< m1 >>
rect 256 348 257 349 
<< m1 >>
rect 257 348 258 349 
<< m2 >>
rect 257 348 258 349 
<< m2c >>
rect 257 348 258 349 
<< m1 >>
rect 257 348 258 349 
<< m2 >>
rect 257 348 258 349 
<< m1 >>
rect 283 348 284 349 
<< m2 >>
rect 283 348 284 349 
<< m2c >>
rect 283 348 284 349 
<< m1 >>
rect 283 348 284 349 
<< m2 >>
rect 283 348 284 349 
<< m1 >>
rect 284 348 285 349 
<< m1 >>
rect 285 348 286 349 
<< m1 >>
rect 286 348 287 349 
<< m1 >>
rect 287 348 288 349 
<< m2 >>
rect 287 348 288 349 
<< m2c >>
rect 287 348 288 349 
<< m1 >>
rect 287 348 288 349 
<< m2 >>
rect 287 348 288 349 
<< m2 >>
rect 288 348 289 349 
<< m1 >>
rect 289 348 290 349 
<< m2 >>
rect 289 348 290 349 
<< m2 >>
rect 290 348 291 349 
<< m1 >>
rect 291 348 292 349 
<< m2 >>
rect 291 348 292 349 
<< m2 >>
rect 292 348 293 349 
<< m1 >>
rect 293 348 294 349 
<< m2 >>
rect 293 348 294 349 
<< m2c >>
rect 293 348 294 349 
<< m1 >>
rect 293 348 294 349 
<< m2 >>
rect 293 348 294 349 
<< m1 >>
rect 325 348 326 349 
<< m1 >>
rect 379 348 380 349 
<< m1 >>
rect 37 349 38 350 
<< m1 >>
rect 91 349 92 350 
<< m1 >>
rect 127 349 128 350 
<< m2 >>
rect 127 349 128 350 
<< m1 >>
rect 172 349 173 350 
<< m1 >>
rect 175 349 176 350 
<< m1 >>
rect 178 349 179 350 
<< m1 >>
rect 192 349 193 350 
<< m1 >>
rect 193 349 194 350 
<< m1 >>
rect 194 349 195 350 
<< m1 >>
rect 195 349 196 350 
<< m1 >>
rect 196 349 197 350 
<< m1 >>
rect 197 349 198 350 
<< m1 >>
rect 198 349 199 350 
<< m1 >>
rect 199 349 200 350 
<< m1 >>
rect 200 349 201 350 
<< m1 >>
rect 201 349 202 350 
<< m1 >>
rect 202 349 203 350 
<< m1 >>
rect 203 349 204 350 
<< m1 >>
rect 204 349 205 350 
<< m1 >>
rect 205 349 206 350 
<< m1 >>
rect 206 349 207 350 
<< m1 >>
rect 207 349 208 350 
<< m1 >>
rect 208 349 209 350 
<< m1 >>
rect 209 349 210 350 
<< m1 >>
rect 210 349 211 350 
<< m1 >>
rect 211 349 212 350 
<< m1 >>
rect 212 349 213 350 
<< m1 >>
rect 214 349 215 350 
<< m1 >>
rect 217 349 218 350 
<< m1 >>
rect 244 349 245 350 
<< m1 >>
rect 246 349 247 350 
<< m1 >>
rect 253 349 254 350 
<< m2 >>
rect 254 349 255 350 
<< m1 >>
rect 289 349 290 350 
<< m1 >>
rect 291 349 292 350 
<< m1 >>
rect 293 349 294 350 
<< m1 >>
rect 325 349 326 350 
<< m1 >>
rect 379 349 380 350 
<< m1 >>
rect 37 350 38 351 
<< m1 >>
rect 91 350 92 351 
<< m1 >>
rect 127 350 128 351 
<< m2 >>
rect 127 350 128 351 
<< m1 >>
rect 172 350 173 351 
<< m1 >>
rect 175 350 176 351 
<< m1 >>
rect 178 350 179 351 
<< m1 >>
rect 212 350 213 351 
<< m1 >>
rect 214 350 215 351 
<< m1 >>
rect 217 350 218 351 
<< m1 >>
rect 244 350 245 351 
<< m1 >>
rect 246 350 247 351 
<< m1 >>
rect 253 350 254 351 
<< m2 >>
rect 254 350 255 351 
<< m1 >>
rect 289 350 290 351 
<< m1 >>
rect 291 350 292 351 
<< m1 >>
rect 293 350 294 351 
<< m1 >>
rect 325 350 326 351 
<< m1 >>
rect 379 350 380 351 
<< m1 >>
rect 37 351 38 352 
<< m1 >>
rect 91 351 92 352 
<< m1 >>
rect 127 351 128 352 
<< m2 >>
rect 127 351 128 352 
<< m1 >>
rect 172 351 173 352 
<< m1 >>
rect 175 351 176 352 
<< m1 >>
rect 178 351 179 352 
<< m1 >>
rect 212 351 213 352 
<< m2 >>
rect 212 351 213 352 
<< m2c >>
rect 212 351 213 352 
<< m1 >>
rect 212 351 213 352 
<< m2 >>
rect 212 351 213 352 
<< m2 >>
rect 213 351 214 352 
<< m1 >>
rect 214 351 215 352 
<< m2 >>
rect 214 351 215 352 
<< m2 >>
rect 215 351 216 352 
<< m2 >>
rect 216 351 217 352 
<< m1 >>
rect 217 351 218 352 
<< m2 >>
rect 217 351 218 352 
<< m2 >>
rect 218 351 219 352 
<< m1 >>
rect 244 351 245 352 
<< m1 >>
rect 246 351 247 352 
<< m1 >>
rect 253 351 254 352 
<< m2 >>
rect 254 351 255 352 
<< m1 >>
rect 289 351 290 352 
<< m1 >>
rect 291 351 292 352 
<< m1 >>
rect 293 351 294 352 
<< m1 >>
rect 325 351 326 352 
<< m1 >>
rect 379 351 380 352 
<< m1 >>
rect 37 352 38 353 
<< m1 >>
rect 91 352 92 353 
<< m1 >>
rect 127 352 128 353 
<< m2 >>
rect 127 352 128 353 
<< m1 >>
rect 172 352 173 353 
<< m1 >>
rect 175 352 176 353 
<< m1 >>
rect 178 352 179 353 
<< m1 >>
rect 214 352 215 353 
<< m1 >>
rect 217 352 218 353 
<< m2 >>
rect 218 352 219 353 
<< m1 >>
rect 219 352 220 353 
<< m2 >>
rect 219 352 220 353 
<< m2c >>
rect 219 352 220 353 
<< m1 >>
rect 219 352 220 353 
<< m2 >>
rect 219 352 220 353 
<< m1 >>
rect 220 352 221 353 
<< m1 >>
rect 221 352 222 353 
<< m1 >>
rect 222 352 223 353 
<< m1 >>
rect 223 352 224 353 
<< m1 >>
rect 224 352 225 353 
<< m1 >>
rect 225 352 226 353 
<< m1 >>
rect 226 352 227 353 
<< m1 >>
rect 227 352 228 353 
<< m1 >>
rect 228 352 229 353 
<< m1 >>
rect 229 352 230 353 
<< m1 >>
rect 232 352 233 353 
<< m1 >>
rect 233 352 234 353 
<< m1 >>
rect 234 352 235 353 
<< m1 >>
rect 235 352 236 353 
<< m1 >>
rect 236 352 237 353 
<< m1 >>
rect 237 352 238 353 
<< m1 >>
rect 238 352 239 353 
<< m1 >>
rect 239 352 240 353 
<< m1 >>
rect 240 352 241 353 
<< m1 >>
rect 241 352 242 353 
<< m1 >>
rect 242 352 243 353 
<< m2 >>
rect 242 352 243 353 
<< m2c >>
rect 242 352 243 353 
<< m1 >>
rect 242 352 243 353 
<< m2 >>
rect 242 352 243 353 
<< m2 >>
rect 243 352 244 353 
<< m1 >>
rect 244 352 245 353 
<< m2 >>
rect 244 352 245 353 
<< m2 >>
rect 245 352 246 353 
<< m1 >>
rect 246 352 247 353 
<< m2 >>
rect 246 352 247 353 
<< m2c >>
rect 246 352 247 353 
<< m1 >>
rect 246 352 247 353 
<< m2 >>
rect 246 352 247 353 
<< m1 >>
rect 253 352 254 353 
<< m2 >>
rect 254 352 255 353 
<< m1 >>
rect 289 352 290 353 
<< m1 >>
rect 291 352 292 353 
<< m1 >>
rect 293 352 294 353 
<< m1 >>
rect 325 352 326 353 
<< m1 >>
rect 379 352 380 353 
<< m1 >>
rect 37 353 38 354 
<< m1 >>
rect 91 353 92 354 
<< m1 >>
rect 127 353 128 354 
<< m2 >>
rect 127 353 128 354 
<< m1 >>
rect 172 353 173 354 
<< m1 >>
rect 175 353 176 354 
<< m1 >>
rect 178 353 179 354 
<< m1 >>
rect 214 353 215 354 
<< m1 >>
rect 217 353 218 354 
<< m1 >>
rect 229 353 230 354 
<< m1 >>
rect 232 353 233 354 
<< m1 >>
rect 244 353 245 354 
<< m1 >>
rect 253 353 254 354 
<< m2 >>
rect 254 353 255 354 
<< m1 >>
rect 289 353 290 354 
<< m1 >>
rect 291 353 292 354 
<< m1 >>
rect 293 353 294 354 
<< m1 >>
rect 325 353 326 354 
<< m1 >>
rect 379 353 380 354 
<< pdiffusion >>
rect 12 354 13 355 
<< pdiffusion >>
rect 13 354 14 355 
<< pdiffusion >>
rect 14 354 15 355 
<< pdiffusion >>
rect 15 354 16 355 
<< pdiffusion >>
rect 16 354 17 355 
<< pdiffusion >>
rect 17 354 18 355 
<< pdiffusion >>
rect 30 354 31 355 
<< pdiffusion >>
rect 31 354 32 355 
<< pdiffusion >>
rect 32 354 33 355 
<< pdiffusion >>
rect 33 354 34 355 
<< pdiffusion >>
rect 34 354 35 355 
<< pdiffusion >>
rect 35 354 36 355 
<< m1 >>
rect 37 354 38 355 
<< pdiffusion >>
rect 48 354 49 355 
<< pdiffusion >>
rect 49 354 50 355 
<< pdiffusion >>
rect 50 354 51 355 
<< pdiffusion >>
rect 51 354 52 355 
<< pdiffusion >>
rect 52 354 53 355 
<< pdiffusion >>
rect 53 354 54 355 
<< pdiffusion >>
rect 66 354 67 355 
<< pdiffusion >>
rect 67 354 68 355 
<< pdiffusion >>
rect 68 354 69 355 
<< pdiffusion >>
rect 69 354 70 355 
<< pdiffusion >>
rect 70 354 71 355 
<< pdiffusion >>
rect 71 354 72 355 
<< pdiffusion >>
rect 84 354 85 355 
<< pdiffusion >>
rect 85 354 86 355 
<< pdiffusion >>
rect 86 354 87 355 
<< pdiffusion >>
rect 87 354 88 355 
<< pdiffusion >>
rect 88 354 89 355 
<< pdiffusion >>
rect 89 354 90 355 
<< m1 >>
rect 91 354 92 355 
<< pdiffusion >>
rect 102 354 103 355 
<< pdiffusion >>
rect 103 354 104 355 
<< pdiffusion >>
rect 104 354 105 355 
<< pdiffusion >>
rect 105 354 106 355 
<< pdiffusion >>
rect 106 354 107 355 
<< pdiffusion >>
rect 107 354 108 355 
<< pdiffusion >>
rect 120 354 121 355 
<< pdiffusion >>
rect 121 354 122 355 
<< pdiffusion >>
rect 122 354 123 355 
<< pdiffusion >>
rect 123 354 124 355 
<< pdiffusion >>
rect 124 354 125 355 
<< pdiffusion >>
rect 125 354 126 355 
<< m1 >>
rect 127 354 128 355 
<< m2 >>
rect 127 354 128 355 
<< pdiffusion >>
rect 138 354 139 355 
<< pdiffusion >>
rect 139 354 140 355 
<< pdiffusion >>
rect 140 354 141 355 
<< pdiffusion >>
rect 141 354 142 355 
<< pdiffusion >>
rect 142 354 143 355 
<< pdiffusion >>
rect 143 354 144 355 
<< pdiffusion >>
rect 156 354 157 355 
<< pdiffusion >>
rect 157 354 158 355 
<< pdiffusion >>
rect 158 354 159 355 
<< pdiffusion >>
rect 159 354 160 355 
<< pdiffusion >>
rect 160 354 161 355 
<< pdiffusion >>
rect 161 354 162 355 
<< m1 >>
rect 172 354 173 355 
<< pdiffusion >>
rect 174 354 175 355 
<< m1 >>
rect 175 354 176 355 
<< pdiffusion >>
rect 175 354 176 355 
<< pdiffusion >>
rect 176 354 177 355 
<< pdiffusion >>
rect 177 354 178 355 
<< m1 >>
rect 178 354 179 355 
<< pdiffusion >>
rect 178 354 179 355 
<< pdiffusion >>
rect 179 354 180 355 
<< pdiffusion >>
rect 192 354 193 355 
<< pdiffusion >>
rect 193 354 194 355 
<< pdiffusion >>
rect 194 354 195 355 
<< pdiffusion >>
rect 195 354 196 355 
<< pdiffusion >>
rect 196 354 197 355 
<< pdiffusion >>
rect 197 354 198 355 
<< pdiffusion >>
rect 210 354 211 355 
<< pdiffusion >>
rect 211 354 212 355 
<< pdiffusion >>
rect 212 354 213 355 
<< pdiffusion >>
rect 213 354 214 355 
<< m1 >>
rect 214 354 215 355 
<< pdiffusion >>
rect 214 354 215 355 
<< pdiffusion >>
rect 215 354 216 355 
<< m1 >>
rect 217 354 218 355 
<< pdiffusion >>
rect 228 354 229 355 
<< m1 >>
rect 229 354 230 355 
<< pdiffusion >>
rect 229 354 230 355 
<< pdiffusion >>
rect 230 354 231 355 
<< pdiffusion >>
rect 231 354 232 355 
<< m1 >>
rect 232 354 233 355 
<< pdiffusion >>
rect 232 354 233 355 
<< pdiffusion >>
rect 233 354 234 355 
<< m1 >>
rect 244 354 245 355 
<< pdiffusion >>
rect 246 354 247 355 
<< pdiffusion >>
rect 247 354 248 355 
<< pdiffusion >>
rect 248 354 249 355 
<< pdiffusion >>
rect 249 354 250 355 
<< pdiffusion >>
rect 250 354 251 355 
<< pdiffusion >>
rect 251 354 252 355 
<< m1 >>
rect 253 354 254 355 
<< m2 >>
rect 254 354 255 355 
<< pdiffusion >>
rect 264 354 265 355 
<< pdiffusion >>
rect 265 354 266 355 
<< pdiffusion >>
rect 266 354 267 355 
<< pdiffusion >>
rect 267 354 268 355 
<< pdiffusion >>
rect 268 354 269 355 
<< pdiffusion >>
rect 269 354 270 355 
<< pdiffusion >>
rect 282 354 283 355 
<< pdiffusion >>
rect 283 354 284 355 
<< pdiffusion >>
rect 284 354 285 355 
<< pdiffusion >>
rect 285 354 286 355 
<< pdiffusion >>
rect 286 354 287 355 
<< pdiffusion >>
rect 287 354 288 355 
<< m1 >>
rect 289 354 290 355 
<< m1 >>
rect 291 354 292 355 
<< m1 >>
rect 293 354 294 355 
<< pdiffusion >>
rect 300 354 301 355 
<< pdiffusion >>
rect 301 354 302 355 
<< pdiffusion >>
rect 302 354 303 355 
<< pdiffusion >>
rect 303 354 304 355 
<< pdiffusion >>
rect 304 354 305 355 
<< pdiffusion >>
rect 305 354 306 355 
<< pdiffusion >>
rect 318 354 319 355 
<< pdiffusion >>
rect 319 354 320 355 
<< pdiffusion >>
rect 320 354 321 355 
<< pdiffusion >>
rect 321 354 322 355 
<< pdiffusion >>
rect 322 354 323 355 
<< pdiffusion >>
rect 323 354 324 355 
<< m1 >>
rect 325 354 326 355 
<< pdiffusion >>
rect 336 354 337 355 
<< pdiffusion >>
rect 337 354 338 355 
<< pdiffusion >>
rect 338 354 339 355 
<< pdiffusion >>
rect 339 354 340 355 
<< pdiffusion >>
rect 340 354 341 355 
<< pdiffusion >>
rect 341 354 342 355 
<< pdiffusion >>
rect 354 354 355 355 
<< pdiffusion >>
rect 355 354 356 355 
<< pdiffusion >>
rect 356 354 357 355 
<< pdiffusion >>
rect 357 354 358 355 
<< pdiffusion >>
rect 358 354 359 355 
<< pdiffusion >>
rect 359 354 360 355 
<< pdiffusion >>
rect 372 354 373 355 
<< pdiffusion >>
rect 373 354 374 355 
<< pdiffusion >>
rect 374 354 375 355 
<< pdiffusion >>
rect 375 354 376 355 
<< pdiffusion >>
rect 376 354 377 355 
<< pdiffusion >>
rect 377 354 378 355 
<< m1 >>
rect 379 354 380 355 
<< pdiffusion >>
rect 390 354 391 355 
<< pdiffusion >>
rect 391 354 392 355 
<< pdiffusion >>
rect 392 354 393 355 
<< pdiffusion >>
rect 393 354 394 355 
<< pdiffusion >>
rect 394 354 395 355 
<< pdiffusion >>
rect 395 354 396 355 
<< pdiffusion >>
rect 408 354 409 355 
<< pdiffusion >>
rect 409 354 410 355 
<< pdiffusion >>
rect 410 354 411 355 
<< pdiffusion >>
rect 411 354 412 355 
<< pdiffusion >>
rect 412 354 413 355 
<< pdiffusion >>
rect 413 354 414 355 
<< pdiffusion >>
rect 444 354 445 355 
<< pdiffusion >>
rect 445 354 446 355 
<< pdiffusion >>
rect 446 354 447 355 
<< pdiffusion >>
rect 447 354 448 355 
<< pdiffusion >>
rect 448 354 449 355 
<< pdiffusion >>
rect 449 354 450 355 
<< pdiffusion >>
rect 12 355 13 356 
<< pdiffusion >>
rect 13 355 14 356 
<< pdiffusion >>
rect 14 355 15 356 
<< pdiffusion >>
rect 15 355 16 356 
<< pdiffusion >>
rect 16 355 17 356 
<< pdiffusion >>
rect 17 355 18 356 
<< pdiffusion >>
rect 30 355 31 356 
<< pdiffusion >>
rect 31 355 32 356 
<< pdiffusion >>
rect 32 355 33 356 
<< pdiffusion >>
rect 33 355 34 356 
<< pdiffusion >>
rect 34 355 35 356 
<< pdiffusion >>
rect 35 355 36 356 
<< m1 >>
rect 37 355 38 356 
<< pdiffusion >>
rect 48 355 49 356 
<< pdiffusion >>
rect 49 355 50 356 
<< pdiffusion >>
rect 50 355 51 356 
<< pdiffusion >>
rect 51 355 52 356 
<< pdiffusion >>
rect 52 355 53 356 
<< pdiffusion >>
rect 53 355 54 356 
<< pdiffusion >>
rect 66 355 67 356 
<< pdiffusion >>
rect 67 355 68 356 
<< pdiffusion >>
rect 68 355 69 356 
<< pdiffusion >>
rect 69 355 70 356 
<< pdiffusion >>
rect 70 355 71 356 
<< pdiffusion >>
rect 71 355 72 356 
<< pdiffusion >>
rect 84 355 85 356 
<< pdiffusion >>
rect 85 355 86 356 
<< pdiffusion >>
rect 86 355 87 356 
<< pdiffusion >>
rect 87 355 88 356 
<< pdiffusion >>
rect 88 355 89 356 
<< pdiffusion >>
rect 89 355 90 356 
<< m1 >>
rect 91 355 92 356 
<< pdiffusion >>
rect 102 355 103 356 
<< pdiffusion >>
rect 103 355 104 356 
<< pdiffusion >>
rect 104 355 105 356 
<< pdiffusion >>
rect 105 355 106 356 
<< pdiffusion >>
rect 106 355 107 356 
<< pdiffusion >>
rect 107 355 108 356 
<< pdiffusion >>
rect 120 355 121 356 
<< pdiffusion >>
rect 121 355 122 356 
<< pdiffusion >>
rect 122 355 123 356 
<< pdiffusion >>
rect 123 355 124 356 
<< pdiffusion >>
rect 124 355 125 356 
<< pdiffusion >>
rect 125 355 126 356 
<< m1 >>
rect 127 355 128 356 
<< m2 >>
rect 127 355 128 356 
<< pdiffusion >>
rect 138 355 139 356 
<< pdiffusion >>
rect 139 355 140 356 
<< pdiffusion >>
rect 140 355 141 356 
<< pdiffusion >>
rect 141 355 142 356 
<< pdiffusion >>
rect 142 355 143 356 
<< pdiffusion >>
rect 143 355 144 356 
<< pdiffusion >>
rect 156 355 157 356 
<< pdiffusion >>
rect 157 355 158 356 
<< pdiffusion >>
rect 158 355 159 356 
<< pdiffusion >>
rect 159 355 160 356 
<< pdiffusion >>
rect 160 355 161 356 
<< pdiffusion >>
rect 161 355 162 356 
<< m1 >>
rect 172 355 173 356 
<< pdiffusion >>
rect 174 355 175 356 
<< pdiffusion >>
rect 175 355 176 356 
<< pdiffusion >>
rect 176 355 177 356 
<< pdiffusion >>
rect 177 355 178 356 
<< pdiffusion >>
rect 178 355 179 356 
<< pdiffusion >>
rect 179 355 180 356 
<< pdiffusion >>
rect 192 355 193 356 
<< pdiffusion >>
rect 193 355 194 356 
<< pdiffusion >>
rect 194 355 195 356 
<< pdiffusion >>
rect 195 355 196 356 
<< pdiffusion >>
rect 196 355 197 356 
<< pdiffusion >>
rect 197 355 198 356 
<< pdiffusion >>
rect 210 355 211 356 
<< pdiffusion >>
rect 211 355 212 356 
<< pdiffusion >>
rect 212 355 213 356 
<< pdiffusion >>
rect 213 355 214 356 
<< pdiffusion >>
rect 214 355 215 356 
<< pdiffusion >>
rect 215 355 216 356 
<< m1 >>
rect 217 355 218 356 
<< pdiffusion >>
rect 228 355 229 356 
<< pdiffusion >>
rect 229 355 230 356 
<< pdiffusion >>
rect 230 355 231 356 
<< pdiffusion >>
rect 231 355 232 356 
<< pdiffusion >>
rect 232 355 233 356 
<< pdiffusion >>
rect 233 355 234 356 
<< m1 >>
rect 244 355 245 356 
<< pdiffusion >>
rect 246 355 247 356 
<< pdiffusion >>
rect 247 355 248 356 
<< pdiffusion >>
rect 248 355 249 356 
<< pdiffusion >>
rect 249 355 250 356 
<< pdiffusion >>
rect 250 355 251 356 
<< pdiffusion >>
rect 251 355 252 356 
<< m1 >>
rect 253 355 254 356 
<< m2 >>
rect 254 355 255 356 
<< pdiffusion >>
rect 264 355 265 356 
<< pdiffusion >>
rect 265 355 266 356 
<< pdiffusion >>
rect 266 355 267 356 
<< pdiffusion >>
rect 267 355 268 356 
<< pdiffusion >>
rect 268 355 269 356 
<< pdiffusion >>
rect 269 355 270 356 
<< pdiffusion >>
rect 282 355 283 356 
<< pdiffusion >>
rect 283 355 284 356 
<< pdiffusion >>
rect 284 355 285 356 
<< pdiffusion >>
rect 285 355 286 356 
<< pdiffusion >>
rect 286 355 287 356 
<< pdiffusion >>
rect 287 355 288 356 
<< m1 >>
rect 289 355 290 356 
<< m1 >>
rect 291 355 292 356 
<< m1 >>
rect 293 355 294 356 
<< pdiffusion >>
rect 300 355 301 356 
<< pdiffusion >>
rect 301 355 302 356 
<< pdiffusion >>
rect 302 355 303 356 
<< pdiffusion >>
rect 303 355 304 356 
<< pdiffusion >>
rect 304 355 305 356 
<< pdiffusion >>
rect 305 355 306 356 
<< pdiffusion >>
rect 318 355 319 356 
<< pdiffusion >>
rect 319 355 320 356 
<< pdiffusion >>
rect 320 355 321 356 
<< pdiffusion >>
rect 321 355 322 356 
<< pdiffusion >>
rect 322 355 323 356 
<< pdiffusion >>
rect 323 355 324 356 
<< m1 >>
rect 325 355 326 356 
<< pdiffusion >>
rect 336 355 337 356 
<< pdiffusion >>
rect 337 355 338 356 
<< pdiffusion >>
rect 338 355 339 356 
<< pdiffusion >>
rect 339 355 340 356 
<< pdiffusion >>
rect 340 355 341 356 
<< pdiffusion >>
rect 341 355 342 356 
<< pdiffusion >>
rect 354 355 355 356 
<< pdiffusion >>
rect 355 355 356 356 
<< pdiffusion >>
rect 356 355 357 356 
<< pdiffusion >>
rect 357 355 358 356 
<< pdiffusion >>
rect 358 355 359 356 
<< pdiffusion >>
rect 359 355 360 356 
<< pdiffusion >>
rect 372 355 373 356 
<< pdiffusion >>
rect 373 355 374 356 
<< pdiffusion >>
rect 374 355 375 356 
<< pdiffusion >>
rect 375 355 376 356 
<< pdiffusion >>
rect 376 355 377 356 
<< pdiffusion >>
rect 377 355 378 356 
<< m1 >>
rect 379 355 380 356 
<< pdiffusion >>
rect 390 355 391 356 
<< pdiffusion >>
rect 391 355 392 356 
<< pdiffusion >>
rect 392 355 393 356 
<< pdiffusion >>
rect 393 355 394 356 
<< pdiffusion >>
rect 394 355 395 356 
<< pdiffusion >>
rect 395 355 396 356 
<< pdiffusion >>
rect 408 355 409 356 
<< pdiffusion >>
rect 409 355 410 356 
<< pdiffusion >>
rect 410 355 411 356 
<< pdiffusion >>
rect 411 355 412 356 
<< pdiffusion >>
rect 412 355 413 356 
<< pdiffusion >>
rect 413 355 414 356 
<< pdiffusion >>
rect 444 355 445 356 
<< pdiffusion >>
rect 445 355 446 356 
<< pdiffusion >>
rect 446 355 447 356 
<< pdiffusion >>
rect 447 355 448 356 
<< pdiffusion >>
rect 448 355 449 356 
<< pdiffusion >>
rect 449 355 450 356 
<< pdiffusion >>
rect 12 356 13 357 
<< pdiffusion >>
rect 13 356 14 357 
<< pdiffusion >>
rect 14 356 15 357 
<< pdiffusion >>
rect 15 356 16 357 
<< pdiffusion >>
rect 16 356 17 357 
<< pdiffusion >>
rect 17 356 18 357 
<< pdiffusion >>
rect 30 356 31 357 
<< pdiffusion >>
rect 31 356 32 357 
<< pdiffusion >>
rect 32 356 33 357 
<< pdiffusion >>
rect 33 356 34 357 
<< pdiffusion >>
rect 34 356 35 357 
<< pdiffusion >>
rect 35 356 36 357 
<< m1 >>
rect 37 356 38 357 
<< pdiffusion >>
rect 48 356 49 357 
<< pdiffusion >>
rect 49 356 50 357 
<< pdiffusion >>
rect 50 356 51 357 
<< pdiffusion >>
rect 51 356 52 357 
<< pdiffusion >>
rect 52 356 53 357 
<< pdiffusion >>
rect 53 356 54 357 
<< pdiffusion >>
rect 66 356 67 357 
<< pdiffusion >>
rect 67 356 68 357 
<< pdiffusion >>
rect 68 356 69 357 
<< pdiffusion >>
rect 69 356 70 357 
<< pdiffusion >>
rect 70 356 71 357 
<< pdiffusion >>
rect 71 356 72 357 
<< pdiffusion >>
rect 84 356 85 357 
<< pdiffusion >>
rect 85 356 86 357 
<< pdiffusion >>
rect 86 356 87 357 
<< pdiffusion >>
rect 87 356 88 357 
<< pdiffusion >>
rect 88 356 89 357 
<< pdiffusion >>
rect 89 356 90 357 
<< m1 >>
rect 91 356 92 357 
<< pdiffusion >>
rect 102 356 103 357 
<< pdiffusion >>
rect 103 356 104 357 
<< pdiffusion >>
rect 104 356 105 357 
<< pdiffusion >>
rect 105 356 106 357 
<< pdiffusion >>
rect 106 356 107 357 
<< pdiffusion >>
rect 107 356 108 357 
<< pdiffusion >>
rect 120 356 121 357 
<< pdiffusion >>
rect 121 356 122 357 
<< pdiffusion >>
rect 122 356 123 357 
<< pdiffusion >>
rect 123 356 124 357 
<< pdiffusion >>
rect 124 356 125 357 
<< pdiffusion >>
rect 125 356 126 357 
<< m1 >>
rect 127 356 128 357 
<< m2 >>
rect 127 356 128 357 
<< pdiffusion >>
rect 138 356 139 357 
<< pdiffusion >>
rect 139 356 140 357 
<< pdiffusion >>
rect 140 356 141 357 
<< pdiffusion >>
rect 141 356 142 357 
<< pdiffusion >>
rect 142 356 143 357 
<< pdiffusion >>
rect 143 356 144 357 
<< pdiffusion >>
rect 156 356 157 357 
<< pdiffusion >>
rect 157 356 158 357 
<< pdiffusion >>
rect 158 356 159 357 
<< pdiffusion >>
rect 159 356 160 357 
<< pdiffusion >>
rect 160 356 161 357 
<< pdiffusion >>
rect 161 356 162 357 
<< m1 >>
rect 172 356 173 357 
<< pdiffusion >>
rect 174 356 175 357 
<< pdiffusion >>
rect 175 356 176 357 
<< pdiffusion >>
rect 176 356 177 357 
<< pdiffusion >>
rect 177 356 178 357 
<< pdiffusion >>
rect 178 356 179 357 
<< pdiffusion >>
rect 179 356 180 357 
<< pdiffusion >>
rect 192 356 193 357 
<< pdiffusion >>
rect 193 356 194 357 
<< pdiffusion >>
rect 194 356 195 357 
<< pdiffusion >>
rect 195 356 196 357 
<< pdiffusion >>
rect 196 356 197 357 
<< pdiffusion >>
rect 197 356 198 357 
<< pdiffusion >>
rect 210 356 211 357 
<< pdiffusion >>
rect 211 356 212 357 
<< pdiffusion >>
rect 212 356 213 357 
<< pdiffusion >>
rect 213 356 214 357 
<< pdiffusion >>
rect 214 356 215 357 
<< pdiffusion >>
rect 215 356 216 357 
<< m1 >>
rect 217 356 218 357 
<< pdiffusion >>
rect 228 356 229 357 
<< pdiffusion >>
rect 229 356 230 357 
<< pdiffusion >>
rect 230 356 231 357 
<< pdiffusion >>
rect 231 356 232 357 
<< pdiffusion >>
rect 232 356 233 357 
<< pdiffusion >>
rect 233 356 234 357 
<< m1 >>
rect 244 356 245 357 
<< pdiffusion >>
rect 246 356 247 357 
<< pdiffusion >>
rect 247 356 248 357 
<< pdiffusion >>
rect 248 356 249 357 
<< pdiffusion >>
rect 249 356 250 357 
<< pdiffusion >>
rect 250 356 251 357 
<< pdiffusion >>
rect 251 356 252 357 
<< m1 >>
rect 253 356 254 357 
<< m2 >>
rect 254 356 255 357 
<< pdiffusion >>
rect 264 356 265 357 
<< pdiffusion >>
rect 265 356 266 357 
<< pdiffusion >>
rect 266 356 267 357 
<< pdiffusion >>
rect 267 356 268 357 
<< pdiffusion >>
rect 268 356 269 357 
<< pdiffusion >>
rect 269 356 270 357 
<< pdiffusion >>
rect 282 356 283 357 
<< pdiffusion >>
rect 283 356 284 357 
<< pdiffusion >>
rect 284 356 285 357 
<< pdiffusion >>
rect 285 356 286 357 
<< pdiffusion >>
rect 286 356 287 357 
<< pdiffusion >>
rect 287 356 288 357 
<< m1 >>
rect 289 356 290 357 
<< m1 >>
rect 291 356 292 357 
<< m1 >>
rect 293 356 294 357 
<< pdiffusion >>
rect 300 356 301 357 
<< pdiffusion >>
rect 301 356 302 357 
<< pdiffusion >>
rect 302 356 303 357 
<< pdiffusion >>
rect 303 356 304 357 
<< pdiffusion >>
rect 304 356 305 357 
<< pdiffusion >>
rect 305 356 306 357 
<< pdiffusion >>
rect 318 356 319 357 
<< pdiffusion >>
rect 319 356 320 357 
<< pdiffusion >>
rect 320 356 321 357 
<< pdiffusion >>
rect 321 356 322 357 
<< pdiffusion >>
rect 322 356 323 357 
<< pdiffusion >>
rect 323 356 324 357 
<< m1 >>
rect 325 356 326 357 
<< pdiffusion >>
rect 336 356 337 357 
<< pdiffusion >>
rect 337 356 338 357 
<< pdiffusion >>
rect 338 356 339 357 
<< pdiffusion >>
rect 339 356 340 357 
<< pdiffusion >>
rect 340 356 341 357 
<< pdiffusion >>
rect 341 356 342 357 
<< pdiffusion >>
rect 354 356 355 357 
<< pdiffusion >>
rect 355 356 356 357 
<< pdiffusion >>
rect 356 356 357 357 
<< pdiffusion >>
rect 357 356 358 357 
<< pdiffusion >>
rect 358 356 359 357 
<< pdiffusion >>
rect 359 356 360 357 
<< pdiffusion >>
rect 372 356 373 357 
<< pdiffusion >>
rect 373 356 374 357 
<< pdiffusion >>
rect 374 356 375 357 
<< pdiffusion >>
rect 375 356 376 357 
<< pdiffusion >>
rect 376 356 377 357 
<< pdiffusion >>
rect 377 356 378 357 
<< m1 >>
rect 379 356 380 357 
<< pdiffusion >>
rect 390 356 391 357 
<< pdiffusion >>
rect 391 356 392 357 
<< pdiffusion >>
rect 392 356 393 357 
<< pdiffusion >>
rect 393 356 394 357 
<< pdiffusion >>
rect 394 356 395 357 
<< pdiffusion >>
rect 395 356 396 357 
<< pdiffusion >>
rect 408 356 409 357 
<< pdiffusion >>
rect 409 356 410 357 
<< pdiffusion >>
rect 410 356 411 357 
<< pdiffusion >>
rect 411 356 412 357 
<< pdiffusion >>
rect 412 356 413 357 
<< pdiffusion >>
rect 413 356 414 357 
<< pdiffusion >>
rect 444 356 445 357 
<< pdiffusion >>
rect 445 356 446 357 
<< pdiffusion >>
rect 446 356 447 357 
<< pdiffusion >>
rect 447 356 448 357 
<< pdiffusion >>
rect 448 356 449 357 
<< pdiffusion >>
rect 449 356 450 357 
<< pdiffusion >>
rect 12 357 13 358 
<< pdiffusion >>
rect 13 357 14 358 
<< pdiffusion >>
rect 14 357 15 358 
<< pdiffusion >>
rect 15 357 16 358 
<< pdiffusion >>
rect 16 357 17 358 
<< pdiffusion >>
rect 17 357 18 358 
<< pdiffusion >>
rect 30 357 31 358 
<< pdiffusion >>
rect 31 357 32 358 
<< pdiffusion >>
rect 32 357 33 358 
<< pdiffusion >>
rect 33 357 34 358 
<< pdiffusion >>
rect 34 357 35 358 
<< pdiffusion >>
rect 35 357 36 358 
<< m1 >>
rect 37 357 38 358 
<< pdiffusion >>
rect 48 357 49 358 
<< pdiffusion >>
rect 49 357 50 358 
<< pdiffusion >>
rect 50 357 51 358 
<< pdiffusion >>
rect 51 357 52 358 
<< pdiffusion >>
rect 52 357 53 358 
<< pdiffusion >>
rect 53 357 54 358 
<< pdiffusion >>
rect 66 357 67 358 
<< pdiffusion >>
rect 67 357 68 358 
<< pdiffusion >>
rect 68 357 69 358 
<< pdiffusion >>
rect 69 357 70 358 
<< pdiffusion >>
rect 70 357 71 358 
<< pdiffusion >>
rect 71 357 72 358 
<< pdiffusion >>
rect 84 357 85 358 
<< pdiffusion >>
rect 85 357 86 358 
<< pdiffusion >>
rect 86 357 87 358 
<< pdiffusion >>
rect 87 357 88 358 
<< pdiffusion >>
rect 88 357 89 358 
<< pdiffusion >>
rect 89 357 90 358 
<< m1 >>
rect 91 357 92 358 
<< pdiffusion >>
rect 102 357 103 358 
<< pdiffusion >>
rect 103 357 104 358 
<< pdiffusion >>
rect 104 357 105 358 
<< pdiffusion >>
rect 105 357 106 358 
<< pdiffusion >>
rect 106 357 107 358 
<< pdiffusion >>
rect 107 357 108 358 
<< pdiffusion >>
rect 120 357 121 358 
<< pdiffusion >>
rect 121 357 122 358 
<< pdiffusion >>
rect 122 357 123 358 
<< pdiffusion >>
rect 123 357 124 358 
<< pdiffusion >>
rect 124 357 125 358 
<< pdiffusion >>
rect 125 357 126 358 
<< m1 >>
rect 127 357 128 358 
<< m2 >>
rect 127 357 128 358 
<< pdiffusion >>
rect 138 357 139 358 
<< pdiffusion >>
rect 139 357 140 358 
<< pdiffusion >>
rect 140 357 141 358 
<< pdiffusion >>
rect 141 357 142 358 
<< pdiffusion >>
rect 142 357 143 358 
<< pdiffusion >>
rect 143 357 144 358 
<< pdiffusion >>
rect 156 357 157 358 
<< pdiffusion >>
rect 157 357 158 358 
<< pdiffusion >>
rect 158 357 159 358 
<< pdiffusion >>
rect 159 357 160 358 
<< pdiffusion >>
rect 160 357 161 358 
<< pdiffusion >>
rect 161 357 162 358 
<< m1 >>
rect 172 357 173 358 
<< pdiffusion >>
rect 174 357 175 358 
<< pdiffusion >>
rect 175 357 176 358 
<< pdiffusion >>
rect 176 357 177 358 
<< pdiffusion >>
rect 177 357 178 358 
<< pdiffusion >>
rect 178 357 179 358 
<< pdiffusion >>
rect 179 357 180 358 
<< pdiffusion >>
rect 192 357 193 358 
<< pdiffusion >>
rect 193 357 194 358 
<< pdiffusion >>
rect 194 357 195 358 
<< pdiffusion >>
rect 195 357 196 358 
<< pdiffusion >>
rect 196 357 197 358 
<< pdiffusion >>
rect 197 357 198 358 
<< pdiffusion >>
rect 210 357 211 358 
<< pdiffusion >>
rect 211 357 212 358 
<< pdiffusion >>
rect 212 357 213 358 
<< pdiffusion >>
rect 213 357 214 358 
<< pdiffusion >>
rect 214 357 215 358 
<< pdiffusion >>
rect 215 357 216 358 
<< m1 >>
rect 217 357 218 358 
<< pdiffusion >>
rect 228 357 229 358 
<< pdiffusion >>
rect 229 357 230 358 
<< pdiffusion >>
rect 230 357 231 358 
<< pdiffusion >>
rect 231 357 232 358 
<< pdiffusion >>
rect 232 357 233 358 
<< pdiffusion >>
rect 233 357 234 358 
<< m1 >>
rect 244 357 245 358 
<< pdiffusion >>
rect 246 357 247 358 
<< pdiffusion >>
rect 247 357 248 358 
<< pdiffusion >>
rect 248 357 249 358 
<< pdiffusion >>
rect 249 357 250 358 
<< pdiffusion >>
rect 250 357 251 358 
<< pdiffusion >>
rect 251 357 252 358 
<< m1 >>
rect 253 357 254 358 
<< m2 >>
rect 254 357 255 358 
<< pdiffusion >>
rect 264 357 265 358 
<< pdiffusion >>
rect 265 357 266 358 
<< pdiffusion >>
rect 266 357 267 358 
<< pdiffusion >>
rect 267 357 268 358 
<< pdiffusion >>
rect 268 357 269 358 
<< pdiffusion >>
rect 269 357 270 358 
<< pdiffusion >>
rect 282 357 283 358 
<< pdiffusion >>
rect 283 357 284 358 
<< pdiffusion >>
rect 284 357 285 358 
<< pdiffusion >>
rect 285 357 286 358 
<< pdiffusion >>
rect 286 357 287 358 
<< pdiffusion >>
rect 287 357 288 358 
<< m1 >>
rect 289 357 290 358 
<< m1 >>
rect 291 357 292 358 
<< m1 >>
rect 293 357 294 358 
<< pdiffusion >>
rect 300 357 301 358 
<< pdiffusion >>
rect 301 357 302 358 
<< pdiffusion >>
rect 302 357 303 358 
<< pdiffusion >>
rect 303 357 304 358 
<< pdiffusion >>
rect 304 357 305 358 
<< pdiffusion >>
rect 305 357 306 358 
<< pdiffusion >>
rect 318 357 319 358 
<< pdiffusion >>
rect 319 357 320 358 
<< pdiffusion >>
rect 320 357 321 358 
<< pdiffusion >>
rect 321 357 322 358 
<< pdiffusion >>
rect 322 357 323 358 
<< pdiffusion >>
rect 323 357 324 358 
<< m1 >>
rect 325 357 326 358 
<< pdiffusion >>
rect 336 357 337 358 
<< pdiffusion >>
rect 337 357 338 358 
<< pdiffusion >>
rect 338 357 339 358 
<< pdiffusion >>
rect 339 357 340 358 
<< pdiffusion >>
rect 340 357 341 358 
<< pdiffusion >>
rect 341 357 342 358 
<< pdiffusion >>
rect 354 357 355 358 
<< pdiffusion >>
rect 355 357 356 358 
<< pdiffusion >>
rect 356 357 357 358 
<< pdiffusion >>
rect 357 357 358 358 
<< pdiffusion >>
rect 358 357 359 358 
<< pdiffusion >>
rect 359 357 360 358 
<< pdiffusion >>
rect 372 357 373 358 
<< pdiffusion >>
rect 373 357 374 358 
<< pdiffusion >>
rect 374 357 375 358 
<< pdiffusion >>
rect 375 357 376 358 
<< pdiffusion >>
rect 376 357 377 358 
<< pdiffusion >>
rect 377 357 378 358 
<< m1 >>
rect 379 357 380 358 
<< pdiffusion >>
rect 390 357 391 358 
<< pdiffusion >>
rect 391 357 392 358 
<< pdiffusion >>
rect 392 357 393 358 
<< pdiffusion >>
rect 393 357 394 358 
<< pdiffusion >>
rect 394 357 395 358 
<< pdiffusion >>
rect 395 357 396 358 
<< pdiffusion >>
rect 408 357 409 358 
<< pdiffusion >>
rect 409 357 410 358 
<< pdiffusion >>
rect 410 357 411 358 
<< pdiffusion >>
rect 411 357 412 358 
<< pdiffusion >>
rect 412 357 413 358 
<< pdiffusion >>
rect 413 357 414 358 
<< pdiffusion >>
rect 444 357 445 358 
<< pdiffusion >>
rect 445 357 446 358 
<< pdiffusion >>
rect 446 357 447 358 
<< pdiffusion >>
rect 447 357 448 358 
<< pdiffusion >>
rect 448 357 449 358 
<< pdiffusion >>
rect 449 357 450 358 
<< pdiffusion >>
rect 12 358 13 359 
<< pdiffusion >>
rect 13 358 14 359 
<< pdiffusion >>
rect 14 358 15 359 
<< pdiffusion >>
rect 15 358 16 359 
<< pdiffusion >>
rect 16 358 17 359 
<< pdiffusion >>
rect 17 358 18 359 
<< pdiffusion >>
rect 30 358 31 359 
<< pdiffusion >>
rect 31 358 32 359 
<< pdiffusion >>
rect 32 358 33 359 
<< pdiffusion >>
rect 33 358 34 359 
<< pdiffusion >>
rect 34 358 35 359 
<< pdiffusion >>
rect 35 358 36 359 
<< m1 >>
rect 37 358 38 359 
<< pdiffusion >>
rect 48 358 49 359 
<< pdiffusion >>
rect 49 358 50 359 
<< pdiffusion >>
rect 50 358 51 359 
<< pdiffusion >>
rect 51 358 52 359 
<< pdiffusion >>
rect 52 358 53 359 
<< pdiffusion >>
rect 53 358 54 359 
<< pdiffusion >>
rect 66 358 67 359 
<< pdiffusion >>
rect 67 358 68 359 
<< pdiffusion >>
rect 68 358 69 359 
<< pdiffusion >>
rect 69 358 70 359 
<< pdiffusion >>
rect 70 358 71 359 
<< pdiffusion >>
rect 71 358 72 359 
<< pdiffusion >>
rect 84 358 85 359 
<< pdiffusion >>
rect 85 358 86 359 
<< pdiffusion >>
rect 86 358 87 359 
<< pdiffusion >>
rect 87 358 88 359 
<< pdiffusion >>
rect 88 358 89 359 
<< pdiffusion >>
rect 89 358 90 359 
<< m1 >>
rect 91 358 92 359 
<< pdiffusion >>
rect 102 358 103 359 
<< pdiffusion >>
rect 103 358 104 359 
<< pdiffusion >>
rect 104 358 105 359 
<< pdiffusion >>
rect 105 358 106 359 
<< pdiffusion >>
rect 106 358 107 359 
<< pdiffusion >>
rect 107 358 108 359 
<< pdiffusion >>
rect 120 358 121 359 
<< pdiffusion >>
rect 121 358 122 359 
<< pdiffusion >>
rect 122 358 123 359 
<< pdiffusion >>
rect 123 358 124 359 
<< pdiffusion >>
rect 124 358 125 359 
<< pdiffusion >>
rect 125 358 126 359 
<< m1 >>
rect 127 358 128 359 
<< m2 >>
rect 127 358 128 359 
<< pdiffusion >>
rect 138 358 139 359 
<< pdiffusion >>
rect 139 358 140 359 
<< pdiffusion >>
rect 140 358 141 359 
<< pdiffusion >>
rect 141 358 142 359 
<< pdiffusion >>
rect 142 358 143 359 
<< pdiffusion >>
rect 143 358 144 359 
<< pdiffusion >>
rect 156 358 157 359 
<< pdiffusion >>
rect 157 358 158 359 
<< pdiffusion >>
rect 158 358 159 359 
<< pdiffusion >>
rect 159 358 160 359 
<< pdiffusion >>
rect 160 358 161 359 
<< pdiffusion >>
rect 161 358 162 359 
<< m1 >>
rect 172 358 173 359 
<< pdiffusion >>
rect 174 358 175 359 
<< pdiffusion >>
rect 175 358 176 359 
<< pdiffusion >>
rect 176 358 177 359 
<< pdiffusion >>
rect 177 358 178 359 
<< pdiffusion >>
rect 178 358 179 359 
<< pdiffusion >>
rect 179 358 180 359 
<< pdiffusion >>
rect 192 358 193 359 
<< pdiffusion >>
rect 193 358 194 359 
<< pdiffusion >>
rect 194 358 195 359 
<< pdiffusion >>
rect 195 358 196 359 
<< pdiffusion >>
rect 196 358 197 359 
<< pdiffusion >>
rect 197 358 198 359 
<< pdiffusion >>
rect 210 358 211 359 
<< pdiffusion >>
rect 211 358 212 359 
<< pdiffusion >>
rect 212 358 213 359 
<< pdiffusion >>
rect 213 358 214 359 
<< pdiffusion >>
rect 214 358 215 359 
<< pdiffusion >>
rect 215 358 216 359 
<< m1 >>
rect 217 358 218 359 
<< pdiffusion >>
rect 228 358 229 359 
<< pdiffusion >>
rect 229 358 230 359 
<< pdiffusion >>
rect 230 358 231 359 
<< pdiffusion >>
rect 231 358 232 359 
<< pdiffusion >>
rect 232 358 233 359 
<< pdiffusion >>
rect 233 358 234 359 
<< m1 >>
rect 244 358 245 359 
<< pdiffusion >>
rect 246 358 247 359 
<< pdiffusion >>
rect 247 358 248 359 
<< pdiffusion >>
rect 248 358 249 359 
<< pdiffusion >>
rect 249 358 250 359 
<< pdiffusion >>
rect 250 358 251 359 
<< pdiffusion >>
rect 251 358 252 359 
<< m1 >>
rect 253 358 254 359 
<< m2 >>
rect 254 358 255 359 
<< pdiffusion >>
rect 264 358 265 359 
<< pdiffusion >>
rect 265 358 266 359 
<< pdiffusion >>
rect 266 358 267 359 
<< pdiffusion >>
rect 267 358 268 359 
<< pdiffusion >>
rect 268 358 269 359 
<< pdiffusion >>
rect 269 358 270 359 
<< pdiffusion >>
rect 282 358 283 359 
<< pdiffusion >>
rect 283 358 284 359 
<< pdiffusion >>
rect 284 358 285 359 
<< pdiffusion >>
rect 285 358 286 359 
<< pdiffusion >>
rect 286 358 287 359 
<< pdiffusion >>
rect 287 358 288 359 
<< m1 >>
rect 289 358 290 359 
<< m1 >>
rect 291 358 292 359 
<< m1 >>
rect 293 358 294 359 
<< pdiffusion >>
rect 300 358 301 359 
<< pdiffusion >>
rect 301 358 302 359 
<< pdiffusion >>
rect 302 358 303 359 
<< pdiffusion >>
rect 303 358 304 359 
<< pdiffusion >>
rect 304 358 305 359 
<< pdiffusion >>
rect 305 358 306 359 
<< pdiffusion >>
rect 318 358 319 359 
<< pdiffusion >>
rect 319 358 320 359 
<< pdiffusion >>
rect 320 358 321 359 
<< pdiffusion >>
rect 321 358 322 359 
<< pdiffusion >>
rect 322 358 323 359 
<< pdiffusion >>
rect 323 358 324 359 
<< m1 >>
rect 325 358 326 359 
<< pdiffusion >>
rect 336 358 337 359 
<< pdiffusion >>
rect 337 358 338 359 
<< pdiffusion >>
rect 338 358 339 359 
<< pdiffusion >>
rect 339 358 340 359 
<< pdiffusion >>
rect 340 358 341 359 
<< pdiffusion >>
rect 341 358 342 359 
<< pdiffusion >>
rect 354 358 355 359 
<< pdiffusion >>
rect 355 358 356 359 
<< pdiffusion >>
rect 356 358 357 359 
<< pdiffusion >>
rect 357 358 358 359 
<< pdiffusion >>
rect 358 358 359 359 
<< pdiffusion >>
rect 359 358 360 359 
<< pdiffusion >>
rect 372 358 373 359 
<< pdiffusion >>
rect 373 358 374 359 
<< pdiffusion >>
rect 374 358 375 359 
<< pdiffusion >>
rect 375 358 376 359 
<< pdiffusion >>
rect 376 358 377 359 
<< pdiffusion >>
rect 377 358 378 359 
<< m1 >>
rect 379 358 380 359 
<< pdiffusion >>
rect 390 358 391 359 
<< pdiffusion >>
rect 391 358 392 359 
<< pdiffusion >>
rect 392 358 393 359 
<< pdiffusion >>
rect 393 358 394 359 
<< pdiffusion >>
rect 394 358 395 359 
<< pdiffusion >>
rect 395 358 396 359 
<< pdiffusion >>
rect 408 358 409 359 
<< pdiffusion >>
rect 409 358 410 359 
<< pdiffusion >>
rect 410 358 411 359 
<< pdiffusion >>
rect 411 358 412 359 
<< pdiffusion >>
rect 412 358 413 359 
<< pdiffusion >>
rect 413 358 414 359 
<< pdiffusion >>
rect 444 358 445 359 
<< pdiffusion >>
rect 445 358 446 359 
<< pdiffusion >>
rect 446 358 447 359 
<< pdiffusion >>
rect 447 358 448 359 
<< pdiffusion >>
rect 448 358 449 359 
<< pdiffusion >>
rect 449 358 450 359 
<< pdiffusion >>
rect 12 359 13 360 
<< pdiffusion >>
rect 13 359 14 360 
<< pdiffusion >>
rect 14 359 15 360 
<< pdiffusion >>
rect 15 359 16 360 
<< pdiffusion >>
rect 16 359 17 360 
<< pdiffusion >>
rect 17 359 18 360 
<< pdiffusion >>
rect 30 359 31 360 
<< pdiffusion >>
rect 31 359 32 360 
<< pdiffusion >>
rect 32 359 33 360 
<< pdiffusion >>
rect 33 359 34 360 
<< pdiffusion >>
rect 34 359 35 360 
<< pdiffusion >>
rect 35 359 36 360 
<< m1 >>
rect 37 359 38 360 
<< pdiffusion >>
rect 48 359 49 360 
<< pdiffusion >>
rect 49 359 50 360 
<< pdiffusion >>
rect 50 359 51 360 
<< pdiffusion >>
rect 51 359 52 360 
<< pdiffusion >>
rect 52 359 53 360 
<< pdiffusion >>
rect 53 359 54 360 
<< pdiffusion >>
rect 66 359 67 360 
<< pdiffusion >>
rect 67 359 68 360 
<< pdiffusion >>
rect 68 359 69 360 
<< pdiffusion >>
rect 69 359 70 360 
<< pdiffusion >>
rect 70 359 71 360 
<< pdiffusion >>
rect 71 359 72 360 
<< pdiffusion >>
rect 84 359 85 360 
<< pdiffusion >>
rect 85 359 86 360 
<< pdiffusion >>
rect 86 359 87 360 
<< pdiffusion >>
rect 87 359 88 360 
<< m1 >>
rect 88 359 89 360 
<< pdiffusion >>
rect 88 359 89 360 
<< pdiffusion >>
rect 89 359 90 360 
<< m1 >>
rect 91 359 92 360 
<< pdiffusion >>
rect 102 359 103 360 
<< pdiffusion >>
rect 103 359 104 360 
<< pdiffusion >>
rect 104 359 105 360 
<< pdiffusion >>
rect 105 359 106 360 
<< pdiffusion >>
rect 106 359 107 360 
<< pdiffusion >>
rect 107 359 108 360 
<< pdiffusion >>
rect 120 359 121 360 
<< pdiffusion >>
rect 121 359 122 360 
<< pdiffusion >>
rect 122 359 123 360 
<< pdiffusion >>
rect 123 359 124 360 
<< pdiffusion >>
rect 124 359 125 360 
<< pdiffusion >>
rect 125 359 126 360 
<< m1 >>
rect 127 359 128 360 
<< m2 >>
rect 127 359 128 360 
<< pdiffusion >>
rect 138 359 139 360 
<< pdiffusion >>
rect 139 359 140 360 
<< pdiffusion >>
rect 140 359 141 360 
<< pdiffusion >>
rect 141 359 142 360 
<< pdiffusion >>
rect 142 359 143 360 
<< pdiffusion >>
rect 143 359 144 360 
<< pdiffusion >>
rect 156 359 157 360 
<< pdiffusion >>
rect 157 359 158 360 
<< pdiffusion >>
rect 158 359 159 360 
<< pdiffusion >>
rect 159 359 160 360 
<< m1 >>
rect 160 359 161 360 
<< pdiffusion >>
rect 160 359 161 360 
<< pdiffusion >>
rect 161 359 162 360 
<< m1 >>
rect 172 359 173 360 
<< pdiffusion >>
rect 174 359 175 360 
<< pdiffusion >>
rect 175 359 176 360 
<< pdiffusion >>
rect 176 359 177 360 
<< pdiffusion >>
rect 177 359 178 360 
<< pdiffusion >>
rect 178 359 179 360 
<< pdiffusion >>
rect 179 359 180 360 
<< pdiffusion >>
rect 192 359 193 360 
<< pdiffusion >>
rect 193 359 194 360 
<< pdiffusion >>
rect 194 359 195 360 
<< pdiffusion >>
rect 195 359 196 360 
<< m1 >>
rect 196 359 197 360 
<< pdiffusion >>
rect 196 359 197 360 
<< pdiffusion >>
rect 197 359 198 360 
<< pdiffusion >>
rect 210 359 211 360 
<< pdiffusion >>
rect 211 359 212 360 
<< pdiffusion >>
rect 212 359 213 360 
<< pdiffusion >>
rect 213 359 214 360 
<< m1 >>
rect 214 359 215 360 
<< pdiffusion >>
rect 214 359 215 360 
<< pdiffusion >>
rect 215 359 216 360 
<< m1 >>
rect 217 359 218 360 
<< pdiffusion >>
rect 228 359 229 360 
<< pdiffusion >>
rect 229 359 230 360 
<< pdiffusion >>
rect 230 359 231 360 
<< pdiffusion >>
rect 231 359 232 360 
<< pdiffusion >>
rect 232 359 233 360 
<< pdiffusion >>
rect 233 359 234 360 
<< m1 >>
rect 244 359 245 360 
<< pdiffusion >>
rect 246 359 247 360 
<< pdiffusion >>
rect 247 359 248 360 
<< pdiffusion >>
rect 248 359 249 360 
<< pdiffusion >>
rect 249 359 250 360 
<< m1 >>
rect 250 359 251 360 
<< pdiffusion >>
rect 250 359 251 360 
<< pdiffusion >>
rect 251 359 252 360 
<< m1 >>
rect 253 359 254 360 
<< m2 >>
rect 254 359 255 360 
<< pdiffusion >>
rect 264 359 265 360 
<< pdiffusion >>
rect 265 359 266 360 
<< pdiffusion >>
rect 266 359 267 360 
<< pdiffusion >>
rect 267 359 268 360 
<< m1 >>
rect 268 359 269 360 
<< pdiffusion >>
rect 268 359 269 360 
<< pdiffusion >>
rect 269 359 270 360 
<< pdiffusion >>
rect 282 359 283 360 
<< pdiffusion >>
rect 283 359 284 360 
<< pdiffusion >>
rect 284 359 285 360 
<< pdiffusion >>
rect 285 359 286 360 
<< pdiffusion >>
rect 286 359 287 360 
<< pdiffusion >>
rect 287 359 288 360 
<< m1 >>
rect 289 359 290 360 
<< m1 >>
rect 291 359 292 360 
<< m1 >>
rect 293 359 294 360 
<< pdiffusion >>
rect 300 359 301 360 
<< pdiffusion >>
rect 301 359 302 360 
<< pdiffusion >>
rect 302 359 303 360 
<< pdiffusion >>
rect 303 359 304 360 
<< pdiffusion >>
rect 304 359 305 360 
<< pdiffusion >>
rect 305 359 306 360 
<< pdiffusion >>
rect 318 359 319 360 
<< pdiffusion >>
rect 319 359 320 360 
<< pdiffusion >>
rect 320 359 321 360 
<< pdiffusion >>
rect 321 359 322 360 
<< pdiffusion >>
rect 322 359 323 360 
<< pdiffusion >>
rect 323 359 324 360 
<< m1 >>
rect 325 359 326 360 
<< pdiffusion >>
rect 336 359 337 360 
<< pdiffusion >>
rect 337 359 338 360 
<< pdiffusion >>
rect 338 359 339 360 
<< pdiffusion >>
rect 339 359 340 360 
<< m1 >>
rect 340 359 341 360 
<< pdiffusion >>
rect 340 359 341 360 
<< pdiffusion >>
rect 341 359 342 360 
<< pdiffusion >>
rect 354 359 355 360 
<< pdiffusion >>
rect 355 359 356 360 
<< pdiffusion >>
rect 356 359 357 360 
<< pdiffusion >>
rect 357 359 358 360 
<< m1 >>
rect 358 359 359 360 
<< pdiffusion >>
rect 358 359 359 360 
<< pdiffusion >>
rect 359 359 360 360 
<< pdiffusion >>
rect 372 359 373 360 
<< pdiffusion >>
rect 373 359 374 360 
<< pdiffusion >>
rect 374 359 375 360 
<< pdiffusion >>
rect 375 359 376 360 
<< pdiffusion >>
rect 376 359 377 360 
<< pdiffusion >>
rect 377 359 378 360 
<< m1 >>
rect 379 359 380 360 
<< pdiffusion >>
rect 390 359 391 360 
<< pdiffusion >>
rect 391 359 392 360 
<< pdiffusion >>
rect 392 359 393 360 
<< pdiffusion >>
rect 393 359 394 360 
<< pdiffusion >>
rect 394 359 395 360 
<< pdiffusion >>
rect 395 359 396 360 
<< pdiffusion >>
rect 408 359 409 360 
<< pdiffusion >>
rect 409 359 410 360 
<< pdiffusion >>
rect 410 359 411 360 
<< pdiffusion >>
rect 411 359 412 360 
<< m1 >>
rect 412 359 413 360 
<< pdiffusion >>
rect 412 359 413 360 
<< pdiffusion >>
rect 413 359 414 360 
<< pdiffusion >>
rect 444 359 445 360 
<< pdiffusion >>
rect 445 359 446 360 
<< pdiffusion >>
rect 446 359 447 360 
<< pdiffusion >>
rect 447 359 448 360 
<< pdiffusion >>
rect 448 359 449 360 
<< pdiffusion >>
rect 449 359 450 360 
<< m1 >>
rect 37 360 38 361 
<< m1 >>
rect 88 360 89 361 
<< m1 >>
rect 91 360 92 361 
<< m1 >>
rect 127 360 128 361 
<< m2 >>
rect 127 360 128 361 
<< m1 >>
rect 160 360 161 361 
<< m2 >>
rect 164 360 165 361 
<< m1 >>
rect 165 360 166 361 
<< m2 >>
rect 165 360 166 361 
<< m2c >>
rect 165 360 166 361 
<< m1 >>
rect 165 360 166 361 
<< m2 >>
rect 165 360 166 361 
<< m1 >>
rect 166 360 167 361 
<< m1 >>
rect 167 360 168 361 
<< m1 >>
rect 168 360 169 361 
<< m1 >>
rect 169 360 170 361 
<< m1 >>
rect 170 360 171 361 
<< m1 >>
rect 171 360 172 361 
<< m1 >>
rect 172 360 173 361 
<< m1 >>
rect 196 360 197 361 
<< m1 >>
rect 214 360 215 361 
<< m1 >>
rect 217 360 218 361 
<< m1 >>
rect 244 360 245 361 
<< m1 >>
rect 250 360 251 361 
<< m1 >>
rect 253 360 254 361 
<< m2 >>
rect 254 360 255 361 
<< m1 >>
rect 268 360 269 361 
<< m1 >>
rect 289 360 290 361 
<< m1 >>
rect 291 360 292 361 
<< m1 >>
rect 293 360 294 361 
<< m1 >>
rect 325 360 326 361 
<< m1 >>
rect 340 360 341 361 
<< m1 >>
rect 358 360 359 361 
<< m1 >>
rect 379 360 380 361 
<< m1 >>
rect 412 360 413 361 
<< m1 >>
rect 37 361 38 362 
<< m1 >>
rect 88 361 89 362 
<< m1 >>
rect 89 361 90 362 
<< m1 >>
rect 90 361 91 362 
<< m1 >>
rect 91 361 92 362 
<< m1 >>
rect 127 361 128 362 
<< m2 >>
rect 127 361 128 362 
<< m1 >>
rect 160 361 161 362 
<< m1 >>
rect 161 361 162 362 
<< m1 >>
rect 162 361 163 362 
<< m1 >>
rect 163 361 164 362 
<< m2 >>
rect 164 361 165 362 
<< m1 >>
rect 196 361 197 362 
<< m1 >>
rect 214 361 215 362 
<< m1 >>
rect 217 361 218 362 
<< m1 >>
rect 244 361 245 362 
<< m1 >>
rect 250 361 251 362 
<< m1 >>
rect 251 361 252 362 
<< m2 >>
rect 251 361 252 362 
<< m2c >>
rect 251 361 252 362 
<< m1 >>
rect 251 361 252 362 
<< m2 >>
rect 251 361 252 362 
<< m2 >>
rect 252 361 253 362 
<< m1 >>
rect 253 361 254 362 
<< m2 >>
rect 253 361 254 362 
<< m2 >>
rect 254 361 255 362 
<< m1 >>
rect 268 361 269 362 
<< m1 >>
rect 289 361 290 362 
<< m1 >>
rect 291 361 292 362 
<< m1 >>
rect 293 361 294 362 
<< m1 >>
rect 325 361 326 362 
<< m1 >>
rect 340 361 341 362 
<< m1 >>
rect 358 361 359 362 
<< m1 >>
rect 379 361 380 362 
<< m1 >>
rect 412 361 413 362 
<< m1 >>
rect 413 361 414 362 
<< m1 >>
rect 414 361 415 362 
<< m1 >>
rect 415 361 416 362 
<< m1 >>
rect 37 362 38 363 
<< m1 >>
rect 127 362 128 363 
<< m2 >>
rect 127 362 128 363 
<< m1 >>
rect 163 362 164 363 
<< m2 >>
rect 164 362 165 363 
<< m1 >>
rect 196 362 197 363 
<< m1 >>
rect 214 362 215 363 
<< m1 >>
rect 217 362 218 363 
<< m1 >>
rect 244 362 245 363 
<< m1 >>
rect 253 362 254 363 
<< m1 >>
rect 268 362 269 363 
<< m1 >>
rect 289 362 290 363 
<< m1 >>
rect 291 362 292 363 
<< m1 >>
rect 293 362 294 363 
<< m1 >>
rect 325 362 326 363 
<< m1 >>
rect 340 362 341 363 
<< m1 >>
rect 341 362 342 363 
<< m1 >>
rect 342 362 343 363 
<< m1 >>
rect 343 362 344 363 
<< m1 >>
rect 344 362 345 363 
<< m1 >>
rect 345 362 346 363 
<< m1 >>
rect 346 362 347 363 
<< m1 >>
rect 347 362 348 363 
<< m1 >>
rect 348 362 349 363 
<< m1 >>
rect 349 362 350 363 
<< m1 >>
rect 350 362 351 363 
<< m1 >>
rect 351 362 352 363 
<< m1 >>
rect 352 362 353 363 
<< m1 >>
rect 353 362 354 363 
<< m1 >>
rect 354 362 355 363 
<< m2 >>
rect 354 362 355 363 
<< m2c >>
rect 354 362 355 363 
<< m1 >>
rect 354 362 355 363 
<< m2 >>
rect 354 362 355 363 
<< m1 >>
rect 358 362 359 363 
<< m2 >>
rect 358 362 359 363 
<< m2c >>
rect 358 362 359 363 
<< m1 >>
rect 358 362 359 363 
<< m2 >>
rect 358 362 359 363 
<< m1 >>
rect 379 362 380 363 
<< m1 >>
rect 415 362 416 363 
<< m1 >>
rect 37 363 38 364 
<< m1 >>
rect 127 363 128 364 
<< m2 >>
rect 127 363 128 364 
<< m1 >>
rect 163 363 164 364 
<< m2 >>
rect 164 363 165 364 
<< m1 >>
rect 196 363 197 364 
<< m1 >>
rect 214 363 215 364 
<< m1 >>
rect 217 363 218 364 
<< m1 >>
rect 244 363 245 364 
<< m1 >>
rect 253 363 254 364 
<< m1 >>
rect 268 363 269 364 
<< m1 >>
rect 289 363 290 364 
<< m1 >>
rect 291 363 292 364 
<< m1 >>
rect 293 363 294 364 
<< m1 >>
rect 325 363 326 364 
<< m2 >>
rect 354 363 355 364 
<< m2 >>
rect 358 363 359 364 
<< m1 >>
rect 379 363 380 364 
<< m1 >>
rect 415 363 416 364 
<< m1 >>
rect 37 364 38 365 
<< m1 >>
rect 38 364 39 365 
<< m1 >>
rect 39 364 40 365 
<< m1 >>
rect 40 364 41 365 
<< m1 >>
rect 41 364 42 365 
<< m1 >>
rect 42 364 43 365 
<< m1 >>
rect 43 364 44 365 
<< m1 >>
rect 44 364 45 365 
<< m1 >>
rect 45 364 46 365 
<< m1 >>
rect 46 364 47 365 
<< m1 >>
rect 47 364 48 365 
<< m1 >>
rect 48 364 49 365 
<< m1 >>
rect 49 364 50 365 
<< m1 >>
rect 50 364 51 365 
<< m1 >>
rect 51 364 52 365 
<< m1 >>
rect 52 364 53 365 
<< m1 >>
rect 53 364 54 365 
<< m1 >>
rect 54 364 55 365 
<< m1 >>
rect 55 364 56 365 
<< m1 >>
rect 56 364 57 365 
<< m1 >>
rect 57 364 58 365 
<< m1 >>
rect 58 364 59 365 
<< m1 >>
rect 59 364 60 365 
<< m1 >>
rect 60 364 61 365 
<< m1 >>
rect 61 364 62 365 
<< m1 >>
rect 62 364 63 365 
<< m1 >>
rect 63 364 64 365 
<< m1 >>
rect 64 364 65 365 
<< m1 >>
rect 65 364 66 365 
<< m1 >>
rect 66 364 67 365 
<< m1 >>
rect 67 364 68 365 
<< m1 >>
rect 68 364 69 365 
<< m1 >>
rect 69 364 70 365 
<< m1 >>
rect 70 364 71 365 
<< m1 >>
rect 127 364 128 365 
<< m2 >>
rect 127 364 128 365 
<< m1 >>
rect 128 364 129 365 
<< m1 >>
rect 129 364 130 365 
<< m1 >>
rect 130 364 131 365 
<< m1 >>
rect 131 364 132 365 
<< m1 >>
rect 132 364 133 365 
<< m1 >>
rect 133 364 134 365 
<< m1 >>
rect 134 364 135 365 
<< m1 >>
rect 135 364 136 365 
<< m1 >>
rect 136 364 137 365 
<< m1 >>
rect 137 364 138 365 
<< m1 >>
rect 138 364 139 365 
<< m1 >>
rect 139 364 140 365 
<< m1 >>
rect 140 364 141 365 
<< m1 >>
rect 141 364 142 365 
<< m1 >>
rect 142 364 143 365 
<< m1 >>
rect 143 364 144 365 
<< m1 >>
rect 144 364 145 365 
<< m1 >>
rect 145 364 146 365 
<< m1 >>
rect 146 364 147 365 
<< m1 >>
rect 147 364 148 365 
<< m1 >>
rect 148 364 149 365 
<< m1 >>
rect 149 364 150 365 
<< m1 >>
rect 150 364 151 365 
<< m1 >>
rect 151 364 152 365 
<< m1 >>
rect 152 364 153 365 
<< m1 >>
rect 153 364 154 365 
<< m1 >>
rect 154 364 155 365 
<< m1 >>
rect 155 364 156 365 
<< m1 >>
rect 156 364 157 365 
<< m1 >>
rect 157 364 158 365 
<< m1 >>
rect 163 364 164 365 
<< m2 >>
rect 164 364 165 365 
<< m1 >>
rect 196 364 197 365 
<< m1 >>
rect 197 364 198 365 
<< m1 >>
rect 198 364 199 365 
<< m1 >>
rect 199 364 200 365 
<< m1 >>
rect 200 364 201 365 
<< m1 >>
rect 201 364 202 365 
<< m1 >>
rect 202 364 203 365 
<< m1 >>
rect 203 364 204 365 
<< m1 >>
rect 204 364 205 365 
<< m1 >>
rect 205 364 206 365 
<< m1 >>
rect 206 364 207 365 
<< m1 >>
rect 207 364 208 365 
<< m1 >>
rect 208 364 209 365 
<< m1 >>
rect 209 364 210 365 
<< m1 >>
rect 210 364 211 365 
<< m1 >>
rect 211 364 212 365 
<< m1 >>
rect 212 364 213 365 
<< m1 >>
rect 213 364 214 365 
<< m1 >>
rect 214 364 215 365 
<< m1 >>
rect 217 364 218 365 
<< m1 >>
rect 244 364 245 365 
<< m1 >>
rect 253 364 254 365 
<< m1 >>
rect 268 364 269 365 
<< m1 >>
rect 289 364 290 365 
<< m1 >>
rect 291 364 292 365 
<< m1 >>
rect 293 364 294 365 
<< m1 >>
rect 325 364 326 365 
<< m1 >>
rect 326 364 327 365 
<< m1 >>
rect 327 364 328 365 
<< m1 >>
rect 328 364 329 365 
<< m1 >>
rect 329 364 330 365 
<< m1 >>
rect 330 364 331 365 
<< m1 >>
rect 331 364 332 365 
<< m1 >>
rect 332 364 333 365 
<< m1 >>
rect 333 364 334 365 
<< m1 >>
rect 334 364 335 365 
<< m1 >>
rect 335 364 336 365 
<< m1 >>
rect 336 364 337 365 
<< m1 >>
rect 337 364 338 365 
<< m1 >>
rect 338 364 339 365 
<< m1 >>
rect 339 364 340 365 
<< m1 >>
rect 340 364 341 365 
<< m1 >>
rect 341 364 342 365 
<< m1 >>
rect 342 364 343 365 
<< m1 >>
rect 343 364 344 365 
<< m1 >>
rect 344 364 345 365 
<< m1 >>
rect 345 364 346 365 
<< m1 >>
rect 346 364 347 365 
<< m1 >>
rect 347 364 348 365 
<< m1 >>
rect 348 364 349 365 
<< m1 >>
rect 349 364 350 365 
<< m1 >>
rect 350 364 351 365 
<< m1 >>
rect 351 364 352 365 
<< m1 >>
rect 352 364 353 365 
<< m1 >>
rect 353 364 354 365 
<< m1 >>
rect 354 364 355 365 
<< m2 >>
rect 354 364 355 365 
<< m1 >>
rect 355 364 356 365 
<< m2 >>
rect 355 364 356 365 
<< m1 >>
rect 356 364 357 365 
<< m2 >>
rect 356 364 357 365 
<< m1 >>
rect 357 364 358 365 
<< m2 >>
rect 357 364 358 365 
<< m1 >>
rect 358 364 359 365 
<< m2 >>
rect 358 364 359 365 
<< m1 >>
rect 379 364 380 365 
<< m1 >>
rect 415 364 416 365 
<< m1 >>
rect 70 365 71 366 
<< m2 >>
rect 127 365 128 366 
<< m1 >>
rect 157 365 158 366 
<< m1 >>
rect 163 365 164 366 
<< m2 >>
rect 164 365 165 366 
<< m1 >>
rect 217 365 218 366 
<< m1 >>
rect 244 365 245 366 
<< m1 >>
rect 253 365 254 366 
<< m1 >>
rect 268 365 269 366 
<< m1 >>
rect 289 365 290 366 
<< m1 >>
rect 291 365 292 366 
<< m1 >>
rect 293 365 294 366 
<< m1 >>
rect 358 365 359 366 
<< m1 >>
rect 379 365 380 366 
<< m1 >>
rect 415 365 416 366 
<< m1 >>
rect 70 366 71 367 
<< m2 >>
rect 127 366 128 367 
<< m1 >>
rect 157 366 158 367 
<< m1 >>
rect 163 366 164 367 
<< m2 >>
rect 164 366 165 367 
<< m1 >>
rect 217 366 218 367 
<< m1 >>
rect 244 366 245 367 
<< m1 >>
rect 253 366 254 367 
<< m1 >>
rect 268 366 269 367 
<< m1 >>
rect 289 366 290 367 
<< m1 >>
rect 291 366 292 367 
<< m1 >>
rect 293 366 294 367 
<< m1 >>
rect 358 366 359 367 
<< m1 >>
rect 379 366 380 367 
<< m1 >>
rect 415 366 416 367 
<< m1 >>
rect 70 367 71 368 
<< m1 >>
rect 100 367 101 368 
<< m1 >>
rect 101 367 102 368 
<< m1 >>
rect 102 367 103 368 
<< m1 >>
rect 103 367 104 368 
<< m1 >>
rect 104 367 105 368 
<< m1 >>
rect 105 367 106 368 
<< m1 >>
rect 106 367 107 368 
<< m1 >>
rect 107 367 108 368 
<< m1 >>
rect 108 367 109 368 
<< m1 >>
rect 109 367 110 368 
<< m1 >>
rect 110 367 111 368 
<< m1 >>
rect 111 367 112 368 
<< m1 >>
rect 112 367 113 368 
<< m1 >>
rect 113 367 114 368 
<< m1 >>
rect 114 367 115 368 
<< m1 >>
rect 115 367 116 368 
<< m1 >>
rect 116 367 117 368 
<< m1 >>
rect 117 367 118 368 
<< m1 >>
rect 118 367 119 368 
<< m1 >>
rect 119 367 120 368 
<< m1 >>
rect 120 367 121 368 
<< m1 >>
rect 121 367 122 368 
<< m1 >>
rect 122 367 123 368 
<< m1 >>
rect 123 367 124 368 
<< m1 >>
rect 124 367 125 368 
<< m1 >>
rect 125 367 126 368 
<< m1 >>
rect 126 367 127 368 
<< m1 >>
rect 127 367 128 368 
<< m2 >>
rect 127 367 128 368 
<< m1 >>
rect 128 367 129 368 
<< m1 >>
rect 129 367 130 368 
<< m1 >>
rect 130 367 131 368 
<< m1 >>
rect 131 367 132 368 
<< m1 >>
rect 132 367 133 368 
<< m1 >>
rect 133 367 134 368 
<< m1 >>
rect 134 367 135 368 
<< m1 >>
rect 135 367 136 368 
<< m1 >>
rect 136 367 137 368 
<< m1 >>
rect 137 367 138 368 
<< m1 >>
rect 138 367 139 368 
<< m1 >>
rect 139 367 140 368 
<< m1 >>
rect 140 367 141 368 
<< m1 >>
rect 141 367 142 368 
<< m1 >>
rect 142 367 143 368 
<< m1 >>
rect 143 367 144 368 
<< m1 >>
rect 144 367 145 368 
<< m1 >>
rect 145 367 146 368 
<< m1 >>
rect 146 367 147 368 
<< m1 >>
rect 147 367 148 368 
<< m1 >>
rect 148 367 149 368 
<< m1 >>
rect 149 367 150 368 
<< m1 >>
rect 150 367 151 368 
<< m1 >>
rect 151 367 152 368 
<< m1 >>
rect 152 367 153 368 
<< m1 >>
rect 153 367 154 368 
<< m1 >>
rect 154 367 155 368 
<< m1 >>
rect 155 367 156 368 
<< m2 >>
rect 155 367 156 368 
<< m2c >>
rect 155 367 156 368 
<< m1 >>
rect 155 367 156 368 
<< m2 >>
rect 155 367 156 368 
<< m2 >>
rect 156 367 157 368 
<< m1 >>
rect 157 367 158 368 
<< m2 >>
rect 157 367 158 368 
<< m2 >>
rect 158 367 159 368 
<< m1 >>
rect 163 367 164 368 
<< m2 >>
rect 164 367 165 368 
<< m1 >>
rect 217 367 218 368 
<< m1 >>
rect 244 367 245 368 
<< m1 >>
rect 253 367 254 368 
<< m1 >>
rect 255 367 256 368 
<< m1 >>
rect 256 367 257 368 
<< m1 >>
rect 257 367 258 368 
<< m1 >>
rect 258 367 259 368 
<< m1 >>
rect 259 367 260 368 
<< m1 >>
rect 260 367 261 368 
<< m1 >>
rect 261 367 262 368 
<< m1 >>
rect 262 367 263 368 
<< m1 >>
rect 263 367 264 368 
<< m1 >>
rect 264 367 265 368 
<< m1 >>
rect 265 367 266 368 
<< m1 >>
rect 266 367 267 368 
<< m1 >>
rect 267 367 268 368 
<< m1 >>
rect 268 367 269 368 
<< m1 >>
rect 289 367 290 368 
<< m1 >>
rect 291 367 292 368 
<< m1 >>
rect 293 367 294 368 
<< m1 >>
rect 358 367 359 368 
<< m1 >>
rect 379 367 380 368 
<< m1 >>
rect 415 367 416 368 
<< m1 >>
rect 70 368 71 369 
<< m1 >>
rect 100 368 101 369 
<< m2 >>
rect 127 368 128 369 
<< m1 >>
rect 157 368 158 369 
<< m2 >>
rect 158 368 159 369 
<< m1 >>
rect 163 368 164 369 
<< m2 >>
rect 164 368 165 369 
<< m1 >>
rect 217 368 218 369 
<< m1 >>
rect 244 368 245 369 
<< m1 >>
rect 253 368 254 369 
<< m1 >>
rect 255 368 256 369 
<< m1 >>
rect 289 368 290 369 
<< m1 >>
rect 291 368 292 369 
<< m1 >>
rect 293 368 294 369 
<< m1 >>
rect 358 368 359 369 
<< m1 >>
rect 379 368 380 369 
<< m1 >>
rect 415 368 416 369 
<< m1 >>
rect 67 369 68 370 
<< m1 >>
rect 68 369 69 370 
<< m2 >>
rect 68 369 69 370 
<< m2c >>
rect 68 369 69 370 
<< m1 >>
rect 68 369 69 370 
<< m2 >>
rect 68 369 69 370 
<< m2 >>
rect 69 369 70 370 
<< m1 >>
rect 70 369 71 370 
<< m2 >>
rect 70 369 71 370 
<< m2 >>
rect 71 369 72 370 
<< m1 >>
rect 100 369 101 370 
<< m1 >>
rect 127 369 128 370 
<< m2 >>
rect 127 369 128 370 
<< m2c >>
rect 127 369 128 370 
<< m1 >>
rect 127 369 128 370 
<< m2 >>
rect 127 369 128 370 
<< m1 >>
rect 157 369 158 370 
<< m2 >>
rect 158 369 159 370 
<< m1 >>
rect 163 369 164 370 
<< m2 >>
rect 164 369 165 370 
<< m1 >>
rect 217 369 218 370 
<< m1 >>
rect 244 369 245 370 
<< m1 >>
rect 253 369 254 370 
<< m1 >>
rect 255 369 256 370 
<< m1 >>
rect 283 369 284 370 
<< m1 >>
rect 284 369 285 370 
<< m1 >>
rect 285 369 286 370 
<< m1 >>
rect 286 369 287 370 
<< m1 >>
rect 287 369 288 370 
<< m2 >>
rect 287 369 288 370 
<< m2c >>
rect 287 369 288 370 
<< m1 >>
rect 287 369 288 370 
<< m2 >>
rect 287 369 288 370 
<< m2 >>
rect 288 369 289 370 
<< m1 >>
rect 289 369 290 370 
<< m2 >>
rect 289 369 290 370 
<< m2 >>
rect 290 369 291 370 
<< m1 >>
rect 291 369 292 370 
<< m2 >>
rect 291 369 292 370 
<< m2c >>
rect 291 369 292 370 
<< m1 >>
rect 291 369 292 370 
<< m2 >>
rect 291 369 292 370 
<< m1 >>
rect 293 369 294 370 
<< m1 >>
rect 358 369 359 370 
<< m1 >>
rect 379 369 380 370 
<< m1 >>
rect 415 369 416 370 
<< m1 >>
rect 67 370 68 371 
<< m1 >>
rect 70 370 71 371 
<< m2 >>
rect 71 370 72 371 
<< m1 >>
rect 72 370 73 371 
<< m2 >>
rect 72 370 73 371 
<< m2c >>
rect 72 370 73 371 
<< m1 >>
rect 72 370 73 371 
<< m2 >>
rect 72 370 73 371 
<< m1 >>
rect 73 370 74 371 
<< m1 >>
rect 74 370 75 371 
<< m1 >>
rect 75 370 76 371 
<< m1 >>
rect 76 370 77 371 
<< m1 >>
rect 77 370 78 371 
<< m1 >>
rect 78 370 79 371 
<< m1 >>
rect 79 370 80 371 
<< m1 >>
rect 80 370 81 371 
<< m1 >>
rect 81 370 82 371 
<< m1 >>
rect 82 370 83 371 
<< m1 >>
rect 100 370 101 371 
<< m1 >>
rect 127 370 128 371 
<< m1 >>
rect 142 370 143 371 
<< m1 >>
rect 143 370 144 371 
<< m1 >>
rect 144 370 145 371 
<< m1 >>
rect 145 370 146 371 
<< m1 >>
rect 157 370 158 371 
<< m2 >>
rect 158 370 159 371 
<< m1 >>
rect 159 370 160 371 
<< m2 >>
rect 159 370 160 371 
<< m2c >>
rect 159 370 160 371 
<< m1 >>
rect 159 370 160 371 
<< m2 >>
rect 159 370 160 371 
<< m1 >>
rect 160 370 161 371 
<< m1 >>
rect 163 370 164 371 
<< m2 >>
rect 164 370 165 371 
<< m1 >>
rect 217 370 218 371 
<< m1 >>
rect 244 370 245 371 
<< m1 >>
rect 253 370 254 371 
<< m1 >>
rect 255 370 256 371 
<< m1 >>
rect 283 370 284 371 
<< m1 >>
rect 289 370 290 371 
<< m1 >>
rect 293 370 294 371 
<< m1 >>
rect 358 370 359 371 
<< m1 >>
rect 379 370 380 371 
<< m1 >>
rect 415 370 416 371 
<< m1 >>
rect 67 371 68 372 
<< m1 >>
rect 70 371 71 372 
<< m1 >>
rect 82 371 83 372 
<< m1 >>
rect 100 371 101 372 
<< m1 >>
rect 127 371 128 372 
<< m1 >>
rect 142 371 143 372 
<< m1 >>
rect 145 371 146 372 
<< m1 >>
rect 157 371 158 372 
<< m1 >>
rect 160 371 161 372 
<< m1 >>
rect 163 371 164 372 
<< m2 >>
rect 164 371 165 372 
<< m1 >>
rect 217 371 218 372 
<< m1 >>
rect 244 371 245 372 
<< m1 >>
rect 253 371 254 372 
<< m1 >>
rect 255 371 256 372 
<< m1 >>
rect 283 371 284 372 
<< m1 >>
rect 289 371 290 372 
<< m1 >>
rect 293 371 294 372 
<< m1 >>
rect 358 371 359 372 
<< m1 >>
rect 379 371 380 372 
<< m1 >>
rect 415 371 416 372 
<< pdiffusion >>
rect 12 372 13 373 
<< pdiffusion >>
rect 13 372 14 373 
<< pdiffusion >>
rect 14 372 15 373 
<< pdiffusion >>
rect 15 372 16 373 
<< pdiffusion >>
rect 16 372 17 373 
<< pdiffusion >>
rect 17 372 18 373 
<< pdiffusion >>
rect 30 372 31 373 
<< pdiffusion >>
rect 31 372 32 373 
<< pdiffusion >>
rect 32 372 33 373 
<< pdiffusion >>
rect 33 372 34 373 
<< pdiffusion >>
rect 34 372 35 373 
<< pdiffusion >>
rect 35 372 36 373 
<< pdiffusion >>
rect 48 372 49 373 
<< pdiffusion >>
rect 49 372 50 373 
<< pdiffusion >>
rect 50 372 51 373 
<< pdiffusion >>
rect 51 372 52 373 
<< pdiffusion >>
rect 52 372 53 373 
<< pdiffusion >>
rect 53 372 54 373 
<< pdiffusion >>
rect 66 372 67 373 
<< m1 >>
rect 67 372 68 373 
<< pdiffusion >>
rect 67 372 68 373 
<< pdiffusion >>
rect 68 372 69 373 
<< pdiffusion >>
rect 69 372 70 373 
<< m1 >>
rect 70 372 71 373 
<< pdiffusion >>
rect 70 372 71 373 
<< pdiffusion >>
rect 71 372 72 373 
<< m1 >>
rect 82 372 83 373 
<< pdiffusion >>
rect 84 372 85 373 
<< pdiffusion >>
rect 85 372 86 373 
<< pdiffusion >>
rect 86 372 87 373 
<< pdiffusion >>
rect 87 372 88 373 
<< pdiffusion >>
rect 88 372 89 373 
<< pdiffusion >>
rect 89 372 90 373 
<< m1 >>
rect 100 372 101 373 
<< pdiffusion >>
rect 102 372 103 373 
<< pdiffusion >>
rect 103 372 104 373 
<< pdiffusion >>
rect 104 372 105 373 
<< pdiffusion >>
rect 105 372 106 373 
<< pdiffusion >>
rect 106 372 107 373 
<< pdiffusion >>
rect 107 372 108 373 
<< pdiffusion >>
rect 120 372 121 373 
<< pdiffusion >>
rect 121 372 122 373 
<< pdiffusion >>
rect 122 372 123 373 
<< pdiffusion >>
rect 123 372 124 373 
<< pdiffusion >>
rect 124 372 125 373 
<< pdiffusion >>
rect 125 372 126 373 
<< m1 >>
rect 127 372 128 373 
<< pdiffusion >>
rect 138 372 139 373 
<< pdiffusion >>
rect 139 372 140 373 
<< pdiffusion >>
rect 140 372 141 373 
<< pdiffusion >>
rect 141 372 142 373 
<< m1 >>
rect 142 372 143 373 
<< pdiffusion >>
rect 142 372 143 373 
<< pdiffusion >>
rect 143 372 144 373 
<< m1 >>
rect 145 372 146 373 
<< pdiffusion >>
rect 156 372 157 373 
<< m1 >>
rect 157 372 158 373 
<< pdiffusion >>
rect 157 372 158 373 
<< pdiffusion >>
rect 158 372 159 373 
<< pdiffusion >>
rect 159 372 160 373 
<< m1 >>
rect 160 372 161 373 
<< pdiffusion >>
rect 160 372 161 373 
<< pdiffusion >>
rect 161 372 162 373 
<< m1 >>
rect 163 372 164 373 
<< m2 >>
rect 164 372 165 373 
<< pdiffusion >>
rect 174 372 175 373 
<< pdiffusion >>
rect 175 372 176 373 
<< pdiffusion >>
rect 176 372 177 373 
<< pdiffusion >>
rect 177 372 178 373 
<< pdiffusion >>
rect 178 372 179 373 
<< pdiffusion >>
rect 179 372 180 373 
<< pdiffusion >>
rect 210 372 211 373 
<< pdiffusion >>
rect 211 372 212 373 
<< pdiffusion >>
rect 212 372 213 373 
<< pdiffusion >>
rect 213 372 214 373 
<< pdiffusion >>
rect 214 372 215 373 
<< pdiffusion >>
rect 215 372 216 373 
<< m1 >>
rect 217 372 218 373 
<< pdiffusion >>
rect 228 372 229 373 
<< pdiffusion >>
rect 229 372 230 373 
<< pdiffusion >>
rect 230 372 231 373 
<< pdiffusion >>
rect 231 372 232 373 
<< pdiffusion >>
rect 232 372 233 373 
<< pdiffusion >>
rect 233 372 234 373 
<< m1 >>
rect 244 372 245 373 
<< pdiffusion >>
rect 246 372 247 373 
<< pdiffusion >>
rect 247 372 248 373 
<< pdiffusion >>
rect 248 372 249 373 
<< pdiffusion >>
rect 249 372 250 373 
<< pdiffusion >>
rect 250 372 251 373 
<< pdiffusion >>
rect 251 372 252 373 
<< m1 >>
rect 253 372 254 373 
<< m1 >>
rect 255 372 256 373 
<< pdiffusion >>
rect 264 372 265 373 
<< pdiffusion >>
rect 265 372 266 373 
<< pdiffusion >>
rect 266 372 267 373 
<< pdiffusion >>
rect 267 372 268 373 
<< pdiffusion >>
rect 268 372 269 373 
<< pdiffusion >>
rect 269 372 270 373 
<< pdiffusion >>
rect 282 372 283 373 
<< m1 >>
rect 283 372 284 373 
<< pdiffusion >>
rect 283 372 284 373 
<< pdiffusion >>
rect 284 372 285 373 
<< pdiffusion >>
rect 285 372 286 373 
<< pdiffusion >>
rect 286 372 287 373 
<< pdiffusion >>
rect 287 372 288 373 
<< m1 >>
rect 289 372 290 373 
<< m1 >>
rect 293 372 294 373 
<< pdiffusion >>
rect 300 372 301 373 
<< pdiffusion >>
rect 301 372 302 373 
<< pdiffusion >>
rect 302 372 303 373 
<< pdiffusion >>
rect 303 372 304 373 
<< pdiffusion >>
rect 304 372 305 373 
<< pdiffusion >>
rect 305 372 306 373 
<< pdiffusion >>
rect 318 372 319 373 
<< pdiffusion >>
rect 319 372 320 373 
<< pdiffusion >>
rect 320 372 321 373 
<< pdiffusion >>
rect 321 372 322 373 
<< pdiffusion >>
rect 322 372 323 373 
<< pdiffusion >>
rect 323 372 324 373 
<< pdiffusion >>
rect 336 372 337 373 
<< pdiffusion >>
rect 337 372 338 373 
<< pdiffusion >>
rect 338 372 339 373 
<< pdiffusion >>
rect 339 372 340 373 
<< pdiffusion >>
rect 340 372 341 373 
<< pdiffusion >>
rect 341 372 342 373 
<< pdiffusion >>
rect 354 372 355 373 
<< pdiffusion >>
rect 355 372 356 373 
<< pdiffusion >>
rect 356 372 357 373 
<< pdiffusion >>
rect 357 372 358 373 
<< m1 >>
rect 358 372 359 373 
<< pdiffusion >>
rect 358 372 359 373 
<< pdiffusion >>
rect 359 372 360 373 
<< pdiffusion >>
rect 372 372 373 373 
<< pdiffusion >>
rect 373 372 374 373 
<< pdiffusion >>
rect 374 372 375 373 
<< pdiffusion >>
rect 375 372 376 373 
<< pdiffusion >>
rect 376 372 377 373 
<< pdiffusion >>
rect 377 372 378 373 
<< m1 >>
rect 379 372 380 373 
<< pdiffusion >>
rect 390 372 391 373 
<< pdiffusion >>
rect 391 372 392 373 
<< pdiffusion >>
rect 392 372 393 373 
<< pdiffusion >>
rect 393 372 394 373 
<< pdiffusion >>
rect 394 372 395 373 
<< pdiffusion >>
rect 395 372 396 373 
<< pdiffusion >>
rect 408 372 409 373 
<< pdiffusion >>
rect 409 372 410 373 
<< pdiffusion >>
rect 410 372 411 373 
<< pdiffusion >>
rect 411 372 412 373 
<< pdiffusion >>
rect 412 372 413 373 
<< pdiffusion >>
rect 413 372 414 373 
<< m1 >>
rect 415 372 416 373 
<< pdiffusion >>
rect 426 372 427 373 
<< pdiffusion >>
rect 427 372 428 373 
<< pdiffusion >>
rect 428 372 429 373 
<< pdiffusion >>
rect 429 372 430 373 
<< pdiffusion >>
rect 430 372 431 373 
<< pdiffusion >>
rect 431 372 432 373 
<< pdiffusion >>
rect 444 372 445 373 
<< pdiffusion >>
rect 445 372 446 373 
<< pdiffusion >>
rect 446 372 447 373 
<< pdiffusion >>
rect 447 372 448 373 
<< pdiffusion >>
rect 448 372 449 373 
<< pdiffusion >>
rect 449 372 450 373 
<< pdiffusion >>
rect 12 373 13 374 
<< pdiffusion >>
rect 13 373 14 374 
<< pdiffusion >>
rect 14 373 15 374 
<< pdiffusion >>
rect 15 373 16 374 
<< pdiffusion >>
rect 16 373 17 374 
<< pdiffusion >>
rect 17 373 18 374 
<< pdiffusion >>
rect 30 373 31 374 
<< pdiffusion >>
rect 31 373 32 374 
<< pdiffusion >>
rect 32 373 33 374 
<< pdiffusion >>
rect 33 373 34 374 
<< pdiffusion >>
rect 34 373 35 374 
<< pdiffusion >>
rect 35 373 36 374 
<< pdiffusion >>
rect 48 373 49 374 
<< pdiffusion >>
rect 49 373 50 374 
<< pdiffusion >>
rect 50 373 51 374 
<< pdiffusion >>
rect 51 373 52 374 
<< pdiffusion >>
rect 52 373 53 374 
<< pdiffusion >>
rect 53 373 54 374 
<< pdiffusion >>
rect 66 373 67 374 
<< pdiffusion >>
rect 67 373 68 374 
<< pdiffusion >>
rect 68 373 69 374 
<< pdiffusion >>
rect 69 373 70 374 
<< pdiffusion >>
rect 70 373 71 374 
<< pdiffusion >>
rect 71 373 72 374 
<< m1 >>
rect 82 373 83 374 
<< pdiffusion >>
rect 84 373 85 374 
<< pdiffusion >>
rect 85 373 86 374 
<< pdiffusion >>
rect 86 373 87 374 
<< pdiffusion >>
rect 87 373 88 374 
<< pdiffusion >>
rect 88 373 89 374 
<< pdiffusion >>
rect 89 373 90 374 
<< m1 >>
rect 100 373 101 374 
<< pdiffusion >>
rect 102 373 103 374 
<< pdiffusion >>
rect 103 373 104 374 
<< pdiffusion >>
rect 104 373 105 374 
<< pdiffusion >>
rect 105 373 106 374 
<< pdiffusion >>
rect 106 373 107 374 
<< pdiffusion >>
rect 107 373 108 374 
<< pdiffusion >>
rect 120 373 121 374 
<< pdiffusion >>
rect 121 373 122 374 
<< pdiffusion >>
rect 122 373 123 374 
<< pdiffusion >>
rect 123 373 124 374 
<< pdiffusion >>
rect 124 373 125 374 
<< pdiffusion >>
rect 125 373 126 374 
<< m1 >>
rect 127 373 128 374 
<< pdiffusion >>
rect 138 373 139 374 
<< pdiffusion >>
rect 139 373 140 374 
<< pdiffusion >>
rect 140 373 141 374 
<< pdiffusion >>
rect 141 373 142 374 
<< pdiffusion >>
rect 142 373 143 374 
<< pdiffusion >>
rect 143 373 144 374 
<< m1 >>
rect 145 373 146 374 
<< pdiffusion >>
rect 156 373 157 374 
<< pdiffusion >>
rect 157 373 158 374 
<< pdiffusion >>
rect 158 373 159 374 
<< pdiffusion >>
rect 159 373 160 374 
<< pdiffusion >>
rect 160 373 161 374 
<< pdiffusion >>
rect 161 373 162 374 
<< m1 >>
rect 163 373 164 374 
<< m2 >>
rect 164 373 165 374 
<< pdiffusion >>
rect 174 373 175 374 
<< pdiffusion >>
rect 175 373 176 374 
<< pdiffusion >>
rect 176 373 177 374 
<< pdiffusion >>
rect 177 373 178 374 
<< pdiffusion >>
rect 178 373 179 374 
<< pdiffusion >>
rect 179 373 180 374 
<< pdiffusion >>
rect 210 373 211 374 
<< pdiffusion >>
rect 211 373 212 374 
<< pdiffusion >>
rect 212 373 213 374 
<< pdiffusion >>
rect 213 373 214 374 
<< pdiffusion >>
rect 214 373 215 374 
<< pdiffusion >>
rect 215 373 216 374 
<< m1 >>
rect 217 373 218 374 
<< pdiffusion >>
rect 228 373 229 374 
<< pdiffusion >>
rect 229 373 230 374 
<< pdiffusion >>
rect 230 373 231 374 
<< pdiffusion >>
rect 231 373 232 374 
<< pdiffusion >>
rect 232 373 233 374 
<< pdiffusion >>
rect 233 373 234 374 
<< m1 >>
rect 244 373 245 374 
<< pdiffusion >>
rect 246 373 247 374 
<< pdiffusion >>
rect 247 373 248 374 
<< pdiffusion >>
rect 248 373 249 374 
<< pdiffusion >>
rect 249 373 250 374 
<< pdiffusion >>
rect 250 373 251 374 
<< pdiffusion >>
rect 251 373 252 374 
<< m1 >>
rect 253 373 254 374 
<< m1 >>
rect 255 373 256 374 
<< pdiffusion >>
rect 264 373 265 374 
<< pdiffusion >>
rect 265 373 266 374 
<< pdiffusion >>
rect 266 373 267 374 
<< pdiffusion >>
rect 267 373 268 374 
<< pdiffusion >>
rect 268 373 269 374 
<< pdiffusion >>
rect 269 373 270 374 
<< pdiffusion >>
rect 282 373 283 374 
<< pdiffusion >>
rect 283 373 284 374 
<< pdiffusion >>
rect 284 373 285 374 
<< pdiffusion >>
rect 285 373 286 374 
<< pdiffusion >>
rect 286 373 287 374 
<< pdiffusion >>
rect 287 373 288 374 
<< m1 >>
rect 289 373 290 374 
<< m1 >>
rect 293 373 294 374 
<< pdiffusion >>
rect 300 373 301 374 
<< pdiffusion >>
rect 301 373 302 374 
<< pdiffusion >>
rect 302 373 303 374 
<< pdiffusion >>
rect 303 373 304 374 
<< pdiffusion >>
rect 304 373 305 374 
<< pdiffusion >>
rect 305 373 306 374 
<< pdiffusion >>
rect 318 373 319 374 
<< pdiffusion >>
rect 319 373 320 374 
<< pdiffusion >>
rect 320 373 321 374 
<< pdiffusion >>
rect 321 373 322 374 
<< pdiffusion >>
rect 322 373 323 374 
<< pdiffusion >>
rect 323 373 324 374 
<< pdiffusion >>
rect 336 373 337 374 
<< pdiffusion >>
rect 337 373 338 374 
<< pdiffusion >>
rect 338 373 339 374 
<< pdiffusion >>
rect 339 373 340 374 
<< pdiffusion >>
rect 340 373 341 374 
<< pdiffusion >>
rect 341 373 342 374 
<< pdiffusion >>
rect 354 373 355 374 
<< pdiffusion >>
rect 355 373 356 374 
<< pdiffusion >>
rect 356 373 357 374 
<< pdiffusion >>
rect 357 373 358 374 
<< pdiffusion >>
rect 358 373 359 374 
<< pdiffusion >>
rect 359 373 360 374 
<< pdiffusion >>
rect 372 373 373 374 
<< pdiffusion >>
rect 373 373 374 374 
<< pdiffusion >>
rect 374 373 375 374 
<< pdiffusion >>
rect 375 373 376 374 
<< pdiffusion >>
rect 376 373 377 374 
<< pdiffusion >>
rect 377 373 378 374 
<< m1 >>
rect 379 373 380 374 
<< pdiffusion >>
rect 390 373 391 374 
<< pdiffusion >>
rect 391 373 392 374 
<< pdiffusion >>
rect 392 373 393 374 
<< pdiffusion >>
rect 393 373 394 374 
<< pdiffusion >>
rect 394 373 395 374 
<< pdiffusion >>
rect 395 373 396 374 
<< pdiffusion >>
rect 408 373 409 374 
<< pdiffusion >>
rect 409 373 410 374 
<< pdiffusion >>
rect 410 373 411 374 
<< pdiffusion >>
rect 411 373 412 374 
<< pdiffusion >>
rect 412 373 413 374 
<< pdiffusion >>
rect 413 373 414 374 
<< m1 >>
rect 415 373 416 374 
<< pdiffusion >>
rect 426 373 427 374 
<< pdiffusion >>
rect 427 373 428 374 
<< pdiffusion >>
rect 428 373 429 374 
<< pdiffusion >>
rect 429 373 430 374 
<< pdiffusion >>
rect 430 373 431 374 
<< pdiffusion >>
rect 431 373 432 374 
<< pdiffusion >>
rect 444 373 445 374 
<< pdiffusion >>
rect 445 373 446 374 
<< pdiffusion >>
rect 446 373 447 374 
<< pdiffusion >>
rect 447 373 448 374 
<< pdiffusion >>
rect 448 373 449 374 
<< pdiffusion >>
rect 449 373 450 374 
<< pdiffusion >>
rect 12 374 13 375 
<< pdiffusion >>
rect 13 374 14 375 
<< pdiffusion >>
rect 14 374 15 375 
<< pdiffusion >>
rect 15 374 16 375 
<< pdiffusion >>
rect 16 374 17 375 
<< pdiffusion >>
rect 17 374 18 375 
<< pdiffusion >>
rect 30 374 31 375 
<< pdiffusion >>
rect 31 374 32 375 
<< pdiffusion >>
rect 32 374 33 375 
<< pdiffusion >>
rect 33 374 34 375 
<< pdiffusion >>
rect 34 374 35 375 
<< pdiffusion >>
rect 35 374 36 375 
<< pdiffusion >>
rect 48 374 49 375 
<< pdiffusion >>
rect 49 374 50 375 
<< pdiffusion >>
rect 50 374 51 375 
<< pdiffusion >>
rect 51 374 52 375 
<< pdiffusion >>
rect 52 374 53 375 
<< pdiffusion >>
rect 53 374 54 375 
<< pdiffusion >>
rect 66 374 67 375 
<< pdiffusion >>
rect 67 374 68 375 
<< pdiffusion >>
rect 68 374 69 375 
<< pdiffusion >>
rect 69 374 70 375 
<< pdiffusion >>
rect 70 374 71 375 
<< pdiffusion >>
rect 71 374 72 375 
<< m1 >>
rect 82 374 83 375 
<< pdiffusion >>
rect 84 374 85 375 
<< pdiffusion >>
rect 85 374 86 375 
<< pdiffusion >>
rect 86 374 87 375 
<< pdiffusion >>
rect 87 374 88 375 
<< pdiffusion >>
rect 88 374 89 375 
<< pdiffusion >>
rect 89 374 90 375 
<< m1 >>
rect 100 374 101 375 
<< pdiffusion >>
rect 102 374 103 375 
<< pdiffusion >>
rect 103 374 104 375 
<< pdiffusion >>
rect 104 374 105 375 
<< pdiffusion >>
rect 105 374 106 375 
<< pdiffusion >>
rect 106 374 107 375 
<< pdiffusion >>
rect 107 374 108 375 
<< pdiffusion >>
rect 120 374 121 375 
<< pdiffusion >>
rect 121 374 122 375 
<< pdiffusion >>
rect 122 374 123 375 
<< pdiffusion >>
rect 123 374 124 375 
<< pdiffusion >>
rect 124 374 125 375 
<< pdiffusion >>
rect 125 374 126 375 
<< m1 >>
rect 127 374 128 375 
<< pdiffusion >>
rect 138 374 139 375 
<< pdiffusion >>
rect 139 374 140 375 
<< pdiffusion >>
rect 140 374 141 375 
<< pdiffusion >>
rect 141 374 142 375 
<< pdiffusion >>
rect 142 374 143 375 
<< pdiffusion >>
rect 143 374 144 375 
<< m1 >>
rect 145 374 146 375 
<< pdiffusion >>
rect 156 374 157 375 
<< pdiffusion >>
rect 157 374 158 375 
<< pdiffusion >>
rect 158 374 159 375 
<< pdiffusion >>
rect 159 374 160 375 
<< pdiffusion >>
rect 160 374 161 375 
<< pdiffusion >>
rect 161 374 162 375 
<< m1 >>
rect 163 374 164 375 
<< m2 >>
rect 164 374 165 375 
<< pdiffusion >>
rect 174 374 175 375 
<< pdiffusion >>
rect 175 374 176 375 
<< pdiffusion >>
rect 176 374 177 375 
<< pdiffusion >>
rect 177 374 178 375 
<< pdiffusion >>
rect 178 374 179 375 
<< pdiffusion >>
rect 179 374 180 375 
<< pdiffusion >>
rect 210 374 211 375 
<< pdiffusion >>
rect 211 374 212 375 
<< pdiffusion >>
rect 212 374 213 375 
<< pdiffusion >>
rect 213 374 214 375 
<< pdiffusion >>
rect 214 374 215 375 
<< pdiffusion >>
rect 215 374 216 375 
<< m1 >>
rect 217 374 218 375 
<< pdiffusion >>
rect 228 374 229 375 
<< pdiffusion >>
rect 229 374 230 375 
<< pdiffusion >>
rect 230 374 231 375 
<< pdiffusion >>
rect 231 374 232 375 
<< pdiffusion >>
rect 232 374 233 375 
<< pdiffusion >>
rect 233 374 234 375 
<< m1 >>
rect 244 374 245 375 
<< pdiffusion >>
rect 246 374 247 375 
<< pdiffusion >>
rect 247 374 248 375 
<< pdiffusion >>
rect 248 374 249 375 
<< pdiffusion >>
rect 249 374 250 375 
<< pdiffusion >>
rect 250 374 251 375 
<< pdiffusion >>
rect 251 374 252 375 
<< m1 >>
rect 253 374 254 375 
<< m1 >>
rect 255 374 256 375 
<< pdiffusion >>
rect 264 374 265 375 
<< pdiffusion >>
rect 265 374 266 375 
<< pdiffusion >>
rect 266 374 267 375 
<< pdiffusion >>
rect 267 374 268 375 
<< pdiffusion >>
rect 268 374 269 375 
<< pdiffusion >>
rect 269 374 270 375 
<< pdiffusion >>
rect 282 374 283 375 
<< pdiffusion >>
rect 283 374 284 375 
<< pdiffusion >>
rect 284 374 285 375 
<< pdiffusion >>
rect 285 374 286 375 
<< pdiffusion >>
rect 286 374 287 375 
<< pdiffusion >>
rect 287 374 288 375 
<< m1 >>
rect 289 374 290 375 
<< m1 >>
rect 293 374 294 375 
<< pdiffusion >>
rect 300 374 301 375 
<< pdiffusion >>
rect 301 374 302 375 
<< pdiffusion >>
rect 302 374 303 375 
<< pdiffusion >>
rect 303 374 304 375 
<< pdiffusion >>
rect 304 374 305 375 
<< pdiffusion >>
rect 305 374 306 375 
<< pdiffusion >>
rect 318 374 319 375 
<< pdiffusion >>
rect 319 374 320 375 
<< pdiffusion >>
rect 320 374 321 375 
<< pdiffusion >>
rect 321 374 322 375 
<< pdiffusion >>
rect 322 374 323 375 
<< pdiffusion >>
rect 323 374 324 375 
<< pdiffusion >>
rect 336 374 337 375 
<< pdiffusion >>
rect 337 374 338 375 
<< pdiffusion >>
rect 338 374 339 375 
<< pdiffusion >>
rect 339 374 340 375 
<< pdiffusion >>
rect 340 374 341 375 
<< pdiffusion >>
rect 341 374 342 375 
<< pdiffusion >>
rect 354 374 355 375 
<< pdiffusion >>
rect 355 374 356 375 
<< pdiffusion >>
rect 356 374 357 375 
<< pdiffusion >>
rect 357 374 358 375 
<< pdiffusion >>
rect 358 374 359 375 
<< pdiffusion >>
rect 359 374 360 375 
<< pdiffusion >>
rect 372 374 373 375 
<< pdiffusion >>
rect 373 374 374 375 
<< pdiffusion >>
rect 374 374 375 375 
<< pdiffusion >>
rect 375 374 376 375 
<< pdiffusion >>
rect 376 374 377 375 
<< pdiffusion >>
rect 377 374 378 375 
<< m1 >>
rect 379 374 380 375 
<< pdiffusion >>
rect 390 374 391 375 
<< pdiffusion >>
rect 391 374 392 375 
<< pdiffusion >>
rect 392 374 393 375 
<< pdiffusion >>
rect 393 374 394 375 
<< pdiffusion >>
rect 394 374 395 375 
<< pdiffusion >>
rect 395 374 396 375 
<< pdiffusion >>
rect 408 374 409 375 
<< pdiffusion >>
rect 409 374 410 375 
<< pdiffusion >>
rect 410 374 411 375 
<< pdiffusion >>
rect 411 374 412 375 
<< pdiffusion >>
rect 412 374 413 375 
<< pdiffusion >>
rect 413 374 414 375 
<< m1 >>
rect 415 374 416 375 
<< pdiffusion >>
rect 426 374 427 375 
<< pdiffusion >>
rect 427 374 428 375 
<< pdiffusion >>
rect 428 374 429 375 
<< pdiffusion >>
rect 429 374 430 375 
<< pdiffusion >>
rect 430 374 431 375 
<< pdiffusion >>
rect 431 374 432 375 
<< pdiffusion >>
rect 444 374 445 375 
<< pdiffusion >>
rect 445 374 446 375 
<< pdiffusion >>
rect 446 374 447 375 
<< pdiffusion >>
rect 447 374 448 375 
<< pdiffusion >>
rect 448 374 449 375 
<< pdiffusion >>
rect 449 374 450 375 
<< pdiffusion >>
rect 12 375 13 376 
<< pdiffusion >>
rect 13 375 14 376 
<< pdiffusion >>
rect 14 375 15 376 
<< pdiffusion >>
rect 15 375 16 376 
<< pdiffusion >>
rect 16 375 17 376 
<< pdiffusion >>
rect 17 375 18 376 
<< pdiffusion >>
rect 30 375 31 376 
<< pdiffusion >>
rect 31 375 32 376 
<< pdiffusion >>
rect 32 375 33 376 
<< pdiffusion >>
rect 33 375 34 376 
<< pdiffusion >>
rect 34 375 35 376 
<< pdiffusion >>
rect 35 375 36 376 
<< pdiffusion >>
rect 48 375 49 376 
<< pdiffusion >>
rect 49 375 50 376 
<< pdiffusion >>
rect 50 375 51 376 
<< pdiffusion >>
rect 51 375 52 376 
<< pdiffusion >>
rect 52 375 53 376 
<< pdiffusion >>
rect 53 375 54 376 
<< pdiffusion >>
rect 66 375 67 376 
<< pdiffusion >>
rect 67 375 68 376 
<< pdiffusion >>
rect 68 375 69 376 
<< pdiffusion >>
rect 69 375 70 376 
<< pdiffusion >>
rect 70 375 71 376 
<< pdiffusion >>
rect 71 375 72 376 
<< m1 >>
rect 82 375 83 376 
<< pdiffusion >>
rect 84 375 85 376 
<< pdiffusion >>
rect 85 375 86 376 
<< pdiffusion >>
rect 86 375 87 376 
<< pdiffusion >>
rect 87 375 88 376 
<< pdiffusion >>
rect 88 375 89 376 
<< pdiffusion >>
rect 89 375 90 376 
<< m1 >>
rect 100 375 101 376 
<< pdiffusion >>
rect 102 375 103 376 
<< pdiffusion >>
rect 103 375 104 376 
<< pdiffusion >>
rect 104 375 105 376 
<< pdiffusion >>
rect 105 375 106 376 
<< pdiffusion >>
rect 106 375 107 376 
<< pdiffusion >>
rect 107 375 108 376 
<< pdiffusion >>
rect 120 375 121 376 
<< pdiffusion >>
rect 121 375 122 376 
<< pdiffusion >>
rect 122 375 123 376 
<< pdiffusion >>
rect 123 375 124 376 
<< pdiffusion >>
rect 124 375 125 376 
<< pdiffusion >>
rect 125 375 126 376 
<< m1 >>
rect 127 375 128 376 
<< pdiffusion >>
rect 138 375 139 376 
<< pdiffusion >>
rect 139 375 140 376 
<< pdiffusion >>
rect 140 375 141 376 
<< pdiffusion >>
rect 141 375 142 376 
<< pdiffusion >>
rect 142 375 143 376 
<< pdiffusion >>
rect 143 375 144 376 
<< m1 >>
rect 145 375 146 376 
<< pdiffusion >>
rect 156 375 157 376 
<< pdiffusion >>
rect 157 375 158 376 
<< pdiffusion >>
rect 158 375 159 376 
<< pdiffusion >>
rect 159 375 160 376 
<< pdiffusion >>
rect 160 375 161 376 
<< pdiffusion >>
rect 161 375 162 376 
<< m1 >>
rect 163 375 164 376 
<< m2 >>
rect 164 375 165 376 
<< pdiffusion >>
rect 174 375 175 376 
<< pdiffusion >>
rect 175 375 176 376 
<< pdiffusion >>
rect 176 375 177 376 
<< pdiffusion >>
rect 177 375 178 376 
<< pdiffusion >>
rect 178 375 179 376 
<< pdiffusion >>
rect 179 375 180 376 
<< pdiffusion >>
rect 210 375 211 376 
<< pdiffusion >>
rect 211 375 212 376 
<< pdiffusion >>
rect 212 375 213 376 
<< pdiffusion >>
rect 213 375 214 376 
<< pdiffusion >>
rect 214 375 215 376 
<< pdiffusion >>
rect 215 375 216 376 
<< m1 >>
rect 217 375 218 376 
<< pdiffusion >>
rect 228 375 229 376 
<< pdiffusion >>
rect 229 375 230 376 
<< pdiffusion >>
rect 230 375 231 376 
<< pdiffusion >>
rect 231 375 232 376 
<< pdiffusion >>
rect 232 375 233 376 
<< pdiffusion >>
rect 233 375 234 376 
<< m1 >>
rect 244 375 245 376 
<< pdiffusion >>
rect 246 375 247 376 
<< pdiffusion >>
rect 247 375 248 376 
<< pdiffusion >>
rect 248 375 249 376 
<< pdiffusion >>
rect 249 375 250 376 
<< pdiffusion >>
rect 250 375 251 376 
<< pdiffusion >>
rect 251 375 252 376 
<< m1 >>
rect 253 375 254 376 
<< m1 >>
rect 255 375 256 376 
<< pdiffusion >>
rect 264 375 265 376 
<< pdiffusion >>
rect 265 375 266 376 
<< pdiffusion >>
rect 266 375 267 376 
<< pdiffusion >>
rect 267 375 268 376 
<< pdiffusion >>
rect 268 375 269 376 
<< pdiffusion >>
rect 269 375 270 376 
<< pdiffusion >>
rect 282 375 283 376 
<< pdiffusion >>
rect 283 375 284 376 
<< pdiffusion >>
rect 284 375 285 376 
<< pdiffusion >>
rect 285 375 286 376 
<< pdiffusion >>
rect 286 375 287 376 
<< pdiffusion >>
rect 287 375 288 376 
<< m1 >>
rect 289 375 290 376 
<< m1 >>
rect 293 375 294 376 
<< pdiffusion >>
rect 300 375 301 376 
<< pdiffusion >>
rect 301 375 302 376 
<< pdiffusion >>
rect 302 375 303 376 
<< pdiffusion >>
rect 303 375 304 376 
<< pdiffusion >>
rect 304 375 305 376 
<< pdiffusion >>
rect 305 375 306 376 
<< pdiffusion >>
rect 318 375 319 376 
<< pdiffusion >>
rect 319 375 320 376 
<< pdiffusion >>
rect 320 375 321 376 
<< pdiffusion >>
rect 321 375 322 376 
<< pdiffusion >>
rect 322 375 323 376 
<< pdiffusion >>
rect 323 375 324 376 
<< pdiffusion >>
rect 336 375 337 376 
<< pdiffusion >>
rect 337 375 338 376 
<< pdiffusion >>
rect 338 375 339 376 
<< pdiffusion >>
rect 339 375 340 376 
<< pdiffusion >>
rect 340 375 341 376 
<< pdiffusion >>
rect 341 375 342 376 
<< pdiffusion >>
rect 354 375 355 376 
<< pdiffusion >>
rect 355 375 356 376 
<< pdiffusion >>
rect 356 375 357 376 
<< pdiffusion >>
rect 357 375 358 376 
<< pdiffusion >>
rect 358 375 359 376 
<< pdiffusion >>
rect 359 375 360 376 
<< pdiffusion >>
rect 372 375 373 376 
<< pdiffusion >>
rect 373 375 374 376 
<< pdiffusion >>
rect 374 375 375 376 
<< pdiffusion >>
rect 375 375 376 376 
<< pdiffusion >>
rect 376 375 377 376 
<< pdiffusion >>
rect 377 375 378 376 
<< m1 >>
rect 379 375 380 376 
<< pdiffusion >>
rect 390 375 391 376 
<< pdiffusion >>
rect 391 375 392 376 
<< pdiffusion >>
rect 392 375 393 376 
<< pdiffusion >>
rect 393 375 394 376 
<< pdiffusion >>
rect 394 375 395 376 
<< pdiffusion >>
rect 395 375 396 376 
<< pdiffusion >>
rect 408 375 409 376 
<< pdiffusion >>
rect 409 375 410 376 
<< pdiffusion >>
rect 410 375 411 376 
<< pdiffusion >>
rect 411 375 412 376 
<< pdiffusion >>
rect 412 375 413 376 
<< pdiffusion >>
rect 413 375 414 376 
<< m1 >>
rect 415 375 416 376 
<< pdiffusion >>
rect 426 375 427 376 
<< pdiffusion >>
rect 427 375 428 376 
<< pdiffusion >>
rect 428 375 429 376 
<< pdiffusion >>
rect 429 375 430 376 
<< pdiffusion >>
rect 430 375 431 376 
<< pdiffusion >>
rect 431 375 432 376 
<< pdiffusion >>
rect 444 375 445 376 
<< pdiffusion >>
rect 445 375 446 376 
<< pdiffusion >>
rect 446 375 447 376 
<< pdiffusion >>
rect 447 375 448 376 
<< pdiffusion >>
rect 448 375 449 376 
<< pdiffusion >>
rect 449 375 450 376 
<< pdiffusion >>
rect 12 376 13 377 
<< pdiffusion >>
rect 13 376 14 377 
<< pdiffusion >>
rect 14 376 15 377 
<< pdiffusion >>
rect 15 376 16 377 
<< pdiffusion >>
rect 16 376 17 377 
<< pdiffusion >>
rect 17 376 18 377 
<< pdiffusion >>
rect 30 376 31 377 
<< pdiffusion >>
rect 31 376 32 377 
<< pdiffusion >>
rect 32 376 33 377 
<< pdiffusion >>
rect 33 376 34 377 
<< pdiffusion >>
rect 34 376 35 377 
<< pdiffusion >>
rect 35 376 36 377 
<< pdiffusion >>
rect 48 376 49 377 
<< pdiffusion >>
rect 49 376 50 377 
<< pdiffusion >>
rect 50 376 51 377 
<< pdiffusion >>
rect 51 376 52 377 
<< pdiffusion >>
rect 52 376 53 377 
<< pdiffusion >>
rect 53 376 54 377 
<< pdiffusion >>
rect 66 376 67 377 
<< pdiffusion >>
rect 67 376 68 377 
<< pdiffusion >>
rect 68 376 69 377 
<< pdiffusion >>
rect 69 376 70 377 
<< pdiffusion >>
rect 70 376 71 377 
<< pdiffusion >>
rect 71 376 72 377 
<< m1 >>
rect 82 376 83 377 
<< pdiffusion >>
rect 84 376 85 377 
<< pdiffusion >>
rect 85 376 86 377 
<< pdiffusion >>
rect 86 376 87 377 
<< pdiffusion >>
rect 87 376 88 377 
<< pdiffusion >>
rect 88 376 89 377 
<< pdiffusion >>
rect 89 376 90 377 
<< m1 >>
rect 100 376 101 377 
<< pdiffusion >>
rect 102 376 103 377 
<< pdiffusion >>
rect 103 376 104 377 
<< pdiffusion >>
rect 104 376 105 377 
<< pdiffusion >>
rect 105 376 106 377 
<< pdiffusion >>
rect 106 376 107 377 
<< pdiffusion >>
rect 107 376 108 377 
<< pdiffusion >>
rect 120 376 121 377 
<< pdiffusion >>
rect 121 376 122 377 
<< pdiffusion >>
rect 122 376 123 377 
<< pdiffusion >>
rect 123 376 124 377 
<< pdiffusion >>
rect 124 376 125 377 
<< pdiffusion >>
rect 125 376 126 377 
<< m1 >>
rect 127 376 128 377 
<< pdiffusion >>
rect 138 376 139 377 
<< pdiffusion >>
rect 139 376 140 377 
<< pdiffusion >>
rect 140 376 141 377 
<< pdiffusion >>
rect 141 376 142 377 
<< pdiffusion >>
rect 142 376 143 377 
<< pdiffusion >>
rect 143 376 144 377 
<< m1 >>
rect 145 376 146 377 
<< pdiffusion >>
rect 156 376 157 377 
<< pdiffusion >>
rect 157 376 158 377 
<< pdiffusion >>
rect 158 376 159 377 
<< pdiffusion >>
rect 159 376 160 377 
<< pdiffusion >>
rect 160 376 161 377 
<< pdiffusion >>
rect 161 376 162 377 
<< m1 >>
rect 163 376 164 377 
<< m2 >>
rect 164 376 165 377 
<< pdiffusion >>
rect 174 376 175 377 
<< pdiffusion >>
rect 175 376 176 377 
<< pdiffusion >>
rect 176 376 177 377 
<< pdiffusion >>
rect 177 376 178 377 
<< pdiffusion >>
rect 178 376 179 377 
<< pdiffusion >>
rect 179 376 180 377 
<< pdiffusion >>
rect 210 376 211 377 
<< pdiffusion >>
rect 211 376 212 377 
<< pdiffusion >>
rect 212 376 213 377 
<< pdiffusion >>
rect 213 376 214 377 
<< pdiffusion >>
rect 214 376 215 377 
<< pdiffusion >>
rect 215 376 216 377 
<< m1 >>
rect 217 376 218 377 
<< pdiffusion >>
rect 228 376 229 377 
<< pdiffusion >>
rect 229 376 230 377 
<< pdiffusion >>
rect 230 376 231 377 
<< pdiffusion >>
rect 231 376 232 377 
<< pdiffusion >>
rect 232 376 233 377 
<< pdiffusion >>
rect 233 376 234 377 
<< m1 >>
rect 244 376 245 377 
<< pdiffusion >>
rect 246 376 247 377 
<< pdiffusion >>
rect 247 376 248 377 
<< pdiffusion >>
rect 248 376 249 377 
<< pdiffusion >>
rect 249 376 250 377 
<< pdiffusion >>
rect 250 376 251 377 
<< pdiffusion >>
rect 251 376 252 377 
<< m1 >>
rect 253 376 254 377 
<< m1 >>
rect 255 376 256 377 
<< pdiffusion >>
rect 264 376 265 377 
<< pdiffusion >>
rect 265 376 266 377 
<< pdiffusion >>
rect 266 376 267 377 
<< pdiffusion >>
rect 267 376 268 377 
<< pdiffusion >>
rect 268 376 269 377 
<< pdiffusion >>
rect 269 376 270 377 
<< pdiffusion >>
rect 282 376 283 377 
<< pdiffusion >>
rect 283 376 284 377 
<< pdiffusion >>
rect 284 376 285 377 
<< pdiffusion >>
rect 285 376 286 377 
<< pdiffusion >>
rect 286 376 287 377 
<< pdiffusion >>
rect 287 376 288 377 
<< m1 >>
rect 289 376 290 377 
<< m1 >>
rect 293 376 294 377 
<< pdiffusion >>
rect 300 376 301 377 
<< pdiffusion >>
rect 301 376 302 377 
<< pdiffusion >>
rect 302 376 303 377 
<< pdiffusion >>
rect 303 376 304 377 
<< pdiffusion >>
rect 304 376 305 377 
<< pdiffusion >>
rect 305 376 306 377 
<< pdiffusion >>
rect 318 376 319 377 
<< pdiffusion >>
rect 319 376 320 377 
<< pdiffusion >>
rect 320 376 321 377 
<< pdiffusion >>
rect 321 376 322 377 
<< pdiffusion >>
rect 322 376 323 377 
<< pdiffusion >>
rect 323 376 324 377 
<< pdiffusion >>
rect 336 376 337 377 
<< pdiffusion >>
rect 337 376 338 377 
<< pdiffusion >>
rect 338 376 339 377 
<< pdiffusion >>
rect 339 376 340 377 
<< pdiffusion >>
rect 340 376 341 377 
<< pdiffusion >>
rect 341 376 342 377 
<< pdiffusion >>
rect 354 376 355 377 
<< pdiffusion >>
rect 355 376 356 377 
<< pdiffusion >>
rect 356 376 357 377 
<< pdiffusion >>
rect 357 376 358 377 
<< pdiffusion >>
rect 358 376 359 377 
<< pdiffusion >>
rect 359 376 360 377 
<< pdiffusion >>
rect 372 376 373 377 
<< pdiffusion >>
rect 373 376 374 377 
<< pdiffusion >>
rect 374 376 375 377 
<< pdiffusion >>
rect 375 376 376 377 
<< pdiffusion >>
rect 376 376 377 377 
<< pdiffusion >>
rect 377 376 378 377 
<< m1 >>
rect 379 376 380 377 
<< pdiffusion >>
rect 390 376 391 377 
<< pdiffusion >>
rect 391 376 392 377 
<< pdiffusion >>
rect 392 376 393 377 
<< pdiffusion >>
rect 393 376 394 377 
<< pdiffusion >>
rect 394 376 395 377 
<< pdiffusion >>
rect 395 376 396 377 
<< pdiffusion >>
rect 408 376 409 377 
<< pdiffusion >>
rect 409 376 410 377 
<< pdiffusion >>
rect 410 376 411 377 
<< pdiffusion >>
rect 411 376 412 377 
<< pdiffusion >>
rect 412 376 413 377 
<< pdiffusion >>
rect 413 376 414 377 
<< m1 >>
rect 415 376 416 377 
<< pdiffusion >>
rect 426 376 427 377 
<< pdiffusion >>
rect 427 376 428 377 
<< pdiffusion >>
rect 428 376 429 377 
<< pdiffusion >>
rect 429 376 430 377 
<< pdiffusion >>
rect 430 376 431 377 
<< pdiffusion >>
rect 431 376 432 377 
<< pdiffusion >>
rect 444 376 445 377 
<< pdiffusion >>
rect 445 376 446 377 
<< pdiffusion >>
rect 446 376 447 377 
<< pdiffusion >>
rect 447 376 448 377 
<< pdiffusion >>
rect 448 376 449 377 
<< pdiffusion >>
rect 449 376 450 377 
<< pdiffusion >>
rect 12 377 13 378 
<< m1 >>
rect 13 377 14 378 
<< pdiffusion >>
rect 13 377 14 378 
<< pdiffusion >>
rect 14 377 15 378 
<< pdiffusion >>
rect 15 377 16 378 
<< pdiffusion >>
rect 16 377 17 378 
<< pdiffusion >>
rect 17 377 18 378 
<< pdiffusion >>
rect 30 377 31 378 
<< pdiffusion >>
rect 31 377 32 378 
<< pdiffusion >>
rect 32 377 33 378 
<< pdiffusion >>
rect 33 377 34 378 
<< m1 >>
rect 34 377 35 378 
<< pdiffusion >>
rect 34 377 35 378 
<< pdiffusion >>
rect 35 377 36 378 
<< pdiffusion >>
rect 48 377 49 378 
<< pdiffusion >>
rect 49 377 50 378 
<< pdiffusion >>
rect 50 377 51 378 
<< pdiffusion >>
rect 51 377 52 378 
<< m1 >>
rect 52 377 53 378 
<< pdiffusion >>
rect 52 377 53 378 
<< pdiffusion >>
rect 53 377 54 378 
<< pdiffusion >>
rect 66 377 67 378 
<< pdiffusion >>
rect 67 377 68 378 
<< pdiffusion >>
rect 68 377 69 378 
<< pdiffusion >>
rect 69 377 70 378 
<< pdiffusion >>
rect 70 377 71 378 
<< pdiffusion >>
rect 71 377 72 378 
<< m1 >>
rect 82 377 83 378 
<< pdiffusion >>
rect 84 377 85 378 
<< m1 >>
rect 85 377 86 378 
<< pdiffusion >>
rect 85 377 86 378 
<< pdiffusion >>
rect 86 377 87 378 
<< pdiffusion >>
rect 87 377 88 378 
<< pdiffusion >>
rect 88 377 89 378 
<< pdiffusion >>
rect 89 377 90 378 
<< m1 >>
rect 100 377 101 378 
<< pdiffusion >>
rect 102 377 103 378 
<< pdiffusion >>
rect 103 377 104 378 
<< pdiffusion >>
rect 104 377 105 378 
<< pdiffusion >>
rect 105 377 106 378 
<< pdiffusion >>
rect 106 377 107 378 
<< pdiffusion >>
rect 107 377 108 378 
<< pdiffusion >>
rect 120 377 121 378 
<< pdiffusion >>
rect 121 377 122 378 
<< pdiffusion >>
rect 122 377 123 378 
<< pdiffusion >>
rect 123 377 124 378 
<< pdiffusion >>
rect 124 377 125 378 
<< pdiffusion >>
rect 125 377 126 378 
<< m1 >>
rect 127 377 128 378 
<< pdiffusion >>
rect 138 377 139 378 
<< pdiffusion >>
rect 139 377 140 378 
<< pdiffusion >>
rect 140 377 141 378 
<< pdiffusion >>
rect 141 377 142 378 
<< pdiffusion >>
rect 142 377 143 378 
<< pdiffusion >>
rect 143 377 144 378 
<< m1 >>
rect 145 377 146 378 
<< pdiffusion >>
rect 156 377 157 378 
<< pdiffusion >>
rect 157 377 158 378 
<< pdiffusion >>
rect 158 377 159 378 
<< pdiffusion >>
rect 159 377 160 378 
<< m1 >>
rect 160 377 161 378 
<< pdiffusion >>
rect 160 377 161 378 
<< pdiffusion >>
rect 161 377 162 378 
<< m1 >>
rect 163 377 164 378 
<< m2 >>
rect 164 377 165 378 
<< pdiffusion >>
rect 174 377 175 378 
<< pdiffusion >>
rect 175 377 176 378 
<< pdiffusion >>
rect 176 377 177 378 
<< pdiffusion >>
rect 177 377 178 378 
<< m1 >>
rect 178 377 179 378 
<< pdiffusion >>
rect 178 377 179 378 
<< pdiffusion >>
rect 179 377 180 378 
<< pdiffusion >>
rect 210 377 211 378 
<< m1 >>
rect 211 377 212 378 
<< pdiffusion >>
rect 211 377 212 378 
<< pdiffusion >>
rect 212 377 213 378 
<< pdiffusion >>
rect 213 377 214 378 
<< pdiffusion >>
rect 214 377 215 378 
<< pdiffusion >>
rect 215 377 216 378 
<< m1 >>
rect 217 377 218 378 
<< pdiffusion >>
rect 228 377 229 378 
<< m1 >>
rect 229 377 230 378 
<< pdiffusion >>
rect 229 377 230 378 
<< pdiffusion >>
rect 230 377 231 378 
<< pdiffusion >>
rect 231 377 232 378 
<< pdiffusion >>
rect 232 377 233 378 
<< pdiffusion >>
rect 233 377 234 378 
<< m1 >>
rect 244 377 245 378 
<< pdiffusion >>
rect 246 377 247 378 
<< m1 >>
rect 247 377 248 378 
<< pdiffusion >>
rect 247 377 248 378 
<< pdiffusion >>
rect 248 377 249 378 
<< pdiffusion >>
rect 249 377 250 378 
<< pdiffusion >>
rect 250 377 251 378 
<< pdiffusion >>
rect 251 377 252 378 
<< m1 >>
rect 253 377 254 378 
<< m1 >>
rect 255 377 256 378 
<< pdiffusion >>
rect 264 377 265 378 
<< pdiffusion >>
rect 265 377 266 378 
<< pdiffusion >>
rect 266 377 267 378 
<< pdiffusion >>
rect 267 377 268 378 
<< m1 >>
rect 268 377 269 378 
<< pdiffusion >>
rect 268 377 269 378 
<< pdiffusion >>
rect 269 377 270 378 
<< pdiffusion >>
rect 282 377 283 378 
<< pdiffusion >>
rect 283 377 284 378 
<< pdiffusion >>
rect 284 377 285 378 
<< pdiffusion >>
rect 285 377 286 378 
<< pdiffusion >>
rect 286 377 287 378 
<< pdiffusion >>
rect 287 377 288 378 
<< m1 >>
rect 289 377 290 378 
<< m1 >>
rect 293 377 294 378 
<< pdiffusion >>
rect 300 377 301 378 
<< pdiffusion >>
rect 301 377 302 378 
<< pdiffusion >>
rect 302 377 303 378 
<< pdiffusion >>
rect 303 377 304 378 
<< pdiffusion >>
rect 304 377 305 378 
<< pdiffusion >>
rect 305 377 306 378 
<< pdiffusion >>
rect 318 377 319 378 
<< pdiffusion >>
rect 319 377 320 378 
<< pdiffusion >>
rect 320 377 321 378 
<< pdiffusion >>
rect 321 377 322 378 
<< m1 >>
rect 322 377 323 378 
<< pdiffusion >>
rect 322 377 323 378 
<< pdiffusion >>
rect 323 377 324 378 
<< pdiffusion >>
rect 336 377 337 378 
<< pdiffusion >>
rect 337 377 338 378 
<< pdiffusion >>
rect 338 377 339 378 
<< pdiffusion >>
rect 339 377 340 378 
<< pdiffusion >>
rect 340 377 341 378 
<< pdiffusion >>
rect 341 377 342 378 
<< pdiffusion >>
rect 354 377 355 378 
<< pdiffusion >>
rect 355 377 356 378 
<< pdiffusion >>
rect 356 377 357 378 
<< pdiffusion >>
rect 357 377 358 378 
<< pdiffusion >>
rect 358 377 359 378 
<< pdiffusion >>
rect 359 377 360 378 
<< pdiffusion >>
rect 372 377 373 378 
<< pdiffusion >>
rect 373 377 374 378 
<< pdiffusion >>
rect 374 377 375 378 
<< pdiffusion >>
rect 375 377 376 378 
<< pdiffusion >>
rect 376 377 377 378 
<< pdiffusion >>
rect 377 377 378 378 
<< m1 >>
rect 379 377 380 378 
<< pdiffusion >>
rect 390 377 391 378 
<< pdiffusion >>
rect 391 377 392 378 
<< pdiffusion >>
rect 392 377 393 378 
<< pdiffusion >>
rect 393 377 394 378 
<< pdiffusion >>
rect 394 377 395 378 
<< pdiffusion >>
rect 395 377 396 378 
<< pdiffusion >>
rect 408 377 409 378 
<< pdiffusion >>
rect 409 377 410 378 
<< pdiffusion >>
rect 410 377 411 378 
<< pdiffusion >>
rect 411 377 412 378 
<< m1 >>
rect 412 377 413 378 
<< pdiffusion >>
rect 412 377 413 378 
<< pdiffusion >>
rect 413 377 414 378 
<< m1 >>
rect 415 377 416 378 
<< pdiffusion >>
rect 426 377 427 378 
<< pdiffusion >>
rect 427 377 428 378 
<< pdiffusion >>
rect 428 377 429 378 
<< pdiffusion >>
rect 429 377 430 378 
<< pdiffusion >>
rect 430 377 431 378 
<< pdiffusion >>
rect 431 377 432 378 
<< pdiffusion >>
rect 444 377 445 378 
<< pdiffusion >>
rect 445 377 446 378 
<< pdiffusion >>
rect 446 377 447 378 
<< pdiffusion >>
rect 447 377 448 378 
<< m1 >>
rect 448 377 449 378 
<< pdiffusion >>
rect 448 377 449 378 
<< pdiffusion >>
rect 449 377 450 378 
<< m1 >>
rect 13 378 14 379 
<< m1 >>
rect 34 378 35 379 
<< m1 >>
rect 52 378 53 379 
<< m1 >>
rect 82 378 83 379 
<< m1 >>
rect 85 378 86 379 
<< m1 >>
rect 100 378 101 379 
<< m1 >>
rect 127 378 128 379 
<< m1 >>
rect 145 378 146 379 
<< m1 >>
rect 160 378 161 379 
<< m1 >>
rect 163 378 164 379 
<< m2 >>
rect 164 378 165 379 
<< m1 >>
rect 178 378 179 379 
<< m1 >>
rect 211 378 212 379 
<< m1 >>
rect 217 378 218 379 
<< m1 >>
rect 229 378 230 379 
<< m1 >>
rect 244 378 245 379 
<< m1 >>
rect 247 378 248 379 
<< m1 >>
rect 253 378 254 379 
<< m1 >>
rect 255 378 256 379 
<< m1 >>
rect 268 378 269 379 
<< m1 >>
rect 289 378 290 379 
<< m1 >>
rect 293 378 294 379 
<< m1 >>
rect 322 378 323 379 
<< m1 >>
rect 379 378 380 379 
<< m1 >>
rect 412 378 413 379 
<< m1 >>
rect 415 378 416 379 
<< m1 >>
rect 448 378 449 379 
<< m1 >>
rect 13 379 14 380 
<< m1 >>
rect 34 379 35 380 
<< m1 >>
rect 52 379 53 380 
<< m1 >>
rect 82 379 83 380 
<< m1 >>
rect 85 379 86 380 
<< m1 >>
rect 100 379 101 380 
<< m1 >>
rect 127 379 128 380 
<< m1 >>
rect 145 379 146 380 
<< m1 >>
rect 160 379 161 380 
<< m1 >>
rect 163 379 164 380 
<< m2 >>
rect 164 379 165 380 
<< m1 >>
rect 178 379 179 380 
<< m1 >>
rect 211 379 212 380 
<< m1 >>
rect 217 379 218 380 
<< m1 >>
rect 229 379 230 380 
<< m1 >>
rect 244 379 245 380 
<< m1 >>
rect 247 379 248 380 
<< m1 >>
rect 253 379 254 380 
<< m1 >>
rect 255 379 256 380 
<< m1 >>
rect 268 379 269 380 
<< m1 >>
rect 289 379 290 380 
<< m1 >>
rect 293 379 294 380 
<< m1 >>
rect 322 379 323 380 
<< m1 >>
rect 379 379 380 380 
<< m1 >>
rect 412 379 413 380 
<< m1 >>
rect 413 379 414 380 
<< m1 >>
rect 414 379 415 380 
<< m1 >>
rect 415 379 416 380 
<< m1 >>
rect 448 379 449 380 
<< m1 >>
rect 13 380 14 381 
<< m1 >>
rect 34 380 35 381 
<< m1 >>
rect 52 380 53 381 
<< m1 >>
rect 82 380 83 381 
<< m2 >>
rect 82 380 83 381 
<< m2c >>
rect 82 380 83 381 
<< m1 >>
rect 82 380 83 381 
<< m2 >>
rect 82 380 83 381 
<< m1 >>
rect 85 380 86 381 
<< m1 >>
rect 86 380 87 381 
<< m1 >>
rect 87 380 88 381 
<< m1 >>
rect 88 380 89 381 
<< m1 >>
rect 89 380 90 381 
<< m1 >>
rect 90 380 91 381 
<< m1 >>
rect 91 380 92 381 
<< m1 >>
rect 92 380 93 381 
<< m1 >>
rect 93 380 94 381 
<< m1 >>
rect 94 380 95 381 
<< m1 >>
rect 95 380 96 381 
<< m1 >>
rect 96 380 97 381 
<< m1 >>
rect 97 380 98 381 
<< m1 >>
rect 98 380 99 381 
<< m1 >>
rect 99 380 100 381 
<< m1 >>
rect 100 380 101 381 
<< m1 >>
rect 127 380 128 381 
<< m2 >>
rect 127 380 128 381 
<< m2c >>
rect 127 380 128 381 
<< m1 >>
rect 127 380 128 381 
<< m2 >>
rect 127 380 128 381 
<< m1 >>
rect 145 380 146 381 
<< m2 >>
rect 145 380 146 381 
<< m2c >>
rect 145 380 146 381 
<< m1 >>
rect 145 380 146 381 
<< m2 >>
rect 145 380 146 381 
<< m1 >>
rect 158 380 159 381 
<< m2 >>
rect 158 380 159 381 
<< m2c >>
rect 158 380 159 381 
<< m1 >>
rect 158 380 159 381 
<< m2 >>
rect 158 380 159 381 
<< m2 >>
rect 159 380 160 381 
<< m1 >>
rect 160 380 161 381 
<< m2 >>
rect 160 380 161 381 
<< m2 >>
rect 161 380 162 381 
<< m2 >>
rect 162 380 163 381 
<< m1 >>
rect 163 380 164 381 
<< m2 >>
rect 163 380 164 381 
<< m2 >>
rect 164 380 165 381 
<< m1 >>
rect 178 380 179 381 
<< m1 >>
rect 211 380 212 381 
<< m1 >>
rect 212 380 213 381 
<< m1 >>
rect 213 380 214 381 
<< m1 >>
rect 214 380 215 381 
<< m1 >>
rect 215 380 216 381 
<< m2 >>
rect 215 380 216 381 
<< m2c >>
rect 215 380 216 381 
<< m1 >>
rect 215 380 216 381 
<< m2 >>
rect 215 380 216 381 
<< m2 >>
rect 216 380 217 381 
<< m1 >>
rect 217 380 218 381 
<< m2 >>
rect 217 380 218 381 
<< m2 >>
rect 218 380 219 381 
<< m1 >>
rect 219 380 220 381 
<< m2 >>
rect 219 380 220 381 
<< m2c >>
rect 219 380 220 381 
<< m1 >>
rect 219 380 220 381 
<< m2 >>
rect 219 380 220 381 
<< m1 >>
rect 220 380 221 381 
<< m1 >>
rect 221 380 222 381 
<< m1 >>
rect 222 380 223 381 
<< m1 >>
rect 223 380 224 381 
<< m1 >>
rect 224 380 225 381 
<< m1 >>
rect 225 380 226 381 
<< m1 >>
rect 226 380 227 381 
<< m1 >>
rect 227 380 228 381 
<< m1 >>
rect 228 380 229 381 
<< m1 >>
rect 229 380 230 381 
<< m1 >>
rect 244 380 245 381 
<< m1 >>
rect 247 380 248 381 
<< m1 >>
rect 248 380 249 381 
<< m1 >>
rect 249 380 250 381 
<< m1 >>
rect 250 380 251 381 
<< m1 >>
rect 251 380 252 381 
<< m2 >>
rect 251 380 252 381 
<< m2c >>
rect 251 380 252 381 
<< m1 >>
rect 251 380 252 381 
<< m2 >>
rect 251 380 252 381 
<< m2 >>
rect 252 380 253 381 
<< m1 >>
rect 253 380 254 381 
<< m2 >>
rect 253 380 254 381 
<< m2 >>
rect 254 380 255 381 
<< m1 >>
rect 255 380 256 381 
<< m2 >>
rect 255 380 256 381 
<< m2c >>
rect 255 380 256 381 
<< m1 >>
rect 255 380 256 381 
<< m2 >>
rect 255 380 256 381 
<< m1 >>
rect 268 380 269 381 
<< m1 >>
rect 289 380 290 381 
<< m1 >>
rect 293 380 294 381 
<< m1 >>
rect 322 380 323 381 
<< m1 >>
rect 379 380 380 381 
<< m1 >>
rect 448 380 449 381 
<< m1 >>
rect 13 381 14 382 
<< m1 >>
rect 34 381 35 382 
<< m1 >>
rect 52 381 53 382 
<< m2 >>
rect 82 381 83 382 
<< m2 >>
rect 127 381 128 382 
<< m2 >>
rect 145 381 146 382 
<< m1 >>
rect 158 381 159 382 
<< m1 >>
rect 160 381 161 382 
<< m1 >>
rect 163 381 164 382 
<< m1 >>
rect 178 381 179 382 
<< m1 >>
rect 217 381 218 382 
<< m1 >>
rect 244 381 245 382 
<< m1 >>
rect 253 381 254 382 
<< m1 >>
rect 268 381 269 382 
<< m1 >>
rect 289 381 290 382 
<< m1 >>
rect 293 381 294 382 
<< m1 >>
rect 322 381 323 382 
<< m1 >>
rect 379 381 380 382 
<< m1 >>
rect 448 381 449 382 
<< m1 >>
rect 13 382 14 383 
<< m1 >>
rect 14 382 15 383 
<< m1 >>
rect 15 382 16 383 
<< m1 >>
rect 16 382 17 383 
<< m1 >>
rect 17 382 18 383 
<< m1 >>
rect 18 382 19 383 
<< m1 >>
rect 19 382 20 383 
<< m1 >>
rect 20 382 21 383 
<< m1 >>
rect 21 382 22 383 
<< m1 >>
rect 22 382 23 383 
<< m1 >>
rect 23 382 24 383 
<< m1 >>
rect 24 382 25 383 
<< m1 >>
rect 25 382 26 383 
<< m1 >>
rect 26 382 27 383 
<< m1 >>
rect 27 382 28 383 
<< m1 >>
rect 28 382 29 383 
<< m1 >>
rect 29 382 30 383 
<< m1 >>
rect 30 382 31 383 
<< m1 >>
rect 31 382 32 383 
<< m1 >>
rect 32 382 33 383 
<< m1 >>
rect 33 382 34 383 
<< m1 >>
rect 34 382 35 383 
<< m1 >>
rect 52 382 53 383 
<< m1 >>
rect 67 382 68 383 
<< m1 >>
rect 68 382 69 383 
<< m1 >>
rect 69 382 70 383 
<< m1 >>
rect 70 382 71 383 
<< m1 >>
rect 71 382 72 383 
<< m1 >>
rect 72 382 73 383 
<< m1 >>
rect 73 382 74 383 
<< m1 >>
rect 74 382 75 383 
<< m1 >>
rect 75 382 76 383 
<< m1 >>
rect 76 382 77 383 
<< m1 >>
rect 77 382 78 383 
<< m1 >>
rect 78 382 79 383 
<< m1 >>
rect 79 382 80 383 
<< m1 >>
rect 80 382 81 383 
<< m1 >>
rect 81 382 82 383 
<< m1 >>
rect 82 382 83 383 
<< m2 >>
rect 82 382 83 383 
<< m1 >>
rect 83 382 84 383 
<< m1 >>
rect 84 382 85 383 
<< m1 >>
rect 85 382 86 383 
<< m1 >>
rect 86 382 87 383 
<< m1 >>
rect 87 382 88 383 
<< m1 >>
rect 88 382 89 383 
<< m1 >>
rect 89 382 90 383 
<< m1 >>
rect 90 382 91 383 
<< m1 >>
rect 91 382 92 383 
<< m1 >>
rect 92 382 93 383 
<< m1 >>
rect 93 382 94 383 
<< m1 >>
rect 94 382 95 383 
<< m1 >>
rect 95 382 96 383 
<< m1 >>
rect 96 382 97 383 
<< m1 >>
rect 97 382 98 383 
<< m1 >>
rect 98 382 99 383 
<< m1 >>
rect 99 382 100 383 
<< m1 >>
rect 100 382 101 383 
<< m1 >>
rect 101 382 102 383 
<< m1 >>
rect 102 382 103 383 
<< m1 >>
rect 103 382 104 383 
<< m1 >>
rect 104 382 105 383 
<< m1 >>
rect 105 382 106 383 
<< m1 >>
rect 106 382 107 383 
<< m1 >>
rect 107 382 108 383 
<< m1 >>
rect 108 382 109 383 
<< m1 >>
rect 109 382 110 383 
<< m1 >>
rect 110 382 111 383 
<< m1 >>
rect 111 382 112 383 
<< m1 >>
rect 112 382 113 383 
<< m1 >>
rect 113 382 114 383 
<< m1 >>
rect 114 382 115 383 
<< m1 >>
rect 115 382 116 383 
<< m1 >>
rect 116 382 117 383 
<< m1 >>
rect 117 382 118 383 
<< m1 >>
rect 118 382 119 383 
<< m1 >>
rect 119 382 120 383 
<< m1 >>
rect 120 382 121 383 
<< m1 >>
rect 121 382 122 383 
<< m1 >>
rect 122 382 123 383 
<< m1 >>
rect 123 382 124 383 
<< m1 >>
rect 124 382 125 383 
<< m1 >>
rect 125 382 126 383 
<< m1 >>
rect 126 382 127 383 
<< m1 >>
rect 127 382 128 383 
<< m2 >>
rect 127 382 128 383 
<< m1 >>
rect 128 382 129 383 
<< m1 >>
rect 129 382 130 383 
<< m1 >>
rect 130 382 131 383 
<< m1 >>
rect 131 382 132 383 
<< m1 >>
rect 132 382 133 383 
<< m1 >>
rect 133 382 134 383 
<< m1 >>
rect 134 382 135 383 
<< m1 >>
rect 135 382 136 383 
<< m1 >>
rect 136 382 137 383 
<< m1 >>
rect 137 382 138 383 
<< m1 >>
rect 138 382 139 383 
<< m1 >>
rect 139 382 140 383 
<< m1 >>
rect 140 382 141 383 
<< m1 >>
rect 141 382 142 383 
<< m1 >>
rect 142 382 143 383 
<< m1 >>
rect 143 382 144 383 
<< m1 >>
rect 144 382 145 383 
<< m1 >>
rect 145 382 146 383 
<< m2 >>
rect 145 382 146 383 
<< m1 >>
rect 146 382 147 383 
<< m1 >>
rect 147 382 148 383 
<< m1 >>
rect 148 382 149 383 
<< m1 >>
rect 149 382 150 383 
<< m1 >>
rect 150 382 151 383 
<< m1 >>
rect 151 382 152 383 
<< m1 >>
rect 152 382 153 383 
<< m1 >>
rect 153 382 154 383 
<< m1 >>
rect 154 382 155 383 
<< m1 >>
rect 155 382 156 383 
<< m1 >>
rect 156 382 157 383 
<< m1 >>
rect 157 382 158 383 
<< m1 >>
rect 158 382 159 383 
<< m1 >>
rect 160 382 161 383 
<< m1 >>
rect 163 382 164 383 
<< m1 >>
rect 164 382 165 383 
<< m1 >>
rect 165 382 166 383 
<< m1 >>
rect 166 382 167 383 
<< m1 >>
rect 167 382 168 383 
<< m1 >>
rect 168 382 169 383 
<< m1 >>
rect 169 382 170 383 
<< m1 >>
rect 170 382 171 383 
<< m1 >>
rect 171 382 172 383 
<< m1 >>
rect 172 382 173 383 
<< m1 >>
rect 173 382 174 383 
<< m1 >>
rect 174 382 175 383 
<< m1 >>
rect 175 382 176 383 
<< m1 >>
rect 176 382 177 383 
<< m1 >>
rect 177 382 178 383 
<< m1 >>
rect 178 382 179 383 
<< m1 >>
rect 217 382 218 383 
<< m1 >>
rect 244 382 245 383 
<< m1 >>
rect 253 382 254 383 
<< m1 >>
rect 254 382 255 383 
<< m1 >>
rect 255 382 256 383 
<< m1 >>
rect 256 382 257 383 
<< m1 >>
rect 257 382 258 383 
<< m1 >>
rect 258 382 259 383 
<< m1 >>
rect 259 382 260 383 
<< m1 >>
rect 260 382 261 383 
<< m1 >>
rect 261 382 262 383 
<< m1 >>
rect 262 382 263 383 
<< m1 >>
rect 263 382 264 383 
<< m1 >>
rect 264 382 265 383 
<< m1 >>
rect 265 382 266 383 
<< m1 >>
rect 266 382 267 383 
<< m1 >>
rect 267 382 268 383 
<< m1 >>
rect 268 382 269 383 
<< m1 >>
rect 289 382 290 383 
<< m1 >>
rect 293 382 294 383 
<< m1 >>
rect 294 382 295 383 
<< m1 >>
rect 295 382 296 383 
<< m1 >>
rect 296 382 297 383 
<< m1 >>
rect 297 382 298 383 
<< m1 >>
rect 298 382 299 383 
<< m1 >>
rect 299 382 300 383 
<< m1 >>
rect 300 382 301 383 
<< m1 >>
rect 301 382 302 383 
<< m1 >>
rect 302 382 303 383 
<< m1 >>
rect 303 382 304 383 
<< m1 >>
rect 304 382 305 383 
<< m1 >>
rect 305 382 306 383 
<< m1 >>
rect 306 382 307 383 
<< m1 >>
rect 307 382 308 383 
<< m1 >>
rect 308 382 309 383 
<< m1 >>
rect 309 382 310 383 
<< m1 >>
rect 310 382 311 383 
<< m1 >>
rect 311 382 312 383 
<< m1 >>
rect 312 382 313 383 
<< m1 >>
rect 313 382 314 383 
<< m1 >>
rect 314 382 315 383 
<< m1 >>
rect 315 382 316 383 
<< m1 >>
rect 316 382 317 383 
<< m1 >>
rect 317 382 318 383 
<< m1 >>
rect 318 382 319 383 
<< m1 >>
rect 319 382 320 383 
<< m1 >>
rect 320 382 321 383 
<< m1 >>
rect 321 382 322 383 
<< m1 >>
rect 322 382 323 383 
<< m1 >>
rect 379 382 380 383 
<< m1 >>
rect 380 382 381 383 
<< m1 >>
rect 381 382 382 383 
<< m1 >>
rect 382 382 383 383 
<< m1 >>
rect 383 382 384 383 
<< m1 >>
rect 384 382 385 383 
<< m1 >>
rect 385 382 386 383 
<< m1 >>
rect 386 382 387 383 
<< m1 >>
rect 387 382 388 383 
<< m1 >>
rect 388 382 389 383 
<< m1 >>
rect 389 382 390 383 
<< m1 >>
rect 390 382 391 383 
<< m1 >>
rect 391 382 392 383 
<< m1 >>
rect 392 382 393 383 
<< m1 >>
rect 393 382 394 383 
<< m1 >>
rect 394 382 395 383 
<< m1 >>
rect 395 382 396 383 
<< m1 >>
rect 396 382 397 383 
<< m1 >>
rect 397 382 398 383 
<< m1 >>
rect 398 382 399 383 
<< m1 >>
rect 399 382 400 383 
<< m1 >>
rect 400 382 401 383 
<< m1 >>
rect 401 382 402 383 
<< m1 >>
rect 402 382 403 383 
<< m1 >>
rect 403 382 404 383 
<< m1 >>
rect 404 382 405 383 
<< m1 >>
rect 405 382 406 383 
<< m1 >>
rect 406 382 407 383 
<< m1 >>
rect 407 382 408 383 
<< m1 >>
rect 408 382 409 383 
<< m1 >>
rect 409 382 410 383 
<< m1 >>
rect 410 382 411 383 
<< m1 >>
rect 411 382 412 383 
<< m1 >>
rect 412 382 413 383 
<< m1 >>
rect 413 382 414 383 
<< m1 >>
rect 414 382 415 383 
<< m1 >>
rect 415 382 416 383 
<< m1 >>
rect 416 382 417 383 
<< m1 >>
rect 417 382 418 383 
<< m1 >>
rect 418 382 419 383 
<< m1 >>
rect 419 382 420 383 
<< m1 >>
rect 420 382 421 383 
<< m1 >>
rect 421 382 422 383 
<< m1 >>
rect 422 382 423 383 
<< m1 >>
rect 423 382 424 383 
<< m1 >>
rect 424 382 425 383 
<< m1 >>
rect 425 382 426 383 
<< m1 >>
rect 426 382 427 383 
<< m1 >>
rect 427 382 428 383 
<< m1 >>
rect 428 382 429 383 
<< m1 >>
rect 429 382 430 383 
<< m1 >>
rect 430 382 431 383 
<< m1 >>
rect 431 382 432 383 
<< m1 >>
rect 432 382 433 383 
<< m1 >>
rect 433 382 434 383 
<< m1 >>
rect 434 382 435 383 
<< m1 >>
rect 435 382 436 383 
<< m1 >>
rect 436 382 437 383 
<< m1 >>
rect 437 382 438 383 
<< m1 >>
rect 438 382 439 383 
<< m1 >>
rect 439 382 440 383 
<< m1 >>
rect 440 382 441 383 
<< m1 >>
rect 441 382 442 383 
<< m1 >>
rect 442 382 443 383 
<< m1 >>
rect 443 382 444 383 
<< m1 >>
rect 444 382 445 383 
<< m1 >>
rect 445 382 446 383 
<< m1 >>
rect 446 382 447 383 
<< m1 >>
rect 447 382 448 383 
<< m1 >>
rect 448 382 449 383 
<< m1 >>
rect 52 383 53 384 
<< m1 >>
rect 67 383 68 384 
<< m2 >>
rect 82 383 83 384 
<< m2 >>
rect 127 383 128 384 
<< m2 >>
rect 145 383 146 384 
<< m1 >>
rect 160 383 161 384 
<< m1 >>
rect 217 383 218 384 
<< m1 >>
rect 244 383 245 384 
<< m1 >>
rect 289 383 290 384 
<< m1 >>
rect 52 384 53 385 
<< m1 >>
rect 67 384 68 385 
<< m1 >>
rect 82 384 83 385 
<< m2 >>
rect 82 384 83 385 
<< m2c >>
rect 82 384 83 385 
<< m1 >>
rect 82 384 83 385 
<< m2 >>
rect 82 384 83 385 
<< m1 >>
rect 127 384 128 385 
<< m2 >>
rect 127 384 128 385 
<< m2c >>
rect 127 384 128 385 
<< m1 >>
rect 127 384 128 385 
<< m2 >>
rect 127 384 128 385 
<< m1 >>
rect 145 384 146 385 
<< m2 >>
rect 145 384 146 385 
<< m2c >>
rect 145 384 146 385 
<< m1 >>
rect 145 384 146 385 
<< m2 >>
rect 145 384 146 385 
<< m1 >>
rect 160 384 161 385 
<< m1 >>
rect 217 384 218 385 
<< m1 >>
rect 244 384 245 385 
<< m1 >>
rect 289 384 290 385 
<< m1 >>
rect 52 385 53 386 
<< m1 >>
rect 67 385 68 386 
<< m1 >>
rect 82 385 83 386 
<< m1 >>
rect 127 385 128 386 
<< m1 >>
rect 145 385 146 386 
<< m1 >>
rect 160 385 161 386 
<< m2 >>
rect 160 385 161 386 
<< m2 >>
rect 161 385 162 386 
<< m1 >>
rect 162 385 163 386 
<< m2 >>
rect 162 385 163 386 
<< m2c >>
rect 162 385 163 386 
<< m1 >>
rect 162 385 163 386 
<< m2 >>
rect 162 385 163 386 
<< m1 >>
rect 163 385 164 386 
<< m1 >>
rect 164 385 165 386 
<< m1 >>
rect 165 385 166 386 
<< m1 >>
rect 166 385 167 386 
<< m1 >>
rect 167 385 168 386 
<< m1 >>
rect 168 385 169 386 
<< m1 >>
rect 169 385 170 386 
<< m1 >>
rect 170 385 171 386 
<< m1 >>
rect 171 385 172 386 
<< m1 >>
rect 172 385 173 386 
<< m1 >>
rect 173 385 174 386 
<< m1 >>
rect 174 385 175 386 
<< m1 >>
rect 175 385 176 386 
<< m1 >>
rect 176 385 177 386 
<< m1 >>
rect 177 385 178 386 
<< m1 >>
rect 178 385 179 386 
<< m1 >>
rect 179 385 180 386 
<< m1 >>
rect 180 385 181 386 
<< m1 >>
rect 181 385 182 386 
<< m1 >>
rect 182 385 183 386 
<< m1 >>
rect 183 385 184 386 
<< m1 >>
rect 184 385 185 386 
<< m1 >>
rect 185 385 186 386 
<< m1 >>
rect 186 385 187 386 
<< m1 >>
rect 187 385 188 386 
<< m1 >>
rect 188 385 189 386 
<< m1 >>
rect 189 385 190 386 
<< m1 >>
rect 190 385 191 386 
<< m1 >>
rect 191 385 192 386 
<< m1 >>
rect 192 385 193 386 
<< m1 >>
rect 193 385 194 386 
<< m1 >>
rect 194 385 195 386 
<< m1 >>
rect 195 385 196 386 
<< m1 >>
rect 196 385 197 386 
<< m1 >>
rect 197 385 198 386 
<< m1 >>
rect 198 385 199 386 
<< m1 >>
rect 199 385 200 386 
<< m1 >>
rect 200 385 201 386 
<< m1 >>
rect 201 385 202 386 
<< m1 >>
rect 202 385 203 386 
<< m1 >>
rect 203 385 204 386 
<< m1 >>
rect 204 385 205 386 
<< m1 >>
rect 205 385 206 386 
<< m1 >>
rect 206 385 207 386 
<< m1 >>
rect 207 385 208 386 
<< m1 >>
rect 208 385 209 386 
<< m1 >>
rect 209 385 210 386 
<< m1 >>
rect 210 385 211 386 
<< m1 >>
rect 211 385 212 386 
<< m1 >>
rect 212 385 213 386 
<< m1 >>
rect 213 385 214 386 
<< m1 >>
rect 214 385 215 386 
<< m1 >>
rect 215 385 216 386 
<< m1 >>
rect 216 385 217 386 
<< m1 >>
rect 217 385 218 386 
<< m1 >>
rect 244 385 245 386 
<< m1 >>
rect 245 385 246 386 
<< m1 >>
rect 246 385 247 386 
<< m1 >>
rect 247 385 248 386 
<< m1 >>
rect 248 385 249 386 
<< m1 >>
rect 249 385 250 386 
<< m1 >>
rect 250 385 251 386 
<< m1 >>
rect 251 385 252 386 
<< m1 >>
rect 252 385 253 386 
<< m1 >>
rect 253 385 254 386 
<< m1 >>
rect 254 385 255 386 
<< m1 >>
rect 255 385 256 386 
<< m1 >>
rect 256 385 257 386 
<< m1 >>
rect 257 385 258 386 
<< m1 >>
rect 258 385 259 386 
<< m1 >>
rect 259 385 260 386 
<< m1 >>
rect 260 385 261 386 
<< m1 >>
rect 261 385 262 386 
<< m1 >>
rect 262 385 263 386 
<< m1 >>
rect 263 385 264 386 
<< m1 >>
rect 264 385 265 386 
<< m1 >>
rect 265 385 266 386 
<< m1 >>
rect 266 385 267 386 
<< m1 >>
rect 267 385 268 386 
<< m1 >>
rect 268 385 269 386 
<< m1 >>
rect 269 385 270 386 
<< m1 >>
rect 270 385 271 386 
<< m1 >>
rect 271 385 272 386 
<< m1 >>
rect 272 385 273 386 
<< m1 >>
rect 273 385 274 386 
<< m1 >>
rect 274 385 275 386 
<< m1 >>
rect 275 385 276 386 
<< m1 >>
rect 276 385 277 386 
<< m1 >>
rect 277 385 278 386 
<< m1 >>
rect 278 385 279 386 
<< m1 >>
rect 279 385 280 386 
<< m1 >>
rect 280 385 281 386 
<< m1 >>
rect 281 385 282 386 
<< m1 >>
rect 282 385 283 386 
<< m1 >>
rect 283 385 284 386 
<< m1 >>
rect 284 385 285 386 
<< m1 >>
rect 285 385 286 386 
<< m1 >>
rect 286 385 287 386 
<< m1 >>
rect 287 385 288 386 
<< m1 >>
rect 289 385 290 386 
<< m1 >>
rect 52 386 53 387 
<< m1 >>
rect 67 386 68 387 
<< m1 >>
rect 82 386 83 387 
<< m1 >>
rect 127 386 128 387 
<< m1 >>
rect 145 386 146 387 
<< m1 >>
rect 160 386 161 387 
<< m2 >>
rect 160 386 161 387 
<< m1 >>
rect 287 386 288 387 
<< m1 >>
rect 289 386 290 387 
<< m1 >>
rect 52 387 53 388 
<< m1 >>
rect 53 387 54 388 
<< m1 >>
rect 54 387 55 388 
<< m1 >>
rect 55 387 56 388 
<< m1 >>
rect 56 387 57 388 
<< m1 >>
rect 57 387 58 388 
<< m1 >>
rect 58 387 59 388 
<< m1 >>
rect 59 387 60 388 
<< m1 >>
rect 60 387 61 388 
<< m1 >>
rect 61 387 62 388 
<< m1 >>
rect 62 387 63 388 
<< m1 >>
rect 63 387 64 388 
<< m1 >>
rect 64 387 65 388 
<< m1 >>
rect 67 387 68 388 
<< m1 >>
rect 82 387 83 388 
<< m1 >>
rect 103 387 104 388 
<< m1 >>
rect 104 387 105 388 
<< m1 >>
rect 105 387 106 388 
<< m1 >>
rect 106 387 107 388 
<< m1 >>
rect 107 387 108 388 
<< m1 >>
rect 108 387 109 388 
<< m1 >>
rect 109 387 110 388 
<< m1 >>
rect 127 387 128 388 
<< m1 >>
rect 145 387 146 388 
<< m1 >>
rect 160 387 161 388 
<< m2 >>
rect 160 387 161 388 
<< m1 >>
rect 161 387 162 388 
<< m1 >>
rect 162 387 163 388 
<< m1 >>
rect 163 387 164 388 
<< m1 >>
rect 164 387 165 388 
<< m1 >>
rect 165 387 166 388 
<< m1 >>
rect 166 387 167 388 
<< m1 >>
rect 167 387 168 388 
<< m1 >>
rect 168 387 169 388 
<< m1 >>
rect 169 387 170 388 
<< m1 >>
rect 170 387 171 388 
<< m1 >>
rect 171 387 172 388 
<< m1 >>
rect 172 387 173 388 
<< m1 >>
rect 287 387 288 388 
<< m1 >>
rect 289 387 290 388 
<< m1 >>
rect 64 388 65 389 
<< m1 >>
rect 67 388 68 389 
<< m1 >>
rect 82 388 83 389 
<< m1 >>
rect 103 388 104 389 
<< m1 >>
rect 109 388 110 389 
<< m1 >>
rect 127 388 128 389 
<< m1 >>
rect 145 388 146 389 
<< m2 >>
rect 160 388 161 389 
<< m1 >>
rect 172 388 173 389 
<< m1 >>
rect 287 388 288 389 
<< m2 >>
rect 287 388 288 389 
<< m2c >>
rect 287 388 288 389 
<< m1 >>
rect 287 388 288 389 
<< m2 >>
rect 287 388 288 389 
<< m2 >>
rect 288 388 289 389 
<< m1 >>
rect 289 388 290 389 
<< m2 >>
rect 289 388 290 389 
<< m2 >>
rect 290 388 291 389 
<< m1 >>
rect 64 389 65 390 
<< m1 >>
rect 67 389 68 390 
<< m1 >>
rect 82 389 83 390 
<< m1 >>
rect 103 389 104 390 
<< m1 >>
rect 109 389 110 390 
<< m1 >>
rect 127 389 128 390 
<< m1 >>
rect 145 389 146 390 
<< m1 >>
rect 160 389 161 390 
<< m2 >>
rect 160 389 161 390 
<< m1 >>
rect 172 389 173 390 
<< m1 >>
rect 289 389 290 390 
<< m2 >>
rect 290 389 291 390 
<< pdiffusion >>
rect 12 390 13 391 
<< pdiffusion >>
rect 13 390 14 391 
<< pdiffusion >>
rect 14 390 15 391 
<< pdiffusion >>
rect 15 390 16 391 
<< pdiffusion >>
rect 16 390 17 391 
<< pdiffusion >>
rect 17 390 18 391 
<< pdiffusion >>
rect 30 390 31 391 
<< pdiffusion >>
rect 31 390 32 391 
<< pdiffusion >>
rect 32 390 33 391 
<< pdiffusion >>
rect 33 390 34 391 
<< pdiffusion >>
rect 34 390 35 391 
<< pdiffusion >>
rect 35 390 36 391 
<< pdiffusion >>
rect 48 390 49 391 
<< pdiffusion >>
rect 49 390 50 391 
<< pdiffusion >>
rect 50 390 51 391 
<< pdiffusion >>
rect 51 390 52 391 
<< pdiffusion >>
rect 52 390 53 391 
<< pdiffusion >>
rect 53 390 54 391 
<< m1 >>
rect 64 390 65 391 
<< pdiffusion >>
rect 66 390 67 391 
<< m1 >>
rect 67 390 68 391 
<< pdiffusion >>
rect 67 390 68 391 
<< pdiffusion >>
rect 68 390 69 391 
<< pdiffusion >>
rect 69 390 70 391 
<< pdiffusion >>
rect 70 390 71 391 
<< pdiffusion >>
rect 71 390 72 391 
<< m1 >>
rect 82 390 83 391 
<< pdiffusion >>
rect 84 390 85 391 
<< pdiffusion >>
rect 85 390 86 391 
<< pdiffusion >>
rect 86 390 87 391 
<< pdiffusion >>
rect 87 390 88 391 
<< pdiffusion >>
rect 88 390 89 391 
<< pdiffusion >>
rect 89 390 90 391 
<< pdiffusion >>
rect 102 390 103 391 
<< m1 >>
rect 103 390 104 391 
<< pdiffusion >>
rect 103 390 104 391 
<< pdiffusion >>
rect 104 390 105 391 
<< pdiffusion >>
rect 105 390 106 391 
<< pdiffusion >>
rect 106 390 107 391 
<< pdiffusion >>
rect 107 390 108 391 
<< m1 >>
rect 109 390 110 391 
<< pdiffusion >>
rect 120 390 121 391 
<< pdiffusion >>
rect 121 390 122 391 
<< pdiffusion >>
rect 122 390 123 391 
<< pdiffusion >>
rect 123 390 124 391 
<< pdiffusion >>
rect 124 390 125 391 
<< pdiffusion >>
rect 125 390 126 391 
<< m1 >>
rect 127 390 128 391 
<< pdiffusion >>
rect 138 390 139 391 
<< pdiffusion >>
rect 139 390 140 391 
<< pdiffusion >>
rect 140 390 141 391 
<< pdiffusion >>
rect 141 390 142 391 
<< pdiffusion >>
rect 142 390 143 391 
<< pdiffusion >>
rect 143 390 144 391 
<< m1 >>
rect 145 390 146 391 
<< pdiffusion >>
rect 156 390 157 391 
<< pdiffusion >>
rect 157 390 158 391 
<< pdiffusion >>
rect 158 390 159 391 
<< m1 >>
rect 159 390 160 391 
<< m2 >>
rect 159 390 160 391 
<< m2c >>
rect 159 390 160 391 
<< m1 >>
rect 159 390 160 391 
<< m2 >>
rect 159 390 160 391 
<< pdiffusion >>
rect 159 390 160 391 
<< m1 >>
rect 160 390 161 391 
<< pdiffusion >>
rect 160 390 161 391 
<< pdiffusion >>
rect 161 390 162 391 
<< m1 >>
rect 172 390 173 391 
<< pdiffusion >>
rect 174 390 175 391 
<< pdiffusion >>
rect 175 390 176 391 
<< pdiffusion >>
rect 176 390 177 391 
<< pdiffusion >>
rect 177 390 178 391 
<< pdiffusion >>
rect 178 390 179 391 
<< pdiffusion >>
rect 179 390 180 391 
<< pdiffusion >>
rect 192 390 193 391 
<< pdiffusion >>
rect 193 390 194 391 
<< pdiffusion >>
rect 194 390 195 391 
<< pdiffusion >>
rect 195 390 196 391 
<< pdiffusion >>
rect 196 390 197 391 
<< pdiffusion >>
rect 197 390 198 391 
<< pdiffusion >>
rect 210 390 211 391 
<< pdiffusion >>
rect 211 390 212 391 
<< pdiffusion >>
rect 212 390 213 391 
<< pdiffusion >>
rect 213 390 214 391 
<< pdiffusion >>
rect 214 390 215 391 
<< pdiffusion >>
rect 215 390 216 391 
<< pdiffusion >>
rect 228 390 229 391 
<< pdiffusion >>
rect 229 390 230 391 
<< pdiffusion >>
rect 230 390 231 391 
<< pdiffusion >>
rect 231 390 232 391 
<< pdiffusion >>
rect 232 390 233 391 
<< pdiffusion >>
rect 233 390 234 391 
<< pdiffusion >>
rect 246 390 247 391 
<< pdiffusion >>
rect 247 390 248 391 
<< pdiffusion >>
rect 248 390 249 391 
<< pdiffusion >>
rect 249 390 250 391 
<< pdiffusion >>
rect 250 390 251 391 
<< pdiffusion >>
rect 251 390 252 391 
<< pdiffusion >>
rect 282 390 283 391 
<< pdiffusion >>
rect 283 390 284 391 
<< pdiffusion >>
rect 284 390 285 391 
<< pdiffusion >>
rect 285 390 286 391 
<< pdiffusion >>
rect 286 390 287 391 
<< pdiffusion >>
rect 287 390 288 391 
<< m1 >>
rect 289 390 290 391 
<< m2 >>
rect 290 390 291 391 
<< pdiffusion >>
rect 300 390 301 391 
<< pdiffusion >>
rect 301 390 302 391 
<< pdiffusion >>
rect 302 390 303 391 
<< pdiffusion >>
rect 303 390 304 391 
<< pdiffusion >>
rect 304 390 305 391 
<< pdiffusion >>
rect 305 390 306 391 
<< pdiffusion >>
rect 318 390 319 391 
<< pdiffusion >>
rect 319 390 320 391 
<< pdiffusion >>
rect 320 390 321 391 
<< pdiffusion >>
rect 321 390 322 391 
<< pdiffusion >>
rect 322 390 323 391 
<< pdiffusion >>
rect 323 390 324 391 
<< pdiffusion >>
rect 336 390 337 391 
<< pdiffusion >>
rect 337 390 338 391 
<< pdiffusion >>
rect 338 390 339 391 
<< pdiffusion >>
rect 339 390 340 391 
<< pdiffusion >>
rect 340 390 341 391 
<< pdiffusion >>
rect 341 390 342 391 
<< pdiffusion >>
rect 354 390 355 391 
<< pdiffusion >>
rect 355 390 356 391 
<< pdiffusion >>
rect 356 390 357 391 
<< pdiffusion >>
rect 357 390 358 391 
<< pdiffusion >>
rect 358 390 359 391 
<< pdiffusion >>
rect 359 390 360 391 
<< pdiffusion >>
rect 372 390 373 391 
<< pdiffusion >>
rect 373 390 374 391 
<< pdiffusion >>
rect 374 390 375 391 
<< pdiffusion >>
rect 375 390 376 391 
<< pdiffusion >>
rect 376 390 377 391 
<< pdiffusion >>
rect 377 390 378 391 
<< pdiffusion >>
rect 390 390 391 391 
<< pdiffusion >>
rect 391 390 392 391 
<< pdiffusion >>
rect 392 390 393 391 
<< pdiffusion >>
rect 393 390 394 391 
<< pdiffusion >>
rect 394 390 395 391 
<< pdiffusion >>
rect 395 390 396 391 
<< pdiffusion >>
rect 408 390 409 391 
<< pdiffusion >>
rect 409 390 410 391 
<< pdiffusion >>
rect 410 390 411 391 
<< pdiffusion >>
rect 411 390 412 391 
<< pdiffusion >>
rect 412 390 413 391 
<< pdiffusion >>
rect 413 390 414 391 
<< pdiffusion >>
rect 426 390 427 391 
<< pdiffusion >>
rect 427 390 428 391 
<< pdiffusion >>
rect 428 390 429 391 
<< pdiffusion >>
rect 429 390 430 391 
<< pdiffusion >>
rect 430 390 431 391 
<< pdiffusion >>
rect 431 390 432 391 
<< pdiffusion >>
rect 444 390 445 391 
<< pdiffusion >>
rect 445 390 446 391 
<< pdiffusion >>
rect 446 390 447 391 
<< pdiffusion >>
rect 447 390 448 391 
<< pdiffusion >>
rect 448 390 449 391 
<< pdiffusion >>
rect 449 390 450 391 
<< pdiffusion >>
rect 12 391 13 392 
<< pdiffusion >>
rect 13 391 14 392 
<< pdiffusion >>
rect 14 391 15 392 
<< pdiffusion >>
rect 15 391 16 392 
<< pdiffusion >>
rect 16 391 17 392 
<< pdiffusion >>
rect 17 391 18 392 
<< pdiffusion >>
rect 30 391 31 392 
<< pdiffusion >>
rect 31 391 32 392 
<< pdiffusion >>
rect 32 391 33 392 
<< pdiffusion >>
rect 33 391 34 392 
<< pdiffusion >>
rect 34 391 35 392 
<< pdiffusion >>
rect 35 391 36 392 
<< pdiffusion >>
rect 48 391 49 392 
<< pdiffusion >>
rect 49 391 50 392 
<< pdiffusion >>
rect 50 391 51 392 
<< pdiffusion >>
rect 51 391 52 392 
<< pdiffusion >>
rect 52 391 53 392 
<< pdiffusion >>
rect 53 391 54 392 
<< m1 >>
rect 64 391 65 392 
<< pdiffusion >>
rect 66 391 67 392 
<< pdiffusion >>
rect 67 391 68 392 
<< pdiffusion >>
rect 68 391 69 392 
<< pdiffusion >>
rect 69 391 70 392 
<< pdiffusion >>
rect 70 391 71 392 
<< pdiffusion >>
rect 71 391 72 392 
<< m1 >>
rect 82 391 83 392 
<< pdiffusion >>
rect 84 391 85 392 
<< pdiffusion >>
rect 85 391 86 392 
<< pdiffusion >>
rect 86 391 87 392 
<< pdiffusion >>
rect 87 391 88 392 
<< pdiffusion >>
rect 88 391 89 392 
<< pdiffusion >>
rect 89 391 90 392 
<< pdiffusion >>
rect 102 391 103 392 
<< pdiffusion >>
rect 103 391 104 392 
<< pdiffusion >>
rect 104 391 105 392 
<< pdiffusion >>
rect 105 391 106 392 
<< pdiffusion >>
rect 106 391 107 392 
<< pdiffusion >>
rect 107 391 108 392 
<< m1 >>
rect 109 391 110 392 
<< pdiffusion >>
rect 120 391 121 392 
<< pdiffusion >>
rect 121 391 122 392 
<< pdiffusion >>
rect 122 391 123 392 
<< pdiffusion >>
rect 123 391 124 392 
<< pdiffusion >>
rect 124 391 125 392 
<< pdiffusion >>
rect 125 391 126 392 
<< m1 >>
rect 127 391 128 392 
<< pdiffusion >>
rect 138 391 139 392 
<< pdiffusion >>
rect 139 391 140 392 
<< pdiffusion >>
rect 140 391 141 392 
<< pdiffusion >>
rect 141 391 142 392 
<< pdiffusion >>
rect 142 391 143 392 
<< pdiffusion >>
rect 143 391 144 392 
<< m1 >>
rect 145 391 146 392 
<< pdiffusion >>
rect 156 391 157 392 
<< pdiffusion >>
rect 157 391 158 392 
<< pdiffusion >>
rect 158 391 159 392 
<< pdiffusion >>
rect 159 391 160 392 
<< pdiffusion >>
rect 160 391 161 392 
<< pdiffusion >>
rect 161 391 162 392 
<< m1 >>
rect 172 391 173 392 
<< pdiffusion >>
rect 174 391 175 392 
<< pdiffusion >>
rect 175 391 176 392 
<< pdiffusion >>
rect 176 391 177 392 
<< pdiffusion >>
rect 177 391 178 392 
<< pdiffusion >>
rect 178 391 179 392 
<< pdiffusion >>
rect 179 391 180 392 
<< pdiffusion >>
rect 192 391 193 392 
<< pdiffusion >>
rect 193 391 194 392 
<< pdiffusion >>
rect 194 391 195 392 
<< pdiffusion >>
rect 195 391 196 392 
<< pdiffusion >>
rect 196 391 197 392 
<< pdiffusion >>
rect 197 391 198 392 
<< pdiffusion >>
rect 210 391 211 392 
<< pdiffusion >>
rect 211 391 212 392 
<< pdiffusion >>
rect 212 391 213 392 
<< pdiffusion >>
rect 213 391 214 392 
<< pdiffusion >>
rect 214 391 215 392 
<< pdiffusion >>
rect 215 391 216 392 
<< pdiffusion >>
rect 228 391 229 392 
<< pdiffusion >>
rect 229 391 230 392 
<< pdiffusion >>
rect 230 391 231 392 
<< pdiffusion >>
rect 231 391 232 392 
<< pdiffusion >>
rect 232 391 233 392 
<< pdiffusion >>
rect 233 391 234 392 
<< pdiffusion >>
rect 246 391 247 392 
<< pdiffusion >>
rect 247 391 248 392 
<< pdiffusion >>
rect 248 391 249 392 
<< pdiffusion >>
rect 249 391 250 392 
<< pdiffusion >>
rect 250 391 251 392 
<< pdiffusion >>
rect 251 391 252 392 
<< pdiffusion >>
rect 282 391 283 392 
<< pdiffusion >>
rect 283 391 284 392 
<< pdiffusion >>
rect 284 391 285 392 
<< pdiffusion >>
rect 285 391 286 392 
<< pdiffusion >>
rect 286 391 287 392 
<< pdiffusion >>
rect 287 391 288 392 
<< m1 >>
rect 289 391 290 392 
<< m2 >>
rect 290 391 291 392 
<< pdiffusion >>
rect 300 391 301 392 
<< pdiffusion >>
rect 301 391 302 392 
<< pdiffusion >>
rect 302 391 303 392 
<< pdiffusion >>
rect 303 391 304 392 
<< pdiffusion >>
rect 304 391 305 392 
<< pdiffusion >>
rect 305 391 306 392 
<< pdiffusion >>
rect 318 391 319 392 
<< pdiffusion >>
rect 319 391 320 392 
<< pdiffusion >>
rect 320 391 321 392 
<< pdiffusion >>
rect 321 391 322 392 
<< pdiffusion >>
rect 322 391 323 392 
<< pdiffusion >>
rect 323 391 324 392 
<< pdiffusion >>
rect 336 391 337 392 
<< pdiffusion >>
rect 337 391 338 392 
<< pdiffusion >>
rect 338 391 339 392 
<< pdiffusion >>
rect 339 391 340 392 
<< pdiffusion >>
rect 340 391 341 392 
<< pdiffusion >>
rect 341 391 342 392 
<< pdiffusion >>
rect 354 391 355 392 
<< pdiffusion >>
rect 355 391 356 392 
<< pdiffusion >>
rect 356 391 357 392 
<< pdiffusion >>
rect 357 391 358 392 
<< pdiffusion >>
rect 358 391 359 392 
<< pdiffusion >>
rect 359 391 360 392 
<< pdiffusion >>
rect 372 391 373 392 
<< pdiffusion >>
rect 373 391 374 392 
<< pdiffusion >>
rect 374 391 375 392 
<< pdiffusion >>
rect 375 391 376 392 
<< pdiffusion >>
rect 376 391 377 392 
<< pdiffusion >>
rect 377 391 378 392 
<< pdiffusion >>
rect 390 391 391 392 
<< pdiffusion >>
rect 391 391 392 392 
<< pdiffusion >>
rect 392 391 393 392 
<< pdiffusion >>
rect 393 391 394 392 
<< pdiffusion >>
rect 394 391 395 392 
<< pdiffusion >>
rect 395 391 396 392 
<< pdiffusion >>
rect 408 391 409 392 
<< pdiffusion >>
rect 409 391 410 392 
<< pdiffusion >>
rect 410 391 411 392 
<< pdiffusion >>
rect 411 391 412 392 
<< pdiffusion >>
rect 412 391 413 392 
<< pdiffusion >>
rect 413 391 414 392 
<< pdiffusion >>
rect 426 391 427 392 
<< pdiffusion >>
rect 427 391 428 392 
<< pdiffusion >>
rect 428 391 429 392 
<< pdiffusion >>
rect 429 391 430 392 
<< pdiffusion >>
rect 430 391 431 392 
<< pdiffusion >>
rect 431 391 432 392 
<< pdiffusion >>
rect 444 391 445 392 
<< pdiffusion >>
rect 445 391 446 392 
<< pdiffusion >>
rect 446 391 447 392 
<< pdiffusion >>
rect 447 391 448 392 
<< pdiffusion >>
rect 448 391 449 392 
<< pdiffusion >>
rect 449 391 450 392 
<< pdiffusion >>
rect 12 392 13 393 
<< pdiffusion >>
rect 13 392 14 393 
<< pdiffusion >>
rect 14 392 15 393 
<< pdiffusion >>
rect 15 392 16 393 
<< pdiffusion >>
rect 16 392 17 393 
<< pdiffusion >>
rect 17 392 18 393 
<< pdiffusion >>
rect 30 392 31 393 
<< pdiffusion >>
rect 31 392 32 393 
<< pdiffusion >>
rect 32 392 33 393 
<< pdiffusion >>
rect 33 392 34 393 
<< pdiffusion >>
rect 34 392 35 393 
<< pdiffusion >>
rect 35 392 36 393 
<< pdiffusion >>
rect 48 392 49 393 
<< pdiffusion >>
rect 49 392 50 393 
<< pdiffusion >>
rect 50 392 51 393 
<< pdiffusion >>
rect 51 392 52 393 
<< pdiffusion >>
rect 52 392 53 393 
<< pdiffusion >>
rect 53 392 54 393 
<< m1 >>
rect 64 392 65 393 
<< pdiffusion >>
rect 66 392 67 393 
<< pdiffusion >>
rect 67 392 68 393 
<< pdiffusion >>
rect 68 392 69 393 
<< pdiffusion >>
rect 69 392 70 393 
<< pdiffusion >>
rect 70 392 71 393 
<< pdiffusion >>
rect 71 392 72 393 
<< m1 >>
rect 82 392 83 393 
<< pdiffusion >>
rect 84 392 85 393 
<< pdiffusion >>
rect 85 392 86 393 
<< pdiffusion >>
rect 86 392 87 393 
<< pdiffusion >>
rect 87 392 88 393 
<< pdiffusion >>
rect 88 392 89 393 
<< pdiffusion >>
rect 89 392 90 393 
<< pdiffusion >>
rect 102 392 103 393 
<< pdiffusion >>
rect 103 392 104 393 
<< pdiffusion >>
rect 104 392 105 393 
<< pdiffusion >>
rect 105 392 106 393 
<< pdiffusion >>
rect 106 392 107 393 
<< pdiffusion >>
rect 107 392 108 393 
<< m1 >>
rect 109 392 110 393 
<< pdiffusion >>
rect 120 392 121 393 
<< pdiffusion >>
rect 121 392 122 393 
<< pdiffusion >>
rect 122 392 123 393 
<< pdiffusion >>
rect 123 392 124 393 
<< pdiffusion >>
rect 124 392 125 393 
<< pdiffusion >>
rect 125 392 126 393 
<< m1 >>
rect 127 392 128 393 
<< pdiffusion >>
rect 138 392 139 393 
<< pdiffusion >>
rect 139 392 140 393 
<< pdiffusion >>
rect 140 392 141 393 
<< pdiffusion >>
rect 141 392 142 393 
<< pdiffusion >>
rect 142 392 143 393 
<< pdiffusion >>
rect 143 392 144 393 
<< m1 >>
rect 145 392 146 393 
<< pdiffusion >>
rect 156 392 157 393 
<< pdiffusion >>
rect 157 392 158 393 
<< pdiffusion >>
rect 158 392 159 393 
<< pdiffusion >>
rect 159 392 160 393 
<< pdiffusion >>
rect 160 392 161 393 
<< pdiffusion >>
rect 161 392 162 393 
<< m1 >>
rect 172 392 173 393 
<< pdiffusion >>
rect 174 392 175 393 
<< pdiffusion >>
rect 175 392 176 393 
<< pdiffusion >>
rect 176 392 177 393 
<< pdiffusion >>
rect 177 392 178 393 
<< pdiffusion >>
rect 178 392 179 393 
<< pdiffusion >>
rect 179 392 180 393 
<< pdiffusion >>
rect 192 392 193 393 
<< pdiffusion >>
rect 193 392 194 393 
<< pdiffusion >>
rect 194 392 195 393 
<< pdiffusion >>
rect 195 392 196 393 
<< pdiffusion >>
rect 196 392 197 393 
<< pdiffusion >>
rect 197 392 198 393 
<< pdiffusion >>
rect 210 392 211 393 
<< pdiffusion >>
rect 211 392 212 393 
<< pdiffusion >>
rect 212 392 213 393 
<< pdiffusion >>
rect 213 392 214 393 
<< pdiffusion >>
rect 214 392 215 393 
<< pdiffusion >>
rect 215 392 216 393 
<< pdiffusion >>
rect 228 392 229 393 
<< pdiffusion >>
rect 229 392 230 393 
<< pdiffusion >>
rect 230 392 231 393 
<< pdiffusion >>
rect 231 392 232 393 
<< pdiffusion >>
rect 232 392 233 393 
<< pdiffusion >>
rect 233 392 234 393 
<< pdiffusion >>
rect 246 392 247 393 
<< pdiffusion >>
rect 247 392 248 393 
<< pdiffusion >>
rect 248 392 249 393 
<< pdiffusion >>
rect 249 392 250 393 
<< pdiffusion >>
rect 250 392 251 393 
<< pdiffusion >>
rect 251 392 252 393 
<< pdiffusion >>
rect 282 392 283 393 
<< pdiffusion >>
rect 283 392 284 393 
<< pdiffusion >>
rect 284 392 285 393 
<< pdiffusion >>
rect 285 392 286 393 
<< pdiffusion >>
rect 286 392 287 393 
<< pdiffusion >>
rect 287 392 288 393 
<< m1 >>
rect 289 392 290 393 
<< m2 >>
rect 290 392 291 393 
<< pdiffusion >>
rect 300 392 301 393 
<< pdiffusion >>
rect 301 392 302 393 
<< pdiffusion >>
rect 302 392 303 393 
<< pdiffusion >>
rect 303 392 304 393 
<< pdiffusion >>
rect 304 392 305 393 
<< pdiffusion >>
rect 305 392 306 393 
<< pdiffusion >>
rect 318 392 319 393 
<< pdiffusion >>
rect 319 392 320 393 
<< pdiffusion >>
rect 320 392 321 393 
<< pdiffusion >>
rect 321 392 322 393 
<< pdiffusion >>
rect 322 392 323 393 
<< pdiffusion >>
rect 323 392 324 393 
<< pdiffusion >>
rect 336 392 337 393 
<< pdiffusion >>
rect 337 392 338 393 
<< pdiffusion >>
rect 338 392 339 393 
<< pdiffusion >>
rect 339 392 340 393 
<< pdiffusion >>
rect 340 392 341 393 
<< pdiffusion >>
rect 341 392 342 393 
<< pdiffusion >>
rect 354 392 355 393 
<< pdiffusion >>
rect 355 392 356 393 
<< pdiffusion >>
rect 356 392 357 393 
<< pdiffusion >>
rect 357 392 358 393 
<< pdiffusion >>
rect 358 392 359 393 
<< pdiffusion >>
rect 359 392 360 393 
<< pdiffusion >>
rect 372 392 373 393 
<< pdiffusion >>
rect 373 392 374 393 
<< pdiffusion >>
rect 374 392 375 393 
<< pdiffusion >>
rect 375 392 376 393 
<< pdiffusion >>
rect 376 392 377 393 
<< pdiffusion >>
rect 377 392 378 393 
<< pdiffusion >>
rect 390 392 391 393 
<< pdiffusion >>
rect 391 392 392 393 
<< pdiffusion >>
rect 392 392 393 393 
<< pdiffusion >>
rect 393 392 394 393 
<< pdiffusion >>
rect 394 392 395 393 
<< pdiffusion >>
rect 395 392 396 393 
<< pdiffusion >>
rect 408 392 409 393 
<< pdiffusion >>
rect 409 392 410 393 
<< pdiffusion >>
rect 410 392 411 393 
<< pdiffusion >>
rect 411 392 412 393 
<< pdiffusion >>
rect 412 392 413 393 
<< pdiffusion >>
rect 413 392 414 393 
<< pdiffusion >>
rect 426 392 427 393 
<< pdiffusion >>
rect 427 392 428 393 
<< pdiffusion >>
rect 428 392 429 393 
<< pdiffusion >>
rect 429 392 430 393 
<< pdiffusion >>
rect 430 392 431 393 
<< pdiffusion >>
rect 431 392 432 393 
<< pdiffusion >>
rect 444 392 445 393 
<< pdiffusion >>
rect 445 392 446 393 
<< pdiffusion >>
rect 446 392 447 393 
<< pdiffusion >>
rect 447 392 448 393 
<< pdiffusion >>
rect 448 392 449 393 
<< pdiffusion >>
rect 449 392 450 393 
<< pdiffusion >>
rect 12 393 13 394 
<< pdiffusion >>
rect 13 393 14 394 
<< pdiffusion >>
rect 14 393 15 394 
<< pdiffusion >>
rect 15 393 16 394 
<< pdiffusion >>
rect 16 393 17 394 
<< pdiffusion >>
rect 17 393 18 394 
<< pdiffusion >>
rect 30 393 31 394 
<< pdiffusion >>
rect 31 393 32 394 
<< pdiffusion >>
rect 32 393 33 394 
<< pdiffusion >>
rect 33 393 34 394 
<< pdiffusion >>
rect 34 393 35 394 
<< pdiffusion >>
rect 35 393 36 394 
<< pdiffusion >>
rect 48 393 49 394 
<< pdiffusion >>
rect 49 393 50 394 
<< pdiffusion >>
rect 50 393 51 394 
<< pdiffusion >>
rect 51 393 52 394 
<< pdiffusion >>
rect 52 393 53 394 
<< pdiffusion >>
rect 53 393 54 394 
<< m1 >>
rect 64 393 65 394 
<< pdiffusion >>
rect 66 393 67 394 
<< pdiffusion >>
rect 67 393 68 394 
<< pdiffusion >>
rect 68 393 69 394 
<< pdiffusion >>
rect 69 393 70 394 
<< pdiffusion >>
rect 70 393 71 394 
<< pdiffusion >>
rect 71 393 72 394 
<< m1 >>
rect 82 393 83 394 
<< pdiffusion >>
rect 84 393 85 394 
<< pdiffusion >>
rect 85 393 86 394 
<< pdiffusion >>
rect 86 393 87 394 
<< pdiffusion >>
rect 87 393 88 394 
<< pdiffusion >>
rect 88 393 89 394 
<< pdiffusion >>
rect 89 393 90 394 
<< pdiffusion >>
rect 102 393 103 394 
<< pdiffusion >>
rect 103 393 104 394 
<< pdiffusion >>
rect 104 393 105 394 
<< pdiffusion >>
rect 105 393 106 394 
<< pdiffusion >>
rect 106 393 107 394 
<< pdiffusion >>
rect 107 393 108 394 
<< m1 >>
rect 109 393 110 394 
<< pdiffusion >>
rect 120 393 121 394 
<< pdiffusion >>
rect 121 393 122 394 
<< pdiffusion >>
rect 122 393 123 394 
<< pdiffusion >>
rect 123 393 124 394 
<< pdiffusion >>
rect 124 393 125 394 
<< pdiffusion >>
rect 125 393 126 394 
<< m1 >>
rect 127 393 128 394 
<< pdiffusion >>
rect 138 393 139 394 
<< pdiffusion >>
rect 139 393 140 394 
<< pdiffusion >>
rect 140 393 141 394 
<< pdiffusion >>
rect 141 393 142 394 
<< pdiffusion >>
rect 142 393 143 394 
<< pdiffusion >>
rect 143 393 144 394 
<< m1 >>
rect 145 393 146 394 
<< pdiffusion >>
rect 156 393 157 394 
<< pdiffusion >>
rect 157 393 158 394 
<< pdiffusion >>
rect 158 393 159 394 
<< pdiffusion >>
rect 159 393 160 394 
<< pdiffusion >>
rect 160 393 161 394 
<< pdiffusion >>
rect 161 393 162 394 
<< m1 >>
rect 172 393 173 394 
<< pdiffusion >>
rect 174 393 175 394 
<< pdiffusion >>
rect 175 393 176 394 
<< pdiffusion >>
rect 176 393 177 394 
<< pdiffusion >>
rect 177 393 178 394 
<< pdiffusion >>
rect 178 393 179 394 
<< pdiffusion >>
rect 179 393 180 394 
<< pdiffusion >>
rect 192 393 193 394 
<< pdiffusion >>
rect 193 393 194 394 
<< pdiffusion >>
rect 194 393 195 394 
<< pdiffusion >>
rect 195 393 196 394 
<< pdiffusion >>
rect 196 393 197 394 
<< pdiffusion >>
rect 197 393 198 394 
<< pdiffusion >>
rect 210 393 211 394 
<< pdiffusion >>
rect 211 393 212 394 
<< pdiffusion >>
rect 212 393 213 394 
<< pdiffusion >>
rect 213 393 214 394 
<< pdiffusion >>
rect 214 393 215 394 
<< pdiffusion >>
rect 215 393 216 394 
<< pdiffusion >>
rect 228 393 229 394 
<< pdiffusion >>
rect 229 393 230 394 
<< pdiffusion >>
rect 230 393 231 394 
<< pdiffusion >>
rect 231 393 232 394 
<< pdiffusion >>
rect 232 393 233 394 
<< pdiffusion >>
rect 233 393 234 394 
<< pdiffusion >>
rect 246 393 247 394 
<< pdiffusion >>
rect 247 393 248 394 
<< pdiffusion >>
rect 248 393 249 394 
<< pdiffusion >>
rect 249 393 250 394 
<< pdiffusion >>
rect 250 393 251 394 
<< pdiffusion >>
rect 251 393 252 394 
<< pdiffusion >>
rect 282 393 283 394 
<< pdiffusion >>
rect 283 393 284 394 
<< pdiffusion >>
rect 284 393 285 394 
<< pdiffusion >>
rect 285 393 286 394 
<< pdiffusion >>
rect 286 393 287 394 
<< pdiffusion >>
rect 287 393 288 394 
<< m1 >>
rect 289 393 290 394 
<< m2 >>
rect 290 393 291 394 
<< pdiffusion >>
rect 300 393 301 394 
<< pdiffusion >>
rect 301 393 302 394 
<< pdiffusion >>
rect 302 393 303 394 
<< pdiffusion >>
rect 303 393 304 394 
<< pdiffusion >>
rect 304 393 305 394 
<< pdiffusion >>
rect 305 393 306 394 
<< pdiffusion >>
rect 318 393 319 394 
<< pdiffusion >>
rect 319 393 320 394 
<< pdiffusion >>
rect 320 393 321 394 
<< pdiffusion >>
rect 321 393 322 394 
<< pdiffusion >>
rect 322 393 323 394 
<< pdiffusion >>
rect 323 393 324 394 
<< pdiffusion >>
rect 336 393 337 394 
<< pdiffusion >>
rect 337 393 338 394 
<< pdiffusion >>
rect 338 393 339 394 
<< pdiffusion >>
rect 339 393 340 394 
<< pdiffusion >>
rect 340 393 341 394 
<< pdiffusion >>
rect 341 393 342 394 
<< pdiffusion >>
rect 354 393 355 394 
<< pdiffusion >>
rect 355 393 356 394 
<< pdiffusion >>
rect 356 393 357 394 
<< pdiffusion >>
rect 357 393 358 394 
<< pdiffusion >>
rect 358 393 359 394 
<< pdiffusion >>
rect 359 393 360 394 
<< pdiffusion >>
rect 372 393 373 394 
<< pdiffusion >>
rect 373 393 374 394 
<< pdiffusion >>
rect 374 393 375 394 
<< pdiffusion >>
rect 375 393 376 394 
<< pdiffusion >>
rect 376 393 377 394 
<< pdiffusion >>
rect 377 393 378 394 
<< pdiffusion >>
rect 390 393 391 394 
<< pdiffusion >>
rect 391 393 392 394 
<< pdiffusion >>
rect 392 393 393 394 
<< pdiffusion >>
rect 393 393 394 394 
<< pdiffusion >>
rect 394 393 395 394 
<< pdiffusion >>
rect 395 393 396 394 
<< pdiffusion >>
rect 408 393 409 394 
<< pdiffusion >>
rect 409 393 410 394 
<< pdiffusion >>
rect 410 393 411 394 
<< pdiffusion >>
rect 411 393 412 394 
<< pdiffusion >>
rect 412 393 413 394 
<< pdiffusion >>
rect 413 393 414 394 
<< pdiffusion >>
rect 426 393 427 394 
<< pdiffusion >>
rect 427 393 428 394 
<< pdiffusion >>
rect 428 393 429 394 
<< pdiffusion >>
rect 429 393 430 394 
<< pdiffusion >>
rect 430 393 431 394 
<< pdiffusion >>
rect 431 393 432 394 
<< pdiffusion >>
rect 444 393 445 394 
<< pdiffusion >>
rect 445 393 446 394 
<< pdiffusion >>
rect 446 393 447 394 
<< pdiffusion >>
rect 447 393 448 394 
<< pdiffusion >>
rect 448 393 449 394 
<< pdiffusion >>
rect 449 393 450 394 
<< pdiffusion >>
rect 12 394 13 395 
<< pdiffusion >>
rect 13 394 14 395 
<< pdiffusion >>
rect 14 394 15 395 
<< pdiffusion >>
rect 15 394 16 395 
<< pdiffusion >>
rect 16 394 17 395 
<< pdiffusion >>
rect 17 394 18 395 
<< pdiffusion >>
rect 30 394 31 395 
<< pdiffusion >>
rect 31 394 32 395 
<< pdiffusion >>
rect 32 394 33 395 
<< pdiffusion >>
rect 33 394 34 395 
<< pdiffusion >>
rect 34 394 35 395 
<< pdiffusion >>
rect 35 394 36 395 
<< pdiffusion >>
rect 48 394 49 395 
<< pdiffusion >>
rect 49 394 50 395 
<< pdiffusion >>
rect 50 394 51 395 
<< pdiffusion >>
rect 51 394 52 395 
<< pdiffusion >>
rect 52 394 53 395 
<< pdiffusion >>
rect 53 394 54 395 
<< m1 >>
rect 64 394 65 395 
<< pdiffusion >>
rect 66 394 67 395 
<< pdiffusion >>
rect 67 394 68 395 
<< pdiffusion >>
rect 68 394 69 395 
<< pdiffusion >>
rect 69 394 70 395 
<< pdiffusion >>
rect 70 394 71 395 
<< pdiffusion >>
rect 71 394 72 395 
<< m1 >>
rect 82 394 83 395 
<< pdiffusion >>
rect 84 394 85 395 
<< pdiffusion >>
rect 85 394 86 395 
<< pdiffusion >>
rect 86 394 87 395 
<< pdiffusion >>
rect 87 394 88 395 
<< pdiffusion >>
rect 88 394 89 395 
<< pdiffusion >>
rect 89 394 90 395 
<< pdiffusion >>
rect 102 394 103 395 
<< pdiffusion >>
rect 103 394 104 395 
<< pdiffusion >>
rect 104 394 105 395 
<< pdiffusion >>
rect 105 394 106 395 
<< pdiffusion >>
rect 106 394 107 395 
<< pdiffusion >>
rect 107 394 108 395 
<< m1 >>
rect 109 394 110 395 
<< pdiffusion >>
rect 120 394 121 395 
<< pdiffusion >>
rect 121 394 122 395 
<< pdiffusion >>
rect 122 394 123 395 
<< pdiffusion >>
rect 123 394 124 395 
<< pdiffusion >>
rect 124 394 125 395 
<< pdiffusion >>
rect 125 394 126 395 
<< m1 >>
rect 127 394 128 395 
<< pdiffusion >>
rect 138 394 139 395 
<< pdiffusion >>
rect 139 394 140 395 
<< pdiffusion >>
rect 140 394 141 395 
<< pdiffusion >>
rect 141 394 142 395 
<< pdiffusion >>
rect 142 394 143 395 
<< pdiffusion >>
rect 143 394 144 395 
<< m1 >>
rect 145 394 146 395 
<< pdiffusion >>
rect 156 394 157 395 
<< pdiffusion >>
rect 157 394 158 395 
<< pdiffusion >>
rect 158 394 159 395 
<< pdiffusion >>
rect 159 394 160 395 
<< pdiffusion >>
rect 160 394 161 395 
<< pdiffusion >>
rect 161 394 162 395 
<< m1 >>
rect 172 394 173 395 
<< pdiffusion >>
rect 174 394 175 395 
<< pdiffusion >>
rect 175 394 176 395 
<< pdiffusion >>
rect 176 394 177 395 
<< pdiffusion >>
rect 177 394 178 395 
<< pdiffusion >>
rect 178 394 179 395 
<< pdiffusion >>
rect 179 394 180 395 
<< pdiffusion >>
rect 192 394 193 395 
<< pdiffusion >>
rect 193 394 194 395 
<< pdiffusion >>
rect 194 394 195 395 
<< pdiffusion >>
rect 195 394 196 395 
<< pdiffusion >>
rect 196 394 197 395 
<< pdiffusion >>
rect 197 394 198 395 
<< pdiffusion >>
rect 210 394 211 395 
<< pdiffusion >>
rect 211 394 212 395 
<< pdiffusion >>
rect 212 394 213 395 
<< pdiffusion >>
rect 213 394 214 395 
<< pdiffusion >>
rect 214 394 215 395 
<< pdiffusion >>
rect 215 394 216 395 
<< pdiffusion >>
rect 228 394 229 395 
<< pdiffusion >>
rect 229 394 230 395 
<< pdiffusion >>
rect 230 394 231 395 
<< pdiffusion >>
rect 231 394 232 395 
<< pdiffusion >>
rect 232 394 233 395 
<< pdiffusion >>
rect 233 394 234 395 
<< pdiffusion >>
rect 246 394 247 395 
<< pdiffusion >>
rect 247 394 248 395 
<< pdiffusion >>
rect 248 394 249 395 
<< pdiffusion >>
rect 249 394 250 395 
<< pdiffusion >>
rect 250 394 251 395 
<< pdiffusion >>
rect 251 394 252 395 
<< pdiffusion >>
rect 282 394 283 395 
<< pdiffusion >>
rect 283 394 284 395 
<< pdiffusion >>
rect 284 394 285 395 
<< pdiffusion >>
rect 285 394 286 395 
<< pdiffusion >>
rect 286 394 287 395 
<< pdiffusion >>
rect 287 394 288 395 
<< m1 >>
rect 289 394 290 395 
<< m2 >>
rect 290 394 291 395 
<< pdiffusion >>
rect 300 394 301 395 
<< pdiffusion >>
rect 301 394 302 395 
<< pdiffusion >>
rect 302 394 303 395 
<< pdiffusion >>
rect 303 394 304 395 
<< pdiffusion >>
rect 304 394 305 395 
<< pdiffusion >>
rect 305 394 306 395 
<< pdiffusion >>
rect 318 394 319 395 
<< pdiffusion >>
rect 319 394 320 395 
<< pdiffusion >>
rect 320 394 321 395 
<< pdiffusion >>
rect 321 394 322 395 
<< pdiffusion >>
rect 322 394 323 395 
<< pdiffusion >>
rect 323 394 324 395 
<< pdiffusion >>
rect 336 394 337 395 
<< pdiffusion >>
rect 337 394 338 395 
<< pdiffusion >>
rect 338 394 339 395 
<< pdiffusion >>
rect 339 394 340 395 
<< pdiffusion >>
rect 340 394 341 395 
<< pdiffusion >>
rect 341 394 342 395 
<< pdiffusion >>
rect 354 394 355 395 
<< pdiffusion >>
rect 355 394 356 395 
<< pdiffusion >>
rect 356 394 357 395 
<< pdiffusion >>
rect 357 394 358 395 
<< pdiffusion >>
rect 358 394 359 395 
<< pdiffusion >>
rect 359 394 360 395 
<< pdiffusion >>
rect 372 394 373 395 
<< pdiffusion >>
rect 373 394 374 395 
<< pdiffusion >>
rect 374 394 375 395 
<< pdiffusion >>
rect 375 394 376 395 
<< pdiffusion >>
rect 376 394 377 395 
<< pdiffusion >>
rect 377 394 378 395 
<< pdiffusion >>
rect 390 394 391 395 
<< pdiffusion >>
rect 391 394 392 395 
<< pdiffusion >>
rect 392 394 393 395 
<< pdiffusion >>
rect 393 394 394 395 
<< pdiffusion >>
rect 394 394 395 395 
<< pdiffusion >>
rect 395 394 396 395 
<< pdiffusion >>
rect 408 394 409 395 
<< pdiffusion >>
rect 409 394 410 395 
<< pdiffusion >>
rect 410 394 411 395 
<< pdiffusion >>
rect 411 394 412 395 
<< pdiffusion >>
rect 412 394 413 395 
<< pdiffusion >>
rect 413 394 414 395 
<< pdiffusion >>
rect 426 394 427 395 
<< pdiffusion >>
rect 427 394 428 395 
<< pdiffusion >>
rect 428 394 429 395 
<< pdiffusion >>
rect 429 394 430 395 
<< pdiffusion >>
rect 430 394 431 395 
<< pdiffusion >>
rect 431 394 432 395 
<< pdiffusion >>
rect 444 394 445 395 
<< pdiffusion >>
rect 445 394 446 395 
<< pdiffusion >>
rect 446 394 447 395 
<< pdiffusion >>
rect 447 394 448 395 
<< pdiffusion >>
rect 448 394 449 395 
<< pdiffusion >>
rect 449 394 450 395 
<< pdiffusion >>
rect 12 395 13 396 
<< pdiffusion >>
rect 13 395 14 396 
<< pdiffusion >>
rect 14 395 15 396 
<< pdiffusion >>
rect 15 395 16 396 
<< pdiffusion >>
rect 16 395 17 396 
<< pdiffusion >>
rect 17 395 18 396 
<< pdiffusion >>
rect 30 395 31 396 
<< pdiffusion >>
rect 31 395 32 396 
<< pdiffusion >>
rect 32 395 33 396 
<< pdiffusion >>
rect 33 395 34 396 
<< pdiffusion >>
rect 34 395 35 396 
<< pdiffusion >>
rect 35 395 36 396 
<< pdiffusion >>
rect 48 395 49 396 
<< pdiffusion >>
rect 49 395 50 396 
<< pdiffusion >>
rect 50 395 51 396 
<< pdiffusion >>
rect 51 395 52 396 
<< pdiffusion >>
rect 52 395 53 396 
<< pdiffusion >>
rect 53 395 54 396 
<< m1 >>
rect 64 395 65 396 
<< pdiffusion >>
rect 66 395 67 396 
<< pdiffusion >>
rect 67 395 68 396 
<< pdiffusion >>
rect 68 395 69 396 
<< pdiffusion >>
rect 69 395 70 396 
<< pdiffusion >>
rect 70 395 71 396 
<< pdiffusion >>
rect 71 395 72 396 
<< m1 >>
rect 82 395 83 396 
<< pdiffusion >>
rect 84 395 85 396 
<< m1 >>
rect 85 395 86 396 
<< pdiffusion >>
rect 85 395 86 396 
<< pdiffusion >>
rect 86 395 87 396 
<< pdiffusion >>
rect 87 395 88 396 
<< pdiffusion >>
rect 88 395 89 396 
<< pdiffusion >>
rect 89 395 90 396 
<< pdiffusion >>
rect 102 395 103 396 
<< pdiffusion >>
rect 103 395 104 396 
<< pdiffusion >>
rect 104 395 105 396 
<< pdiffusion >>
rect 105 395 106 396 
<< pdiffusion >>
rect 106 395 107 396 
<< pdiffusion >>
rect 107 395 108 396 
<< m1 >>
rect 109 395 110 396 
<< pdiffusion >>
rect 120 395 121 396 
<< pdiffusion >>
rect 121 395 122 396 
<< pdiffusion >>
rect 122 395 123 396 
<< pdiffusion >>
rect 123 395 124 396 
<< m1 >>
rect 124 395 125 396 
<< pdiffusion >>
rect 124 395 125 396 
<< pdiffusion >>
rect 125 395 126 396 
<< m1 >>
rect 127 395 128 396 
<< pdiffusion >>
rect 138 395 139 396 
<< pdiffusion >>
rect 139 395 140 396 
<< pdiffusion >>
rect 140 395 141 396 
<< pdiffusion >>
rect 141 395 142 396 
<< pdiffusion >>
rect 142 395 143 396 
<< pdiffusion >>
rect 143 395 144 396 
<< m1 >>
rect 145 395 146 396 
<< pdiffusion >>
rect 156 395 157 396 
<< pdiffusion >>
rect 157 395 158 396 
<< pdiffusion >>
rect 158 395 159 396 
<< pdiffusion >>
rect 159 395 160 396 
<< pdiffusion >>
rect 160 395 161 396 
<< pdiffusion >>
rect 161 395 162 396 
<< m1 >>
rect 172 395 173 396 
<< pdiffusion >>
rect 174 395 175 396 
<< pdiffusion >>
rect 175 395 176 396 
<< pdiffusion >>
rect 176 395 177 396 
<< pdiffusion >>
rect 177 395 178 396 
<< pdiffusion >>
rect 178 395 179 396 
<< pdiffusion >>
rect 179 395 180 396 
<< pdiffusion >>
rect 192 395 193 396 
<< pdiffusion >>
rect 193 395 194 396 
<< pdiffusion >>
rect 194 395 195 396 
<< pdiffusion >>
rect 195 395 196 396 
<< pdiffusion >>
rect 196 395 197 396 
<< pdiffusion >>
rect 197 395 198 396 
<< pdiffusion >>
rect 210 395 211 396 
<< pdiffusion >>
rect 211 395 212 396 
<< pdiffusion >>
rect 212 395 213 396 
<< pdiffusion >>
rect 213 395 214 396 
<< pdiffusion >>
rect 214 395 215 396 
<< pdiffusion >>
rect 215 395 216 396 
<< pdiffusion >>
rect 228 395 229 396 
<< pdiffusion >>
rect 229 395 230 396 
<< pdiffusion >>
rect 230 395 231 396 
<< pdiffusion >>
rect 231 395 232 396 
<< pdiffusion >>
rect 232 395 233 396 
<< pdiffusion >>
rect 233 395 234 396 
<< pdiffusion >>
rect 246 395 247 396 
<< pdiffusion >>
rect 247 395 248 396 
<< pdiffusion >>
rect 248 395 249 396 
<< pdiffusion >>
rect 249 395 250 396 
<< pdiffusion >>
rect 250 395 251 396 
<< pdiffusion >>
rect 251 395 252 396 
<< pdiffusion >>
rect 282 395 283 396 
<< pdiffusion >>
rect 283 395 284 396 
<< pdiffusion >>
rect 284 395 285 396 
<< pdiffusion >>
rect 285 395 286 396 
<< pdiffusion >>
rect 286 395 287 396 
<< pdiffusion >>
rect 287 395 288 396 
<< m1 >>
rect 289 395 290 396 
<< m2 >>
rect 290 395 291 396 
<< pdiffusion >>
rect 300 395 301 396 
<< m1 >>
rect 301 395 302 396 
<< pdiffusion >>
rect 301 395 302 396 
<< pdiffusion >>
rect 302 395 303 396 
<< pdiffusion >>
rect 303 395 304 396 
<< pdiffusion >>
rect 304 395 305 396 
<< pdiffusion >>
rect 305 395 306 396 
<< pdiffusion >>
rect 318 395 319 396 
<< pdiffusion >>
rect 319 395 320 396 
<< pdiffusion >>
rect 320 395 321 396 
<< pdiffusion >>
rect 321 395 322 396 
<< pdiffusion >>
rect 322 395 323 396 
<< pdiffusion >>
rect 323 395 324 396 
<< pdiffusion >>
rect 336 395 337 396 
<< pdiffusion >>
rect 337 395 338 396 
<< pdiffusion >>
rect 338 395 339 396 
<< pdiffusion >>
rect 339 395 340 396 
<< pdiffusion >>
rect 340 395 341 396 
<< pdiffusion >>
rect 341 395 342 396 
<< pdiffusion >>
rect 354 395 355 396 
<< pdiffusion >>
rect 355 395 356 396 
<< pdiffusion >>
rect 356 395 357 396 
<< pdiffusion >>
rect 357 395 358 396 
<< pdiffusion >>
rect 358 395 359 396 
<< pdiffusion >>
rect 359 395 360 396 
<< pdiffusion >>
rect 372 395 373 396 
<< pdiffusion >>
rect 373 395 374 396 
<< pdiffusion >>
rect 374 395 375 396 
<< pdiffusion >>
rect 375 395 376 396 
<< pdiffusion >>
rect 376 395 377 396 
<< pdiffusion >>
rect 377 395 378 396 
<< pdiffusion >>
rect 390 395 391 396 
<< pdiffusion >>
rect 391 395 392 396 
<< pdiffusion >>
rect 392 395 393 396 
<< pdiffusion >>
rect 393 395 394 396 
<< pdiffusion >>
rect 394 395 395 396 
<< pdiffusion >>
rect 395 395 396 396 
<< pdiffusion >>
rect 408 395 409 396 
<< pdiffusion >>
rect 409 395 410 396 
<< pdiffusion >>
rect 410 395 411 396 
<< pdiffusion >>
rect 411 395 412 396 
<< pdiffusion >>
rect 412 395 413 396 
<< pdiffusion >>
rect 413 395 414 396 
<< pdiffusion >>
rect 426 395 427 396 
<< pdiffusion >>
rect 427 395 428 396 
<< pdiffusion >>
rect 428 395 429 396 
<< pdiffusion >>
rect 429 395 430 396 
<< pdiffusion >>
rect 430 395 431 396 
<< pdiffusion >>
rect 431 395 432 396 
<< pdiffusion >>
rect 444 395 445 396 
<< pdiffusion >>
rect 445 395 446 396 
<< pdiffusion >>
rect 446 395 447 396 
<< pdiffusion >>
rect 447 395 448 396 
<< pdiffusion >>
rect 448 395 449 396 
<< pdiffusion >>
rect 449 395 450 396 
<< m1 >>
rect 64 396 65 397 
<< m1 >>
rect 82 396 83 397 
<< m1 >>
rect 85 396 86 397 
<< m1 >>
rect 109 396 110 397 
<< m1 >>
rect 124 396 125 397 
<< m1 >>
rect 127 396 128 397 
<< m1 >>
rect 145 396 146 397 
<< m1 >>
rect 172 396 173 397 
<< m1 >>
rect 289 396 290 397 
<< m2 >>
rect 290 396 291 397 
<< m1 >>
rect 301 396 302 397 
<< m1 >>
rect 64 397 65 398 
<< m1 >>
rect 82 397 83 398 
<< m1 >>
rect 83 397 84 398 
<< m1 >>
rect 84 397 85 398 
<< m1 >>
rect 85 397 86 398 
<< m1 >>
rect 109 397 110 398 
<< m1 >>
rect 124 397 125 398 
<< m1 >>
rect 127 397 128 398 
<< m1 >>
rect 145 397 146 398 
<< m1 >>
rect 172 397 173 398 
<< m1 >>
rect 289 397 290 398 
<< m2 >>
rect 290 397 291 398 
<< m1 >>
rect 291 397 292 398 
<< m2 >>
rect 291 397 292 398 
<< m2c >>
rect 291 397 292 398 
<< m1 >>
rect 291 397 292 398 
<< m2 >>
rect 291 397 292 398 
<< m1 >>
rect 292 397 293 398 
<< m1 >>
rect 293 397 294 398 
<< m1 >>
rect 294 397 295 398 
<< m1 >>
rect 295 397 296 398 
<< m1 >>
rect 296 397 297 398 
<< m1 >>
rect 297 397 298 398 
<< m1 >>
rect 298 397 299 398 
<< m1 >>
rect 299 397 300 398 
<< m1 >>
rect 300 397 301 398 
<< m1 >>
rect 301 397 302 398 
<< m1 >>
rect 64 398 65 399 
<< m1 >>
rect 109 398 110 399 
<< m1 >>
rect 124 398 125 399 
<< m1 >>
rect 127 398 128 399 
<< m1 >>
rect 145 398 146 399 
<< m1 >>
rect 172 398 173 399 
<< m1 >>
rect 289 398 290 399 
<< m1 >>
rect 64 399 65 400 
<< m1 >>
rect 109 399 110 400 
<< m1 >>
rect 124 399 125 400 
<< m1 >>
rect 127 399 128 400 
<< m1 >>
rect 145 399 146 400 
<< m1 >>
rect 172 399 173 400 
<< m1 >>
rect 289 399 290 400 
<< m1 >>
rect 64 400 65 401 
<< m1 >>
rect 109 400 110 401 
<< m1 >>
rect 110 400 111 401 
<< m1 >>
rect 111 400 112 401 
<< m1 >>
rect 112 400 113 401 
<< m1 >>
rect 113 400 114 401 
<< m1 >>
rect 114 400 115 401 
<< m1 >>
rect 115 400 116 401 
<< m1 >>
rect 116 400 117 401 
<< m1 >>
rect 117 400 118 401 
<< m1 >>
rect 118 400 119 401 
<< m1 >>
rect 119 400 120 401 
<< m1 >>
rect 120 400 121 401 
<< m1 >>
rect 121 400 122 401 
<< m1 >>
rect 122 400 123 401 
<< m1 >>
rect 123 400 124 401 
<< m1 >>
rect 124 400 125 401 
<< m1 >>
rect 127 400 128 401 
<< m2 >>
rect 127 400 128 401 
<< m2c >>
rect 127 400 128 401 
<< m1 >>
rect 127 400 128 401 
<< m2 >>
rect 127 400 128 401 
<< m1 >>
rect 145 400 146 401 
<< m1 >>
rect 172 400 173 401 
<< m1 >>
rect 289 400 290 401 
<< m1 >>
rect 64 401 65 402 
<< m2 >>
rect 127 401 128 402 
<< m1 >>
rect 145 401 146 402 
<< m1 >>
rect 172 401 173 402 
<< m1 >>
rect 289 401 290 402 
<< m1 >>
rect 64 402 65 403 
<< m1 >>
rect 121 402 122 403 
<< m1 >>
rect 122 402 123 403 
<< m1 >>
rect 123 402 124 403 
<< m1 >>
rect 124 402 125 403 
<< m1 >>
rect 125 402 126 403 
<< m1 >>
rect 126 402 127 403 
<< m1 >>
rect 127 402 128 403 
<< m2 >>
rect 127 402 128 403 
<< m1 >>
rect 128 402 129 403 
<< m1 >>
rect 129 402 130 403 
<< m1 >>
rect 130 402 131 403 
<< m1 >>
rect 131 402 132 403 
<< m1 >>
rect 132 402 133 403 
<< m1 >>
rect 133 402 134 403 
<< m1 >>
rect 134 402 135 403 
<< m1 >>
rect 135 402 136 403 
<< m1 >>
rect 136 402 137 403 
<< m1 >>
rect 137 402 138 403 
<< m1 >>
rect 138 402 139 403 
<< m1 >>
rect 139 402 140 403 
<< m1 >>
rect 140 402 141 403 
<< m1 >>
rect 141 402 142 403 
<< m1 >>
rect 142 402 143 403 
<< m1 >>
rect 143 402 144 403 
<< m1 >>
rect 144 402 145 403 
<< m1 >>
rect 145 402 146 403 
<< m1 >>
rect 172 402 173 403 
<< m1 >>
rect 289 402 290 403 
<< m1 >>
rect 64 403 65 404 
<< m1 >>
rect 121 403 122 404 
<< m2 >>
rect 127 403 128 404 
<< m1 >>
rect 172 403 173 404 
<< m1 >>
rect 173 403 174 404 
<< m1 >>
rect 174 403 175 404 
<< m1 >>
rect 175 403 176 404 
<< m1 >>
rect 176 403 177 404 
<< m1 >>
rect 177 403 178 404 
<< m1 >>
rect 178 403 179 404 
<< m1 >>
rect 179 403 180 404 
<< m1 >>
rect 180 403 181 404 
<< m1 >>
rect 181 403 182 404 
<< m1 >>
rect 182 403 183 404 
<< m1 >>
rect 183 403 184 404 
<< m1 >>
rect 184 403 185 404 
<< m1 >>
rect 185 403 186 404 
<< m1 >>
rect 186 403 187 404 
<< m1 >>
rect 187 403 188 404 
<< m1 >>
rect 188 403 189 404 
<< m1 >>
rect 189 403 190 404 
<< m1 >>
rect 190 403 191 404 
<< m1 >>
rect 191 403 192 404 
<< m1 >>
rect 192 403 193 404 
<< m1 >>
rect 193 403 194 404 
<< m1 >>
rect 194 403 195 404 
<< m1 >>
rect 195 403 196 404 
<< m1 >>
rect 196 403 197 404 
<< m1 >>
rect 289 403 290 404 
<< m1 >>
rect 64 404 65 405 
<< m1 >>
rect 121 404 122 405 
<< m1 >>
rect 127 404 128 405 
<< m2 >>
rect 127 404 128 405 
<< m2c >>
rect 127 404 128 405 
<< m1 >>
rect 127 404 128 405 
<< m2 >>
rect 127 404 128 405 
<< m1 >>
rect 196 404 197 405 
<< m1 >>
rect 289 404 290 405 
<< m1 >>
rect 49 405 50 406 
<< m1 >>
rect 50 405 51 406 
<< m1 >>
rect 51 405 52 406 
<< m1 >>
rect 52 405 53 406 
<< m1 >>
rect 53 405 54 406 
<< m1 >>
rect 54 405 55 406 
<< m1 >>
rect 55 405 56 406 
<< m1 >>
rect 56 405 57 406 
<< m1 >>
rect 57 405 58 406 
<< m1 >>
rect 58 405 59 406 
<< m1 >>
rect 59 405 60 406 
<< m1 >>
rect 60 405 61 406 
<< m1 >>
rect 61 405 62 406 
<< m1 >>
rect 62 405 63 406 
<< m2 >>
rect 62 405 63 406 
<< m2c >>
rect 62 405 63 406 
<< m1 >>
rect 62 405 63 406 
<< m2 >>
rect 62 405 63 406 
<< m2 >>
rect 63 405 64 406 
<< m1 >>
rect 64 405 65 406 
<< m2 >>
rect 64 405 65 406 
<< m2 >>
rect 65 405 66 406 
<< m1 >>
rect 66 405 67 406 
<< m2 >>
rect 66 405 67 406 
<< m2c >>
rect 66 405 67 406 
<< m1 >>
rect 66 405 67 406 
<< m2 >>
rect 66 405 67 406 
<< m1 >>
rect 67 405 68 406 
<< m1 >>
rect 121 405 122 406 
<< m1 >>
rect 127 405 128 406 
<< m1 >>
rect 196 405 197 406 
<< m1 >>
rect 289 405 290 406 
<< m1 >>
rect 49 406 50 407 
<< m1 >>
rect 64 406 65 407 
<< m1 >>
rect 67 406 68 407 
<< m1 >>
rect 121 406 122 407 
<< m1 >>
rect 127 406 128 407 
<< m1 >>
rect 196 406 197 407 
<< m1 >>
rect 289 406 290 407 
<< m1 >>
rect 49 407 50 408 
<< m1 >>
rect 64 407 65 408 
<< m1 >>
rect 67 407 68 408 
<< m1 >>
rect 121 407 122 408 
<< m1 >>
rect 127 407 128 408 
<< m1 >>
rect 196 407 197 408 
<< m1 >>
rect 289 407 290 408 
<< pdiffusion >>
rect 12 408 13 409 
<< pdiffusion >>
rect 13 408 14 409 
<< pdiffusion >>
rect 14 408 15 409 
<< pdiffusion >>
rect 15 408 16 409 
<< pdiffusion >>
rect 16 408 17 409 
<< pdiffusion >>
rect 17 408 18 409 
<< pdiffusion >>
rect 30 408 31 409 
<< pdiffusion >>
rect 31 408 32 409 
<< pdiffusion >>
rect 32 408 33 409 
<< pdiffusion >>
rect 33 408 34 409 
<< pdiffusion >>
rect 34 408 35 409 
<< pdiffusion >>
rect 35 408 36 409 
<< pdiffusion >>
rect 48 408 49 409 
<< m1 >>
rect 49 408 50 409 
<< pdiffusion >>
rect 49 408 50 409 
<< pdiffusion >>
rect 50 408 51 409 
<< pdiffusion >>
rect 51 408 52 409 
<< pdiffusion >>
rect 52 408 53 409 
<< pdiffusion >>
rect 53 408 54 409 
<< m1 >>
rect 64 408 65 409 
<< pdiffusion >>
rect 66 408 67 409 
<< m1 >>
rect 67 408 68 409 
<< pdiffusion >>
rect 67 408 68 409 
<< pdiffusion >>
rect 68 408 69 409 
<< pdiffusion >>
rect 69 408 70 409 
<< pdiffusion >>
rect 70 408 71 409 
<< pdiffusion >>
rect 71 408 72 409 
<< pdiffusion >>
rect 84 408 85 409 
<< pdiffusion >>
rect 85 408 86 409 
<< pdiffusion >>
rect 86 408 87 409 
<< pdiffusion >>
rect 87 408 88 409 
<< pdiffusion >>
rect 88 408 89 409 
<< pdiffusion >>
rect 89 408 90 409 
<< pdiffusion >>
rect 102 408 103 409 
<< pdiffusion >>
rect 103 408 104 409 
<< pdiffusion >>
rect 104 408 105 409 
<< pdiffusion >>
rect 105 408 106 409 
<< pdiffusion >>
rect 106 408 107 409 
<< pdiffusion >>
rect 107 408 108 409 
<< pdiffusion >>
rect 120 408 121 409 
<< m1 >>
rect 121 408 122 409 
<< pdiffusion >>
rect 121 408 122 409 
<< pdiffusion >>
rect 122 408 123 409 
<< pdiffusion >>
rect 123 408 124 409 
<< pdiffusion >>
rect 124 408 125 409 
<< pdiffusion >>
rect 125 408 126 409 
<< m1 >>
rect 127 408 128 409 
<< pdiffusion >>
rect 138 408 139 409 
<< pdiffusion >>
rect 139 408 140 409 
<< pdiffusion >>
rect 140 408 141 409 
<< pdiffusion >>
rect 141 408 142 409 
<< pdiffusion >>
rect 142 408 143 409 
<< pdiffusion >>
rect 143 408 144 409 
<< pdiffusion >>
rect 156 408 157 409 
<< pdiffusion >>
rect 157 408 158 409 
<< pdiffusion >>
rect 158 408 159 409 
<< pdiffusion >>
rect 159 408 160 409 
<< pdiffusion >>
rect 160 408 161 409 
<< pdiffusion >>
rect 161 408 162 409 
<< pdiffusion >>
rect 174 408 175 409 
<< pdiffusion >>
rect 175 408 176 409 
<< pdiffusion >>
rect 176 408 177 409 
<< pdiffusion >>
rect 177 408 178 409 
<< pdiffusion >>
rect 178 408 179 409 
<< pdiffusion >>
rect 179 408 180 409 
<< pdiffusion >>
rect 192 408 193 409 
<< pdiffusion >>
rect 193 408 194 409 
<< pdiffusion >>
rect 194 408 195 409 
<< pdiffusion >>
rect 195 408 196 409 
<< m1 >>
rect 196 408 197 409 
<< pdiffusion >>
rect 196 408 197 409 
<< pdiffusion >>
rect 197 408 198 409 
<< pdiffusion >>
rect 210 408 211 409 
<< pdiffusion >>
rect 211 408 212 409 
<< pdiffusion >>
rect 212 408 213 409 
<< pdiffusion >>
rect 213 408 214 409 
<< pdiffusion >>
rect 214 408 215 409 
<< pdiffusion >>
rect 215 408 216 409 
<< pdiffusion >>
rect 228 408 229 409 
<< pdiffusion >>
rect 229 408 230 409 
<< pdiffusion >>
rect 230 408 231 409 
<< pdiffusion >>
rect 231 408 232 409 
<< pdiffusion >>
rect 232 408 233 409 
<< pdiffusion >>
rect 233 408 234 409 
<< pdiffusion >>
rect 246 408 247 409 
<< pdiffusion >>
rect 247 408 248 409 
<< pdiffusion >>
rect 248 408 249 409 
<< pdiffusion >>
rect 249 408 250 409 
<< pdiffusion >>
rect 250 408 251 409 
<< pdiffusion >>
rect 251 408 252 409 
<< pdiffusion >>
rect 264 408 265 409 
<< pdiffusion >>
rect 265 408 266 409 
<< pdiffusion >>
rect 266 408 267 409 
<< pdiffusion >>
rect 267 408 268 409 
<< pdiffusion >>
rect 268 408 269 409 
<< pdiffusion >>
rect 269 408 270 409 
<< pdiffusion >>
rect 282 408 283 409 
<< pdiffusion >>
rect 283 408 284 409 
<< pdiffusion >>
rect 284 408 285 409 
<< pdiffusion >>
rect 285 408 286 409 
<< pdiffusion >>
rect 286 408 287 409 
<< pdiffusion >>
rect 287 408 288 409 
<< m1 >>
rect 289 408 290 409 
<< pdiffusion >>
rect 300 408 301 409 
<< pdiffusion >>
rect 301 408 302 409 
<< pdiffusion >>
rect 302 408 303 409 
<< pdiffusion >>
rect 303 408 304 409 
<< pdiffusion >>
rect 304 408 305 409 
<< pdiffusion >>
rect 305 408 306 409 
<< pdiffusion >>
rect 336 408 337 409 
<< pdiffusion >>
rect 337 408 338 409 
<< pdiffusion >>
rect 338 408 339 409 
<< pdiffusion >>
rect 339 408 340 409 
<< pdiffusion >>
rect 340 408 341 409 
<< pdiffusion >>
rect 341 408 342 409 
<< pdiffusion >>
rect 354 408 355 409 
<< pdiffusion >>
rect 355 408 356 409 
<< pdiffusion >>
rect 356 408 357 409 
<< pdiffusion >>
rect 357 408 358 409 
<< pdiffusion >>
rect 358 408 359 409 
<< pdiffusion >>
rect 359 408 360 409 
<< pdiffusion >>
rect 372 408 373 409 
<< pdiffusion >>
rect 373 408 374 409 
<< pdiffusion >>
rect 374 408 375 409 
<< pdiffusion >>
rect 375 408 376 409 
<< pdiffusion >>
rect 376 408 377 409 
<< pdiffusion >>
rect 377 408 378 409 
<< pdiffusion >>
rect 390 408 391 409 
<< pdiffusion >>
rect 391 408 392 409 
<< pdiffusion >>
rect 392 408 393 409 
<< pdiffusion >>
rect 393 408 394 409 
<< pdiffusion >>
rect 394 408 395 409 
<< pdiffusion >>
rect 395 408 396 409 
<< pdiffusion >>
rect 408 408 409 409 
<< pdiffusion >>
rect 409 408 410 409 
<< pdiffusion >>
rect 410 408 411 409 
<< pdiffusion >>
rect 411 408 412 409 
<< pdiffusion >>
rect 412 408 413 409 
<< pdiffusion >>
rect 413 408 414 409 
<< pdiffusion >>
rect 426 408 427 409 
<< pdiffusion >>
rect 427 408 428 409 
<< pdiffusion >>
rect 428 408 429 409 
<< pdiffusion >>
rect 429 408 430 409 
<< pdiffusion >>
rect 430 408 431 409 
<< pdiffusion >>
rect 431 408 432 409 
<< pdiffusion >>
rect 444 408 445 409 
<< pdiffusion >>
rect 445 408 446 409 
<< pdiffusion >>
rect 446 408 447 409 
<< pdiffusion >>
rect 447 408 448 409 
<< pdiffusion >>
rect 448 408 449 409 
<< pdiffusion >>
rect 449 408 450 409 
<< pdiffusion >>
rect 12 409 13 410 
<< pdiffusion >>
rect 13 409 14 410 
<< pdiffusion >>
rect 14 409 15 410 
<< pdiffusion >>
rect 15 409 16 410 
<< pdiffusion >>
rect 16 409 17 410 
<< pdiffusion >>
rect 17 409 18 410 
<< pdiffusion >>
rect 30 409 31 410 
<< pdiffusion >>
rect 31 409 32 410 
<< pdiffusion >>
rect 32 409 33 410 
<< pdiffusion >>
rect 33 409 34 410 
<< pdiffusion >>
rect 34 409 35 410 
<< pdiffusion >>
rect 35 409 36 410 
<< pdiffusion >>
rect 48 409 49 410 
<< pdiffusion >>
rect 49 409 50 410 
<< pdiffusion >>
rect 50 409 51 410 
<< pdiffusion >>
rect 51 409 52 410 
<< pdiffusion >>
rect 52 409 53 410 
<< pdiffusion >>
rect 53 409 54 410 
<< m1 >>
rect 64 409 65 410 
<< pdiffusion >>
rect 66 409 67 410 
<< pdiffusion >>
rect 67 409 68 410 
<< pdiffusion >>
rect 68 409 69 410 
<< pdiffusion >>
rect 69 409 70 410 
<< pdiffusion >>
rect 70 409 71 410 
<< pdiffusion >>
rect 71 409 72 410 
<< pdiffusion >>
rect 84 409 85 410 
<< pdiffusion >>
rect 85 409 86 410 
<< pdiffusion >>
rect 86 409 87 410 
<< pdiffusion >>
rect 87 409 88 410 
<< pdiffusion >>
rect 88 409 89 410 
<< pdiffusion >>
rect 89 409 90 410 
<< pdiffusion >>
rect 102 409 103 410 
<< pdiffusion >>
rect 103 409 104 410 
<< pdiffusion >>
rect 104 409 105 410 
<< pdiffusion >>
rect 105 409 106 410 
<< pdiffusion >>
rect 106 409 107 410 
<< pdiffusion >>
rect 107 409 108 410 
<< pdiffusion >>
rect 120 409 121 410 
<< pdiffusion >>
rect 121 409 122 410 
<< pdiffusion >>
rect 122 409 123 410 
<< pdiffusion >>
rect 123 409 124 410 
<< pdiffusion >>
rect 124 409 125 410 
<< pdiffusion >>
rect 125 409 126 410 
<< m1 >>
rect 127 409 128 410 
<< pdiffusion >>
rect 138 409 139 410 
<< pdiffusion >>
rect 139 409 140 410 
<< pdiffusion >>
rect 140 409 141 410 
<< pdiffusion >>
rect 141 409 142 410 
<< pdiffusion >>
rect 142 409 143 410 
<< pdiffusion >>
rect 143 409 144 410 
<< pdiffusion >>
rect 156 409 157 410 
<< pdiffusion >>
rect 157 409 158 410 
<< pdiffusion >>
rect 158 409 159 410 
<< pdiffusion >>
rect 159 409 160 410 
<< pdiffusion >>
rect 160 409 161 410 
<< pdiffusion >>
rect 161 409 162 410 
<< pdiffusion >>
rect 174 409 175 410 
<< pdiffusion >>
rect 175 409 176 410 
<< pdiffusion >>
rect 176 409 177 410 
<< pdiffusion >>
rect 177 409 178 410 
<< pdiffusion >>
rect 178 409 179 410 
<< pdiffusion >>
rect 179 409 180 410 
<< pdiffusion >>
rect 192 409 193 410 
<< pdiffusion >>
rect 193 409 194 410 
<< pdiffusion >>
rect 194 409 195 410 
<< pdiffusion >>
rect 195 409 196 410 
<< pdiffusion >>
rect 196 409 197 410 
<< pdiffusion >>
rect 197 409 198 410 
<< pdiffusion >>
rect 210 409 211 410 
<< pdiffusion >>
rect 211 409 212 410 
<< pdiffusion >>
rect 212 409 213 410 
<< pdiffusion >>
rect 213 409 214 410 
<< pdiffusion >>
rect 214 409 215 410 
<< pdiffusion >>
rect 215 409 216 410 
<< pdiffusion >>
rect 228 409 229 410 
<< pdiffusion >>
rect 229 409 230 410 
<< pdiffusion >>
rect 230 409 231 410 
<< pdiffusion >>
rect 231 409 232 410 
<< pdiffusion >>
rect 232 409 233 410 
<< pdiffusion >>
rect 233 409 234 410 
<< pdiffusion >>
rect 246 409 247 410 
<< pdiffusion >>
rect 247 409 248 410 
<< pdiffusion >>
rect 248 409 249 410 
<< pdiffusion >>
rect 249 409 250 410 
<< pdiffusion >>
rect 250 409 251 410 
<< pdiffusion >>
rect 251 409 252 410 
<< pdiffusion >>
rect 264 409 265 410 
<< pdiffusion >>
rect 265 409 266 410 
<< pdiffusion >>
rect 266 409 267 410 
<< pdiffusion >>
rect 267 409 268 410 
<< pdiffusion >>
rect 268 409 269 410 
<< pdiffusion >>
rect 269 409 270 410 
<< pdiffusion >>
rect 282 409 283 410 
<< pdiffusion >>
rect 283 409 284 410 
<< pdiffusion >>
rect 284 409 285 410 
<< pdiffusion >>
rect 285 409 286 410 
<< pdiffusion >>
rect 286 409 287 410 
<< pdiffusion >>
rect 287 409 288 410 
<< m1 >>
rect 289 409 290 410 
<< pdiffusion >>
rect 300 409 301 410 
<< pdiffusion >>
rect 301 409 302 410 
<< pdiffusion >>
rect 302 409 303 410 
<< pdiffusion >>
rect 303 409 304 410 
<< pdiffusion >>
rect 304 409 305 410 
<< pdiffusion >>
rect 305 409 306 410 
<< pdiffusion >>
rect 336 409 337 410 
<< pdiffusion >>
rect 337 409 338 410 
<< pdiffusion >>
rect 338 409 339 410 
<< pdiffusion >>
rect 339 409 340 410 
<< pdiffusion >>
rect 340 409 341 410 
<< pdiffusion >>
rect 341 409 342 410 
<< pdiffusion >>
rect 354 409 355 410 
<< pdiffusion >>
rect 355 409 356 410 
<< pdiffusion >>
rect 356 409 357 410 
<< pdiffusion >>
rect 357 409 358 410 
<< pdiffusion >>
rect 358 409 359 410 
<< pdiffusion >>
rect 359 409 360 410 
<< pdiffusion >>
rect 372 409 373 410 
<< pdiffusion >>
rect 373 409 374 410 
<< pdiffusion >>
rect 374 409 375 410 
<< pdiffusion >>
rect 375 409 376 410 
<< pdiffusion >>
rect 376 409 377 410 
<< pdiffusion >>
rect 377 409 378 410 
<< pdiffusion >>
rect 390 409 391 410 
<< pdiffusion >>
rect 391 409 392 410 
<< pdiffusion >>
rect 392 409 393 410 
<< pdiffusion >>
rect 393 409 394 410 
<< pdiffusion >>
rect 394 409 395 410 
<< pdiffusion >>
rect 395 409 396 410 
<< pdiffusion >>
rect 408 409 409 410 
<< pdiffusion >>
rect 409 409 410 410 
<< pdiffusion >>
rect 410 409 411 410 
<< pdiffusion >>
rect 411 409 412 410 
<< pdiffusion >>
rect 412 409 413 410 
<< pdiffusion >>
rect 413 409 414 410 
<< pdiffusion >>
rect 426 409 427 410 
<< pdiffusion >>
rect 427 409 428 410 
<< pdiffusion >>
rect 428 409 429 410 
<< pdiffusion >>
rect 429 409 430 410 
<< pdiffusion >>
rect 430 409 431 410 
<< pdiffusion >>
rect 431 409 432 410 
<< pdiffusion >>
rect 444 409 445 410 
<< pdiffusion >>
rect 445 409 446 410 
<< pdiffusion >>
rect 446 409 447 410 
<< pdiffusion >>
rect 447 409 448 410 
<< pdiffusion >>
rect 448 409 449 410 
<< pdiffusion >>
rect 449 409 450 410 
<< pdiffusion >>
rect 12 410 13 411 
<< pdiffusion >>
rect 13 410 14 411 
<< pdiffusion >>
rect 14 410 15 411 
<< pdiffusion >>
rect 15 410 16 411 
<< pdiffusion >>
rect 16 410 17 411 
<< pdiffusion >>
rect 17 410 18 411 
<< pdiffusion >>
rect 30 410 31 411 
<< pdiffusion >>
rect 31 410 32 411 
<< pdiffusion >>
rect 32 410 33 411 
<< pdiffusion >>
rect 33 410 34 411 
<< pdiffusion >>
rect 34 410 35 411 
<< pdiffusion >>
rect 35 410 36 411 
<< pdiffusion >>
rect 48 410 49 411 
<< pdiffusion >>
rect 49 410 50 411 
<< pdiffusion >>
rect 50 410 51 411 
<< pdiffusion >>
rect 51 410 52 411 
<< pdiffusion >>
rect 52 410 53 411 
<< pdiffusion >>
rect 53 410 54 411 
<< m1 >>
rect 64 410 65 411 
<< pdiffusion >>
rect 66 410 67 411 
<< pdiffusion >>
rect 67 410 68 411 
<< pdiffusion >>
rect 68 410 69 411 
<< pdiffusion >>
rect 69 410 70 411 
<< pdiffusion >>
rect 70 410 71 411 
<< pdiffusion >>
rect 71 410 72 411 
<< pdiffusion >>
rect 84 410 85 411 
<< pdiffusion >>
rect 85 410 86 411 
<< pdiffusion >>
rect 86 410 87 411 
<< pdiffusion >>
rect 87 410 88 411 
<< pdiffusion >>
rect 88 410 89 411 
<< pdiffusion >>
rect 89 410 90 411 
<< pdiffusion >>
rect 102 410 103 411 
<< pdiffusion >>
rect 103 410 104 411 
<< pdiffusion >>
rect 104 410 105 411 
<< pdiffusion >>
rect 105 410 106 411 
<< pdiffusion >>
rect 106 410 107 411 
<< pdiffusion >>
rect 107 410 108 411 
<< pdiffusion >>
rect 120 410 121 411 
<< pdiffusion >>
rect 121 410 122 411 
<< pdiffusion >>
rect 122 410 123 411 
<< pdiffusion >>
rect 123 410 124 411 
<< pdiffusion >>
rect 124 410 125 411 
<< pdiffusion >>
rect 125 410 126 411 
<< m1 >>
rect 127 410 128 411 
<< pdiffusion >>
rect 138 410 139 411 
<< pdiffusion >>
rect 139 410 140 411 
<< pdiffusion >>
rect 140 410 141 411 
<< pdiffusion >>
rect 141 410 142 411 
<< pdiffusion >>
rect 142 410 143 411 
<< pdiffusion >>
rect 143 410 144 411 
<< pdiffusion >>
rect 156 410 157 411 
<< pdiffusion >>
rect 157 410 158 411 
<< pdiffusion >>
rect 158 410 159 411 
<< pdiffusion >>
rect 159 410 160 411 
<< pdiffusion >>
rect 160 410 161 411 
<< pdiffusion >>
rect 161 410 162 411 
<< pdiffusion >>
rect 174 410 175 411 
<< pdiffusion >>
rect 175 410 176 411 
<< pdiffusion >>
rect 176 410 177 411 
<< pdiffusion >>
rect 177 410 178 411 
<< pdiffusion >>
rect 178 410 179 411 
<< pdiffusion >>
rect 179 410 180 411 
<< pdiffusion >>
rect 192 410 193 411 
<< pdiffusion >>
rect 193 410 194 411 
<< pdiffusion >>
rect 194 410 195 411 
<< pdiffusion >>
rect 195 410 196 411 
<< pdiffusion >>
rect 196 410 197 411 
<< pdiffusion >>
rect 197 410 198 411 
<< pdiffusion >>
rect 210 410 211 411 
<< pdiffusion >>
rect 211 410 212 411 
<< pdiffusion >>
rect 212 410 213 411 
<< pdiffusion >>
rect 213 410 214 411 
<< pdiffusion >>
rect 214 410 215 411 
<< pdiffusion >>
rect 215 410 216 411 
<< pdiffusion >>
rect 228 410 229 411 
<< pdiffusion >>
rect 229 410 230 411 
<< pdiffusion >>
rect 230 410 231 411 
<< pdiffusion >>
rect 231 410 232 411 
<< pdiffusion >>
rect 232 410 233 411 
<< pdiffusion >>
rect 233 410 234 411 
<< pdiffusion >>
rect 246 410 247 411 
<< pdiffusion >>
rect 247 410 248 411 
<< pdiffusion >>
rect 248 410 249 411 
<< pdiffusion >>
rect 249 410 250 411 
<< pdiffusion >>
rect 250 410 251 411 
<< pdiffusion >>
rect 251 410 252 411 
<< pdiffusion >>
rect 264 410 265 411 
<< pdiffusion >>
rect 265 410 266 411 
<< pdiffusion >>
rect 266 410 267 411 
<< pdiffusion >>
rect 267 410 268 411 
<< pdiffusion >>
rect 268 410 269 411 
<< pdiffusion >>
rect 269 410 270 411 
<< pdiffusion >>
rect 282 410 283 411 
<< pdiffusion >>
rect 283 410 284 411 
<< pdiffusion >>
rect 284 410 285 411 
<< pdiffusion >>
rect 285 410 286 411 
<< pdiffusion >>
rect 286 410 287 411 
<< pdiffusion >>
rect 287 410 288 411 
<< m1 >>
rect 289 410 290 411 
<< pdiffusion >>
rect 300 410 301 411 
<< pdiffusion >>
rect 301 410 302 411 
<< pdiffusion >>
rect 302 410 303 411 
<< pdiffusion >>
rect 303 410 304 411 
<< pdiffusion >>
rect 304 410 305 411 
<< pdiffusion >>
rect 305 410 306 411 
<< pdiffusion >>
rect 336 410 337 411 
<< pdiffusion >>
rect 337 410 338 411 
<< pdiffusion >>
rect 338 410 339 411 
<< pdiffusion >>
rect 339 410 340 411 
<< pdiffusion >>
rect 340 410 341 411 
<< pdiffusion >>
rect 341 410 342 411 
<< pdiffusion >>
rect 354 410 355 411 
<< pdiffusion >>
rect 355 410 356 411 
<< pdiffusion >>
rect 356 410 357 411 
<< pdiffusion >>
rect 357 410 358 411 
<< pdiffusion >>
rect 358 410 359 411 
<< pdiffusion >>
rect 359 410 360 411 
<< pdiffusion >>
rect 372 410 373 411 
<< pdiffusion >>
rect 373 410 374 411 
<< pdiffusion >>
rect 374 410 375 411 
<< pdiffusion >>
rect 375 410 376 411 
<< pdiffusion >>
rect 376 410 377 411 
<< pdiffusion >>
rect 377 410 378 411 
<< pdiffusion >>
rect 390 410 391 411 
<< pdiffusion >>
rect 391 410 392 411 
<< pdiffusion >>
rect 392 410 393 411 
<< pdiffusion >>
rect 393 410 394 411 
<< pdiffusion >>
rect 394 410 395 411 
<< pdiffusion >>
rect 395 410 396 411 
<< pdiffusion >>
rect 408 410 409 411 
<< pdiffusion >>
rect 409 410 410 411 
<< pdiffusion >>
rect 410 410 411 411 
<< pdiffusion >>
rect 411 410 412 411 
<< pdiffusion >>
rect 412 410 413 411 
<< pdiffusion >>
rect 413 410 414 411 
<< pdiffusion >>
rect 426 410 427 411 
<< pdiffusion >>
rect 427 410 428 411 
<< pdiffusion >>
rect 428 410 429 411 
<< pdiffusion >>
rect 429 410 430 411 
<< pdiffusion >>
rect 430 410 431 411 
<< pdiffusion >>
rect 431 410 432 411 
<< pdiffusion >>
rect 444 410 445 411 
<< pdiffusion >>
rect 445 410 446 411 
<< pdiffusion >>
rect 446 410 447 411 
<< pdiffusion >>
rect 447 410 448 411 
<< pdiffusion >>
rect 448 410 449 411 
<< pdiffusion >>
rect 449 410 450 411 
<< pdiffusion >>
rect 12 411 13 412 
<< pdiffusion >>
rect 13 411 14 412 
<< pdiffusion >>
rect 14 411 15 412 
<< pdiffusion >>
rect 15 411 16 412 
<< pdiffusion >>
rect 16 411 17 412 
<< pdiffusion >>
rect 17 411 18 412 
<< pdiffusion >>
rect 30 411 31 412 
<< pdiffusion >>
rect 31 411 32 412 
<< pdiffusion >>
rect 32 411 33 412 
<< pdiffusion >>
rect 33 411 34 412 
<< pdiffusion >>
rect 34 411 35 412 
<< pdiffusion >>
rect 35 411 36 412 
<< pdiffusion >>
rect 48 411 49 412 
<< pdiffusion >>
rect 49 411 50 412 
<< pdiffusion >>
rect 50 411 51 412 
<< pdiffusion >>
rect 51 411 52 412 
<< pdiffusion >>
rect 52 411 53 412 
<< pdiffusion >>
rect 53 411 54 412 
<< m1 >>
rect 64 411 65 412 
<< pdiffusion >>
rect 66 411 67 412 
<< pdiffusion >>
rect 67 411 68 412 
<< pdiffusion >>
rect 68 411 69 412 
<< pdiffusion >>
rect 69 411 70 412 
<< pdiffusion >>
rect 70 411 71 412 
<< pdiffusion >>
rect 71 411 72 412 
<< pdiffusion >>
rect 84 411 85 412 
<< pdiffusion >>
rect 85 411 86 412 
<< pdiffusion >>
rect 86 411 87 412 
<< pdiffusion >>
rect 87 411 88 412 
<< pdiffusion >>
rect 88 411 89 412 
<< pdiffusion >>
rect 89 411 90 412 
<< pdiffusion >>
rect 102 411 103 412 
<< pdiffusion >>
rect 103 411 104 412 
<< pdiffusion >>
rect 104 411 105 412 
<< pdiffusion >>
rect 105 411 106 412 
<< pdiffusion >>
rect 106 411 107 412 
<< pdiffusion >>
rect 107 411 108 412 
<< pdiffusion >>
rect 120 411 121 412 
<< pdiffusion >>
rect 121 411 122 412 
<< pdiffusion >>
rect 122 411 123 412 
<< pdiffusion >>
rect 123 411 124 412 
<< pdiffusion >>
rect 124 411 125 412 
<< pdiffusion >>
rect 125 411 126 412 
<< m1 >>
rect 127 411 128 412 
<< pdiffusion >>
rect 138 411 139 412 
<< pdiffusion >>
rect 139 411 140 412 
<< pdiffusion >>
rect 140 411 141 412 
<< pdiffusion >>
rect 141 411 142 412 
<< pdiffusion >>
rect 142 411 143 412 
<< pdiffusion >>
rect 143 411 144 412 
<< pdiffusion >>
rect 156 411 157 412 
<< pdiffusion >>
rect 157 411 158 412 
<< pdiffusion >>
rect 158 411 159 412 
<< pdiffusion >>
rect 159 411 160 412 
<< pdiffusion >>
rect 160 411 161 412 
<< pdiffusion >>
rect 161 411 162 412 
<< pdiffusion >>
rect 174 411 175 412 
<< pdiffusion >>
rect 175 411 176 412 
<< pdiffusion >>
rect 176 411 177 412 
<< pdiffusion >>
rect 177 411 178 412 
<< pdiffusion >>
rect 178 411 179 412 
<< pdiffusion >>
rect 179 411 180 412 
<< pdiffusion >>
rect 192 411 193 412 
<< pdiffusion >>
rect 193 411 194 412 
<< pdiffusion >>
rect 194 411 195 412 
<< pdiffusion >>
rect 195 411 196 412 
<< pdiffusion >>
rect 196 411 197 412 
<< pdiffusion >>
rect 197 411 198 412 
<< pdiffusion >>
rect 210 411 211 412 
<< pdiffusion >>
rect 211 411 212 412 
<< pdiffusion >>
rect 212 411 213 412 
<< pdiffusion >>
rect 213 411 214 412 
<< pdiffusion >>
rect 214 411 215 412 
<< pdiffusion >>
rect 215 411 216 412 
<< pdiffusion >>
rect 228 411 229 412 
<< pdiffusion >>
rect 229 411 230 412 
<< pdiffusion >>
rect 230 411 231 412 
<< pdiffusion >>
rect 231 411 232 412 
<< pdiffusion >>
rect 232 411 233 412 
<< pdiffusion >>
rect 233 411 234 412 
<< pdiffusion >>
rect 246 411 247 412 
<< pdiffusion >>
rect 247 411 248 412 
<< pdiffusion >>
rect 248 411 249 412 
<< pdiffusion >>
rect 249 411 250 412 
<< pdiffusion >>
rect 250 411 251 412 
<< pdiffusion >>
rect 251 411 252 412 
<< pdiffusion >>
rect 264 411 265 412 
<< pdiffusion >>
rect 265 411 266 412 
<< pdiffusion >>
rect 266 411 267 412 
<< pdiffusion >>
rect 267 411 268 412 
<< pdiffusion >>
rect 268 411 269 412 
<< pdiffusion >>
rect 269 411 270 412 
<< pdiffusion >>
rect 282 411 283 412 
<< pdiffusion >>
rect 283 411 284 412 
<< pdiffusion >>
rect 284 411 285 412 
<< pdiffusion >>
rect 285 411 286 412 
<< pdiffusion >>
rect 286 411 287 412 
<< pdiffusion >>
rect 287 411 288 412 
<< m1 >>
rect 289 411 290 412 
<< pdiffusion >>
rect 300 411 301 412 
<< pdiffusion >>
rect 301 411 302 412 
<< pdiffusion >>
rect 302 411 303 412 
<< pdiffusion >>
rect 303 411 304 412 
<< pdiffusion >>
rect 304 411 305 412 
<< pdiffusion >>
rect 305 411 306 412 
<< pdiffusion >>
rect 336 411 337 412 
<< pdiffusion >>
rect 337 411 338 412 
<< pdiffusion >>
rect 338 411 339 412 
<< pdiffusion >>
rect 339 411 340 412 
<< pdiffusion >>
rect 340 411 341 412 
<< pdiffusion >>
rect 341 411 342 412 
<< pdiffusion >>
rect 354 411 355 412 
<< pdiffusion >>
rect 355 411 356 412 
<< pdiffusion >>
rect 356 411 357 412 
<< pdiffusion >>
rect 357 411 358 412 
<< pdiffusion >>
rect 358 411 359 412 
<< pdiffusion >>
rect 359 411 360 412 
<< pdiffusion >>
rect 372 411 373 412 
<< pdiffusion >>
rect 373 411 374 412 
<< pdiffusion >>
rect 374 411 375 412 
<< pdiffusion >>
rect 375 411 376 412 
<< pdiffusion >>
rect 376 411 377 412 
<< pdiffusion >>
rect 377 411 378 412 
<< pdiffusion >>
rect 390 411 391 412 
<< pdiffusion >>
rect 391 411 392 412 
<< pdiffusion >>
rect 392 411 393 412 
<< pdiffusion >>
rect 393 411 394 412 
<< pdiffusion >>
rect 394 411 395 412 
<< pdiffusion >>
rect 395 411 396 412 
<< pdiffusion >>
rect 408 411 409 412 
<< pdiffusion >>
rect 409 411 410 412 
<< pdiffusion >>
rect 410 411 411 412 
<< pdiffusion >>
rect 411 411 412 412 
<< pdiffusion >>
rect 412 411 413 412 
<< pdiffusion >>
rect 413 411 414 412 
<< pdiffusion >>
rect 426 411 427 412 
<< pdiffusion >>
rect 427 411 428 412 
<< pdiffusion >>
rect 428 411 429 412 
<< pdiffusion >>
rect 429 411 430 412 
<< pdiffusion >>
rect 430 411 431 412 
<< pdiffusion >>
rect 431 411 432 412 
<< pdiffusion >>
rect 444 411 445 412 
<< pdiffusion >>
rect 445 411 446 412 
<< pdiffusion >>
rect 446 411 447 412 
<< pdiffusion >>
rect 447 411 448 412 
<< pdiffusion >>
rect 448 411 449 412 
<< pdiffusion >>
rect 449 411 450 412 
<< pdiffusion >>
rect 12 412 13 413 
<< pdiffusion >>
rect 13 412 14 413 
<< pdiffusion >>
rect 14 412 15 413 
<< pdiffusion >>
rect 15 412 16 413 
<< pdiffusion >>
rect 16 412 17 413 
<< pdiffusion >>
rect 17 412 18 413 
<< pdiffusion >>
rect 30 412 31 413 
<< pdiffusion >>
rect 31 412 32 413 
<< pdiffusion >>
rect 32 412 33 413 
<< pdiffusion >>
rect 33 412 34 413 
<< pdiffusion >>
rect 34 412 35 413 
<< pdiffusion >>
rect 35 412 36 413 
<< pdiffusion >>
rect 48 412 49 413 
<< pdiffusion >>
rect 49 412 50 413 
<< pdiffusion >>
rect 50 412 51 413 
<< pdiffusion >>
rect 51 412 52 413 
<< pdiffusion >>
rect 52 412 53 413 
<< pdiffusion >>
rect 53 412 54 413 
<< m1 >>
rect 64 412 65 413 
<< pdiffusion >>
rect 66 412 67 413 
<< pdiffusion >>
rect 67 412 68 413 
<< pdiffusion >>
rect 68 412 69 413 
<< pdiffusion >>
rect 69 412 70 413 
<< pdiffusion >>
rect 70 412 71 413 
<< pdiffusion >>
rect 71 412 72 413 
<< pdiffusion >>
rect 84 412 85 413 
<< pdiffusion >>
rect 85 412 86 413 
<< pdiffusion >>
rect 86 412 87 413 
<< pdiffusion >>
rect 87 412 88 413 
<< pdiffusion >>
rect 88 412 89 413 
<< pdiffusion >>
rect 89 412 90 413 
<< pdiffusion >>
rect 102 412 103 413 
<< pdiffusion >>
rect 103 412 104 413 
<< pdiffusion >>
rect 104 412 105 413 
<< pdiffusion >>
rect 105 412 106 413 
<< pdiffusion >>
rect 106 412 107 413 
<< pdiffusion >>
rect 107 412 108 413 
<< pdiffusion >>
rect 120 412 121 413 
<< pdiffusion >>
rect 121 412 122 413 
<< pdiffusion >>
rect 122 412 123 413 
<< pdiffusion >>
rect 123 412 124 413 
<< pdiffusion >>
rect 124 412 125 413 
<< pdiffusion >>
rect 125 412 126 413 
<< m1 >>
rect 127 412 128 413 
<< pdiffusion >>
rect 138 412 139 413 
<< pdiffusion >>
rect 139 412 140 413 
<< pdiffusion >>
rect 140 412 141 413 
<< pdiffusion >>
rect 141 412 142 413 
<< pdiffusion >>
rect 142 412 143 413 
<< pdiffusion >>
rect 143 412 144 413 
<< pdiffusion >>
rect 156 412 157 413 
<< pdiffusion >>
rect 157 412 158 413 
<< pdiffusion >>
rect 158 412 159 413 
<< pdiffusion >>
rect 159 412 160 413 
<< pdiffusion >>
rect 160 412 161 413 
<< pdiffusion >>
rect 161 412 162 413 
<< pdiffusion >>
rect 174 412 175 413 
<< pdiffusion >>
rect 175 412 176 413 
<< pdiffusion >>
rect 176 412 177 413 
<< pdiffusion >>
rect 177 412 178 413 
<< pdiffusion >>
rect 178 412 179 413 
<< pdiffusion >>
rect 179 412 180 413 
<< pdiffusion >>
rect 192 412 193 413 
<< pdiffusion >>
rect 193 412 194 413 
<< pdiffusion >>
rect 194 412 195 413 
<< pdiffusion >>
rect 195 412 196 413 
<< pdiffusion >>
rect 196 412 197 413 
<< pdiffusion >>
rect 197 412 198 413 
<< pdiffusion >>
rect 210 412 211 413 
<< pdiffusion >>
rect 211 412 212 413 
<< pdiffusion >>
rect 212 412 213 413 
<< pdiffusion >>
rect 213 412 214 413 
<< pdiffusion >>
rect 214 412 215 413 
<< pdiffusion >>
rect 215 412 216 413 
<< pdiffusion >>
rect 228 412 229 413 
<< pdiffusion >>
rect 229 412 230 413 
<< pdiffusion >>
rect 230 412 231 413 
<< pdiffusion >>
rect 231 412 232 413 
<< pdiffusion >>
rect 232 412 233 413 
<< pdiffusion >>
rect 233 412 234 413 
<< pdiffusion >>
rect 246 412 247 413 
<< pdiffusion >>
rect 247 412 248 413 
<< pdiffusion >>
rect 248 412 249 413 
<< pdiffusion >>
rect 249 412 250 413 
<< pdiffusion >>
rect 250 412 251 413 
<< pdiffusion >>
rect 251 412 252 413 
<< pdiffusion >>
rect 264 412 265 413 
<< pdiffusion >>
rect 265 412 266 413 
<< pdiffusion >>
rect 266 412 267 413 
<< pdiffusion >>
rect 267 412 268 413 
<< pdiffusion >>
rect 268 412 269 413 
<< pdiffusion >>
rect 269 412 270 413 
<< pdiffusion >>
rect 282 412 283 413 
<< pdiffusion >>
rect 283 412 284 413 
<< pdiffusion >>
rect 284 412 285 413 
<< pdiffusion >>
rect 285 412 286 413 
<< pdiffusion >>
rect 286 412 287 413 
<< pdiffusion >>
rect 287 412 288 413 
<< m1 >>
rect 289 412 290 413 
<< pdiffusion >>
rect 300 412 301 413 
<< pdiffusion >>
rect 301 412 302 413 
<< pdiffusion >>
rect 302 412 303 413 
<< pdiffusion >>
rect 303 412 304 413 
<< pdiffusion >>
rect 304 412 305 413 
<< pdiffusion >>
rect 305 412 306 413 
<< pdiffusion >>
rect 336 412 337 413 
<< pdiffusion >>
rect 337 412 338 413 
<< pdiffusion >>
rect 338 412 339 413 
<< pdiffusion >>
rect 339 412 340 413 
<< pdiffusion >>
rect 340 412 341 413 
<< pdiffusion >>
rect 341 412 342 413 
<< pdiffusion >>
rect 354 412 355 413 
<< pdiffusion >>
rect 355 412 356 413 
<< pdiffusion >>
rect 356 412 357 413 
<< pdiffusion >>
rect 357 412 358 413 
<< pdiffusion >>
rect 358 412 359 413 
<< pdiffusion >>
rect 359 412 360 413 
<< pdiffusion >>
rect 372 412 373 413 
<< pdiffusion >>
rect 373 412 374 413 
<< pdiffusion >>
rect 374 412 375 413 
<< pdiffusion >>
rect 375 412 376 413 
<< pdiffusion >>
rect 376 412 377 413 
<< pdiffusion >>
rect 377 412 378 413 
<< pdiffusion >>
rect 390 412 391 413 
<< pdiffusion >>
rect 391 412 392 413 
<< pdiffusion >>
rect 392 412 393 413 
<< pdiffusion >>
rect 393 412 394 413 
<< pdiffusion >>
rect 394 412 395 413 
<< pdiffusion >>
rect 395 412 396 413 
<< pdiffusion >>
rect 408 412 409 413 
<< pdiffusion >>
rect 409 412 410 413 
<< pdiffusion >>
rect 410 412 411 413 
<< pdiffusion >>
rect 411 412 412 413 
<< pdiffusion >>
rect 412 412 413 413 
<< pdiffusion >>
rect 413 412 414 413 
<< pdiffusion >>
rect 426 412 427 413 
<< pdiffusion >>
rect 427 412 428 413 
<< pdiffusion >>
rect 428 412 429 413 
<< pdiffusion >>
rect 429 412 430 413 
<< pdiffusion >>
rect 430 412 431 413 
<< pdiffusion >>
rect 431 412 432 413 
<< pdiffusion >>
rect 444 412 445 413 
<< pdiffusion >>
rect 445 412 446 413 
<< pdiffusion >>
rect 446 412 447 413 
<< pdiffusion >>
rect 447 412 448 413 
<< pdiffusion >>
rect 448 412 449 413 
<< pdiffusion >>
rect 449 412 450 413 
<< pdiffusion >>
rect 12 413 13 414 
<< pdiffusion >>
rect 13 413 14 414 
<< pdiffusion >>
rect 14 413 15 414 
<< pdiffusion >>
rect 15 413 16 414 
<< pdiffusion >>
rect 16 413 17 414 
<< pdiffusion >>
rect 17 413 18 414 
<< pdiffusion >>
rect 30 413 31 414 
<< pdiffusion >>
rect 31 413 32 414 
<< pdiffusion >>
rect 32 413 33 414 
<< pdiffusion >>
rect 33 413 34 414 
<< pdiffusion >>
rect 34 413 35 414 
<< pdiffusion >>
rect 35 413 36 414 
<< pdiffusion >>
rect 48 413 49 414 
<< pdiffusion >>
rect 49 413 50 414 
<< pdiffusion >>
rect 50 413 51 414 
<< pdiffusion >>
rect 51 413 52 414 
<< m1 >>
rect 52 413 53 414 
<< pdiffusion >>
rect 52 413 53 414 
<< pdiffusion >>
rect 53 413 54 414 
<< m1 >>
rect 64 413 65 414 
<< pdiffusion >>
rect 66 413 67 414 
<< pdiffusion >>
rect 67 413 68 414 
<< pdiffusion >>
rect 68 413 69 414 
<< pdiffusion >>
rect 69 413 70 414 
<< m1 >>
rect 70 413 71 414 
<< pdiffusion >>
rect 70 413 71 414 
<< pdiffusion >>
rect 71 413 72 414 
<< pdiffusion >>
rect 84 413 85 414 
<< pdiffusion >>
rect 85 413 86 414 
<< pdiffusion >>
rect 86 413 87 414 
<< pdiffusion >>
rect 87 413 88 414 
<< pdiffusion >>
rect 88 413 89 414 
<< pdiffusion >>
rect 89 413 90 414 
<< pdiffusion >>
rect 102 413 103 414 
<< pdiffusion >>
rect 103 413 104 414 
<< pdiffusion >>
rect 104 413 105 414 
<< pdiffusion >>
rect 105 413 106 414 
<< pdiffusion >>
rect 106 413 107 414 
<< pdiffusion >>
rect 107 413 108 414 
<< pdiffusion >>
rect 120 413 121 414 
<< pdiffusion >>
rect 121 413 122 414 
<< pdiffusion >>
rect 122 413 123 414 
<< pdiffusion >>
rect 123 413 124 414 
<< m1 >>
rect 124 413 125 414 
<< pdiffusion >>
rect 124 413 125 414 
<< pdiffusion >>
rect 125 413 126 414 
<< m1 >>
rect 127 413 128 414 
<< pdiffusion >>
rect 138 413 139 414 
<< pdiffusion >>
rect 139 413 140 414 
<< pdiffusion >>
rect 140 413 141 414 
<< pdiffusion >>
rect 141 413 142 414 
<< pdiffusion >>
rect 142 413 143 414 
<< pdiffusion >>
rect 143 413 144 414 
<< pdiffusion >>
rect 156 413 157 414 
<< pdiffusion >>
rect 157 413 158 414 
<< pdiffusion >>
rect 158 413 159 414 
<< pdiffusion >>
rect 159 413 160 414 
<< pdiffusion >>
rect 160 413 161 414 
<< pdiffusion >>
rect 161 413 162 414 
<< pdiffusion >>
rect 174 413 175 414 
<< pdiffusion >>
rect 175 413 176 414 
<< pdiffusion >>
rect 176 413 177 414 
<< pdiffusion >>
rect 177 413 178 414 
<< pdiffusion >>
rect 178 413 179 414 
<< pdiffusion >>
rect 179 413 180 414 
<< pdiffusion >>
rect 192 413 193 414 
<< pdiffusion >>
rect 193 413 194 414 
<< pdiffusion >>
rect 194 413 195 414 
<< pdiffusion >>
rect 195 413 196 414 
<< pdiffusion >>
rect 196 413 197 414 
<< pdiffusion >>
rect 197 413 198 414 
<< pdiffusion >>
rect 210 413 211 414 
<< pdiffusion >>
rect 211 413 212 414 
<< pdiffusion >>
rect 212 413 213 414 
<< pdiffusion >>
rect 213 413 214 414 
<< pdiffusion >>
rect 214 413 215 414 
<< pdiffusion >>
rect 215 413 216 414 
<< pdiffusion >>
rect 228 413 229 414 
<< pdiffusion >>
rect 229 413 230 414 
<< pdiffusion >>
rect 230 413 231 414 
<< pdiffusion >>
rect 231 413 232 414 
<< pdiffusion >>
rect 232 413 233 414 
<< pdiffusion >>
rect 233 413 234 414 
<< pdiffusion >>
rect 246 413 247 414 
<< pdiffusion >>
rect 247 413 248 414 
<< pdiffusion >>
rect 248 413 249 414 
<< pdiffusion >>
rect 249 413 250 414 
<< pdiffusion >>
rect 250 413 251 414 
<< pdiffusion >>
rect 251 413 252 414 
<< pdiffusion >>
rect 264 413 265 414 
<< pdiffusion >>
rect 265 413 266 414 
<< pdiffusion >>
rect 266 413 267 414 
<< pdiffusion >>
rect 267 413 268 414 
<< pdiffusion >>
rect 268 413 269 414 
<< pdiffusion >>
rect 269 413 270 414 
<< pdiffusion >>
rect 282 413 283 414 
<< pdiffusion >>
rect 283 413 284 414 
<< pdiffusion >>
rect 284 413 285 414 
<< pdiffusion >>
rect 285 413 286 414 
<< pdiffusion >>
rect 286 413 287 414 
<< pdiffusion >>
rect 287 413 288 414 
<< m1 >>
rect 289 413 290 414 
<< pdiffusion >>
rect 300 413 301 414 
<< pdiffusion >>
rect 301 413 302 414 
<< pdiffusion >>
rect 302 413 303 414 
<< pdiffusion >>
rect 303 413 304 414 
<< pdiffusion >>
rect 304 413 305 414 
<< pdiffusion >>
rect 305 413 306 414 
<< pdiffusion >>
rect 336 413 337 414 
<< pdiffusion >>
rect 337 413 338 414 
<< pdiffusion >>
rect 338 413 339 414 
<< pdiffusion >>
rect 339 413 340 414 
<< pdiffusion >>
rect 340 413 341 414 
<< pdiffusion >>
rect 341 413 342 414 
<< pdiffusion >>
rect 354 413 355 414 
<< pdiffusion >>
rect 355 413 356 414 
<< pdiffusion >>
rect 356 413 357 414 
<< pdiffusion >>
rect 357 413 358 414 
<< pdiffusion >>
rect 358 413 359 414 
<< pdiffusion >>
rect 359 413 360 414 
<< pdiffusion >>
rect 372 413 373 414 
<< pdiffusion >>
rect 373 413 374 414 
<< pdiffusion >>
rect 374 413 375 414 
<< pdiffusion >>
rect 375 413 376 414 
<< pdiffusion >>
rect 376 413 377 414 
<< pdiffusion >>
rect 377 413 378 414 
<< pdiffusion >>
rect 390 413 391 414 
<< pdiffusion >>
rect 391 413 392 414 
<< pdiffusion >>
rect 392 413 393 414 
<< pdiffusion >>
rect 393 413 394 414 
<< pdiffusion >>
rect 394 413 395 414 
<< pdiffusion >>
rect 395 413 396 414 
<< pdiffusion >>
rect 408 413 409 414 
<< pdiffusion >>
rect 409 413 410 414 
<< pdiffusion >>
rect 410 413 411 414 
<< pdiffusion >>
rect 411 413 412 414 
<< pdiffusion >>
rect 412 413 413 414 
<< pdiffusion >>
rect 413 413 414 414 
<< pdiffusion >>
rect 426 413 427 414 
<< pdiffusion >>
rect 427 413 428 414 
<< pdiffusion >>
rect 428 413 429 414 
<< pdiffusion >>
rect 429 413 430 414 
<< pdiffusion >>
rect 430 413 431 414 
<< pdiffusion >>
rect 431 413 432 414 
<< pdiffusion >>
rect 444 413 445 414 
<< pdiffusion >>
rect 445 413 446 414 
<< pdiffusion >>
rect 446 413 447 414 
<< pdiffusion >>
rect 447 413 448 414 
<< pdiffusion >>
rect 448 413 449 414 
<< pdiffusion >>
rect 449 413 450 414 
<< m1 >>
rect 52 414 53 415 
<< m1 >>
rect 64 414 65 415 
<< m1 >>
rect 70 414 71 415 
<< m1 >>
rect 124 414 125 415 
<< m1 >>
rect 127 414 128 415 
<< m1 >>
rect 289 414 290 415 
<< m1 >>
rect 52 415 53 416 
<< m1 >>
rect 64 415 65 416 
<< m1 >>
rect 70 415 71 416 
<< m1 >>
rect 124 415 125 416 
<< m1 >>
rect 125 415 126 416 
<< m1 >>
rect 126 415 127 416 
<< m1 >>
rect 127 415 128 416 
<< m1 >>
rect 289 415 290 416 
<< m1 >>
rect 52 416 53 417 
<< m1 >>
rect 64 416 65 417 
<< m1 >>
rect 70 416 71 417 
<< m1 >>
rect 289 416 290 417 
<< m1 >>
rect 52 417 53 418 
<< m1 >>
rect 64 417 65 418 
<< m1 >>
rect 70 417 71 418 
<< m1 >>
rect 289 417 290 418 
<< m1 >>
rect 46 418 47 419 
<< m1 >>
rect 47 418 48 419 
<< m1 >>
rect 48 418 49 419 
<< m1 >>
rect 49 418 50 419 
<< m1 >>
rect 50 418 51 419 
<< m1 >>
rect 51 418 52 419 
<< m1 >>
rect 52 418 53 419 
<< m1 >>
rect 64 418 65 419 
<< m1 >>
rect 65 418 66 419 
<< m1 >>
rect 66 418 67 419 
<< m1 >>
rect 67 418 68 419 
<< m1 >>
rect 68 418 69 419 
<< m1 >>
rect 69 418 70 419 
<< m1 >>
rect 70 418 71 419 
<< m1 >>
rect 289 418 290 419 
<< m1 >>
rect 46 419 47 420 
<< m1 >>
rect 289 419 290 420 
<< m1 >>
rect 46 420 47 421 
<< m1 >>
rect 289 420 290 421 
<< m1 >>
rect 46 421 47 422 
<< m1 >>
rect 289 421 290 422 
<< m1 >>
rect 46 422 47 423 
<< m1 >>
rect 289 422 290 423 
<< m1 >>
rect 46 423 47 424 
<< m1 >>
rect 139 423 140 424 
<< m1 >>
rect 140 423 141 424 
<< m1 >>
rect 141 423 142 424 
<< m1 >>
rect 142 423 143 424 
<< m1 >>
rect 143 423 144 424 
<< m1 >>
rect 144 423 145 424 
<< m1 >>
rect 145 423 146 424 
<< m1 >>
rect 146 423 147 424 
<< m1 >>
rect 147 423 148 424 
<< m1 >>
rect 148 423 149 424 
<< m1 >>
rect 149 423 150 424 
<< m1 >>
rect 150 423 151 424 
<< m1 >>
rect 151 423 152 424 
<< m1 >>
rect 152 423 153 424 
<< m1 >>
rect 153 423 154 424 
<< m1 >>
rect 154 423 155 424 
<< m1 >>
rect 289 423 290 424 
<< m1 >>
rect 301 423 302 424 
<< m1 >>
rect 302 423 303 424 
<< m1 >>
rect 303 423 304 424 
<< m1 >>
rect 304 423 305 424 
<< m1 >>
rect 305 423 306 424 
<< m1 >>
rect 306 423 307 424 
<< m1 >>
rect 307 423 308 424 
<< m1 >>
rect 46 424 47 425 
<< m1 >>
rect 52 424 53 425 
<< m1 >>
rect 53 424 54 425 
<< m1 >>
rect 54 424 55 425 
<< m1 >>
rect 55 424 56 425 
<< m1 >>
rect 56 424 57 425 
<< m1 >>
rect 57 424 58 425 
<< m1 >>
rect 58 424 59 425 
<< m1 >>
rect 59 424 60 425 
<< m1 >>
rect 60 424 61 425 
<< m1 >>
rect 61 424 62 425 
<< m1 >>
rect 62 424 63 425 
<< m1 >>
rect 63 424 64 425 
<< m1 >>
rect 64 424 65 425 
<< m1 >>
rect 139 424 140 425 
<< m2 >>
rect 145 424 146 425 
<< m2 >>
rect 146 424 147 425 
<< m2 >>
rect 147 424 148 425 
<< m2 >>
rect 148 424 149 425 
<< m2 >>
rect 149 424 150 425 
<< m2 >>
rect 150 424 151 425 
<< m2 >>
rect 151 424 152 425 
<< m2 >>
rect 152 424 153 425 
<< m2 >>
rect 153 424 154 425 
<< m1 >>
rect 154 424 155 425 
<< m2 >>
rect 154 424 155 425 
<< m2 >>
rect 155 424 156 425 
<< m1 >>
rect 156 424 157 425 
<< m2 >>
rect 156 424 157 425 
<< m2c >>
rect 156 424 157 425 
<< m1 >>
rect 156 424 157 425 
<< m2 >>
rect 156 424 157 425 
<< m1 >>
rect 157 424 158 425 
<< m1 >>
rect 226 424 227 425 
<< m1 >>
rect 227 424 228 425 
<< m1 >>
rect 228 424 229 425 
<< m1 >>
rect 229 424 230 425 
<< m1 >>
rect 289 424 290 425 
<< m1 >>
rect 301 424 302 425 
<< m1 >>
rect 307 424 308 425 
<< m1 >>
rect 46 425 47 426 
<< m1 >>
rect 52 425 53 426 
<< m1 >>
rect 64 425 65 426 
<< m1 >>
rect 139 425 140 426 
<< m1 >>
rect 145 425 146 426 
<< m2 >>
rect 145 425 146 426 
<< m2c >>
rect 145 425 146 426 
<< m1 >>
rect 145 425 146 426 
<< m2 >>
rect 145 425 146 426 
<< m1 >>
rect 154 425 155 426 
<< m1 >>
rect 157 425 158 426 
<< m1 >>
rect 226 425 227 426 
<< m1 >>
rect 229 425 230 426 
<< m1 >>
rect 289 425 290 426 
<< m1 >>
rect 301 425 302 426 
<< m1 >>
rect 307 425 308 426 
<< pdiffusion >>
rect 12 426 13 427 
<< pdiffusion >>
rect 13 426 14 427 
<< pdiffusion >>
rect 14 426 15 427 
<< pdiffusion >>
rect 15 426 16 427 
<< pdiffusion >>
rect 16 426 17 427 
<< pdiffusion >>
rect 17 426 18 427 
<< pdiffusion >>
rect 30 426 31 427 
<< pdiffusion >>
rect 31 426 32 427 
<< pdiffusion >>
rect 32 426 33 427 
<< pdiffusion >>
rect 33 426 34 427 
<< pdiffusion >>
rect 34 426 35 427 
<< pdiffusion >>
rect 35 426 36 427 
<< m1 >>
rect 46 426 47 427 
<< pdiffusion >>
rect 48 426 49 427 
<< pdiffusion >>
rect 49 426 50 427 
<< pdiffusion >>
rect 50 426 51 427 
<< pdiffusion >>
rect 51 426 52 427 
<< m1 >>
rect 52 426 53 427 
<< pdiffusion >>
rect 52 426 53 427 
<< pdiffusion >>
rect 53 426 54 427 
<< m1 >>
rect 64 426 65 427 
<< pdiffusion >>
rect 66 426 67 427 
<< pdiffusion >>
rect 67 426 68 427 
<< pdiffusion >>
rect 68 426 69 427 
<< pdiffusion >>
rect 69 426 70 427 
<< pdiffusion >>
rect 70 426 71 427 
<< pdiffusion >>
rect 71 426 72 427 
<< pdiffusion >>
rect 84 426 85 427 
<< pdiffusion >>
rect 85 426 86 427 
<< pdiffusion >>
rect 86 426 87 427 
<< pdiffusion >>
rect 87 426 88 427 
<< pdiffusion >>
rect 88 426 89 427 
<< pdiffusion >>
rect 89 426 90 427 
<< pdiffusion >>
rect 120 426 121 427 
<< pdiffusion >>
rect 121 426 122 427 
<< pdiffusion >>
rect 122 426 123 427 
<< pdiffusion >>
rect 123 426 124 427 
<< pdiffusion >>
rect 124 426 125 427 
<< pdiffusion >>
rect 125 426 126 427 
<< pdiffusion >>
rect 138 426 139 427 
<< m1 >>
rect 139 426 140 427 
<< pdiffusion >>
rect 139 426 140 427 
<< pdiffusion >>
rect 140 426 141 427 
<< pdiffusion >>
rect 141 426 142 427 
<< pdiffusion >>
rect 142 426 143 427 
<< pdiffusion >>
rect 143 426 144 427 
<< m1 >>
rect 145 426 146 427 
<< m1 >>
rect 154 426 155 427 
<< pdiffusion >>
rect 156 426 157 427 
<< m1 >>
rect 157 426 158 427 
<< pdiffusion >>
rect 157 426 158 427 
<< pdiffusion >>
rect 158 426 159 427 
<< pdiffusion >>
rect 159 426 160 427 
<< pdiffusion >>
rect 160 426 161 427 
<< pdiffusion >>
rect 161 426 162 427 
<< pdiffusion >>
rect 174 426 175 427 
<< pdiffusion >>
rect 175 426 176 427 
<< pdiffusion >>
rect 176 426 177 427 
<< pdiffusion >>
rect 177 426 178 427 
<< pdiffusion >>
rect 178 426 179 427 
<< pdiffusion >>
rect 179 426 180 427 
<< pdiffusion >>
rect 192 426 193 427 
<< pdiffusion >>
rect 193 426 194 427 
<< pdiffusion >>
rect 194 426 195 427 
<< pdiffusion >>
rect 195 426 196 427 
<< pdiffusion >>
rect 196 426 197 427 
<< pdiffusion >>
rect 197 426 198 427 
<< pdiffusion >>
rect 210 426 211 427 
<< pdiffusion >>
rect 211 426 212 427 
<< pdiffusion >>
rect 212 426 213 427 
<< pdiffusion >>
rect 213 426 214 427 
<< pdiffusion >>
rect 214 426 215 427 
<< pdiffusion >>
rect 215 426 216 427 
<< m1 >>
rect 226 426 227 427 
<< pdiffusion >>
rect 228 426 229 427 
<< m1 >>
rect 229 426 230 427 
<< pdiffusion >>
rect 229 426 230 427 
<< pdiffusion >>
rect 230 426 231 427 
<< pdiffusion >>
rect 231 426 232 427 
<< pdiffusion >>
rect 232 426 233 427 
<< pdiffusion >>
rect 233 426 234 427 
<< pdiffusion >>
rect 246 426 247 427 
<< pdiffusion >>
rect 247 426 248 427 
<< pdiffusion >>
rect 248 426 249 427 
<< pdiffusion >>
rect 249 426 250 427 
<< pdiffusion >>
rect 250 426 251 427 
<< pdiffusion >>
rect 251 426 252 427 
<< pdiffusion >>
rect 264 426 265 427 
<< pdiffusion >>
rect 265 426 266 427 
<< pdiffusion >>
rect 266 426 267 427 
<< pdiffusion >>
rect 267 426 268 427 
<< pdiffusion >>
rect 268 426 269 427 
<< pdiffusion >>
rect 269 426 270 427 
<< pdiffusion >>
rect 282 426 283 427 
<< pdiffusion >>
rect 283 426 284 427 
<< pdiffusion >>
rect 284 426 285 427 
<< pdiffusion >>
rect 285 426 286 427 
<< pdiffusion >>
rect 286 426 287 427 
<< pdiffusion >>
rect 287 426 288 427 
<< m1 >>
rect 289 426 290 427 
<< pdiffusion >>
rect 300 426 301 427 
<< m1 >>
rect 301 426 302 427 
<< pdiffusion >>
rect 301 426 302 427 
<< pdiffusion >>
rect 302 426 303 427 
<< pdiffusion >>
rect 303 426 304 427 
<< pdiffusion >>
rect 304 426 305 427 
<< pdiffusion >>
rect 305 426 306 427 
<< m1 >>
rect 307 426 308 427 
<< pdiffusion >>
rect 318 426 319 427 
<< pdiffusion >>
rect 319 426 320 427 
<< pdiffusion >>
rect 320 426 321 427 
<< pdiffusion >>
rect 321 426 322 427 
<< pdiffusion >>
rect 322 426 323 427 
<< pdiffusion >>
rect 323 426 324 427 
<< pdiffusion >>
rect 336 426 337 427 
<< pdiffusion >>
rect 337 426 338 427 
<< pdiffusion >>
rect 338 426 339 427 
<< pdiffusion >>
rect 339 426 340 427 
<< pdiffusion >>
rect 340 426 341 427 
<< pdiffusion >>
rect 341 426 342 427 
<< pdiffusion >>
rect 354 426 355 427 
<< pdiffusion >>
rect 355 426 356 427 
<< pdiffusion >>
rect 356 426 357 427 
<< pdiffusion >>
rect 357 426 358 427 
<< pdiffusion >>
rect 358 426 359 427 
<< pdiffusion >>
rect 359 426 360 427 
<< pdiffusion >>
rect 372 426 373 427 
<< pdiffusion >>
rect 373 426 374 427 
<< pdiffusion >>
rect 374 426 375 427 
<< pdiffusion >>
rect 375 426 376 427 
<< pdiffusion >>
rect 376 426 377 427 
<< pdiffusion >>
rect 377 426 378 427 
<< pdiffusion >>
rect 390 426 391 427 
<< pdiffusion >>
rect 391 426 392 427 
<< pdiffusion >>
rect 392 426 393 427 
<< pdiffusion >>
rect 393 426 394 427 
<< pdiffusion >>
rect 394 426 395 427 
<< pdiffusion >>
rect 395 426 396 427 
<< pdiffusion >>
rect 408 426 409 427 
<< pdiffusion >>
rect 409 426 410 427 
<< pdiffusion >>
rect 410 426 411 427 
<< pdiffusion >>
rect 411 426 412 427 
<< pdiffusion >>
rect 412 426 413 427 
<< pdiffusion >>
rect 413 426 414 427 
<< pdiffusion >>
rect 426 426 427 427 
<< pdiffusion >>
rect 427 426 428 427 
<< pdiffusion >>
rect 428 426 429 427 
<< pdiffusion >>
rect 429 426 430 427 
<< pdiffusion >>
rect 430 426 431 427 
<< pdiffusion >>
rect 431 426 432 427 
<< pdiffusion >>
rect 444 426 445 427 
<< pdiffusion >>
rect 445 426 446 427 
<< pdiffusion >>
rect 446 426 447 427 
<< pdiffusion >>
rect 447 426 448 427 
<< pdiffusion >>
rect 448 426 449 427 
<< pdiffusion >>
rect 449 426 450 427 
<< pdiffusion >>
rect 12 427 13 428 
<< pdiffusion >>
rect 13 427 14 428 
<< pdiffusion >>
rect 14 427 15 428 
<< pdiffusion >>
rect 15 427 16 428 
<< pdiffusion >>
rect 16 427 17 428 
<< pdiffusion >>
rect 17 427 18 428 
<< pdiffusion >>
rect 30 427 31 428 
<< pdiffusion >>
rect 31 427 32 428 
<< pdiffusion >>
rect 32 427 33 428 
<< pdiffusion >>
rect 33 427 34 428 
<< pdiffusion >>
rect 34 427 35 428 
<< pdiffusion >>
rect 35 427 36 428 
<< m1 >>
rect 46 427 47 428 
<< pdiffusion >>
rect 48 427 49 428 
<< pdiffusion >>
rect 49 427 50 428 
<< pdiffusion >>
rect 50 427 51 428 
<< pdiffusion >>
rect 51 427 52 428 
<< pdiffusion >>
rect 52 427 53 428 
<< pdiffusion >>
rect 53 427 54 428 
<< m1 >>
rect 64 427 65 428 
<< pdiffusion >>
rect 66 427 67 428 
<< pdiffusion >>
rect 67 427 68 428 
<< pdiffusion >>
rect 68 427 69 428 
<< pdiffusion >>
rect 69 427 70 428 
<< pdiffusion >>
rect 70 427 71 428 
<< pdiffusion >>
rect 71 427 72 428 
<< pdiffusion >>
rect 84 427 85 428 
<< pdiffusion >>
rect 85 427 86 428 
<< pdiffusion >>
rect 86 427 87 428 
<< pdiffusion >>
rect 87 427 88 428 
<< pdiffusion >>
rect 88 427 89 428 
<< pdiffusion >>
rect 89 427 90 428 
<< pdiffusion >>
rect 120 427 121 428 
<< pdiffusion >>
rect 121 427 122 428 
<< pdiffusion >>
rect 122 427 123 428 
<< pdiffusion >>
rect 123 427 124 428 
<< pdiffusion >>
rect 124 427 125 428 
<< pdiffusion >>
rect 125 427 126 428 
<< pdiffusion >>
rect 138 427 139 428 
<< pdiffusion >>
rect 139 427 140 428 
<< pdiffusion >>
rect 140 427 141 428 
<< pdiffusion >>
rect 141 427 142 428 
<< pdiffusion >>
rect 142 427 143 428 
<< pdiffusion >>
rect 143 427 144 428 
<< m1 >>
rect 145 427 146 428 
<< m1 >>
rect 154 427 155 428 
<< pdiffusion >>
rect 156 427 157 428 
<< pdiffusion >>
rect 157 427 158 428 
<< pdiffusion >>
rect 158 427 159 428 
<< pdiffusion >>
rect 159 427 160 428 
<< pdiffusion >>
rect 160 427 161 428 
<< pdiffusion >>
rect 161 427 162 428 
<< pdiffusion >>
rect 174 427 175 428 
<< pdiffusion >>
rect 175 427 176 428 
<< pdiffusion >>
rect 176 427 177 428 
<< pdiffusion >>
rect 177 427 178 428 
<< pdiffusion >>
rect 178 427 179 428 
<< pdiffusion >>
rect 179 427 180 428 
<< pdiffusion >>
rect 192 427 193 428 
<< pdiffusion >>
rect 193 427 194 428 
<< pdiffusion >>
rect 194 427 195 428 
<< pdiffusion >>
rect 195 427 196 428 
<< pdiffusion >>
rect 196 427 197 428 
<< pdiffusion >>
rect 197 427 198 428 
<< pdiffusion >>
rect 210 427 211 428 
<< pdiffusion >>
rect 211 427 212 428 
<< pdiffusion >>
rect 212 427 213 428 
<< pdiffusion >>
rect 213 427 214 428 
<< pdiffusion >>
rect 214 427 215 428 
<< pdiffusion >>
rect 215 427 216 428 
<< m1 >>
rect 226 427 227 428 
<< pdiffusion >>
rect 228 427 229 428 
<< pdiffusion >>
rect 229 427 230 428 
<< pdiffusion >>
rect 230 427 231 428 
<< pdiffusion >>
rect 231 427 232 428 
<< pdiffusion >>
rect 232 427 233 428 
<< pdiffusion >>
rect 233 427 234 428 
<< pdiffusion >>
rect 246 427 247 428 
<< pdiffusion >>
rect 247 427 248 428 
<< pdiffusion >>
rect 248 427 249 428 
<< pdiffusion >>
rect 249 427 250 428 
<< pdiffusion >>
rect 250 427 251 428 
<< pdiffusion >>
rect 251 427 252 428 
<< pdiffusion >>
rect 264 427 265 428 
<< pdiffusion >>
rect 265 427 266 428 
<< pdiffusion >>
rect 266 427 267 428 
<< pdiffusion >>
rect 267 427 268 428 
<< pdiffusion >>
rect 268 427 269 428 
<< pdiffusion >>
rect 269 427 270 428 
<< pdiffusion >>
rect 282 427 283 428 
<< pdiffusion >>
rect 283 427 284 428 
<< pdiffusion >>
rect 284 427 285 428 
<< pdiffusion >>
rect 285 427 286 428 
<< pdiffusion >>
rect 286 427 287 428 
<< pdiffusion >>
rect 287 427 288 428 
<< m1 >>
rect 289 427 290 428 
<< pdiffusion >>
rect 300 427 301 428 
<< pdiffusion >>
rect 301 427 302 428 
<< pdiffusion >>
rect 302 427 303 428 
<< pdiffusion >>
rect 303 427 304 428 
<< pdiffusion >>
rect 304 427 305 428 
<< pdiffusion >>
rect 305 427 306 428 
<< m1 >>
rect 307 427 308 428 
<< pdiffusion >>
rect 318 427 319 428 
<< pdiffusion >>
rect 319 427 320 428 
<< pdiffusion >>
rect 320 427 321 428 
<< pdiffusion >>
rect 321 427 322 428 
<< pdiffusion >>
rect 322 427 323 428 
<< pdiffusion >>
rect 323 427 324 428 
<< pdiffusion >>
rect 336 427 337 428 
<< pdiffusion >>
rect 337 427 338 428 
<< pdiffusion >>
rect 338 427 339 428 
<< pdiffusion >>
rect 339 427 340 428 
<< pdiffusion >>
rect 340 427 341 428 
<< pdiffusion >>
rect 341 427 342 428 
<< pdiffusion >>
rect 354 427 355 428 
<< pdiffusion >>
rect 355 427 356 428 
<< pdiffusion >>
rect 356 427 357 428 
<< pdiffusion >>
rect 357 427 358 428 
<< pdiffusion >>
rect 358 427 359 428 
<< pdiffusion >>
rect 359 427 360 428 
<< pdiffusion >>
rect 372 427 373 428 
<< pdiffusion >>
rect 373 427 374 428 
<< pdiffusion >>
rect 374 427 375 428 
<< pdiffusion >>
rect 375 427 376 428 
<< pdiffusion >>
rect 376 427 377 428 
<< pdiffusion >>
rect 377 427 378 428 
<< pdiffusion >>
rect 390 427 391 428 
<< pdiffusion >>
rect 391 427 392 428 
<< pdiffusion >>
rect 392 427 393 428 
<< pdiffusion >>
rect 393 427 394 428 
<< pdiffusion >>
rect 394 427 395 428 
<< pdiffusion >>
rect 395 427 396 428 
<< pdiffusion >>
rect 408 427 409 428 
<< pdiffusion >>
rect 409 427 410 428 
<< pdiffusion >>
rect 410 427 411 428 
<< pdiffusion >>
rect 411 427 412 428 
<< pdiffusion >>
rect 412 427 413 428 
<< pdiffusion >>
rect 413 427 414 428 
<< pdiffusion >>
rect 426 427 427 428 
<< pdiffusion >>
rect 427 427 428 428 
<< pdiffusion >>
rect 428 427 429 428 
<< pdiffusion >>
rect 429 427 430 428 
<< pdiffusion >>
rect 430 427 431 428 
<< pdiffusion >>
rect 431 427 432 428 
<< pdiffusion >>
rect 444 427 445 428 
<< pdiffusion >>
rect 445 427 446 428 
<< pdiffusion >>
rect 446 427 447 428 
<< pdiffusion >>
rect 447 427 448 428 
<< pdiffusion >>
rect 448 427 449 428 
<< pdiffusion >>
rect 449 427 450 428 
<< pdiffusion >>
rect 12 428 13 429 
<< pdiffusion >>
rect 13 428 14 429 
<< pdiffusion >>
rect 14 428 15 429 
<< pdiffusion >>
rect 15 428 16 429 
<< pdiffusion >>
rect 16 428 17 429 
<< pdiffusion >>
rect 17 428 18 429 
<< pdiffusion >>
rect 30 428 31 429 
<< pdiffusion >>
rect 31 428 32 429 
<< pdiffusion >>
rect 32 428 33 429 
<< pdiffusion >>
rect 33 428 34 429 
<< pdiffusion >>
rect 34 428 35 429 
<< pdiffusion >>
rect 35 428 36 429 
<< m1 >>
rect 46 428 47 429 
<< pdiffusion >>
rect 48 428 49 429 
<< pdiffusion >>
rect 49 428 50 429 
<< pdiffusion >>
rect 50 428 51 429 
<< pdiffusion >>
rect 51 428 52 429 
<< pdiffusion >>
rect 52 428 53 429 
<< pdiffusion >>
rect 53 428 54 429 
<< m1 >>
rect 64 428 65 429 
<< pdiffusion >>
rect 66 428 67 429 
<< pdiffusion >>
rect 67 428 68 429 
<< pdiffusion >>
rect 68 428 69 429 
<< pdiffusion >>
rect 69 428 70 429 
<< pdiffusion >>
rect 70 428 71 429 
<< pdiffusion >>
rect 71 428 72 429 
<< pdiffusion >>
rect 84 428 85 429 
<< pdiffusion >>
rect 85 428 86 429 
<< pdiffusion >>
rect 86 428 87 429 
<< pdiffusion >>
rect 87 428 88 429 
<< pdiffusion >>
rect 88 428 89 429 
<< pdiffusion >>
rect 89 428 90 429 
<< pdiffusion >>
rect 120 428 121 429 
<< pdiffusion >>
rect 121 428 122 429 
<< pdiffusion >>
rect 122 428 123 429 
<< pdiffusion >>
rect 123 428 124 429 
<< pdiffusion >>
rect 124 428 125 429 
<< pdiffusion >>
rect 125 428 126 429 
<< pdiffusion >>
rect 138 428 139 429 
<< pdiffusion >>
rect 139 428 140 429 
<< pdiffusion >>
rect 140 428 141 429 
<< pdiffusion >>
rect 141 428 142 429 
<< pdiffusion >>
rect 142 428 143 429 
<< pdiffusion >>
rect 143 428 144 429 
<< m1 >>
rect 145 428 146 429 
<< m1 >>
rect 154 428 155 429 
<< pdiffusion >>
rect 156 428 157 429 
<< pdiffusion >>
rect 157 428 158 429 
<< pdiffusion >>
rect 158 428 159 429 
<< pdiffusion >>
rect 159 428 160 429 
<< pdiffusion >>
rect 160 428 161 429 
<< pdiffusion >>
rect 161 428 162 429 
<< pdiffusion >>
rect 174 428 175 429 
<< pdiffusion >>
rect 175 428 176 429 
<< pdiffusion >>
rect 176 428 177 429 
<< pdiffusion >>
rect 177 428 178 429 
<< pdiffusion >>
rect 178 428 179 429 
<< pdiffusion >>
rect 179 428 180 429 
<< pdiffusion >>
rect 192 428 193 429 
<< pdiffusion >>
rect 193 428 194 429 
<< pdiffusion >>
rect 194 428 195 429 
<< pdiffusion >>
rect 195 428 196 429 
<< pdiffusion >>
rect 196 428 197 429 
<< pdiffusion >>
rect 197 428 198 429 
<< pdiffusion >>
rect 210 428 211 429 
<< pdiffusion >>
rect 211 428 212 429 
<< pdiffusion >>
rect 212 428 213 429 
<< pdiffusion >>
rect 213 428 214 429 
<< pdiffusion >>
rect 214 428 215 429 
<< pdiffusion >>
rect 215 428 216 429 
<< m1 >>
rect 226 428 227 429 
<< pdiffusion >>
rect 228 428 229 429 
<< pdiffusion >>
rect 229 428 230 429 
<< pdiffusion >>
rect 230 428 231 429 
<< pdiffusion >>
rect 231 428 232 429 
<< pdiffusion >>
rect 232 428 233 429 
<< pdiffusion >>
rect 233 428 234 429 
<< pdiffusion >>
rect 246 428 247 429 
<< pdiffusion >>
rect 247 428 248 429 
<< pdiffusion >>
rect 248 428 249 429 
<< pdiffusion >>
rect 249 428 250 429 
<< pdiffusion >>
rect 250 428 251 429 
<< pdiffusion >>
rect 251 428 252 429 
<< pdiffusion >>
rect 264 428 265 429 
<< pdiffusion >>
rect 265 428 266 429 
<< pdiffusion >>
rect 266 428 267 429 
<< pdiffusion >>
rect 267 428 268 429 
<< pdiffusion >>
rect 268 428 269 429 
<< pdiffusion >>
rect 269 428 270 429 
<< pdiffusion >>
rect 282 428 283 429 
<< pdiffusion >>
rect 283 428 284 429 
<< pdiffusion >>
rect 284 428 285 429 
<< pdiffusion >>
rect 285 428 286 429 
<< pdiffusion >>
rect 286 428 287 429 
<< pdiffusion >>
rect 287 428 288 429 
<< m1 >>
rect 289 428 290 429 
<< pdiffusion >>
rect 300 428 301 429 
<< pdiffusion >>
rect 301 428 302 429 
<< pdiffusion >>
rect 302 428 303 429 
<< pdiffusion >>
rect 303 428 304 429 
<< pdiffusion >>
rect 304 428 305 429 
<< pdiffusion >>
rect 305 428 306 429 
<< m1 >>
rect 307 428 308 429 
<< pdiffusion >>
rect 318 428 319 429 
<< pdiffusion >>
rect 319 428 320 429 
<< pdiffusion >>
rect 320 428 321 429 
<< pdiffusion >>
rect 321 428 322 429 
<< pdiffusion >>
rect 322 428 323 429 
<< pdiffusion >>
rect 323 428 324 429 
<< pdiffusion >>
rect 336 428 337 429 
<< pdiffusion >>
rect 337 428 338 429 
<< pdiffusion >>
rect 338 428 339 429 
<< pdiffusion >>
rect 339 428 340 429 
<< pdiffusion >>
rect 340 428 341 429 
<< pdiffusion >>
rect 341 428 342 429 
<< pdiffusion >>
rect 354 428 355 429 
<< pdiffusion >>
rect 355 428 356 429 
<< pdiffusion >>
rect 356 428 357 429 
<< pdiffusion >>
rect 357 428 358 429 
<< pdiffusion >>
rect 358 428 359 429 
<< pdiffusion >>
rect 359 428 360 429 
<< pdiffusion >>
rect 372 428 373 429 
<< pdiffusion >>
rect 373 428 374 429 
<< pdiffusion >>
rect 374 428 375 429 
<< pdiffusion >>
rect 375 428 376 429 
<< pdiffusion >>
rect 376 428 377 429 
<< pdiffusion >>
rect 377 428 378 429 
<< pdiffusion >>
rect 390 428 391 429 
<< pdiffusion >>
rect 391 428 392 429 
<< pdiffusion >>
rect 392 428 393 429 
<< pdiffusion >>
rect 393 428 394 429 
<< pdiffusion >>
rect 394 428 395 429 
<< pdiffusion >>
rect 395 428 396 429 
<< pdiffusion >>
rect 408 428 409 429 
<< pdiffusion >>
rect 409 428 410 429 
<< pdiffusion >>
rect 410 428 411 429 
<< pdiffusion >>
rect 411 428 412 429 
<< pdiffusion >>
rect 412 428 413 429 
<< pdiffusion >>
rect 413 428 414 429 
<< pdiffusion >>
rect 426 428 427 429 
<< pdiffusion >>
rect 427 428 428 429 
<< pdiffusion >>
rect 428 428 429 429 
<< pdiffusion >>
rect 429 428 430 429 
<< pdiffusion >>
rect 430 428 431 429 
<< pdiffusion >>
rect 431 428 432 429 
<< pdiffusion >>
rect 444 428 445 429 
<< pdiffusion >>
rect 445 428 446 429 
<< pdiffusion >>
rect 446 428 447 429 
<< pdiffusion >>
rect 447 428 448 429 
<< pdiffusion >>
rect 448 428 449 429 
<< pdiffusion >>
rect 449 428 450 429 
<< pdiffusion >>
rect 12 429 13 430 
<< pdiffusion >>
rect 13 429 14 430 
<< pdiffusion >>
rect 14 429 15 430 
<< pdiffusion >>
rect 15 429 16 430 
<< pdiffusion >>
rect 16 429 17 430 
<< pdiffusion >>
rect 17 429 18 430 
<< pdiffusion >>
rect 30 429 31 430 
<< pdiffusion >>
rect 31 429 32 430 
<< pdiffusion >>
rect 32 429 33 430 
<< pdiffusion >>
rect 33 429 34 430 
<< pdiffusion >>
rect 34 429 35 430 
<< pdiffusion >>
rect 35 429 36 430 
<< m1 >>
rect 46 429 47 430 
<< pdiffusion >>
rect 48 429 49 430 
<< pdiffusion >>
rect 49 429 50 430 
<< pdiffusion >>
rect 50 429 51 430 
<< pdiffusion >>
rect 51 429 52 430 
<< pdiffusion >>
rect 52 429 53 430 
<< pdiffusion >>
rect 53 429 54 430 
<< m1 >>
rect 64 429 65 430 
<< pdiffusion >>
rect 66 429 67 430 
<< pdiffusion >>
rect 67 429 68 430 
<< pdiffusion >>
rect 68 429 69 430 
<< pdiffusion >>
rect 69 429 70 430 
<< pdiffusion >>
rect 70 429 71 430 
<< pdiffusion >>
rect 71 429 72 430 
<< pdiffusion >>
rect 84 429 85 430 
<< pdiffusion >>
rect 85 429 86 430 
<< pdiffusion >>
rect 86 429 87 430 
<< pdiffusion >>
rect 87 429 88 430 
<< pdiffusion >>
rect 88 429 89 430 
<< pdiffusion >>
rect 89 429 90 430 
<< pdiffusion >>
rect 120 429 121 430 
<< pdiffusion >>
rect 121 429 122 430 
<< pdiffusion >>
rect 122 429 123 430 
<< pdiffusion >>
rect 123 429 124 430 
<< pdiffusion >>
rect 124 429 125 430 
<< pdiffusion >>
rect 125 429 126 430 
<< pdiffusion >>
rect 138 429 139 430 
<< pdiffusion >>
rect 139 429 140 430 
<< pdiffusion >>
rect 140 429 141 430 
<< pdiffusion >>
rect 141 429 142 430 
<< pdiffusion >>
rect 142 429 143 430 
<< pdiffusion >>
rect 143 429 144 430 
<< m1 >>
rect 145 429 146 430 
<< m1 >>
rect 154 429 155 430 
<< pdiffusion >>
rect 156 429 157 430 
<< pdiffusion >>
rect 157 429 158 430 
<< pdiffusion >>
rect 158 429 159 430 
<< pdiffusion >>
rect 159 429 160 430 
<< pdiffusion >>
rect 160 429 161 430 
<< pdiffusion >>
rect 161 429 162 430 
<< pdiffusion >>
rect 174 429 175 430 
<< pdiffusion >>
rect 175 429 176 430 
<< pdiffusion >>
rect 176 429 177 430 
<< pdiffusion >>
rect 177 429 178 430 
<< pdiffusion >>
rect 178 429 179 430 
<< pdiffusion >>
rect 179 429 180 430 
<< pdiffusion >>
rect 192 429 193 430 
<< pdiffusion >>
rect 193 429 194 430 
<< pdiffusion >>
rect 194 429 195 430 
<< pdiffusion >>
rect 195 429 196 430 
<< pdiffusion >>
rect 196 429 197 430 
<< pdiffusion >>
rect 197 429 198 430 
<< pdiffusion >>
rect 210 429 211 430 
<< pdiffusion >>
rect 211 429 212 430 
<< pdiffusion >>
rect 212 429 213 430 
<< pdiffusion >>
rect 213 429 214 430 
<< pdiffusion >>
rect 214 429 215 430 
<< pdiffusion >>
rect 215 429 216 430 
<< m1 >>
rect 226 429 227 430 
<< pdiffusion >>
rect 228 429 229 430 
<< pdiffusion >>
rect 229 429 230 430 
<< pdiffusion >>
rect 230 429 231 430 
<< pdiffusion >>
rect 231 429 232 430 
<< pdiffusion >>
rect 232 429 233 430 
<< pdiffusion >>
rect 233 429 234 430 
<< pdiffusion >>
rect 246 429 247 430 
<< pdiffusion >>
rect 247 429 248 430 
<< pdiffusion >>
rect 248 429 249 430 
<< pdiffusion >>
rect 249 429 250 430 
<< pdiffusion >>
rect 250 429 251 430 
<< pdiffusion >>
rect 251 429 252 430 
<< pdiffusion >>
rect 264 429 265 430 
<< pdiffusion >>
rect 265 429 266 430 
<< pdiffusion >>
rect 266 429 267 430 
<< pdiffusion >>
rect 267 429 268 430 
<< pdiffusion >>
rect 268 429 269 430 
<< pdiffusion >>
rect 269 429 270 430 
<< pdiffusion >>
rect 282 429 283 430 
<< pdiffusion >>
rect 283 429 284 430 
<< pdiffusion >>
rect 284 429 285 430 
<< pdiffusion >>
rect 285 429 286 430 
<< pdiffusion >>
rect 286 429 287 430 
<< pdiffusion >>
rect 287 429 288 430 
<< m1 >>
rect 289 429 290 430 
<< pdiffusion >>
rect 300 429 301 430 
<< pdiffusion >>
rect 301 429 302 430 
<< pdiffusion >>
rect 302 429 303 430 
<< pdiffusion >>
rect 303 429 304 430 
<< pdiffusion >>
rect 304 429 305 430 
<< pdiffusion >>
rect 305 429 306 430 
<< m1 >>
rect 307 429 308 430 
<< pdiffusion >>
rect 318 429 319 430 
<< pdiffusion >>
rect 319 429 320 430 
<< pdiffusion >>
rect 320 429 321 430 
<< pdiffusion >>
rect 321 429 322 430 
<< pdiffusion >>
rect 322 429 323 430 
<< pdiffusion >>
rect 323 429 324 430 
<< pdiffusion >>
rect 336 429 337 430 
<< pdiffusion >>
rect 337 429 338 430 
<< pdiffusion >>
rect 338 429 339 430 
<< pdiffusion >>
rect 339 429 340 430 
<< pdiffusion >>
rect 340 429 341 430 
<< pdiffusion >>
rect 341 429 342 430 
<< pdiffusion >>
rect 354 429 355 430 
<< pdiffusion >>
rect 355 429 356 430 
<< pdiffusion >>
rect 356 429 357 430 
<< pdiffusion >>
rect 357 429 358 430 
<< pdiffusion >>
rect 358 429 359 430 
<< pdiffusion >>
rect 359 429 360 430 
<< pdiffusion >>
rect 372 429 373 430 
<< pdiffusion >>
rect 373 429 374 430 
<< pdiffusion >>
rect 374 429 375 430 
<< pdiffusion >>
rect 375 429 376 430 
<< pdiffusion >>
rect 376 429 377 430 
<< pdiffusion >>
rect 377 429 378 430 
<< pdiffusion >>
rect 390 429 391 430 
<< pdiffusion >>
rect 391 429 392 430 
<< pdiffusion >>
rect 392 429 393 430 
<< pdiffusion >>
rect 393 429 394 430 
<< pdiffusion >>
rect 394 429 395 430 
<< pdiffusion >>
rect 395 429 396 430 
<< pdiffusion >>
rect 408 429 409 430 
<< pdiffusion >>
rect 409 429 410 430 
<< pdiffusion >>
rect 410 429 411 430 
<< pdiffusion >>
rect 411 429 412 430 
<< pdiffusion >>
rect 412 429 413 430 
<< pdiffusion >>
rect 413 429 414 430 
<< pdiffusion >>
rect 426 429 427 430 
<< pdiffusion >>
rect 427 429 428 430 
<< pdiffusion >>
rect 428 429 429 430 
<< pdiffusion >>
rect 429 429 430 430 
<< pdiffusion >>
rect 430 429 431 430 
<< pdiffusion >>
rect 431 429 432 430 
<< pdiffusion >>
rect 444 429 445 430 
<< pdiffusion >>
rect 445 429 446 430 
<< pdiffusion >>
rect 446 429 447 430 
<< pdiffusion >>
rect 447 429 448 430 
<< pdiffusion >>
rect 448 429 449 430 
<< pdiffusion >>
rect 449 429 450 430 
<< pdiffusion >>
rect 12 430 13 431 
<< pdiffusion >>
rect 13 430 14 431 
<< pdiffusion >>
rect 14 430 15 431 
<< pdiffusion >>
rect 15 430 16 431 
<< pdiffusion >>
rect 16 430 17 431 
<< pdiffusion >>
rect 17 430 18 431 
<< pdiffusion >>
rect 30 430 31 431 
<< pdiffusion >>
rect 31 430 32 431 
<< pdiffusion >>
rect 32 430 33 431 
<< pdiffusion >>
rect 33 430 34 431 
<< pdiffusion >>
rect 34 430 35 431 
<< pdiffusion >>
rect 35 430 36 431 
<< m1 >>
rect 46 430 47 431 
<< pdiffusion >>
rect 48 430 49 431 
<< pdiffusion >>
rect 49 430 50 431 
<< pdiffusion >>
rect 50 430 51 431 
<< pdiffusion >>
rect 51 430 52 431 
<< pdiffusion >>
rect 52 430 53 431 
<< pdiffusion >>
rect 53 430 54 431 
<< m1 >>
rect 64 430 65 431 
<< pdiffusion >>
rect 66 430 67 431 
<< pdiffusion >>
rect 67 430 68 431 
<< pdiffusion >>
rect 68 430 69 431 
<< pdiffusion >>
rect 69 430 70 431 
<< pdiffusion >>
rect 70 430 71 431 
<< pdiffusion >>
rect 71 430 72 431 
<< pdiffusion >>
rect 84 430 85 431 
<< pdiffusion >>
rect 85 430 86 431 
<< pdiffusion >>
rect 86 430 87 431 
<< pdiffusion >>
rect 87 430 88 431 
<< pdiffusion >>
rect 88 430 89 431 
<< pdiffusion >>
rect 89 430 90 431 
<< pdiffusion >>
rect 120 430 121 431 
<< pdiffusion >>
rect 121 430 122 431 
<< pdiffusion >>
rect 122 430 123 431 
<< pdiffusion >>
rect 123 430 124 431 
<< pdiffusion >>
rect 124 430 125 431 
<< pdiffusion >>
rect 125 430 126 431 
<< pdiffusion >>
rect 138 430 139 431 
<< pdiffusion >>
rect 139 430 140 431 
<< pdiffusion >>
rect 140 430 141 431 
<< pdiffusion >>
rect 141 430 142 431 
<< pdiffusion >>
rect 142 430 143 431 
<< pdiffusion >>
rect 143 430 144 431 
<< m1 >>
rect 145 430 146 431 
<< m1 >>
rect 154 430 155 431 
<< pdiffusion >>
rect 156 430 157 431 
<< pdiffusion >>
rect 157 430 158 431 
<< pdiffusion >>
rect 158 430 159 431 
<< pdiffusion >>
rect 159 430 160 431 
<< pdiffusion >>
rect 160 430 161 431 
<< pdiffusion >>
rect 161 430 162 431 
<< pdiffusion >>
rect 174 430 175 431 
<< pdiffusion >>
rect 175 430 176 431 
<< pdiffusion >>
rect 176 430 177 431 
<< pdiffusion >>
rect 177 430 178 431 
<< pdiffusion >>
rect 178 430 179 431 
<< pdiffusion >>
rect 179 430 180 431 
<< pdiffusion >>
rect 192 430 193 431 
<< pdiffusion >>
rect 193 430 194 431 
<< pdiffusion >>
rect 194 430 195 431 
<< pdiffusion >>
rect 195 430 196 431 
<< pdiffusion >>
rect 196 430 197 431 
<< pdiffusion >>
rect 197 430 198 431 
<< pdiffusion >>
rect 210 430 211 431 
<< pdiffusion >>
rect 211 430 212 431 
<< pdiffusion >>
rect 212 430 213 431 
<< pdiffusion >>
rect 213 430 214 431 
<< pdiffusion >>
rect 214 430 215 431 
<< pdiffusion >>
rect 215 430 216 431 
<< m1 >>
rect 226 430 227 431 
<< pdiffusion >>
rect 228 430 229 431 
<< pdiffusion >>
rect 229 430 230 431 
<< pdiffusion >>
rect 230 430 231 431 
<< pdiffusion >>
rect 231 430 232 431 
<< pdiffusion >>
rect 232 430 233 431 
<< pdiffusion >>
rect 233 430 234 431 
<< pdiffusion >>
rect 246 430 247 431 
<< pdiffusion >>
rect 247 430 248 431 
<< pdiffusion >>
rect 248 430 249 431 
<< pdiffusion >>
rect 249 430 250 431 
<< pdiffusion >>
rect 250 430 251 431 
<< pdiffusion >>
rect 251 430 252 431 
<< pdiffusion >>
rect 264 430 265 431 
<< pdiffusion >>
rect 265 430 266 431 
<< pdiffusion >>
rect 266 430 267 431 
<< pdiffusion >>
rect 267 430 268 431 
<< pdiffusion >>
rect 268 430 269 431 
<< pdiffusion >>
rect 269 430 270 431 
<< pdiffusion >>
rect 282 430 283 431 
<< pdiffusion >>
rect 283 430 284 431 
<< pdiffusion >>
rect 284 430 285 431 
<< pdiffusion >>
rect 285 430 286 431 
<< pdiffusion >>
rect 286 430 287 431 
<< pdiffusion >>
rect 287 430 288 431 
<< m1 >>
rect 289 430 290 431 
<< pdiffusion >>
rect 300 430 301 431 
<< pdiffusion >>
rect 301 430 302 431 
<< pdiffusion >>
rect 302 430 303 431 
<< pdiffusion >>
rect 303 430 304 431 
<< pdiffusion >>
rect 304 430 305 431 
<< pdiffusion >>
rect 305 430 306 431 
<< m1 >>
rect 307 430 308 431 
<< pdiffusion >>
rect 318 430 319 431 
<< pdiffusion >>
rect 319 430 320 431 
<< pdiffusion >>
rect 320 430 321 431 
<< pdiffusion >>
rect 321 430 322 431 
<< pdiffusion >>
rect 322 430 323 431 
<< pdiffusion >>
rect 323 430 324 431 
<< pdiffusion >>
rect 336 430 337 431 
<< pdiffusion >>
rect 337 430 338 431 
<< pdiffusion >>
rect 338 430 339 431 
<< pdiffusion >>
rect 339 430 340 431 
<< pdiffusion >>
rect 340 430 341 431 
<< pdiffusion >>
rect 341 430 342 431 
<< pdiffusion >>
rect 354 430 355 431 
<< pdiffusion >>
rect 355 430 356 431 
<< pdiffusion >>
rect 356 430 357 431 
<< pdiffusion >>
rect 357 430 358 431 
<< pdiffusion >>
rect 358 430 359 431 
<< pdiffusion >>
rect 359 430 360 431 
<< pdiffusion >>
rect 372 430 373 431 
<< pdiffusion >>
rect 373 430 374 431 
<< pdiffusion >>
rect 374 430 375 431 
<< pdiffusion >>
rect 375 430 376 431 
<< pdiffusion >>
rect 376 430 377 431 
<< pdiffusion >>
rect 377 430 378 431 
<< pdiffusion >>
rect 390 430 391 431 
<< pdiffusion >>
rect 391 430 392 431 
<< pdiffusion >>
rect 392 430 393 431 
<< pdiffusion >>
rect 393 430 394 431 
<< pdiffusion >>
rect 394 430 395 431 
<< pdiffusion >>
rect 395 430 396 431 
<< pdiffusion >>
rect 408 430 409 431 
<< pdiffusion >>
rect 409 430 410 431 
<< pdiffusion >>
rect 410 430 411 431 
<< pdiffusion >>
rect 411 430 412 431 
<< pdiffusion >>
rect 412 430 413 431 
<< pdiffusion >>
rect 413 430 414 431 
<< pdiffusion >>
rect 426 430 427 431 
<< pdiffusion >>
rect 427 430 428 431 
<< pdiffusion >>
rect 428 430 429 431 
<< pdiffusion >>
rect 429 430 430 431 
<< pdiffusion >>
rect 430 430 431 431 
<< pdiffusion >>
rect 431 430 432 431 
<< pdiffusion >>
rect 444 430 445 431 
<< pdiffusion >>
rect 445 430 446 431 
<< pdiffusion >>
rect 446 430 447 431 
<< pdiffusion >>
rect 447 430 448 431 
<< pdiffusion >>
rect 448 430 449 431 
<< pdiffusion >>
rect 449 430 450 431 
<< pdiffusion >>
rect 12 431 13 432 
<< pdiffusion >>
rect 13 431 14 432 
<< pdiffusion >>
rect 14 431 15 432 
<< pdiffusion >>
rect 15 431 16 432 
<< pdiffusion >>
rect 16 431 17 432 
<< pdiffusion >>
rect 17 431 18 432 
<< pdiffusion >>
rect 30 431 31 432 
<< pdiffusion >>
rect 31 431 32 432 
<< pdiffusion >>
rect 32 431 33 432 
<< pdiffusion >>
rect 33 431 34 432 
<< pdiffusion >>
rect 34 431 35 432 
<< pdiffusion >>
rect 35 431 36 432 
<< m1 >>
rect 46 431 47 432 
<< pdiffusion >>
rect 48 431 49 432 
<< pdiffusion >>
rect 49 431 50 432 
<< pdiffusion >>
rect 50 431 51 432 
<< pdiffusion >>
rect 51 431 52 432 
<< pdiffusion >>
rect 52 431 53 432 
<< pdiffusion >>
rect 53 431 54 432 
<< m1 >>
rect 64 431 65 432 
<< pdiffusion >>
rect 66 431 67 432 
<< m1 >>
rect 67 431 68 432 
<< pdiffusion >>
rect 67 431 68 432 
<< pdiffusion >>
rect 68 431 69 432 
<< pdiffusion >>
rect 69 431 70 432 
<< pdiffusion >>
rect 70 431 71 432 
<< pdiffusion >>
rect 71 431 72 432 
<< pdiffusion >>
rect 84 431 85 432 
<< pdiffusion >>
rect 85 431 86 432 
<< pdiffusion >>
rect 86 431 87 432 
<< pdiffusion >>
rect 87 431 88 432 
<< pdiffusion >>
rect 88 431 89 432 
<< pdiffusion >>
rect 89 431 90 432 
<< pdiffusion >>
rect 120 431 121 432 
<< pdiffusion >>
rect 121 431 122 432 
<< pdiffusion >>
rect 122 431 123 432 
<< pdiffusion >>
rect 123 431 124 432 
<< pdiffusion >>
rect 124 431 125 432 
<< pdiffusion >>
rect 125 431 126 432 
<< pdiffusion >>
rect 138 431 139 432 
<< pdiffusion >>
rect 139 431 140 432 
<< pdiffusion >>
rect 140 431 141 432 
<< pdiffusion >>
rect 141 431 142 432 
<< pdiffusion >>
rect 142 431 143 432 
<< pdiffusion >>
rect 143 431 144 432 
<< m1 >>
rect 145 431 146 432 
<< m1 >>
rect 154 431 155 432 
<< pdiffusion >>
rect 156 431 157 432 
<< pdiffusion >>
rect 157 431 158 432 
<< pdiffusion >>
rect 158 431 159 432 
<< pdiffusion >>
rect 159 431 160 432 
<< pdiffusion >>
rect 160 431 161 432 
<< pdiffusion >>
rect 161 431 162 432 
<< pdiffusion >>
rect 174 431 175 432 
<< pdiffusion >>
rect 175 431 176 432 
<< pdiffusion >>
rect 176 431 177 432 
<< pdiffusion >>
rect 177 431 178 432 
<< pdiffusion >>
rect 178 431 179 432 
<< pdiffusion >>
rect 179 431 180 432 
<< pdiffusion >>
rect 192 431 193 432 
<< pdiffusion >>
rect 193 431 194 432 
<< pdiffusion >>
rect 194 431 195 432 
<< pdiffusion >>
rect 195 431 196 432 
<< pdiffusion >>
rect 196 431 197 432 
<< pdiffusion >>
rect 197 431 198 432 
<< pdiffusion >>
rect 210 431 211 432 
<< pdiffusion >>
rect 211 431 212 432 
<< pdiffusion >>
rect 212 431 213 432 
<< pdiffusion >>
rect 213 431 214 432 
<< pdiffusion >>
rect 214 431 215 432 
<< pdiffusion >>
rect 215 431 216 432 
<< m1 >>
rect 226 431 227 432 
<< pdiffusion >>
rect 228 431 229 432 
<< pdiffusion >>
rect 229 431 230 432 
<< pdiffusion >>
rect 230 431 231 432 
<< pdiffusion >>
rect 231 431 232 432 
<< pdiffusion >>
rect 232 431 233 432 
<< pdiffusion >>
rect 233 431 234 432 
<< pdiffusion >>
rect 246 431 247 432 
<< pdiffusion >>
rect 247 431 248 432 
<< pdiffusion >>
rect 248 431 249 432 
<< pdiffusion >>
rect 249 431 250 432 
<< pdiffusion >>
rect 250 431 251 432 
<< pdiffusion >>
rect 251 431 252 432 
<< pdiffusion >>
rect 264 431 265 432 
<< pdiffusion >>
rect 265 431 266 432 
<< pdiffusion >>
rect 266 431 267 432 
<< pdiffusion >>
rect 267 431 268 432 
<< pdiffusion >>
rect 268 431 269 432 
<< pdiffusion >>
rect 269 431 270 432 
<< pdiffusion >>
rect 282 431 283 432 
<< pdiffusion >>
rect 283 431 284 432 
<< pdiffusion >>
rect 284 431 285 432 
<< pdiffusion >>
rect 285 431 286 432 
<< pdiffusion >>
rect 286 431 287 432 
<< pdiffusion >>
rect 287 431 288 432 
<< m1 >>
rect 289 431 290 432 
<< pdiffusion >>
rect 300 431 301 432 
<< pdiffusion >>
rect 301 431 302 432 
<< pdiffusion >>
rect 302 431 303 432 
<< pdiffusion >>
rect 303 431 304 432 
<< pdiffusion >>
rect 304 431 305 432 
<< pdiffusion >>
rect 305 431 306 432 
<< m1 >>
rect 307 431 308 432 
<< pdiffusion >>
rect 318 431 319 432 
<< pdiffusion >>
rect 319 431 320 432 
<< pdiffusion >>
rect 320 431 321 432 
<< pdiffusion >>
rect 321 431 322 432 
<< pdiffusion >>
rect 322 431 323 432 
<< pdiffusion >>
rect 323 431 324 432 
<< pdiffusion >>
rect 336 431 337 432 
<< pdiffusion >>
rect 337 431 338 432 
<< pdiffusion >>
rect 338 431 339 432 
<< pdiffusion >>
rect 339 431 340 432 
<< m1 >>
rect 340 431 341 432 
<< pdiffusion >>
rect 340 431 341 432 
<< pdiffusion >>
rect 341 431 342 432 
<< pdiffusion >>
rect 354 431 355 432 
<< pdiffusion >>
rect 355 431 356 432 
<< pdiffusion >>
rect 356 431 357 432 
<< pdiffusion >>
rect 357 431 358 432 
<< pdiffusion >>
rect 358 431 359 432 
<< pdiffusion >>
rect 359 431 360 432 
<< pdiffusion >>
rect 372 431 373 432 
<< pdiffusion >>
rect 373 431 374 432 
<< pdiffusion >>
rect 374 431 375 432 
<< pdiffusion >>
rect 375 431 376 432 
<< pdiffusion >>
rect 376 431 377 432 
<< pdiffusion >>
rect 377 431 378 432 
<< pdiffusion >>
rect 390 431 391 432 
<< pdiffusion >>
rect 391 431 392 432 
<< pdiffusion >>
rect 392 431 393 432 
<< pdiffusion >>
rect 393 431 394 432 
<< pdiffusion >>
rect 394 431 395 432 
<< pdiffusion >>
rect 395 431 396 432 
<< pdiffusion >>
rect 408 431 409 432 
<< pdiffusion >>
rect 409 431 410 432 
<< pdiffusion >>
rect 410 431 411 432 
<< pdiffusion >>
rect 411 431 412 432 
<< pdiffusion >>
rect 412 431 413 432 
<< pdiffusion >>
rect 413 431 414 432 
<< pdiffusion >>
rect 426 431 427 432 
<< pdiffusion >>
rect 427 431 428 432 
<< pdiffusion >>
rect 428 431 429 432 
<< pdiffusion >>
rect 429 431 430 432 
<< pdiffusion >>
rect 430 431 431 432 
<< pdiffusion >>
rect 431 431 432 432 
<< pdiffusion >>
rect 444 431 445 432 
<< pdiffusion >>
rect 445 431 446 432 
<< pdiffusion >>
rect 446 431 447 432 
<< pdiffusion >>
rect 447 431 448 432 
<< pdiffusion >>
rect 448 431 449 432 
<< pdiffusion >>
rect 449 431 450 432 
<< m1 >>
rect 46 432 47 433 
<< m1 >>
rect 64 432 65 433 
<< m1 >>
rect 67 432 68 433 
<< m1 >>
rect 145 432 146 433 
<< m1 >>
rect 154 432 155 433 
<< m1 >>
rect 226 432 227 433 
<< m1 >>
rect 289 432 290 433 
<< m1 >>
rect 307 432 308 433 
<< m1 >>
rect 340 432 341 433 
<< m1 >>
rect 46 433 47 434 
<< m1 >>
rect 64 433 65 434 
<< m1 >>
rect 65 433 66 434 
<< m1 >>
rect 66 433 67 434 
<< m1 >>
rect 67 433 68 434 
<< m1 >>
rect 145 433 146 434 
<< m1 >>
rect 154 433 155 434 
<< m1 >>
rect 226 433 227 434 
<< m1 >>
rect 289 433 290 434 
<< m1 >>
rect 307 433 308 434 
<< m1 >>
rect 340 433 341 434 
<< m1 >>
rect 341 433 342 434 
<< m1 >>
rect 342 433 343 434 
<< m1 >>
rect 343 433 344 434 
<< m1 >>
rect 46 434 47 435 
<< m1 >>
rect 145 434 146 435 
<< m1 >>
rect 154 434 155 435 
<< m1 >>
rect 226 434 227 435 
<< m1 >>
rect 289 434 290 435 
<< m1 >>
rect 307 434 308 435 
<< m1 >>
rect 343 434 344 435 
<< m1 >>
rect 46 435 47 436 
<< m1 >>
rect 145 435 146 436 
<< m1 >>
rect 154 435 155 436 
<< m1 >>
rect 226 435 227 436 
<< m1 >>
rect 289 435 290 436 
<< m1 >>
rect 307 435 308 436 
<< m1 >>
rect 343 435 344 436 
<< m1 >>
rect 13 436 14 437 
<< m1 >>
rect 14 436 15 437 
<< m1 >>
rect 15 436 16 437 
<< m1 >>
rect 16 436 17 437 
<< m1 >>
rect 17 436 18 437 
<< m1 >>
rect 18 436 19 437 
<< m1 >>
rect 19 436 20 437 
<< m1 >>
rect 20 436 21 437 
<< m1 >>
rect 21 436 22 437 
<< m1 >>
rect 22 436 23 437 
<< m1 >>
rect 23 436 24 437 
<< m1 >>
rect 24 436 25 437 
<< m1 >>
rect 25 436 26 437 
<< m1 >>
rect 26 436 27 437 
<< m1 >>
rect 27 436 28 437 
<< m1 >>
rect 28 436 29 437 
<< m1 >>
rect 29 436 30 437 
<< m1 >>
rect 30 436 31 437 
<< m1 >>
rect 31 436 32 437 
<< m1 >>
rect 32 436 33 437 
<< m1 >>
rect 33 436 34 437 
<< m1 >>
rect 34 436 35 437 
<< m1 >>
rect 35 436 36 437 
<< m1 >>
rect 36 436 37 437 
<< m1 >>
rect 37 436 38 437 
<< m1 >>
rect 38 436 39 437 
<< m1 >>
rect 39 436 40 437 
<< m1 >>
rect 40 436 41 437 
<< m1 >>
rect 41 436 42 437 
<< m1 >>
rect 42 436 43 437 
<< m1 >>
rect 43 436 44 437 
<< m1 >>
rect 44 436 45 437 
<< m1 >>
rect 45 436 46 437 
<< m1 >>
rect 46 436 47 437 
<< m1 >>
rect 145 436 146 437 
<< m1 >>
rect 154 436 155 437 
<< m1 >>
rect 226 436 227 437 
<< m1 >>
rect 289 436 290 437 
<< m1 >>
rect 307 436 308 437 
<< m1 >>
rect 343 436 344 437 
<< m1 >>
rect 13 437 14 438 
<< m1 >>
rect 145 437 146 438 
<< m1 >>
rect 154 437 155 438 
<< m1 >>
rect 226 437 227 438 
<< m1 >>
rect 289 437 290 438 
<< m1 >>
rect 307 437 308 438 
<< m1 >>
rect 343 437 344 438 
<< m1 >>
rect 13 438 14 439 
<< m1 >>
rect 145 438 146 439 
<< m1 >>
rect 154 438 155 439 
<< m1 >>
rect 226 438 227 439 
<< m1 >>
rect 289 438 290 439 
<< m1 >>
rect 307 438 308 439 
<< m1 >>
rect 343 438 344 439 
<< m1 >>
rect 13 439 14 440 
<< m1 >>
rect 145 439 146 440 
<< m1 >>
rect 154 439 155 440 
<< m1 >>
rect 155 439 156 440 
<< m1 >>
rect 156 439 157 440 
<< m1 >>
rect 157 439 158 440 
<< m1 >>
rect 158 439 159 440 
<< m1 >>
rect 159 439 160 440 
<< m1 >>
rect 160 439 161 440 
<< m1 >>
rect 161 439 162 440 
<< m1 >>
rect 162 439 163 440 
<< m1 >>
rect 163 439 164 440 
<< m1 >>
rect 164 439 165 440 
<< m1 >>
rect 165 439 166 440 
<< m1 >>
rect 166 439 167 440 
<< m1 >>
rect 167 439 168 440 
<< m1 >>
rect 168 439 169 440 
<< m1 >>
rect 169 439 170 440 
<< m1 >>
rect 170 439 171 440 
<< m1 >>
rect 171 439 172 440 
<< m1 >>
rect 172 439 173 440 
<< m1 >>
rect 226 439 227 440 
<< m1 >>
rect 283 439 284 440 
<< m1 >>
rect 284 439 285 440 
<< m1 >>
rect 285 439 286 440 
<< m1 >>
rect 286 439 287 440 
<< m1 >>
rect 287 439 288 440 
<< m2 >>
rect 287 439 288 440 
<< m2c >>
rect 287 439 288 440 
<< m1 >>
rect 287 439 288 440 
<< m2 >>
rect 287 439 288 440 
<< m2 >>
rect 288 439 289 440 
<< m1 >>
rect 289 439 290 440 
<< m2 >>
rect 289 439 290 440 
<< m2 >>
rect 290 439 291 440 
<< m1 >>
rect 291 439 292 440 
<< m2 >>
rect 291 439 292 440 
<< m2c >>
rect 291 439 292 440 
<< m1 >>
rect 291 439 292 440 
<< m2 >>
rect 291 439 292 440 
<< m1 >>
rect 292 439 293 440 
<< m1 >>
rect 293 439 294 440 
<< m1 >>
rect 294 439 295 440 
<< m1 >>
rect 295 439 296 440 
<< m1 >>
rect 296 439 297 440 
<< m1 >>
rect 297 439 298 440 
<< m1 >>
rect 298 439 299 440 
<< m1 >>
rect 299 439 300 440 
<< m1 >>
rect 300 439 301 440 
<< m1 >>
rect 301 439 302 440 
<< m1 >>
rect 302 439 303 440 
<< m1 >>
rect 303 439 304 440 
<< m1 >>
rect 304 439 305 440 
<< m1 >>
rect 307 439 308 440 
<< m1 >>
rect 343 439 344 440 
<< m1 >>
rect 13 440 14 441 
<< m1 >>
rect 145 440 146 441 
<< m1 >>
rect 172 440 173 441 
<< m1 >>
rect 226 440 227 441 
<< m1 >>
rect 283 440 284 441 
<< m1 >>
rect 289 440 290 441 
<< m1 >>
rect 304 440 305 441 
<< m1 >>
rect 307 440 308 441 
<< m1 >>
rect 343 440 344 441 
<< m1 >>
rect 13 441 14 442 
<< m1 >>
rect 145 441 146 442 
<< m1 >>
rect 172 441 173 442 
<< m1 >>
rect 226 441 227 442 
<< m1 >>
rect 283 441 284 442 
<< m1 >>
rect 289 441 290 442 
<< m1 >>
rect 304 441 305 442 
<< m1 >>
rect 307 441 308 442 
<< m1 >>
rect 343 441 344 442 
<< m1 >>
rect 13 442 14 443 
<< m1 >>
rect 142 442 143 443 
<< m1 >>
rect 143 442 144 443 
<< m1 >>
rect 144 442 145 443 
<< m1 >>
rect 145 442 146 443 
<< m1 >>
rect 172 442 173 443 
<< m1 >>
rect 226 442 227 443 
<< m1 >>
rect 283 442 284 443 
<< m1 >>
rect 289 442 290 443 
<< m1 >>
rect 304 442 305 443 
<< m1 >>
rect 307 442 308 443 
<< m1 >>
rect 343 442 344 443 
<< m1 >>
rect 13 443 14 444 
<< m1 >>
rect 142 443 143 444 
<< m1 >>
rect 172 443 173 444 
<< m1 >>
rect 226 443 227 444 
<< m1 >>
rect 283 443 284 444 
<< m1 >>
rect 289 443 290 444 
<< m1 >>
rect 304 443 305 444 
<< m1 >>
rect 307 443 308 444 
<< m1 >>
rect 343 443 344 444 
<< pdiffusion >>
rect 12 444 13 445 
<< m1 >>
rect 13 444 14 445 
<< pdiffusion >>
rect 13 444 14 445 
<< pdiffusion >>
rect 14 444 15 445 
<< pdiffusion >>
rect 15 444 16 445 
<< pdiffusion >>
rect 16 444 17 445 
<< pdiffusion >>
rect 17 444 18 445 
<< pdiffusion >>
rect 30 444 31 445 
<< pdiffusion >>
rect 31 444 32 445 
<< pdiffusion >>
rect 32 444 33 445 
<< pdiffusion >>
rect 33 444 34 445 
<< pdiffusion >>
rect 34 444 35 445 
<< pdiffusion >>
rect 35 444 36 445 
<< pdiffusion >>
rect 48 444 49 445 
<< pdiffusion >>
rect 49 444 50 445 
<< pdiffusion >>
rect 50 444 51 445 
<< pdiffusion >>
rect 51 444 52 445 
<< pdiffusion >>
rect 52 444 53 445 
<< pdiffusion >>
rect 53 444 54 445 
<< pdiffusion >>
rect 66 444 67 445 
<< pdiffusion >>
rect 67 444 68 445 
<< pdiffusion >>
rect 68 444 69 445 
<< pdiffusion >>
rect 69 444 70 445 
<< pdiffusion >>
rect 70 444 71 445 
<< pdiffusion >>
rect 71 444 72 445 
<< pdiffusion >>
rect 84 444 85 445 
<< pdiffusion >>
rect 85 444 86 445 
<< pdiffusion >>
rect 86 444 87 445 
<< pdiffusion >>
rect 87 444 88 445 
<< pdiffusion >>
rect 88 444 89 445 
<< pdiffusion >>
rect 89 444 90 445 
<< pdiffusion >>
rect 102 444 103 445 
<< pdiffusion >>
rect 103 444 104 445 
<< pdiffusion >>
rect 104 444 105 445 
<< pdiffusion >>
rect 105 444 106 445 
<< pdiffusion >>
rect 106 444 107 445 
<< pdiffusion >>
rect 107 444 108 445 
<< pdiffusion >>
rect 120 444 121 445 
<< pdiffusion >>
rect 121 444 122 445 
<< pdiffusion >>
rect 122 444 123 445 
<< pdiffusion >>
rect 123 444 124 445 
<< pdiffusion >>
rect 124 444 125 445 
<< pdiffusion >>
rect 125 444 126 445 
<< pdiffusion >>
rect 138 444 139 445 
<< pdiffusion >>
rect 139 444 140 445 
<< pdiffusion >>
rect 140 444 141 445 
<< pdiffusion >>
rect 141 444 142 445 
<< m1 >>
rect 142 444 143 445 
<< pdiffusion >>
rect 142 444 143 445 
<< pdiffusion >>
rect 143 444 144 445 
<< pdiffusion >>
rect 156 444 157 445 
<< pdiffusion >>
rect 157 444 158 445 
<< pdiffusion >>
rect 158 444 159 445 
<< pdiffusion >>
rect 159 444 160 445 
<< pdiffusion >>
rect 160 444 161 445 
<< pdiffusion >>
rect 161 444 162 445 
<< m1 >>
rect 172 444 173 445 
<< pdiffusion >>
rect 174 444 175 445 
<< pdiffusion >>
rect 175 444 176 445 
<< pdiffusion >>
rect 176 444 177 445 
<< pdiffusion >>
rect 177 444 178 445 
<< pdiffusion >>
rect 178 444 179 445 
<< pdiffusion >>
rect 179 444 180 445 
<< pdiffusion >>
rect 192 444 193 445 
<< pdiffusion >>
rect 193 444 194 445 
<< pdiffusion >>
rect 194 444 195 445 
<< pdiffusion >>
rect 195 444 196 445 
<< pdiffusion >>
rect 196 444 197 445 
<< pdiffusion >>
rect 197 444 198 445 
<< pdiffusion >>
rect 210 444 211 445 
<< pdiffusion >>
rect 211 444 212 445 
<< pdiffusion >>
rect 212 444 213 445 
<< pdiffusion >>
rect 213 444 214 445 
<< pdiffusion >>
rect 214 444 215 445 
<< pdiffusion >>
rect 215 444 216 445 
<< m1 >>
rect 226 444 227 445 
<< pdiffusion >>
rect 228 444 229 445 
<< pdiffusion >>
rect 229 444 230 445 
<< pdiffusion >>
rect 230 444 231 445 
<< pdiffusion >>
rect 231 444 232 445 
<< pdiffusion >>
rect 232 444 233 445 
<< pdiffusion >>
rect 233 444 234 445 
<< pdiffusion >>
rect 246 444 247 445 
<< pdiffusion >>
rect 247 444 248 445 
<< pdiffusion >>
rect 248 444 249 445 
<< pdiffusion >>
rect 249 444 250 445 
<< pdiffusion >>
rect 250 444 251 445 
<< pdiffusion >>
rect 251 444 252 445 
<< pdiffusion >>
rect 264 444 265 445 
<< pdiffusion >>
rect 265 444 266 445 
<< pdiffusion >>
rect 266 444 267 445 
<< pdiffusion >>
rect 267 444 268 445 
<< pdiffusion >>
rect 268 444 269 445 
<< pdiffusion >>
rect 269 444 270 445 
<< pdiffusion >>
rect 282 444 283 445 
<< m1 >>
rect 283 444 284 445 
<< pdiffusion >>
rect 283 444 284 445 
<< pdiffusion >>
rect 284 444 285 445 
<< pdiffusion >>
rect 285 444 286 445 
<< pdiffusion >>
rect 286 444 287 445 
<< pdiffusion >>
rect 287 444 288 445 
<< m1 >>
rect 289 444 290 445 
<< pdiffusion >>
rect 300 444 301 445 
<< pdiffusion >>
rect 301 444 302 445 
<< pdiffusion >>
rect 302 444 303 445 
<< pdiffusion >>
rect 303 444 304 445 
<< m1 >>
rect 304 444 305 445 
<< pdiffusion >>
rect 304 444 305 445 
<< pdiffusion >>
rect 305 444 306 445 
<< m1 >>
rect 307 444 308 445 
<< pdiffusion >>
rect 318 444 319 445 
<< pdiffusion >>
rect 319 444 320 445 
<< pdiffusion >>
rect 320 444 321 445 
<< pdiffusion >>
rect 321 444 322 445 
<< pdiffusion >>
rect 322 444 323 445 
<< pdiffusion >>
rect 323 444 324 445 
<< pdiffusion >>
rect 336 444 337 445 
<< pdiffusion >>
rect 337 444 338 445 
<< pdiffusion >>
rect 338 444 339 445 
<< pdiffusion >>
rect 339 444 340 445 
<< pdiffusion >>
rect 340 444 341 445 
<< pdiffusion >>
rect 341 444 342 445 
<< m1 >>
rect 343 444 344 445 
<< pdiffusion >>
rect 354 444 355 445 
<< pdiffusion >>
rect 355 444 356 445 
<< pdiffusion >>
rect 356 444 357 445 
<< pdiffusion >>
rect 357 444 358 445 
<< pdiffusion >>
rect 358 444 359 445 
<< pdiffusion >>
rect 359 444 360 445 
<< pdiffusion >>
rect 372 444 373 445 
<< pdiffusion >>
rect 373 444 374 445 
<< pdiffusion >>
rect 374 444 375 445 
<< pdiffusion >>
rect 375 444 376 445 
<< pdiffusion >>
rect 376 444 377 445 
<< pdiffusion >>
rect 377 444 378 445 
<< pdiffusion >>
rect 390 444 391 445 
<< pdiffusion >>
rect 391 444 392 445 
<< pdiffusion >>
rect 392 444 393 445 
<< pdiffusion >>
rect 393 444 394 445 
<< pdiffusion >>
rect 394 444 395 445 
<< pdiffusion >>
rect 395 444 396 445 
<< pdiffusion >>
rect 408 444 409 445 
<< pdiffusion >>
rect 409 444 410 445 
<< pdiffusion >>
rect 410 444 411 445 
<< pdiffusion >>
rect 411 444 412 445 
<< pdiffusion >>
rect 412 444 413 445 
<< pdiffusion >>
rect 413 444 414 445 
<< pdiffusion >>
rect 426 444 427 445 
<< pdiffusion >>
rect 427 444 428 445 
<< pdiffusion >>
rect 428 444 429 445 
<< pdiffusion >>
rect 429 444 430 445 
<< pdiffusion >>
rect 430 444 431 445 
<< pdiffusion >>
rect 431 444 432 445 
<< pdiffusion >>
rect 444 444 445 445 
<< pdiffusion >>
rect 445 444 446 445 
<< pdiffusion >>
rect 446 444 447 445 
<< pdiffusion >>
rect 447 444 448 445 
<< pdiffusion >>
rect 448 444 449 445 
<< pdiffusion >>
rect 449 444 450 445 
<< pdiffusion >>
rect 12 445 13 446 
<< pdiffusion >>
rect 13 445 14 446 
<< pdiffusion >>
rect 14 445 15 446 
<< pdiffusion >>
rect 15 445 16 446 
<< pdiffusion >>
rect 16 445 17 446 
<< pdiffusion >>
rect 17 445 18 446 
<< pdiffusion >>
rect 30 445 31 446 
<< pdiffusion >>
rect 31 445 32 446 
<< pdiffusion >>
rect 32 445 33 446 
<< pdiffusion >>
rect 33 445 34 446 
<< pdiffusion >>
rect 34 445 35 446 
<< pdiffusion >>
rect 35 445 36 446 
<< pdiffusion >>
rect 48 445 49 446 
<< pdiffusion >>
rect 49 445 50 446 
<< pdiffusion >>
rect 50 445 51 446 
<< pdiffusion >>
rect 51 445 52 446 
<< pdiffusion >>
rect 52 445 53 446 
<< pdiffusion >>
rect 53 445 54 446 
<< pdiffusion >>
rect 66 445 67 446 
<< pdiffusion >>
rect 67 445 68 446 
<< pdiffusion >>
rect 68 445 69 446 
<< pdiffusion >>
rect 69 445 70 446 
<< pdiffusion >>
rect 70 445 71 446 
<< pdiffusion >>
rect 71 445 72 446 
<< pdiffusion >>
rect 84 445 85 446 
<< pdiffusion >>
rect 85 445 86 446 
<< pdiffusion >>
rect 86 445 87 446 
<< pdiffusion >>
rect 87 445 88 446 
<< pdiffusion >>
rect 88 445 89 446 
<< pdiffusion >>
rect 89 445 90 446 
<< pdiffusion >>
rect 102 445 103 446 
<< pdiffusion >>
rect 103 445 104 446 
<< pdiffusion >>
rect 104 445 105 446 
<< pdiffusion >>
rect 105 445 106 446 
<< pdiffusion >>
rect 106 445 107 446 
<< pdiffusion >>
rect 107 445 108 446 
<< pdiffusion >>
rect 120 445 121 446 
<< pdiffusion >>
rect 121 445 122 446 
<< pdiffusion >>
rect 122 445 123 446 
<< pdiffusion >>
rect 123 445 124 446 
<< pdiffusion >>
rect 124 445 125 446 
<< pdiffusion >>
rect 125 445 126 446 
<< pdiffusion >>
rect 138 445 139 446 
<< pdiffusion >>
rect 139 445 140 446 
<< pdiffusion >>
rect 140 445 141 446 
<< pdiffusion >>
rect 141 445 142 446 
<< pdiffusion >>
rect 142 445 143 446 
<< pdiffusion >>
rect 143 445 144 446 
<< pdiffusion >>
rect 156 445 157 446 
<< pdiffusion >>
rect 157 445 158 446 
<< pdiffusion >>
rect 158 445 159 446 
<< pdiffusion >>
rect 159 445 160 446 
<< pdiffusion >>
rect 160 445 161 446 
<< pdiffusion >>
rect 161 445 162 446 
<< m1 >>
rect 172 445 173 446 
<< pdiffusion >>
rect 174 445 175 446 
<< pdiffusion >>
rect 175 445 176 446 
<< pdiffusion >>
rect 176 445 177 446 
<< pdiffusion >>
rect 177 445 178 446 
<< pdiffusion >>
rect 178 445 179 446 
<< pdiffusion >>
rect 179 445 180 446 
<< pdiffusion >>
rect 192 445 193 446 
<< pdiffusion >>
rect 193 445 194 446 
<< pdiffusion >>
rect 194 445 195 446 
<< pdiffusion >>
rect 195 445 196 446 
<< pdiffusion >>
rect 196 445 197 446 
<< pdiffusion >>
rect 197 445 198 446 
<< pdiffusion >>
rect 210 445 211 446 
<< pdiffusion >>
rect 211 445 212 446 
<< pdiffusion >>
rect 212 445 213 446 
<< pdiffusion >>
rect 213 445 214 446 
<< pdiffusion >>
rect 214 445 215 446 
<< pdiffusion >>
rect 215 445 216 446 
<< m1 >>
rect 226 445 227 446 
<< pdiffusion >>
rect 228 445 229 446 
<< pdiffusion >>
rect 229 445 230 446 
<< pdiffusion >>
rect 230 445 231 446 
<< pdiffusion >>
rect 231 445 232 446 
<< pdiffusion >>
rect 232 445 233 446 
<< pdiffusion >>
rect 233 445 234 446 
<< pdiffusion >>
rect 246 445 247 446 
<< pdiffusion >>
rect 247 445 248 446 
<< pdiffusion >>
rect 248 445 249 446 
<< pdiffusion >>
rect 249 445 250 446 
<< pdiffusion >>
rect 250 445 251 446 
<< pdiffusion >>
rect 251 445 252 446 
<< pdiffusion >>
rect 264 445 265 446 
<< pdiffusion >>
rect 265 445 266 446 
<< pdiffusion >>
rect 266 445 267 446 
<< pdiffusion >>
rect 267 445 268 446 
<< pdiffusion >>
rect 268 445 269 446 
<< pdiffusion >>
rect 269 445 270 446 
<< pdiffusion >>
rect 282 445 283 446 
<< pdiffusion >>
rect 283 445 284 446 
<< pdiffusion >>
rect 284 445 285 446 
<< pdiffusion >>
rect 285 445 286 446 
<< pdiffusion >>
rect 286 445 287 446 
<< pdiffusion >>
rect 287 445 288 446 
<< m1 >>
rect 289 445 290 446 
<< pdiffusion >>
rect 300 445 301 446 
<< pdiffusion >>
rect 301 445 302 446 
<< pdiffusion >>
rect 302 445 303 446 
<< pdiffusion >>
rect 303 445 304 446 
<< pdiffusion >>
rect 304 445 305 446 
<< pdiffusion >>
rect 305 445 306 446 
<< m1 >>
rect 307 445 308 446 
<< pdiffusion >>
rect 318 445 319 446 
<< pdiffusion >>
rect 319 445 320 446 
<< pdiffusion >>
rect 320 445 321 446 
<< pdiffusion >>
rect 321 445 322 446 
<< pdiffusion >>
rect 322 445 323 446 
<< pdiffusion >>
rect 323 445 324 446 
<< pdiffusion >>
rect 336 445 337 446 
<< pdiffusion >>
rect 337 445 338 446 
<< pdiffusion >>
rect 338 445 339 446 
<< pdiffusion >>
rect 339 445 340 446 
<< pdiffusion >>
rect 340 445 341 446 
<< pdiffusion >>
rect 341 445 342 446 
<< m1 >>
rect 343 445 344 446 
<< pdiffusion >>
rect 354 445 355 446 
<< pdiffusion >>
rect 355 445 356 446 
<< pdiffusion >>
rect 356 445 357 446 
<< pdiffusion >>
rect 357 445 358 446 
<< pdiffusion >>
rect 358 445 359 446 
<< pdiffusion >>
rect 359 445 360 446 
<< pdiffusion >>
rect 372 445 373 446 
<< pdiffusion >>
rect 373 445 374 446 
<< pdiffusion >>
rect 374 445 375 446 
<< pdiffusion >>
rect 375 445 376 446 
<< pdiffusion >>
rect 376 445 377 446 
<< pdiffusion >>
rect 377 445 378 446 
<< pdiffusion >>
rect 390 445 391 446 
<< pdiffusion >>
rect 391 445 392 446 
<< pdiffusion >>
rect 392 445 393 446 
<< pdiffusion >>
rect 393 445 394 446 
<< pdiffusion >>
rect 394 445 395 446 
<< pdiffusion >>
rect 395 445 396 446 
<< pdiffusion >>
rect 408 445 409 446 
<< pdiffusion >>
rect 409 445 410 446 
<< pdiffusion >>
rect 410 445 411 446 
<< pdiffusion >>
rect 411 445 412 446 
<< pdiffusion >>
rect 412 445 413 446 
<< pdiffusion >>
rect 413 445 414 446 
<< pdiffusion >>
rect 426 445 427 446 
<< pdiffusion >>
rect 427 445 428 446 
<< pdiffusion >>
rect 428 445 429 446 
<< pdiffusion >>
rect 429 445 430 446 
<< pdiffusion >>
rect 430 445 431 446 
<< pdiffusion >>
rect 431 445 432 446 
<< pdiffusion >>
rect 444 445 445 446 
<< pdiffusion >>
rect 445 445 446 446 
<< pdiffusion >>
rect 446 445 447 446 
<< pdiffusion >>
rect 447 445 448 446 
<< pdiffusion >>
rect 448 445 449 446 
<< pdiffusion >>
rect 449 445 450 446 
<< pdiffusion >>
rect 12 446 13 447 
<< pdiffusion >>
rect 13 446 14 447 
<< pdiffusion >>
rect 14 446 15 447 
<< pdiffusion >>
rect 15 446 16 447 
<< pdiffusion >>
rect 16 446 17 447 
<< pdiffusion >>
rect 17 446 18 447 
<< pdiffusion >>
rect 30 446 31 447 
<< pdiffusion >>
rect 31 446 32 447 
<< pdiffusion >>
rect 32 446 33 447 
<< pdiffusion >>
rect 33 446 34 447 
<< pdiffusion >>
rect 34 446 35 447 
<< pdiffusion >>
rect 35 446 36 447 
<< pdiffusion >>
rect 48 446 49 447 
<< pdiffusion >>
rect 49 446 50 447 
<< pdiffusion >>
rect 50 446 51 447 
<< pdiffusion >>
rect 51 446 52 447 
<< pdiffusion >>
rect 52 446 53 447 
<< pdiffusion >>
rect 53 446 54 447 
<< pdiffusion >>
rect 66 446 67 447 
<< pdiffusion >>
rect 67 446 68 447 
<< pdiffusion >>
rect 68 446 69 447 
<< pdiffusion >>
rect 69 446 70 447 
<< pdiffusion >>
rect 70 446 71 447 
<< pdiffusion >>
rect 71 446 72 447 
<< pdiffusion >>
rect 84 446 85 447 
<< pdiffusion >>
rect 85 446 86 447 
<< pdiffusion >>
rect 86 446 87 447 
<< pdiffusion >>
rect 87 446 88 447 
<< pdiffusion >>
rect 88 446 89 447 
<< pdiffusion >>
rect 89 446 90 447 
<< pdiffusion >>
rect 102 446 103 447 
<< pdiffusion >>
rect 103 446 104 447 
<< pdiffusion >>
rect 104 446 105 447 
<< pdiffusion >>
rect 105 446 106 447 
<< pdiffusion >>
rect 106 446 107 447 
<< pdiffusion >>
rect 107 446 108 447 
<< pdiffusion >>
rect 120 446 121 447 
<< pdiffusion >>
rect 121 446 122 447 
<< pdiffusion >>
rect 122 446 123 447 
<< pdiffusion >>
rect 123 446 124 447 
<< pdiffusion >>
rect 124 446 125 447 
<< pdiffusion >>
rect 125 446 126 447 
<< pdiffusion >>
rect 138 446 139 447 
<< pdiffusion >>
rect 139 446 140 447 
<< pdiffusion >>
rect 140 446 141 447 
<< pdiffusion >>
rect 141 446 142 447 
<< pdiffusion >>
rect 142 446 143 447 
<< pdiffusion >>
rect 143 446 144 447 
<< pdiffusion >>
rect 156 446 157 447 
<< pdiffusion >>
rect 157 446 158 447 
<< pdiffusion >>
rect 158 446 159 447 
<< pdiffusion >>
rect 159 446 160 447 
<< pdiffusion >>
rect 160 446 161 447 
<< pdiffusion >>
rect 161 446 162 447 
<< m1 >>
rect 172 446 173 447 
<< pdiffusion >>
rect 174 446 175 447 
<< pdiffusion >>
rect 175 446 176 447 
<< pdiffusion >>
rect 176 446 177 447 
<< pdiffusion >>
rect 177 446 178 447 
<< pdiffusion >>
rect 178 446 179 447 
<< pdiffusion >>
rect 179 446 180 447 
<< pdiffusion >>
rect 192 446 193 447 
<< pdiffusion >>
rect 193 446 194 447 
<< pdiffusion >>
rect 194 446 195 447 
<< pdiffusion >>
rect 195 446 196 447 
<< pdiffusion >>
rect 196 446 197 447 
<< pdiffusion >>
rect 197 446 198 447 
<< pdiffusion >>
rect 210 446 211 447 
<< pdiffusion >>
rect 211 446 212 447 
<< pdiffusion >>
rect 212 446 213 447 
<< pdiffusion >>
rect 213 446 214 447 
<< pdiffusion >>
rect 214 446 215 447 
<< pdiffusion >>
rect 215 446 216 447 
<< m1 >>
rect 226 446 227 447 
<< pdiffusion >>
rect 228 446 229 447 
<< pdiffusion >>
rect 229 446 230 447 
<< pdiffusion >>
rect 230 446 231 447 
<< pdiffusion >>
rect 231 446 232 447 
<< pdiffusion >>
rect 232 446 233 447 
<< pdiffusion >>
rect 233 446 234 447 
<< pdiffusion >>
rect 246 446 247 447 
<< pdiffusion >>
rect 247 446 248 447 
<< pdiffusion >>
rect 248 446 249 447 
<< pdiffusion >>
rect 249 446 250 447 
<< pdiffusion >>
rect 250 446 251 447 
<< pdiffusion >>
rect 251 446 252 447 
<< pdiffusion >>
rect 264 446 265 447 
<< pdiffusion >>
rect 265 446 266 447 
<< pdiffusion >>
rect 266 446 267 447 
<< pdiffusion >>
rect 267 446 268 447 
<< pdiffusion >>
rect 268 446 269 447 
<< pdiffusion >>
rect 269 446 270 447 
<< pdiffusion >>
rect 282 446 283 447 
<< pdiffusion >>
rect 283 446 284 447 
<< pdiffusion >>
rect 284 446 285 447 
<< pdiffusion >>
rect 285 446 286 447 
<< pdiffusion >>
rect 286 446 287 447 
<< pdiffusion >>
rect 287 446 288 447 
<< m1 >>
rect 289 446 290 447 
<< pdiffusion >>
rect 300 446 301 447 
<< pdiffusion >>
rect 301 446 302 447 
<< pdiffusion >>
rect 302 446 303 447 
<< pdiffusion >>
rect 303 446 304 447 
<< pdiffusion >>
rect 304 446 305 447 
<< pdiffusion >>
rect 305 446 306 447 
<< m1 >>
rect 307 446 308 447 
<< pdiffusion >>
rect 318 446 319 447 
<< pdiffusion >>
rect 319 446 320 447 
<< pdiffusion >>
rect 320 446 321 447 
<< pdiffusion >>
rect 321 446 322 447 
<< pdiffusion >>
rect 322 446 323 447 
<< pdiffusion >>
rect 323 446 324 447 
<< pdiffusion >>
rect 336 446 337 447 
<< pdiffusion >>
rect 337 446 338 447 
<< pdiffusion >>
rect 338 446 339 447 
<< pdiffusion >>
rect 339 446 340 447 
<< pdiffusion >>
rect 340 446 341 447 
<< pdiffusion >>
rect 341 446 342 447 
<< m1 >>
rect 343 446 344 447 
<< pdiffusion >>
rect 354 446 355 447 
<< pdiffusion >>
rect 355 446 356 447 
<< pdiffusion >>
rect 356 446 357 447 
<< pdiffusion >>
rect 357 446 358 447 
<< pdiffusion >>
rect 358 446 359 447 
<< pdiffusion >>
rect 359 446 360 447 
<< pdiffusion >>
rect 372 446 373 447 
<< pdiffusion >>
rect 373 446 374 447 
<< pdiffusion >>
rect 374 446 375 447 
<< pdiffusion >>
rect 375 446 376 447 
<< pdiffusion >>
rect 376 446 377 447 
<< pdiffusion >>
rect 377 446 378 447 
<< pdiffusion >>
rect 390 446 391 447 
<< pdiffusion >>
rect 391 446 392 447 
<< pdiffusion >>
rect 392 446 393 447 
<< pdiffusion >>
rect 393 446 394 447 
<< pdiffusion >>
rect 394 446 395 447 
<< pdiffusion >>
rect 395 446 396 447 
<< pdiffusion >>
rect 408 446 409 447 
<< pdiffusion >>
rect 409 446 410 447 
<< pdiffusion >>
rect 410 446 411 447 
<< pdiffusion >>
rect 411 446 412 447 
<< pdiffusion >>
rect 412 446 413 447 
<< pdiffusion >>
rect 413 446 414 447 
<< pdiffusion >>
rect 426 446 427 447 
<< pdiffusion >>
rect 427 446 428 447 
<< pdiffusion >>
rect 428 446 429 447 
<< pdiffusion >>
rect 429 446 430 447 
<< pdiffusion >>
rect 430 446 431 447 
<< pdiffusion >>
rect 431 446 432 447 
<< pdiffusion >>
rect 444 446 445 447 
<< pdiffusion >>
rect 445 446 446 447 
<< pdiffusion >>
rect 446 446 447 447 
<< pdiffusion >>
rect 447 446 448 447 
<< pdiffusion >>
rect 448 446 449 447 
<< pdiffusion >>
rect 449 446 450 447 
<< pdiffusion >>
rect 12 447 13 448 
<< pdiffusion >>
rect 13 447 14 448 
<< pdiffusion >>
rect 14 447 15 448 
<< pdiffusion >>
rect 15 447 16 448 
<< pdiffusion >>
rect 16 447 17 448 
<< pdiffusion >>
rect 17 447 18 448 
<< pdiffusion >>
rect 30 447 31 448 
<< pdiffusion >>
rect 31 447 32 448 
<< pdiffusion >>
rect 32 447 33 448 
<< pdiffusion >>
rect 33 447 34 448 
<< pdiffusion >>
rect 34 447 35 448 
<< pdiffusion >>
rect 35 447 36 448 
<< pdiffusion >>
rect 48 447 49 448 
<< pdiffusion >>
rect 49 447 50 448 
<< pdiffusion >>
rect 50 447 51 448 
<< pdiffusion >>
rect 51 447 52 448 
<< pdiffusion >>
rect 52 447 53 448 
<< pdiffusion >>
rect 53 447 54 448 
<< pdiffusion >>
rect 66 447 67 448 
<< pdiffusion >>
rect 67 447 68 448 
<< pdiffusion >>
rect 68 447 69 448 
<< pdiffusion >>
rect 69 447 70 448 
<< pdiffusion >>
rect 70 447 71 448 
<< pdiffusion >>
rect 71 447 72 448 
<< pdiffusion >>
rect 84 447 85 448 
<< pdiffusion >>
rect 85 447 86 448 
<< pdiffusion >>
rect 86 447 87 448 
<< pdiffusion >>
rect 87 447 88 448 
<< pdiffusion >>
rect 88 447 89 448 
<< pdiffusion >>
rect 89 447 90 448 
<< pdiffusion >>
rect 102 447 103 448 
<< pdiffusion >>
rect 103 447 104 448 
<< pdiffusion >>
rect 104 447 105 448 
<< pdiffusion >>
rect 105 447 106 448 
<< pdiffusion >>
rect 106 447 107 448 
<< pdiffusion >>
rect 107 447 108 448 
<< pdiffusion >>
rect 120 447 121 448 
<< pdiffusion >>
rect 121 447 122 448 
<< pdiffusion >>
rect 122 447 123 448 
<< pdiffusion >>
rect 123 447 124 448 
<< pdiffusion >>
rect 124 447 125 448 
<< pdiffusion >>
rect 125 447 126 448 
<< pdiffusion >>
rect 138 447 139 448 
<< pdiffusion >>
rect 139 447 140 448 
<< pdiffusion >>
rect 140 447 141 448 
<< pdiffusion >>
rect 141 447 142 448 
<< pdiffusion >>
rect 142 447 143 448 
<< pdiffusion >>
rect 143 447 144 448 
<< pdiffusion >>
rect 156 447 157 448 
<< pdiffusion >>
rect 157 447 158 448 
<< pdiffusion >>
rect 158 447 159 448 
<< pdiffusion >>
rect 159 447 160 448 
<< pdiffusion >>
rect 160 447 161 448 
<< pdiffusion >>
rect 161 447 162 448 
<< m1 >>
rect 172 447 173 448 
<< pdiffusion >>
rect 174 447 175 448 
<< pdiffusion >>
rect 175 447 176 448 
<< pdiffusion >>
rect 176 447 177 448 
<< pdiffusion >>
rect 177 447 178 448 
<< pdiffusion >>
rect 178 447 179 448 
<< pdiffusion >>
rect 179 447 180 448 
<< pdiffusion >>
rect 192 447 193 448 
<< pdiffusion >>
rect 193 447 194 448 
<< pdiffusion >>
rect 194 447 195 448 
<< pdiffusion >>
rect 195 447 196 448 
<< pdiffusion >>
rect 196 447 197 448 
<< pdiffusion >>
rect 197 447 198 448 
<< pdiffusion >>
rect 210 447 211 448 
<< pdiffusion >>
rect 211 447 212 448 
<< pdiffusion >>
rect 212 447 213 448 
<< pdiffusion >>
rect 213 447 214 448 
<< pdiffusion >>
rect 214 447 215 448 
<< pdiffusion >>
rect 215 447 216 448 
<< m1 >>
rect 226 447 227 448 
<< pdiffusion >>
rect 228 447 229 448 
<< pdiffusion >>
rect 229 447 230 448 
<< pdiffusion >>
rect 230 447 231 448 
<< pdiffusion >>
rect 231 447 232 448 
<< pdiffusion >>
rect 232 447 233 448 
<< pdiffusion >>
rect 233 447 234 448 
<< pdiffusion >>
rect 246 447 247 448 
<< pdiffusion >>
rect 247 447 248 448 
<< pdiffusion >>
rect 248 447 249 448 
<< pdiffusion >>
rect 249 447 250 448 
<< pdiffusion >>
rect 250 447 251 448 
<< pdiffusion >>
rect 251 447 252 448 
<< pdiffusion >>
rect 264 447 265 448 
<< pdiffusion >>
rect 265 447 266 448 
<< pdiffusion >>
rect 266 447 267 448 
<< pdiffusion >>
rect 267 447 268 448 
<< pdiffusion >>
rect 268 447 269 448 
<< pdiffusion >>
rect 269 447 270 448 
<< pdiffusion >>
rect 282 447 283 448 
<< pdiffusion >>
rect 283 447 284 448 
<< pdiffusion >>
rect 284 447 285 448 
<< pdiffusion >>
rect 285 447 286 448 
<< pdiffusion >>
rect 286 447 287 448 
<< pdiffusion >>
rect 287 447 288 448 
<< m1 >>
rect 289 447 290 448 
<< pdiffusion >>
rect 300 447 301 448 
<< pdiffusion >>
rect 301 447 302 448 
<< pdiffusion >>
rect 302 447 303 448 
<< pdiffusion >>
rect 303 447 304 448 
<< pdiffusion >>
rect 304 447 305 448 
<< pdiffusion >>
rect 305 447 306 448 
<< m1 >>
rect 307 447 308 448 
<< pdiffusion >>
rect 318 447 319 448 
<< pdiffusion >>
rect 319 447 320 448 
<< pdiffusion >>
rect 320 447 321 448 
<< pdiffusion >>
rect 321 447 322 448 
<< pdiffusion >>
rect 322 447 323 448 
<< pdiffusion >>
rect 323 447 324 448 
<< pdiffusion >>
rect 336 447 337 448 
<< pdiffusion >>
rect 337 447 338 448 
<< pdiffusion >>
rect 338 447 339 448 
<< pdiffusion >>
rect 339 447 340 448 
<< pdiffusion >>
rect 340 447 341 448 
<< pdiffusion >>
rect 341 447 342 448 
<< m1 >>
rect 343 447 344 448 
<< pdiffusion >>
rect 354 447 355 448 
<< pdiffusion >>
rect 355 447 356 448 
<< pdiffusion >>
rect 356 447 357 448 
<< pdiffusion >>
rect 357 447 358 448 
<< pdiffusion >>
rect 358 447 359 448 
<< pdiffusion >>
rect 359 447 360 448 
<< pdiffusion >>
rect 372 447 373 448 
<< pdiffusion >>
rect 373 447 374 448 
<< pdiffusion >>
rect 374 447 375 448 
<< pdiffusion >>
rect 375 447 376 448 
<< pdiffusion >>
rect 376 447 377 448 
<< pdiffusion >>
rect 377 447 378 448 
<< pdiffusion >>
rect 390 447 391 448 
<< pdiffusion >>
rect 391 447 392 448 
<< pdiffusion >>
rect 392 447 393 448 
<< pdiffusion >>
rect 393 447 394 448 
<< pdiffusion >>
rect 394 447 395 448 
<< pdiffusion >>
rect 395 447 396 448 
<< pdiffusion >>
rect 408 447 409 448 
<< pdiffusion >>
rect 409 447 410 448 
<< pdiffusion >>
rect 410 447 411 448 
<< pdiffusion >>
rect 411 447 412 448 
<< pdiffusion >>
rect 412 447 413 448 
<< pdiffusion >>
rect 413 447 414 448 
<< pdiffusion >>
rect 426 447 427 448 
<< pdiffusion >>
rect 427 447 428 448 
<< pdiffusion >>
rect 428 447 429 448 
<< pdiffusion >>
rect 429 447 430 448 
<< pdiffusion >>
rect 430 447 431 448 
<< pdiffusion >>
rect 431 447 432 448 
<< pdiffusion >>
rect 444 447 445 448 
<< pdiffusion >>
rect 445 447 446 448 
<< pdiffusion >>
rect 446 447 447 448 
<< pdiffusion >>
rect 447 447 448 448 
<< pdiffusion >>
rect 448 447 449 448 
<< pdiffusion >>
rect 449 447 450 448 
<< pdiffusion >>
rect 12 448 13 449 
<< pdiffusion >>
rect 13 448 14 449 
<< pdiffusion >>
rect 14 448 15 449 
<< pdiffusion >>
rect 15 448 16 449 
<< pdiffusion >>
rect 16 448 17 449 
<< pdiffusion >>
rect 17 448 18 449 
<< pdiffusion >>
rect 30 448 31 449 
<< pdiffusion >>
rect 31 448 32 449 
<< pdiffusion >>
rect 32 448 33 449 
<< pdiffusion >>
rect 33 448 34 449 
<< pdiffusion >>
rect 34 448 35 449 
<< pdiffusion >>
rect 35 448 36 449 
<< pdiffusion >>
rect 48 448 49 449 
<< pdiffusion >>
rect 49 448 50 449 
<< pdiffusion >>
rect 50 448 51 449 
<< pdiffusion >>
rect 51 448 52 449 
<< pdiffusion >>
rect 52 448 53 449 
<< pdiffusion >>
rect 53 448 54 449 
<< pdiffusion >>
rect 66 448 67 449 
<< pdiffusion >>
rect 67 448 68 449 
<< pdiffusion >>
rect 68 448 69 449 
<< pdiffusion >>
rect 69 448 70 449 
<< pdiffusion >>
rect 70 448 71 449 
<< pdiffusion >>
rect 71 448 72 449 
<< pdiffusion >>
rect 84 448 85 449 
<< pdiffusion >>
rect 85 448 86 449 
<< pdiffusion >>
rect 86 448 87 449 
<< pdiffusion >>
rect 87 448 88 449 
<< pdiffusion >>
rect 88 448 89 449 
<< pdiffusion >>
rect 89 448 90 449 
<< pdiffusion >>
rect 102 448 103 449 
<< pdiffusion >>
rect 103 448 104 449 
<< pdiffusion >>
rect 104 448 105 449 
<< pdiffusion >>
rect 105 448 106 449 
<< pdiffusion >>
rect 106 448 107 449 
<< pdiffusion >>
rect 107 448 108 449 
<< pdiffusion >>
rect 120 448 121 449 
<< pdiffusion >>
rect 121 448 122 449 
<< pdiffusion >>
rect 122 448 123 449 
<< pdiffusion >>
rect 123 448 124 449 
<< pdiffusion >>
rect 124 448 125 449 
<< pdiffusion >>
rect 125 448 126 449 
<< pdiffusion >>
rect 138 448 139 449 
<< pdiffusion >>
rect 139 448 140 449 
<< pdiffusion >>
rect 140 448 141 449 
<< pdiffusion >>
rect 141 448 142 449 
<< pdiffusion >>
rect 142 448 143 449 
<< pdiffusion >>
rect 143 448 144 449 
<< pdiffusion >>
rect 156 448 157 449 
<< pdiffusion >>
rect 157 448 158 449 
<< pdiffusion >>
rect 158 448 159 449 
<< pdiffusion >>
rect 159 448 160 449 
<< pdiffusion >>
rect 160 448 161 449 
<< pdiffusion >>
rect 161 448 162 449 
<< m1 >>
rect 172 448 173 449 
<< pdiffusion >>
rect 174 448 175 449 
<< pdiffusion >>
rect 175 448 176 449 
<< pdiffusion >>
rect 176 448 177 449 
<< pdiffusion >>
rect 177 448 178 449 
<< pdiffusion >>
rect 178 448 179 449 
<< pdiffusion >>
rect 179 448 180 449 
<< pdiffusion >>
rect 192 448 193 449 
<< pdiffusion >>
rect 193 448 194 449 
<< pdiffusion >>
rect 194 448 195 449 
<< pdiffusion >>
rect 195 448 196 449 
<< pdiffusion >>
rect 196 448 197 449 
<< pdiffusion >>
rect 197 448 198 449 
<< pdiffusion >>
rect 210 448 211 449 
<< pdiffusion >>
rect 211 448 212 449 
<< pdiffusion >>
rect 212 448 213 449 
<< pdiffusion >>
rect 213 448 214 449 
<< pdiffusion >>
rect 214 448 215 449 
<< pdiffusion >>
rect 215 448 216 449 
<< m1 >>
rect 226 448 227 449 
<< pdiffusion >>
rect 228 448 229 449 
<< pdiffusion >>
rect 229 448 230 449 
<< pdiffusion >>
rect 230 448 231 449 
<< pdiffusion >>
rect 231 448 232 449 
<< pdiffusion >>
rect 232 448 233 449 
<< pdiffusion >>
rect 233 448 234 449 
<< pdiffusion >>
rect 246 448 247 449 
<< pdiffusion >>
rect 247 448 248 449 
<< pdiffusion >>
rect 248 448 249 449 
<< pdiffusion >>
rect 249 448 250 449 
<< pdiffusion >>
rect 250 448 251 449 
<< pdiffusion >>
rect 251 448 252 449 
<< pdiffusion >>
rect 264 448 265 449 
<< pdiffusion >>
rect 265 448 266 449 
<< pdiffusion >>
rect 266 448 267 449 
<< pdiffusion >>
rect 267 448 268 449 
<< pdiffusion >>
rect 268 448 269 449 
<< pdiffusion >>
rect 269 448 270 449 
<< pdiffusion >>
rect 282 448 283 449 
<< pdiffusion >>
rect 283 448 284 449 
<< pdiffusion >>
rect 284 448 285 449 
<< pdiffusion >>
rect 285 448 286 449 
<< pdiffusion >>
rect 286 448 287 449 
<< pdiffusion >>
rect 287 448 288 449 
<< m1 >>
rect 289 448 290 449 
<< pdiffusion >>
rect 300 448 301 449 
<< pdiffusion >>
rect 301 448 302 449 
<< pdiffusion >>
rect 302 448 303 449 
<< pdiffusion >>
rect 303 448 304 449 
<< pdiffusion >>
rect 304 448 305 449 
<< pdiffusion >>
rect 305 448 306 449 
<< m1 >>
rect 307 448 308 449 
<< pdiffusion >>
rect 318 448 319 449 
<< pdiffusion >>
rect 319 448 320 449 
<< pdiffusion >>
rect 320 448 321 449 
<< pdiffusion >>
rect 321 448 322 449 
<< pdiffusion >>
rect 322 448 323 449 
<< pdiffusion >>
rect 323 448 324 449 
<< pdiffusion >>
rect 336 448 337 449 
<< pdiffusion >>
rect 337 448 338 449 
<< pdiffusion >>
rect 338 448 339 449 
<< pdiffusion >>
rect 339 448 340 449 
<< pdiffusion >>
rect 340 448 341 449 
<< pdiffusion >>
rect 341 448 342 449 
<< m1 >>
rect 343 448 344 449 
<< pdiffusion >>
rect 354 448 355 449 
<< pdiffusion >>
rect 355 448 356 449 
<< pdiffusion >>
rect 356 448 357 449 
<< pdiffusion >>
rect 357 448 358 449 
<< pdiffusion >>
rect 358 448 359 449 
<< pdiffusion >>
rect 359 448 360 449 
<< pdiffusion >>
rect 372 448 373 449 
<< pdiffusion >>
rect 373 448 374 449 
<< pdiffusion >>
rect 374 448 375 449 
<< pdiffusion >>
rect 375 448 376 449 
<< pdiffusion >>
rect 376 448 377 449 
<< pdiffusion >>
rect 377 448 378 449 
<< pdiffusion >>
rect 390 448 391 449 
<< pdiffusion >>
rect 391 448 392 449 
<< pdiffusion >>
rect 392 448 393 449 
<< pdiffusion >>
rect 393 448 394 449 
<< pdiffusion >>
rect 394 448 395 449 
<< pdiffusion >>
rect 395 448 396 449 
<< pdiffusion >>
rect 408 448 409 449 
<< pdiffusion >>
rect 409 448 410 449 
<< pdiffusion >>
rect 410 448 411 449 
<< pdiffusion >>
rect 411 448 412 449 
<< pdiffusion >>
rect 412 448 413 449 
<< pdiffusion >>
rect 413 448 414 449 
<< pdiffusion >>
rect 426 448 427 449 
<< pdiffusion >>
rect 427 448 428 449 
<< pdiffusion >>
rect 428 448 429 449 
<< pdiffusion >>
rect 429 448 430 449 
<< pdiffusion >>
rect 430 448 431 449 
<< pdiffusion >>
rect 431 448 432 449 
<< pdiffusion >>
rect 444 448 445 449 
<< pdiffusion >>
rect 445 448 446 449 
<< pdiffusion >>
rect 446 448 447 449 
<< pdiffusion >>
rect 447 448 448 449 
<< pdiffusion >>
rect 448 448 449 449 
<< pdiffusion >>
rect 449 448 450 449 
<< pdiffusion >>
rect 12 449 13 450 
<< pdiffusion >>
rect 13 449 14 450 
<< pdiffusion >>
rect 14 449 15 450 
<< pdiffusion >>
rect 15 449 16 450 
<< pdiffusion >>
rect 16 449 17 450 
<< pdiffusion >>
rect 17 449 18 450 
<< pdiffusion >>
rect 30 449 31 450 
<< pdiffusion >>
rect 31 449 32 450 
<< pdiffusion >>
rect 32 449 33 450 
<< pdiffusion >>
rect 33 449 34 450 
<< pdiffusion >>
rect 34 449 35 450 
<< pdiffusion >>
rect 35 449 36 450 
<< pdiffusion >>
rect 48 449 49 450 
<< pdiffusion >>
rect 49 449 50 450 
<< pdiffusion >>
rect 50 449 51 450 
<< pdiffusion >>
rect 51 449 52 450 
<< pdiffusion >>
rect 52 449 53 450 
<< pdiffusion >>
rect 53 449 54 450 
<< pdiffusion >>
rect 66 449 67 450 
<< m1 >>
rect 67 449 68 450 
<< pdiffusion >>
rect 67 449 68 450 
<< pdiffusion >>
rect 68 449 69 450 
<< pdiffusion >>
rect 69 449 70 450 
<< pdiffusion >>
rect 70 449 71 450 
<< pdiffusion >>
rect 71 449 72 450 
<< pdiffusion >>
rect 84 449 85 450 
<< pdiffusion >>
rect 85 449 86 450 
<< pdiffusion >>
rect 86 449 87 450 
<< pdiffusion >>
rect 87 449 88 450 
<< m1 >>
rect 88 449 89 450 
<< pdiffusion >>
rect 88 449 89 450 
<< pdiffusion >>
rect 89 449 90 450 
<< pdiffusion >>
rect 102 449 103 450 
<< pdiffusion >>
rect 103 449 104 450 
<< pdiffusion >>
rect 104 449 105 450 
<< pdiffusion >>
rect 105 449 106 450 
<< pdiffusion >>
rect 106 449 107 450 
<< pdiffusion >>
rect 107 449 108 450 
<< pdiffusion >>
rect 120 449 121 450 
<< pdiffusion >>
rect 121 449 122 450 
<< pdiffusion >>
rect 122 449 123 450 
<< pdiffusion >>
rect 123 449 124 450 
<< pdiffusion >>
rect 124 449 125 450 
<< pdiffusion >>
rect 125 449 126 450 
<< pdiffusion >>
rect 138 449 139 450 
<< pdiffusion >>
rect 139 449 140 450 
<< pdiffusion >>
rect 140 449 141 450 
<< pdiffusion >>
rect 141 449 142 450 
<< pdiffusion >>
rect 142 449 143 450 
<< pdiffusion >>
rect 143 449 144 450 
<< pdiffusion >>
rect 156 449 157 450 
<< pdiffusion >>
rect 157 449 158 450 
<< pdiffusion >>
rect 158 449 159 450 
<< pdiffusion >>
rect 159 449 160 450 
<< pdiffusion >>
rect 160 449 161 450 
<< pdiffusion >>
rect 161 449 162 450 
<< m1 >>
rect 172 449 173 450 
<< pdiffusion >>
rect 174 449 175 450 
<< m1 >>
rect 175 449 176 450 
<< pdiffusion >>
rect 175 449 176 450 
<< pdiffusion >>
rect 176 449 177 450 
<< pdiffusion >>
rect 177 449 178 450 
<< pdiffusion >>
rect 178 449 179 450 
<< pdiffusion >>
rect 179 449 180 450 
<< pdiffusion >>
rect 192 449 193 450 
<< pdiffusion >>
rect 193 449 194 450 
<< pdiffusion >>
rect 194 449 195 450 
<< pdiffusion >>
rect 195 449 196 450 
<< pdiffusion >>
rect 196 449 197 450 
<< pdiffusion >>
rect 197 449 198 450 
<< pdiffusion >>
rect 210 449 211 450 
<< m1 >>
rect 211 449 212 450 
<< pdiffusion >>
rect 211 449 212 450 
<< pdiffusion >>
rect 212 449 213 450 
<< pdiffusion >>
rect 213 449 214 450 
<< pdiffusion >>
rect 214 449 215 450 
<< pdiffusion >>
rect 215 449 216 450 
<< m1 >>
rect 226 449 227 450 
<< pdiffusion >>
rect 228 449 229 450 
<< pdiffusion >>
rect 229 449 230 450 
<< pdiffusion >>
rect 230 449 231 450 
<< pdiffusion >>
rect 231 449 232 450 
<< pdiffusion >>
rect 232 449 233 450 
<< pdiffusion >>
rect 233 449 234 450 
<< pdiffusion >>
rect 246 449 247 450 
<< pdiffusion >>
rect 247 449 248 450 
<< pdiffusion >>
rect 248 449 249 450 
<< pdiffusion >>
rect 249 449 250 450 
<< pdiffusion >>
rect 250 449 251 450 
<< pdiffusion >>
rect 251 449 252 450 
<< pdiffusion >>
rect 264 449 265 450 
<< pdiffusion >>
rect 265 449 266 450 
<< pdiffusion >>
rect 266 449 267 450 
<< pdiffusion >>
rect 267 449 268 450 
<< pdiffusion >>
rect 268 449 269 450 
<< pdiffusion >>
rect 269 449 270 450 
<< pdiffusion >>
rect 282 449 283 450 
<< pdiffusion >>
rect 283 449 284 450 
<< pdiffusion >>
rect 284 449 285 450 
<< pdiffusion >>
rect 285 449 286 450 
<< pdiffusion >>
rect 286 449 287 450 
<< pdiffusion >>
rect 287 449 288 450 
<< m1 >>
rect 289 449 290 450 
<< pdiffusion >>
rect 300 449 301 450 
<< pdiffusion >>
rect 301 449 302 450 
<< pdiffusion >>
rect 302 449 303 450 
<< pdiffusion >>
rect 303 449 304 450 
<< pdiffusion >>
rect 304 449 305 450 
<< pdiffusion >>
rect 305 449 306 450 
<< m1 >>
rect 307 449 308 450 
<< pdiffusion >>
rect 318 449 319 450 
<< pdiffusion >>
rect 319 449 320 450 
<< pdiffusion >>
rect 320 449 321 450 
<< pdiffusion >>
rect 321 449 322 450 
<< m1 >>
rect 322 449 323 450 
<< pdiffusion >>
rect 322 449 323 450 
<< pdiffusion >>
rect 323 449 324 450 
<< pdiffusion >>
rect 336 449 337 450 
<< pdiffusion >>
rect 337 449 338 450 
<< pdiffusion >>
rect 338 449 339 450 
<< pdiffusion >>
rect 339 449 340 450 
<< pdiffusion >>
rect 340 449 341 450 
<< pdiffusion >>
rect 341 449 342 450 
<< m1 >>
rect 343 449 344 450 
<< pdiffusion >>
rect 354 449 355 450 
<< pdiffusion >>
rect 355 449 356 450 
<< pdiffusion >>
rect 356 449 357 450 
<< pdiffusion >>
rect 357 449 358 450 
<< m1 >>
rect 358 449 359 450 
<< pdiffusion >>
rect 358 449 359 450 
<< pdiffusion >>
rect 359 449 360 450 
<< pdiffusion >>
rect 372 449 373 450 
<< pdiffusion >>
rect 373 449 374 450 
<< pdiffusion >>
rect 374 449 375 450 
<< pdiffusion >>
rect 375 449 376 450 
<< pdiffusion >>
rect 376 449 377 450 
<< pdiffusion >>
rect 377 449 378 450 
<< pdiffusion >>
rect 390 449 391 450 
<< pdiffusion >>
rect 391 449 392 450 
<< pdiffusion >>
rect 392 449 393 450 
<< pdiffusion >>
rect 393 449 394 450 
<< pdiffusion >>
rect 394 449 395 450 
<< pdiffusion >>
rect 395 449 396 450 
<< pdiffusion >>
rect 408 449 409 450 
<< pdiffusion >>
rect 409 449 410 450 
<< pdiffusion >>
rect 410 449 411 450 
<< pdiffusion >>
rect 411 449 412 450 
<< pdiffusion >>
rect 412 449 413 450 
<< pdiffusion >>
rect 413 449 414 450 
<< pdiffusion >>
rect 426 449 427 450 
<< pdiffusion >>
rect 427 449 428 450 
<< pdiffusion >>
rect 428 449 429 450 
<< pdiffusion >>
rect 429 449 430 450 
<< pdiffusion >>
rect 430 449 431 450 
<< pdiffusion >>
rect 431 449 432 450 
<< pdiffusion >>
rect 444 449 445 450 
<< pdiffusion >>
rect 445 449 446 450 
<< pdiffusion >>
rect 446 449 447 450 
<< pdiffusion >>
rect 447 449 448 450 
<< m1 >>
rect 448 449 449 450 
<< pdiffusion >>
rect 448 449 449 450 
<< pdiffusion >>
rect 449 449 450 450 
<< m1 >>
rect 67 450 68 451 
<< m1 >>
rect 88 450 89 451 
<< m1 >>
rect 172 450 173 451 
<< m1 >>
rect 175 450 176 451 
<< m1 >>
rect 211 450 212 451 
<< m1 >>
rect 226 450 227 451 
<< m1 >>
rect 289 450 290 451 
<< m1 >>
rect 307 450 308 451 
<< m1 >>
rect 322 450 323 451 
<< m1 >>
rect 343 450 344 451 
<< m1 >>
rect 358 450 359 451 
<< m1 >>
rect 448 450 449 451 
<< m1 >>
rect 67 451 68 452 
<< m1 >>
rect 88 451 89 452 
<< m1 >>
rect 172 451 173 452 
<< m1 >>
rect 173 451 174 452 
<< m1 >>
rect 174 451 175 452 
<< m1 >>
rect 175 451 176 452 
<< m1 >>
rect 211 451 212 452 
<< m1 >>
rect 226 451 227 452 
<< m1 >>
rect 289 451 290 452 
<< m1 >>
rect 307 451 308 452 
<< m1 >>
rect 322 451 323 452 
<< m1 >>
rect 343 451 344 452 
<< m1 >>
rect 358 451 359 452 
<< m1 >>
rect 448 451 449 452 
<< m1 >>
rect 67 452 68 453 
<< m1 >>
rect 88 452 89 453 
<< m1 >>
rect 211 452 212 453 
<< m1 >>
rect 212 452 213 453 
<< m1 >>
rect 213 452 214 453 
<< m1 >>
rect 214 452 215 453 
<< m1 >>
rect 215 452 216 453 
<< m1 >>
rect 216 452 217 453 
<< m1 >>
rect 217 452 218 453 
<< m1 >>
rect 218 452 219 453 
<< m1 >>
rect 219 452 220 453 
<< m1 >>
rect 220 452 221 453 
<< m1 >>
rect 221 452 222 453 
<< m1 >>
rect 222 452 223 453 
<< m1 >>
rect 223 452 224 453 
<< m1 >>
rect 224 452 225 453 
<< m1 >>
rect 225 452 226 453 
<< m1 >>
rect 226 452 227 453 
<< m1 >>
rect 289 452 290 453 
<< m1 >>
rect 307 452 308 453 
<< m2 >>
rect 307 452 308 453 
<< m2c >>
rect 307 452 308 453 
<< m1 >>
rect 307 452 308 453 
<< m2 >>
rect 307 452 308 453 
<< m1 >>
rect 320 452 321 453 
<< m2 >>
rect 320 452 321 453 
<< m2c >>
rect 320 452 321 453 
<< m1 >>
rect 320 452 321 453 
<< m2 >>
rect 320 452 321 453 
<< m1 >>
rect 321 452 322 453 
<< m1 >>
rect 322 452 323 453 
<< m1 >>
rect 343 452 344 453 
<< m1 >>
rect 358 452 359 453 
<< m1 >>
rect 448 452 449 453 
<< m1 >>
rect 67 453 68 454 
<< m1 >>
rect 88 453 89 454 
<< m1 >>
rect 289 453 290 454 
<< m2 >>
rect 307 453 308 454 
<< m2 >>
rect 320 453 321 454 
<< m1 >>
rect 343 453 344 454 
<< m1 >>
rect 358 453 359 454 
<< m1 >>
rect 448 453 449 454 
<< m1 >>
rect 67 454 68 455 
<< m1 >>
rect 68 454 69 455 
<< m1 >>
rect 69 454 70 455 
<< m1 >>
rect 70 454 71 455 
<< m1 >>
rect 71 454 72 455 
<< m1 >>
rect 72 454 73 455 
<< m1 >>
rect 73 454 74 455 
<< m1 >>
rect 74 454 75 455 
<< m1 >>
rect 75 454 76 455 
<< m1 >>
rect 76 454 77 455 
<< m1 >>
rect 77 454 78 455 
<< m1 >>
rect 78 454 79 455 
<< m1 >>
rect 79 454 80 455 
<< m1 >>
rect 80 454 81 455 
<< m1 >>
rect 81 454 82 455 
<< m1 >>
rect 82 454 83 455 
<< m1 >>
rect 83 454 84 455 
<< m1 >>
rect 84 454 85 455 
<< m1 >>
rect 85 454 86 455 
<< m1 >>
rect 86 454 87 455 
<< m1 >>
rect 87 454 88 455 
<< m1 >>
rect 88 454 89 455 
<< m1 >>
rect 289 454 290 455 
<< m1 >>
rect 290 454 291 455 
<< m1 >>
rect 291 454 292 455 
<< m1 >>
rect 292 454 293 455 
<< m1 >>
rect 293 454 294 455 
<< m1 >>
rect 294 454 295 455 
<< m1 >>
rect 295 454 296 455 
<< m1 >>
rect 296 454 297 455 
<< m1 >>
rect 297 454 298 455 
<< m1 >>
rect 298 454 299 455 
<< m1 >>
rect 299 454 300 455 
<< m1 >>
rect 300 454 301 455 
<< m1 >>
rect 301 454 302 455 
<< m1 >>
rect 302 454 303 455 
<< m1 >>
rect 303 454 304 455 
<< m1 >>
rect 304 454 305 455 
<< m1 >>
rect 305 454 306 455 
<< m1 >>
rect 306 454 307 455 
<< m1 >>
rect 307 454 308 455 
<< m2 >>
rect 307 454 308 455 
<< m1 >>
rect 308 454 309 455 
<< m2 >>
rect 308 454 309 455 
<< m1 >>
rect 309 454 310 455 
<< m2 >>
rect 309 454 310 455 
<< m1 >>
rect 310 454 311 455 
<< m2 >>
rect 310 454 311 455 
<< m1 >>
rect 311 454 312 455 
<< m2 >>
rect 311 454 312 455 
<< m1 >>
rect 312 454 313 455 
<< m2 >>
rect 312 454 313 455 
<< m1 >>
rect 313 454 314 455 
<< m2 >>
rect 313 454 314 455 
<< m1 >>
rect 314 454 315 455 
<< m2 >>
rect 314 454 315 455 
<< m1 >>
rect 315 454 316 455 
<< m2 >>
rect 315 454 316 455 
<< m1 >>
rect 316 454 317 455 
<< m2 >>
rect 316 454 317 455 
<< m1 >>
rect 317 454 318 455 
<< m2 >>
rect 317 454 318 455 
<< m1 >>
rect 318 454 319 455 
<< m2 >>
rect 318 454 319 455 
<< m1 >>
rect 319 454 320 455 
<< m2 >>
rect 319 454 320 455 
<< m1 >>
rect 320 454 321 455 
<< m2 >>
rect 320 454 321 455 
<< m1 >>
rect 321 454 322 455 
<< m1 >>
rect 322 454 323 455 
<< m1 >>
rect 323 454 324 455 
<< m1 >>
rect 324 454 325 455 
<< m1 >>
rect 325 454 326 455 
<< m1 >>
rect 326 454 327 455 
<< m1 >>
rect 327 454 328 455 
<< m1 >>
rect 328 454 329 455 
<< m1 >>
rect 329 454 330 455 
<< m1 >>
rect 330 454 331 455 
<< m1 >>
rect 331 454 332 455 
<< m1 >>
rect 332 454 333 455 
<< m1 >>
rect 333 454 334 455 
<< m1 >>
rect 334 454 335 455 
<< m1 >>
rect 335 454 336 455 
<< m1 >>
rect 336 454 337 455 
<< m1 >>
rect 337 454 338 455 
<< m1 >>
rect 338 454 339 455 
<< m1 >>
rect 339 454 340 455 
<< m1 >>
rect 340 454 341 455 
<< m1 >>
rect 341 454 342 455 
<< m2 >>
rect 341 454 342 455 
<< m2c >>
rect 341 454 342 455 
<< m1 >>
rect 341 454 342 455 
<< m2 >>
rect 341 454 342 455 
<< m2 >>
rect 342 454 343 455 
<< m1 >>
rect 343 454 344 455 
<< m2 >>
rect 343 454 344 455 
<< m1 >>
rect 344 454 345 455 
<< m2 >>
rect 344 454 345 455 
<< m1 >>
rect 345 454 346 455 
<< m2 >>
rect 345 454 346 455 
<< m1 >>
rect 346 454 347 455 
<< m2 >>
rect 346 454 347 455 
<< m1 >>
rect 347 454 348 455 
<< m2 >>
rect 347 454 348 455 
<< m1 >>
rect 348 454 349 455 
<< m2 >>
rect 348 454 349 455 
<< m1 >>
rect 349 454 350 455 
<< m2 >>
rect 349 454 350 455 
<< m1 >>
rect 350 454 351 455 
<< m2 >>
rect 350 454 351 455 
<< m1 >>
rect 351 454 352 455 
<< m2 >>
rect 351 454 352 455 
<< m1 >>
rect 352 454 353 455 
<< m2 >>
rect 352 454 353 455 
<< m1 >>
rect 353 454 354 455 
<< m2 >>
rect 353 454 354 455 
<< m1 >>
rect 354 454 355 455 
<< m2 >>
rect 354 454 355 455 
<< m1 >>
rect 355 454 356 455 
<< m2 >>
rect 355 454 356 455 
<< m1 >>
rect 356 454 357 455 
<< m2 >>
rect 356 454 357 455 
<< m1 >>
rect 357 454 358 455 
<< m2 >>
rect 357 454 358 455 
<< m1 >>
rect 358 454 359 455 
<< m2 >>
rect 358 454 359 455 
<< m2 >>
rect 359 454 360 455 
<< m1 >>
rect 360 454 361 455 
<< m2 >>
rect 360 454 361 455 
<< m2c >>
rect 360 454 361 455 
<< m1 >>
rect 360 454 361 455 
<< m2 >>
rect 360 454 361 455 
<< m1 >>
rect 361 454 362 455 
<< m1 >>
rect 362 454 363 455 
<< m1 >>
rect 363 454 364 455 
<< m1 >>
rect 364 454 365 455 
<< m1 >>
rect 365 454 366 455 
<< m1 >>
rect 366 454 367 455 
<< m1 >>
rect 367 454 368 455 
<< m1 >>
rect 368 454 369 455 
<< m1 >>
rect 369 454 370 455 
<< m1 >>
rect 370 454 371 455 
<< m1 >>
rect 371 454 372 455 
<< m1 >>
rect 372 454 373 455 
<< m1 >>
rect 373 454 374 455 
<< m1 >>
rect 374 454 375 455 
<< m1 >>
rect 375 454 376 455 
<< m1 >>
rect 376 454 377 455 
<< m1 >>
rect 377 454 378 455 
<< m1 >>
rect 378 454 379 455 
<< m1 >>
rect 379 454 380 455 
<< m1 >>
rect 380 454 381 455 
<< m1 >>
rect 381 454 382 455 
<< m1 >>
rect 382 454 383 455 
<< m1 >>
rect 383 454 384 455 
<< m1 >>
rect 384 454 385 455 
<< m1 >>
rect 385 454 386 455 
<< m1 >>
rect 386 454 387 455 
<< m1 >>
rect 387 454 388 455 
<< m1 >>
rect 388 454 389 455 
<< m1 >>
rect 389 454 390 455 
<< m1 >>
rect 390 454 391 455 
<< m1 >>
rect 391 454 392 455 
<< m1 >>
rect 392 454 393 455 
<< m1 >>
rect 393 454 394 455 
<< m1 >>
rect 394 454 395 455 
<< m1 >>
rect 395 454 396 455 
<< m1 >>
rect 396 454 397 455 
<< m1 >>
rect 397 454 398 455 
<< m1 >>
rect 398 454 399 455 
<< m1 >>
rect 399 454 400 455 
<< m1 >>
rect 400 454 401 455 
<< m1 >>
rect 401 454 402 455 
<< m1 >>
rect 402 454 403 455 
<< m1 >>
rect 403 454 404 455 
<< m1 >>
rect 404 454 405 455 
<< m1 >>
rect 405 454 406 455 
<< m1 >>
rect 406 454 407 455 
<< m1 >>
rect 407 454 408 455 
<< m1 >>
rect 408 454 409 455 
<< m1 >>
rect 409 454 410 455 
<< m1 >>
rect 410 454 411 455 
<< m1 >>
rect 411 454 412 455 
<< m1 >>
rect 412 454 413 455 
<< m1 >>
rect 413 454 414 455 
<< m1 >>
rect 414 454 415 455 
<< m1 >>
rect 415 454 416 455 
<< m1 >>
rect 416 454 417 455 
<< m1 >>
rect 417 454 418 455 
<< m1 >>
rect 418 454 419 455 
<< m1 >>
rect 419 454 420 455 
<< m1 >>
rect 420 454 421 455 
<< m1 >>
rect 421 454 422 455 
<< m1 >>
rect 422 454 423 455 
<< m1 >>
rect 423 454 424 455 
<< m1 >>
rect 424 454 425 455 
<< m1 >>
rect 425 454 426 455 
<< m1 >>
rect 426 454 427 455 
<< m1 >>
rect 427 454 428 455 
<< m1 >>
rect 428 454 429 455 
<< m1 >>
rect 429 454 430 455 
<< m1 >>
rect 430 454 431 455 
<< m1 >>
rect 431 454 432 455 
<< m1 >>
rect 432 454 433 455 
<< m1 >>
rect 433 454 434 455 
<< m1 >>
rect 434 454 435 455 
<< m1 >>
rect 435 454 436 455 
<< m1 >>
rect 436 454 437 455 
<< m1 >>
rect 437 454 438 455 
<< m1 >>
rect 438 454 439 455 
<< m1 >>
rect 439 454 440 455 
<< m1 >>
rect 440 454 441 455 
<< m1 >>
rect 441 454 442 455 
<< m1 >>
rect 442 454 443 455 
<< m1 >>
rect 443 454 444 455 
<< m1 >>
rect 444 454 445 455 
<< m1 >>
rect 445 454 446 455 
<< m1 >>
rect 446 454 447 455 
<< m1 >>
rect 447 454 448 455 
<< m1 >>
rect 448 454 449 455 
<< labels >>
rlabel pdiffusion 283 102 284 103  0 t = 1
rlabel pdiffusion 286 102 287 103  0 t = 2
rlabel pdiffusion 283 107 284 108  0 t = 3
rlabel pdiffusion 286 107 287 108  0 t = 4
rlabel pdiffusion 282 102 288 108 0 cell no = 1
<< m1 >>
rect 283 102 284 103 
rect 286 102 287 103 
rect 283 107 284 108 
rect 286 107 287 108 
<< m2 >>
rect 283 102 284 103 
rect 286 102 287 103 
rect 283 107 284 108 
rect 286 107 287 108 
<< m2c >>
rect 283 102 284 103 
rect 286 102 287 103 
rect 283 107 284 108 
rect 286 107 287 108 
<< labels >>
rlabel pdiffusion 67 30 68 31  0 t = 1
rlabel pdiffusion 70 30 71 31  0 t = 2
rlabel pdiffusion 67 35 68 36  0 t = 3
rlabel pdiffusion 70 35 71 36  0 t = 4
rlabel pdiffusion 66 30 72 36 0 cell no = 2
<< m1 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2c >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< labels >>
rlabel pdiffusion 319 12 320 13  0 t = 1
rlabel pdiffusion 322 12 323 13  0 t = 2
rlabel pdiffusion 319 17 320 18  0 t = 3
rlabel pdiffusion 322 17 323 18  0 t = 4
rlabel pdiffusion 318 12 324 18 0 cell no = 3
<< m1 >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< m2 >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< m2c >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< labels >>
rlabel pdiffusion 49 246 50 247  0 t = 1
rlabel pdiffusion 52 246 53 247  0 t = 2
rlabel pdiffusion 49 251 50 252  0 t = 3
rlabel pdiffusion 52 251 53 252  0 t = 4
rlabel pdiffusion 48 246 54 252 0 cell no = 4
<< m1 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2c >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 5
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 6
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 175 138 176 139  0 t = 1
rlabel pdiffusion 178 138 179 139  0 t = 2
rlabel pdiffusion 175 143 176 144  0 t = 3
rlabel pdiffusion 178 143 179 144  0 t = 4
rlabel pdiffusion 174 138 180 144 0 cell no = 7
<< m1 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2c >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< labels >>
rlabel pdiffusion 193 174 194 175  0 t = 1
rlabel pdiffusion 196 174 197 175  0 t = 2
rlabel pdiffusion 193 179 194 180  0 t = 3
rlabel pdiffusion 196 179 197 180  0 t = 4
rlabel pdiffusion 192 174 198 180 0 cell no = 8
<< m1 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2c >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< labels >>
rlabel pdiffusion 157 12 158 13  0 t = 1
rlabel pdiffusion 160 12 161 13  0 t = 2
rlabel pdiffusion 157 17 158 18  0 t = 3
rlabel pdiffusion 160 17 161 18  0 t = 4
rlabel pdiffusion 156 12 162 18 0 cell no = 9
<< m1 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2c >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< labels >>
rlabel pdiffusion 157 30 158 31  0 t = 1
rlabel pdiffusion 160 30 161 31  0 t = 2
rlabel pdiffusion 157 35 158 36  0 t = 3
rlabel pdiffusion 160 35 161 36  0 t = 4
rlabel pdiffusion 156 30 162 36 0 cell no = 10
<< m1 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2c >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< labels >>
rlabel pdiffusion 355 120 356 121  0 t = 1
rlabel pdiffusion 358 120 359 121  0 t = 2
rlabel pdiffusion 355 125 356 126  0 t = 3
rlabel pdiffusion 358 125 359 126  0 t = 4
rlabel pdiffusion 354 120 360 126 0 cell no = 11
<< m1 >>
rect 355 120 356 121 
rect 358 120 359 121 
rect 355 125 356 126 
rect 358 125 359 126 
<< m2 >>
rect 355 120 356 121 
rect 358 120 359 121 
rect 355 125 356 126 
rect 358 125 359 126 
<< m2c >>
rect 355 120 356 121 
rect 358 120 359 121 
rect 355 125 356 126 
rect 358 125 359 126 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 12
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 301 264 302 265  0 t = 1
rlabel pdiffusion 304 264 305 265  0 t = 2
rlabel pdiffusion 301 269 302 270  0 t = 3
rlabel pdiffusion 304 269 305 270  0 t = 4
rlabel pdiffusion 300 264 306 270 0 cell no = 13
<< m1 >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< m2 >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< m2c >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< labels >>
rlabel pdiffusion 139 12 140 13  0 t = 1
rlabel pdiffusion 142 12 143 13  0 t = 2
rlabel pdiffusion 139 17 140 18  0 t = 3
rlabel pdiffusion 142 17 143 18  0 t = 4
rlabel pdiffusion 138 12 144 18 0 cell no = 14
<< m1 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2c >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< labels >>
rlabel pdiffusion 265 12 266 13  0 t = 1
rlabel pdiffusion 268 12 269 13  0 t = 2
rlabel pdiffusion 265 17 266 18  0 t = 3
rlabel pdiffusion 268 17 269 18  0 t = 4
rlabel pdiffusion 264 12 270 18 0 cell no = 15
<< m1 >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< m2 >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< m2c >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< labels >>
rlabel pdiffusion 211 84 212 85  0 t = 1
rlabel pdiffusion 214 84 215 85  0 t = 2
rlabel pdiffusion 211 89 212 90  0 t = 3
rlabel pdiffusion 214 89 215 90  0 t = 4
rlabel pdiffusion 210 84 216 90 0 cell no = 16
<< m1 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2c >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< labels >>
rlabel pdiffusion 355 66 356 67  0 t = 1
rlabel pdiffusion 358 66 359 67  0 t = 2
rlabel pdiffusion 355 71 356 72  0 t = 3
rlabel pdiffusion 358 71 359 72  0 t = 4
rlabel pdiffusion 354 66 360 72 0 cell no = 17
<< m1 >>
rect 355 66 356 67 
rect 358 66 359 67 
rect 355 71 356 72 
rect 358 71 359 72 
<< m2 >>
rect 355 66 356 67 
rect 358 66 359 67 
rect 355 71 356 72 
rect 358 71 359 72 
<< m2c >>
rect 355 66 356 67 
rect 358 66 359 67 
rect 355 71 356 72 
rect 358 71 359 72 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 18
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 157 138 158 139  0 t = 1
rlabel pdiffusion 160 138 161 139  0 t = 2
rlabel pdiffusion 157 143 158 144  0 t = 3
rlabel pdiffusion 160 143 161 144  0 t = 4
rlabel pdiffusion 156 138 162 144 0 cell no = 19
<< m1 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2c >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< labels >>
rlabel pdiffusion 391 66 392 67  0 t = 1
rlabel pdiffusion 394 66 395 67  0 t = 2
rlabel pdiffusion 391 71 392 72  0 t = 3
rlabel pdiffusion 394 71 395 72  0 t = 4
rlabel pdiffusion 390 66 396 72 0 cell no = 20
<< m1 >>
rect 391 66 392 67 
rect 394 66 395 67 
rect 391 71 392 72 
rect 394 71 395 72 
<< m2 >>
rect 391 66 392 67 
rect 394 66 395 67 
rect 391 71 392 72 
rect 394 71 395 72 
<< m2c >>
rect 391 66 392 67 
rect 394 66 395 67 
rect 391 71 392 72 
rect 394 71 395 72 
<< labels >>
rlabel pdiffusion 409 30 410 31  0 t = 1
rlabel pdiffusion 412 30 413 31  0 t = 2
rlabel pdiffusion 409 35 410 36  0 t = 3
rlabel pdiffusion 412 35 413 36  0 t = 4
rlabel pdiffusion 408 30 414 36 0 cell no = 21
<< m1 >>
rect 409 30 410 31 
rect 412 30 413 31 
rect 409 35 410 36 
rect 412 35 413 36 
<< m2 >>
rect 409 30 410 31 
rect 412 30 413 31 
rect 409 35 410 36 
rect 412 35 413 36 
<< m2c >>
rect 409 30 410 31 
rect 412 30 413 31 
rect 409 35 410 36 
rect 412 35 413 36 
<< labels >>
rlabel pdiffusion 103 30 104 31  0 t = 1
rlabel pdiffusion 106 30 107 31  0 t = 2
rlabel pdiffusion 103 35 104 36  0 t = 3
rlabel pdiffusion 106 35 107 36  0 t = 4
rlabel pdiffusion 102 30 108 36 0 cell no = 22
<< m1 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2c >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< labels >>
rlabel pdiffusion 319 48 320 49  0 t = 1
rlabel pdiffusion 322 48 323 49  0 t = 2
rlabel pdiffusion 319 53 320 54  0 t = 3
rlabel pdiffusion 322 53 323 54  0 t = 4
rlabel pdiffusion 318 48 324 54 0 cell no = 23
<< m1 >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< m2 >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< m2c >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< labels >>
rlabel pdiffusion 301 84 302 85  0 t = 1
rlabel pdiffusion 304 84 305 85  0 t = 2
rlabel pdiffusion 301 89 302 90  0 t = 3
rlabel pdiffusion 304 89 305 90  0 t = 4
rlabel pdiffusion 300 84 306 90 0 cell no = 24
<< m1 >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< m2 >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< m2c >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< labels >>
rlabel pdiffusion 391 30 392 31  0 t = 1
rlabel pdiffusion 394 30 395 31  0 t = 2
rlabel pdiffusion 391 35 392 36  0 t = 3
rlabel pdiffusion 394 35 395 36  0 t = 4
rlabel pdiffusion 390 30 396 36 0 cell no = 25
<< m1 >>
rect 391 30 392 31 
rect 394 30 395 31 
rect 391 35 392 36 
rect 394 35 395 36 
<< m2 >>
rect 391 30 392 31 
rect 394 30 395 31 
rect 391 35 392 36 
rect 394 35 395 36 
<< m2c >>
rect 391 30 392 31 
rect 394 30 395 31 
rect 391 35 392 36 
rect 394 35 395 36 
<< labels >>
rlabel pdiffusion 103 84 104 85  0 t = 1
rlabel pdiffusion 106 84 107 85  0 t = 2
rlabel pdiffusion 103 89 104 90  0 t = 3
rlabel pdiffusion 106 89 107 90  0 t = 4
rlabel pdiffusion 102 84 108 90 0 cell no = 26
<< m1 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2c >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< labels >>
rlabel pdiffusion 13 228 14 229  0 t = 1
rlabel pdiffusion 16 228 17 229  0 t = 2
rlabel pdiffusion 13 233 14 234  0 t = 3
rlabel pdiffusion 16 233 17 234  0 t = 4
rlabel pdiffusion 12 228 18 234 0 cell no = 27
<< m1 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2c >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< labels >>
rlabel pdiffusion 31 138 32 139  0 t = 1
rlabel pdiffusion 34 138 35 139  0 t = 2
rlabel pdiffusion 31 143 32 144  0 t = 3
rlabel pdiffusion 34 143 35 144  0 t = 4
rlabel pdiffusion 30 138 36 144 0 cell no = 28
<< m1 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2c >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< labels >>
rlabel pdiffusion 283 228 284 229  0 t = 1
rlabel pdiffusion 286 228 287 229  0 t = 2
rlabel pdiffusion 283 233 284 234  0 t = 3
rlabel pdiffusion 286 233 287 234  0 t = 4
rlabel pdiffusion 282 228 288 234 0 cell no = 29
<< m1 >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< m2 >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< m2c >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< labels >>
rlabel pdiffusion 229 84 230 85  0 t = 1
rlabel pdiffusion 232 84 233 85  0 t = 2
rlabel pdiffusion 229 89 230 90  0 t = 3
rlabel pdiffusion 232 89 233 90  0 t = 4
rlabel pdiffusion 228 84 234 90 0 cell no = 30
<< m1 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2c >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< labels >>
rlabel pdiffusion 445 210 446 211  0 t = 1
rlabel pdiffusion 448 210 449 211  0 t = 2
rlabel pdiffusion 445 215 446 216  0 t = 3
rlabel pdiffusion 448 215 449 216  0 t = 4
rlabel pdiffusion 444 210 450 216 0 cell no = 31
<< m1 >>
rect 445 210 446 211 
rect 448 210 449 211 
rect 445 215 446 216 
rect 448 215 449 216 
<< m2 >>
rect 445 210 446 211 
rect 448 210 449 211 
rect 445 215 446 216 
rect 448 215 449 216 
<< m2c >>
rect 445 210 446 211 
rect 448 210 449 211 
rect 445 215 446 216 
rect 448 215 449 216 
<< labels >>
rlabel pdiffusion 193 246 194 247  0 t = 1
rlabel pdiffusion 196 246 197 247  0 t = 2
rlabel pdiffusion 193 251 194 252  0 t = 3
rlabel pdiffusion 196 251 197 252  0 t = 4
rlabel pdiffusion 192 246 198 252 0 cell no = 32
<< m1 >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< m2 >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< m2c >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 33
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 319 30 320 31  0 t = 1
rlabel pdiffusion 322 30 323 31  0 t = 2
rlabel pdiffusion 319 35 320 36  0 t = 3
rlabel pdiffusion 322 35 323 36  0 t = 4
rlabel pdiffusion 318 30 324 36 0 cell no = 34
<< m1 >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< m2 >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< m2c >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< labels >>
rlabel pdiffusion 229 12 230 13  0 t = 1
rlabel pdiffusion 232 12 233 13  0 t = 2
rlabel pdiffusion 229 17 230 18  0 t = 3
rlabel pdiffusion 232 17 233 18  0 t = 4
rlabel pdiffusion 228 12 234 18 0 cell no = 35
<< m1 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2c >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< labels >>
rlabel pdiffusion 301 246 302 247  0 t = 1
rlabel pdiffusion 304 246 305 247  0 t = 2
rlabel pdiffusion 301 251 302 252  0 t = 3
rlabel pdiffusion 304 251 305 252  0 t = 4
rlabel pdiffusion 300 246 306 252 0 cell no = 36
<< m1 >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< m2 >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< m2c >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< labels >>
rlabel pdiffusion 49 156 50 157  0 t = 1
rlabel pdiffusion 52 156 53 157  0 t = 2
rlabel pdiffusion 49 161 50 162  0 t = 3
rlabel pdiffusion 52 161 53 162  0 t = 4
rlabel pdiffusion 48 156 54 162 0 cell no = 37
<< m1 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2c >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< labels >>
rlabel pdiffusion 175 120 176 121  0 t = 1
rlabel pdiffusion 178 120 179 121  0 t = 2
rlabel pdiffusion 175 125 176 126  0 t = 3
rlabel pdiffusion 178 125 179 126  0 t = 4
rlabel pdiffusion 174 120 180 126 0 cell no = 38
<< m1 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2c >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< labels >>
rlabel pdiffusion 139 120 140 121  0 t = 1
rlabel pdiffusion 142 120 143 121  0 t = 2
rlabel pdiffusion 139 125 140 126  0 t = 3
rlabel pdiffusion 142 125 143 126  0 t = 4
rlabel pdiffusion 138 120 144 126 0 cell no = 39
<< m1 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2c >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< labels >>
rlabel pdiffusion 373 102 374 103  0 t = 1
rlabel pdiffusion 376 102 377 103  0 t = 2
rlabel pdiffusion 373 107 374 108  0 t = 3
rlabel pdiffusion 376 107 377 108  0 t = 4
rlabel pdiffusion 372 102 378 108 0 cell no = 40
<< m1 >>
rect 373 102 374 103 
rect 376 102 377 103 
rect 373 107 374 108 
rect 376 107 377 108 
<< m2 >>
rect 373 102 374 103 
rect 376 102 377 103 
rect 373 107 374 108 
rect 376 107 377 108 
<< m2c >>
rect 373 102 374 103 
rect 376 102 377 103 
rect 373 107 374 108 
rect 376 107 377 108 
<< labels >>
rlabel pdiffusion 427 12 428 13  0 t = 1
rlabel pdiffusion 430 12 431 13  0 t = 2
rlabel pdiffusion 427 17 428 18  0 t = 3
rlabel pdiffusion 430 17 431 18  0 t = 4
rlabel pdiffusion 426 12 432 18 0 cell no = 41
<< m1 >>
rect 427 12 428 13 
rect 430 12 431 13 
rect 427 17 428 18 
rect 430 17 431 18 
<< m2 >>
rect 427 12 428 13 
rect 430 12 431 13 
rect 427 17 428 18 
rect 430 17 431 18 
<< m2c >>
rect 427 12 428 13 
rect 430 12 431 13 
rect 427 17 428 18 
rect 430 17 431 18 
<< labels >>
rlabel pdiffusion 211 66 212 67  0 t = 1
rlabel pdiffusion 214 66 215 67  0 t = 2
rlabel pdiffusion 211 71 212 72  0 t = 3
rlabel pdiffusion 214 71 215 72  0 t = 4
rlabel pdiffusion 210 66 216 72 0 cell no = 42
<< m1 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2c >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< labels >>
rlabel pdiffusion 445 102 446 103  0 t = 1
rlabel pdiffusion 448 102 449 103  0 t = 2
rlabel pdiffusion 445 107 446 108  0 t = 3
rlabel pdiffusion 448 107 449 108  0 t = 4
rlabel pdiffusion 444 102 450 108 0 cell no = 43
<< m1 >>
rect 445 102 446 103 
rect 448 102 449 103 
rect 445 107 446 108 
rect 448 107 449 108 
<< m2 >>
rect 445 102 446 103 
rect 448 102 449 103 
rect 445 107 446 108 
rect 448 107 449 108 
<< m2c >>
rect 445 102 446 103 
rect 448 102 449 103 
rect 445 107 446 108 
rect 448 107 449 108 
<< labels >>
rlabel pdiffusion 247 12 248 13  0 t = 1
rlabel pdiffusion 250 12 251 13  0 t = 2
rlabel pdiffusion 247 17 248 18  0 t = 3
rlabel pdiffusion 250 17 251 18  0 t = 4
rlabel pdiffusion 246 12 252 18 0 cell no = 44
<< m1 >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< m2 >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< m2c >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< labels >>
rlabel pdiffusion 301 30 302 31  0 t = 1
rlabel pdiffusion 304 30 305 31  0 t = 2
rlabel pdiffusion 301 35 302 36  0 t = 3
rlabel pdiffusion 304 35 305 36  0 t = 4
rlabel pdiffusion 300 30 306 36 0 cell no = 45
<< m1 >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< m2 >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< m2c >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< labels >>
rlabel pdiffusion 445 12 446 13  0 t = 1
rlabel pdiffusion 448 12 449 13  0 t = 2
rlabel pdiffusion 445 17 446 18  0 t = 3
rlabel pdiffusion 448 17 449 18  0 t = 4
rlabel pdiffusion 444 12 450 18 0 cell no = 46
<< m1 >>
rect 445 12 446 13 
rect 448 12 449 13 
rect 445 17 446 18 
rect 448 17 449 18 
<< m2 >>
rect 445 12 446 13 
rect 448 12 449 13 
rect 445 17 446 18 
rect 448 17 449 18 
<< m2c >>
rect 445 12 446 13 
rect 448 12 449 13 
rect 445 17 446 18 
rect 448 17 449 18 
<< labels >>
rlabel pdiffusion 337 66 338 67  0 t = 1
rlabel pdiffusion 340 66 341 67  0 t = 2
rlabel pdiffusion 337 71 338 72  0 t = 3
rlabel pdiffusion 340 71 341 72  0 t = 4
rlabel pdiffusion 336 66 342 72 0 cell no = 47
<< m1 >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< m2 >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< m2c >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< labels >>
rlabel pdiffusion 301 102 302 103  0 t = 1
rlabel pdiffusion 304 102 305 103  0 t = 2
rlabel pdiffusion 301 107 302 108  0 t = 3
rlabel pdiffusion 304 107 305 108  0 t = 4
rlabel pdiffusion 300 102 306 108 0 cell no = 48
<< m1 >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< m2 >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< m2c >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< labels >>
rlabel pdiffusion 175 66 176 67  0 t = 1
rlabel pdiffusion 178 66 179 67  0 t = 2
rlabel pdiffusion 175 71 176 72  0 t = 3
rlabel pdiffusion 178 71 179 72  0 t = 4
rlabel pdiffusion 174 66 180 72 0 cell no = 49
<< m1 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2c >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< labels >>
rlabel pdiffusion 283 372 284 373  0 t = 1
rlabel pdiffusion 286 372 287 373  0 t = 2
rlabel pdiffusion 283 377 284 378  0 t = 3
rlabel pdiffusion 286 377 287 378  0 t = 4
rlabel pdiffusion 282 372 288 378 0 cell no = 50
<< m1 >>
rect 283 372 284 373 
rect 286 372 287 373 
rect 283 377 284 378 
rect 286 377 287 378 
<< m2 >>
rect 283 372 284 373 
rect 286 372 287 373 
rect 283 377 284 378 
rect 286 377 287 378 
<< m2c >>
rect 283 372 284 373 
rect 286 372 287 373 
rect 283 377 284 378 
rect 286 377 287 378 
<< labels >>
rlabel pdiffusion 67 336 68 337  0 t = 1
rlabel pdiffusion 70 336 71 337  0 t = 2
rlabel pdiffusion 67 341 68 342  0 t = 3
rlabel pdiffusion 70 341 71 342  0 t = 4
rlabel pdiffusion 66 336 72 342 0 cell no = 51
<< m1 >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< m2 >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< m2c >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< labels >>
rlabel pdiffusion 283 138 284 139  0 t = 1
rlabel pdiffusion 286 138 287 139  0 t = 2
rlabel pdiffusion 283 143 284 144  0 t = 3
rlabel pdiffusion 286 143 287 144  0 t = 4
rlabel pdiffusion 282 138 288 144 0 cell no = 52
<< m1 >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< m2 >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< m2c >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 53
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 54
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 121 300 122 301  0 t = 1
rlabel pdiffusion 124 300 125 301  0 t = 2
rlabel pdiffusion 121 305 122 306  0 t = 3
rlabel pdiffusion 124 305 125 306  0 t = 4
rlabel pdiffusion 120 300 126 306 0 cell no = 55
<< m1 >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< m2 >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< m2c >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< labels >>
rlabel pdiffusion 175 156 176 157  0 t = 1
rlabel pdiffusion 178 156 179 157  0 t = 2
rlabel pdiffusion 175 161 176 162  0 t = 3
rlabel pdiffusion 178 161 179 162  0 t = 4
rlabel pdiffusion 174 156 180 162 0 cell no = 56
<< m1 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2c >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< labels >>
rlabel pdiffusion 67 156 68 157  0 t = 1
rlabel pdiffusion 70 156 71 157  0 t = 2
rlabel pdiffusion 67 161 68 162  0 t = 3
rlabel pdiffusion 70 161 71 162  0 t = 4
rlabel pdiffusion 66 156 72 162 0 cell no = 57
<< m1 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2c >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 58
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 67 264 68 265  0 t = 1
rlabel pdiffusion 70 264 71 265  0 t = 2
rlabel pdiffusion 67 269 68 270  0 t = 3
rlabel pdiffusion 70 269 71 270  0 t = 4
rlabel pdiffusion 66 264 72 270 0 cell no = 59
<< m1 >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< m2 >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< m2c >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< labels >>
rlabel pdiffusion 247 102 248 103  0 t = 1
rlabel pdiffusion 250 102 251 103  0 t = 2
rlabel pdiffusion 247 107 248 108  0 t = 3
rlabel pdiffusion 250 107 251 108  0 t = 4
rlabel pdiffusion 246 102 252 108 0 cell no = 60
<< m1 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2c >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< labels >>
rlabel pdiffusion 355 354 356 355  0 t = 1
rlabel pdiffusion 358 354 359 355  0 t = 2
rlabel pdiffusion 355 359 356 360  0 t = 3
rlabel pdiffusion 358 359 359 360  0 t = 4
rlabel pdiffusion 354 354 360 360 0 cell no = 61
<< m1 >>
rect 355 354 356 355 
rect 358 354 359 355 
rect 355 359 356 360 
rect 358 359 359 360 
<< m2 >>
rect 355 354 356 355 
rect 358 354 359 355 
rect 355 359 356 360 
rect 358 359 359 360 
<< m2c >>
rect 355 354 356 355 
rect 358 354 359 355 
rect 355 359 356 360 
rect 358 359 359 360 
<< labels >>
rlabel pdiffusion 301 120 302 121  0 t = 1
rlabel pdiffusion 304 120 305 121  0 t = 2
rlabel pdiffusion 301 125 302 126  0 t = 3
rlabel pdiffusion 304 125 305 126  0 t = 4
rlabel pdiffusion 300 120 306 126 0 cell no = 62
<< m1 >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< m2 >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< m2c >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< labels >>
rlabel pdiffusion 373 66 374 67  0 t = 1
rlabel pdiffusion 376 66 377 67  0 t = 2
rlabel pdiffusion 373 71 374 72  0 t = 3
rlabel pdiffusion 376 71 377 72  0 t = 4
rlabel pdiffusion 372 66 378 72 0 cell no = 63
<< m1 >>
rect 373 66 374 67 
rect 376 66 377 67 
rect 373 71 374 72 
rect 376 71 377 72 
<< m2 >>
rect 373 66 374 67 
rect 376 66 377 67 
rect 373 71 374 72 
rect 376 71 377 72 
<< m2c >>
rect 373 66 374 67 
rect 376 66 377 67 
rect 373 71 374 72 
rect 376 71 377 72 
<< labels >>
rlabel pdiffusion 229 354 230 355  0 t = 1
rlabel pdiffusion 232 354 233 355  0 t = 2
rlabel pdiffusion 229 359 230 360  0 t = 3
rlabel pdiffusion 232 359 233 360  0 t = 4
rlabel pdiffusion 228 354 234 360 0 cell no = 64
<< m1 >>
rect 229 354 230 355 
rect 232 354 233 355 
rect 229 359 230 360 
rect 232 359 233 360 
<< m2 >>
rect 229 354 230 355 
rect 232 354 233 355 
rect 229 359 230 360 
rect 232 359 233 360 
<< m2c >>
rect 229 354 230 355 
rect 232 354 233 355 
rect 229 359 230 360 
rect 232 359 233 360 
<< labels >>
rlabel pdiffusion 445 66 446 67  0 t = 1
rlabel pdiffusion 448 66 449 67  0 t = 2
rlabel pdiffusion 445 71 446 72  0 t = 3
rlabel pdiffusion 448 71 449 72  0 t = 4
rlabel pdiffusion 444 66 450 72 0 cell no = 65
<< m1 >>
rect 445 66 446 67 
rect 448 66 449 67 
rect 445 71 446 72 
rect 448 71 449 72 
<< m2 >>
rect 445 66 446 67 
rect 448 66 449 67 
rect 445 71 446 72 
rect 448 71 449 72 
<< m2c >>
rect 445 66 446 67 
rect 448 66 449 67 
rect 445 71 446 72 
rect 448 71 449 72 
<< labels >>
rlabel pdiffusion 139 66 140 67  0 t = 1
rlabel pdiffusion 142 66 143 67  0 t = 2
rlabel pdiffusion 139 71 140 72  0 t = 3
rlabel pdiffusion 142 71 143 72  0 t = 4
rlabel pdiffusion 138 66 144 72 0 cell no = 66
<< m1 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2c >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< labels >>
rlabel pdiffusion 283 30 284 31  0 t = 1
rlabel pdiffusion 286 30 287 31  0 t = 2
rlabel pdiffusion 283 35 284 36  0 t = 3
rlabel pdiffusion 286 35 287 36  0 t = 4
rlabel pdiffusion 282 30 288 36 0 cell no = 67
<< m1 >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< m2 >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< m2c >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< labels >>
rlabel pdiffusion 409 48 410 49  0 t = 1
rlabel pdiffusion 412 48 413 49  0 t = 2
rlabel pdiffusion 409 53 410 54  0 t = 3
rlabel pdiffusion 412 53 413 54  0 t = 4
rlabel pdiffusion 408 48 414 54 0 cell no = 68
<< m1 >>
rect 409 48 410 49 
rect 412 48 413 49 
rect 409 53 410 54 
rect 412 53 413 54 
<< m2 >>
rect 409 48 410 49 
rect 412 48 413 49 
rect 409 53 410 54 
rect 412 53 413 54 
<< m2c >>
rect 409 48 410 49 
rect 412 48 413 49 
rect 409 53 410 54 
rect 412 53 413 54 
<< labels >>
rlabel pdiffusion 391 12 392 13  0 t = 1
rlabel pdiffusion 394 12 395 13  0 t = 2
rlabel pdiffusion 391 17 392 18  0 t = 3
rlabel pdiffusion 394 17 395 18  0 t = 4
rlabel pdiffusion 390 12 396 18 0 cell no = 69
<< m1 >>
rect 391 12 392 13 
rect 394 12 395 13 
rect 391 17 392 18 
rect 394 17 395 18 
<< m2 >>
rect 391 12 392 13 
rect 394 12 395 13 
rect 391 17 392 18 
rect 394 17 395 18 
<< m2c >>
rect 391 12 392 13 
rect 394 12 395 13 
rect 391 17 392 18 
rect 394 17 395 18 
<< labels >>
rlabel pdiffusion 427 48 428 49  0 t = 1
rlabel pdiffusion 430 48 431 49  0 t = 2
rlabel pdiffusion 427 53 428 54  0 t = 3
rlabel pdiffusion 430 53 431 54  0 t = 4
rlabel pdiffusion 426 48 432 54 0 cell no = 70
<< m1 >>
rect 427 48 428 49 
rect 430 48 431 49 
rect 427 53 428 54 
rect 430 53 431 54 
<< m2 >>
rect 427 48 428 49 
rect 430 48 431 49 
rect 427 53 428 54 
rect 430 53 431 54 
<< m2c >>
rect 427 48 428 49 
rect 430 48 431 49 
rect 427 53 428 54 
rect 430 53 431 54 
<< labels >>
rlabel pdiffusion 427 30 428 31  0 t = 1
rlabel pdiffusion 430 30 431 31  0 t = 2
rlabel pdiffusion 427 35 428 36  0 t = 3
rlabel pdiffusion 430 35 431 36  0 t = 4
rlabel pdiffusion 426 30 432 36 0 cell no = 71
<< m1 >>
rect 427 30 428 31 
rect 430 30 431 31 
rect 427 35 428 36 
rect 430 35 431 36 
<< m2 >>
rect 427 30 428 31 
rect 430 30 431 31 
rect 427 35 428 36 
rect 430 35 431 36 
<< m2c >>
rect 427 30 428 31 
rect 430 30 431 31 
rect 427 35 428 36 
rect 430 35 431 36 
<< labels >>
rlabel pdiffusion 355 12 356 13  0 t = 1
rlabel pdiffusion 358 12 359 13  0 t = 2
rlabel pdiffusion 355 17 356 18  0 t = 3
rlabel pdiffusion 358 17 359 18  0 t = 4
rlabel pdiffusion 354 12 360 18 0 cell no = 72
<< m1 >>
rect 355 12 356 13 
rect 358 12 359 13 
rect 355 17 356 18 
rect 358 17 359 18 
<< m2 >>
rect 355 12 356 13 
rect 358 12 359 13 
rect 355 17 356 18 
rect 358 17 359 18 
<< m2c >>
rect 355 12 356 13 
rect 358 12 359 13 
rect 355 17 356 18 
rect 358 17 359 18 
<< labels >>
rlabel pdiffusion 175 192 176 193  0 t = 1
rlabel pdiffusion 178 192 179 193  0 t = 2
rlabel pdiffusion 175 197 176 198  0 t = 3
rlabel pdiffusion 178 197 179 198  0 t = 4
rlabel pdiffusion 174 192 180 198 0 cell no = 73
<< m1 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2c >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< labels >>
rlabel pdiffusion 319 102 320 103  0 t = 1
rlabel pdiffusion 322 102 323 103  0 t = 2
rlabel pdiffusion 319 107 320 108  0 t = 3
rlabel pdiffusion 322 107 323 108  0 t = 4
rlabel pdiffusion 318 102 324 108 0 cell no = 74
<< m1 >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< m2 >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< m2c >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< labels >>
rlabel pdiffusion 427 66 428 67  0 t = 1
rlabel pdiffusion 430 66 431 67  0 t = 2
rlabel pdiffusion 427 71 428 72  0 t = 3
rlabel pdiffusion 430 71 431 72  0 t = 4
rlabel pdiffusion 426 66 432 72 0 cell no = 75
<< m1 >>
rect 427 66 428 67 
rect 430 66 431 67 
rect 427 71 428 72 
rect 430 71 431 72 
<< m2 >>
rect 427 66 428 67 
rect 430 66 431 67 
rect 427 71 428 72 
rect 430 71 431 72 
<< m2c >>
rect 427 66 428 67 
rect 430 66 431 67 
rect 427 71 428 72 
rect 430 71 431 72 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 76
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 157 66 158 67  0 t = 1
rlabel pdiffusion 160 66 161 67  0 t = 2
rlabel pdiffusion 157 71 158 72  0 t = 3
rlabel pdiffusion 160 71 161 72  0 t = 4
rlabel pdiffusion 156 66 162 72 0 cell no = 77
<< m1 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2c >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 78
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 337 336 338 337  0 t = 1
rlabel pdiffusion 340 336 341 337  0 t = 2
rlabel pdiffusion 337 341 338 342  0 t = 3
rlabel pdiffusion 340 341 341 342  0 t = 4
rlabel pdiffusion 336 336 342 342 0 cell no = 79
<< m1 >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< m2 >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< m2c >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 80
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 81
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 82
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< labels >>
rlabel pdiffusion 247 174 248 175  0 t = 1
rlabel pdiffusion 250 174 251 175  0 t = 2
rlabel pdiffusion 247 179 248 180  0 t = 3
rlabel pdiffusion 250 179 251 180  0 t = 4
rlabel pdiffusion 246 174 252 180 0 cell no = 83
<< m1 >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< m2 >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< m2c >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< labels >>
rlabel pdiffusion 283 264 284 265  0 t = 1
rlabel pdiffusion 286 264 287 265  0 t = 2
rlabel pdiffusion 283 269 284 270  0 t = 3
rlabel pdiffusion 286 269 287 270  0 t = 4
rlabel pdiffusion 282 264 288 270 0 cell no = 84
<< m1 >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< m2 >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< m2c >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< labels >>
rlabel pdiffusion 31 372 32 373  0 t = 1
rlabel pdiffusion 34 372 35 373  0 t = 2
rlabel pdiffusion 31 377 32 378  0 t = 3
rlabel pdiffusion 34 377 35 378  0 t = 4
rlabel pdiffusion 30 372 36 378 0 cell no = 85
<< m1 >>
rect 31 372 32 373 
rect 34 372 35 373 
rect 31 377 32 378 
rect 34 377 35 378 
<< m2 >>
rect 31 372 32 373 
rect 34 372 35 373 
rect 31 377 32 378 
rect 34 377 35 378 
<< m2c >>
rect 31 372 32 373 
rect 34 372 35 373 
rect 31 377 32 378 
rect 34 377 35 378 
<< labels >>
rlabel pdiffusion 337 156 338 157  0 t = 1
rlabel pdiffusion 340 156 341 157  0 t = 2
rlabel pdiffusion 337 161 338 162  0 t = 3
rlabel pdiffusion 340 161 341 162  0 t = 4
rlabel pdiffusion 336 156 342 162 0 cell no = 86
<< m1 >>
rect 337 156 338 157 
rect 340 156 341 157 
rect 337 161 338 162 
rect 340 161 341 162 
<< m2 >>
rect 337 156 338 157 
rect 340 156 341 157 
rect 337 161 338 162 
rect 340 161 341 162 
<< m2c >>
rect 337 156 338 157 
rect 340 156 341 157 
rect 337 161 338 162 
rect 340 161 341 162 
<< labels >>
rlabel pdiffusion 193 66 194 67  0 t = 1
rlabel pdiffusion 196 66 197 67  0 t = 2
rlabel pdiffusion 193 71 194 72  0 t = 3
rlabel pdiffusion 196 71 197 72  0 t = 4
rlabel pdiffusion 192 66 198 72 0 cell no = 87
<< m1 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2c >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 88
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 265 282 266 283  0 t = 1
rlabel pdiffusion 268 282 269 283  0 t = 2
rlabel pdiffusion 265 287 266 288  0 t = 3
rlabel pdiffusion 268 287 269 288  0 t = 4
rlabel pdiffusion 264 282 270 288 0 cell no = 89
<< m1 >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< m2 >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< m2c >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< labels >>
rlabel pdiffusion 337 30 338 31  0 t = 1
rlabel pdiffusion 340 30 341 31  0 t = 2
rlabel pdiffusion 337 35 338 36  0 t = 3
rlabel pdiffusion 340 35 341 36  0 t = 4
rlabel pdiffusion 336 30 342 36 0 cell no = 90
<< m1 >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< m2 >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< m2c >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< labels >>
rlabel pdiffusion 139 156 140 157  0 t = 1
rlabel pdiffusion 142 156 143 157  0 t = 2
rlabel pdiffusion 139 161 140 162  0 t = 3
rlabel pdiffusion 142 161 143 162  0 t = 4
rlabel pdiffusion 138 156 144 162 0 cell no = 91
<< m1 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2c >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< labels >>
rlabel pdiffusion 283 84 284 85  0 t = 1
rlabel pdiffusion 286 84 287 85  0 t = 2
rlabel pdiffusion 283 89 284 90  0 t = 3
rlabel pdiffusion 286 89 287 90  0 t = 4
rlabel pdiffusion 282 84 288 90 0 cell no = 92
<< m1 >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< m2 >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< m2c >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< labels >>
rlabel pdiffusion 85 138 86 139  0 t = 1
rlabel pdiffusion 88 138 89 139  0 t = 2
rlabel pdiffusion 85 143 86 144  0 t = 3
rlabel pdiffusion 88 143 89 144  0 t = 4
rlabel pdiffusion 84 138 90 144 0 cell no = 93
<< m1 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2c >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< labels >>
rlabel pdiffusion 409 282 410 283  0 t = 1
rlabel pdiffusion 412 282 413 283  0 t = 2
rlabel pdiffusion 409 287 410 288  0 t = 3
rlabel pdiffusion 412 287 413 288  0 t = 4
rlabel pdiffusion 408 282 414 288 0 cell no = 94
<< m1 >>
rect 409 282 410 283 
rect 412 282 413 283 
rect 409 287 410 288 
rect 412 287 413 288 
<< m2 >>
rect 409 282 410 283 
rect 412 282 413 283 
rect 409 287 410 288 
rect 412 287 413 288 
<< m2c >>
rect 409 282 410 283 
rect 412 282 413 283 
rect 409 287 410 288 
rect 412 287 413 288 
<< labels >>
rlabel pdiffusion 265 84 266 85  0 t = 1
rlabel pdiffusion 268 84 269 85  0 t = 2
rlabel pdiffusion 265 89 266 90  0 t = 3
rlabel pdiffusion 268 89 269 90  0 t = 4
rlabel pdiffusion 264 84 270 90 0 cell no = 95
<< m1 >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< m2 >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< m2c >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< labels >>
rlabel pdiffusion 391 48 392 49  0 t = 1
rlabel pdiffusion 394 48 395 49  0 t = 2
rlabel pdiffusion 391 53 392 54  0 t = 3
rlabel pdiffusion 394 53 395 54  0 t = 4
rlabel pdiffusion 390 48 396 54 0 cell no = 96
<< m1 >>
rect 391 48 392 49 
rect 394 48 395 49 
rect 391 53 392 54 
rect 394 53 395 54 
<< m2 >>
rect 391 48 392 49 
rect 394 48 395 49 
rect 391 53 392 54 
rect 394 53 395 54 
<< m2c >>
rect 391 48 392 49 
rect 394 48 395 49 
rect 391 53 392 54 
rect 394 53 395 54 
<< labels >>
rlabel pdiffusion 427 192 428 193  0 t = 1
rlabel pdiffusion 430 192 431 193  0 t = 2
rlabel pdiffusion 427 197 428 198  0 t = 3
rlabel pdiffusion 430 197 431 198  0 t = 4
rlabel pdiffusion 426 192 432 198 0 cell no = 97
<< m1 >>
rect 427 192 428 193 
rect 430 192 431 193 
rect 427 197 428 198 
rect 430 197 431 198 
<< m2 >>
rect 427 192 428 193 
rect 430 192 431 193 
rect 427 197 428 198 
rect 430 197 431 198 
<< m2c >>
rect 427 192 428 193 
rect 430 192 431 193 
rect 427 197 428 198 
rect 430 197 431 198 
<< labels >>
rlabel pdiffusion 409 102 410 103  0 t = 1
rlabel pdiffusion 412 102 413 103  0 t = 2
rlabel pdiffusion 409 107 410 108  0 t = 3
rlabel pdiffusion 412 107 413 108  0 t = 4
rlabel pdiffusion 408 102 414 108 0 cell no = 98
<< m1 >>
rect 409 102 410 103 
rect 412 102 413 103 
rect 409 107 410 108 
rect 412 107 413 108 
<< m2 >>
rect 409 102 410 103 
rect 412 102 413 103 
rect 409 107 410 108 
rect 412 107 413 108 
<< m2c >>
rect 409 102 410 103 
rect 412 102 413 103 
rect 409 107 410 108 
rect 412 107 413 108 
<< labels >>
rlabel pdiffusion 373 30 374 31  0 t = 1
rlabel pdiffusion 376 30 377 31  0 t = 2
rlabel pdiffusion 373 35 374 36  0 t = 3
rlabel pdiffusion 376 35 377 36  0 t = 4
rlabel pdiffusion 372 30 378 36 0 cell no = 99
<< m1 >>
rect 373 30 374 31 
rect 376 30 377 31 
rect 373 35 374 36 
rect 376 35 377 36 
<< m2 >>
rect 373 30 374 31 
rect 376 30 377 31 
rect 373 35 374 36 
rect 376 35 377 36 
<< m2c >>
rect 373 30 374 31 
rect 376 30 377 31 
rect 373 35 374 36 
rect 376 35 377 36 
<< labels >>
rlabel pdiffusion 67 138 68 139  0 t = 1
rlabel pdiffusion 70 138 71 139  0 t = 2
rlabel pdiffusion 67 143 68 144  0 t = 3
rlabel pdiffusion 70 143 71 144  0 t = 4
rlabel pdiffusion 66 138 72 144 0 cell no = 100
<< m1 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2c >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< labels >>
rlabel pdiffusion 67 318 68 319  0 t = 1
rlabel pdiffusion 70 318 71 319  0 t = 2
rlabel pdiffusion 67 323 68 324  0 t = 3
rlabel pdiffusion 70 323 71 324  0 t = 4
rlabel pdiffusion 66 318 72 324 0 cell no = 101
<< m1 >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< m2 >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< m2c >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< labels >>
rlabel pdiffusion 49 120 50 121  0 t = 1
rlabel pdiffusion 52 120 53 121  0 t = 2
rlabel pdiffusion 49 125 50 126  0 t = 3
rlabel pdiffusion 52 125 53 126  0 t = 4
rlabel pdiffusion 48 120 54 126 0 cell no = 102
<< m1 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2c >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< labels >>
rlabel pdiffusion 103 174 104 175  0 t = 1
rlabel pdiffusion 106 174 107 175  0 t = 2
rlabel pdiffusion 103 179 104 180  0 t = 3
rlabel pdiffusion 106 179 107 180  0 t = 4
rlabel pdiffusion 102 174 108 180 0 cell no = 103
<< m1 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2c >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< labels >>
rlabel pdiffusion 247 228 248 229  0 t = 1
rlabel pdiffusion 250 228 251 229  0 t = 2
rlabel pdiffusion 247 233 248 234  0 t = 3
rlabel pdiffusion 250 233 251 234  0 t = 4
rlabel pdiffusion 246 228 252 234 0 cell no = 104
<< m1 >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< m2 >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< m2c >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< labels >>
rlabel pdiffusion 85 12 86 13  0 t = 1
rlabel pdiffusion 88 12 89 13  0 t = 2
rlabel pdiffusion 85 17 86 18  0 t = 3
rlabel pdiffusion 88 17 89 18  0 t = 4
rlabel pdiffusion 84 12 90 18 0 cell no = 105
<< m1 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2c >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< labels >>
rlabel pdiffusion 283 48 284 49  0 t = 1
rlabel pdiffusion 286 48 287 49  0 t = 2
rlabel pdiffusion 283 53 284 54  0 t = 3
rlabel pdiffusion 286 53 287 54  0 t = 4
rlabel pdiffusion 282 48 288 54 0 cell no = 106
<< m1 >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< m2 >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< m2c >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 107
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 157 102 158 103  0 t = 1
rlabel pdiffusion 160 102 161 103  0 t = 2
rlabel pdiffusion 157 107 158 108  0 t = 3
rlabel pdiffusion 160 107 161 108  0 t = 4
rlabel pdiffusion 156 102 162 108 0 cell no = 108
<< m1 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2c >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< labels >>
rlabel pdiffusion 103 300 104 301  0 t = 1
rlabel pdiffusion 106 300 107 301  0 t = 2
rlabel pdiffusion 103 305 104 306  0 t = 3
rlabel pdiffusion 106 305 107 306  0 t = 4
rlabel pdiffusion 102 300 108 306 0 cell no = 109
<< m1 >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< m2 >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< m2c >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< labels >>
rlabel pdiffusion 283 210 284 211  0 t = 1
rlabel pdiffusion 286 210 287 211  0 t = 2
rlabel pdiffusion 283 215 284 216  0 t = 3
rlabel pdiffusion 286 215 287 216  0 t = 4
rlabel pdiffusion 282 210 288 216 0 cell no = 110
<< m1 >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< m2 >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< m2c >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< labels >>
rlabel pdiffusion 211 12 212 13  0 t = 1
rlabel pdiffusion 214 12 215 13  0 t = 2
rlabel pdiffusion 211 17 212 18  0 t = 3
rlabel pdiffusion 214 17 215 18  0 t = 4
rlabel pdiffusion 210 12 216 18 0 cell no = 111
<< m1 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2c >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< labels >>
rlabel pdiffusion 121 174 122 175  0 t = 1
rlabel pdiffusion 124 174 125 175  0 t = 2
rlabel pdiffusion 121 179 122 180  0 t = 3
rlabel pdiffusion 124 179 125 180  0 t = 4
rlabel pdiffusion 120 174 126 180 0 cell no = 112
<< m1 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2c >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< labels >>
rlabel pdiffusion 175 12 176 13  0 t = 1
rlabel pdiffusion 178 12 179 13  0 t = 2
rlabel pdiffusion 175 17 176 18  0 t = 3
rlabel pdiffusion 178 17 179 18  0 t = 4
rlabel pdiffusion 174 12 180 18 0 cell no = 113
<< m1 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2c >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< labels >>
rlabel pdiffusion 49 192 50 193  0 t = 1
rlabel pdiffusion 52 192 53 193  0 t = 2
rlabel pdiffusion 49 197 50 198  0 t = 3
rlabel pdiffusion 52 197 53 198  0 t = 4
rlabel pdiffusion 48 192 54 198 0 cell no = 114
<< m1 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2c >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< labels >>
rlabel pdiffusion 427 84 428 85  0 t = 1
rlabel pdiffusion 430 84 431 85  0 t = 2
rlabel pdiffusion 427 89 428 90  0 t = 3
rlabel pdiffusion 430 89 431 90  0 t = 4
rlabel pdiffusion 426 84 432 90 0 cell no = 115
<< m1 >>
rect 427 84 428 85 
rect 430 84 431 85 
rect 427 89 428 90 
rect 430 89 431 90 
<< m2 >>
rect 427 84 428 85 
rect 430 84 431 85 
rect 427 89 428 90 
rect 430 89 431 90 
<< m2c >>
rect 427 84 428 85 
rect 430 84 431 85 
rect 427 89 428 90 
rect 430 89 431 90 
<< labels >>
rlabel pdiffusion 301 66 302 67  0 t = 1
rlabel pdiffusion 304 66 305 67  0 t = 2
rlabel pdiffusion 301 71 302 72  0 t = 3
rlabel pdiffusion 304 71 305 72  0 t = 4
rlabel pdiffusion 300 66 306 72 0 cell no = 116
<< m1 >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< m2 >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< m2c >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< labels >>
rlabel pdiffusion 391 120 392 121  0 t = 1
rlabel pdiffusion 394 120 395 121  0 t = 2
rlabel pdiffusion 391 125 392 126  0 t = 3
rlabel pdiffusion 394 125 395 126  0 t = 4
rlabel pdiffusion 390 120 396 126 0 cell no = 117
<< m1 >>
rect 391 120 392 121 
rect 394 120 395 121 
rect 391 125 392 126 
rect 394 125 395 126 
<< m2 >>
rect 391 120 392 121 
rect 394 120 395 121 
rect 391 125 392 126 
rect 394 125 395 126 
<< m2c >>
rect 391 120 392 121 
rect 394 120 395 121 
rect 391 125 392 126 
rect 394 125 395 126 
<< labels >>
rlabel pdiffusion 211 156 212 157  0 t = 1
rlabel pdiffusion 214 156 215 157  0 t = 2
rlabel pdiffusion 211 161 212 162  0 t = 3
rlabel pdiffusion 214 161 215 162  0 t = 4
rlabel pdiffusion 210 156 216 162 0 cell no = 118
<< m1 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2c >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< labels >>
rlabel pdiffusion 121 138 122 139  0 t = 1
rlabel pdiffusion 124 138 125 139  0 t = 2
rlabel pdiffusion 121 143 122 144  0 t = 3
rlabel pdiffusion 124 143 125 144  0 t = 4
rlabel pdiffusion 120 138 126 144 0 cell no = 119
<< m1 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2c >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< labels >>
rlabel pdiffusion 283 66 284 67  0 t = 1
rlabel pdiffusion 286 66 287 67  0 t = 2
rlabel pdiffusion 283 71 284 72  0 t = 3
rlabel pdiffusion 286 71 287 72  0 t = 4
rlabel pdiffusion 282 66 288 72 0 cell no = 120
<< m1 >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< m2 >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< m2c >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< labels >>
rlabel pdiffusion 301 48 302 49  0 t = 1
rlabel pdiffusion 304 48 305 49  0 t = 2
rlabel pdiffusion 301 53 302 54  0 t = 3
rlabel pdiffusion 304 53 305 54  0 t = 4
rlabel pdiffusion 300 48 306 54 0 cell no = 121
<< m1 >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< m2 >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< m2c >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< labels >>
rlabel pdiffusion 427 156 428 157  0 t = 1
rlabel pdiffusion 430 156 431 157  0 t = 2
rlabel pdiffusion 427 161 428 162  0 t = 3
rlabel pdiffusion 430 161 431 162  0 t = 4
rlabel pdiffusion 426 156 432 162 0 cell no = 122
<< m1 >>
rect 427 156 428 157 
rect 430 156 431 157 
rect 427 161 428 162 
rect 430 161 431 162 
<< m2 >>
rect 427 156 428 157 
rect 430 156 431 157 
rect 427 161 428 162 
rect 430 161 431 162 
<< m2c >>
rect 427 156 428 157 
rect 430 156 431 157 
rect 427 161 428 162 
rect 430 161 431 162 
<< labels >>
rlabel pdiffusion 355 102 356 103  0 t = 1
rlabel pdiffusion 358 102 359 103  0 t = 2
rlabel pdiffusion 355 107 356 108  0 t = 3
rlabel pdiffusion 358 107 359 108  0 t = 4
rlabel pdiffusion 354 102 360 108 0 cell no = 123
<< m1 >>
rect 355 102 356 103 
rect 358 102 359 103 
rect 355 107 356 108 
rect 358 107 359 108 
<< m2 >>
rect 355 102 356 103 
rect 358 102 359 103 
rect 355 107 356 108 
rect 358 107 359 108 
<< m2c >>
rect 355 102 356 103 
rect 358 102 359 103 
rect 355 107 356 108 
rect 358 107 359 108 
<< labels >>
rlabel pdiffusion 409 120 410 121  0 t = 1
rlabel pdiffusion 412 120 413 121  0 t = 2
rlabel pdiffusion 409 125 410 126  0 t = 3
rlabel pdiffusion 412 125 413 126  0 t = 4
rlabel pdiffusion 408 120 414 126 0 cell no = 124
<< m1 >>
rect 409 120 410 121 
rect 412 120 413 121 
rect 409 125 410 126 
rect 412 125 413 126 
<< m2 >>
rect 409 120 410 121 
rect 412 120 413 121 
rect 409 125 410 126 
rect 412 125 413 126 
<< m2c >>
rect 409 120 410 121 
rect 412 120 413 121 
rect 409 125 410 126 
rect 412 125 413 126 
<< labels >>
rlabel pdiffusion 445 84 446 85  0 t = 1
rlabel pdiffusion 448 84 449 85  0 t = 2
rlabel pdiffusion 445 89 446 90  0 t = 3
rlabel pdiffusion 448 89 449 90  0 t = 4
rlabel pdiffusion 444 84 450 90 0 cell no = 125
<< m1 >>
rect 445 84 446 85 
rect 448 84 449 85 
rect 445 89 446 90 
rect 448 89 449 90 
<< m2 >>
rect 445 84 446 85 
rect 448 84 449 85 
rect 445 89 446 90 
rect 448 89 449 90 
<< m2c >>
rect 445 84 446 85 
rect 448 84 449 85 
rect 445 89 446 90 
rect 448 89 449 90 
<< labels >>
rlabel pdiffusion 193 120 194 121  0 t = 1
rlabel pdiffusion 196 120 197 121  0 t = 2
rlabel pdiffusion 193 125 194 126  0 t = 3
rlabel pdiffusion 196 125 197 126  0 t = 4
rlabel pdiffusion 192 120 198 126 0 cell no = 126
<< m1 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2c >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< labels >>
rlabel pdiffusion 175 246 176 247  0 t = 1
rlabel pdiffusion 178 246 179 247  0 t = 2
rlabel pdiffusion 175 251 176 252  0 t = 3
rlabel pdiffusion 178 251 179 252  0 t = 4
rlabel pdiffusion 174 246 180 252 0 cell no = 127
<< m1 >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< m2 >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< m2c >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 128
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 301 210 302 211  0 t = 1
rlabel pdiffusion 304 210 305 211  0 t = 2
rlabel pdiffusion 301 215 302 216  0 t = 3
rlabel pdiffusion 304 215 305 216  0 t = 4
rlabel pdiffusion 300 210 306 216 0 cell no = 129
<< m1 >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< m2 >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< m2c >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 130
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 121 102 122 103  0 t = 1
rlabel pdiffusion 124 102 125 103  0 t = 2
rlabel pdiffusion 121 107 122 108  0 t = 3
rlabel pdiffusion 124 107 125 108  0 t = 4
rlabel pdiffusion 120 102 126 108 0 cell no = 131
<< m1 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2c >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< labels >>
rlabel pdiffusion 157 84 158 85  0 t = 1
rlabel pdiffusion 160 84 161 85  0 t = 2
rlabel pdiffusion 157 89 158 90  0 t = 3
rlabel pdiffusion 160 89 161 90  0 t = 4
rlabel pdiffusion 156 84 162 90 0 cell no = 132
<< m1 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2c >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< labels >>
rlabel pdiffusion 13 336 14 337  0 t = 1
rlabel pdiffusion 16 336 17 337  0 t = 2
rlabel pdiffusion 13 341 14 342  0 t = 3
rlabel pdiffusion 16 341 17 342  0 t = 4
rlabel pdiffusion 12 336 18 342 0 cell no = 133
<< m1 >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< m2 >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< m2c >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< labels >>
rlabel pdiffusion 31 192 32 193  0 t = 1
rlabel pdiffusion 34 192 35 193  0 t = 2
rlabel pdiffusion 31 197 32 198  0 t = 3
rlabel pdiffusion 34 197 35 198  0 t = 4
rlabel pdiffusion 30 192 36 198 0 cell no = 134
<< m1 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2c >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< labels >>
rlabel pdiffusion 229 192 230 193  0 t = 1
rlabel pdiffusion 232 192 233 193  0 t = 2
rlabel pdiffusion 229 197 230 198  0 t = 3
rlabel pdiffusion 232 197 233 198  0 t = 4
rlabel pdiffusion 228 192 234 198 0 cell no = 135
<< m1 >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< m2 >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< m2c >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< labels >>
rlabel pdiffusion 211 138 212 139  0 t = 1
rlabel pdiffusion 214 138 215 139  0 t = 2
rlabel pdiffusion 211 143 212 144  0 t = 3
rlabel pdiffusion 214 143 215 144  0 t = 4
rlabel pdiffusion 210 138 216 144 0 cell no = 136
<< m1 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2c >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< labels >>
rlabel pdiffusion 139 282 140 283  0 t = 1
rlabel pdiffusion 142 282 143 283  0 t = 2
rlabel pdiffusion 139 287 140 288  0 t = 3
rlabel pdiffusion 142 287 143 288  0 t = 4
rlabel pdiffusion 138 282 144 288 0 cell no = 137
<< m1 >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< m2 >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< m2c >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< labels >>
rlabel pdiffusion 319 84 320 85  0 t = 1
rlabel pdiffusion 322 84 323 85  0 t = 2
rlabel pdiffusion 319 89 320 90  0 t = 3
rlabel pdiffusion 322 89 323 90  0 t = 4
rlabel pdiffusion 318 84 324 90 0 cell no = 138
<< m1 >>
rect 319 84 320 85 
rect 322 84 323 85 
rect 319 89 320 90 
rect 322 89 323 90 
<< m2 >>
rect 319 84 320 85 
rect 322 84 323 85 
rect 319 89 320 90 
rect 322 89 323 90 
<< m2c >>
rect 319 84 320 85 
rect 322 84 323 85 
rect 319 89 320 90 
rect 322 89 323 90 
<< labels >>
rlabel pdiffusion 265 102 266 103  0 t = 1
rlabel pdiffusion 268 102 269 103  0 t = 2
rlabel pdiffusion 265 107 266 108  0 t = 3
rlabel pdiffusion 268 107 269 108  0 t = 4
rlabel pdiffusion 264 102 270 108 0 cell no = 139
<< m1 >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< m2 >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< m2c >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< labels >>
rlabel pdiffusion 337 138 338 139  0 t = 1
rlabel pdiffusion 340 138 341 139  0 t = 2
rlabel pdiffusion 337 143 338 144  0 t = 3
rlabel pdiffusion 340 143 341 144  0 t = 4
rlabel pdiffusion 336 138 342 144 0 cell no = 140
<< m1 >>
rect 337 138 338 139 
rect 340 138 341 139 
rect 337 143 338 144 
rect 340 143 341 144 
<< m2 >>
rect 337 138 338 139 
rect 340 138 341 139 
rect 337 143 338 144 
rect 340 143 341 144 
<< m2c >>
rect 337 138 338 139 
rect 340 138 341 139 
rect 337 143 338 144 
rect 340 143 341 144 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 141
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 229 30 230 31  0 t = 1
rlabel pdiffusion 232 30 233 31  0 t = 2
rlabel pdiffusion 229 35 230 36  0 t = 3
rlabel pdiffusion 232 35 233 36  0 t = 4
rlabel pdiffusion 228 30 234 36 0 cell no = 142
<< m1 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2c >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< labels >>
rlabel pdiffusion 391 174 392 175  0 t = 1
rlabel pdiffusion 394 174 395 175  0 t = 2
rlabel pdiffusion 391 179 392 180  0 t = 3
rlabel pdiffusion 394 179 395 180  0 t = 4
rlabel pdiffusion 390 174 396 180 0 cell no = 143
<< m1 >>
rect 391 174 392 175 
rect 394 174 395 175 
rect 391 179 392 180 
rect 394 179 395 180 
<< m2 >>
rect 391 174 392 175 
rect 394 174 395 175 
rect 391 179 392 180 
rect 394 179 395 180 
<< m2c >>
rect 391 174 392 175 
rect 394 174 395 175 
rect 391 179 392 180 
rect 394 179 395 180 
<< labels >>
rlabel pdiffusion 409 138 410 139  0 t = 1
rlabel pdiffusion 412 138 413 139  0 t = 2
rlabel pdiffusion 409 143 410 144  0 t = 3
rlabel pdiffusion 412 143 413 144  0 t = 4
rlabel pdiffusion 408 138 414 144 0 cell no = 144
<< m1 >>
rect 409 138 410 139 
rect 412 138 413 139 
rect 409 143 410 144 
rect 412 143 413 144 
<< m2 >>
rect 409 138 410 139 
rect 412 138 413 139 
rect 409 143 410 144 
rect 412 143 413 144 
<< m2c >>
rect 409 138 410 139 
rect 412 138 413 139 
rect 409 143 410 144 
rect 412 143 413 144 
<< labels >>
rlabel pdiffusion 337 48 338 49  0 t = 1
rlabel pdiffusion 340 48 341 49  0 t = 2
rlabel pdiffusion 337 53 338 54  0 t = 3
rlabel pdiffusion 340 53 341 54  0 t = 4
rlabel pdiffusion 336 48 342 54 0 cell no = 145
<< m1 >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< m2 >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< m2c >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< labels >>
rlabel pdiffusion 157 228 158 229  0 t = 1
rlabel pdiffusion 160 228 161 229  0 t = 2
rlabel pdiffusion 157 233 158 234  0 t = 3
rlabel pdiffusion 160 233 161 234  0 t = 4
rlabel pdiffusion 156 228 162 234 0 cell no = 146
<< m1 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2c >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< labels >>
rlabel pdiffusion 445 228 446 229  0 t = 1
rlabel pdiffusion 448 228 449 229  0 t = 2
rlabel pdiffusion 445 233 446 234  0 t = 3
rlabel pdiffusion 448 233 449 234  0 t = 4
rlabel pdiffusion 444 228 450 234 0 cell no = 147
<< m1 >>
rect 445 228 446 229 
rect 448 228 449 229 
rect 445 233 446 234 
rect 448 233 449 234 
<< m2 >>
rect 445 228 446 229 
rect 448 228 449 229 
rect 445 233 446 234 
rect 448 233 449 234 
<< m2c >>
rect 445 228 446 229 
rect 448 228 449 229 
rect 445 233 446 234 
rect 448 233 449 234 
<< labels >>
rlabel pdiffusion 355 48 356 49  0 t = 1
rlabel pdiffusion 358 48 359 49  0 t = 2
rlabel pdiffusion 355 53 356 54  0 t = 3
rlabel pdiffusion 358 53 359 54  0 t = 4
rlabel pdiffusion 354 48 360 54 0 cell no = 148
<< m1 >>
rect 355 48 356 49 
rect 358 48 359 49 
rect 355 53 356 54 
rect 358 53 359 54 
<< m2 >>
rect 355 48 356 49 
rect 358 48 359 49 
rect 355 53 356 54 
rect 358 53 359 54 
<< m2c >>
rect 355 48 356 49 
rect 358 48 359 49 
rect 355 53 356 54 
rect 358 53 359 54 
<< labels >>
rlabel pdiffusion 427 228 428 229  0 t = 1
rlabel pdiffusion 430 228 431 229  0 t = 2
rlabel pdiffusion 427 233 428 234  0 t = 3
rlabel pdiffusion 430 233 431 234  0 t = 4
rlabel pdiffusion 426 228 432 234 0 cell no = 149
<< m1 >>
rect 427 228 428 229 
rect 430 228 431 229 
rect 427 233 428 234 
rect 430 233 431 234 
<< m2 >>
rect 427 228 428 229 
rect 430 228 431 229 
rect 427 233 428 234 
rect 430 233 431 234 
<< m2c >>
rect 427 228 428 229 
rect 430 228 431 229 
rect 427 233 428 234 
rect 430 233 431 234 
<< labels >>
rlabel pdiffusion 409 66 410 67  0 t = 1
rlabel pdiffusion 412 66 413 67  0 t = 2
rlabel pdiffusion 409 71 410 72  0 t = 3
rlabel pdiffusion 412 71 413 72  0 t = 4
rlabel pdiffusion 408 66 414 72 0 cell no = 150
<< m1 >>
rect 409 66 410 67 
rect 412 66 413 67 
rect 409 71 410 72 
rect 412 71 413 72 
<< m2 >>
rect 409 66 410 67 
rect 412 66 413 67 
rect 409 71 410 72 
rect 412 71 413 72 
<< m2c >>
rect 409 66 410 67 
rect 412 66 413 67 
rect 409 71 410 72 
rect 412 71 413 72 
<< labels >>
rlabel pdiffusion 139 210 140 211  0 t = 1
rlabel pdiffusion 142 210 143 211  0 t = 2
rlabel pdiffusion 139 215 140 216  0 t = 3
rlabel pdiffusion 142 215 143 216  0 t = 4
rlabel pdiffusion 138 210 144 216 0 cell no = 151
<< m1 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2c >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< labels >>
rlabel pdiffusion 265 192 266 193  0 t = 1
rlabel pdiffusion 268 192 269 193  0 t = 2
rlabel pdiffusion 265 197 266 198  0 t = 3
rlabel pdiffusion 268 197 269 198  0 t = 4
rlabel pdiffusion 264 192 270 198 0 cell no = 152
<< m1 >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< m2 >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< m2c >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 153
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 49 174 50 175  0 t = 1
rlabel pdiffusion 52 174 53 175  0 t = 2
rlabel pdiffusion 49 179 50 180  0 t = 3
rlabel pdiffusion 52 179 53 180  0 t = 4
rlabel pdiffusion 48 174 54 180 0 cell no = 154
<< m1 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2c >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< labels >>
rlabel pdiffusion 85 120 86 121  0 t = 1
rlabel pdiffusion 88 120 89 121  0 t = 2
rlabel pdiffusion 85 125 86 126  0 t = 3
rlabel pdiffusion 88 125 89 126  0 t = 4
rlabel pdiffusion 84 120 90 126 0 cell no = 155
<< m1 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2c >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< labels >>
rlabel pdiffusion 85 174 86 175  0 t = 1
rlabel pdiffusion 88 174 89 175  0 t = 2
rlabel pdiffusion 85 179 86 180  0 t = 3
rlabel pdiffusion 88 179 89 180  0 t = 4
rlabel pdiffusion 84 174 90 180 0 cell no = 156
<< m1 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2c >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< labels >>
rlabel pdiffusion 211 372 212 373  0 t = 1
rlabel pdiffusion 214 372 215 373  0 t = 2
rlabel pdiffusion 211 377 212 378  0 t = 3
rlabel pdiffusion 214 377 215 378  0 t = 4
rlabel pdiffusion 210 372 216 378 0 cell no = 157
<< m1 >>
rect 211 372 212 373 
rect 214 372 215 373 
rect 211 377 212 378 
rect 214 377 215 378 
<< m2 >>
rect 211 372 212 373 
rect 214 372 215 373 
rect 211 377 212 378 
rect 214 377 215 378 
<< m2c >>
rect 211 372 212 373 
rect 214 372 215 373 
rect 211 377 212 378 
rect 214 377 215 378 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 158
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 67 120 68 121  0 t = 1
rlabel pdiffusion 70 120 71 121  0 t = 2
rlabel pdiffusion 67 125 68 126  0 t = 3
rlabel pdiffusion 70 125 71 126  0 t = 4
rlabel pdiffusion 66 120 72 126 0 cell no = 159
<< m1 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2c >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< labels >>
rlabel pdiffusion 31 210 32 211  0 t = 1
rlabel pdiffusion 34 210 35 211  0 t = 2
rlabel pdiffusion 31 215 32 216  0 t = 3
rlabel pdiffusion 34 215 35 216  0 t = 4
rlabel pdiffusion 30 210 36 216 0 cell no = 160
<< m1 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2c >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< labels >>
rlabel pdiffusion 175 84 176 85  0 t = 1
rlabel pdiffusion 178 84 179 85  0 t = 2
rlabel pdiffusion 175 89 176 90  0 t = 3
rlabel pdiffusion 178 89 179 90  0 t = 4
rlabel pdiffusion 174 84 180 90 0 cell no = 161
<< m1 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2c >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< labels >>
rlabel pdiffusion 211 210 212 211  0 t = 1
rlabel pdiffusion 214 210 215 211  0 t = 2
rlabel pdiffusion 211 215 212 216  0 t = 3
rlabel pdiffusion 214 215 215 216  0 t = 4
rlabel pdiffusion 210 210 216 216 0 cell no = 162
<< m1 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2c >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< labels >>
rlabel pdiffusion 85 282 86 283  0 t = 1
rlabel pdiffusion 88 282 89 283  0 t = 2
rlabel pdiffusion 85 287 86 288  0 t = 3
rlabel pdiffusion 88 287 89 288  0 t = 4
rlabel pdiffusion 84 282 90 288 0 cell no = 163
<< m1 >>
rect 85 282 86 283 
rect 88 282 89 283 
rect 85 287 86 288 
rect 88 287 89 288 
<< m2 >>
rect 85 282 86 283 
rect 88 282 89 283 
rect 85 287 86 288 
rect 88 287 89 288 
<< m2c >>
rect 85 282 86 283 
rect 88 282 89 283 
rect 85 287 86 288 
rect 88 287 89 288 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 164
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 373 84 374 85  0 t = 1
rlabel pdiffusion 376 84 377 85  0 t = 2
rlabel pdiffusion 373 89 374 90  0 t = 3
rlabel pdiffusion 376 89 377 90  0 t = 4
rlabel pdiffusion 372 84 378 90 0 cell no = 165
<< m1 >>
rect 373 84 374 85 
rect 376 84 377 85 
rect 373 89 374 90 
rect 376 89 377 90 
<< m2 >>
rect 373 84 374 85 
rect 376 84 377 85 
rect 373 89 374 90 
rect 376 89 377 90 
<< m2c >>
rect 373 84 374 85 
rect 376 84 377 85 
rect 373 89 374 90 
rect 376 89 377 90 
<< labels >>
rlabel pdiffusion 391 156 392 157  0 t = 1
rlabel pdiffusion 394 156 395 157  0 t = 2
rlabel pdiffusion 391 161 392 162  0 t = 3
rlabel pdiffusion 394 161 395 162  0 t = 4
rlabel pdiffusion 390 156 396 162 0 cell no = 166
<< m1 >>
rect 391 156 392 157 
rect 394 156 395 157 
rect 391 161 392 162 
rect 394 161 395 162 
<< m2 >>
rect 391 156 392 157 
rect 394 156 395 157 
rect 391 161 392 162 
rect 394 161 395 162 
<< m2c >>
rect 391 156 392 157 
rect 394 156 395 157 
rect 391 161 392 162 
rect 394 161 395 162 
<< labels >>
rlabel pdiffusion 301 138 302 139  0 t = 1
rlabel pdiffusion 304 138 305 139  0 t = 2
rlabel pdiffusion 301 143 302 144  0 t = 3
rlabel pdiffusion 304 143 305 144  0 t = 4
rlabel pdiffusion 300 138 306 144 0 cell no = 167
<< m1 >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< m2 >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< m2c >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< labels >>
rlabel pdiffusion 85 156 86 157  0 t = 1
rlabel pdiffusion 88 156 89 157  0 t = 2
rlabel pdiffusion 85 161 86 162  0 t = 3
rlabel pdiffusion 88 161 89 162  0 t = 4
rlabel pdiffusion 84 156 90 162 0 cell no = 168
<< m1 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2c >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< labels >>
rlabel pdiffusion 391 192 392 193  0 t = 1
rlabel pdiffusion 394 192 395 193  0 t = 2
rlabel pdiffusion 391 197 392 198  0 t = 3
rlabel pdiffusion 394 197 395 198  0 t = 4
rlabel pdiffusion 390 192 396 198 0 cell no = 169
<< m1 >>
rect 391 192 392 193 
rect 394 192 395 193 
rect 391 197 392 198 
rect 394 197 395 198 
<< m2 >>
rect 391 192 392 193 
rect 394 192 395 193 
rect 391 197 392 198 
rect 394 197 395 198 
<< m2c >>
rect 391 192 392 193 
rect 394 192 395 193 
rect 391 197 392 198 
rect 394 197 395 198 
<< labels >>
rlabel pdiffusion 265 210 266 211  0 t = 1
rlabel pdiffusion 268 210 269 211  0 t = 2
rlabel pdiffusion 265 215 266 216  0 t = 3
rlabel pdiffusion 268 215 269 216  0 t = 4
rlabel pdiffusion 264 210 270 216 0 cell no = 170
<< m1 >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< m2 >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< m2c >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< labels >>
rlabel pdiffusion 247 210 248 211  0 t = 1
rlabel pdiffusion 250 210 251 211  0 t = 2
rlabel pdiffusion 247 215 248 216  0 t = 3
rlabel pdiffusion 250 215 251 216  0 t = 4
rlabel pdiffusion 246 210 252 216 0 cell no = 171
<< m1 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2c >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< labels >>
rlabel pdiffusion 391 102 392 103  0 t = 1
rlabel pdiffusion 394 102 395 103  0 t = 2
rlabel pdiffusion 391 107 392 108  0 t = 3
rlabel pdiffusion 394 107 395 108  0 t = 4
rlabel pdiffusion 390 102 396 108 0 cell no = 172
<< m1 >>
rect 391 102 392 103 
rect 394 102 395 103 
rect 391 107 392 108 
rect 394 107 395 108 
<< m2 >>
rect 391 102 392 103 
rect 394 102 395 103 
rect 391 107 392 108 
rect 394 107 395 108 
<< m2c >>
rect 391 102 392 103 
rect 394 102 395 103 
rect 391 107 392 108 
rect 394 107 395 108 
<< labels >>
rlabel pdiffusion 373 192 374 193  0 t = 1
rlabel pdiffusion 376 192 377 193  0 t = 2
rlabel pdiffusion 373 197 374 198  0 t = 3
rlabel pdiffusion 376 197 377 198  0 t = 4
rlabel pdiffusion 372 192 378 198 0 cell no = 173
<< m1 >>
rect 373 192 374 193 
rect 376 192 377 193 
rect 373 197 374 198 
rect 376 197 377 198 
<< m2 >>
rect 373 192 374 193 
rect 376 192 377 193 
rect 373 197 374 198 
rect 376 197 377 198 
<< m2c >>
rect 373 192 374 193 
rect 376 192 377 193 
rect 373 197 374 198 
rect 376 197 377 198 
<< labels >>
rlabel pdiffusion 301 228 302 229  0 t = 1
rlabel pdiffusion 304 228 305 229  0 t = 2
rlabel pdiffusion 301 233 302 234  0 t = 3
rlabel pdiffusion 304 233 305 234  0 t = 4
rlabel pdiffusion 300 228 306 234 0 cell no = 174
<< m1 >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< m2 >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< m2c >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< labels >>
rlabel pdiffusion 373 156 374 157  0 t = 1
rlabel pdiffusion 376 156 377 157  0 t = 2
rlabel pdiffusion 373 161 374 162  0 t = 3
rlabel pdiffusion 376 161 377 162  0 t = 4
rlabel pdiffusion 372 156 378 162 0 cell no = 175
<< m1 >>
rect 373 156 374 157 
rect 376 156 377 157 
rect 373 161 374 162 
rect 376 161 377 162 
<< m2 >>
rect 373 156 374 157 
rect 376 156 377 157 
rect 373 161 374 162 
rect 376 161 377 162 
<< m2c >>
rect 373 156 374 157 
rect 376 156 377 157 
rect 373 161 374 162 
rect 376 161 377 162 
<< labels >>
rlabel pdiffusion 67 228 68 229  0 t = 1
rlabel pdiffusion 70 228 71 229  0 t = 2
rlabel pdiffusion 67 233 68 234  0 t = 3
rlabel pdiffusion 70 233 71 234  0 t = 4
rlabel pdiffusion 66 228 72 234 0 cell no = 176
<< m1 >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< m2 >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< m2c >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< labels >>
rlabel pdiffusion 265 156 266 157  0 t = 1
rlabel pdiffusion 268 156 269 157  0 t = 2
rlabel pdiffusion 265 161 266 162  0 t = 3
rlabel pdiffusion 268 161 269 162  0 t = 4
rlabel pdiffusion 264 156 270 162 0 cell no = 177
<< m1 >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< m2 >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< m2c >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< labels >>
rlabel pdiffusion 49 138 50 139  0 t = 1
rlabel pdiffusion 52 138 53 139  0 t = 2
rlabel pdiffusion 49 143 50 144  0 t = 3
rlabel pdiffusion 52 143 53 144  0 t = 4
rlabel pdiffusion 48 138 54 144 0 cell no = 178
<< m1 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2c >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< labels >>
rlabel pdiffusion 265 30 266 31  0 t = 1
rlabel pdiffusion 268 30 269 31  0 t = 2
rlabel pdiffusion 265 35 266 36  0 t = 3
rlabel pdiffusion 268 35 269 36  0 t = 4
rlabel pdiffusion 264 30 270 36 0 cell no = 179
<< m1 >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< m2 >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< m2c >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< labels >>
rlabel pdiffusion 229 48 230 49  0 t = 1
rlabel pdiffusion 232 48 233 49  0 t = 2
rlabel pdiffusion 229 53 230 54  0 t = 3
rlabel pdiffusion 232 53 233 54  0 t = 4
rlabel pdiffusion 228 48 234 54 0 cell no = 180
<< m1 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2c >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< labels >>
rlabel pdiffusion 373 246 374 247  0 t = 1
rlabel pdiffusion 376 246 377 247  0 t = 2
rlabel pdiffusion 373 251 374 252  0 t = 3
rlabel pdiffusion 376 251 377 252  0 t = 4
rlabel pdiffusion 372 246 378 252 0 cell no = 181
<< m1 >>
rect 373 246 374 247 
rect 376 246 377 247 
rect 373 251 374 252 
rect 376 251 377 252 
<< m2 >>
rect 373 246 374 247 
rect 376 246 377 247 
rect 373 251 374 252 
rect 376 251 377 252 
<< m2c >>
rect 373 246 374 247 
rect 376 246 377 247 
rect 373 251 374 252 
rect 376 251 377 252 
<< labels >>
rlabel pdiffusion 175 174 176 175  0 t = 1
rlabel pdiffusion 178 174 179 175  0 t = 2
rlabel pdiffusion 175 179 176 180  0 t = 3
rlabel pdiffusion 178 179 179 180  0 t = 4
rlabel pdiffusion 174 174 180 180 0 cell no = 182
<< m1 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2c >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< labels >>
rlabel pdiffusion 139 84 140 85  0 t = 1
rlabel pdiffusion 142 84 143 85  0 t = 2
rlabel pdiffusion 139 89 140 90  0 t = 3
rlabel pdiffusion 142 89 143 90  0 t = 4
rlabel pdiffusion 138 84 144 90 0 cell no = 183
<< m1 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2c >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< labels >>
rlabel pdiffusion 31 228 32 229  0 t = 1
rlabel pdiffusion 34 228 35 229  0 t = 2
rlabel pdiffusion 31 233 32 234  0 t = 3
rlabel pdiffusion 34 233 35 234  0 t = 4
rlabel pdiffusion 30 228 36 234 0 cell no = 184
<< m1 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2c >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< labels >>
rlabel pdiffusion 31 30 32 31  0 t = 1
rlabel pdiffusion 34 30 35 31  0 t = 2
rlabel pdiffusion 31 35 32 36  0 t = 3
rlabel pdiffusion 34 35 35 36  0 t = 4
rlabel pdiffusion 30 30 36 36 0 cell no = 185
<< m1 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2c >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< labels >>
rlabel pdiffusion 427 210 428 211  0 t = 1
rlabel pdiffusion 430 210 431 211  0 t = 2
rlabel pdiffusion 427 215 428 216  0 t = 3
rlabel pdiffusion 430 215 431 216  0 t = 4
rlabel pdiffusion 426 210 432 216 0 cell no = 186
<< m1 >>
rect 427 210 428 211 
rect 430 210 431 211 
rect 427 215 428 216 
rect 430 215 431 216 
<< m2 >>
rect 427 210 428 211 
rect 430 210 431 211 
rect 427 215 428 216 
rect 430 215 431 216 
<< m2c >>
rect 427 210 428 211 
rect 430 210 431 211 
rect 427 215 428 216 
rect 430 215 431 216 
<< labels >>
rlabel pdiffusion 283 336 284 337  0 t = 1
rlabel pdiffusion 286 336 287 337  0 t = 2
rlabel pdiffusion 283 341 284 342  0 t = 3
rlabel pdiffusion 286 341 287 342  0 t = 4
rlabel pdiffusion 282 336 288 342 0 cell no = 187
<< m1 >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< m2 >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< m2c >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< labels >>
rlabel pdiffusion 283 120 284 121  0 t = 1
rlabel pdiffusion 286 120 287 121  0 t = 2
rlabel pdiffusion 283 125 284 126  0 t = 3
rlabel pdiffusion 286 125 287 126  0 t = 4
rlabel pdiffusion 282 120 288 126 0 cell no = 188
<< m1 >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< m2 >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< m2c >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< labels >>
rlabel pdiffusion 409 192 410 193  0 t = 1
rlabel pdiffusion 412 192 413 193  0 t = 2
rlabel pdiffusion 409 197 410 198  0 t = 3
rlabel pdiffusion 412 197 413 198  0 t = 4
rlabel pdiffusion 408 192 414 198 0 cell no = 189
<< m1 >>
rect 409 192 410 193 
rect 412 192 413 193 
rect 409 197 410 198 
rect 412 197 413 198 
<< m2 >>
rect 409 192 410 193 
rect 412 192 413 193 
rect 409 197 410 198 
rect 412 197 413 198 
<< m2c >>
rect 409 192 410 193 
rect 412 192 413 193 
rect 409 197 410 198 
rect 412 197 413 198 
<< labels >>
rlabel pdiffusion 355 264 356 265  0 t = 1
rlabel pdiffusion 358 264 359 265  0 t = 2
rlabel pdiffusion 355 269 356 270  0 t = 3
rlabel pdiffusion 358 269 359 270  0 t = 4
rlabel pdiffusion 354 264 360 270 0 cell no = 190
<< m1 >>
rect 355 264 356 265 
rect 358 264 359 265 
rect 355 269 356 270 
rect 358 269 359 270 
<< m2 >>
rect 355 264 356 265 
rect 358 264 359 265 
rect 355 269 356 270 
rect 358 269 359 270 
<< m2c >>
rect 355 264 356 265 
rect 358 264 359 265 
rect 355 269 356 270 
rect 358 269 359 270 
<< labels >>
rlabel pdiffusion 355 228 356 229  0 t = 1
rlabel pdiffusion 358 228 359 229  0 t = 2
rlabel pdiffusion 355 233 356 234  0 t = 3
rlabel pdiffusion 358 233 359 234  0 t = 4
rlabel pdiffusion 354 228 360 234 0 cell no = 191
<< m1 >>
rect 355 228 356 229 
rect 358 228 359 229 
rect 355 233 356 234 
rect 358 233 359 234 
<< m2 >>
rect 355 228 356 229 
rect 358 228 359 229 
rect 355 233 356 234 
rect 358 233 359 234 
<< m2c >>
rect 355 228 356 229 
rect 358 228 359 229 
rect 355 233 356 234 
rect 358 233 359 234 
<< labels >>
rlabel pdiffusion 193 102 194 103  0 t = 1
rlabel pdiffusion 196 102 197 103  0 t = 2
rlabel pdiffusion 193 107 194 108  0 t = 3
rlabel pdiffusion 196 107 197 108  0 t = 4
rlabel pdiffusion 192 102 198 108 0 cell no = 192
<< m1 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2c >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< labels >>
rlabel pdiffusion 337 12 338 13  0 t = 1
rlabel pdiffusion 340 12 341 13  0 t = 2
rlabel pdiffusion 337 17 338 18  0 t = 3
rlabel pdiffusion 340 17 341 18  0 t = 4
rlabel pdiffusion 336 12 342 18 0 cell no = 193
<< m1 >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< m2 >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< m2c >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< labels >>
rlabel pdiffusion 283 156 284 157  0 t = 1
rlabel pdiffusion 286 156 287 157  0 t = 2
rlabel pdiffusion 283 161 284 162  0 t = 3
rlabel pdiffusion 286 161 287 162  0 t = 4
rlabel pdiffusion 282 156 288 162 0 cell no = 194
<< m1 >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< m2 >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< m2c >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< labels >>
rlabel pdiffusion 427 174 428 175  0 t = 1
rlabel pdiffusion 430 174 431 175  0 t = 2
rlabel pdiffusion 427 179 428 180  0 t = 3
rlabel pdiffusion 430 179 431 180  0 t = 4
rlabel pdiffusion 426 174 432 180 0 cell no = 195
<< m1 >>
rect 427 174 428 175 
rect 430 174 431 175 
rect 427 179 428 180 
rect 430 179 431 180 
<< m2 >>
rect 427 174 428 175 
rect 430 174 431 175 
rect 427 179 428 180 
rect 430 179 431 180 
<< m2c >>
rect 427 174 428 175 
rect 430 174 431 175 
rect 427 179 428 180 
rect 430 179 431 180 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 196
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 373 174 374 175  0 t = 1
rlabel pdiffusion 376 174 377 175  0 t = 2
rlabel pdiffusion 373 179 374 180  0 t = 3
rlabel pdiffusion 376 179 377 180  0 t = 4
rlabel pdiffusion 372 174 378 180 0 cell no = 197
<< m1 >>
rect 373 174 374 175 
rect 376 174 377 175 
rect 373 179 374 180 
rect 376 179 377 180 
<< m2 >>
rect 373 174 374 175 
rect 376 174 377 175 
rect 373 179 374 180 
rect 376 179 377 180 
<< m2c >>
rect 373 174 374 175 
rect 376 174 377 175 
rect 373 179 374 180 
rect 376 179 377 180 
<< labels >>
rlabel pdiffusion 211 336 212 337  0 t = 1
rlabel pdiffusion 214 336 215 337  0 t = 2
rlabel pdiffusion 211 341 212 342  0 t = 3
rlabel pdiffusion 214 341 215 342  0 t = 4
rlabel pdiffusion 210 336 216 342 0 cell no = 198
<< m1 >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< m2 >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< m2c >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< labels >>
rlabel pdiffusion 301 156 302 157  0 t = 1
rlabel pdiffusion 304 156 305 157  0 t = 2
rlabel pdiffusion 301 161 302 162  0 t = 3
rlabel pdiffusion 304 161 305 162  0 t = 4
rlabel pdiffusion 300 156 306 162 0 cell no = 199
<< m1 >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< m2 >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< m2c >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< labels >>
rlabel pdiffusion 193 48 194 49  0 t = 1
rlabel pdiffusion 196 48 197 49  0 t = 2
rlabel pdiffusion 193 53 194 54  0 t = 3
rlabel pdiffusion 196 53 197 54  0 t = 4
rlabel pdiffusion 192 48 198 54 0 cell no = 200
<< m1 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2c >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< labels >>
rlabel pdiffusion 103 228 104 229  0 t = 1
rlabel pdiffusion 106 228 107 229  0 t = 2
rlabel pdiffusion 103 233 104 234  0 t = 3
rlabel pdiffusion 106 233 107 234  0 t = 4
rlabel pdiffusion 102 228 108 234 0 cell no = 201
<< m1 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2c >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< labels >>
rlabel pdiffusion 85 246 86 247  0 t = 1
rlabel pdiffusion 88 246 89 247  0 t = 2
rlabel pdiffusion 85 251 86 252  0 t = 3
rlabel pdiffusion 88 251 89 252  0 t = 4
rlabel pdiffusion 84 246 90 252 0 cell no = 202
<< m1 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2c >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< labels >>
rlabel pdiffusion 49 408 50 409  0 t = 1
rlabel pdiffusion 52 408 53 409  0 t = 2
rlabel pdiffusion 49 413 50 414  0 t = 3
rlabel pdiffusion 52 413 53 414  0 t = 4
rlabel pdiffusion 48 408 54 414 0 cell no = 203
<< m1 >>
rect 49 408 50 409 
rect 52 408 53 409 
rect 49 413 50 414 
rect 52 413 53 414 
<< m2 >>
rect 49 408 50 409 
rect 52 408 53 409 
rect 49 413 50 414 
rect 52 413 53 414 
<< m2c >>
rect 49 408 50 409 
rect 52 408 53 409 
rect 49 413 50 414 
rect 52 413 53 414 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 204
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 247 138 248 139  0 t = 1
rlabel pdiffusion 250 138 251 139  0 t = 2
rlabel pdiffusion 247 143 248 144  0 t = 3
rlabel pdiffusion 250 143 251 144  0 t = 4
rlabel pdiffusion 246 138 252 144 0 cell no = 205
<< m1 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2c >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< labels >>
rlabel pdiffusion 139 444 140 445  0 t = 1
rlabel pdiffusion 142 444 143 445  0 t = 2
rlabel pdiffusion 139 449 140 450  0 t = 3
rlabel pdiffusion 142 449 143 450  0 t = 4
rlabel pdiffusion 138 444 144 450 0 cell no = 206
<< m1 >>
rect 139 444 140 445 
rect 142 444 143 445 
rect 139 449 140 450 
rect 142 449 143 450 
<< m2 >>
rect 139 444 140 445 
rect 142 444 143 445 
rect 139 449 140 450 
rect 142 449 143 450 
<< m2c >>
rect 139 444 140 445 
rect 142 444 143 445 
rect 139 449 140 450 
rect 142 449 143 450 
<< labels >>
rlabel pdiffusion 31 12 32 13  0 t = 1
rlabel pdiffusion 34 12 35 13  0 t = 2
rlabel pdiffusion 31 17 32 18  0 t = 3
rlabel pdiffusion 34 17 35 18  0 t = 4
rlabel pdiffusion 30 12 36 18 0 cell no = 207
<< m1 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2c >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< labels >>
rlabel pdiffusion 157 174 158 175  0 t = 1
rlabel pdiffusion 160 174 161 175  0 t = 2
rlabel pdiffusion 157 179 158 180  0 t = 3
rlabel pdiffusion 160 179 161 180  0 t = 4
rlabel pdiffusion 156 174 162 180 0 cell no = 208
<< m1 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2c >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< labels >>
rlabel pdiffusion 85 264 86 265  0 t = 1
rlabel pdiffusion 88 264 89 265  0 t = 2
rlabel pdiffusion 85 269 86 270  0 t = 3
rlabel pdiffusion 88 269 89 270  0 t = 4
rlabel pdiffusion 84 264 90 270 0 cell no = 209
<< m1 >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< m2 >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< m2c >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< labels >>
rlabel pdiffusion 175 210 176 211  0 t = 1
rlabel pdiffusion 178 210 179 211  0 t = 2
rlabel pdiffusion 175 215 176 216  0 t = 3
rlabel pdiffusion 178 215 179 216  0 t = 4
rlabel pdiffusion 174 210 180 216 0 cell no = 210
<< m1 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2c >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< labels >>
rlabel pdiffusion 121 318 122 319  0 t = 1
rlabel pdiffusion 124 318 125 319  0 t = 2
rlabel pdiffusion 121 323 122 324  0 t = 3
rlabel pdiffusion 124 323 125 324  0 t = 4
rlabel pdiffusion 120 318 126 324 0 cell no = 211
<< m1 >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< m2 >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< m2c >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< labels >>
rlabel pdiffusion 139 174 140 175  0 t = 1
rlabel pdiffusion 142 174 143 175  0 t = 2
rlabel pdiffusion 139 179 140 180  0 t = 3
rlabel pdiffusion 142 179 143 180  0 t = 4
rlabel pdiffusion 138 174 144 180 0 cell no = 212
<< m1 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2c >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< labels >>
rlabel pdiffusion 211 318 212 319  0 t = 1
rlabel pdiffusion 214 318 215 319  0 t = 2
rlabel pdiffusion 211 323 212 324  0 t = 3
rlabel pdiffusion 214 323 215 324  0 t = 4
rlabel pdiffusion 210 318 216 324 0 cell no = 213
<< m1 >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< m2 >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< m2c >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< labels >>
rlabel pdiffusion 229 174 230 175  0 t = 1
rlabel pdiffusion 232 174 233 175  0 t = 2
rlabel pdiffusion 229 179 230 180  0 t = 3
rlabel pdiffusion 232 179 233 180  0 t = 4
rlabel pdiffusion 228 174 234 180 0 cell no = 214
<< m1 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2c >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< labels >>
rlabel pdiffusion 355 84 356 85  0 t = 1
rlabel pdiffusion 358 84 359 85  0 t = 2
rlabel pdiffusion 355 89 356 90  0 t = 3
rlabel pdiffusion 358 89 359 90  0 t = 4
rlabel pdiffusion 354 84 360 90 0 cell no = 215
<< m1 >>
rect 355 84 356 85 
rect 358 84 359 85 
rect 355 89 356 90 
rect 358 89 359 90 
<< m2 >>
rect 355 84 356 85 
rect 358 84 359 85 
rect 355 89 356 90 
rect 358 89 359 90 
<< m2c >>
rect 355 84 356 85 
rect 358 84 359 85 
rect 355 89 356 90 
rect 358 89 359 90 
<< labels >>
rlabel pdiffusion 301 390 302 391  0 t = 1
rlabel pdiffusion 304 390 305 391  0 t = 2
rlabel pdiffusion 301 395 302 396  0 t = 3
rlabel pdiffusion 304 395 305 396  0 t = 4
rlabel pdiffusion 300 390 306 396 0 cell no = 216
<< m1 >>
rect 301 390 302 391 
rect 304 390 305 391 
rect 301 395 302 396 
rect 304 395 305 396 
<< m2 >>
rect 301 390 302 391 
rect 304 390 305 391 
rect 301 395 302 396 
rect 304 395 305 396 
<< m2c >>
rect 301 390 302 391 
rect 304 390 305 391 
rect 301 395 302 396 
rect 304 395 305 396 
<< labels >>
rlabel pdiffusion 319 192 320 193  0 t = 1
rlabel pdiffusion 322 192 323 193  0 t = 2
rlabel pdiffusion 319 197 320 198  0 t = 3
rlabel pdiffusion 322 197 323 198  0 t = 4
rlabel pdiffusion 318 192 324 198 0 cell no = 217
<< m1 >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< m2 >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< m2c >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< labels >>
rlabel pdiffusion 193 12 194 13  0 t = 1
rlabel pdiffusion 196 12 197 13  0 t = 2
rlabel pdiffusion 193 17 194 18  0 t = 3
rlabel pdiffusion 196 17 197 18  0 t = 4
rlabel pdiffusion 192 12 198 18 0 cell no = 218
<< m1 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2c >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< labels >>
rlabel pdiffusion 373 300 374 301  0 t = 1
rlabel pdiffusion 376 300 377 301  0 t = 2
rlabel pdiffusion 373 305 374 306  0 t = 3
rlabel pdiffusion 376 305 377 306  0 t = 4
rlabel pdiffusion 372 300 378 306 0 cell no = 219
<< m1 >>
rect 373 300 374 301 
rect 376 300 377 301 
rect 373 305 374 306 
rect 376 305 377 306 
<< m2 >>
rect 373 300 374 301 
rect 376 300 377 301 
rect 373 305 374 306 
rect 376 305 377 306 
<< m2c >>
rect 373 300 374 301 
rect 376 300 377 301 
rect 373 305 374 306 
rect 376 305 377 306 
<< labels >>
rlabel pdiffusion 445 156 446 157  0 t = 1
rlabel pdiffusion 448 156 449 157  0 t = 2
rlabel pdiffusion 445 161 446 162  0 t = 3
rlabel pdiffusion 448 161 449 162  0 t = 4
rlabel pdiffusion 444 156 450 162 0 cell no = 220
<< m1 >>
rect 445 156 446 157 
rect 448 156 449 157 
rect 445 161 446 162 
rect 448 161 449 162 
<< m2 >>
rect 445 156 446 157 
rect 448 156 449 157 
rect 445 161 446 162 
rect 448 161 449 162 
<< m2c >>
rect 445 156 446 157 
rect 448 156 449 157 
rect 445 161 446 162 
rect 448 161 449 162 
<< labels >>
rlabel pdiffusion 301 12 302 13  0 t = 1
rlabel pdiffusion 304 12 305 13  0 t = 2
rlabel pdiffusion 301 17 302 18  0 t = 3
rlabel pdiffusion 304 17 305 18  0 t = 4
rlabel pdiffusion 300 12 306 18 0 cell no = 221
<< m1 >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< m2 >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< m2c >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< labels >>
rlabel pdiffusion 13 138 14 139  0 t = 1
rlabel pdiffusion 16 138 17 139  0 t = 2
rlabel pdiffusion 13 143 14 144  0 t = 3
rlabel pdiffusion 16 143 17 144  0 t = 4
rlabel pdiffusion 12 138 18 144 0 cell no = 222
<< m1 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2c >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< labels >>
rlabel pdiffusion 283 192 284 193  0 t = 1
rlabel pdiffusion 286 192 287 193  0 t = 2
rlabel pdiffusion 283 197 284 198  0 t = 3
rlabel pdiffusion 286 197 287 198  0 t = 4
rlabel pdiffusion 282 192 288 198 0 cell no = 223
<< m1 >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< m2 >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< m2c >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< labels >>
rlabel pdiffusion 337 102 338 103  0 t = 1
rlabel pdiffusion 340 102 341 103  0 t = 2
rlabel pdiffusion 337 107 338 108  0 t = 3
rlabel pdiffusion 340 107 341 108  0 t = 4
rlabel pdiffusion 336 102 342 108 0 cell no = 224
<< m1 >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< m2 >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< m2c >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< labels >>
rlabel pdiffusion 157 48 158 49  0 t = 1
rlabel pdiffusion 160 48 161 49  0 t = 2
rlabel pdiffusion 157 53 158 54  0 t = 3
rlabel pdiffusion 160 53 161 54  0 t = 4
rlabel pdiffusion 156 48 162 54 0 cell no = 225
<< m1 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2c >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< labels >>
rlabel pdiffusion 31 246 32 247  0 t = 1
rlabel pdiffusion 34 246 35 247  0 t = 2
rlabel pdiffusion 31 251 32 252  0 t = 3
rlabel pdiffusion 34 251 35 252  0 t = 4
rlabel pdiffusion 30 246 36 252 0 cell no = 226
<< m1 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2c >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< labels >>
rlabel pdiffusion 13 210 14 211  0 t = 1
rlabel pdiffusion 16 210 17 211  0 t = 2
rlabel pdiffusion 13 215 14 216  0 t = 3
rlabel pdiffusion 16 215 17 216  0 t = 4
rlabel pdiffusion 12 210 18 216 0 cell no = 227
<< m1 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2c >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 228
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 85 210 86 211  0 t = 1
rlabel pdiffusion 88 210 89 211  0 t = 2
rlabel pdiffusion 85 215 86 216  0 t = 3
rlabel pdiffusion 88 215 89 216  0 t = 4
rlabel pdiffusion 84 210 90 216 0 cell no = 229
<< m1 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2c >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< labels >>
rlabel pdiffusion 85 228 86 229  0 t = 1
rlabel pdiffusion 88 228 89 229  0 t = 2
rlabel pdiffusion 85 233 86 234  0 t = 3
rlabel pdiffusion 88 233 89 234  0 t = 4
rlabel pdiffusion 84 228 90 234 0 cell no = 230
<< m1 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2c >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< labels >>
rlabel pdiffusion 13 120 14 121  0 t = 1
rlabel pdiffusion 16 120 17 121  0 t = 2
rlabel pdiffusion 13 125 14 126  0 t = 3
rlabel pdiffusion 16 125 17 126  0 t = 4
rlabel pdiffusion 12 120 18 126 0 cell no = 231
<< m1 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2c >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< labels >>
rlabel pdiffusion 211 102 212 103  0 t = 1
rlabel pdiffusion 214 102 215 103  0 t = 2
rlabel pdiffusion 211 107 212 108  0 t = 3
rlabel pdiffusion 214 107 215 108  0 t = 4
rlabel pdiffusion 210 102 216 108 0 cell no = 232
<< m1 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2c >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< labels >>
rlabel pdiffusion 409 354 410 355  0 t = 1
rlabel pdiffusion 412 354 413 355  0 t = 2
rlabel pdiffusion 409 359 410 360  0 t = 3
rlabel pdiffusion 412 359 413 360  0 t = 4
rlabel pdiffusion 408 354 414 360 0 cell no = 233
<< m1 >>
rect 409 354 410 355 
rect 412 354 413 355 
rect 409 359 410 360 
rect 412 359 413 360 
<< m2 >>
rect 409 354 410 355 
rect 412 354 413 355 
rect 409 359 410 360 
rect 412 359 413 360 
<< m2c >>
rect 409 354 410 355 
rect 412 354 413 355 
rect 409 359 410 360 
rect 412 359 413 360 
<< labels >>
rlabel pdiffusion 139 48 140 49  0 t = 1
rlabel pdiffusion 142 48 143 49  0 t = 2
rlabel pdiffusion 139 53 140 54  0 t = 3
rlabel pdiffusion 142 53 143 54  0 t = 4
rlabel pdiffusion 138 48 144 54 0 cell no = 234
<< m1 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2c >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< labels >>
rlabel pdiffusion 193 192 194 193  0 t = 1
rlabel pdiffusion 196 192 197 193  0 t = 2
rlabel pdiffusion 193 197 194 198  0 t = 3
rlabel pdiffusion 196 197 197 198  0 t = 4
rlabel pdiffusion 192 192 198 198 0 cell no = 235
<< m1 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2c >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< labels >>
rlabel pdiffusion 229 138 230 139  0 t = 1
rlabel pdiffusion 232 138 233 139  0 t = 2
rlabel pdiffusion 229 143 230 144  0 t = 3
rlabel pdiffusion 232 143 233 144  0 t = 4
rlabel pdiffusion 228 138 234 144 0 cell no = 236
<< m1 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2c >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< labels >>
rlabel pdiffusion 319 246 320 247  0 t = 1
rlabel pdiffusion 322 246 323 247  0 t = 2
rlabel pdiffusion 319 251 320 252  0 t = 3
rlabel pdiffusion 322 251 323 252  0 t = 4
rlabel pdiffusion 318 246 324 252 0 cell no = 237
<< m1 >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< m2 >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< m2c >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< labels >>
rlabel pdiffusion 175 318 176 319  0 t = 1
rlabel pdiffusion 178 318 179 319  0 t = 2
rlabel pdiffusion 175 323 176 324  0 t = 3
rlabel pdiffusion 178 323 179 324  0 t = 4
rlabel pdiffusion 174 318 180 324 0 cell no = 238
<< m1 >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< m2 >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< m2c >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< labels >>
rlabel pdiffusion 283 318 284 319  0 t = 1
rlabel pdiffusion 286 318 287 319  0 t = 2
rlabel pdiffusion 283 323 284 324  0 t = 3
rlabel pdiffusion 286 323 287 324  0 t = 4
rlabel pdiffusion 282 318 288 324 0 cell no = 239
<< m1 >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< m2 >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< m2c >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< labels >>
rlabel pdiffusion 211 192 212 193  0 t = 1
rlabel pdiffusion 214 192 215 193  0 t = 2
rlabel pdiffusion 211 197 212 198  0 t = 3
rlabel pdiffusion 214 197 215 198  0 t = 4
rlabel pdiffusion 210 192 216 198 0 cell no = 240
<< m1 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2c >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< labels >>
rlabel pdiffusion 445 138 446 139  0 t = 1
rlabel pdiffusion 448 138 449 139  0 t = 2
rlabel pdiffusion 445 143 446 144  0 t = 3
rlabel pdiffusion 448 143 449 144  0 t = 4
rlabel pdiffusion 444 138 450 144 0 cell no = 241
<< m1 >>
rect 445 138 446 139 
rect 448 138 449 139 
rect 445 143 446 144 
rect 448 143 449 144 
<< m2 >>
rect 445 138 446 139 
rect 448 138 449 139 
rect 445 143 446 144 
rect 448 143 449 144 
<< m2c >>
rect 445 138 446 139 
rect 448 138 449 139 
rect 445 143 446 144 
rect 448 143 449 144 
<< labels >>
rlabel pdiffusion 391 84 392 85  0 t = 1
rlabel pdiffusion 394 84 395 85  0 t = 2
rlabel pdiffusion 391 89 392 90  0 t = 3
rlabel pdiffusion 394 89 395 90  0 t = 4
rlabel pdiffusion 390 84 396 90 0 cell no = 242
<< m1 >>
rect 391 84 392 85 
rect 394 84 395 85 
rect 391 89 392 90 
rect 394 89 395 90 
<< m2 >>
rect 391 84 392 85 
rect 394 84 395 85 
rect 391 89 392 90 
rect 394 89 395 90 
<< m2c >>
rect 391 84 392 85 
rect 394 84 395 85 
rect 391 89 392 90 
rect 394 89 395 90 
<< labels >>
rlabel pdiffusion 121 336 122 337  0 t = 1
rlabel pdiffusion 124 336 125 337  0 t = 2
rlabel pdiffusion 121 341 122 342  0 t = 3
rlabel pdiffusion 124 341 125 342  0 t = 4
rlabel pdiffusion 120 336 126 342 0 cell no = 243
<< m1 >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< m2 >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< m2c >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< labels >>
rlabel pdiffusion 283 174 284 175  0 t = 1
rlabel pdiffusion 286 174 287 175  0 t = 2
rlabel pdiffusion 283 179 284 180  0 t = 3
rlabel pdiffusion 286 179 287 180  0 t = 4
rlabel pdiffusion 282 174 288 180 0 cell no = 244
<< m1 >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< m2 >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< m2c >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< labels >>
rlabel pdiffusion 427 138 428 139  0 t = 1
rlabel pdiffusion 430 138 431 139  0 t = 2
rlabel pdiffusion 427 143 428 144  0 t = 3
rlabel pdiffusion 430 143 431 144  0 t = 4
rlabel pdiffusion 426 138 432 144 0 cell no = 245
<< m1 >>
rect 427 138 428 139 
rect 430 138 431 139 
rect 427 143 428 144 
rect 430 143 431 144 
<< m2 >>
rect 427 138 428 139 
rect 430 138 431 139 
rect 427 143 428 144 
rect 430 143 431 144 
<< m2c >>
rect 427 138 428 139 
rect 430 138 431 139 
rect 427 143 428 144 
rect 430 143 431 144 
<< labels >>
rlabel pdiffusion 319 156 320 157  0 t = 1
rlabel pdiffusion 322 156 323 157  0 t = 2
rlabel pdiffusion 319 161 320 162  0 t = 3
rlabel pdiffusion 322 161 323 162  0 t = 4
rlabel pdiffusion 318 156 324 162 0 cell no = 246
<< m1 >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< m2 >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< m2c >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< labels >>
rlabel pdiffusion 427 282 428 283  0 t = 1
rlabel pdiffusion 430 282 431 283  0 t = 2
rlabel pdiffusion 427 287 428 288  0 t = 3
rlabel pdiffusion 430 287 431 288  0 t = 4
rlabel pdiffusion 426 282 432 288 0 cell no = 247
<< m1 >>
rect 427 282 428 283 
rect 430 282 431 283 
rect 427 287 428 288 
rect 430 287 431 288 
<< m2 >>
rect 427 282 428 283 
rect 430 282 431 283 
rect 427 287 428 288 
rect 430 287 431 288 
<< m2c >>
rect 427 282 428 283 
rect 430 282 431 283 
rect 427 287 428 288 
rect 430 287 431 288 
<< labels >>
rlabel pdiffusion 355 210 356 211  0 t = 1
rlabel pdiffusion 358 210 359 211  0 t = 2
rlabel pdiffusion 355 215 356 216  0 t = 3
rlabel pdiffusion 358 215 359 216  0 t = 4
rlabel pdiffusion 354 210 360 216 0 cell no = 248
<< m1 >>
rect 355 210 356 211 
rect 358 210 359 211 
rect 355 215 356 216 
rect 358 215 359 216 
<< m2 >>
rect 355 210 356 211 
rect 358 210 359 211 
rect 355 215 356 216 
rect 358 215 359 216 
<< m2c >>
rect 355 210 356 211 
rect 358 210 359 211 
rect 355 215 356 216 
rect 358 215 359 216 
<< labels >>
rlabel pdiffusion 301 444 302 445  0 t = 1
rlabel pdiffusion 304 444 305 445  0 t = 2
rlabel pdiffusion 301 449 302 450  0 t = 3
rlabel pdiffusion 304 449 305 450  0 t = 4
rlabel pdiffusion 300 444 306 450 0 cell no = 249
<< m1 >>
rect 301 444 302 445 
rect 304 444 305 445 
rect 301 449 302 450 
rect 304 449 305 450 
<< m2 >>
rect 301 444 302 445 
rect 304 444 305 445 
rect 301 449 302 450 
rect 304 449 305 450 
<< m2c >>
rect 301 444 302 445 
rect 304 444 305 445 
rect 301 449 302 450 
rect 304 449 305 450 
<< labels >>
rlabel pdiffusion 373 12 374 13  0 t = 1
rlabel pdiffusion 376 12 377 13  0 t = 2
rlabel pdiffusion 373 17 374 18  0 t = 3
rlabel pdiffusion 376 17 377 18  0 t = 4
rlabel pdiffusion 372 12 378 18 0 cell no = 250
<< m1 >>
rect 373 12 374 13 
rect 376 12 377 13 
rect 373 17 374 18 
rect 376 17 377 18 
<< m2 >>
rect 373 12 374 13 
rect 376 12 377 13 
rect 373 17 374 18 
rect 376 17 377 18 
<< m2c >>
rect 373 12 374 13 
rect 376 12 377 13 
rect 373 17 374 18 
rect 376 17 377 18 
<< labels >>
rlabel pdiffusion 13 174 14 175  0 t = 1
rlabel pdiffusion 16 174 17 175  0 t = 2
rlabel pdiffusion 13 179 14 180  0 t = 3
rlabel pdiffusion 16 179 17 180  0 t = 4
rlabel pdiffusion 12 174 18 180 0 cell no = 251
<< m1 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2c >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 252
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 193 210 194 211  0 t = 1
rlabel pdiffusion 196 210 197 211  0 t = 2
rlabel pdiffusion 193 215 194 216  0 t = 3
rlabel pdiffusion 196 215 197 216  0 t = 4
rlabel pdiffusion 192 210 198 216 0 cell no = 253
<< m1 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2c >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< labels >>
rlabel pdiffusion 13 300 14 301  0 t = 1
rlabel pdiffusion 16 300 17 301  0 t = 2
rlabel pdiffusion 13 305 14 306  0 t = 3
rlabel pdiffusion 16 305 17 306  0 t = 4
rlabel pdiffusion 12 300 18 306 0 cell no = 254
<< m1 >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< m2 >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< m2c >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< labels >>
rlabel pdiffusion 31 336 32 337  0 t = 1
rlabel pdiffusion 34 336 35 337  0 t = 2
rlabel pdiffusion 31 341 32 342  0 t = 3
rlabel pdiffusion 34 341 35 342  0 t = 4
rlabel pdiffusion 30 336 36 342 0 cell no = 255
<< m1 >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< m2 >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< m2c >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< labels >>
rlabel pdiffusion 13 156 14 157  0 t = 1
rlabel pdiffusion 16 156 17 157  0 t = 2
rlabel pdiffusion 13 161 14 162  0 t = 3
rlabel pdiffusion 16 161 17 162  0 t = 4
rlabel pdiffusion 12 156 18 162 0 cell no = 256
<< m1 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2c >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 257
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 373 228 374 229  0 t = 1
rlabel pdiffusion 376 228 377 229  0 t = 2
rlabel pdiffusion 373 233 374 234  0 t = 3
rlabel pdiffusion 376 233 377 234  0 t = 4
rlabel pdiffusion 372 228 378 234 0 cell no = 258
<< m1 >>
rect 373 228 374 229 
rect 376 228 377 229 
rect 373 233 374 234 
rect 376 233 377 234 
<< m2 >>
rect 373 228 374 229 
rect 376 228 377 229 
rect 373 233 374 234 
rect 376 233 377 234 
<< m2c >>
rect 373 228 374 229 
rect 376 228 377 229 
rect 373 233 374 234 
rect 376 233 377 234 
<< labels >>
rlabel pdiffusion 103 444 104 445  0 t = 1
rlabel pdiffusion 106 444 107 445  0 t = 2
rlabel pdiffusion 103 449 104 450  0 t = 3
rlabel pdiffusion 106 449 107 450  0 t = 4
rlabel pdiffusion 102 444 108 450 0 cell no = 259
<< m1 >>
rect 103 444 104 445 
rect 106 444 107 445 
rect 103 449 104 450 
rect 106 449 107 450 
<< m2 >>
rect 103 444 104 445 
rect 106 444 107 445 
rect 103 449 104 450 
rect 106 449 107 450 
<< m2c >>
rect 103 444 104 445 
rect 106 444 107 445 
rect 103 449 104 450 
rect 106 449 107 450 
<< labels >>
rlabel pdiffusion 211 30 212 31  0 t = 1
rlabel pdiffusion 214 30 215 31  0 t = 2
rlabel pdiffusion 211 35 212 36  0 t = 3
rlabel pdiffusion 214 35 215 36  0 t = 4
rlabel pdiffusion 210 30 216 36 0 cell no = 260
<< m1 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2c >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< labels >>
rlabel pdiffusion 355 30 356 31  0 t = 1
rlabel pdiffusion 358 30 359 31  0 t = 2
rlabel pdiffusion 355 35 356 36  0 t = 3
rlabel pdiffusion 358 35 359 36  0 t = 4
rlabel pdiffusion 354 30 360 36 0 cell no = 261
<< m1 >>
rect 355 30 356 31 
rect 358 30 359 31 
rect 355 35 356 36 
rect 358 35 359 36 
<< m2 >>
rect 355 30 356 31 
rect 358 30 359 31 
rect 355 35 356 36 
rect 358 35 359 36 
<< m2c >>
rect 355 30 356 31 
rect 358 30 359 31 
rect 355 35 356 36 
rect 358 35 359 36 
<< labels >>
rlabel pdiffusion 193 138 194 139  0 t = 1
rlabel pdiffusion 196 138 197 139  0 t = 2
rlabel pdiffusion 193 143 194 144  0 t = 3
rlabel pdiffusion 196 143 197 144  0 t = 4
rlabel pdiffusion 192 138 198 144 0 cell no = 262
<< m1 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2c >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< labels >>
rlabel pdiffusion 229 102 230 103  0 t = 1
rlabel pdiffusion 232 102 233 103  0 t = 2
rlabel pdiffusion 229 107 230 108  0 t = 3
rlabel pdiffusion 232 107 233 108  0 t = 4
rlabel pdiffusion 228 102 234 108 0 cell no = 263
<< m1 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2c >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< labels >>
rlabel pdiffusion 229 246 230 247  0 t = 1
rlabel pdiffusion 232 246 233 247  0 t = 2
rlabel pdiffusion 229 251 230 252  0 t = 3
rlabel pdiffusion 232 251 233 252  0 t = 4
rlabel pdiffusion 228 246 234 252 0 cell no = 264
<< m1 >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< m2 >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< m2c >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< labels >>
rlabel pdiffusion 337 264 338 265  0 t = 1
rlabel pdiffusion 340 264 341 265  0 t = 2
rlabel pdiffusion 337 269 338 270  0 t = 3
rlabel pdiffusion 340 269 341 270  0 t = 4
rlabel pdiffusion 336 264 342 270 0 cell no = 265
<< m1 >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< m2 >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< m2c >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< labels >>
rlabel pdiffusion 139 246 140 247  0 t = 1
rlabel pdiffusion 142 246 143 247  0 t = 2
rlabel pdiffusion 139 251 140 252  0 t = 3
rlabel pdiffusion 142 251 143 252  0 t = 4
rlabel pdiffusion 138 246 144 252 0 cell no = 266
<< m1 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2c >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< labels >>
rlabel pdiffusion 265 66 266 67  0 t = 1
rlabel pdiffusion 268 66 269 67  0 t = 2
rlabel pdiffusion 265 71 266 72  0 t = 3
rlabel pdiffusion 268 71 269 72  0 t = 4
rlabel pdiffusion 264 66 270 72 0 cell no = 267
<< m1 >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< m2 >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< m2c >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< labels >>
rlabel pdiffusion 283 246 284 247  0 t = 1
rlabel pdiffusion 286 246 287 247  0 t = 2
rlabel pdiffusion 283 251 284 252  0 t = 3
rlabel pdiffusion 286 251 287 252  0 t = 4
rlabel pdiffusion 282 246 288 252 0 cell no = 268
<< m1 >>
rect 283 246 284 247 
rect 286 246 287 247 
rect 283 251 284 252 
rect 286 251 287 252 
<< m2 >>
rect 283 246 284 247 
rect 286 246 287 247 
rect 283 251 284 252 
rect 286 251 287 252 
<< m2c >>
rect 283 246 284 247 
rect 286 246 287 247 
rect 283 251 284 252 
rect 286 251 287 252 
<< labels >>
rlabel pdiffusion 409 156 410 157  0 t = 1
rlabel pdiffusion 412 156 413 157  0 t = 2
rlabel pdiffusion 409 161 410 162  0 t = 3
rlabel pdiffusion 412 161 413 162  0 t = 4
rlabel pdiffusion 408 156 414 162 0 cell no = 269
<< m1 >>
rect 409 156 410 157 
rect 412 156 413 157 
rect 409 161 410 162 
rect 412 161 413 162 
<< m2 >>
rect 409 156 410 157 
rect 412 156 413 157 
rect 409 161 410 162 
rect 412 161 413 162 
<< m2c >>
rect 409 156 410 157 
rect 412 156 413 157 
rect 409 161 410 162 
rect 412 161 413 162 
<< labels >>
rlabel pdiffusion 67 444 68 445  0 t = 1
rlabel pdiffusion 70 444 71 445  0 t = 2
rlabel pdiffusion 67 449 68 450  0 t = 3
rlabel pdiffusion 70 449 71 450  0 t = 4
rlabel pdiffusion 66 444 72 450 0 cell no = 270
<< m1 >>
rect 67 444 68 445 
rect 70 444 71 445 
rect 67 449 68 450 
rect 70 449 71 450 
<< m2 >>
rect 67 444 68 445 
rect 70 444 71 445 
rect 67 449 68 450 
rect 70 449 71 450 
<< m2c >>
rect 67 444 68 445 
rect 70 444 71 445 
rect 67 449 68 450 
rect 70 449 71 450 
<< labels >>
rlabel pdiffusion 193 84 194 85  0 t = 1
rlabel pdiffusion 196 84 197 85  0 t = 2
rlabel pdiffusion 193 89 194 90  0 t = 3
rlabel pdiffusion 196 89 197 90  0 t = 4
rlabel pdiffusion 192 84 198 90 0 cell no = 271
<< m1 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2c >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< labels >>
rlabel pdiffusion 283 12 284 13  0 t = 1
rlabel pdiffusion 286 12 287 13  0 t = 2
rlabel pdiffusion 283 17 284 18  0 t = 3
rlabel pdiffusion 286 17 287 18  0 t = 4
rlabel pdiffusion 282 12 288 18 0 cell no = 272
<< m1 >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< m2 >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< m2c >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< labels >>
rlabel pdiffusion 229 228 230 229  0 t = 1
rlabel pdiffusion 232 228 233 229  0 t = 2
rlabel pdiffusion 229 233 230 234  0 t = 3
rlabel pdiffusion 232 233 233 234  0 t = 4
rlabel pdiffusion 228 228 234 234 0 cell no = 273
<< m1 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2c >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< labels >>
rlabel pdiffusion 121 156 122 157  0 t = 1
rlabel pdiffusion 124 156 125 157  0 t = 2
rlabel pdiffusion 121 161 122 162  0 t = 3
rlabel pdiffusion 124 161 125 162  0 t = 4
rlabel pdiffusion 120 156 126 162 0 cell no = 274
<< m1 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2c >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< labels >>
rlabel pdiffusion 445 408 446 409  0 t = 1
rlabel pdiffusion 448 408 449 409  0 t = 2
rlabel pdiffusion 445 413 446 414  0 t = 3
rlabel pdiffusion 448 413 449 414  0 t = 4
rlabel pdiffusion 444 408 450 414 0 cell no = 275
<< m1 >>
rect 445 408 446 409 
rect 448 408 449 409 
rect 445 413 446 414 
rect 448 413 449 414 
<< m2 >>
rect 445 408 446 409 
rect 448 408 449 409 
rect 445 413 446 414 
rect 448 413 449 414 
<< m2c >>
rect 445 408 446 409 
rect 448 408 449 409 
rect 445 413 446 414 
rect 448 413 449 414 
<< labels >>
rlabel pdiffusion 103 264 104 265  0 t = 1
rlabel pdiffusion 106 264 107 265  0 t = 2
rlabel pdiffusion 103 269 104 270  0 t = 3
rlabel pdiffusion 106 269 107 270  0 t = 4
rlabel pdiffusion 102 264 108 270 0 cell no = 276
<< m1 >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< m2 >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< m2c >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< labels >>
rlabel pdiffusion 319 138 320 139  0 t = 1
rlabel pdiffusion 322 138 323 139  0 t = 2
rlabel pdiffusion 319 143 320 144  0 t = 3
rlabel pdiffusion 322 143 323 144  0 t = 4
rlabel pdiffusion 318 138 324 144 0 cell no = 277
<< m1 >>
rect 319 138 320 139 
rect 322 138 323 139 
rect 319 143 320 144 
rect 322 143 323 144 
<< m2 >>
rect 319 138 320 139 
rect 322 138 323 139 
rect 319 143 320 144 
rect 322 143 323 144 
<< m2c >>
rect 319 138 320 139 
rect 322 138 323 139 
rect 319 143 320 144 
rect 322 143 323 144 
<< labels >>
rlabel pdiffusion 175 48 176 49  0 t = 1
rlabel pdiffusion 178 48 179 49  0 t = 2
rlabel pdiffusion 175 53 176 54  0 t = 3
rlabel pdiffusion 178 53 179 54  0 t = 4
rlabel pdiffusion 174 48 180 54 0 cell no = 278
<< m1 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2c >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< labels >>
rlabel pdiffusion 67 192 68 193  0 t = 1
rlabel pdiffusion 70 192 71 193  0 t = 2
rlabel pdiffusion 67 197 68 198  0 t = 3
rlabel pdiffusion 70 197 71 198  0 t = 4
rlabel pdiffusion 66 192 72 198 0 cell no = 279
<< m1 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2c >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< labels >>
rlabel pdiffusion 121 228 122 229  0 t = 1
rlabel pdiffusion 124 228 125 229  0 t = 2
rlabel pdiffusion 121 233 122 234  0 t = 3
rlabel pdiffusion 124 233 125 234  0 t = 4
rlabel pdiffusion 120 228 126 234 0 cell no = 280
<< m1 >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< m2 >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< m2c >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< labels >>
rlabel pdiffusion 157 408 158 409  0 t = 1
rlabel pdiffusion 160 408 161 409  0 t = 2
rlabel pdiffusion 157 413 158 414  0 t = 3
rlabel pdiffusion 160 413 161 414  0 t = 4
rlabel pdiffusion 156 408 162 414 0 cell no = 281
<< m1 >>
rect 157 408 158 409 
rect 160 408 161 409 
rect 157 413 158 414 
rect 160 413 161 414 
<< m2 >>
rect 157 408 158 409 
rect 160 408 161 409 
rect 157 413 158 414 
rect 160 413 161 414 
<< m2c >>
rect 157 408 158 409 
rect 160 408 161 409 
rect 157 413 158 414 
rect 160 413 161 414 
<< labels >>
rlabel pdiffusion 157 210 158 211  0 t = 1
rlabel pdiffusion 160 210 161 211  0 t = 2
rlabel pdiffusion 157 215 158 216  0 t = 3
rlabel pdiffusion 160 215 161 216  0 t = 4
rlabel pdiffusion 156 210 162 216 0 cell no = 282
<< m1 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2c >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< labels >>
rlabel pdiffusion 193 426 194 427  0 t = 1
rlabel pdiffusion 196 426 197 427  0 t = 2
rlabel pdiffusion 193 431 194 432  0 t = 3
rlabel pdiffusion 196 431 197 432  0 t = 4
rlabel pdiffusion 192 426 198 432 0 cell no = 283
<< m1 >>
rect 193 426 194 427 
rect 196 426 197 427 
rect 193 431 194 432 
rect 196 431 197 432 
<< m2 >>
rect 193 426 194 427 
rect 196 426 197 427 
rect 193 431 194 432 
rect 196 431 197 432 
<< m2c >>
rect 193 426 194 427 
rect 196 426 197 427 
rect 193 431 194 432 
rect 196 431 197 432 
<< labels >>
rlabel pdiffusion 229 282 230 283  0 t = 1
rlabel pdiffusion 232 282 233 283  0 t = 2
rlabel pdiffusion 229 287 230 288  0 t = 3
rlabel pdiffusion 232 287 233 288  0 t = 4
rlabel pdiffusion 228 282 234 288 0 cell no = 284
<< m1 >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< m2 >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< m2c >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< labels >>
rlabel pdiffusion 229 426 230 427  0 t = 1
rlabel pdiffusion 232 426 233 427  0 t = 2
rlabel pdiffusion 229 431 230 432  0 t = 3
rlabel pdiffusion 232 431 233 432  0 t = 4
rlabel pdiffusion 228 426 234 432 0 cell no = 285
<< m1 >>
rect 229 426 230 427 
rect 232 426 233 427 
rect 229 431 230 432 
rect 232 431 233 432 
<< m2 >>
rect 229 426 230 427 
rect 232 426 233 427 
rect 229 431 230 432 
rect 232 431 233 432 
<< m2c >>
rect 229 426 230 427 
rect 232 426 233 427 
rect 229 431 230 432 
rect 232 431 233 432 
<< labels >>
rlabel pdiffusion 121 246 122 247  0 t = 1
rlabel pdiffusion 124 246 125 247  0 t = 2
rlabel pdiffusion 121 251 122 252  0 t = 3
rlabel pdiffusion 124 251 125 252  0 t = 4
rlabel pdiffusion 120 246 126 252 0 cell no = 286
<< m1 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2c >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< labels >>
rlabel pdiffusion 373 210 374 211  0 t = 1
rlabel pdiffusion 376 210 377 211  0 t = 2
rlabel pdiffusion 373 215 374 216  0 t = 3
rlabel pdiffusion 376 215 377 216  0 t = 4
rlabel pdiffusion 372 210 378 216 0 cell no = 287
<< m1 >>
rect 373 210 374 211 
rect 376 210 377 211 
rect 373 215 374 216 
rect 376 215 377 216 
<< m2 >>
rect 373 210 374 211 
rect 376 210 377 211 
rect 373 215 374 216 
rect 376 215 377 216 
<< m2c >>
rect 373 210 374 211 
rect 376 210 377 211 
rect 373 215 374 216 
rect 376 215 377 216 
<< labels >>
rlabel pdiffusion 445 246 446 247  0 t = 1
rlabel pdiffusion 448 246 449 247  0 t = 2
rlabel pdiffusion 445 251 446 252  0 t = 3
rlabel pdiffusion 448 251 449 252  0 t = 4
rlabel pdiffusion 444 246 450 252 0 cell no = 288
<< m1 >>
rect 445 246 446 247 
rect 448 246 449 247 
rect 445 251 446 252 
rect 448 251 449 252 
<< m2 >>
rect 445 246 446 247 
rect 448 246 449 247 
rect 445 251 446 252 
rect 448 251 449 252 
<< m2c >>
rect 445 246 446 247 
rect 448 246 449 247 
rect 445 251 446 252 
rect 448 251 449 252 
<< labels >>
rlabel pdiffusion 157 192 158 193  0 t = 1
rlabel pdiffusion 160 192 161 193  0 t = 2
rlabel pdiffusion 157 197 158 198  0 t = 3
rlabel pdiffusion 160 197 161 198  0 t = 4
rlabel pdiffusion 156 192 162 198 0 cell no = 289
<< m1 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2c >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< labels >>
rlabel pdiffusion 337 426 338 427  0 t = 1
rlabel pdiffusion 340 426 341 427  0 t = 2
rlabel pdiffusion 337 431 338 432  0 t = 3
rlabel pdiffusion 340 431 341 432  0 t = 4
rlabel pdiffusion 336 426 342 432 0 cell no = 290
<< m1 >>
rect 337 426 338 427 
rect 340 426 341 427 
rect 337 431 338 432 
rect 340 431 341 432 
<< m2 >>
rect 337 426 338 427 
rect 340 426 341 427 
rect 337 431 338 432 
rect 340 431 341 432 
<< m2c >>
rect 337 426 338 427 
rect 340 426 341 427 
rect 337 431 338 432 
rect 340 431 341 432 
<< labels >>
rlabel pdiffusion 319 318 320 319  0 t = 1
rlabel pdiffusion 322 318 323 319  0 t = 2
rlabel pdiffusion 319 323 320 324  0 t = 3
rlabel pdiffusion 322 323 323 324  0 t = 4
rlabel pdiffusion 318 318 324 324 0 cell no = 291
<< m1 >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< m2 >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< m2c >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 292
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 409 174 410 175  0 t = 1
rlabel pdiffusion 412 174 413 175  0 t = 2
rlabel pdiffusion 409 179 410 180  0 t = 3
rlabel pdiffusion 412 179 413 180  0 t = 4
rlabel pdiffusion 408 174 414 180 0 cell no = 293
<< m1 >>
rect 409 174 410 175 
rect 412 174 413 175 
rect 409 179 410 180 
rect 412 179 413 180 
<< m2 >>
rect 409 174 410 175 
rect 412 174 413 175 
rect 409 179 410 180 
rect 412 179 413 180 
<< m2c >>
rect 409 174 410 175 
rect 412 174 413 175 
rect 409 179 410 180 
rect 412 179 413 180 
<< labels >>
rlabel pdiffusion 427 246 428 247  0 t = 1
rlabel pdiffusion 430 246 431 247  0 t = 2
rlabel pdiffusion 427 251 428 252  0 t = 3
rlabel pdiffusion 430 251 431 252  0 t = 4
rlabel pdiffusion 426 246 432 252 0 cell no = 294
<< m1 >>
rect 427 246 428 247 
rect 430 246 431 247 
rect 427 251 428 252 
rect 430 251 431 252 
<< m2 >>
rect 427 246 428 247 
rect 430 246 431 247 
rect 427 251 428 252 
rect 430 251 431 252 
<< m2c >>
rect 427 246 428 247 
rect 430 246 431 247 
rect 427 251 428 252 
rect 430 251 431 252 
<< labels >>
rlabel pdiffusion 265 48 266 49  0 t = 1
rlabel pdiffusion 268 48 269 49  0 t = 2
rlabel pdiffusion 265 53 266 54  0 t = 3
rlabel pdiffusion 268 53 269 54  0 t = 4
rlabel pdiffusion 264 48 270 54 0 cell no = 295
<< m1 >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< m2 >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< m2c >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< labels >>
rlabel pdiffusion 247 390 248 391  0 t = 1
rlabel pdiffusion 250 390 251 391  0 t = 2
rlabel pdiffusion 247 395 248 396  0 t = 3
rlabel pdiffusion 250 395 251 396  0 t = 4
rlabel pdiffusion 246 390 252 396 0 cell no = 296
<< m1 >>
rect 247 390 248 391 
rect 250 390 251 391 
rect 247 395 248 396 
rect 250 395 251 396 
<< m2 >>
rect 247 390 248 391 
rect 250 390 251 391 
rect 247 395 248 396 
rect 250 395 251 396 
<< m2c >>
rect 247 390 248 391 
rect 250 390 251 391 
rect 247 395 248 396 
rect 250 395 251 396 
<< labels >>
rlabel pdiffusion 157 120 158 121  0 t = 1
rlabel pdiffusion 160 120 161 121  0 t = 2
rlabel pdiffusion 157 125 158 126  0 t = 3
rlabel pdiffusion 160 125 161 126  0 t = 4
rlabel pdiffusion 156 120 162 126 0 cell no = 297
<< m1 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2c >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< labels >>
rlabel pdiffusion 13 192 14 193  0 t = 1
rlabel pdiffusion 16 192 17 193  0 t = 2
rlabel pdiffusion 13 197 14 198  0 t = 3
rlabel pdiffusion 16 197 17 198  0 t = 4
rlabel pdiffusion 12 192 18 198 0 cell no = 298
<< m1 >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< m2 >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< m2c >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< labels >>
rlabel pdiffusion 121 210 122 211  0 t = 1
rlabel pdiffusion 124 210 125 211  0 t = 2
rlabel pdiffusion 121 215 122 216  0 t = 3
rlabel pdiffusion 124 215 125 216  0 t = 4
rlabel pdiffusion 120 210 126 216 0 cell no = 299
<< m1 >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< m2 >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< m2c >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< labels >>
rlabel pdiffusion 265 174 266 175  0 t = 1
rlabel pdiffusion 268 174 269 175  0 t = 2
rlabel pdiffusion 265 179 266 180  0 t = 3
rlabel pdiffusion 268 179 269 180  0 t = 4
rlabel pdiffusion 264 174 270 180 0 cell no = 300
<< m1 >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< m2 >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< m2c >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 301
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 175 30 176 31  0 t = 1
rlabel pdiffusion 178 30 179 31  0 t = 2
rlabel pdiffusion 175 35 176 36  0 t = 3
rlabel pdiffusion 178 35 179 36  0 t = 4
rlabel pdiffusion 174 30 180 36 0 cell no = 302
<< m1 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2c >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< labels >>
rlabel pdiffusion 49 228 50 229  0 t = 1
rlabel pdiffusion 52 228 53 229  0 t = 2
rlabel pdiffusion 49 233 50 234  0 t = 3
rlabel pdiffusion 52 233 53 234  0 t = 4
rlabel pdiffusion 48 228 54 234 0 cell no = 303
<< m1 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2c >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< labels >>
rlabel pdiffusion 139 102 140 103  0 t = 1
rlabel pdiffusion 142 102 143 103  0 t = 2
rlabel pdiffusion 139 107 140 108  0 t = 3
rlabel pdiffusion 142 107 143 108  0 t = 4
rlabel pdiffusion 138 102 144 108 0 cell no = 304
<< m1 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2c >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< labels >>
rlabel pdiffusion 301 336 302 337  0 t = 1
rlabel pdiffusion 304 336 305 337  0 t = 2
rlabel pdiffusion 301 341 302 342  0 t = 3
rlabel pdiffusion 304 341 305 342  0 t = 4
rlabel pdiffusion 300 336 306 342 0 cell no = 305
<< m1 >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< m2 >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< m2c >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< labels >>
rlabel pdiffusion 67 174 68 175  0 t = 1
rlabel pdiffusion 70 174 71 175  0 t = 2
rlabel pdiffusion 67 179 68 180  0 t = 3
rlabel pdiffusion 70 179 71 180  0 t = 4
rlabel pdiffusion 66 174 72 180 0 cell no = 306
<< m1 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2c >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< labels >>
rlabel pdiffusion 103 192 104 193  0 t = 1
rlabel pdiffusion 106 192 107 193  0 t = 2
rlabel pdiffusion 103 197 104 198  0 t = 3
rlabel pdiffusion 106 197 107 198  0 t = 4
rlabel pdiffusion 102 192 108 198 0 cell no = 307
<< m1 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2c >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< labels >>
rlabel pdiffusion 85 192 86 193  0 t = 1
rlabel pdiffusion 88 192 89 193  0 t = 2
rlabel pdiffusion 85 197 86 198  0 t = 3
rlabel pdiffusion 88 197 89 198  0 t = 4
rlabel pdiffusion 84 192 90 198 0 cell no = 308
<< m1 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2c >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< labels >>
rlabel pdiffusion 355 174 356 175  0 t = 1
rlabel pdiffusion 358 174 359 175  0 t = 2
rlabel pdiffusion 355 179 356 180  0 t = 3
rlabel pdiffusion 358 179 359 180  0 t = 4
rlabel pdiffusion 354 174 360 180 0 cell no = 309
<< m1 >>
rect 355 174 356 175 
rect 358 174 359 175 
rect 355 179 356 180 
rect 358 179 359 180 
<< m2 >>
rect 355 174 356 175 
rect 358 174 359 175 
rect 355 179 356 180 
rect 358 179 359 180 
<< m2c >>
rect 355 174 356 175 
rect 358 174 359 175 
rect 355 179 356 180 
rect 358 179 359 180 
<< labels >>
rlabel pdiffusion 175 228 176 229  0 t = 1
rlabel pdiffusion 178 228 179 229  0 t = 2
rlabel pdiffusion 175 233 176 234  0 t = 3
rlabel pdiffusion 178 233 179 234  0 t = 4
rlabel pdiffusion 174 228 180 234 0 cell no = 310
<< m1 >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< m2 >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< m2c >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< labels >>
rlabel pdiffusion 247 372 248 373  0 t = 1
rlabel pdiffusion 250 372 251 373  0 t = 2
rlabel pdiffusion 247 377 248 378  0 t = 3
rlabel pdiffusion 250 377 251 378  0 t = 4
rlabel pdiffusion 246 372 252 378 0 cell no = 311
<< m1 >>
rect 247 372 248 373 
rect 250 372 251 373 
rect 247 377 248 378 
rect 250 377 251 378 
<< m2 >>
rect 247 372 248 373 
rect 250 372 251 373 
rect 247 377 248 378 
rect 250 377 251 378 
<< m2c >>
rect 247 372 248 373 
rect 250 372 251 373 
rect 247 377 248 378 
rect 250 377 251 378 
<< labels >>
rlabel pdiffusion 49 264 50 265  0 t = 1
rlabel pdiffusion 52 264 53 265  0 t = 2
rlabel pdiffusion 49 269 50 270  0 t = 3
rlabel pdiffusion 52 269 53 270  0 t = 4
rlabel pdiffusion 48 264 54 270 0 cell no = 312
<< m1 >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< m2 >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< m2c >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< labels >>
rlabel pdiffusion 445 192 446 193  0 t = 1
rlabel pdiffusion 448 192 449 193  0 t = 2
rlabel pdiffusion 445 197 446 198  0 t = 3
rlabel pdiffusion 448 197 449 198  0 t = 4
rlabel pdiffusion 444 192 450 198 0 cell no = 313
<< m1 >>
rect 445 192 446 193 
rect 448 192 449 193 
rect 445 197 446 198 
rect 448 197 449 198 
<< m2 >>
rect 445 192 446 193 
rect 448 192 449 193 
rect 445 197 446 198 
rect 448 197 449 198 
<< m2c >>
rect 445 192 446 193 
rect 448 192 449 193 
rect 445 197 446 198 
rect 448 197 449 198 
<< labels >>
rlabel pdiffusion 409 246 410 247  0 t = 1
rlabel pdiffusion 412 246 413 247  0 t = 2
rlabel pdiffusion 409 251 410 252  0 t = 3
rlabel pdiffusion 412 251 413 252  0 t = 4
rlabel pdiffusion 408 246 414 252 0 cell no = 314
<< m1 >>
rect 409 246 410 247 
rect 412 246 413 247 
rect 409 251 410 252 
rect 412 251 413 252 
<< m2 >>
rect 409 246 410 247 
rect 412 246 413 247 
rect 409 251 410 252 
rect 412 251 413 252 
<< m2c >>
rect 409 246 410 247 
rect 412 246 413 247 
rect 409 251 410 252 
rect 412 251 413 252 
<< labels >>
rlabel pdiffusion 247 30 248 31  0 t = 1
rlabel pdiffusion 250 30 251 31  0 t = 2
rlabel pdiffusion 247 35 248 36  0 t = 3
rlabel pdiffusion 250 35 251 36  0 t = 4
rlabel pdiffusion 246 30 252 36 0 cell no = 315
<< m1 >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< m2 >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< m2c >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< labels >>
rlabel pdiffusion 13 246 14 247  0 t = 1
rlabel pdiffusion 16 246 17 247  0 t = 2
rlabel pdiffusion 13 251 14 252  0 t = 3
rlabel pdiffusion 16 251 17 252  0 t = 4
rlabel pdiffusion 12 246 18 252 0 cell no = 316
<< m1 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2c >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< labels >>
rlabel pdiffusion 247 84 248 85  0 t = 1
rlabel pdiffusion 250 84 251 85  0 t = 2
rlabel pdiffusion 247 89 248 90  0 t = 3
rlabel pdiffusion 250 89 251 90  0 t = 4
rlabel pdiffusion 246 84 252 90 0 cell no = 317
<< m1 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2c >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< labels >>
rlabel pdiffusion 445 48 446 49  0 t = 1
rlabel pdiffusion 448 48 449 49  0 t = 2
rlabel pdiffusion 445 53 446 54  0 t = 3
rlabel pdiffusion 448 53 449 54  0 t = 4
rlabel pdiffusion 444 48 450 54 0 cell no = 318
<< m1 >>
rect 445 48 446 49 
rect 448 48 449 49 
rect 445 53 446 54 
rect 448 53 449 54 
<< m2 >>
rect 445 48 446 49 
rect 448 48 449 49 
rect 445 53 446 54 
rect 448 53 449 54 
<< m2c >>
rect 445 48 446 49 
rect 448 48 449 49 
rect 445 53 446 54 
rect 448 53 449 54 
<< labels >>
rlabel pdiffusion 103 390 104 391  0 t = 1
rlabel pdiffusion 106 390 107 391  0 t = 2
rlabel pdiffusion 103 395 104 396  0 t = 3
rlabel pdiffusion 106 395 107 396  0 t = 4
rlabel pdiffusion 102 390 108 396 0 cell no = 319
<< m1 >>
rect 103 390 104 391 
rect 106 390 107 391 
rect 103 395 104 396 
rect 106 395 107 396 
<< m2 >>
rect 103 390 104 391 
rect 106 390 107 391 
rect 103 395 104 396 
rect 106 395 107 396 
<< m2c >>
rect 103 390 104 391 
rect 106 390 107 391 
rect 103 395 104 396 
rect 106 395 107 396 
<< labels >>
rlabel pdiffusion 427 264 428 265  0 t = 1
rlabel pdiffusion 430 264 431 265  0 t = 2
rlabel pdiffusion 427 269 428 270  0 t = 3
rlabel pdiffusion 430 269 431 270  0 t = 4
rlabel pdiffusion 426 264 432 270 0 cell no = 320
<< m1 >>
rect 427 264 428 265 
rect 430 264 431 265 
rect 427 269 428 270 
rect 430 269 431 270 
<< m2 >>
rect 427 264 428 265 
rect 430 264 431 265 
rect 427 269 428 270 
rect 430 269 431 270 
<< m2c >>
rect 427 264 428 265 
rect 430 264 431 265 
rect 427 269 428 270 
rect 430 269 431 270 
<< labels >>
rlabel pdiffusion 391 264 392 265  0 t = 1
rlabel pdiffusion 394 264 395 265  0 t = 2
rlabel pdiffusion 391 269 392 270  0 t = 3
rlabel pdiffusion 394 269 395 270  0 t = 4
rlabel pdiffusion 390 264 396 270 0 cell no = 321
<< m1 >>
rect 391 264 392 265 
rect 394 264 395 265 
rect 391 269 392 270 
rect 394 269 395 270 
<< m2 >>
rect 391 264 392 265 
rect 394 264 395 265 
rect 391 269 392 270 
rect 394 269 395 270 
<< m2c >>
rect 391 264 392 265 
rect 394 264 395 265 
rect 391 269 392 270 
rect 394 269 395 270 
<< labels >>
rlabel pdiffusion 445 282 446 283  0 t = 1
rlabel pdiffusion 448 282 449 283  0 t = 2
rlabel pdiffusion 445 287 446 288  0 t = 3
rlabel pdiffusion 448 287 449 288  0 t = 4
rlabel pdiffusion 444 282 450 288 0 cell no = 322
<< m1 >>
rect 445 282 446 283 
rect 448 282 449 283 
rect 445 287 446 288 
rect 448 287 449 288 
<< m2 >>
rect 445 282 446 283 
rect 448 282 449 283 
rect 445 287 446 288 
rect 448 287 449 288 
<< m2c >>
rect 445 282 446 283 
rect 448 282 449 283 
rect 445 287 446 288 
rect 448 287 449 288 
<< labels >>
rlabel pdiffusion 445 264 446 265  0 t = 1
rlabel pdiffusion 448 264 449 265  0 t = 2
rlabel pdiffusion 445 269 446 270  0 t = 3
rlabel pdiffusion 448 269 449 270  0 t = 4
rlabel pdiffusion 444 264 450 270 0 cell no = 323
<< m1 >>
rect 445 264 446 265 
rect 448 264 449 265 
rect 445 269 446 270 
rect 448 269 449 270 
<< m2 >>
rect 445 264 446 265 
rect 448 264 449 265 
rect 445 269 446 270 
rect 448 269 449 270 
<< m2c >>
rect 445 264 446 265 
rect 448 264 449 265 
rect 445 269 446 270 
rect 448 269 449 270 
<< labels >>
rlabel pdiffusion 337 372 338 373  0 t = 1
rlabel pdiffusion 340 372 341 373  0 t = 2
rlabel pdiffusion 337 377 338 378  0 t = 3
rlabel pdiffusion 340 377 341 378  0 t = 4
rlabel pdiffusion 336 372 342 378 0 cell no = 324
<< m1 >>
rect 337 372 338 373 
rect 340 372 341 373 
rect 337 377 338 378 
rect 340 377 341 378 
<< m2 >>
rect 337 372 338 373 
rect 340 372 341 373 
rect 337 377 338 378 
rect 340 377 341 378 
<< m2c >>
rect 337 372 338 373 
rect 340 372 341 373 
rect 337 377 338 378 
rect 340 377 341 378 
<< labels >>
rlabel pdiffusion 373 120 374 121  0 t = 1
rlabel pdiffusion 376 120 377 121  0 t = 2
rlabel pdiffusion 373 125 374 126  0 t = 3
rlabel pdiffusion 376 125 377 126  0 t = 4
rlabel pdiffusion 372 120 378 126 0 cell no = 325
<< m1 >>
rect 373 120 374 121 
rect 376 120 377 121 
rect 373 125 374 126 
rect 376 125 377 126 
<< m2 >>
rect 373 120 374 121 
rect 376 120 377 121 
rect 373 125 374 126 
rect 376 125 377 126 
<< m2c >>
rect 373 120 374 121 
rect 376 120 377 121 
rect 373 125 374 126 
rect 376 125 377 126 
<< labels >>
rlabel pdiffusion 121 282 122 283  0 t = 1
rlabel pdiffusion 124 282 125 283  0 t = 2
rlabel pdiffusion 121 287 122 288  0 t = 3
rlabel pdiffusion 124 287 125 288  0 t = 4
rlabel pdiffusion 120 282 126 288 0 cell no = 326
<< m1 >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< m2 >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< m2c >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< labels >>
rlabel pdiffusion 13 264 14 265  0 t = 1
rlabel pdiffusion 16 264 17 265  0 t = 2
rlabel pdiffusion 13 269 14 270  0 t = 3
rlabel pdiffusion 16 269 17 270  0 t = 4
rlabel pdiffusion 12 264 18 270 0 cell no = 327
<< m1 >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< m2 >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< m2c >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 328
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 85 390 86 391  0 t = 1
rlabel pdiffusion 88 390 89 391  0 t = 2
rlabel pdiffusion 85 395 86 396  0 t = 3
rlabel pdiffusion 88 395 89 396  0 t = 4
rlabel pdiffusion 84 390 90 396 0 cell no = 329
<< m1 >>
rect 85 390 86 391 
rect 88 390 89 391 
rect 85 395 86 396 
rect 88 395 89 396 
<< m2 >>
rect 85 390 86 391 
rect 88 390 89 391 
rect 85 395 86 396 
rect 88 395 89 396 
<< m2c >>
rect 85 390 86 391 
rect 88 390 89 391 
rect 85 395 86 396 
rect 88 395 89 396 
<< labels >>
rlabel pdiffusion 139 300 140 301  0 t = 1
rlabel pdiffusion 142 300 143 301  0 t = 2
rlabel pdiffusion 139 305 140 306  0 t = 3
rlabel pdiffusion 142 305 143 306  0 t = 4
rlabel pdiffusion 138 300 144 306 0 cell no = 330
<< m1 >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< m2 >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< m2c >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< labels >>
rlabel pdiffusion 229 120 230 121  0 t = 1
rlabel pdiffusion 232 120 233 121  0 t = 2
rlabel pdiffusion 229 125 230 126  0 t = 3
rlabel pdiffusion 232 125 233 126  0 t = 4
rlabel pdiffusion 228 120 234 126 0 cell no = 331
<< m1 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2c >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< labels >>
rlabel pdiffusion 157 282 158 283  0 t = 1
rlabel pdiffusion 160 282 161 283  0 t = 2
rlabel pdiffusion 157 287 158 288  0 t = 3
rlabel pdiffusion 160 287 161 288  0 t = 4
rlabel pdiffusion 156 282 162 288 0 cell no = 332
<< m1 >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< m2 >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< m2c >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< labels >>
rlabel pdiffusion 337 120 338 121  0 t = 1
rlabel pdiffusion 340 120 341 121  0 t = 2
rlabel pdiffusion 337 125 338 126  0 t = 3
rlabel pdiffusion 340 125 341 126  0 t = 4
rlabel pdiffusion 336 120 342 126 0 cell no = 333
<< m1 >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< m2 >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< m2c >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< labels >>
rlabel pdiffusion 265 120 266 121  0 t = 1
rlabel pdiffusion 268 120 269 121  0 t = 2
rlabel pdiffusion 265 125 266 126  0 t = 3
rlabel pdiffusion 268 125 269 126  0 t = 4
rlabel pdiffusion 264 120 270 126 0 cell no = 334
<< m1 >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< m2 >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< m2c >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 335
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 336
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 175 336 176 337  0 t = 1
rlabel pdiffusion 178 336 179 337  0 t = 2
rlabel pdiffusion 175 341 176 342  0 t = 3
rlabel pdiffusion 178 341 179 342  0 t = 4
rlabel pdiffusion 174 336 180 342 0 cell no = 337
<< m1 >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< m2 >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< m2c >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< labels >>
rlabel pdiffusion 319 210 320 211  0 t = 1
rlabel pdiffusion 322 210 323 211  0 t = 2
rlabel pdiffusion 319 215 320 216  0 t = 3
rlabel pdiffusion 322 215 323 216  0 t = 4
rlabel pdiffusion 318 210 324 216 0 cell no = 338
<< m1 >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< m2 >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< m2c >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< labels >>
rlabel pdiffusion 103 354 104 355  0 t = 1
rlabel pdiffusion 106 354 107 355  0 t = 2
rlabel pdiffusion 103 359 104 360  0 t = 3
rlabel pdiffusion 106 359 107 360  0 t = 4
rlabel pdiffusion 102 354 108 360 0 cell no = 339
<< m1 >>
rect 103 354 104 355 
rect 106 354 107 355 
rect 103 359 104 360 
rect 106 359 107 360 
<< m2 >>
rect 103 354 104 355 
rect 106 354 107 355 
rect 103 359 104 360 
rect 106 359 107 360 
<< m2c >>
rect 103 354 104 355 
rect 106 354 107 355 
rect 103 359 104 360 
rect 106 359 107 360 
<< labels >>
rlabel pdiffusion 355 246 356 247  0 t = 1
rlabel pdiffusion 358 246 359 247  0 t = 2
rlabel pdiffusion 355 251 356 252  0 t = 3
rlabel pdiffusion 358 251 359 252  0 t = 4
rlabel pdiffusion 354 246 360 252 0 cell no = 340
<< m1 >>
rect 355 246 356 247 
rect 358 246 359 247 
rect 355 251 356 252 
rect 358 251 359 252 
<< m2 >>
rect 355 246 356 247 
rect 358 246 359 247 
rect 355 251 356 252 
rect 358 251 359 252 
<< m2c >>
rect 355 246 356 247 
rect 358 246 359 247 
rect 355 251 356 252 
rect 358 251 359 252 
<< labels >>
rlabel pdiffusion 157 390 158 391  0 t = 1
rlabel pdiffusion 160 390 161 391  0 t = 2
rlabel pdiffusion 157 395 158 396  0 t = 3
rlabel pdiffusion 160 395 161 396  0 t = 4
rlabel pdiffusion 156 390 162 396 0 cell no = 341
<< m1 >>
rect 157 390 158 391 
rect 160 390 161 391 
rect 157 395 158 396 
rect 160 395 161 396 
<< m2 >>
rect 157 390 158 391 
rect 160 390 161 391 
rect 157 395 158 396 
rect 160 395 161 396 
<< m2c >>
rect 157 390 158 391 
rect 160 390 161 391 
rect 157 395 158 396 
rect 160 395 161 396 
<< labels >>
rlabel pdiffusion 211 48 212 49  0 t = 1
rlabel pdiffusion 214 48 215 49  0 t = 2
rlabel pdiffusion 211 53 212 54  0 t = 3
rlabel pdiffusion 214 53 215 54  0 t = 4
rlabel pdiffusion 210 48 216 54 0 cell no = 342
<< m1 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2c >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< labels >>
rlabel pdiffusion 409 264 410 265  0 t = 1
rlabel pdiffusion 412 264 413 265  0 t = 2
rlabel pdiffusion 409 269 410 270  0 t = 3
rlabel pdiffusion 412 269 413 270  0 t = 4
rlabel pdiffusion 408 264 414 270 0 cell no = 343
<< m1 >>
rect 409 264 410 265 
rect 412 264 413 265 
rect 409 269 410 270 
rect 412 269 413 270 
<< m2 >>
rect 409 264 410 265 
rect 412 264 413 265 
rect 409 269 410 270 
rect 412 269 413 270 
<< m2c >>
rect 409 264 410 265 
rect 412 264 413 265 
rect 409 269 410 270 
rect 412 269 413 270 
<< labels >>
rlabel pdiffusion 139 336 140 337  0 t = 1
rlabel pdiffusion 142 336 143 337  0 t = 2
rlabel pdiffusion 139 341 140 342  0 t = 3
rlabel pdiffusion 142 341 143 342  0 t = 4
rlabel pdiffusion 138 336 144 342 0 cell no = 344
<< m1 >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< m2 >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< m2c >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< labels >>
rlabel pdiffusion 445 444 446 445  0 t = 1
rlabel pdiffusion 448 444 449 445  0 t = 2
rlabel pdiffusion 445 449 446 450  0 t = 3
rlabel pdiffusion 448 449 449 450  0 t = 4
rlabel pdiffusion 444 444 450 450 0 cell no = 345
<< m1 >>
rect 445 444 446 445 
rect 448 444 449 445 
rect 445 449 446 450 
rect 448 449 449 450 
<< m2 >>
rect 445 444 446 445 
rect 448 444 449 445 
rect 445 449 446 450 
rect 448 449 449 450 
<< m2c >>
rect 445 444 446 445 
rect 448 444 449 445 
rect 445 449 446 450 
rect 448 449 449 450 
<< labels >>
rlabel pdiffusion 409 300 410 301  0 t = 1
rlabel pdiffusion 412 300 413 301  0 t = 2
rlabel pdiffusion 409 305 410 306  0 t = 3
rlabel pdiffusion 412 305 413 306  0 t = 4
rlabel pdiffusion 408 300 414 306 0 cell no = 346
<< m1 >>
rect 409 300 410 301 
rect 412 300 413 301 
rect 409 305 410 306 
rect 412 305 413 306 
<< m2 >>
rect 409 300 410 301 
rect 412 300 413 301 
rect 409 305 410 306 
rect 412 305 413 306 
<< m2c >>
rect 409 300 410 301 
rect 412 300 413 301 
rect 409 305 410 306 
rect 412 305 413 306 
<< labels >>
rlabel pdiffusion 337 228 338 229  0 t = 1
rlabel pdiffusion 340 228 341 229  0 t = 2
rlabel pdiffusion 337 233 338 234  0 t = 3
rlabel pdiffusion 340 233 341 234  0 t = 4
rlabel pdiffusion 336 228 342 234 0 cell no = 347
<< m1 >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< m2 >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< m2c >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< labels >>
rlabel pdiffusion 427 102 428 103  0 t = 1
rlabel pdiffusion 430 102 431 103  0 t = 2
rlabel pdiffusion 427 107 428 108  0 t = 3
rlabel pdiffusion 430 107 431 108  0 t = 4
rlabel pdiffusion 426 102 432 108 0 cell no = 348
<< m1 >>
rect 427 102 428 103 
rect 430 102 431 103 
rect 427 107 428 108 
rect 430 107 431 108 
<< m2 >>
rect 427 102 428 103 
rect 430 102 431 103 
rect 427 107 428 108 
rect 430 107 431 108 
<< m2c >>
rect 427 102 428 103 
rect 430 102 431 103 
rect 427 107 428 108 
rect 430 107 431 108 
<< labels >>
rlabel pdiffusion 247 66 248 67  0 t = 1
rlabel pdiffusion 250 66 251 67  0 t = 2
rlabel pdiffusion 247 71 248 72  0 t = 3
rlabel pdiffusion 250 71 251 72  0 t = 4
rlabel pdiffusion 246 66 252 72 0 cell no = 349
<< m1 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2c >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< labels >>
rlabel pdiffusion 355 336 356 337  0 t = 1
rlabel pdiffusion 358 336 359 337  0 t = 2
rlabel pdiffusion 355 341 356 342  0 t = 3
rlabel pdiffusion 358 341 359 342  0 t = 4
rlabel pdiffusion 354 336 360 342 0 cell no = 350
<< m1 >>
rect 355 336 356 337 
rect 358 336 359 337 
rect 355 341 356 342 
rect 358 341 359 342 
<< m2 >>
rect 355 336 356 337 
rect 358 336 359 337 
rect 355 341 356 342 
rect 358 341 359 342 
<< m2c >>
rect 355 336 356 337 
rect 358 336 359 337 
rect 355 341 356 342 
rect 358 341 359 342 
<< labels >>
rlabel pdiffusion 67 282 68 283  0 t = 1
rlabel pdiffusion 70 282 71 283  0 t = 2
rlabel pdiffusion 67 287 68 288  0 t = 3
rlabel pdiffusion 70 287 71 288  0 t = 4
rlabel pdiffusion 66 282 72 288 0 cell no = 351
<< m1 >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< m2 >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< m2c >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< labels >>
rlabel pdiffusion 67 300 68 301  0 t = 1
rlabel pdiffusion 70 300 71 301  0 t = 2
rlabel pdiffusion 67 305 68 306  0 t = 3
rlabel pdiffusion 70 305 71 306  0 t = 4
rlabel pdiffusion 66 300 72 306 0 cell no = 352
<< m1 >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< m2 >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< m2c >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< labels >>
rlabel pdiffusion 31 300 32 301  0 t = 1
rlabel pdiffusion 34 300 35 301  0 t = 2
rlabel pdiffusion 31 305 32 306  0 t = 3
rlabel pdiffusion 34 305 35 306  0 t = 4
rlabel pdiffusion 30 300 36 306 0 cell no = 353
<< m1 >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< m2 >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< m2c >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< labels >>
rlabel pdiffusion 49 300 50 301  0 t = 1
rlabel pdiffusion 52 300 53 301  0 t = 2
rlabel pdiffusion 49 305 50 306  0 t = 3
rlabel pdiffusion 52 305 53 306  0 t = 4
rlabel pdiffusion 48 300 54 306 0 cell no = 354
<< m1 >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< m2 >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< m2c >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< labels >>
rlabel pdiffusion 247 48 248 49  0 t = 1
rlabel pdiffusion 250 48 251 49  0 t = 2
rlabel pdiffusion 247 53 248 54  0 t = 3
rlabel pdiffusion 250 53 251 54  0 t = 4
rlabel pdiffusion 246 48 252 54 0 cell no = 355
<< m1 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2c >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 356
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 157 246 158 247  0 t = 1
rlabel pdiffusion 160 246 161 247  0 t = 2
rlabel pdiffusion 157 251 158 252  0 t = 3
rlabel pdiffusion 160 251 161 252  0 t = 4
rlabel pdiffusion 156 246 162 252 0 cell no = 357
<< m1 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2c >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< labels >>
rlabel pdiffusion 139 228 140 229  0 t = 1
rlabel pdiffusion 142 228 143 229  0 t = 2
rlabel pdiffusion 139 233 140 234  0 t = 3
rlabel pdiffusion 142 233 143 234  0 t = 4
rlabel pdiffusion 138 228 144 234 0 cell no = 358
<< m1 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2c >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< labels >>
rlabel pdiffusion 211 300 212 301  0 t = 1
rlabel pdiffusion 214 300 215 301  0 t = 2
rlabel pdiffusion 211 305 212 306  0 t = 3
rlabel pdiffusion 214 305 215 306  0 t = 4
rlabel pdiffusion 210 300 216 306 0 cell no = 359
<< m1 >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< m2 >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< m2c >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< labels >>
rlabel pdiffusion 193 30 194 31  0 t = 1
rlabel pdiffusion 196 30 197 31  0 t = 2
rlabel pdiffusion 193 35 194 36  0 t = 3
rlabel pdiffusion 196 35 197 36  0 t = 4
rlabel pdiffusion 192 30 198 36 0 cell no = 360
<< m1 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2c >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< labels >>
rlabel pdiffusion 193 300 194 301  0 t = 1
rlabel pdiffusion 196 300 197 301  0 t = 2
rlabel pdiffusion 193 305 194 306  0 t = 3
rlabel pdiffusion 196 305 197 306  0 t = 4
rlabel pdiffusion 192 300 198 306 0 cell no = 361
<< m1 >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< m2 >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< m2c >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< labels >>
rlabel pdiffusion 175 102 176 103  0 t = 1
rlabel pdiffusion 178 102 179 103  0 t = 2
rlabel pdiffusion 175 107 176 108  0 t = 3
rlabel pdiffusion 178 107 179 108  0 t = 4
rlabel pdiffusion 174 102 180 108 0 cell no = 362
<< m1 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2c >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 363
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 409 12 410 13  0 t = 1
rlabel pdiffusion 412 12 413 13  0 t = 2
rlabel pdiffusion 409 17 410 18  0 t = 3
rlabel pdiffusion 412 17 413 18  0 t = 4
rlabel pdiffusion 408 12 414 18 0 cell no = 364
<< m1 >>
rect 409 12 410 13 
rect 412 12 413 13 
rect 409 17 410 18 
rect 412 17 413 18 
<< m2 >>
rect 409 12 410 13 
rect 412 12 413 13 
rect 409 17 410 18 
rect 412 17 413 18 
<< m2c >>
rect 409 12 410 13 
rect 412 12 413 13 
rect 409 17 410 18 
rect 412 17 413 18 
<< labels >>
rlabel pdiffusion 427 300 428 301  0 t = 1
rlabel pdiffusion 430 300 431 301  0 t = 2
rlabel pdiffusion 427 305 428 306  0 t = 3
rlabel pdiffusion 430 305 431 306  0 t = 4
rlabel pdiffusion 426 300 432 306 0 cell no = 365
<< m1 >>
rect 427 300 428 301 
rect 430 300 431 301 
rect 427 305 428 306 
rect 430 305 431 306 
<< m2 >>
rect 427 300 428 301 
rect 430 300 431 301 
rect 427 305 428 306 
rect 430 305 431 306 
<< m2c >>
rect 427 300 428 301 
rect 430 300 431 301 
rect 427 305 428 306 
rect 430 305 431 306 
<< labels >>
rlabel pdiffusion 373 336 374 337  0 t = 1
rlabel pdiffusion 376 336 377 337  0 t = 2
rlabel pdiffusion 373 341 374 342  0 t = 3
rlabel pdiffusion 376 341 377 342  0 t = 4
rlabel pdiffusion 372 336 378 342 0 cell no = 366
<< m1 >>
rect 373 336 374 337 
rect 376 336 377 337 
rect 373 341 374 342 
rect 376 341 377 342 
<< m2 >>
rect 373 336 374 337 
rect 376 336 377 337 
rect 373 341 374 342 
rect 376 341 377 342 
<< m2c >>
rect 373 336 374 337 
rect 376 336 377 337 
rect 373 341 374 342 
rect 376 341 377 342 
<< labels >>
rlabel pdiffusion 319 264 320 265  0 t = 1
rlabel pdiffusion 322 264 323 265  0 t = 2
rlabel pdiffusion 319 269 320 270  0 t = 3
rlabel pdiffusion 322 269 323 270  0 t = 4
rlabel pdiffusion 318 264 324 270 0 cell no = 367
<< m1 >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< m2 >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< m2c >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< labels >>
rlabel pdiffusion 391 390 392 391  0 t = 1
rlabel pdiffusion 394 390 395 391  0 t = 2
rlabel pdiffusion 391 395 392 396  0 t = 3
rlabel pdiffusion 394 395 395 396  0 t = 4
rlabel pdiffusion 390 390 396 396 0 cell no = 368
<< m1 >>
rect 391 390 392 391 
rect 394 390 395 391 
rect 391 395 392 396 
rect 394 395 395 396 
<< m2 >>
rect 391 390 392 391 
rect 394 390 395 391 
rect 391 395 392 396 
rect 394 395 395 396 
<< m2c >>
rect 391 390 392 391 
rect 394 390 395 391 
rect 391 395 392 396 
rect 394 395 395 396 
<< labels >>
rlabel pdiffusion 355 156 356 157  0 t = 1
rlabel pdiffusion 358 156 359 157  0 t = 2
rlabel pdiffusion 355 161 356 162  0 t = 3
rlabel pdiffusion 358 161 359 162  0 t = 4
rlabel pdiffusion 354 156 360 162 0 cell no = 369
<< m1 >>
rect 355 156 356 157 
rect 358 156 359 157 
rect 355 161 356 162 
rect 358 161 359 162 
<< m2 >>
rect 355 156 356 157 
rect 358 156 359 157 
rect 355 161 356 162 
rect 358 161 359 162 
<< m2c >>
rect 355 156 356 157 
rect 358 156 359 157 
rect 355 161 356 162 
rect 358 161 359 162 
<< labels >>
rlabel pdiffusion 337 174 338 175  0 t = 1
rlabel pdiffusion 340 174 341 175  0 t = 2
rlabel pdiffusion 337 179 338 180  0 t = 3
rlabel pdiffusion 340 179 341 180  0 t = 4
rlabel pdiffusion 336 174 342 180 0 cell no = 370
<< m1 >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< m2 >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< m2c >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< labels >>
rlabel pdiffusion 355 300 356 301  0 t = 1
rlabel pdiffusion 358 300 359 301  0 t = 2
rlabel pdiffusion 355 305 356 306  0 t = 3
rlabel pdiffusion 358 305 359 306  0 t = 4
rlabel pdiffusion 354 300 360 306 0 cell no = 371
<< m1 >>
rect 355 300 356 301 
rect 358 300 359 301 
rect 355 305 356 306 
rect 358 305 359 306 
<< m2 >>
rect 355 300 356 301 
rect 358 300 359 301 
rect 355 305 356 306 
rect 358 305 359 306 
<< m2c >>
rect 355 300 356 301 
rect 358 300 359 301 
rect 355 305 356 306 
rect 358 305 359 306 
<< labels >>
rlabel pdiffusion 373 264 374 265  0 t = 1
rlabel pdiffusion 376 264 377 265  0 t = 2
rlabel pdiffusion 373 269 374 270  0 t = 3
rlabel pdiffusion 376 269 377 270  0 t = 4
rlabel pdiffusion 372 264 378 270 0 cell no = 372
<< m1 >>
rect 373 264 374 265 
rect 376 264 377 265 
rect 373 269 374 270 
rect 376 269 377 270 
<< m2 >>
rect 373 264 374 265 
rect 376 264 377 265 
rect 373 269 374 270 
rect 376 269 377 270 
<< m2c >>
rect 373 264 374 265 
rect 376 264 377 265 
rect 373 269 374 270 
rect 376 269 377 270 
<< labels >>
rlabel pdiffusion 319 372 320 373  0 t = 1
rlabel pdiffusion 322 372 323 373  0 t = 2
rlabel pdiffusion 319 377 320 378  0 t = 3
rlabel pdiffusion 322 377 323 378  0 t = 4
rlabel pdiffusion 318 372 324 378 0 cell no = 373
<< m1 >>
rect 319 372 320 373 
rect 322 372 323 373 
rect 319 377 320 378 
rect 322 377 323 378 
<< m2 >>
rect 319 372 320 373 
rect 322 372 323 373 
rect 319 377 320 378 
rect 322 377 323 378 
<< m2c >>
rect 319 372 320 373 
rect 322 372 323 373 
rect 319 377 320 378 
rect 322 377 323 378 
<< labels >>
rlabel pdiffusion 121 426 122 427  0 t = 1
rlabel pdiffusion 124 426 125 427  0 t = 2
rlabel pdiffusion 121 431 122 432  0 t = 3
rlabel pdiffusion 124 431 125 432  0 t = 4
rlabel pdiffusion 120 426 126 432 0 cell no = 374
<< m1 >>
rect 121 426 122 427 
rect 124 426 125 427 
rect 121 431 122 432 
rect 124 431 125 432 
<< m2 >>
rect 121 426 122 427 
rect 124 426 125 427 
rect 121 431 122 432 
rect 124 431 125 432 
<< m2c >>
rect 121 426 122 427 
rect 124 426 125 427 
rect 121 431 122 432 
rect 124 431 125 432 
<< labels >>
rlabel pdiffusion 319 354 320 355  0 t = 1
rlabel pdiffusion 322 354 323 355  0 t = 2
rlabel pdiffusion 319 359 320 360  0 t = 3
rlabel pdiffusion 322 359 323 360  0 t = 4
rlabel pdiffusion 318 354 324 360 0 cell no = 375
<< m1 >>
rect 319 354 320 355 
rect 322 354 323 355 
rect 319 359 320 360 
rect 322 359 323 360 
<< m2 >>
rect 319 354 320 355 
rect 322 354 323 355 
rect 319 359 320 360 
rect 322 359 323 360 
<< m2c >>
rect 319 354 320 355 
rect 322 354 323 355 
rect 319 359 320 360 
rect 322 359 323 360 
<< labels >>
rlabel pdiffusion 211 228 212 229  0 t = 1
rlabel pdiffusion 214 228 215 229  0 t = 2
rlabel pdiffusion 211 233 212 234  0 t = 3
rlabel pdiffusion 214 233 215 234  0 t = 4
rlabel pdiffusion 210 228 216 234 0 cell no = 376
<< m1 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2c >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< labels >>
rlabel pdiffusion 49 336 50 337  0 t = 1
rlabel pdiffusion 52 336 53 337  0 t = 2
rlabel pdiffusion 49 341 50 342  0 t = 3
rlabel pdiffusion 52 341 53 342  0 t = 4
rlabel pdiffusion 48 336 54 342 0 cell no = 377
<< m1 >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< m2 >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< m2c >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< labels >>
rlabel pdiffusion 31 174 32 175  0 t = 1
rlabel pdiffusion 34 174 35 175  0 t = 2
rlabel pdiffusion 31 179 32 180  0 t = 3
rlabel pdiffusion 34 179 35 180  0 t = 4
rlabel pdiffusion 30 174 36 180 0 cell no = 378
<< m1 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2c >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< labels >>
rlabel pdiffusion 13 282 14 283  0 t = 1
rlabel pdiffusion 16 282 17 283  0 t = 2
rlabel pdiffusion 13 287 14 288  0 t = 3
rlabel pdiffusion 16 287 17 288  0 t = 4
rlabel pdiffusion 12 282 18 288 0 cell no = 379
<< m1 >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< m2 >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< m2c >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< labels >>
rlabel pdiffusion 157 156 158 157  0 t = 1
rlabel pdiffusion 160 156 161 157  0 t = 2
rlabel pdiffusion 157 161 158 162  0 t = 3
rlabel pdiffusion 160 161 161 162  0 t = 4
rlabel pdiffusion 156 156 162 162 0 cell no = 380
<< m1 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2c >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< labels >>
rlabel pdiffusion 31 390 32 391  0 t = 1
rlabel pdiffusion 34 390 35 391  0 t = 2
rlabel pdiffusion 31 395 32 396  0 t = 3
rlabel pdiffusion 34 395 35 396  0 t = 4
rlabel pdiffusion 30 390 36 396 0 cell no = 381
<< m1 >>
rect 31 390 32 391 
rect 34 390 35 391 
rect 31 395 32 396 
rect 34 395 35 396 
<< m2 >>
rect 31 390 32 391 
rect 34 390 35 391 
rect 31 395 32 396 
rect 34 395 35 396 
<< m2c >>
rect 31 390 32 391 
rect 34 390 35 391 
rect 31 395 32 396 
rect 34 395 35 396 
<< labels >>
rlabel pdiffusion 139 354 140 355  0 t = 1
rlabel pdiffusion 142 354 143 355  0 t = 2
rlabel pdiffusion 139 359 140 360  0 t = 3
rlabel pdiffusion 142 359 143 360  0 t = 4
rlabel pdiffusion 138 354 144 360 0 cell no = 382
<< m1 >>
rect 139 354 140 355 
rect 142 354 143 355 
rect 139 359 140 360 
rect 142 359 143 360 
<< m2 >>
rect 139 354 140 355 
rect 142 354 143 355 
rect 139 359 140 360 
rect 142 359 143 360 
<< m2c >>
rect 139 354 140 355 
rect 142 354 143 355 
rect 139 359 140 360 
rect 142 359 143 360 
<< labels >>
rlabel pdiffusion 103 156 104 157  0 t = 1
rlabel pdiffusion 106 156 107 157  0 t = 2
rlabel pdiffusion 103 161 104 162  0 t = 3
rlabel pdiffusion 106 161 107 162  0 t = 4
rlabel pdiffusion 102 156 108 162 0 cell no = 383
<< m1 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2c >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< labels >>
rlabel pdiffusion 157 318 158 319  0 t = 1
rlabel pdiffusion 160 318 161 319  0 t = 2
rlabel pdiffusion 157 323 158 324  0 t = 3
rlabel pdiffusion 160 323 161 324  0 t = 4
rlabel pdiffusion 156 318 162 324 0 cell no = 384
<< m1 >>
rect 157 318 158 319 
rect 160 318 161 319 
rect 157 323 158 324 
rect 160 323 161 324 
<< m2 >>
rect 157 318 158 319 
rect 160 318 161 319 
rect 157 323 158 324 
rect 160 323 161 324 
<< m2c >>
rect 157 318 158 319 
rect 160 318 161 319 
rect 157 323 158 324 
rect 160 323 161 324 
<< labels >>
rlabel pdiffusion 301 354 302 355  0 t = 1
rlabel pdiffusion 304 354 305 355  0 t = 2
rlabel pdiffusion 301 359 302 360  0 t = 3
rlabel pdiffusion 304 359 305 360  0 t = 4
rlabel pdiffusion 300 354 306 360 0 cell no = 385
<< m1 >>
rect 301 354 302 355 
rect 304 354 305 355 
rect 301 359 302 360 
rect 304 359 305 360 
<< m2 >>
rect 301 354 302 355 
rect 304 354 305 355 
rect 301 359 302 360 
rect 304 359 305 360 
<< m2c >>
rect 301 354 302 355 
rect 304 354 305 355 
rect 301 359 302 360 
rect 304 359 305 360 
<< labels >>
rlabel pdiffusion 193 354 194 355  0 t = 1
rlabel pdiffusion 196 354 197 355  0 t = 2
rlabel pdiffusion 193 359 194 360  0 t = 3
rlabel pdiffusion 196 359 197 360  0 t = 4
rlabel pdiffusion 192 354 198 360 0 cell no = 386
<< m1 >>
rect 193 354 194 355 
rect 196 354 197 355 
rect 193 359 194 360 
rect 196 359 197 360 
<< m2 >>
rect 193 354 194 355 
rect 196 354 197 355 
rect 193 359 194 360 
rect 196 359 197 360 
<< m2c >>
rect 193 354 194 355 
rect 196 354 197 355 
rect 193 359 194 360 
rect 196 359 197 360 
<< labels >>
rlabel pdiffusion 157 264 158 265  0 t = 1
rlabel pdiffusion 160 264 161 265  0 t = 2
rlabel pdiffusion 157 269 158 270  0 t = 3
rlabel pdiffusion 160 269 161 270  0 t = 4
rlabel pdiffusion 156 264 162 270 0 cell no = 387
<< m1 >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< m2 >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< m2c >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< labels >>
rlabel pdiffusion 247 318 248 319  0 t = 1
rlabel pdiffusion 250 318 251 319  0 t = 2
rlabel pdiffusion 247 323 248 324  0 t = 3
rlabel pdiffusion 250 323 251 324  0 t = 4
rlabel pdiffusion 246 318 252 324 0 cell no = 388
<< m1 >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< m2 >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< m2c >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< labels >>
rlabel pdiffusion 67 390 68 391  0 t = 1
rlabel pdiffusion 70 390 71 391  0 t = 2
rlabel pdiffusion 67 395 68 396  0 t = 3
rlabel pdiffusion 70 395 71 396  0 t = 4
rlabel pdiffusion 66 390 72 396 0 cell no = 389
<< m1 >>
rect 67 390 68 391 
rect 70 390 71 391 
rect 67 395 68 396 
rect 70 395 71 396 
<< m2 >>
rect 67 390 68 391 
rect 70 390 71 391 
rect 67 395 68 396 
rect 70 395 71 396 
<< m2c >>
rect 67 390 68 391 
rect 70 390 71 391 
rect 67 395 68 396 
rect 70 395 71 396 
<< labels >>
rlabel pdiffusion 229 264 230 265  0 t = 1
rlabel pdiffusion 232 264 233 265  0 t = 2
rlabel pdiffusion 229 269 230 270  0 t = 3
rlabel pdiffusion 232 269 233 270  0 t = 4
rlabel pdiffusion 228 264 234 270 0 cell no = 390
<< m1 >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< m2 >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< m2c >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< labels >>
rlabel pdiffusion 265 426 266 427  0 t = 1
rlabel pdiffusion 268 426 269 427  0 t = 2
rlabel pdiffusion 265 431 266 432  0 t = 3
rlabel pdiffusion 268 431 269 432  0 t = 4
rlabel pdiffusion 264 426 270 432 0 cell no = 391
<< m1 >>
rect 265 426 266 427 
rect 268 426 269 427 
rect 265 431 266 432 
rect 268 431 269 432 
<< m2 >>
rect 265 426 266 427 
rect 268 426 269 427 
rect 265 431 266 432 
rect 268 431 269 432 
<< m2c >>
rect 265 426 266 427 
rect 268 426 269 427 
rect 265 431 266 432 
rect 268 431 269 432 
<< labels >>
rlabel pdiffusion 319 228 320 229  0 t = 1
rlabel pdiffusion 322 228 323 229  0 t = 2
rlabel pdiffusion 319 233 320 234  0 t = 3
rlabel pdiffusion 322 233 323 234  0 t = 4
rlabel pdiffusion 318 228 324 234 0 cell no = 392
<< m1 >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< m2 >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< m2c >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< labels >>
rlabel pdiffusion 193 228 194 229  0 t = 1
rlabel pdiffusion 196 228 197 229  0 t = 2
rlabel pdiffusion 193 233 194 234  0 t = 3
rlabel pdiffusion 196 233 197 234  0 t = 4
rlabel pdiffusion 192 228 198 234 0 cell no = 393
<< m1 >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< m2 >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< m2c >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< labels >>
rlabel pdiffusion 265 300 266 301  0 t = 1
rlabel pdiffusion 268 300 269 301  0 t = 2
rlabel pdiffusion 265 305 266 306  0 t = 3
rlabel pdiffusion 268 305 269 306  0 t = 4
rlabel pdiffusion 264 300 270 306 0 cell no = 394
<< m1 >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< m2 >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< m2c >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< labels >>
rlabel pdiffusion 391 228 392 229  0 t = 1
rlabel pdiffusion 394 228 395 229  0 t = 2
rlabel pdiffusion 391 233 392 234  0 t = 3
rlabel pdiffusion 394 233 395 234  0 t = 4
rlabel pdiffusion 390 228 396 234 0 cell no = 395
<< m1 >>
rect 391 228 392 229 
rect 394 228 395 229 
rect 391 233 392 234 
rect 394 233 395 234 
<< m2 >>
rect 391 228 392 229 
rect 394 228 395 229 
rect 391 233 392 234 
rect 394 233 395 234 
<< m2c >>
rect 391 228 392 229 
rect 394 228 395 229 
rect 391 233 392 234 
rect 394 233 395 234 
<< labels >>
rlabel pdiffusion 373 426 374 427  0 t = 1
rlabel pdiffusion 376 426 377 427  0 t = 2
rlabel pdiffusion 373 431 374 432  0 t = 3
rlabel pdiffusion 376 431 377 432  0 t = 4
rlabel pdiffusion 372 426 378 432 0 cell no = 396
<< m1 >>
rect 373 426 374 427 
rect 376 426 377 427 
rect 373 431 374 432 
rect 376 431 377 432 
<< m2 >>
rect 373 426 374 427 
rect 376 426 377 427 
rect 373 431 374 432 
rect 376 431 377 432 
<< m2c >>
rect 373 426 374 427 
rect 376 426 377 427 
rect 373 431 374 432 
rect 376 431 377 432 
<< labels >>
rlabel pdiffusion 373 282 374 283  0 t = 1
rlabel pdiffusion 376 282 377 283  0 t = 2
rlabel pdiffusion 373 287 374 288  0 t = 3
rlabel pdiffusion 376 287 377 288  0 t = 4
rlabel pdiffusion 372 282 378 288 0 cell no = 397
<< m1 >>
rect 373 282 374 283 
rect 376 282 377 283 
rect 373 287 374 288 
rect 376 287 377 288 
<< m2 >>
rect 373 282 374 283 
rect 376 282 377 283 
rect 373 287 374 288 
rect 376 287 377 288 
<< m2c >>
rect 373 282 374 283 
rect 376 282 377 283 
rect 373 287 374 288 
rect 376 287 377 288 
<< labels >>
rlabel pdiffusion 445 372 446 373  0 t = 1
rlabel pdiffusion 448 372 449 373  0 t = 2
rlabel pdiffusion 445 377 446 378  0 t = 3
rlabel pdiffusion 448 377 449 378  0 t = 4
rlabel pdiffusion 444 372 450 378 0 cell no = 398
<< m1 >>
rect 445 372 446 373 
rect 448 372 449 373 
rect 445 377 446 378 
rect 448 377 449 378 
<< m2 >>
rect 445 372 446 373 
rect 448 372 449 373 
rect 445 377 446 378 
rect 448 377 449 378 
<< m2c >>
rect 445 372 446 373 
rect 448 372 449 373 
rect 445 377 446 378 
rect 448 377 449 378 
<< labels >>
rlabel pdiffusion 337 282 338 283  0 t = 1
rlabel pdiffusion 340 282 341 283  0 t = 2
rlabel pdiffusion 337 287 338 288  0 t = 3
rlabel pdiffusion 340 287 341 288  0 t = 4
rlabel pdiffusion 336 282 342 288 0 cell no = 399
<< m1 >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< m2 >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< m2c >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< labels >>
rlabel pdiffusion 427 318 428 319  0 t = 1
rlabel pdiffusion 430 318 431 319  0 t = 2
rlabel pdiffusion 427 323 428 324  0 t = 3
rlabel pdiffusion 430 323 431 324  0 t = 4
rlabel pdiffusion 426 318 432 324 0 cell no = 400
<< m1 >>
rect 427 318 428 319 
rect 430 318 431 319 
rect 427 323 428 324 
rect 430 323 431 324 
<< m2 >>
rect 427 318 428 319 
rect 430 318 431 319 
rect 427 323 428 324 
rect 430 323 431 324 
<< m2c >>
rect 427 318 428 319 
rect 430 318 431 319 
rect 427 323 428 324 
rect 430 323 431 324 
<< labels >>
rlabel pdiffusion 247 246 248 247  0 t = 1
rlabel pdiffusion 250 246 251 247  0 t = 2
rlabel pdiffusion 247 251 248 252  0 t = 3
rlabel pdiffusion 250 251 251 252  0 t = 4
rlabel pdiffusion 246 246 252 252 0 cell no = 401
<< m1 >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< m2 >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< m2c >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< labels >>
rlabel pdiffusion 13 318 14 319  0 t = 1
rlabel pdiffusion 16 318 17 319  0 t = 2
rlabel pdiffusion 13 323 14 324  0 t = 3
rlabel pdiffusion 16 323 17 324  0 t = 4
rlabel pdiffusion 12 318 18 324 0 cell no = 402
<< m1 >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< m2 >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< m2c >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< labels >>
rlabel pdiffusion 67 354 68 355  0 t = 1
rlabel pdiffusion 70 354 71 355  0 t = 2
rlabel pdiffusion 67 359 68 360  0 t = 3
rlabel pdiffusion 70 359 71 360  0 t = 4
rlabel pdiffusion 66 354 72 360 0 cell no = 403
<< m1 >>
rect 67 354 68 355 
rect 70 354 71 355 
rect 67 359 68 360 
rect 70 359 71 360 
<< m2 >>
rect 67 354 68 355 
rect 70 354 71 355 
rect 67 359 68 360 
rect 70 359 71 360 
<< m2c >>
rect 67 354 68 355 
rect 70 354 71 355 
rect 67 359 68 360 
rect 70 359 71 360 
<< labels >>
rlabel pdiffusion 49 210 50 211  0 t = 1
rlabel pdiffusion 52 210 53 211  0 t = 2
rlabel pdiffusion 49 215 50 216  0 t = 3
rlabel pdiffusion 52 215 53 216  0 t = 4
rlabel pdiffusion 48 210 54 216 0 cell no = 404
<< m1 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2c >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< labels >>
rlabel pdiffusion 103 246 104 247  0 t = 1
rlabel pdiffusion 106 246 107 247  0 t = 2
rlabel pdiffusion 103 251 104 252  0 t = 3
rlabel pdiffusion 106 251 107 252  0 t = 4
rlabel pdiffusion 102 246 108 252 0 cell no = 405
<< m1 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2c >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< labels >>
rlabel pdiffusion 157 354 158 355  0 t = 1
rlabel pdiffusion 160 354 161 355  0 t = 2
rlabel pdiffusion 157 359 158 360  0 t = 3
rlabel pdiffusion 160 359 161 360  0 t = 4
rlabel pdiffusion 156 354 162 360 0 cell no = 406
<< m1 >>
rect 157 354 158 355 
rect 160 354 161 355 
rect 157 359 158 360 
rect 160 359 161 360 
<< m2 >>
rect 157 354 158 355 
rect 160 354 161 355 
rect 157 359 158 360 
rect 160 359 161 360 
<< m2c >>
rect 157 354 158 355 
rect 160 354 161 355 
rect 157 359 158 360 
rect 160 359 161 360 
<< labels >>
rlabel pdiffusion 211 282 212 283  0 t = 1
rlabel pdiffusion 214 282 215 283  0 t = 2
rlabel pdiffusion 211 287 212 288  0 t = 3
rlabel pdiffusion 214 287 215 288  0 t = 4
rlabel pdiffusion 210 282 216 288 0 cell no = 407
<< m1 >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< m2 >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< m2c >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< labels >>
rlabel pdiffusion 211 264 212 265  0 t = 1
rlabel pdiffusion 214 264 215 265  0 t = 2
rlabel pdiffusion 211 269 212 270  0 t = 3
rlabel pdiffusion 214 269 215 270  0 t = 4
rlabel pdiffusion 210 264 216 270 0 cell no = 408
<< m1 >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< m2 >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< m2c >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< labels >>
rlabel pdiffusion 139 408 140 409  0 t = 1
rlabel pdiffusion 142 408 143 409  0 t = 2
rlabel pdiffusion 139 413 140 414  0 t = 3
rlabel pdiffusion 142 413 143 414  0 t = 4
rlabel pdiffusion 138 408 144 414 0 cell no = 409
<< m1 >>
rect 139 408 140 409 
rect 142 408 143 409 
rect 139 413 140 414 
rect 142 413 143 414 
<< m2 >>
rect 139 408 140 409 
rect 142 408 143 409 
rect 139 413 140 414 
rect 142 413 143 414 
<< m2c >>
rect 139 408 140 409 
rect 142 408 143 409 
rect 139 413 140 414 
rect 142 413 143 414 
<< labels >>
rlabel pdiffusion 31 84 32 85  0 t = 1
rlabel pdiffusion 34 84 35 85  0 t = 2
rlabel pdiffusion 31 89 32 90  0 t = 3
rlabel pdiffusion 34 89 35 90  0 t = 4
rlabel pdiffusion 30 84 36 90 0 cell no = 410
<< m1 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2c >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< labels >>
rlabel pdiffusion 355 390 356 391  0 t = 1
rlabel pdiffusion 358 390 359 391  0 t = 2
rlabel pdiffusion 355 395 356 396  0 t = 3
rlabel pdiffusion 358 395 359 396  0 t = 4
rlabel pdiffusion 354 390 360 396 0 cell no = 411
<< m1 >>
rect 355 390 356 391 
rect 358 390 359 391 
rect 355 395 356 396 
rect 358 395 359 396 
<< m2 >>
rect 355 390 356 391 
rect 358 390 359 391 
rect 355 395 356 396 
rect 358 395 359 396 
<< m2c >>
rect 355 390 356 391 
rect 358 390 359 391 
rect 355 395 356 396 
rect 358 395 359 396 
<< labels >>
rlabel pdiffusion 175 444 176 445  0 t = 1
rlabel pdiffusion 178 444 179 445  0 t = 2
rlabel pdiffusion 175 449 176 450  0 t = 3
rlabel pdiffusion 178 449 179 450  0 t = 4
rlabel pdiffusion 174 444 180 450 0 cell no = 412
<< m1 >>
rect 175 444 176 445 
rect 178 444 179 445 
rect 175 449 176 450 
rect 178 449 179 450 
<< m2 >>
rect 175 444 176 445 
rect 178 444 179 445 
rect 175 449 176 450 
rect 178 449 179 450 
<< m2c >>
rect 175 444 176 445 
rect 178 444 179 445 
rect 175 449 176 450 
rect 178 449 179 450 
<< labels >>
rlabel pdiffusion 319 336 320 337  0 t = 1
rlabel pdiffusion 322 336 323 337  0 t = 2
rlabel pdiffusion 319 341 320 342  0 t = 3
rlabel pdiffusion 322 341 323 342  0 t = 4
rlabel pdiffusion 318 336 324 342 0 cell no = 413
<< m1 >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< m2 >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< m2c >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< labels >>
rlabel pdiffusion 211 120 212 121  0 t = 1
rlabel pdiffusion 214 120 215 121  0 t = 2
rlabel pdiffusion 211 125 212 126  0 t = 3
rlabel pdiffusion 214 125 215 126  0 t = 4
rlabel pdiffusion 210 120 216 126 0 cell no = 414
<< m1 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2c >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< labels >>
rlabel pdiffusion 175 426 176 427  0 t = 1
rlabel pdiffusion 178 426 179 427  0 t = 2
rlabel pdiffusion 175 431 176 432  0 t = 3
rlabel pdiffusion 178 431 179 432  0 t = 4
rlabel pdiffusion 174 426 180 432 0 cell no = 415
<< m1 >>
rect 175 426 176 427 
rect 178 426 179 427 
rect 175 431 176 432 
rect 178 431 179 432 
<< m2 >>
rect 175 426 176 427 
rect 178 426 179 427 
rect 175 431 176 432 
rect 178 431 179 432 
<< m2c >>
rect 175 426 176 427 
rect 178 426 179 427 
rect 175 431 176 432 
rect 178 431 179 432 
<< labels >>
rlabel pdiffusion 445 318 446 319  0 t = 1
rlabel pdiffusion 448 318 449 319  0 t = 2
rlabel pdiffusion 445 323 446 324  0 t = 3
rlabel pdiffusion 448 323 449 324  0 t = 4
rlabel pdiffusion 444 318 450 324 0 cell no = 416
<< m1 >>
rect 445 318 446 319 
rect 448 318 449 319 
rect 445 323 446 324 
rect 448 323 449 324 
<< m2 >>
rect 445 318 446 319 
rect 448 318 449 319 
rect 445 323 446 324 
rect 448 323 449 324 
<< m2c >>
rect 445 318 446 319 
rect 448 318 449 319 
rect 445 323 446 324 
rect 448 323 449 324 
<< labels >>
rlabel pdiffusion 373 354 374 355  0 t = 1
rlabel pdiffusion 376 354 377 355  0 t = 2
rlabel pdiffusion 373 359 374 360  0 t = 3
rlabel pdiffusion 376 359 377 360  0 t = 4
rlabel pdiffusion 372 354 378 360 0 cell no = 417
<< m1 >>
rect 373 354 374 355 
rect 376 354 377 355 
rect 373 359 374 360 
rect 376 359 377 360 
<< m2 >>
rect 373 354 374 355 
rect 376 354 377 355 
rect 373 359 374 360 
rect 376 359 377 360 
<< m2c >>
rect 373 354 374 355 
rect 376 354 377 355 
rect 373 359 374 360 
rect 376 359 377 360 
<< labels >>
rlabel pdiffusion 391 246 392 247  0 t = 1
rlabel pdiffusion 394 246 395 247  0 t = 2
rlabel pdiffusion 391 251 392 252  0 t = 3
rlabel pdiffusion 394 251 395 252  0 t = 4
rlabel pdiffusion 390 246 396 252 0 cell no = 418
<< m1 >>
rect 391 246 392 247 
rect 394 246 395 247 
rect 391 251 392 252 
rect 394 251 395 252 
<< m2 >>
rect 391 246 392 247 
rect 394 246 395 247 
rect 391 251 392 252 
rect 394 251 395 252 
<< m2c >>
rect 391 246 392 247 
rect 394 246 395 247 
rect 391 251 392 252 
rect 394 251 395 252 
<< labels >>
rlabel pdiffusion 337 300 338 301  0 t = 1
rlabel pdiffusion 340 300 341 301  0 t = 2
rlabel pdiffusion 337 305 338 306  0 t = 3
rlabel pdiffusion 340 305 341 306  0 t = 4
rlabel pdiffusion 336 300 342 306 0 cell no = 419
<< m1 >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< m2 >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< m2c >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< labels >>
rlabel pdiffusion 211 246 212 247  0 t = 1
rlabel pdiffusion 214 246 215 247  0 t = 2
rlabel pdiffusion 211 251 212 252  0 t = 3
rlabel pdiffusion 214 251 215 252  0 t = 4
rlabel pdiffusion 210 246 216 252 0 cell no = 420
<< m1 >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< m2 >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< m2c >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< labels >>
rlabel pdiffusion 391 354 392 355  0 t = 1
rlabel pdiffusion 394 354 395 355  0 t = 2
rlabel pdiffusion 391 359 392 360  0 t = 3
rlabel pdiffusion 394 359 395 360  0 t = 4
rlabel pdiffusion 390 354 396 360 0 cell no = 421
<< m1 >>
rect 391 354 392 355 
rect 394 354 395 355 
rect 391 359 392 360 
rect 394 359 395 360 
<< m2 >>
rect 391 354 392 355 
rect 394 354 395 355 
rect 391 359 392 360 
rect 394 359 395 360 
<< m2c >>
rect 391 354 392 355 
rect 394 354 395 355 
rect 391 359 392 360 
rect 394 359 395 360 
<< labels >>
rlabel pdiffusion 409 372 410 373  0 t = 1
rlabel pdiffusion 412 372 413 373  0 t = 2
rlabel pdiffusion 409 377 410 378  0 t = 3
rlabel pdiffusion 412 377 413 378  0 t = 4
rlabel pdiffusion 408 372 414 378 0 cell no = 422
<< m1 >>
rect 409 372 410 373 
rect 412 372 413 373 
rect 409 377 410 378 
rect 412 377 413 378 
<< m2 >>
rect 409 372 410 373 
rect 412 372 413 373 
rect 409 377 410 378 
rect 412 377 413 378 
<< m2c >>
rect 409 372 410 373 
rect 412 372 413 373 
rect 409 377 410 378 
rect 412 377 413 378 
<< labels >>
rlabel pdiffusion 373 390 374 391  0 t = 1
rlabel pdiffusion 376 390 377 391  0 t = 2
rlabel pdiffusion 373 395 374 396  0 t = 3
rlabel pdiffusion 376 395 377 396  0 t = 4
rlabel pdiffusion 372 390 378 396 0 cell no = 423
<< m1 >>
rect 373 390 374 391 
rect 376 390 377 391 
rect 373 395 374 396 
rect 376 395 377 396 
<< m2 >>
rect 373 390 374 391 
rect 376 390 377 391 
rect 373 395 374 396 
rect 376 395 377 396 
<< m2c >>
rect 373 390 374 391 
rect 376 390 377 391 
rect 373 395 374 396 
rect 376 395 377 396 
<< labels >>
rlabel pdiffusion 427 372 428 373  0 t = 1
rlabel pdiffusion 430 372 431 373  0 t = 2
rlabel pdiffusion 427 377 428 378  0 t = 3
rlabel pdiffusion 430 377 431 378  0 t = 4
rlabel pdiffusion 426 372 432 378 0 cell no = 424
<< m1 >>
rect 427 372 428 373 
rect 430 372 431 373 
rect 427 377 428 378 
rect 430 377 431 378 
<< m2 >>
rect 427 372 428 373 
rect 430 372 431 373 
rect 427 377 428 378 
rect 430 377 431 378 
<< m2c >>
rect 427 372 428 373 
rect 430 372 431 373 
rect 427 377 428 378 
rect 430 377 431 378 
<< labels >>
rlabel pdiffusion 283 300 284 301  0 t = 1
rlabel pdiffusion 286 300 287 301  0 t = 2
rlabel pdiffusion 283 305 284 306  0 t = 3
rlabel pdiffusion 286 305 287 306  0 t = 4
rlabel pdiffusion 282 300 288 306 0 cell no = 425
<< m1 >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< m2 >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< m2c >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< labels >>
rlabel pdiffusion 13 372 14 373  0 t = 1
rlabel pdiffusion 16 372 17 373  0 t = 2
rlabel pdiffusion 13 377 14 378  0 t = 3
rlabel pdiffusion 16 377 17 378  0 t = 4
rlabel pdiffusion 12 372 18 378 0 cell no = 426
<< m1 >>
rect 13 372 14 373 
rect 16 372 17 373 
rect 13 377 14 378 
rect 16 377 17 378 
<< m2 >>
rect 13 372 14 373 
rect 16 372 17 373 
rect 13 377 14 378 
rect 16 377 17 378 
<< m2c >>
rect 13 372 14 373 
rect 16 372 17 373 
rect 13 377 14 378 
rect 16 377 17 378 
<< labels >>
rlabel pdiffusion 85 354 86 355  0 t = 1
rlabel pdiffusion 88 354 89 355  0 t = 2
rlabel pdiffusion 85 359 86 360  0 t = 3
rlabel pdiffusion 88 359 89 360  0 t = 4
rlabel pdiffusion 84 354 90 360 0 cell no = 427
<< m1 >>
rect 85 354 86 355 
rect 88 354 89 355 
rect 85 359 86 360 
rect 88 359 89 360 
<< m2 >>
rect 85 354 86 355 
rect 88 354 89 355 
rect 85 359 86 360 
rect 88 359 89 360 
<< m2c >>
rect 85 354 86 355 
rect 88 354 89 355 
rect 85 359 86 360 
rect 88 359 89 360 
<< labels >>
rlabel pdiffusion 31 426 32 427  0 t = 1
rlabel pdiffusion 34 426 35 427  0 t = 2
rlabel pdiffusion 31 431 32 432  0 t = 3
rlabel pdiffusion 34 431 35 432  0 t = 4
rlabel pdiffusion 30 426 36 432 0 cell no = 428
<< m1 >>
rect 31 426 32 427 
rect 34 426 35 427 
rect 31 431 32 432 
rect 34 431 35 432 
<< m2 >>
rect 31 426 32 427 
rect 34 426 35 427 
rect 31 431 32 432 
rect 34 431 35 432 
<< m2c >>
rect 31 426 32 427 
rect 34 426 35 427 
rect 31 431 32 432 
rect 34 431 35 432 
<< labels >>
rlabel pdiffusion 121 372 122 373  0 t = 1
rlabel pdiffusion 124 372 125 373  0 t = 2
rlabel pdiffusion 121 377 122 378  0 t = 3
rlabel pdiffusion 124 377 125 378  0 t = 4
rlabel pdiffusion 120 372 126 378 0 cell no = 429
<< m1 >>
rect 121 372 122 373 
rect 124 372 125 373 
rect 121 377 122 378 
rect 124 377 125 378 
<< m2 >>
rect 121 372 122 373 
rect 124 372 125 373 
rect 121 377 122 378 
rect 124 377 125 378 
<< m2c >>
rect 121 372 122 373 
rect 124 372 125 373 
rect 121 377 122 378 
rect 124 377 125 378 
<< labels >>
rlabel pdiffusion 283 354 284 355  0 t = 1
rlabel pdiffusion 286 354 287 355  0 t = 2
rlabel pdiffusion 283 359 284 360  0 t = 3
rlabel pdiffusion 286 359 287 360  0 t = 4
rlabel pdiffusion 282 354 288 360 0 cell no = 430
<< m1 >>
rect 283 354 284 355 
rect 286 354 287 355 
rect 283 359 284 360 
rect 286 359 287 360 
<< m2 >>
rect 283 354 284 355 
rect 286 354 287 355 
rect 283 359 284 360 
rect 286 359 287 360 
<< m2c >>
rect 283 354 284 355 
rect 286 354 287 355 
rect 283 359 284 360 
rect 286 359 287 360 
<< labels >>
rlabel pdiffusion 103 372 104 373  0 t = 1
rlabel pdiffusion 106 372 107 373  0 t = 2
rlabel pdiffusion 103 377 104 378  0 t = 3
rlabel pdiffusion 106 377 107 378  0 t = 4
rlabel pdiffusion 102 372 108 378 0 cell no = 431
<< m1 >>
rect 103 372 104 373 
rect 106 372 107 373 
rect 103 377 104 378 
rect 106 377 107 378 
<< m2 >>
rect 103 372 104 373 
rect 106 372 107 373 
rect 103 377 104 378 
rect 106 377 107 378 
<< m2c >>
rect 103 372 104 373 
rect 106 372 107 373 
rect 103 377 104 378 
rect 106 377 107 378 
<< labels >>
rlabel pdiffusion 67 372 68 373  0 t = 1
rlabel pdiffusion 70 372 71 373  0 t = 2
rlabel pdiffusion 67 377 68 378  0 t = 3
rlabel pdiffusion 70 377 71 378  0 t = 4
rlabel pdiffusion 66 372 72 378 0 cell no = 432
<< m1 >>
rect 67 372 68 373 
rect 70 372 71 373 
rect 67 377 68 378 
rect 70 377 71 378 
<< m2 >>
rect 67 372 68 373 
rect 70 372 71 373 
rect 67 377 68 378 
rect 70 377 71 378 
<< m2c >>
rect 67 372 68 373 
rect 70 372 71 373 
rect 67 377 68 378 
rect 70 377 71 378 
<< labels >>
rlabel pdiffusion 337 210 338 211  0 t = 1
rlabel pdiffusion 340 210 341 211  0 t = 2
rlabel pdiffusion 337 215 338 216  0 t = 3
rlabel pdiffusion 340 215 341 216  0 t = 4
rlabel pdiffusion 336 210 342 216 0 cell no = 433
<< m1 >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< m2 >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< m2c >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< labels >>
rlabel pdiffusion 139 390 140 391  0 t = 1
rlabel pdiffusion 142 390 143 391  0 t = 2
rlabel pdiffusion 139 395 140 396  0 t = 3
rlabel pdiffusion 142 395 143 396  0 t = 4
rlabel pdiffusion 138 390 144 396 0 cell no = 434
<< m1 >>
rect 139 390 140 391 
rect 142 390 143 391 
rect 139 395 140 396 
rect 142 395 143 396 
<< m2 >>
rect 139 390 140 391 
rect 142 390 143 391 
rect 139 395 140 396 
rect 142 395 143 396 
<< m2c >>
rect 139 390 140 391 
rect 142 390 143 391 
rect 139 395 140 396 
rect 142 395 143 396 
<< labels >>
rlabel pdiffusion 193 336 194 337  0 t = 1
rlabel pdiffusion 196 336 197 337  0 t = 2
rlabel pdiffusion 193 341 194 342  0 t = 3
rlabel pdiffusion 196 341 197 342  0 t = 4
rlabel pdiffusion 192 336 198 342 0 cell no = 435
<< m1 >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< m2 >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< m2c >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< labels >>
rlabel pdiffusion 31 408 32 409  0 t = 1
rlabel pdiffusion 34 408 35 409  0 t = 2
rlabel pdiffusion 31 413 32 414  0 t = 3
rlabel pdiffusion 34 413 35 414  0 t = 4
rlabel pdiffusion 30 408 36 414 0 cell no = 436
<< m1 >>
rect 31 408 32 409 
rect 34 408 35 409 
rect 31 413 32 414 
rect 34 413 35 414 
<< m2 >>
rect 31 408 32 409 
rect 34 408 35 409 
rect 31 413 32 414 
rect 34 413 35 414 
<< m2c >>
rect 31 408 32 409 
rect 34 408 35 409 
rect 31 413 32 414 
rect 34 413 35 414 
<< labels >>
rlabel pdiffusion 247 156 248 157  0 t = 1
rlabel pdiffusion 250 156 251 157  0 t = 2
rlabel pdiffusion 247 161 248 162  0 t = 3
rlabel pdiffusion 250 161 251 162  0 t = 4
rlabel pdiffusion 246 156 252 162 0 cell no = 437
<< m1 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2c >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< labels >>
rlabel pdiffusion 103 282 104 283  0 t = 1
rlabel pdiffusion 106 282 107 283  0 t = 2
rlabel pdiffusion 103 287 104 288  0 t = 3
rlabel pdiffusion 106 287 107 288  0 t = 4
rlabel pdiffusion 102 282 108 288 0 cell no = 438
<< m1 >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< m2 >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< m2c >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< labels >>
rlabel pdiffusion 121 264 122 265  0 t = 1
rlabel pdiffusion 124 264 125 265  0 t = 2
rlabel pdiffusion 121 269 122 270  0 t = 3
rlabel pdiffusion 124 269 125 270  0 t = 4
rlabel pdiffusion 120 264 126 270 0 cell no = 439
<< m1 >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< m2 >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< m2c >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< labels >>
rlabel pdiffusion 319 300 320 301  0 t = 1
rlabel pdiffusion 322 300 323 301  0 t = 2
rlabel pdiffusion 319 305 320 306  0 t = 3
rlabel pdiffusion 322 305 323 306  0 t = 4
rlabel pdiffusion 318 300 324 306 0 cell no = 440
<< m1 >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< m2 >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< m2c >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< labels >>
rlabel pdiffusion 391 426 392 427  0 t = 1
rlabel pdiffusion 394 426 395 427  0 t = 2
rlabel pdiffusion 391 431 392 432  0 t = 3
rlabel pdiffusion 394 431 395 432  0 t = 4
rlabel pdiffusion 390 426 396 432 0 cell no = 441
<< m1 >>
rect 391 426 392 427 
rect 394 426 395 427 
rect 391 431 392 432 
rect 394 431 395 432 
<< m2 >>
rect 391 426 392 427 
rect 394 426 395 427 
rect 391 431 392 432 
rect 394 431 395 432 
<< m2c >>
rect 391 426 392 427 
rect 394 426 395 427 
rect 391 431 392 432 
rect 394 431 395 432 
<< labels >>
rlabel pdiffusion 391 210 392 211  0 t = 1
rlabel pdiffusion 394 210 395 211  0 t = 2
rlabel pdiffusion 391 215 392 216  0 t = 3
rlabel pdiffusion 394 215 395 216  0 t = 4
rlabel pdiffusion 390 210 396 216 0 cell no = 442
<< m1 >>
rect 391 210 392 211 
rect 394 210 395 211 
rect 391 215 392 216 
rect 394 215 395 216 
<< m2 >>
rect 391 210 392 211 
rect 394 210 395 211 
rect 391 215 392 216 
rect 394 215 395 216 
<< m2c >>
rect 391 210 392 211 
rect 394 210 395 211 
rect 391 215 392 216 
rect 394 215 395 216 
<< labels >>
rlabel pdiffusion 391 282 392 283  0 t = 1
rlabel pdiffusion 394 282 395 283  0 t = 2
rlabel pdiffusion 391 287 392 288  0 t = 3
rlabel pdiffusion 394 287 395 288  0 t = 4
rlabel pdiffusion 390 282 396 288 0 cell no = 443
<< m1 >>
rect 391 282 392 283 
rect 394 282 395 283 
rect 391 287 392 288 
rect 394 287 395 288 
<< m2 >>
rect 391 282 392 283 
rect 394 282 395 283 
rect 391 287 392 288 
rect 394 287 395 288 
<< m2c >>
rect 391 282 392 283 
rect 394 282 395 283 
rect 391 287 392 288 
rect 394 287 395 288 
<< labels >>
rlabel pdiffusion 13 444 14 445  0 t = 1
rlabel pdiffusion 16 444 17 445  0 t = 2
rlabel pdiffusion 13 449 14 450  0 t = 3
rlabel pdiffusion 16 449 17 450  0 t = 4
rlabel pdiffusion 12 444 18 450 0 cell no = 444
<< m1 >>
rect 13 444 14 445 
rect 16 444 17 445 
rect 13 449 14 450 
rect 16 449 17 450 
<< m2 >>
rect 13 444 14 445 
rect 16 444 17 445 
rect 13 449 14 450 
rect 16 449 17 450 
<< m2c >>
rect 13 444 14 445 
rect 16 444 17 445 
rect 13 449 14 450 
rect 16 449 17 450 
<< labels >>
rlabel pdiffusion 283 426 284 427  0 t = 1
rlabel pdiffusion 286 426 287 427  0 t = 2
rlabel pdiffusion 283 431 284 432  0 t = 3
rlabel pdiffusion 286 431 287 432  0 t = 4
rlabel pdiffusion 282 426 288 432 0 cell no = 445
<< m1 >>
rect 283 426 284 427 
rect 286 426 287 427 
rect 283 431 284 432 
rect 286 431 287 432 
<< m2 >>
rect 283 426 284 427 
rect 286 426 287 427 
rect 283 431 284 432 
rect 286 431 287 432 
<< m2c >>
rect 283 426 284 427 
rect 286 426 287 427 
rect 283 431 284 432 
rect 286 431 287 432 
<< labels >>
rlabel pdiffusion 373 318 374 319  0 t = 1
rlabel pdiffusion 376 318 377 319  0 t = 2
rlabel pdiffusion 373 323 374 324  0 t = 3
rlabel pdiffusion 376 323 377 324  0 t = 4
rlabel pdiffusion 372 318 378 324 0 cell no = 446
<< m1 >>
rect 373 318 374 319 
rect 376 318 377 319 
rect 373 323 374 324 
rect 376 323 377 324 
<< m2 >>
rect 373 318 374 319 
rect 376 318 377 319 
rect 373 323 374 324 
rect 376 323 377 324 
<< m2c >>
rect 373 318 374 319 
rect 376 318 377 319 
rect 373 323 374 324 
rect 376 323 377 324 
<< labels >>
rlabel pdiffusion 409 228 410 229  0 t = 1
rlabel pdiffusion 412 228 413 229  0 t = 2
rlabel pdiffusion 409 233 410 234  0 t = 3
rlabel pdiffusion 412 233 413 234  0 t = 4
rlabel pdiffusion 408 228 414 234 0 cell no = 447
<< m1 >>
rect 409 228 410 229 
rect 412 228 413 229 
rect 409 233 410 234 
rect 412 233 413 234 
<< m2 >>
rect 409 228 410 229 
rect 412 228 413 229 
rect 409 233 410 234 
rect 412 233 413 234 
<< m2c >>
rect 409 228 410 229 
rect 412 228 413 229 
rect 409 233 410 234 
rect 412 233 413 234 
<< labels >>
rlabel pdiffusion 121 84 122 85  0 t = 1
rlabel pdiffusion 124 84 125 85  0 t = 2
rlabel pdiffusion 121 89 122 90  0 t = 3
rlabel pdiffusion 124 89 125 90  0 t = 4
rlabel pdiffusion 120 84 126 90 0 cell no = 448
<< m1 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2c >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< labels >>
rlabel pdiffusion 391 300 392 301  0 t = 1
rlabel pdiffusion 394 300 395 301  0 t = 2
rlabel pdiffusion 391 305 392 306  0 t = 3
rlabel pdiffusion 394 305 395 306  0 t = 4
rlabel pdiffusion 390 300 396 306 0 cell no = 449
<< m1 >>
rect 391 300 392 301 
rect 394 300 395 301 
rect 391 305 392 306 
rect 394 305 395 306 
<< m2 >>
rect 391 300 392 301 
rect 394 300 395 301 
rect 391 305 392 306 
rect 394 305 395 306 
<< m2c >>
rect 391 300 392 301 
rect 394 300 395 301 
rect 391 305 392 306 
rect 394 305 395 306 
<< labels >>
rlabel pdiffusion 445 354 446 355  0 t = 1
rlabel pdiffusion 448 354 449 355  0 t = 2
rlabel pdiffusion 445 359 446 360  0 t = 3
rlabel pdiffusion 448 359 449 360  0 t = 4
rlabel pdiffusion 444 354 450 360 0 cell no = 450
<< m1 >>
rect 445 354 446 355 
rect 448 354 449 355 
rect 445 359 446 360 
rect 448 359 449 360 
<< m2 >>
rect 445 354 446 355 
rect 448 354 449 355 
rect 445 359 446 360 
rect 448 359 449 360 
<< m2c >>
rect 445 354 446 355 
rect 448 354 449 355 
rect 445 359 446 360 
rect 448 359 449 360 
<< labels >>
rlabel pdiffusion 337 84 338 85  0 t = 1
rlabel pdiffusion 340 84 341 85  0 t = 2
rlabel pdiffusion 337 89 338 90  0 t = 3
rlabel pdiffusion 340 89 341 90  0 t = 4
rlabel pdiffusion 336 84 342 90 0 cell no = 451
<< m1 >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< m2 >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< m2c >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< labels >>
rlabel pdiffusion 157 336 158 337  0 t = 1
rlabel pdiffusion 160 336 161 337  0 t = 2
rlabel pdiffusion 157 341 158 342  0 t = 3
rlabel pdiffusion 160 341 161 342  0 t = 4
rlabel pdiffusion 156 336 162 342 0 cell no = 452
<< m1 >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< m2 >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< m2c >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< labels >>
rlabel pdiffusion 49 282 50 283  0 t = 1
rlabel pdiffusion 52 282 53 283  0 t = 2
rlabel pdiffusion 49 287 50 288  0 t = 3
rlabel pdiffusion 52 287 53 288  0 t = 4
rlabel pdiffusion 48 282 54 288 0 cell no = 453
<< m1 >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< m2 >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< m2c >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< labels >>
rlabel pdiffusion 67 408 68 409  0 t = 1
rlabel pdiffusion 70 408 71 409  0 t = 2
rlabel pdiffusion 67 413 68 414  0 t = 3
rlabel pdiffusion 70 413 71 414  0 t = 4
rlabel pdiffusion 66 408 72 414 0 cell no = 454
<< m1 >>
rect 67 408 68 409 
rect 70 408 71 409 
rect 67 413 68 414 
rect 70 413 71 414 
<< m2 >>
rect 67 408 68 409 
rect 70 408 71 409 
rect 67 413 68 414 
rect 70 413 71 414 
<< m2c >>
rect 67 408 68 409 
rect 70 408 71 409 
rect 67 413 68 414 
rect 70 413 71 414 
<< labels >>
rlabel pdiffusion 85 300 86 301  0 t = 1
rlabel pdiffusion 88 300 89 301  0 t = 2
rlabel pdiffusion 85 305 86 306  0 t = 3
rlabel pdiffusion 88 305 89 306  0 t = 4
rlabel pdiffusion 84 300 90 306 0 cell no = 455
<< m1 >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< m2 >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< m2c >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< labels >>
rlabel pdiffusion 67 426 68 427  0 t = 1
rlabel pdiffusion 70 426 71 427  0 t = 2
rlabel pdiffusion 67 431 68 432  0 t = 3
rlabel pdiffusion 70 431 71 432  0 t = 4
rlabel pdiffusion 66 426 72 432 0 cell no = 456
<< m1 >>
rect 67 426 68 427 
rect 70 426 71 427 
rect 67 431 68 432 
rect 70 431 71 432 
<< m2 >>
rect 67 426 68 427 
rect 70 426 71 427 
rect 67 431 68 432 
rect 70 431 71 432 
<< m2c >>
rect 67 426 68 427 
rect 70 426 71 427 
rect 67 431 68 432 
rect 70 431 71 432 
<< labels >>
rlabel pdiffusion 103 336 104 337  0 t = 1
rlabel pdiffusion 106 336 107 337  0 t = 2
rlabel pdiffusion 103 341 104 342  0 t = 3
rlabel pdiffusion 106 341 107 342  0 t = 4
rlabel pdiffusion 102 336 108 342 0 cell no = 457
<< m1 >>
rect 103 336 104 337 
rect 106 336 107 337 
rect 103 341 104 342 
rect 106 341 107 342 
<< m2 >>
rect 103 336 104 337 
rect 106 336 107 337 
rect 103 341 104 342 
rect 106 341 107 342 
<< m2c >>
rect 103 336 104 337 
rect 106 336 107 337 
rect 103 341 104 342 
rect 106 341 107 342 
<< labels >>
rlabel pdiffusion 121 390 122 391  0 t = 1
rlabel pdiffusion 124 390 125 391  0 t = 2
rlabel pdiffusion 121 395 122 396  0 t = 3
rlabel pdiffusion 124 395 125 396  0 t = 4
rlabel pdiffusion 120 390 126 396 0 cell no = 458
<< m1 >>
rect 121 390 122 391 
rect 124 390 125 391 
rect 121 395 122 396 
rect 124 395 125 396 
<< m2 >>
rect 121 390 122 391 
rect 124 390 125 391 
rect 121 395 122 396 
rect 124 395 125 396 
<< m2c >>
rect 121 390 122 391 
rect 124 390 125 391 
rect 121 395 122 396 
rect 124 395 125 396 
<< labels >>
rlabel pdiffusion 337 246 338 247  0 t = 1
rlabel pdiffusion 340 246 341 247  0 t = 2
rlabel pdiffusion 337 251 338 252  0 t = 3
rlabel pdiffusion 340 251 341 252  0 t = 4
rlabel pdiffusion 336 246 342 252 0 cell no = 459
<< m1 >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< m2 >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< m2c >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< labels >>
rlabel pdiffusion 427 336 428 337  0 t = 1
rlabel pdiffusion 430 336 431 337  0 t = 2
rlabel pdiffusion 427 341 428 342  0 t = 3
rlabel pdiffusion 430 341 431 342  0 t = 4
rlabel pdiffusion 426 336 432 342 0 cell no = 460
<< m1 >>
rect 427 336 428 337 
rect 430 336 431 337 
rect 427 341 428 342 
rect 430 341 431 342 
<< m2 >>
rect 427 336 428 337 
rect 430 336 431 337 
rect 427 341 428 342 
rect 430 341 431 342 
<< m2c >>
rect 427 336 428 337 
rect 430 336 431 337 
rect 427 341 428 342 
rect 430 341 431 342 
<< labels >>
rlabel pdiffusion 193 408 194 409  0 t = 1
rlabel pdiffusion 196 408 197 409  0 t = 2
rlabel pdiffusion 193 413 194 414  0 t = 3
rlabel pdiffusion 196 413 197 414  0 t = 4
rlabel pdiffusion 192 408 198 414 0 cell no = 461
<< m1 >>
rect 193 408 194 409 
rect 196 408 197 409 
rect 193 413 194 414 
rect 196 413 197 414 
<< m2 >>
rect 193 408 194 409 
rect 196 408 197 409 
rect 193 413 194 414 
rect 196 413 197 414 
<< m2c >>
rect 193 408 194 409 
rect 196 408 197 409 
rect 193 413 194 414 
rect 196 413 197 414 
<< labels >>
rlabel pdiffusion 319 282 320 283  0 t = 1
rlabel pdiffusion 322 282 323 283  0 t = 2
rlabel pdiffusion 319 287 320 288  0 t = 3
rlabel pdiffusion 322 287 323 288  0 t = 4
rlabel pdiffusion 318 282 324 288 0 cell no = 462
<< m1 >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< m2 >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< m2c >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< labels >>
rlabel pdiffusion 229 318 230 319  0 t = 1
rlabel pdiffusion 232 318 233 319  0 t = 2
rlabel pdiffusion 229 323 230 324  0 t = 3
rlabel pdiffusion 232 323 233 324  0 t = 4
rlabel pdiffusion 228 318 234 324 0 cell no = 463
<< m1 >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< m2 >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< m2c >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< labels >>
rlabel pdiffusion 193 444 194 445  0 t = 1
rlabel pdiffusion 196 444 197 445  0 t = 2
rlabel pdiffusion 193 449 194 450  0 t = 3
rlabel pdiffusion 196 449 197 450  0 t = 4
rlabel pdiffusion 192 444 198 450 0 cell no = 464
<< m1 >>
rect 193 444 194 445 
rect 196 444 197 445 
rect 193 449 194 450 
rect 196 449 197 450 
<< m2 >>
rect 193 444 194 445 
rect 196 444 197 445 
rect 193 449 194 450 
rect 196 449 197 450 
<< m2c >>
rect 193 444 194 445 
rect 196 444 197 445 
rect 193 449 194 450 
rect 196 449 197 450 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 465
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 247 264 248 265  0 t = 1
rlabel pdiffusion 250 264 251 265  0 t = 2
rlabel pdiffusion 247 269 248 270  0 t = 3
rlabel pdiffusion 250 269 251 270  0 t = 4
rlabel pdiffusion 246 264 252 270 0 cell no = 466
<< m1 >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< m2 >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< m2c >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< labels >>
rlabel pdiffusion 49 372 50 373  0 t = 1
rlabel pdiffusion 52 372 53 373  0 t = 2
rlabel pdiffusion 49 377 50 378  0 t = 3
rlabel pdiffusion 52 377 53 378  0 t = 4
rlabel pdiffusion 48 372 54 378 0 cell no = 467
<< m1 >>
rect 49 372 50 373 
rect 52 372 53 373 
rect 49 377 50 378 
rect 52 377 53 378 
<< m2 >>
rect 49 372 50 373 
rect 52 372 53 373 
rect 49 377 50 378 
rect 52 377 53 378 
<< m2c >>
rect 49 372 50 373 
rect 52 372 53 373 
rect 49 377 50 378 
rect 52 377 53 378 
<< labels >>
rlabel pdiffusion 247 354 248 355  0 t = 1
rlabel pdiffusion 250 354 251 355  0 t = 2
rlabel pdiffusion 247 359 248 360  0 t = 3
rlabel pdiffusion 250 359 251 360  0 t = 4
rlabel pdiffusion 246 354 252 360 0 cell no = 468
<< m1 >>
rect 247 354 248 355 
rect 250 354 251 355 
rect 247 359 248 360 
rect 250 359 251 360 
<< m2 >>
rect 247 354 248 355 
rect 250 354 251 355 
rect 247 359 248 360 
rect 250 359 251 360 
<< m2c >>
rect 247 354 248 355 
rect 250 354 251 355 
rect 247 359 248 360 
rect 250 359 251 360 
<< labels >>
rlabel pdiffusion 409 408 410 409  0 t = 1
rlabel pdiffusion 412 408 413 409  0 t = 2
rlabel pdiffusion 409 413 410 414  0 t = 3
rlabel pdiffusion 412 413 413 414  0 t = 4
rlabel pdiffusion 408 408 414 414 0 cell no = 469
<< m1 >>
rect 409 408 410 409 
rect 412 408 413 409 
rect 409 413 410 414 
rect 412 413 413 414 
<< m2 >>
rect 409 408 410 409 
rect 412 408 413 409 
rect 409 413 410 414 
rect 412 413 413 414 
<< m2c >>
rect 409 408 410 409 
rect 412 408 413 409 
rect 409 413 410 414 
rect 412 413 413 414 
<< labels >>
rlabel pdiffusion 301 426 302 427  0 t = 1
rlabel pdiffusion 304 426 305 427  0 t = 2
rlabel pdiffusion 301 431 302 432  0 t = 3
rlabel pdiffusion 304 431 305 432  0 t = 4
rlabel pdiffusion 300 426 306 432 0 cell no = 470
<< m1 >>
rect 301 426 302 427 
rect 304 426 305 427 
rect 301 431 302 432 
rect 304 431 305 432 
<< m2 >>
rect 301 426 302 427 
rect 304 426 305 427 
rect 301 431 302 432 
rect 304 431 305 432 
<< m2c >>
rect 301 426 302 427 
rect 304 426 305 427 
rect 301 431 302 432 
rect 304 431 305 432 
<< labels >>
rlabel pdiffusion 355 282 356 283  0 t = 1
rlabel pdiffusion 358 282 359 283  0 t = 2
rlabel pdiffusion 355 287 356 288  0 t = 3
rlabel pdiffusion 358 287 359 288  0 t = 4
rlabel pdiffusion 354 282 360 288 0 cell no = 471
<< m1 >>
rect 355 282 356 283 
rect 358 282 359 283 
rect 355 287 356 288 
rect 358 287 359 288 
<< m2 >>
rect 355 282 356 283 
rect 358 282 359 283 
rect 355 287 356 288 
rect 358 287 359 288 
<< m2c >>
rect 355 282 356 283 
rect 358 282 359 283 
rect 355 287 356 288 
rect 358 287 359 288 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 472
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 247 282 248 283  0 t = 1
rlabel pdiffusion 250 282 251 283  0 t = 2
rlabel pdiffusion 247 287 248 288  0 t = 3
rlabel pdiffusion 250 287 251 288  0 t = 4
rlabel pdiffusion 246 282 252 288 0 cell no = 473
<< m1 >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< m2 >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< m2c >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< labels >>
rlabel pdiffusion 103 138 104 139  0 t = 1
rlabel pdiffusion 106 138 107 139  0 t = 2
rlabel pdiffusion 103 143 104 144  0 t = 3
rlabel pdiffusion 106 143 107 144  0 t = 4
rlabel pdiffusion 102 138 108 144 0 cell no = 474
<< m1 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2c >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< labels >>
rlabel pdiffusion 373 444 374 445  0 t = 1
rlabel pdiffusion 376 444 377 445  0 t = 2
rlabel pdiffusion 373 449 374 450  0 t = 3
rlabel pdiffusion 376 449 377 450  0 t = 4
rlabel pdiffusion 372 444 378 450 0 cell no = 475
<< m1 >>
rect 373 444 374 445 
rect 376 444 377 445 
rect 373 449 374 450 
rect 376 449 377 450 
<< m2 >>
rect 373 444 374 445 
rect 376 444 377 445 
rect 373 449 374 450 
rect 376 449 377 450 
<< m2c >>
rect 373 444 374 445 
rect 376 444 377 445 
rect 373 449 374 450 
rect 376 449 377 450 
<< labels >>
rlabel pdiffusion 175 264 176 265  0 t = 1
rlabel pdiffusion 178 264 179 265  0 t = 2
rlabel pdiffusion 175 269 176 270  0 t = 3
rlabel pdiffusion 178 269 179 270  0 t = 4
rlabel pdiffusion 174 264 180 270 0 cell no = 476
<< m1 >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< m2 >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< m2c >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< labels >>
rlabel pdiffusion 409 84 410 85  0 t = 1
rlabel pdiffusion 412 84 413 85  0 t = 2
rlabel pdiffusion 409 89 410 90  0 t = 3
rlabel pdiffusion 412 89 413 90  0 t = 4
rlabel pdiffusion 408 84 414 90 0 cell no = 477
<< m1 >>
rect 409 84 410 85 
rect 412 84 413 85 
rect 409 89 410 90 
rect 412 89 413 90 
<< m2 >>
rect 409 84 410 85 
rect 412 84 413 85 
rect 409 89 410 90 
rect 412 89 413 90 
<< m2c >>
rect 409 84 410 85 
rect 412 84 413 85 
rect 409 89 410 90 
rect 412 89 413 90 
<< labels >>
rlabel pdiffusion 31 318 32 319  0 t = 1
rlabel pdiffusion 34 318 35 319  0 t = 2
rlabel pdiffusion 31 323 32 324  0 t = 3
rlabel pdiffusion 34 323 35 324  0 t = 4
rlabel pdiffusion 30 318 36 324 0 cell no = 478
<< m1 >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< m2 >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< m2c >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< labels >>
rlabel pdiffusion 49 390 50 391  0 t = 1
rlabel pdiffusion 52 390 53 391  0 t = 2
rlabel pdiffusion 49 395 50 396  0 t = 3
rlabel pdiffusion 52 395 53 396  0 t = 4
rlabel pdiffusion 48 390 54 396 0 cell no = 479
<< m1 >>
rect 49 390 50 391 
rect 52 390 53 391 
rect 49 395 50 396 
rect 52 395 53 396 
<< m2 >>
rect 49 390 50 391 
rect 52 390 53 391 
rect 49 395 50 396 
rect 52 395 53 396 
<< m2c >>
rect 49 390 50 391 
rect 52 390 53 391 
rect 49 395 50 396 
rect 52 395 53 396 
<< labels >>
rlabel pdiffusion 175 300 176 301  0 t = 1
rlabel pdiffusion 178 300 179 301  0 t = 2
rlabel pdiffusion 175 305 176 306  0 t = 3
rlabel pdiffusion 178 305 179 306  0 t = 4
rlabel pdiffusion 174 300 180 306 0 cell no = 480
<< m1 >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< m2 >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< m2c >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< labels >>
rlabel pdiffusion 49 354 50 355  0 t = 1
rlabel pdiffusion 52 354 53 355  0 t = 2
rlabel pdiffusion 49 359 50 360  0 t = 3
rlabel pdiffusion 52 359 53 360  0 t = 4
rlabel pdiffusion 48 354 54 360 0 cell no = 481
<< m1 >>
rect 49 354 50 355 
rect 52 354 53 355 
rect 49 359 50 360 
rect 52 359 53 360 
<< m2 >>
rect 49 354 50 355 
rect 52 354 53 355 
rect 49 359 50 360 
rect 52 359 53 360 
<< m2c >>
rect 49 354 50 355 
rect 52 354 53 355 
rect 49 359 50 360 
rect 52 359 53 360 
<< labels >>
rlabel pdiffusion 157 372 158 373  0 t = 1
rlabel pdiffusion 160 372 161 373  0 t = 2
rlabel pdiffusion 157 377 158 378  0 t = 3
rlabel pdiffusion 160 377 161 378  0 t = 4
rlabel pdiffusion 156 372 162 378 0 cell no = 482
<< m1 >>
rect 157 372 158 373 
rect 160 372 161 373 
rect 157 377 158 378 
rect 160 377 161 378 
<< m2 >>
rect 157 372 158 373 
rect 160 372 161 373 
rect 157 377 158 378 
rect 160 377 161 378 
<< m2c >>
rect 157 372 158 373 
rect 160 372 161 373 
rect 157 377 158 378 
rect 160 377 161 378 
<< labels >>
rlabel pdiffusion 301 282 302 283  0 t = 1
rlabel pdiffusion 304 282 305 283  0 t = 2
rlabel pdiffusion 301 287 302 288  0 t = 3
rlabel pdiffusion 304 287 305 288  0 t = 4
rlabel pdiffusion 300 282 306 288 0 cell no = 483
<< m1 >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< m2 >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< m2c >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< labels >>
rlabel pdiffusion 139 372 140 373  0 t = 1
rlabel pdiffusion 142 372 143 373  0 t = 2
rlabel pdiffusion 139 377 140 378  0 t = 3
rlabel pdiffusion 142 377 143 378  0 t = 4
rlabel pdiffusion 138 372 144 378 0 cell no = 484
<< m1 >>
rect 139 372 140 373 
rect 142 372 143 373 
rect 139 377 140 378 
rect 142 377 143 378 
<< m2 >>
rect 139 372 140 373 
rect 142 372 143 373 
rect 139 377 140 378 
rect 142 377 143 378 
<< m2c >>
rect 139 372 140 373 
rect 142 372 143 373 
rect 139 377 140 378 
rect 142 377 143 378 
<< labels >>
rlabel pdiffusion 13 354 14 355  0 t = 1
rlabel pdiffusion 16 354 17 355  0 t = 2
rlabel pdiffusion 13 359 14 360  0 t = 3
rlabel pdiffusion 16 359 17 360  0 t = 4
rlabel pdiffusion 12 354 18 360 0 cell no = 485
<< m1 >>
rect 13 354 14 355 
rect 16 354 17 355 
rect 13 359 14 360 
rect 16 359 17 360 
<< m2 >>
rect 13 354 14 355 
rect 16 354 17 355 
rect 13 359 14 360 
rect 16 359 17 360 
<< m2c >>
rect 13 354 14 355 
rect 16 354 17 355 
rect 13 359 14 360 
rect 16 359 17 360 
<< labels >>
rlabel pdiffusion 193 390 194 391  0 t = 1
rlabel pdiffusion 196 390 197 391  0 t = 2
rlabel pdiffusion 193 395 194 396  0 t = 3
rlabel pdiffusion 196 395 197 396  0 t = 4
rlabel pdiffusion 192 390 198 396 0 cell no = 486
<< m1 >>
rect 193 390 194 391 
rect 196 390 197 391 
rect 193 395 194 396 
rect 196 395 197 396 
<< m2 >>
rect 193 390 194 391 
rect 196 390 197 391 
rect 193 395 194 396 
rect 196 395 197 396 
<< m2c >>
rect 193 390 194 391 
rect 196 390 197 391 
rect 193 395 194 396 
rect 196 395 197 396 
<< labels >>
rlabel pdiffusion 301 318 302 319  0 t = 1
rlabel pdiffusion 304 318 305 319  0 t = 2
rlabel pdiffusion 301 323 302 324  0 t = 3
rlabel pdiffusion 304 323 305 324  0 t = 4
rlabel pdiffusion 300 318 306 324 0 cell no = 487
<< m1 >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< m2 >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< m2c >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< labels >>
rlabel pdiffusion 121 354 122 355  0 t = 1
rlabel pdiffusion 124 354 125 355  0 t = 2
rlabel pdiffusion 121 359 122 360  0 t = 3
rlabel pdiffusion 124 359 125 360  0 t = 4
rlabel pdiffusion 120 354 126 360 0 cell no = 488
<< m1 >>
rect 121 354 122 355 
rect 124 354 125 355 
rect 121 359 122 360 
rect 124 359 125 360 
<< m2 >>
rect 121 354 122 355 
rect 124 354 125 355 
rect 121 359 122 360 
rect 124 359 125 360 
<< m2c >>
rect 121 354 122 355 
rect 124 354 125 355 
rect 121 359 122 360 
rect 124 359 125 360 
<< labels >>
rlabel pdiffusion 139 192 140 193  0 t = 1
rlabel pdiffusion 142 192 143 193  0 t = 2
rlabel pdiffusion 139 197 140 198  0 t = 3
rlabel pdiffusion 142 197 143 198  0 t = 4
rlabel pdiffusion 138 192 144 198 0 cell no = 489
<< m1 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2c >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< labels >>
rlabel pdiffusion 175 390 176 391  0 t = 1
rlabel pdiffusion 178 390 179 391  0 t = 2
rlabel pdiffusion 175 395 176 396  0 t = 3
rlabel pdiffusion 178 395 179 396  0 t = 4
rlabel pdiffusion 174 390 180 396 0 cell no = 490
<< m1 >>
rect 175 390 176 391 
rect 178 390 179 391 
rect 175 395 176 396 
rect 178 395 179 396 
<< m2 >>
rect 175 390 176 391 
rect 178 390 179 391 
rect 175 395 176 396 
rect 178 395 179 396 
<< m2c >>
rect 175 390 176 391 
rect 178 390 179 391 
rect 175 395 176 396 
rect 178 395 179 396 
<< labels >>
rlabel pdiffusion 121 192 122 193  0 t = 1
rlabel pdiffusion 124 192 125 193  0 t = 2
rlabel pdiffusion 121 197 122 198  0 t = 3
rlabel pdiffusion 124 197 125 198  0 t = 4
rlabel pdiffusion 120 192 126 198 0 cell no = 491
<< m1 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2c >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< labels >>
rlabel pdiffusion 337 444 338 445  0 t = 1
rlabel pdiffusion 340 444 341 445  0 t = 2
rlabel pdiffusion 337 449 338 450  0 t = 3
rlabel pdiffusion 340 449 341 450  0 t = 4
rlabel pdiffusion 336 444 342 450 0 cell no = 492
<< m1 >>
rect 337 444 338 445 
rect 340 444 341 445 
rect 337 449 338 450 
rect 340 449 341 450 
<< m2 >>
rect 337 444 338 445 
rect 340 444 341 445 
rect 337 449 338 450 
rect 340 449 341 450 
<< m2c >>
rect 337 444 338 445 
rect 340 444 341 445 
rect 337 449 338 450 
rect 340 449 341 450 
<< labels >>
rlabel pdiffusion 85 372 86 373  0 t = 1
rlabel pdiffusion 88 372 89 373  0 t = 2
rlabel pdiffusion 85 377 86 378  0 t = 3
rlabel pdiffusion 88 377 89 378  0 t = 4
rlabel pdiffusion 84 372 90 378 0 cell no = 493
<< m1 >>
rect 85 372 86 373 
rect 88 372 89 373 
rect 85 377 86 378 
rect 88 377 89 378 
<< m2 >>
rect 85 372 86 373 
rect 88 372 89 373 
rect 85 377 86 378 
rect 88 377 89 378 
<< m2c >>
rect 85 372 86 373 
rect 88 372 89 373 
rect 85 377 86 378 
rect 88 377 89 378 
<< labels >>
rlabel pdiffusion 355 444 356 445  0 t = 1
rlabel pdiffusion 358 444 359 445  0 t = 2
rlabel pdiffusion 355 449 356 450  0 t = 3
rlabel pdiffusion 358 449 359 450  0 t = 4
rlabel pdiffusion 354 444 360 450 0 cell no = 494
<< m1 >>
rect 355 444 356 445 
rect 358 444 359 445 
rect 355 449 356 450 
rect 358 449 359 450 
<< m2 >>
rect 355 444 356 445 
rect 358 444 359 445 
rect 355 449 356 450 
rect 358 449 359 450 
<< m2c >>
rect 355 444 356 445 
rect 358 444 359 445 
rect 355 449 356 450 
rect 358 449 359 450 
<< labels >>
rlabel pdiffusion 229 300 230 301  0 t = 1
rlabel pdiffusion 232 300 233 301  0 t = 2
rlabel pdiffusion 229 305 230 306  0 t = 3
rlabel pdiffusion 232 305 233 306  0 t = 4
rlabel pdiffusion 228 300 234 306 0 cell no = 495
<< m1 >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< m2 >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< m2c >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< labels >>
rlabel pdiffusion 409 210 410 211  0 t = 1
rlabel pdiffusion 412 210 413 211  0 t = 2
rlabel pdiffusion 409 215 410 216  0 t = 3
rlabel pdiffusion 412 215 413 216  0 t = 4
rlabel pdiffusion 408 210 414 216 0 cell no = 496
<< m1 >>
rect 409 210 410 211 
rect 412 210 413 211 
rect 409 215 410 216 
rect 412 215 413 216 
<< m2 >>
rect 409 210 410 211 
rect 412 210 413 211 
rect 409 215 410 216 
rect 412 215 413 216 
<< m2c >>
rect 409 210 410 211 
rect 412 210 413 211 
rect 409 215 410 216 
rect 412 215 413 216 
<< labels >>
rlabel pdiffusion 409 390 410 391  0 t = 1
rlabel pdiffusion 412 390 413 391  0 t = 2
rlabel pdiffusion 409 395 410 396  0 t = 3
rlabel pdiffusion 412 395 413 396  0 t = 4
rlabel pdiffusion 408 390 414 396 0 cell no = 497
<< m1 >>
rect 409 390 410 391 
rect 412 390 413 391 
rect 409 395 410 396 
rect 412 395 413 396 
<< m2 >>
rect 409 390 410 391 
rect 412 390 413 391 
rect 409 395 410 396 
rect 412 395 413 396 
<< m2c >>
rect 409 390 410 391 
rect 412 390 413 391 
rect 409 395 410 396 
rect 412 395 413 396 
<< labels >>
rlabel pdiffusion 265 228 266 229  0 t = 1
rlabel pdiffusion 268 228 269 229  0 t = 2
rlabel pdiffusion 265 233 266 234  0 t = 3
rlabel pdiffusion 268 233 269 234  0 t = 4
rlabel pdiffusion 264 228 270 234 0 cell no = 498
<< m1 >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< m2 >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< m2c >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< labels >>
rlabel pdiffusion 445 390 446 391  0 t = 1
rlabel pdiffusion 448 390 449 391  0 t = 2
rlabel pdiffusion 445 395 446 396  0 t = 3
rlabel pdiffusion 448 395 449 396  0 t = 4
rlabel pdiffusion 444 390 450 396 0 cell no = 499
<< m1 >>
rect 445 390 446 391 
rect 448 390 449 391 
rect 445 395 446 396 
rect 448 395 449 396 
<< m2 >>
rect 445 390 446 391 
rect 448 390 449 391 
rect 445 395 446 396 
rect 448 395 449 396 
<< m2c >>
rect 445 390 446 391 
rect 448 390 449 391 
rect 445 395 446 396 
rect 448 395 449 396 
<< labels >>
rlabel pdiffusion 211 174 212 175  0 t = 1
rlabel pdiffusion 214 174 215 175  0 t = 2
rlabel pdiffusion 211 179 212 180  0 t = 3
rlabel pdiffusion 214 179 215 180  0 t = 4
rlabel pdiffusion 210 174 216 180 0 cell no = 500
<< m1 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2c >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< labels >>
rlabel pdiffusion 319 444 320 445  0 t = 1
rlabel pdiffusion 322 444 323 445  0 t = 2
rlabel pdiffusion 319 449 320 450  0 t = 3
rlabel pdiffusion 322 449 323 450  0 t = 4
rlabel pdiffusion 318 444 324 450 0 cell no = 501
<< m1 >>
rect 319 444 320 445 
rect 322 444 323 445 
rect 319 449 320 450 
rect 322 449 323 450 
<< m2 >>
rect 319 444 320 445 
rect 322 444 323 445 
rect 319 449 320 450 
rect 322 449 323 450 
<< m2c >>
rect 319 444 320 445 
rect 322 444 323 445 
rect 319 449 320 450 
rect 322 449 323 450 
<< labels >>
rlabel pdiffusion 13 426 14 427  0 t = 1
rlabel pdiffusion 16 426 17 427  0 t = 2
rlabel pdiffusion 13 431 14 432  0 t = 3
rlabel pdiffusion 16 431 17 432  0 t = 4
rlabel pdiffusion 12 426 18 432 0 cell no = 502
<< m1 >>
rect 13 426 14 427 
rect 16 426 17 427 
rect 13 431 14 432 
rect 16 431 17 432 
<< m2 >>
rect 13 426 14 427 
rect 16 426 17 427 
rect 13 431 14 432 
rect 16 431 17 432 
<< m2c >>
rect 13 426 14 427 
rect 16 426 17 427 
rect 13 431 14 432 
rect 16 431 17 432 
<< labels >>
rlabel pdiffusion 13 390 14 391  0 t = 1
rlabel pdiffusion 16 390 17 391  0 t = 2
rlabel pdiffusion 13 395 14 396  0 t = 3
rlabel pdiffusion 16 395 17 396  0 t = 4
rlabel pdiffusion 12 390 18 396 0 cell no = 503
<< m1 >>
rect 13 390 14 391 
rect 16 390 17 391 
rect 13 395 14 396 
rect 16 395 17 396 
<< m2 >>
rect 13 390 14 391 
rect 16 390 17 391 
rect 13 395 14 396 
rect 16 395 17 396 
<< m2c >>
rect 13 390 14 391 
rect 16 390 17 391 
rect 13 395 14 396 
rect 16 395 17 396 
<< labels >>
rlabel pdiffusion 139 318 140 319  0 t = 1
rlabel pdiffusion 142 318 143 319  0 t = 2
rlabel pdiffusion 139 323 140 324  0 t = 3
rlabel pdiffusion 142 323 143 324  0 t = 4
rlabel pdiffusion 138 318 144 324 0 cell no = 504
<< m1 >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< m2 >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< m2c >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< labels >>
rlabel pdiffusion 193 264 194 265  0 t = 1
rlabel pdiffusion 196 264 197 265  0 t = 2
rlabel pdiffusion 193 269 194 270  0 t = 3
rlabel pdiffusion 196 269 197 270  0 t = 4
rlabel pdiffusion 192 264 198 270 0 cell no = 505
<< m1 >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< m2 >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< m2c >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< labels >>
rlabel pdiffusion 49 318 50 319  0 t = 1
rlabel pdiffusion 52 318 53 319  0 t = 2
rlabel pdiffusion 49 323 50 324  0 t = 3
rlabel pdiffusion 52 323 53 324  0 t = 4
rlabel pdiffusion 48 318 54 324 0 cell no = 506
<< m1 >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< m2 >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< m2c >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< labels >>
rlabel pdiffusion 265 372 266 373  0 t = 1
rlabel pdiffusion 268 372 269 373  0 t = 2
rlabel pdiffusion 265 377 266 378  0 t = 3
rlabel pdiffusion 268 377 269 378  0 t = 4
rlabel pdiffusion 264 372 270 378 0 cell no = 507
<< m1 >>
rect 265 372 266 373 
rect 268 372 269 373 
rect 265 377 266 378 
rect 268 377 269 378 
<< m2 >>
rect 265 372 266 373 
rect 268 372 269 373 
rect 265 377 266 378 
rect 268 377 269 378 
<< m2c >>
rect 265 372 266 373 
rect 268 372 269 373 
rect 265 377 266 378 
rect 268 377 269 378 
<< labels >>
rlabel pdiffusion 175 282 176 283  0 t = 1
rlabel pdiffusion 178 282 179 283  0 t = 2
rlabel pdiffusion 175 287 176 288  0 t = 3
rlabel pdiffusion 178 287 179 288  0 t = 4
rlabel pdiffusion 174 282 180 288 0 cell no = 508
<< m1 >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< m2 >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< m2c >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< labels >>
rlabel pdiffusion 355 192 356 193  0 t = 1
rlabel pdiffusion 358 192 359 193  0 t = 2
rlabel pdiffusion 355 197 356 198  0 t = 3
rlabel pdiffusion 358 197 359 198  0 t = 4
rlabel pdiffusion 354 192 360 198 0 cell no = 509
<< m1 >>
rect 355 192 356 193 
rect 358 192 359 193 
rect 355 197 356 198 
rect 358 197 359 198 
<< m2 >>
rect 355 192 356 193 
rect 358 192 359 193 
rect 355 197 356 198 
rect 358 197 359 198 
<< m2c >>
rect 355 192 356 193 
rect 358 192 359 193 
rect 355 197 356 198 
rect 358 197 359 198 
<< labels >>
rlabel pdiffusion 157 300 158 301  0 t = 1
rlabel pdiffusion 160 300 161 301  0 t = 2
rlabel pdiffusion 157 305 158 306  0 t = 3
rlabel pdiffusion 160 305 161 306  0 t = 4
rlabel pdiffusion 156 300 162 306 0 cell no = 510
<< m1 >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< m2 >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< m2c >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< labels >>
rlabel pdiffusion 427 120 428 121  0 t = 1
rlabel pdiffusion 430 120 431 121  0 t = 2
rlabel pdiffusion 427 125 428 126  0 t = 3
rlabel pdiffusion 430 125 431 126  0 t = 4
rlabel pdiffusion 426 120 432 126 0 cell no = 511
<< m1 >>
rect 427 120 428 121 
rect 430 120 431 121 
rect 427 125 428 126 
rect 430 125 431 126 
<< m2 >>
rect 427 120 428 121 
rect 430 120 431 121 
rect 427 125 428 126 
rect 430 125 431 126 
<< m2c >>
rect 427 120 428 121 
rect 430 120 431 121 
rect 427 125 428 126 
rect 430 125 431 126 
<< labels >>
rlabel pdiffusion 355 138 356 139  0 t = 1
rlabel pdiffusion 358 138 359 139  0 t = 2
rlabel pdiffusion 355 143 356 144  0 t = 3
rlabel pdiffusion 358 143 359 144  0 t = 4
rlabel pdiffusion 354 138 360 144 0 cell no = 512
<< m1 >>
rect 355 138 356 139 
rect 358 138 359 139 
rect 355 143 356 144 
rect 358 143 359 144 
<< m2 >>
rect 355 138 356 139 
rect 358 138 359 139 
rect 355 143 356 144 
rect 358 143 359 144 
<< m2c >>
rect 355 138 356 139 
rect 358 138 359 139 
rect 355 143 356 144 
rect 358 143 359 144 
<< labels >>
rlabel pdiffusion 229 372 230 373  0 t = 1
rlabel pdiffusion 232 372 233 373  0 t = 2
rlabel pdiffusion 229 377 230 378  0 t = 3
rlabel pdiffusion 232 377 233 378  0 t = 4
rlabel pdiffusion 228 372 234 378 0 cell no = 513
<< m1 >>
rect 229 372 230 373 
rect 232 372 233 373 
rect 229 377 230 378 
rect 232 377 233 378 
<< m2 >>
rect 229 372 230 373 
rect 232 372 233 373 
rect 229 377 230 378 
rect 232 377 233 378 
<< m2c >>
rect 229 372 230 373 
rect 232 372 233 373 
rect 229 377 230 378 
rect 232 377 233 378 
<< labels >>
rlabel pdiffusion 175 354 176 355  0 t = 1
rlabel pdiffusion 178 354 179 355  0 t = 2
rlabel pdiffusion 175 359 176 360  0 t = 3
rlabel pdiffusion 178 359 179 360  0 t = 4
rlabel pdiffusion 174 354 180 360 0 cell no = 514
<< m1 >>
rect 175 354 176 355 
rect 178 354 179 355 
rect 175 359 176 360 
rect 178 359 179 360 
<< m2 >>
rect 175 354 176 355 
rect 178 354 179 355 
rect 175 359 176 360 
rect 178 359 179 360 
<< m2c >>
rect 175 354 176 355 
rect 178 354 179 355 
rect 175 359 176 360 
rect 178 359 179 360 
<< labels >>
rlabel pdiffusion 85 318 86 319  0 t = 1
rlabel pdiffusion 88 318 89 319  0 t = 2
rlabel pdiffusion 85 323 86 324  0 t = 3
rlabel pdiffusion 88 323 89 324  0 t = 4
rlabel pdiffusion 84 318 90 324 0 cell no = 515
<< m1 >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< m2 >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< m2c >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< labels >>
rlabel pdiffusion 409 426 410 427  0 t = 1
rlabel pdiffusion 412 426 413 427  0 t = 2
rlabel pdiffusion 409 431 410 432  0 t = 3
rlabel pdiffusion 412 431 413 432  0 t = 4
rlabel pdiffusion 408 426 414 432 0 cell no = 516
<< m1 >>
rect 409 426 410 427 
rect 412 426 413 427 
rect 409 431 410 432 
rect 412 431 413 432 
<< m2 >>
rect 409 426 410 427 
rect 412 426 413 427 
rect 409 431 410 432 
rect 412 431 413 432 
<< m2c >>
rect 409 426 410 427 
rect 412 426 413 427 
rect 409 431 410 432 
rect 412 431 413 432 
<< labels >>
rlabel pdiffusion 355 408 356 409  0 t = 1
rlabel pdiffusion 358 408 359 409  0 t = 2
rlabel pdiffusion 355 413 356 414  0 t = 3
rlabel pdiffusion 358 413 359 414  0 t = 4
rlabel pdiffusion 354 408 360 414 0 cell no = 517
<< m1 >>
rect 355 408 356 409 
rect 358 408 359 409 
rect 355 413 356 414 
rect 358 413 359 414 
<< m2 >>
rect 355 408 356 409 
rect 358 408 359 409 
rect 355 413 356 414 
rect 358 413 359 414 
<< m2c >>
rect 355 408 356 409 
rect 358 408 359 409 
rect 355 413 356 414 
rect 358 413 359 414 
<< labels >>
rlabel pdiffusion 337 192 338 193  0 t = 1
rlabel pdiffusion 340 192 341 193  0 t = 2
rlabel pdiffusion 337 197 338 198  0 t = 3
rlabel pdiffusion 340 197 341 198  0 t = 4
rlabel pdiffusion 336 192 342 198 0 cell no = 518
<< m1 >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< m2 >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< m2c >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< labels >>
rlabel pdiffusion 427 426 428 427  0 t = 1
rlabel pdiffusion 430 426 431 427  0 t = 2
rlabel pdiffusion 427 431 428 432  0 t = 3
rlabel pdiffusion 430 431 431 432  0 t = 4
rlabel pdiffusion 426 426 432 432 0 cell no = 519
<< m1 >>
rect 427 426 428 427 
rect 430 426 431 427 
rect 427 431 428 432 
rect 430 431 431 432 
<< m2 >>
rect 427 426 428 427 
rect 430 426 431 427 
rect 427 431 428 432 
rect 430 431 431 432 
<< m2c >>
rect 427 426 428 427 
rect 430 426 431 427 
rect 427 431 428 432 
rect 430 431 431 432 
<< labels >>
rlabel pdiffusion 391 444 392 445  0 t = 1
rlabel pdiffusion 394 444 395 445  0 t = 2
rlabel pdiffusion 391 449 392 450  0 t = 3
rlabel pdiffusion 394 449 395 450  0 t = 4
rlabel pdiffusion 390 444 396 450 0 cell no = 520
<< m1 >>
rect 391 444 392 445 
rect 394 444 395 445 
rect 391 449 392 450 
rect 394 449 395 450 
<< m2 >>
rect 391 444 392 445 
rect 394 444 395 445 
rect 391 449 392 450 
rect 394 449 395 450 
<< m2c >>
rect 391 444 392 445 
rect 394 444 395 445 
rect 391 449 392 450 
rect 394 449 395 450 
<< labels >>
rlabel pdiffusion 427 408 428 409  0 t = 1
rlabel pdiffusion 430 408 431 409  0 t = 2
rlabel pdiffusion 427 413 428 414  0 t = 3
rlabel pdiffusion 430 413 431 414  0 t = 4
rlabel pdiffusion 426 408 432 414 0 cell no = 521
<< m1 >>
rect 427 408 428 409 
rect 430 408 431 409 
rect 427 413 428 414 
rect 430 413 431 414 
<< m2 >>
rect 427 408 428 409 
rect 430 408 431 409 
rect 427 413 428 414 
rect 430 413 431 414 
<< m2c >>
rect 427 408 428 409 
rect 430 408 431 409 
rect 427 413 428 414 
rect 430 413 431 414 
<< labels >>
rlabel pdiffusion 409 444 410 445  0 t = 1
rlabel pdiffusion 412 444 413 445  0 t = 2
rlabel pdiffusion 409 449 410 450  0 t = 3
rlabel pdiffusion 412 449 413 450  0 t = 4
rlabel pdiffusion 408 444 414 450 0 cell no = 522
<< m1 >>
rect 409 444 410 445 
rect 412 444 413 445 
rect 409 449 410 450 
rect 412 449 413 450 
<< m2 >>
rect 409 444 410 445 
rect 412 444 413 445 
rect 409 449 410 450 
rect 412 449 413 450 
<< m2c >>
rect 409 444 410 445 
rect 412 444 413 445 
rect 409 449 410 450 
rect 412 449 413 450 
<< labels >>
rlabel pdiffusion 211 354 212 355  0 t = 1
rlabel pdiffusion 214 354 215 355  0 t = 2
rlabel pdiffusion 211 359 212 360  0 t = 3
rlabel pdiffusion 214 359 215 360  0 t = 4
rlabel pdiffusion 210 354 216 360 0 cell no = 523
<< m1 >>
rect 211 354 212 355 
rect 214 354 215 355 
rect 211 359 212 360 
rect 214 359 215 360 
<< m2 >>
rect 211 354 212 355 
rect 214 354 215 355 
rect 211 359 212 360 
rect 214 359 215 360 
<< m2c >>
rect 211 354 212 355 
rect 214 354 215 355 
rect 211 359 212 360 
rect 214 359 215 360 
<< labels >>
rlabel pdiffusion 265 246 266 247  0 t = 1
rlabel pdiffusion 268 246 269 247  0 t = 2
rlabel pdiffusion 265 251 266 252  0 t = 3
rlabel pdiffusion 268 251 269 252  0 t = 4
rlabel pdiffusion 264 246 270 252 0 cell no = 524
<< m1 >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< m2 >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< m2c >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< labels >>
rlabel pdiffusion 337 390 338 391  0 t = 1
rlabel pdiffusion 340 390 341 391  0 t = 2
rlabel pdiffusion 337 395 338 396  0 t = 3
rlabel pdiffusion 340 395 341 396  0 t = 4
rlabel pdiffusion 336 390 342 396 0 cell no = 525
<< m1 >>
rect 337 390 338 391 
rect 340 390 341 391 
rect 337 395 338 396 
rect 340 395 341 396 
<< m2 >>
rect 337 390 338 391 
rect 340 390 341 391 
rect 337 395 338 396 
rect 340 395 341 396 
<< m2c >>
rect 337 390 338 391 
rect 340 390 341 391 
rect 337 395 338 396 
rect 340 395 341 396 
<< labels >>
rlabel pdiffusion 49 444 50 445  0 t = 1
rlabel pdiffusion 52 444 53 445  0 t = 2
rlabel pdiffusion 49 449 50 450  0 t = 3
rlabel pdiffusion 52 449 53 450  0 t = 4
rlabel pdiffusion 48 444 54 450 0 cell no = 526
<< m1 >>
rect 49 444 50 445 
rect 52 444 53 445 
rect 49 449 50 450 
rect 52 449 53 450 
<< m2 >>
rect 49 444 50 445 
rect 52 444 53 445 
rect 49 449 50 450 
rect 52 449 53 450 
<< m2c >>
rect 49 444 50 445 
rect 52 444 53 445 
rect 49 449 50 450 
rect 52 449 53 450 
<< labels >>
rlabel pdiffusion 85 426 86 427  0 t = 1
rlabel pdiffusion 88 426 89 427  0 t = 2
rlabel pdiffusion 85 431 86 432  0 t = 3
rlabel pdiffusion 88 431 89 432  0 t = 4
rlabel pdiffusion 84 426 90 432 0 cell no = 527
<< m1 >>
rect 85 426 86 427 
rect 88 426 89 427 
rect 85 431 86 432 
rect 88 431 89 432 
<< m2 >>
rect 85 426 86 427 
rect 88 426 89 427 
rect 85 431 86 432 
rect 88 431 89 432 
<< m2c >>
rect 85 426 86 427 
rect 88 426 89 427 
rect 85 431 86 432 
rect 88 431 89 432 
<< labels >>
rlabel pdiffusion 193 156 194 157  0 t = 1
rlabel pdiffusion 196 156 197 157  0 t = 2
rlabel pdiffusion 193 161 194 162  0 t = 3
rlabel pdiffusion 196 161 197 162  0 t = 4
rlabel pdiffusion 192 156 198 162 0 cell no = 528
<< m1 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2c >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< labels >>
rlabel pdiffusion 301 174 302 175  0 t = 1
rlabel pdiffusion 304 174 305 175  0 t = 2
rlabel pdiffusion 301 179 302 180  0 t = 3
rlabel pdiffusion 304 179 305 180  0 t = 4
rlabel pdiffusion 300 174 306 180 0 cell no = 529
<< m1 >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< m2 >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< m2c >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< labels >>
rlabel pdiffusion 211 426 212 427  0 t = 1
rlabel pdiffusion 214 426 215 427  0 t = 2
rlabel pdiffusion 211 431 212 432  0 t = 3
rlabel pdiffusion 214 431 215 432  0 t = 4
rlabel pdiffusion 210 426 216 432 0 cell no = 530
<< m1 >>
rect 211 426 212 427 
rect 214 426 215 427 
rect 211 431 212 432 
rect 214 431 215 432 
<< m2 >>
rect 211 426 212 427 
rect 214 426 215 427 
rect 211 431 212 432 
rect 214 431 215 432 
<< m2c >>
rect 211 426 212 427 
rect 214 426 215 427 
rect 211 431 212 432 
rect 214 431 215 432 
<< labels >>
rlabel pdiffusion 121 444 122 445  0 t = 1
rlabel pdiffusion 124 444 125 445  0 t = 2
rlabel pdiffusion 121 449 122 450  0 t = 3
rlabel pdiffusion 124 449 125 450  0 t = 4
rlabel pdiffusion 120 444 126 450 0 cell no = 531
<< m1 >>
rect 121 444 122 445 
rect 124 444 125 445 
rect 121 449 122 450 
rect 124 449 125 450 
<< m2 >>
rect 121 444 122 445 
rect 124 444 125 445 
rect 121 449 122 450 
rect 124 449 125 450 
<< m2c >>
rect 121 444 122 445 
rect 124 444 125 445 
rect 121 449 122 450 
rect 124 449 125 450 
<< labels >>
rlabel pdiffusion 247 426 248 427  0 t = 1
rlabel pdiffusion 250 426 251 427  0 t = 2
rlabel pdiffusion 247 431 248 432  0 t = 3
rlabel pdiffusion 250 431 251 432  0 t = 4
rlabel pdiffusion 246 426 252 432 0 cell no = 532
<< m1 >>
rect 247 426 248 427 
rect 250 426 251 427 
rect 247 431 248 432 
rect 250 431 251 432 
<< m2 >>
rect 247 426 248 427 
rect 250 426 251 427 
rect 247 431 248 432 
rect 250 431 251 432 
<< m2c >>
rect 247 426 248 427 
rect 250 426 251 427 
rect 247 431 248 432 
rect 250 431 251 432 
<< labels >>
rlabel pdiffusion 211 444 212 445  0 t = 1
rlabel pdiffusion 214 444 215 445  0 t = 2
rlabel pdiffusion 211 449 212 450  0 t = 3
rlabel pdiffusion 214 449 215 450  0 t = 4
rlabel pdiffusion 210 444 216 450 0 cell no = 533
<< m1 >>
rect 211 444 212 445 
rect 214 444 215 445 
rect 211 449 212 450 
rect 214 449 215 450 
<< m2 >>
rect 211 444 212 445 
rect 214 444 215 445 
rect 211 449 212 450 
rect 214 449 215 450 
<< m2c >>
rect 211 444 212 445 
rect 214 444 215 445 
rect 211 449 212 450 
rect 214 449 215 450 
<< labels >>
rlabel pdiffusion 229 444 230 445  0 t = 1
rlabel pdiffusion 232 444 233 445  0 t = 2
rlabel pdiffusion 229 449 230 450  0 t = 3
rlabel pdiffusion 232 449 233 450  0 t = 4
rlabel pdiffusion 228 444 234 450 0 cell no = 534
<< m1 >>
rect 229 444 230 445 
rect 232 444 233 445 
rect 229 449 230 450 
rect 232 449 233 450 
<< m2 >>
rect 229 444 230 445 
rect 232 444 233 445 
rect 229 449 230 450 
rect 232 449 233 450 
<< m2c >>
rect 229 444 230 445 
rect 232 444 233 445 
rect 229 449 230 450 
rect 232 449 233 450 
<< labels >>
rlabel pdiffusion 157 444 158 445  0 t = 1
rlabel pdiffusion 160 444 161 445  0 t = 2
rlabel pdiffusion 157 449 158 450  0 t = 3
rlabel pdiffusion 160 449 161 450  0 t = 4
rlabel pdiffusion 156 444 162 450 0 cell no = 535
<< m1 >>
rect 157 444 158 445 
rect 160 444 161 445 
rect 157 449 158 450 
rect 160 449 161 450 
<< m2 >>
rect 157 444 158 445 
rect 160 444 161 445 
rect 157 449 158 450 
rect 160 449 161 450 
<< m2c >>
rect 157 444 158 445 
rect 160 444 161 445 
rect 157 449 158 450 
rect 160 449 161 450 
<< labels >>
rlabel pdiffusion 103 408 104 409  0 t = 1
rlabel pdiffusion 106 408 107 409  0 t = 2
rlabel pdiffusion 103 413 104 414  0 t = 3
rlabel pdiffusion 106 413 107 414  0 t = 4
rlabel pdiffusion 102 408 108 414 0 cell no = 536
<< m1 >>
rect 103 408 104 409 
rect 106 408 107 409 
rect 103 413 104 414 
rect 106 413 107 414 
<< m2 >>
rect 103 408 104 409 
rect 106 408 107 409 
rect 103 413 104 414 
rect 106 413 107 414 
<< m2c >>
rect 103 408 104 409 
rect 106 408 107 409 
rect 103 413 104 414 
rect 106 413 107 414 
<< labels >>
rlabel pdiffusion 229 66 230 67  0 t = 1
rlabel pdiffusion 232 66 233 67  0 t = 2
rlabel pdiffusion 229 71 230 72  0 t = 3
rlabel pdiffusion 232 71 233 72  0 t = 4
rlabel pdiffusion 228 66 234 72 0 cell no = 537
<< m1 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2c >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< labels >>
rlabel pdiffusion 247 336 248 337  0 t = 1
rlabel pdiffusion 250 336 251 337  0 t = 2
rlabel pdiffusion 247 341 248 342  0 t = 3
rlabel pdiffusion 250 341 251 342  0 t = 4
rlabel pdiffusion 246 336 252 342 0 cell no = 538
<< m1 >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< m2 >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< m2c >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< labels >>
rlabel pdiffusion 391 336 392 337  0 t = 1
rlabel pdiffusion 394 336 395 337  0 t = 2
rlabel pdiffusion 391 341 392 342  0 t = 3
rlabel pdiffusion 394 341 395 342  0 t = 4
rlabel pdiffusion 390 336 396 342 0 cell no = 539
<< m1 >>
rect 391 336 392 337 
rect 394 336 395 337 
rect 391 341 392 342 
rect 394 341 395 342 
<< m2 >>
rect 391 336 392 337 
rect 394 336 395 337 
rect 391 341 392 342 
rect 394 341 395 342 
<< m2c >>
rect 391 336 392 337 
rect 394 336 395 337 
rect 391 341 392 342 
rect 394 341 395 342 
<< labels >>
rlabel pdiffusion 301 300 302 301  0 t = 1
rlabel pdiffusion 304 300 305 301  0 t = 2
rlabel pdiffusion 301 305 302 306  0 t = 3
rlabel pdiffusion 304 305 305 306  0 t = 4
rlabel pdiffusion 300 300 306 306 0 cell no = 540
<< m1 >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< m2 >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< m2c >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< labels >>
rlabel pdiffusion 247 300 248 301  0 t = 1
rlabel pdiffusion 250 300 251 301  0 t = 2
rlabel pdiffusion 247 305 248 306  0 t = 3
rlabel pdiffusion 250 305 251 306  0 t = 4
rlabel pdiffusion 246 300 252 306 0 cell no = 541
<< m1 >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< m2 >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< m2c >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< labels >>
rlabel pdiffusion 445 300 446 301  0 t = 1
rlabel pdiffusion 448 300 449 301  0 t = 2
rlabel pdiffusion 445 305 446 306  0 t = 3
rlabel pdiffusion 448 305 449 306  0 t = 4
rlabel pdiffusion 444 300 450 306 0 cell no = 542
<< m1 >>
rect 445 300 446 301 
rect 448 300 449 301 
rect 445 305 446 306 
rect 448 305 449 306 
<< m2 >>
rect 445 300 446 301 
rect 448 300 449 301 
rect 445 305 446 306 
rect 448 305 449 306 
<< m2c >>
rect 445 300 446 301 
rect 448 300 449 301 
rect 445 305 446 306 
rect 448 305 449 306 
<< labels >>
rlabel pdiffusion 373 372 374 373  0 t = 1
rlabel pdiffusion 376 372 377 373  0 t = 2
rlabel pdiffusion 373 377 374 378  0 t = 3
rlabel pdiffusion 376 377 377 378  0 t = 4
rlabel pdiffusion 372 372 378 378 0 cell no = 543
<< m1 >>
rect 373 372 374 373 
rect 376 372 377 373 
rect 373 377 374 378 
rect 376 377 377 378 
<< m2 >>
rect 373 372 374 373 
rect 376 372 377 373 
rect 373 377 374 378 
rect 376 377 377 378 
<< m2c >>
rect 373 372 374 373 
rect 376 372 377 373 
rect 373 377 374 378 
rect 376 377 377 378 
<< labels >>
rlabel pdiffusion 265 318 266 319  0 t = 1
rlabel pdiffusion 268 318 269 319  0 t = 2
rlabel pdiffusion 265 323 266 324  0 t = 3
rlabel pdiffusion 268 323 269 324  0 t = 4
rlabel pdiffusion 264 318 270 324 0 cell no = 544
<< m1 >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< m2 >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< m2c >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< labels >>
rlabel pdiffusion 355 318 356 319  0 t = 1
rlabel pdiffusion 358 318 359 319  0 t = 2
rlabel pdiffusion 355 323 356 324  0 t = 3
rlabel pdiffusion 358 323 359 324  0 t = 4
rlabel pdiffusion 354 318 360 324 0 cell no = 545
<< m1 >>
rect 355 318 356 319 
rect 358 318 359 319 
rect 355 323 356 324 
rect 358 323 359 324 
<< m2 >>
rect 355 318 356 319 
rect 358 318 359 319 
rect 355 323 356 324 
rect 358 323 359 324 
<< m2c >>
rect 355 318 356 319 
rect 358 318 359 319 
rect 355 323 356 324 
rect 358 323 359 324 
<< labels >>
rlabel pdiffusion 391 372 392 373  0 t = 1
rlabel pdiffusion 394 372 395 373  0 t = 2
rlabel pdiffusion 391 377 392 378  0 t = 3
rlabel pdiffusion 394 377 395 378  0 t = 4
rlabel pdiffusion 390 372 396 378 0 cell no = 546
<< m1 >>
rect 391 372 392 373 
rect 394 372 395 373 
rect 391 377 392 378 
rect 394 377 395 378 
<< m2 >>
rect 391 372 392 373 
rect 394 372 395 373 
rect 391 377 392 378 
rect 394 377 395 378 
<< m2c >>
rect 391 372 392 373 
rect 394 372 395 373 
rect 391 377 392 378 
rect 394 377 395 378 
<< labels >>
rlabel pdiffusion 337 318 338 319  0 t = 1
rlabel pdiffusion 340 318 341 319  0 t = 2
rlabel pdiffusion 337 323 338 324  0 t = 3
rlabel pdiffusion 340 323 341 324  0 t = 4
rlabel pdiffusion 336 318 342 324 0 cell no = 547
<< m1 >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< m2 >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< m2c >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< labels >>
rlabel pdiffusion 391 408 392 409  0 t = 1
rlabel pdiffusion 394 408 395 409  0 t = 2
rlabel pdiffusion 391 413 392 414  0 t = 3
rlabel pdiffusion 394 413 395 414  0 t = 4
rlabel pdiffusion 390 408 396 414 0 cell no = 548
<< m1 >>
rect 391 408 392 409 
rect 394 408 395 409 
rect 391 413 392 414 
rect 394 413 395 414 
<< m2 >>
rect 391 408 392 409 
rect 394 408 395 409 
rect 391 413 392 414 
rect 394 413 395 414 
<< m2c >>
rect 391 408 392 409 
rect 394 408 395 409 
rect 391 413 392 414 
rect 394 413 395 414 
<< labels >>
rlabel pdiffusion 355 372 356 373  0 t = 1
rlabel pdiffusion 358 372 359 373  0 t = 2
rlabel pdiffusion 355 377 356 378  0 t = 3
rlabel pdiffusion 358 377 359 378  0 t = 4
rlabel pdiffusion 354 372 360 378 0 cell no = 549
<< m1 >>
rect 355 372 356 373 
rect 358 372 359 373 
rect 355 377 356 378 
rect 358 377 359 378 
<< m2 >>
rect 355 372 356 373 
rect 358 372 359 373 
rect 355 377 356 378 
rect 358 377 359 378 
<< m2c >>
rect 355 372 356 373 
rect 358 372 359 373 
rect 355 377 356 378 
rect 358 377 359 378 
<< labels >>
rlabel pdiffusion 301 372 302 373  0 t = 1
rlabel pdiffusion 304 372 305 373  0 t = 2
rlabel pdiffusion 301 377 302 378  0 t = 3
rlabel pdiffusion 304 377 305 378  0 t = 4
rlabel pdiffusion 300 372 306 378 0 cell no = 550
<< m1 >>
rect 301 372 302 373 
rect 304 372 305 373 
rect 301 377 302 378 
rect 304 377 305 378 
<< m2 >>
rect 301 372 302 373 
rect 304 372 305 373 
rect 301 377 302 378 
rect 304 377 305 378 
<< m2c >>
rect 301 372 302 373 
rect 304 372 305 373 
rect 301 377 302 378 
rect 304 377 305 378 
<< labels >>
rlabel pdiffusion 31 354 32 355  0 t = 1
rlabel pdiffusion 34 354 35 355  0 t = 2
rlabel pdiffusion 31 359 32 360  0 t = 3
rlabel pdiffusion 34 359 35 360  0 t = 4
rlabel pdiffusion 30 354 36 360 0 cell no = 551
<< m1 >>
rect 31 354 32 355 
rect 34 354 35 355 
rect 31 359 32 360 
rect 34 359 35 360 
<< m2 >>
rect 31 354 32 355 
rect 34 354 35 355 
rect 31 359 32 360 
rect 34 359 35 360 
<< m2c >>
rect 31 354 32 355 
rect 34 354 35 355 
rect 31 359 32 360 
rect 34 359 35 360 
<< labels >>
rlabel pdiffusion 13 408 14 409  0 t = 1
rlabel pdiffusion 16 408 17 409  0 t = 2
rlabel pdiffusion 13 413 14 414  0 t = 3
rlabel pdiffusion 16 413 17 414  0 t = 4
rlabel pdiffusion 12 408 18 414 0 cell no = 552
<< m1 >>
rect 13 408 14 409 
rect 16 408 17 409 
rect 13 413 14 414 
rect 16 413 17 414 
<< m2 >>
rect 13 408 14 409 
rect 16 408 17 409 
rect 13 413 14 414 
rect 16 413 17 414 
<< m2c >>
rect 13 408 14 409 
rect 16 408 17 409 
rect 13 413 14 414 
rect 16 413 17 414 
<< labels >>
rlabel pdiffusion 337 354 338 355  0 t = 1
rlabel pdiffusion 340 354 341 355  0 t = 2
rlabel pdiffusion 337 359 338 360  0 t = 3
rlabel pdiffusion 340 359 341 360  0 t = 4
rlabel pdiffusion 336 354 342 360 0 cell no = 553
<< m1 >>
rect 337 354 338 355 
rect 340 354 341 355 
rect 337 359 338 360 
rect 340 359 341 360 
<< m2 >>
rect 337 354 338 355 
rect 340 354 341 355 
rect 337 359 338 360 
rect 340 359 341 360 
<< m2c >>
rect 337 354 338 355 
rect 340 354 341 355 
rect 337 359 338 360 
rect 340 359 341 360 
<< labels >>
rlabel pdiffusion 373 138 374 139  0 t = 1
rlabel pdiffusion 376 138 377 139  0 t = 2
rlabel pdiffusion 373 143 374 144  0 t = 3
rlabel pdiffusion 376 143 377 144  0 t = 4
rlabel pdiffusion 372 138 378 144 0 cell no = 554
<< m1 >>
rect 373 138 374 139 
rect 376 138 377 139 
rect 373 143 374 144 
rect 376 143 377 144 
<< m2 >>
rect 373 138 374 139 
rect 376 138 377 139 
rect 373 143 374 144 
rect 376 143 377 144 
<< m2c >>
rect 373 138 374 139 
rect 376 138 377 139 
rect 373 143 374 144 
rect 376 143 377 144 
<< labels >>
rlabel pdiffusion 265 264 266 265  0 t = 1
rlabel pdiffusion 268 264 269 265  0 t = 2
rlabel pdiffusion 265 269 266 270  0 t = 3
rlabel pdiffusion 268 269 269 270  0 t = 4
rlabel pdiffusion 264 264 270 270 0 cell no = 555
<< m1 >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< m2 >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< m2c >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< labels >>
rlabel pdiffusion 157 426 158 427  0 t = 1
rlabel pdiffusion 160 426 161 427  0 t = 2
rlabel pdiffusion 157 431 158 432  0 t = 3
rlabel pdiffusion 160 431 161 432  0 t = 4
rlabel pdiffusion 156 426 162 432 0 cell no = 556
<< m1 >>
rect 157 426 158 427 
rect 160 426 161 427 
rect 157 431 158 432 
rect 160 431 161 432 
<< m2 >>
rect 157 426 158 427 
rect 160 426 161 427 
rect 157 431 158 432 
rect 160 431 161 432 
<< m2c >>
rect 157 426 158 427 
rect 160 426 161 427 
rect 157 431 158 432 
rect 160 431 161 432 
<< labels >>
rlabel pdiffusion 445 30 446 31  0 t = 1
rlabel pdiffusion 448 30 449 31  0 t = 2
rlabel pdiffusion 445 35 446 36  0 t = 3
rlabel pdiffusion 448 35 449 36  0 t = 4
rlabel pdiffusion 444 30 450 36 0 cell no = 557
<< m1 >>
rect 445 30 446 31 
rect 448 30 449 31 
rect 445 35 446 36 
rect 448 35 449 36 
<< m2 >>
rect 445 30 446 31 
rect 448 30 449 31 
rect 445 35 446 36 
rect 448 35 449 36 
<< m2c >>
rect 445 30 446 31 
rect 448 30 449 31 
rect 445 35 446 36 
rect 448 35 449 36 
<< labels >>
rlabel pdiffusion 175 408 176 409  0 t = 1
rlabel pdiffusion 178 408 179 409  0 t = 2
rlabel pdiffusion 175 413 176 414  0 t = 3
rlabel pdiffusion 178 413 179 414  0 t = 4
rlabel pdiffusion 174 408 180 414 0 cell no = 558
<< m1 >>
rect 175 408 176 409 
rect 178 408 179 409 
rect 175 413 176 414 
rect 178 413 179 414 
<< m2 >>
rect 175 408 176 409 
rect 178 408 179 409 
rect 175 413 176 414 
rect 178 413 179 414 
<< m2c >>
rect 175 408 176 409 
rect 178 408 179 409 
rect 175 413 176 414 
rect 178 413 179 414 
<< labels >>
rlabel pdiffusion 319 390 320 391  0 t = 1
rlabel pdiffusion 322 390 323 391  0 t = 2
rlabel pdiffusion 319 395 320 396  0 t = 3
rlabel pdiffusion 322 395 323 396  0 t = 4
rlabel pdiffusion 318 390 324 396 0 cell no = 559
<< m1 >>
rect 319 390 320 391 
rect 322 390 323 391 
rect 319 395 320 396 
rect 322 395 323 396 
<< m2 >>
rect 319 390 320 391 
rect 322 390 323 391 
rect 319 395 320 396 
rect 322 395 323 396 
<< m2c >>
rect 319 390 320 391 
rect 322 390 323 391 
rect 319 395 320 396 
rect 322 395 323 396 
<< labels >>
rlabel pdiffusion 229 156 230 157  0 t = 1
rlabel pdiffusion 232 156 233 157  0 t = 2
rlabel pdiffusion 229 161 230 162  0 t = 3
rlabel pdiffusion 232 161 233 162  0 t = 4
rlabel pdiffusion 228 156 234 162 0 cell no = 560
<< m1 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2c >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< labels >>
rlabel pdiffusion 265 444 266 445  0 t = 1
rlabel pdiffusion 268 444 269 445  0 t = 2
rlabel pdiffusion 265 449 266 450  0 t = 3
rlabel pdiffusion 268 449 269 450  0 t = 4
rlabel pdiffusion 264 444 270 450 0 cell no = 561
<< m1 >>
rect 265 444 266 445 
rect 268 444 269 445 
rect 265 449 266 450 
rect 268 449 269 450 
<< m2 >>
rect 265 444 266 445 
rect 268 444 269 445 
rect 265 449 266 450 
rect 268 449 269 450 
<< m2c >>
rect 265 444 266 445 
rect 268 444 269 445 
rect 265 449 266 450 
rect 268 449 269 450 
<< labels >>
rlabel pdiffusion 229 336 230 337  0 t = 1
rlabel pdiffusion 232 336 233 337  0 t = 2
rlabel pdiffusion 229 341 230 342  0 t = 3
rlabel pdiffusion 232 341 233 342  0 t = 4
rlabel pdiffusion 228 336 234 342 0 cell no = 562
<< m1 >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< m2 >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< m2c >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< labels >>
rlabel pdiffusion 445 120 446 121  0 t = 1
rlabel pdiffusion 448 120 449 121  0 t = 2
rlabel pdiffusion 445 125 446 126  0 t = 3
rlabel pdiffusion 448 125 449 126  0 t = 4
rlabel pdiffusion 444 120 450 126 0 cell no = 563
<< m1 >>
rect 445 120 446 121 
rect 448 120 449 121 
rect 445 125 446 126 
rect 448 125 449 126 
<< m2 >>
rect 445 120 446 121 
rect 448 120 449 121 
rect 445 125 446 126 
rect 448 125 449 126 
<< m2c >>
rect 445 120 446 121 
rect 448 120 449 121 
rect 445 125 446 126 
rect 448 125 449 126 
<< labels >>
rlabel pdiffusion 301 192 302 193  0 t = 1
rlabel pdiffusion 304 192 305 193  0 t = 2
rlabel pdiffusion 301 197 302 198  0 t = 3
rlabel pdiffusion 304 197 305 198  0 t = 4
rlabel pdiffusion 300 192 306 198 0 cell no = 564
<< m1 >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< m2 >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< m2c >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< labels >>
rlabel pdiffusion 283 390 284 391  0 t = 1
rlabel pdiffusion 286 390 287 391  0 t = 2
rlabel pdiffusion 283 395 284 396  0 t = 3
rlabel pdiffusion 286 395 287 396  0 t = 4
rlabel pdiffusion 282 390 288 396 0 cell no = 565
<< m1 >>
rect 283 390 284 391 
rect 286 390 287 391 
rect 283 395 284 396 
rect 286 395 287 396 
<< m2 >>
rect 283 390 284 391 
rect 286 390 287 391 
rect 283 395 284 396 
rect 286 395 287 396 
<< m2c >>
rect 283 390 284 391 
rect 286 390 287 391 
rect 283 395 284 396 
rect 286 395 287 396 
<< labels >>
rlabel pdiffusion 85 408 86 409  0 t = 1
rlabel pdiffusion 88 408 89 409  0 t = 2
rlabel pdiffusion 85 413 86 414  0 t = 3
rlabel pdiffusion 88 413 89 414  0 t = 4
rlabel pdiffusion 84 408 90 414 0 cell no = 566
<< m1 >>
rect 85 408 86 409 
rect 88 408 89 409 
rect 85 413 86 414 
rect 88 413 89 414 
<< m2 >>
rect 85 408 86 409 
rect 88 408 89 409 
rect 85 413 86 414 
rect 88 413 89 414 
<< m2c >>
rect 85 408 86 409 
rect 88 408 89 409 
rect 85 413 86 414 
rect 88 413 89 414 
<< labels >>
rlabel pdiffusion 355 426 356 427  0 t = 1
rlabel pdiffusion 358 426 359 427  0 t = 2
rlabel pdiffusion 355 431 356 432  0 t = 3
rlabel pdiffusion 358 431 359 432  0 t = 4
rlabel pdiffusion 354 426 360 432 0 cell no = 567
<< m1 >>
rect 355 426 356 427 
rect 358 426 359 427 
rect 355 431 356 432 
rect 358 431 359 432 
<< m2 >>
rect 355 426 356 427 
rect 358 426 359 427 
rect 355 431 356 432 
rect 358 431 359 432 
<< m2c >>
rect 355 426 356 427 
rect 358 426 359 427 
rect 355 431 356 432 
rect 358 431 359 432 
<< labels >>
rlabel pdiffusion 427 390 428 391  0 t = 1
rlabel pdiffusion 430 390 431 391  0 t = 2
rlabel pdiffusion 427 395 428 396  0 t = 3
rlabel pdiffusion 430 395 431 396  0 t = 4
rlabel pdiffusion 426 390 432 396 0 cell no = 568
<< m1 >>
rect 427 390 428 391 
rect 430 390 431 391 
rect 427 395 428 396 
rect 430 395 431 396 
<< m2 >>
rect 427 390 428 391 
rect 430 390 431 391 
rect 427 395 428 396 
rect 430 395 431 396 
<< m2c >>
rect 427 390 428 391 
rect 430 390 431 391 
rect 427 395 428 396 
rect 430 395 431 396 
<< labels >>
rlabel pdiffusion 409 336 410 337  0 t = 1
rlabel pdiffusion 412 336 413 337  0 t = 2
rlabel pdiffusion 409 341 410 342  0 t = 3
rlabel pdiffusion 412 341 413 342  0 t = 4
rlabel pdiffusion 408 336 414 342 0 cell no = 569
<< m1 >>
rect 409 336 410 337 
rect 412 336 413 337 
rect 409 341 410 342 
rect 412 341 413 342 
<< m2 >>
rect 409 336 410 337 
rect 412 336 413 337 
rect 409 341 410 342 
rect 412 341 413 342 
<< m2c >>
rect 409 336 410 337 
rect 412 336 413 337 
rect 409 341 410 342 
rect 412 341 413 342 
<< labels >>
rlabel pdiffusion 409 318 410 319  0 t = 1
rlabel pdiffusion 412 318 413 319  0 t = 2
rlabel pdiffusion 409 323 410 324  0 t = 3
rlabel pdiffusion 412 323 413 324  0 t = 4
rlabel pdiffusion 408 318 414 324 0 cell no = 570
<< m1 >>
rect 409 318 410 319 
rect 412 318 413 319 
rect 409 323 410 324 
rect 412 323 413 324 
<< m2 >>
rect 409 318 410 319 
rect 412 318 413 319 
rect 409 323 410 324 
rect 412 323 413 324 
<< m2c >>
rect 409 318 410 319 
rect 412 318 413 319 
rect 409 323 410 324 
rect 412 323 413 324 
<< labels >>
rlabel pdiffusion 391 318 392 319  0 t = 1
rlabel pdiffusion 394 318 395 319  0 t = 2
rlabel pdiffusion 391 323 392 324  0 t = 3
rlabel pdiffusion 394 323 395 324  0 t = 4
rlabel pdiffusion 390 318 396 324 0 cell no = 571
<< m1 >>
rect 391 318 392 319 
rect 394 318 395 319 
rect 391 323 392 324 
rect 394 323 395 324 
<< m2 >>
rect 391 318 392 319 
rect 394 318 395 319 
rect 391 323 392 324 
rect 394 323 395 324 
<< m2c >>
rect 391 318 392 319 
rect 394 318 395 319 
rect 391 323 392 324 
rect 394 323 395 324 
<< labels >>
rlabel pdiffusion 445 336 446 337  0 t = 1
rlabel pdiffusion 448 336 449 337  0 t = 2
rlabel pdiffusion 445 341 446 342  0 t = 3
rlabel pdiffusion 448 341 449 342  0 t = 4
rlabel pdiffusion 444 336 450 342 0 cell no = 572
<< m1 >>
rect 445 336 446 337 
rect 448 336 449 337 
rect 445 341 446 342 
rect 448 341 449 342 
<< m2 >>
rect 445 336 446 337 
rect 448 336 449 337 
rect 445 341 446 342 
rect 448 341 449 342 
<< m2c >>
rect 445 336 446 337 
rect 448 336 449 337 
rect 445 341 446 342 
rect 448 341 449 342 
<< labels >>
rlabel pdiffusion 265 354 266 355  0 t = 1
rlabel pdiffusion 268 354 269 355  0 t = 2
rlabel pdiffusion 265 359 266 360  0 t = 3
rlabel pdiffusion 268 359 269 360  0 t = 4
rlabel pdiffusion 264 354 270 360 0 cell no = 573
<< m1 >>
rect 265 354 266 355 
rect 268 354 269 355 
rect 265 359 266 360 
rect 268 359 269 360 
<< m2 >>
rect 265 354 266 355 
rect 268 354 269 355 
rect 265 359 266 360 
rect 268 359 269 360 
<< m2c >>
rect 265 354 266 355 
rect 268 354 269 355 
rect 265 359 266 360 
rect 268 359 269 360 
<< labels >>
rlabel pdiffusion 445 426 446 427  0 t = 1
rlabel pdiffusion 448 426 449 427  0 t = 2
rlabel pdiffusion 445 431 446 432  0 t = 3
rlabel pdiffusion 448 431 449 432  0 t = 4
rlabel pdiffusion 444 426 450 432 0 cell no = 574
<< m1 >>
rect 445 426 446 427 
rect 448 426 449 427 
rect 445 431 446 432 
rect 448 431 449 432 
<< m2 >>
rect 445 426 446 427 
rect 448 426 449 427 
rect 445 431 446 432 
rect 448 431 449 432 
<< m2c >>
rect 445 426 446 427 
rect 448 426 449 427 
rect 445 431 446 432 
rect 448 431 449 432 
<< labels >>
rlabel pdiffusion 373 408 374 409  0 t = 1
rlabel pdiffusion 376 408 377 409  0 t = 2
rlabel pdiffusion 373 413 374 414  0 t = 3
rlabel pdiffusion 376 413 377 414  0 t = 4
rlabel pdiffusion 372 408 378 414 0 cell no = 575
<< m1 >>
rect 373 408 374 409 
rect 376 408 377 409 
rect 373 413 374 414 
rect 376 413 377 414 
<< m2 >>
rect 373 408 374 409 
rect 376 408 377 409 
rect 373 413 374 414 
rect 376 413 377 414 
<< m2c >>
rect 373 408 374 409 
rect 376 408 377 409 
rect 373 413 374 414 
rect 376 413 377 414 
<< labels >>
rlabel pdiffusion 85 336 86 337  0 t = 1
rlabel pdiffusion 88 336 89 337  0 t = 2
rlabel pdiffusion 85 341 86 342  0 t = 3
rlabel pdiffusion 88 341 89 342  0 t = 4
rlabel pdiffusion 84 336 90 342 0 cell no = 576
<< m1 >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< m2 >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< m2c >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< labels >>
rlabel pdiffusion 175 372 176 373  0 t = 1
rlabel pdiffusion 178 372 179 373  0 t = 2
rlabel pdiffusion 175 377 176 378  0 t = 3
rlabel pdiffusion 178 377 179 378  0 t = 4
rlabel pdiffusion 174 372 180 378 0 cell no = 577
<< m1 >>
rect 175 372 176 373 
rect 178 372 179 373 
rect 175 377 176 378 
rect 178 377 179 378 
<< m2 >>
rect 175 372 176 373 
rect 178 372 179 373 
rect 175 377 176 378 
rect 178 377 179 378 
<< m2c >>
rect 175 372 176 373 
rect 178 372 179 373 
rect 175 377 176 378 
rect 178 377 179 378 
<< labels >>
rlabel pdiffusion 85 444 86 445  0 t = 1
rlabel pdiffusion 88 444 89 445  0 t = 2
rlabel pdiffusion 85 449 86 450  0 t = 3
rlabel pdiffusion 88 449 89 450  0 t = 4
rlabel pdiffusion 84 444 90 450 0 cell no = 578
<< m1 >>
rect 85 444 86 445 
rect 88 444 89 445 
rect 85 449 86 450 
rect 88 449 89 450 
<< m2 >>
rect 85 444 86 445 
rect 88 444 89 445 
rect 85 449 86 450 
rect 88 449 89 450 
<< m2c >>
rect 85 444 86 445 
rect 88 444 89 445 
rect 85 449 86 450 
rect 88 449 89 450 
<< labels >>
rlabel pdiffusion 265 138 266 139  0 t = 1
rlabel pdiffusion 268 138 269 139  0 t = 2
rlabel pdiffusion 265 143 266 144  0 t = 3
rlabel pdiffusion 268 143 269 144  0 t = 4
rlabel pdiffusion 264 138 270 144 0 cell no = 579
<< m1 >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< m2 >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< m2c >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< labels >>
rlabel pdiffusion 265 408 266 409  0 t = 1
rlabel pdiffusion 268 408 269 409  0 t = 2
rlabel pdiffusion 265 413 266 414  0 t = 3
rlabel pdiffusion 268 413 269 414  0 t = 4
rlabel pdiffusion 264 408 270 414 0 cell no = 580
<< m1 >>
rect 265 408 266 409 
rect 268 408 269 409 
rect 265 413 266 414 
rect 268 413 269 414 
<< m2 >>
rect 265 408 266 409 
rect 268 408 269 409 
rect 265 413 266 414 
rect 268 413 269 414 
<< m2c >>
rect 265 408 266 409 
rect 268 408 269 409 
rect 265 413 266 414 
rect 268 413 269 414 
<< labels >>
rlabel pdiffusion 283 408 284 409  0 t = 1
rlabel pdiffusion 286 408 287 409  0 t = 2
rlabel pdiffusion 283 413 284 414  0 t = 3
rlabel pdiffusion 286 413 287 414  0 t = 4
rlabel pdiffusion 282 408 288 414 0 cell no = 581
<< m1 >>
rect 283 408 284 409 
rect 286 408 287 409 
rect 283 413 284 414 
rect 286 413 287 414 
<< m2 >>
rect 283 408 284 409 
rect 286 408 287 409 
rect 283 413 284 414 
rect 286 413 287 414 
<< m2c >>
rect 283 408 284 409 
rect 286 408 287 409 
rect 283 413 284 414 
rect 286 413 287 414 
<< labels >>
rlabel pdiffusion 31 444 32 445  0 t = 1
rlabel pdiffusion 34 444 35 445  0 t = 2
rlabel pdiffusion 31 449 32 450  0 t = 3
rlabel pdiffusion 34 449 35 450  0 t = 4
rlabel pdiffusion 30 444 36 450 0 cell no = 582
<< m1 >>
rect 31 444 32 445 
rect 34 444 35 445 
rect 31 449 32 450 
rect 34 449 35 450 
<< m2 >>
rect 31 444 32 445 
rect 34 444 35 445 
rect 31 449 32 450 
rect 34 449 35 450 
<< m2c >>
rect 31 444 32 445 
rect 34 444 35 445 
rect 31 449 32 450 
rect 34 449 35 450 
<< labels >>
rlabel pdiffusion 31 282 32 283  0 t = 1
rlabel pdiffusion 34 282 35 283  0 t = 2
rlabel pdiffusion 31 287 32 288  0 t = 3
rlabel pdiffusion 34 287 35 288  0 t = 4
rlabel pdiffusion 30 282 36 288 0 cell no = 583
<< m1 >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< m2 >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< m2c >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< labels >>
rlabel pdiffusion 301 408 302 409  0 t = 1
rlabel pdiffusion 304 408 305 409  0 t = 2
rlabel pdiffusion 301 413 302 414  0 t = 3
rlabel pdiffusion 304 413 305 414  0 t = 4
rlabel pdiffusion 300 408 306 414 0 cell no = 584
<< m1 >>
rect 301 408 302 409 
rect 304 408 305 409 
rect 301 413 302 414 
rect 304 413 305 414 
<< m2 >>
rect 301 408 302 409 
rect 304 408 305 409 
rect 301 413 302 414 
rect 304 413 305 414 
<< m2c >>
rect 301 408 302 409 
rect 304 408 305 409 
rect 301 413 302 414 
rect 304 413 305 414 
<< labels >>
rlabel pdiffusion 337 408 338 409  0 t = 1
rlabel pdiffusion 340 408 341 409  0 t = 2
rlabel pdiffusion 337 413 338 414  0 t = 3
rlabel pdiffusion 340 413 341 414  0 t = 4
rlabel pdiffusion 336 408 342 414 0 cell no = 585
<< m1 >>
rect 337 408 338 409 
rect 340 408 341 409 
rect 337 413 338 414 
rect 340 413 341 414 
<< m2 >>
rect 337 408 338 409 
rect 340 408 341 409 
rect 337 413 338 414 
rect 340 413 341 414 
<< m2c >>
rect 337 408 338 409 
rect 340 408 341 409 
rect 337 413 338 414 
rect 340 413 341 414 
<< labels >>
rlabel pdiffusion 211 408 212 409  0 t = 1
rlabel pdiffusion 214 408 215 409  0 t = 2
rlabel pdiffusion 211 413 212 414  0 t = 3
rlabel pdiffusion 214 413 215 414  0 t = 4
rlabel pdiffusion 210 408 216 414 0 cell no = 586
<< m1 >>
rect 211 408 212 409 
rect 214 408 215 409 
rect 211 413 212 414 
rect 214 413 215 414 
<< m2 >>
rect 211 408 212 409 
rect 214 408 215 409 
rect 211 413 212 414 
rect 214 413 215 414 
<< m2c >>
rect 211 408 212 409 
rect 214 408 215 409 
rect 211 413 212 414 
rect 214 413 215 414 
<< labels >>
rlabel pdiffusion 229 408 230 409  0 t = 1
rlabel pdiffusion 232 408 233 409  0 t = 2
rlabel pdiffusion 229 413 230 414  0 t = 3
rlabel pdiffusion 232 413 233 414  0 t = 4
rlabel pdiffusion 228 408 234 414 0 cell no = 587
<< m1 >>
rect 229 408 230 409 
rect 232 408 233 409 
rect 229 413 230 414 
rect 232 413 233 414 
<< m2 >>
rect 229 408 230 409 
rect 232 408 233 409 
rect 229 413 230 414 
rect 232 413 233 414 
<< m2c >>
rect 229 408 230 409 
rect 232 408 233 409 
rect 229 413 230 414 
rect 232 413 233 414 
<< labels >>
rlabel pdiffusion 211 390 212 391  0 t = 1
rlabel pdiffusion 214 390 215 391  0 t = 2
rlabel pdiffusion 211 395 212 396  0 t = 3
rlabel pdiffusion 214 395 215 396  0 t = 4
rlabel pdiffusion 210 390 216 396 0 cell no = 588
<< m1 >>
rect 211 390 212 391 
rect 214 390 215 391 
rect 211 395 212 396 
rect 214 395 215 396 
<< m2 >>
rect 211 390 212 391 
rect 214 390 215 391 
rect 211 395 212 396 
rect 214 395 215 396 
<< m2c >>
rect 211 390 212 391 
rect 214 390 215 391 
rect 211 395 212 396 
rect 214 395 215 396 
<< labels >>
rlabel pdiffusion 247 444 248 445  0 t = 1
rlabel pdiffusion 250 444 251 445  0 t = 2
rlabel pdiffusion 247 449 248 450  0 t = 3
rlabel pdiffusion 250 449 251 450  0 t = 4
rlabel pdiffusion 246 444 252 450 0 cell no = 589
<< m1 >>
rect 247 444 248 445 
rect 250 444 251 445 
rect 247 449 248 450 
rect 250 449 251 450 
<< m2 >>
rect 247 444 248 445 
rect 250 444 251 445 
rect 247 449 248 450 
rect 250 449 251 450 
<< m2c >>
rect 247 444 248 445 
rect 250 444 251 445 
rect 247 449 248 450 
rect 250 449 251 450 
<< labels >>
rlabel pdiffusion 247 408 248 409  0 t = 1
rlabel pdiffusion 250 408 251 409  0 t = 2
rlabel pdiffusion 247 413 248 414  0 t = 3
rlabel pdiffusion 250 413 251 414  0 t = 4
rlabel pdiffusion 246 408 252 414 0 cell no = 590
<< m1 >>
rect 247 408 248 409 
rect 250 408 251 409 
rect 247 413 248 414 
rect 250 413 251 414 
<< m2 >>
rect 247 408 248 409 
rect 250 408 251 409 
rect 247 413 248 414 
rect 250 413 251 414 
<< m2c >>
rect 247 408 248 409 
rect 250 408 251 409 
rect 247 413 248 414 
rect 250 413 251 414 
<< labels >>
rlabel pdiffusion 283 444 284 445  0 t = 1
rlabel pdiffusion 286 444 287 445  0 t = 2
rlabel pdiffusion 283 449 284 450  0 t = 3
rlabel pdiffusion 286 449 287 450  0 t = 4
rlabel pdiffusion 282 444 288 450 0 cell no = 591
<< m1 >>
rect 283 444 284 445 
rect 286 444 287 445 
rect 283 449 284 450 
rect 286 449 287 450 
<< m2 >>
rect 283 444 284 445 
rect 286 444 287 445 
rect 283 449 284 450 
rect 286 449 287 450 
<< m2c >>
rect 283 444 284 445 
rect 286 444 287 445 
rect 283 449 284 450 
rect 286 449 287 450 
<< labels >>
rlabel pdiffusion 265 336 266 337  0 t = 1
rlabel pdiffusion 268 336 269 337  0 t = 2
rlabel pdiffusion 265 341 266 342  0 t = 3
rlabel pdiffusion 268 341 269 342  0 t = 4
rlabel pdiffusion 264 336 270 342 0 cell no = 592
<< m1 >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< m2 >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< m2c >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< labels >>
rlabel pdiffusion 193 282 194 283  0 t = 1
rlabel pdiffusion 196 282 197 283  0 t = 2
rlabel pdiffusion 193 287 194 288  0 t = 3
rlabel pdiffusion 196 287 197 288  0 t = 4
rlabel pdiffusion 192 282 198 288 0 cell no = 593
<< m1 >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< m2 >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< m2c >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< labels >>
rlabel pdiffusion 121 408 122 409  0 t = 1
rlabel pdiffusion 124 408 125 409  0 t = 2
rlabel pdiffusion 121 413 122 414  0 t = 3
rlabel pdiffusion 124 413 125 414  0 t = 4
rlabel pdiffusion 120 408 126 414 0 cell no = 594
<< m1 >>
rect 121 408 122 409 
rect 124 408 125 409 
rect 121 413 122 414 
rect 124 413 125 414 
<< m2 >>
rect 121 408 122 409 
rect 124 408 125 409 
rect 121 413 122 414 
rect 124 413 125 414 
<< m2c >>
rect 121 408 122 409 
rect 124 408 125 409 
rect 121 413 122 414 
rect 124 413 125 414 
<< labels >>
rlabel pdiffusion 247 192 248 193  0 t = 1
rlabel pdiffusion 250 192 251 193  0 t = 2
rlabel pdiffusion 247 197 248 198  0 t = 3
rlabel pdiffusion 250 197 251 198  0 t = 4
rlabel pdiffusion 246 192 252 198 0 cell no = 595
<< m1 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2c >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< labels >>
rlabel pdiffusion 427 444 428 445  0 t = 1
rlabel pdiffusion 430 444 431 445  0 t = 2
rlabel pdiffusion 427 449 428 450  0 t = 3
rlabel pdiffusion 430 449 431 450  0 t = 4
rlabel pdiffusion 426 444 432 450 0 cell no = 596
<< m1 >>
rect 427 444 428 445 
rect 430 444 431 445 
rect 427 449 428 450 
rect 430 449 431 450 
<< m2 >>
rect 427 444 428 445 
rect 430 444 431 445 
rect 427 449 428 450 
rect 430 449 431 450 
<< m2c >>
rect 427 444 428 445 
rect 430 444 431 445 
rect 427 449 428 450 
rect 430 449 431 450 
<< labels >>
rlabel pdiffusion 139 426 140 427  0 t = 1
rlabel pdiffusion 142 426 143 427  0 t = 2
rlabel pdiffusion 139 431 140 432  0 t = 3
rlabel pdiffusion 142 431 143 432  0 t = 4
rlabel pdiffusion 138 426 144 432 0 cell no = 597
<< m1 >>
rect 139 426 140 427 
rect 142 426 143 427 
rect 139 431 140 432 
rect 142 431 143 432 
<< m2 >>
rect 139 426 140 427 
rect 142 426 143 427 
rect 139 431 140 432 
rect 142 431 143 432 
<< m2c >>
rect 139 426 140 427 
rect 142 426 143 427 
rect 139 431 140 432 
rect 142 431 143 432 
<< labels >>
rlabel pdiffusion 319 426 320 427  0 t = 1
rlabel pdiffusion 322 426 323 427  0 t = 2
rlabel pdiffusion 319 431 320 432  0 t = 3
rlabel pdiffusion 322 431 323 432  0 t = 4
rlabel pdiffusion 318 426 324 432 0 cell no = 598
<< m1 >>
rect 319 426 320 427 
rect 322 426 323 427 
rect 319 431 320 432 
rect 322 431 323 432 
<< m2 >>
rect 319 426 320 427 
rect 322 426 323 427 
rect 319 431 320 432 
rect 322 431 323 432 
<< m2c >>
rect 319 426 320 427 
rect 322 426 323 427 
rect 319 431 320 432 
rect 322 431 323 432 
<< labels >>
rlabel pdiffusion 229 390 230 391  0 t = 1
rlabel pdiffusion 232 390 233 391  0 t = 2
rlabel pdiffusion 229 395 230 396  0 t = 3
rlabel pdiffusion 232 395 233 396  0 t = 4
rlabel pdiffusion 228 390 234 396 0 cell no = 599
<< m1 >>
rect 229 390 230 391 
rect 232 390 233 391 
rect 229 395 230 396 
rect 232 395 233 396 
<< m2 >>
rect 229 390 230 391 
rect 232 390 233 391 
rect 229 395 230 396 
rect 232 395 233 396 
<< m2c >>
rect 229 390 230 391 
rect 232 390 233 391 
rect 229 395 230 396 
rect 232 395 233 396 
<< labels >>
rlabel pdiffusion 49 426 50 427  0 t = 1
rlabel pdiffusion 52 426 53 427  0 t = 2
rlabel pdiffusion 49 431 50 432  0 t = 3
rlabel pdiffusion 52 431 53 432  0 t = 4
rlabel pdiffusion 48 426 54 432 0 cell no = 600
<< m1 >>
rect 49 426 50 427 
rect 52 426 53 427 
rect 49 431 50 432 
rect 52 431 53 432 
<< m2 >>
rect 49 426 50 427 
rect 52 426 53 427 
rect 49 431 50 432 
rect 52 431 53 432 
<< m2c >>
rect 49 426 50 427 
rect 52 426 53 427 
rect 49 431 50 432 
rect 52 431 53 432 
<< end >> 
