magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 23 0 24 1 
<< m2 >>
rect 23 0 24 1 
<< m2c >>
rect 23 0 24 1 
<< m1 >>
rect 23 0 24 1 
<< m2 >>
rect 23 0 24 1 
<< m1 >>
rect 24 0 25 1 
<< m1 >>
rect 25 0 26 1 
<< m1 >>
rect 26 0 27 1 
<< m1 >>
rect 27 0 28 1 
<< m1 >>
rect 28 0 29 1 
<< m1 >>
rect 29 0 30 1 
<< m1 >>
rect 30 0 31 1 
<< m1 >>
rect 31 0 32 1 
<< m1 >>
rect 32 0 33 1 
<< m1 >>
rect 33 0 34 1 
<< m1 >>
rect 34 0 35 1 
<< m1 >>
rect 35 0 36 1 
<< m1 >>
rect 36 0 37 1 
<< m1 >>
rect 37 0 38 1 
<< m1 >>
rect 38 0 39 1 
<< m1 >>
rect 39 0 40 1 
<< m1 >>
rect 40 0 41 1 
<< m1 >>
rect 41 0 42 1 
<< m1 >>
rect 42 0 43 1 
<< m1 >>
rect 43 0 44 1 
<< m1 >>
rect 44 0 45 1 
<< m1 >>
rect 45 0 46 1 
<< m1 >>
rect 46 0 47 1 
<< m1 >>
rect 47 0 48 1 
<< m1 >>
rect 48 0 49 1 
<< m1 >>
rect 49 0 50 1 
<< m1 >>
rect 50 0 51 1 
<< m1 >>
rect 51 0 52 1 
<< m1 >>
rect 52 0 53 1 
<< m1 >>
rect 53 0 54 1 
<< m1 >>
rect 54 0 55 1 
<< m1 >>
rect 55 0 56 1 
<< m1 >>
rect 56 0 57 1 
<< m1 >>
rect 57 0 58 1 
<< m1 >>
rect 58 0 59 1 
<< m1 >>
rect 59 0 60 1 
<< m1 >>
rect 60 0 61 1 
<< m1 >>
rect 61 0 62 1 
<< m1 >>
rect 62 0 63 1 
<< m1 >>
rect 63 0 64 1 
<< m1 >>
rect 64 0 65 1 
<< m1 >>
rect 65 0 66 1 
<< m1 >>
rect 66 0 67 1 
<< m1 >>
rect 67 0 68 1 
<< m1 >>
rect 68 0 69 1 
<< m1 >>
rect 69 0 70 1 
<< m1 >>
rect 70 0 71 1 
<< m1 >>
rect 71 0 72 1 
<< m1 >>
rect 72 0 73 1 
<< m1 >>
rect 73 0 74 1 
<< m1 >>
rect 74 0 75 1 
<< m1 >>
rect 75 0 76 1 
<< m1 >>
rect 76 0 77 1 
<< m1 >>
rect 77 0 78 1 
<< m1 >>
rect 78 0 79 1 
<< m1 >>
rect 79 0 80 1 
<< m1 >>
rect 80 0 81 1 
<< m1 >>
rect 81 0 82 1 
<< m1 >>
rect 82 0 83 1 
<< m1 >>
rect 83 0 84 1 
<< m1 >>
rect 84 0 85 1 
<< m1 >>
rect 85 0 86 1 
<< m1 >>
rect 86 0 87 1 
<< m1 >>
rect 87 0 88 1 
<< m1 >>
rect 88 0 89 1 
<< m1 >>
rect 89 0 90 1 
<< m1 >>
rect 90 0 91 1 
<< m1 >>
rect 91 0 92 1 
<< m1 >>
rect 92 0 93 1 
<< m1 >>
rect 93 0 94 1 
<< m1 >>
rect 94 0 95 1 
<< m1 >>
rect 95 0 96 1 
<< m1 >>
rect 96 0 97 1 
<< m1 >>
rect 97 0 98 1 
<< m1 >>
rect 98 0 99 1 
<< m1 >>
rect 99 0 100 1 
<< m1 >>
rect 100 0 101 1 
<< m1 >>
rect 101 0 102 1 
<< m1 >>
rect 102 0 103 1 
<< m1 >>
rect 103 0 104 1 
<< m1 >>
rect 104 0 105 1 
<< m1 >>
rect 105 0 106 1 
<< m1 >>
rect 106 0 107 1 
<< m1 >>
rect 107 0 108 1 
<< m1 >>
rect 108 0 109 1 
<< m1 >>
rect 109 0 110 1 
<< m1 >>
rect 110 0 111 1 
<< m1 >>
rect 111 0 112 1 
<< m1 >>
rect 112 0 113 1 
<< m1 >>
rect 113 0 114 1 
<< m1 >>
rect 114 0 115 1 
<< m1 >>
rect 115 0 116 1 
<< m1 >>
rect 116 0 117 1 
<< m1 >>
rect 117 0 118 1 
<< m1 >>
rect 118 0 119 1 
<< m1 >>
rect 119 0 120 1 
<< m1 >>
rect 120 0 121 1 
<< m1 >>
rect 121 0 122 1 
<< m1 >>
rect 122 0 123 1 
<< m1 >>
rect 123 0 124 1 
<< m1 >>
rect 124 0 125 1 
<< m1 >>
rect 125 0 126 1 
<< m1 >>
rect 126 0 127 1 
<< m1 >>
rect 127 0 128 1 
<< m1 >>
rect 128 0 129 1 
<< m1 >>
rect 129 0 130 1 
<< m1 >>
rect 130 0 131 1 
<< m1 >>
rect 131 0 132 1 
<< m1 >>
rect 132 0 133 1 
<< m1 >>
rect 133 0 134 1 
<< m1 >>
rect 134 0 135 1 
<< m1 >>
rect 135 0 136 1 
<< m1 >>
rect 136 0 137 1 
<< m1 >>
rect 137 0 138 1 
<< m1 >>
rect 138 0 139 1 
<< m1 >>
rect 139 0 140 1 
<< m1 >>
rect 140 0 141 1 
<< m1 >>
rect 141 0 142 1 
<< m1 >>
rect 142 0 143 1 
<< m1 >>
rect 143 0 144 1 
<< m1 >>
rect 144 0 145 1 
<< m1 >>
rect 145 0 146 1 
<< m1 >>
rect 146 0 147 1 
<< m1 >>
rect 147 0 148 1 
<< m1 >>
rect 148 0 149 1 
<< m1 >>
rect 149 0 150 1 
<< m1 >>
rect 150 0 151 1 
<< m1 >>
rect 151 0 152 1 
<< m1 >>
rect 152 0 153 1 
<< m1 >>
rect 153 0 154 1 
<< m1 >>
rect 154 0 155 1 
<< m1 >>
rect 155 0 156 1 
<< m1 >>
rect 156 0 157 1 
<< m1 >>
rect 157 0 158 1 
<< m1 >>
rect 158 0 159 1 
<< m1 >>
rect 159 0 160 1 
<< m1 >>
rect 160 0 161 1 
<< m1 >>
rect 161 0 162 1 
<< m1 >>
rect 162 0 163 1 
<< m1 >>
rect 163 0 164 1 
<< m1 >>
rect 164 0 165 1 
<< m1 >>
rect 165 0 166 1 
<< m1 >>
rect 166 0 167 1 
<< m1 >>
rect 167 0 168 1 
<< m1 >>
rect 168 0 169 1 
<< m1 >>
rect 169 0 170 1 
<< m1 >>
rect 170 0 171 1 
<< m1 >>
rect 171 0 172 1 
<< m1 >>
rect 172 0 173 1 
<< m1 >>
rect 173 0 174 1 
<< m1 >>
rect 174 0 175 1 
<< m1 >>
rect 175 0 176 1 
<< m1 >>
rect 176 0 177 1 
<< m1 >>
rect 177 0 178 1 
<< m1 >>
rect 178 0 179 1 
<< m1 >>
rect 179 0 180 1 
<< m1 >>
rect 180 0 181 1 
<< m1 >>
rect 181 0 182 1 
<< m1 >>
rect 182 0 183 1 
<< m1 >>
rect 183 0 184 1 
<< m1 >>
rect 184 0 185 1 
<< m1 >>
rect 185 0 186 1 
<< m1 >>
rect 186 0 187 1 
<< m1 >>
rect 187 0 188 1 
<< m1 >>
rect 188 0 189 1 
<< m1 >>
rect 189 0 190 1 
<< m1 >>
rect 190 0 191 1 
<< m1 >>
rect 191 0 192 1 
<< m1 >>
rect 192 0 193 1 
<< m1 >>
rect 193 0 194 1 
<< m1 >>
rect 194 0 195 1 
<< m1 >>
rect 195 0 196 1 
<< m1 >>
rect 196 0 197 1 
<< m1 >>
rect 197 0 198 1 
<< m1 >>
rect 198 0 199 1 
<< m1 >>
rect 199 0 200 1 
<< m1 >>
rect 200 0 201 1 
<< m1 >>
rect 201 0 202 1 
<< m1 >>
rect 202 0 203 1 
<< m1 >>
rect 203 0 204 1 
<< m1 >>
rect 204 0 205 1 
<< m1 >>
rect 205 0 206 1 
<< m1 >>
rect 206 0 207 1 
<< m1 >>
rect 207 0 208 1 
<< m1 >>
rect 208 0 209 1 
<< m1 >>
rect 209 0 210 1 
<< m1 >>
rect 210 0 211 1 
<< m1 >>
rect 211 0 212 1 
<< m1 >>
rect 212 0 213 1 
<< m1 >>
rect 213 0 214 1 
<< m1 >>
rect 214 0 215 1 
<< m1 >>
rect 215 0 216 1 
<< m1 >>
rect 216 0 217 1 
<< m1 >>
rect 217 0 218 1 
<< m1 >>
rect 218 0 219 1 
<< m1 >>
rect 219 0 220 1 
<< m1 >>
rect 220 0 221 1 
<< m1 >>
rect 221 0 222 1 
<< m1 >>
rect 222 0 223 1 
<< m1 >>
rect 223 0 224 1 
<< m1 >>
rect 224 0 225 1 
<< m1 >>
rect 225 0 226 1 
<< m1 >>
rect 226 0 227 1 
<< m1 >>
rect 227 0 228 1 
<< m1 >>
rect 228 0 229 1 
<< m1 >>
rect 229 0 230 1 
<< m1 >>
rect 230 0 231 1 
<< m1 >>
rect 231 0 232 1 
<< m1 >>
rect 232 0 233 1 
<< m1 >>
rect 233 0 234 1 
<< m1 >>
rect 234 0 235 1 
<< m1 >>
rect 235 0 236 1 
<< m1 >>
rect 236 0 237 1 
<< m1 >>
rect 237 0 238 1 
<< m1 >>
rect 238 0 239 1 
<< m1 >>
rect 239 0 240 1 
<< m1 >>
rect 240 0 241 1 
<< m1 >>
rect 241 0 242 1 
<< m1 >>
rect 242 0 243 1 
<< m1 >>
rect 243 0 244 1 
<< m1 >>
rect 244 0 245 1 
<< m1 >>
rect 245 0 246 1 
<< m1 >>
rect 246 0 247 1 
<< m1 >>
rect 247 0 248 1 
<< m1 >>
rect 248 0 249 1 
<< m1 >>
rect 249 0 250 1 
<< m1 >>
rect 250 0 251 1 
<< m1 >>
rect 251 0 252 1 
<< m1 >>
rect 252 0 253 1 
<< m1 >>
rect 253 0 254 1 
<< m1 >>
rect 254 0 255 1 
<< m1 >>
rect 255 0 256 1 
<< m1 >>
rect 256 0 257 1 
<< m1 >>
rect 257 0 258 1 
<< m1 >>
rect 258 0 259 1 
<< m1 >>
rect 259 0 260 1 
<< m1 >>
rect 260 0 261 1 
<< m1 >>
rect 261 0 262 1 
<< m1 >>
rect 262 0 263 1 
<< m1 >>
rect 263 0 264 1 
<< m1 >>
rect 264 0 265 1 
<< m1 >>
rect 265 0 266 1 
<< m1 >>
rect 266 0 267 1 
<< m1 >>
rect 267 0 268 1 
<< m1 >>
rect 268 0 269 1 
<< m1 >>
rect 269 0 270 1 
<< m1 >>
rect 270 0 271 1 
<< m1 >>
rect 271 0 272 1 
<< m1 >>
rect 272 0 273 1 
<< m2 >>
rect 272 0 273 1 
<< m2c >>
rect 272 0 273 1 
<< m1 >>
rect 272 0 273 1 
<< m2 >>
rect 272 0 273 1 
<< m2 >>
rect 23 1 24 2 
<< m2 >>
rect 272 1 273 2 
<< m1 >>
rect 21 2 22 3 
<< m1 >>
rect 22 2 23 3 
<< m1 >>
rect 23 2 24 3 
<< m2 >>
rect 23 2 24 3 
<< m1 >>
rect 24 2 25 3 
<< m1 >>
rect 25 2 26 3 
<< m1 >>
rect 26 2 27 3 
<< m1 >>
rect 27 2 28 3 
<< m1 >>
rect 28 2 29 3 
<< m1 >>
rect 29 2 30 3 
<< m1 >>
rect 30 2 31 3 
<< m1 >>
rect 31 2 32 3 
<< m1 >>
rect 32 2 33 3 
<< m1 >>
rect 33 2 34 3 
<< m1 >>
rect 34 2 35 3 
<< m1 >>
rect 35 2 36 3 
<< m1 >>
rect 36 2 37 3 
<< m1 >>
rect 37 2 38 3 
<< m1 >>
rect 38 2 39 3 
<< m1 >>
rect 39 2 40 3 
<< m1 >>
rect 40 2 41 3 
<< m1 >>
rect 41 2 42 3 
<< m1 >>
rect 42 2 43 3 
<< m1 >>
rect 43 2 44 3 
<< m1 >>
rect 44 2 45 3 
<< m1 >>
rect 45 2 46 3 
<< m1 >>
rect 46 2 47 3 
<< m2 >>
rect 46 2 47 3 
<< m1 >>
rect 47 2 48 3 
<< m2 >>
rect 47 2 48 3 
<< m1 >>
rect 48 2 49 3 
<< m2 >>
rect 48 2 49 3 
<< m1 >>
rect 49 2 50 3 
<< m2 >>
rect 49 2 50 3 
<< m1 >>
rect 50 2 51 3 
<< m2 >>
rect 50 2 51 3 
<< m1 >>
rect 51 2 52 3 
<< m2 >>
rect 51 2 52 3 
<< m1 >>
rect 52 2 53 3 
<< m2 >>
rect 52 2 53 3 
<< m1 >>
rect 53 2 54 3 
<< m2 >>
rect 53 2 54 3 
<< m1 >>
rect 54 2 55 3 
<< m2 >>
rect 54 2 55 3 
<< m1 >>
rect 55 2 56 3 
<< m2 >>
rect 55 2 56 3 
<< m1 >>
rect 56 2 57 3 
<< m2 >>
rect 56 2 57 3 
<< m1 >>
rect 57 2 58 3 
<< m2 >>
rect 57 2 58 3 
<< m1 >>
rect 58 2 59 3 
<< m2 >>
rect 58 2 59 3 
<< m1 >>
rect 59 2 60 3 
<< m2 >>
rect 59 2 60 3 
<< m1 >>
rect 60 2 61 3 
<< m2 >>
rect 60 2 61 3 
<< m1 >>
rect 61 2 62 3 
<< m2 >>
rect 61 2 62 3 
<< m1 >>
rect 62 2 63 3 
<< m2 >>
rect 62 2 63 3 
<< m1 >>
rect 63 2 64 3 
<< m2 >>
rect 63 2 64 3 
<< m1 >>
rect 64 2 65 3 
<< m2 >>
rect 64 2 65 3 
<< m1 >>
rect 65 2 66 3 
<< m2 >>
rect 65 2 66 3 
<< m1 >>
rect 66 2 67 3 
<< m2 >>
rect 66 2 67 3 
<< m1 >>
rect 67 2 68 3 
<< m2 >>
rect 67 2 68 3 
<< m1 >>
rect 68 2 69 3 
<< m2 >>
rect 68 2 69 3 
<< m1 >>
rect 69 2 70 3 
<< m2 >>
rect 69 2 70 3 
<< m1 >>
rect 70 2 71 3 
<< m2 >>
rect 70 2 71 3 
<< m1 >>
rect 71 2 72 3 
<< m2 >>
rect 71 2 72 3 
<< m1 >>
rect 72 2 73 3 
<< m2 >>
rect 72 2 73 3 
<< m1 >>
rect 73 2 74 3 
<< m2 >>
rect 73 2 74 3 
<< m1 >>
rect 74 2 75 3 
<< m2 >>
rect 74 2 75 3 
<< m1 >>
rect 75 2 76 3 
<< m2 >>
rect 75 2 76 3 
<< m1 >>
rect 76 2 77 3 
<< m2 >>
rect 76 2 77 3 
<< m1 >>
rect 77 2 78 3 
<< m2 >>
rect 77 2 78 3 
<< m1 >>
rect 78 2 79 3 
<< m2 >>
rect 78 2 79 3 
<< m1 >>
rect 79 2 80 3 
<< m2 >>
rect 79 2 80 3 
<< m1 >>
rect 80 2 81 3 
<< m2 >>
rect 80 2 81 3 
<< m1 >>
rect 81 2 82 3 
<< m2 >>
rect 81 2 82 3 
<< m1 >>
rect 82 2 83 3 
<< m2 >>
rect 82 2 83 3 
<< m1 >>
rect 83 2 84 3 
<< m2 >>
rect 83 2 84 3 
<< m1 >>
rect 84 2 85 3 
<< m2 >>
rect 84 2 85 3 
<< m1 >>
rect 85 2 86 3 
<< m2 >>
rect 85 2 86 3 
<< m1 >>
rect 86 2 87 3 
<< m2 >>
rect 86 2 87 3 
<< m1 >>
rect 87 2 88 3 
<< m2 >>
rect 87 2 88 3 
<< m1 >>
rect 88 2 89 3 
<< m2 >>
rect 88 2 89 3 
<< m1 >>
rect 89 2 90 3 
<< m2 >>
rect 89 2 90 3 
<< m1 >>
rect 90 2 91 3 
<< m2 >>
rect 90 2 91 3 
<< m1 >>
rect 91 2 92 3 
<< m2 >>
rect 91 2 92 3 
<< m1 >>
rect 92 2 93 3 
<< m2 >>
rect 92 2 93 3 
<< m1 >>
rect 93 2 94 3 
<< m2 >>
rect 93 2 94 3 
<< m1 >>
rect 94 2 95 3 
<< m2 >>
rect 94 2 95 3 
<< m1 >>
rect 95 2 96 3 
<< m2 >>
rect 95 2 96 3 
<< m1 >>
rect 96 2 97 3 
<< m2 >>
rect 96 2 97 3 
<< m1 >>
rect 97 2 98 3 
<< m2 >>
rect 97 2 98 3 
<< m1 >>
rect 98 2 99 3 
<< m2 >>
rect 98 2 99 3 
<< m1 >>
rect 99 2 100 3 
<< m2 >>
rect 99 2 100 3 
<< m1 >>
rect 100 2 101 3 
<< m2 >>
rect 100 2 101 3 
<< m1 >>
rect 101 2 102 3 
<< m2 >>
rect 101 2 102 3 
<< m1 >>
rect 102 2 103 3 
<< m2 >>
rect 102 2 103 3 
<< m1 >>
rect 103 2 104 3 
<< m2 >>
rect 103 2 104 3 
<< m1 >>
rect 104 2 105 3 
<< m2 >>
rect 104 2 105 3 
<< m1 >>
rect 105 2 106 3 
<< m2 >>
rect 105 2 106 3 
<< m1 >>
rect 106 2 107 3 
<< m2 >>
rect 106 2 107 3 
<< m1 >>
rect 107 2 108 3 
<< m2 >>
rect 107 2 108 3 
<< m1 >>
rect 108 2 109 3 
<< m2 >>
rect 108 2 109 3 
<< m1 >>
rect 109 2 110 3 
<< m2 >>
rect 109 2 110 3 
<< m1 >>
rect 110 2 111 3 
<< m2 >>
rect 110 2 111 3 
<< m1 >>
rect 111 2 112 3 
<< m2 >>
rect 111 2 112 3 
<< m1 >>
rect 112 2 113 3 
<< m2 >>
rect 112 2 113 3 
<< m1 >>
rect 113 2 114 3 
<< m2 >>
rect 113 2 114 3 
<< m1 >>
rect 114 2 115 3 
<< m2 >>
rect 114 2 115 3 
<< m1 >>
rect 115 2 116 3 
<< m2 >>
rect 115 2 116 3 
<< m1 >>
rect 116 2 117 3 
<< m2 >>
rect 116 2 117 3 
<< m1 >>
rect 117 2 118 3 
<< m2 >>
rect 117 2 118 3 
<< m1 >>
rect 118 2 119 3 
<< m2 >>
rect 118 2 119 3 
<< m1 >>
rect 119 2 120 3 
<< m2 >>
rect 119 2 120 3 
<< m1 >>
rect 120 2 121 3 
<< m2 >>
rect 120 2 121 3 
<< m1 >>
rect 121 2 122 3 
<< m2 >>
rect 121 2 122 3 
<< m1 >>
rect 122 2 123 3 
<< m2 >>
rect 122 2 123 3 
<< m1 >>
rect 123 2 124 3 
<< m2 >>
rect 123 2 124 3 
<< m1 >>
rect 124 2 125 3 
<< m2 >>
rect 124 2 125 3 
<< m1 >>
rect 125 2 126 3 
<< m2 >>
rect 125 2 126 3 
<< m1 >>
rect 126 2 127 3 
<< m2 >>
rect 126 2 127 3 
<< m1 >>
rect 127 2 128 3 
<< m2 >>
rect 127 2 128 3 
<< m1 >>
rect 128 2 129 3 
<< m2 >>
rect 128 2 129 3 
<< m1 >>
rect 129 2 130 3 
<< m2 >>
rect 129 2 130 3 
<< m1 >>
rect 130 2 131 3 
<< m2 >>
rect 130 2 131 3 
<< m1 >>
rect 131 2 132 3 
<< m2 >>
rect 131 2 132 3 
<< m1 >>
rect 132 2 133 3 
<< m2 >>
rect 132 2 133 3 
<< m1 >>
rect 133 2 134 3 
<< m2 >>
rect 133 2 134 3 
<< m1 >>
rect 134 2 135 3 
<< m2 >>
rect 134 2 135 3 
<< m1 >>
rect 135 2 136 3 
<< m2 >>
rect 135 2 136 3 
<< m1 >>
rect 136 2 137 3 
<< m2 >>
rect 136 2 137 3 
<< m1 >>
rect 137 2 138 3 
<< m2 >>
rect 137 2 138 3 
<< m1 >>
rect 138 2 139 3 
<< m2 >>
rect 138 2 139 3 
<< m1 >>
rect 139 2 140 3 
<< m2 >>
rect 139 2 140 3 
<< m1 >>
rect 140 2 141 3 
<< m2 >>
rect 140 2 141 3 
<< m1 >>
rect 141 2 142 3 
<< m2 >>
rect 141 2 142 3 
<< m1 >>
rect 142 2 143 3 
<< m2 >>
rect 142 2 143 3 
<< m1 >>
rect 143 2 144 3 
<< m2 >>
rect 143 2 144 3 
<< m1 >>
rect 144 2 145 3 
<< m2 >>
rect 144 2 145 3 
<< m1 >>
rect 145 2 146 3 
<< m2 >>
rect 145 2 146 3 
<< m1 >>
rect 146 2 147 3 
<< m2 >>
rect 146 2 147 3 
<< m1 >>
rect 147 2 148 3 
<< m2 >>
rect 147 2 148 3 
<< m1 >>
rect 148 2 149 3 
<< m2 >>
rect 148 2 149 3 
<< m1 >>
rect 149 2 150 3 
<< m2 >>
rect 149 2 150 3 
<< m1 >>
rect 150 2 151 3 
<< m2 >>
rect 150 2 151 3 
<< m1 >>
rect 151 2 152 3 
<< m2 >>
rect 151 2 152 3 
<< m1 >>
rect 152 2 153 3 
<< m2 >>
rect 152 2 153 3 
<< m1 >>
rect 153 2 154 3 
<< m2 >>
rect 153 2 154 3 
<< m1 >>
rect 154 2 155 3 
<< m2 >>
rect 154 2 155 3 
<< m1 >>
rect 155 2 156 3 
<< m2 >>
rect 155 2 156 3 
<< m1 >>
rect 156 2 157 3 
<< m2 >>
rect 156 2 157 3 
<< m1 >>
rect 157 2 158 3 
<< m2 >>
rect 157 2 158 3 
<< m1 >>
rect 158 2 159 3 
<< m2 >>
rect 158 2 159 3 
<< m1 >>
rect 159 2 160 3 
<< m2 >>
rect 159 2 160 3 
<< m1 >>
rect 160 2 161 3 
<< m2 >>
rect 160 2 161 3 
<< m1 >>
rect 161 2 162 3 
<< m2 >>
rect 161 2 162 3 
<< m1 >>
rect 162 2 163 3 
<< m2 >>
rect 162 2 163 3 
<< m1 >>
rect 163 2 164 3 
<< m2 >>
rect 163 2 164 3 
<< m1 >>
rect 164 2 165 3 
<< m2 >>
rect 164 2 165 3 
<< m1 >>
rect 165 2 166 3 
<< m2 >>
rect 165 2 166 3 
<< m1 >>
rect 166 2 167 3 
<< m2 >>
rect 166 2 167 3 
<< m1 >>
rect 167 2 168 3 
<< m2 >>
rect 167 2 168 3 
<< m1 >>
rect 168 2 169 3 
<< m2 >>
rect 168 2 169 3 
<< m1 >>
rect 169 2 170 3 
<< m2 >>
rect 169 2 170 3 
<< m1 >>
rect 170 2 171 3 
<< m2 >>
rect 170 2 171 3 
<< m1 >>
rect 171 2 172 3 
<< m2 >>
rect 171 2 172 3 
<< m1 >>
rect 172 2 173 3 
<< m2 >>
rect 172 2 173 3 
<< m1 >>
rect 173 2 174 3 
<< m2 >>
rect 173 2 174 3 
<< m1 >>
rect 174 2 175 3 
<< m2 >>
rect 174 2 175 3 
<< m1 >>
rect 175 2 176 3 
<< m2 >>
rect 175 2 176 3 
<< m1 >>
rect 176 2 177 3 
<< m2 >>
rect 176 2 177 3 
<< m1 >>
rect 177 2 178 3 
<< m2 >>
rect 177 2 178 3 
<< m1 >>
rect 178 2 179 3 
<< m2 >>
rect 178 2 179 3 
<< m1 >>
rect 179 2 180 3 
<< m2 >>
rect 179 2 180 3 
<< m1 >>
rect 180 2 181 3 
<< m2 >>
rect 180 2 181 3 
<< m1 >>
rect 181 2 182 3 
<< m2 >>
rect 181 2 182 3 
<< m1 >>
rect 182 2 183 3 
<< m2 >>
rect 182 2 183 3 
<< m1 >>
rect 183 2 184 3 
<< m2 >>
rect 183 2 184 3 
<< m1 >>
rect 184 2 185 3 
<< m2 >>
rect 184 2 185 3 
<< m1 >>
rect 185 2 186 3 
<< m2 >>
rect 185 2 186 3 
<< m1 >>
rect 186 2 187 3 
<< m2 >>
rect 186 2 187 3 
<< m1 >>
rect 187 2 188 3 
<< m2 >>
rect 187 2 188 3 
<< m1 >>
rect 188 2 189 3 
<< m2 >>
rect 188 2 189 3 
<< m1 >>
rect 189 2 190 3 
<< m2 >>
rect 189 2 190 3 
<< m1 >>
rect 190 2 191 3 
<< m2 >>
rect 190 2 191 3 
<< m1 >>
rect 191 2 192 3 
<< m2 >>
rect 191 2 192 3 
<< m1 >>
rect 192 2 193 3 
<< m2 >>
rect 192 2 193 3 
<< m1 >>
rect 193 2 194 3 
<< m2 >>
rect 193 2 194 3 
<< m1 >>
rect 194 2 195 3 
<< m2 >>
rect 194 2 195 3 
<< m1 >>
rect 195 2 196 3 
<< m2 >>
rect 195 2 196 3 
<< m1 >>
rect 196 2 197 3 
<< m2 >>
rect 196 2 197 3 
<< m1 >>
rect 197 2 198 3 
<< m2 >>
rect 197 2 198 3 
<< m1 >>
rect 198 2 199 3 
<< m2 >>
rect 198 2 199 3 
<< m1 >>
rect 199 2 200 3 
<< m2 >>
rect 199 2 200 3 
<< m1 >>
rect 200 2 201 3 
<< m2 >>
rect 200 2 201 3 
<< m1 >>
rect 201 2 202 3 
<< m2 >>
rect 201 2 202 3 
<< m1 >>
rect 202 2 203 3 
<< m2 >>
rect 202 2 203 3 
<< m1 >>
rect 203 2 204 3 
<< m2 >>
rect 203 2 204 3 
<< m1 >>
rect 204 2 205 3 
<< m2 >>
rect 204 2 205 3 
<< m1 >>
rect 205 2 206 3 
<< m2 >>
rect 205 2 206 3 
<< m1 >>
rect 206 2 207 3 
<< m2 >>
rect 206 2 207 3 
<< m1 >>
rect 207 2 208 3 
<< m2 >>
rect 207 2 208 3 
<< m1 >>
rect 208 2 209 3 
<< m2 >>
rect 208 2 209 3 
<< m1 >>
rect 209 2 210 3 
<< m2 >>
rect 209 2 210 3 
<< m1 >>
rect 210 2 211 3 
<< m2 >>
rect 210 2 211 3 
<< m1 >>
rect 211 2 212 3 
<< m2 >>
rect 211 2 212 3 
<< m1 >>
rect 212 2 213 3 
<< m2 >>
rect 212 2 213 3 
<< m1 >>
rect 213 2 214 3 
<< m2 >>
rect 213 2 214 3 
<< m1 >>
rect 214 2 215 3 
<< m2 >>
rect 214 2 215 3 
<< m1 >>
rect 215 2 216 3 
<< m2 >>
rect 215 2 216 3 
<< m1 >>
rect 216 2 217 3 
<< m2 >>
rect 216 2 217 3 
<< m1 >>
rect 217 2 218 3 
<< m2 >>
rect 217 2 218 3 
<< m1 >>
rect 218 2 219 3 
<< m2 >>
rect 218 2 219 3 
<< m1 >>
rect 219 2 220 3 
<< m2 >>
rect 219 2 220 3 
<< m1 >>
rect 220 2 221 3 
<< m2 >>
rect 220 2 221 3 
<< m1 >>
rect 221 2 222 3 
<< m2 >>
rect 221 2 222 3 
<< m1 >>
rect 222 2 223 3 
<< m2 >>
rect 222 2 223 3 
<< m1 >>
rect 223 2 224 3 
<< m2 >>
rect 223 2 224 3 
<< m1 >>
rect 224 2 225 3 
<< m2 >>
rect 224 2 225 3 
<< m1 >>
rect 225 2 226 3 
<< m2 >>
rect 225 2 226 3 
<< m1 >>
rect 226 2 227 3 
<< m2 >>
rect 226 2 227 3 
<< m1 >>
rect 227 2 228 3 
<< m2 >>
rect 227 2 228 3 
<< m1 >>
rect 228 2 229 3 
<< m2 >>
rect 228 2 229 3 
<< m1 >>
rect 229 2 230 3 
<< m2 >>
rect 229 2 230 3 
<< m1 >>
rect 230 2 231 3 
<< m2 >>
rect 230 2 231 3 
<< m1 >>
rect 231 2 232 3 
<< m2 >>
rect 231 2 232 3 
<< m1 >>
rect 232 2 233 3 
<< m2 >>
rect 232 2 233 3 
<< m1 >>
rect 233 2 234 3 
<< m2 >>
rect 233 2 234 3 
<< m1 >>
rect 234 2 235 3 
<< m2 >>
rect 234 2 235 3 
<< m1 >>
rect 235 2 236 3 
<< m2 >>
rect 235 2 236 3 
<< m1 >>
rect 236 2 237 3 
<< m2 >>
rect 236 2 237 3 
<< m1 >>
rect 237 2 238 3 
<< m2 >>
rect 237 2 238 3 
<< m1 >>
rect 238 2 239 3 
<< m2 >>
rect 238 2 239 3 
<< m1 >>
rect 239 2 240 3 
<< m2 >>
rect 239 2 240 3 
<< m1 >>
rect 240 2 241 3 
<< m2 >>
rect 240 2 241 3 
<< m1 >>
rect 241 2 242 3 
<< m2 >>
rect 241 2 242 3 
<< m1 >>
rect 242 2 243 3 
<< m2 >>
rect 242 2 243 3 
<< m1 >>
rect 243 2 244 3 
<< m2 >>
rect 243 2 244 3 
<< m1 >>
rect 244 2 245 3 
<< m2 >>
rect 244 2 245 3 
<< m1 >>
rect 245 2 246 3 
<< m2 >>
rect 245 2 246 3 
<< m1 >>
rect 246 2 247 3 
<< m2 >>
rect 246 2 247 3 
<< m1 >>
rect 247 2 248 3 
<< m2 >>
rect 247 2 248 3 
<< m1 >>
rect 248 2 249 3 
<< m2 >>
rect 248 2 249 3 
<< m1 >>
rect 249 2 250 3 
<< m2 >>
rect 249 2 250 3 
<< m1 >>
rect 250 2 251 3 
<< m2 >>
rect 250 2 251 3 
<< m1 >>
rect 251 2 252 3 
<< m2 >>
rect 251 2 252 3 
<< m1 >>
rect 252 2 253 3 
<< m2 >>
rect 252 2 253 3 
<< m1 >>
rect 253 2 254 3 
<< m2 >>
rect 253 2 254 3 
<< m1 >>
rect 254 2 255 3 
<< m2 >>
rect 254 2 255 3 
<< m1 >>
rect 255 2 256 3 
<< m2 >>
rect 255 2 256 3 
<< m1 >>
rect 256 2 257 3 
<< m2 >>
rect 256 2 257 3 
<< m1 >>
rect 257 2 258 3 
<< m2 >>
rect 257 2 258 3 
<< m1 >>
rect 258 2 259 3 
<< m2 >>
rect 258 2 259 3 
<< m1 >>
rect 259 2 260 3 
<< m2 >>
rect 259 2 260 3 
<< m1 >>
rect 260 2 261 3 
<< m2 >>
rect 260 2 261 3 
<< m1 >>
rect 261 2 262 3 
<< m2 >>
rect 261 2 262 3 
<< m1 >>
rect 262 2 263 3 
<< m2 >>
rect 262 2 263 3 
<< m1 >>
rect 263 2 264 3 
<< m2 >>
rect 263 2 264 3 
<< m1 >>
rect 264 2 265 3 
<< m2 >>
rect 264 2 265 3 
<< m1 >>
rect 265 2 266 3 
<< m2 >>
rect 265 2 266 3 
<< m1 >>
rect 266 2 267 3 
<< m2 >>
rect 266 2 267 3 
<< m1 >>
rect 267 2 268 3 
<< m2 >>
rect 267 2 268 3 
<< m1 >>
rect 268 2 269 3 
<< m2 >>
rect 268 2 269 3 
<< m1 >>
rect 269 2 270 3 
<< m2 >>
rect 269 2 270 3 
<< m1 >>
rect 270 2 271 3 
<< m2 >>
rect 270 2 271 3 
<< m1 >>
rect 271 2 272 3 
<< m1 >>
rect 272 2 273 3 
<< m2 >>
rect 272 2 273 3 
<< m1 >>
rect 273 2 274 3 
<< m1 >>
rect 274 2 275 3 
<< m1 >>
rect 275 2 276 3 
<< m1 >>
rect 276 2 277 3 
<< m1 >>
rect 277 2 278 3 
<< m1 >>
rect 278 2 279 3 
<< m1 >>
rect 279 2 280 3 
<< m1 >>
rect 280 2 281 3 
<< m1 >>
rect 281 2 282 3 
<< m1 >>
rect 282 2 283 3 
<< m1 >>
rect 283 2 284 3 
<< m1 >>
rect 284 2 285 3 
<< m1 >>
rect 285 2 286 3 
<< m1 >>
rect 286 2 287 3 
<< m1 >>
rect 287 2 288 3 
<< m1 >>
rect 288 2 289 3 
<< m1 >>
rect 289 2 290 3 
<< m1 >>
rect 290 2 291 3 
<< m1 >>
rect 291 2 292 3 
<< m1 >>
rect 292 2 293 3 
<< m1 >>
rect 293 2 294 3 
<< m1 >>
rect 294 2 295 3 
<< m1 >>
rect 295 2 296 3 
<< m1 >>
rect 296 2 297 3 
<< m1 >>
rect 297 2 298 3 
<< m1 >>
rect 298 2 299 3 
<< m1 >>
rect 299 2 300 3 
<< m1 >>
rect 300 2 301 3 
<< m1 >>
rect 301 2 302 3 
<< m1 >>
rect 302 2 303 3 
<< m1 >>
rect 303 2 304 3 
<< m1 >>
rect 304 2 305 3 
<< m1 >>
rect 305 2 306 3 
<< m1 >>
rect 306 2 307 3 
<< m1 >>
rect 307 2 308 3 
<< m1 >>
rect 308 2 309 3 
<< m1 >>
rect 309 2 310 3 
<< m1 >>
rect 310 2 311 3 
<< m1 >>
rect 311 2 312 3 
<< m1 >>
rect 312 2 313 3 
<< m1 >>
rect 313 2 314 3 
<< m1 >>
rect 314 2 315 3 
<< m1 >>
rect 315 2 316 3 
<< m1 >>
rect 316 2 317 3 
<< m1 >>
rect 317 2 318 3 
<< m1 >>
rect 318 2 319 3 
<< m1 >>
rect 319 2 320 3 
<< m1 >>
rect 320 2 321 3 
<< m1 >>
rect 321 2 322 3 
<< m1 >>
rect 322 2 323 3 
<< m1 >>
rect 323 2 324 3 
<< m1 >>
rect 324 2 325 3 
<< m1 >>
rect 325 2 326 3 
<< m1 >>
rect 326 2 327 3 
<< m1 >>
rect 327 2 328 3 
<< m1 >>
rect 328 2 329 3 
<< m1 >>
rect 329 2 330 3 
<< m1 >>
rect 330 2 331 3 
<< m1 >>
rect 331 2 332 3 
<< m1 >>
rect 332 2 333 3 
<< m1 >>
rect 333 2 334 3 
<< m1 >>
rect 334 2 335 3 
<< m1 >>
rect 335 2 336 3 
<< m1 >>
rect 336 2 337 3 
<< m1 >>
rect 337 2 338 3 
<< m1 >>
rect 338 2 339 3 
<< m1 >>
rect 339 2 340 3 
<< m1 >>
rect 340 2 341 3 
<< m1 >>
rect 341 2 342 3 
<< m1 >>
rect 342 2 343 3 
<< m1 >>
rect 343 2 344 3 
<< m1 >>
rect 21 3 22 4 
<< m2 >>
rect 23 3 24 4 
<< m2 >>
rect 46 3 47 4 
<< m2 >>
rect 270 3 271 4 
<< m2 >>
rect 272 3 273 4 
<< m1 >>
rect 343 3 344 4 
<< m1 >>
rect 21 4 22 5 
<< m1 >>
rect 23 4 24 5 
<< m2 >>
rect 23 4 24 5 
<< m2c >>
rect 23 4 24 5 
<< m1 >>
rect 23 4 24 5 
<< m2 >>
rect 23 4 24 5 
<< m1 >>
rect 46 4 47 5 
<< m2 >>
rect 46 4 47 5 
<< m2c >>
rect 46 4 47 5 
<< m1 >>
rect 46 4 47 5 
<< m2 >>
rect 46 4 47 5 
<< m1 >>
rect 62 4 63 5 
<< m2 >>
rect 62 4 63 5 
<< m2c >>
rect 62 4 63 5 
<< m1 >>
rect 62 4 63 5 
<< m2 >>
rect 62 4 63 5 
<< m1 >>
rect 63 4 64 5 
<< m1 >>
rect 64 4 65 5 
<< m1 >>
rect 65 4 66 5 
<< m1 >>
rect 66 4 67 5 
<< m1 >>
rect 67 4 68 5 
<< m1 >>
rect 68 4 69 5 
<< m1 >>
rect 69 4 70 5 
<< m1 >>
rect 70 4 71 5 
<< m1 >>
rect 71 4 72 5 
<< m1 >>
rect 72 4 73 5 
<< m1 >>
rect 73 4 74 5 
<< m1 >>
rect 74 4 75 5 
<< m1 >>
rect 75 4 76 5 
<< m1 >>
rect 76 4 77 5 
<< m1 >>
rect 77 4 78 5 
<< m1 >>
rect 78 4 79 5 
<< m1 >>
rect 79 4 80 5 
<< m1 >>
rect 80 4 81 5 
<< m1 >>
rect 81 4 82 5 
<< m1 >>
rect 82 4 83 5 
<< m1 >>
rect 83 4 84 5 
<< m1 >>
rect 84 4 85 5 
<< m1 >>
rect 85 4 86 5 
<< m1 >>
rect 86 4 87 5 
<< m1 >>
rect 87 4 88 5 
<< m1 >>
rect 88 4 89 5 
<< m1 >>
rect 89 4 90 5 
<< m1 >>
rect 90 4 91 5 
<< m1 >>
rect 91 4 92 5 
<< m1 >>
rect 92 4 93 5 
<< m1 >>
rect 93 4 94 5 
<< m1 >>
rect 94 4 95 5 
<< m1 >>
rect 95 4 96 5 
<< m1 >>
rect 96 4 97 5 
<< m1 >>
rect 97 4 98 5 
<< m1 >>
rect 98 4 99 5 
<< m1 >>
rect 99 4 100 5 
<< m1 >>
rect 100 4 101 5 
<< m1 >>
rect 101 4 102 5 
<< m1 >>
rect 102 4 103 5 
<< m1 >>
rect 103 4 104 5 
<< m1 >>
rect 104 4 105 5 
<< m1 >>
rect 105 4 106 5 
<< m1 >>
rect 106 4 107 5 
<< m1 >>
rect 107 4 108 5 
<< m1 >>
rect 108 4 109 5 
<< m1 >>
rect 109 4 110 5 
<< m1 >>
rect 110 4 111 5 
<< m1 >>
rect 111 4 112 5 
<< m1 >>
rect 112 4 113 5 
<< m1 >>
rect 113 4 114 5 
<< m1 >>
rect 114 4 115 5 
<< m1 >>
rect 115 4 116 5 
<< m1 >>
rect 116 4 117 5 
<< m1 >>
rect 117 4 118 5 
<< m1 >>
rect 118 4 119 5 
<< m1 >>
rect 119 4 120 5 
<< m1 >>
rect 120 4 121 5 
<< m1 >>
rect 121 4 122 5 
<< m1 >>
rect 122 4 123 5 
<< m1 >>
rect 123 4 124 5 
<< m1 >>
rect 124 4 125 5 
<< m1 >>
rect 125 4 126 5 
<< m1 >>
rect 126 4 127 5 
<< m1 >>
rect 127 4 128 5 
<< m1 >>
rect 128 4 129 5 
<< m1 >>
rect 129 4 130 5 
<< m1 >>
rect 130 4 131 5 
<< m1 >>
rect 131 4 132 5 
<< m1 >>
rect 132 4 133 5 
<< m1 >>
rect 133 4 134 5 
<< m1 >>
rect 134 4 135 5 
<< m1 >>
rect 135 4 136 5 
<< m1 >>
rect 136 4 137 5 
<< m1 >>
rect 137 4 138 5 
<< m1 >>
rect 138 4 139 5 
<< m1 >>
rect 139 4 140 5 
<< m1 >>
rect 140 4 141 5 
<< m1 >>
rect 141 4 142 5 
<< m1 >>
rect 142 4 143 5 
<< m1 >>
rect 143 4 144 5 
<< m1 >>
rect 144 4 145 5 
<< m1 >>
rect 145 4 146 5 
<< m1 >>
rect 146 4 147 5 
<< m1 >>
rect 147 4 148 5 
<< m1 >>
rect 148 4 149 5 
<< m1 >>
rect 149 4 150 5 
<< m1 >>
rect 150 4 151 5 
<< m1 >>
rect 151 4 152 5 
<< m1 >>
rect 152 4 153 5 
<< m1 >>
rect 153 4 154 5 
<< m1 >>
rect 154 4 155 5 
<< m1 >>
rect 155 4 156 5 
<< m1 >>
rect 156 4 157 5 
<< m1 >>
rect 157 4 158 5 
<< m1 >>
rect 158 4 159 5 
<< m1 >>
rect 159 4 160 5 
<< m1 >>
rect 160 4 161 5 
<< m1 >>
rect 161 4 162 5 
<< m1 >>
rect 162 4 163 5 
<< m1 >>
rect 163 4 164 5 
<< m1 >>
rect 164 4 165 5 
<< m1 >>
rect 165 4 166 5 
<< m1 >>
rect 166 4 167 5 
<< m1 >>
rect 167 4 168 5 
<< m1 >>
rect 168 4 169 5 
<< m1 >>
rect 169 4 170 5 
<< m1 >>
rect 170 4 171 5 
<< m1 >>
rect 171 4 172 5 
<< m1 >>
rect 172 4 173 5 
<< m1 >>
rect 173 4 174 5 
<< m1 >>
rect 174 4 175 5 
<< m1 >>
rect 175 4 176 5 
<< m1 >>
rect 176 4 177 5 
<< m1 >>
rect 177 4 178 5 
<< m1 >>
rect 178 4 179 5 
<< m1 >>
rect 179 4 180 5 
<< m1 >>
rect 180 4 181 5 
<< m1 >>
rect 181 4 182 5 
<< m1 >>
rect 182 4 183 5 
<< m1 >>
rect 183 4 184 5 
<< m1 >>
rect 184 4 185 5 
<< m1 >>
rect 185 4 186 5 
<< m1 >>
rect 186 4 187 5 
<< m1 >>
rect 187 4 188 5 
<< m1 >>
rect 188 4 189 5 
<< m1 >>
rect 189 4 190 5 
<< m1 >>
rect 190 4 191 5 
<< m1 >>
rect 191 4 192 5 
<< m1 >>
rect 192 4 193 5 
<< m1 >>
rect 193 4 194 5 
<< m1 >>
rect 194 4 195 5 
<< m1 >>
rect 195 4 196 5 
<< m1 >>
rect 196 4 197 5 
<< m1 >>
rect 197 4 198 5 
<< m1 >>
rect 198 4 199 5 
<< m1 >>
rect 199 4 200 5 
<< m1 >>
rect 200 4 201 5 
<< m1 >>
rect 201 4 202 5 
<< m1 >>
rect 202 4 203 5 
<< m1 >>
rect 203 4 204 5 
<< m1 >>
rect 204 4 205 5 
<< m1 >>
rect 205 4 206 5 
<< m1 >>
rect 206 4 207 5 
<< m1 >>
rect 207 4 208 5 
<< m1 >>
rect 208 4 209 5 
<< m1 >>
rect 209 4 210 5 
<< m1 >>
rect 210 4 211 5 
<< m1 >>
rect 211 4 212 5 
<< m1 >>
rect 212 4 213 5 
<< m1 >>
rect 213 4 214 5 
<< m1 >>
rect 214 4 215 5 
<< m1 >>
rect 215 4 216 5 
<< m1 >>
rect 216 4 217 5 
<< m1 >>
rect 217 4 218 5 
<< m1 >>
rect 218 4 219 5 
<< m1 >>
rect 219 4 220 5 
<< m1 >>
rect 220 4 221 5 
<< m1 >>
rect 221 4 222 5 
<< m1 >>
rect 222 4 223 5 
<< m1 >>
rect 223 4 224 5 
<< m1 >>
rect 224 4 225 5 
<< m1 >>
rect 225 4 226 5 
<< m1 >>
rect 226 4 227 5 
<< m1 >>
rect 227 4 228 5 
<< m1 >>
rect 228 4 229 5 
<< m1 >>
rect 229 4 230 5 
<< m1 >>
rect 230 4 231 5 
<< m1 >>
rect 231 4 232 5 
<< m1 >>
rect 232 4 233 5 
<< m1 >>
rect 233 4 234 5 
<< m1 >>
rect 234 4 235 5 
<< m1 >>
rect 235 4 236 5 
<< m1 >>
rect 236 4 237 5 
<< m1 >>
rect 237 4 238 5 
<< m1 >>
rect 238 4 239 5 
<< m1 >>
rect 239 4 240 5 
<< m1 >>
rect 240 4 241 5 
<< m1 >>
rect 241 4 242 5 
<< m1 >>
rect 242 4 243 5 
<< m1 >>
rect 243 4 244 5 
<< m1 >>
rect 244 4 245 5 
<< m1 >>
rect 245 4 246 5 
<< m1 >>
rect 246 4 247 5 
<< m1 >>
rect 247 4 248 5 
<< m1 >>
rect 248 4 249 5 
<< m1 >>
rect 249 4 250 5 
<< m1 >>
rect 250 4 251 5 
<< m1 >>
rect 251 4 252 5 
<< m1 >>
rect 252 4 253 5 
<< m1 >>
rect 253 4 254 5 
<< m1 >>
rect 254 4 255 5 
<< m1 >>
rect 255 4 256 5 
<< m1 >>
rect 256 4 257 5 
<< m1 >>
rect 257 4 258 5 
<< m1 >>
rect 258 4 259 5 
<< m1 >>
rect 259 4 260 5 
<< m1 >>
rect 260 4 261 5 
<< m1 >>
rect 261 4 262 5 
<< m1 >>
rect 262 4 263 5 
<< m1 >>
rect 263 4 264 5 
<< m1 >>
rect 264 4 265 5 
<< m1 >>
rect 265 4 266 5 
<< m1 >>
rect 266 4 267 5 
<< m1 >>
rect 267 4 268 5 
<< m1 >>
rect 268 4 269 5 
<< m1 >>
rect 270 4 271 5 
<< m2 >>
rect 270 4 271 5 
<< m2c >>
rect 270 4 271 5 
<< m1 >>
rect 270 4 271 5 
<< m2 >>
rect 270 4 271 5 
<< m1 >>
rect 272 4 273 5 
<< m2 >>
rect 272 4 273 5 
<< m2c >>
rect 272 4 273 5 
<< m1 >>
rect 272 4 273 5 
<< m2 >>
rect 272 4 273 5 
<< m1 >>
rect 273 4 274 5 
<< m1 >>
rect 274 4 275 5 
<< m1 >>
rect 275 4 276 5 
<< m1 >>
rect 276 4 277 5 
<< m1 >>
rect 277 4 278 5 
<< m1 >>
rect 278 4 279 5 
<< m1 >>
rect 279 4 280 5 
<< m1 >>
rect 343 4 344 5 
<< m1 >>
rect 21 5 22 6 
<< m1 >>
rect 23 5 24 6 
<< m1 >>
rect 46 5 47 6 
<< m2 >>
rect 62 5 63 6 
<< m1 >>
rect 268 5 269 6 
<< m2 >>
rect 268 5 269 6 
<< m2c >>
rect 268 5 269 6 
<< m1 >>
rect 268 5 269 6 
<< m2 >>
rect 268 5 269 6 
<< m1 >>
rect 270 5 271 6 
<< m2 >>
rect 270 5 271 6 
<< m1 >>
rect 279 5 280 6 
<< m2 >>
rect 279 5 280 6 
<< m2c >>
rect 279 5 280 6 
<< m1 >>
rect 279 5 280 6 
<< m2 >>
rect 279 5 280 6 
<< m1 >>
rect 343 5 344 6 
<< m1 >>
rect 21 6 22 7 
<< m1 >>
rect 23 6 24 7 
<< m1 >>
rect 46 6 47 7 
<< m1 >>
rect 52 6 53 7 
<< m1 >>
rect 53 6 54 7 
<< m1 >>
rect 54 6 55 7 
<< m1 >>
rect 55 6 56 7 
<< m1 >>
rect 56 6 57 7 
<< m1 >>
rect 57 6 58 7 
<< m1 >>
rect 58 6 59 7 
<< m1 >>
rect 59 6 60 7 
<< m1 >>
rect 60 6 61 7 
<< m1 >>
rect 61 6 62 7 
<< m1 >>
rect 62 6 63 7 
<< m2 >>
rect 62 6 63 7 
<< m1 >>
rect 63 6 64 7 
<< m1 >>
rect 64 6 65 7 
<< m2 >>
rect 64 6 65 7 
<< m2c >>
rect 64 6 65 7 
<< m1 >>
rect 64 6 65 7 
<< m2 >>
rect 64 6 65 7 
<< m2 >>
rect 65 6 66 7 
<< m2 >>
rect 66 6 67 7 
<< m2 >>
rect 67 6 68 7 
<< m2 >>
rect 68 6 69 7 
<< m2 >>
rect 69 6 70 7 
<< m2 >>
rect 70 6 71 7 
<< m2 >>
rect 71 6 72 7 
<< m2 >>
rect 72 6 73 7 
<< m2 >>
rect 73 6 74 7 
<< m2 >>
rect 74 6 75 7 
<< m2 >>
rect 75 6 76 7 
<< m2 >>
rect 76 6 77 7 
<< m2 >>
rect 77 6 78 7 
<< m2 >>
rect 78 6 79 7 
<< m2 >>
rect 79 6 80 7 
<< m2 >>
rect 80 6 81 7 
<< m2 >>
rect 81 6 82 7 
<< m2 >>
rect 82 6 83 7 
<< m2 >>
rect 83 6 84 7 
<< m2 >>
rect 84 6 85 7 
<< m2 >>
rect 85 6 86 7 
<< m2 >>
rect 86 6 87 7 
<< m2 >>
rect 87 6 88 7 
<< m2 >>
rect 88 6 89 7 
<< m2 >>
rect 89 6 90 7 
<< m2 >>
rect 90 6 91 7 
<< m2 >>
rect 91 6 92 7 
<< m2 >>
rect 92 6 93 7 
<< m2 >>
rect 93 6 94 7 
<< m2 >>
rect 94 6 95 7 
<< m2 >>
rect 95 6 96 7 
<< m2 >>
rect 96 6 97 7 
<< m2 >>
rect 97 6 98 7 
<< m2 >>
rect 98 6 99 7 
<< m2 >>
rect 99 6 100 7 
<< m2 >>
rect 100 6 101 7 
<< m2 >>
rect 101 6 102 7 
<< m2 >>
rect 102 6 103 7 
<< m2 >>
rect 103 6 104 7 
<< m2 >>
rect 104 6 105 7 
<< m2 >>
rect 105 6 106 7 
<< m2 >>
rect 106 6 107 7 
<< m2 >>
rect 107 6 108 7 
<< m2 >>
rect 108 6 109 7 
<< m2 >>
rect 109 6 110 7 
<< m2 >>
rect 110 6 111 7 
<< m2 >>
rect 111 6 112 7 
<< m2 >>
rect 112 6 113 7 
<< m2 >>
rect 113 6 114 7 
<< m2 >>
rect 114 6 115 7 
<< m2 >>
rect 115 6 116 7 
<< m2 >>
rect 116 6 117 7 
<< m2 >>
rect 117 6 118 7 
<< m2 >>
rect 118 6 119 7 
<< m2 >>
rect 119 6 120 7 
<< m2 >>
rect 120 6 121 7 
<< m2 >>
rect 121 6 122 7 
<< m2 >>
rect 122 6 123 7 
<< m2 >>
rect 123 6 124 7 
<< m2 >>
rect 124 6 125 7 
<< m2 >>
rect 125 6 126 7 
<< m2 >>
rect 126 6 127 7 
<< m2 >>
rect 127 6 128 7 
<< m2 >>
rect 128 6 129 7 
<< m2 >>
rect 129 6 130 7 
<< m2 >>
rect 130 6 131 7 
<< m2 >>
rect 131 6 132 7 
<< m2 >>
rect 132 6 133 7 
<< m2 >>
rect 133 6 134 7 
<< m2 >>
rect 134 6 135 7 
<< m2 >>
rect 135 6 136 7 
<< m2 >>
rect 136 6 137 7 
<< m2 >>
rect 137 6 138 7 
<< m2 >>
rect 138 6 139 7 
<< m2 >>
rect 139 6 140 7 
<< m2 >>
rect 140 6 141 7 
<< m2 >>
rect 141 6 142 7 
<< m2 >>
rect 142 6 143 7 
<< m2 >>
rect 143 6 144 7 
<< m2 >>
rect 144 6 145 7 
<< m2 >>
rect 145 6 146 7 
<< m2 >>
rect 146 6 147 7 
<< m2 >>
rect 147 6 148 7 
<< m2 >>
rect 148 6 149 7 
<< m2 >>
rect 149 6 150 7 
<< m2 >>
rect 150 6 151 7 
<< m2 >>
rect 151 6 152 7 
<< m2 >>
rect 152 6 153 7 
<< m2 >>
rect 153 6 154 7 
<< m2 >>
rect 154 6 155 7 
<< m2 >>
rect 155 6 156 7 
<< m2 >>
rect 156 6 157 7 
<< m2 >>
rect 157 6 158 7 
<< m2 >>
rect 158 6 159 7 
<< m2 >>
rect 159 6 160 7 
<< m2 >>
rect 160 6 161 7 
<< m2 >>
rect 161 6 162 7 
<< m2 >>
rect 162 6 163 7 
<< m2 >>
rect 163 6 164 7 
<< m2 >>
rect 164 6 165 7 
<< m2 >>
rect 165 6 166 7 
<< m2 >>
rect 166 6 167 7 
<< m2 >>
rect 167 6 168 7 
<< m2 >>
rect 168 6 169 7 
<< m2 >>
rect 169 6 170 7 
<< m2 >>
rect 170 6 171 7 
<< m2 >>
rect 171 6 172 7 
<< m2 >>
rect 172 6 173 7 
<< m2 >>
rect 173 6 174 7 
<< m2 >>
rect 174 6 175 7 
<< m2 >>
rect 175 6 176 7 
<< m2 >>
rect 176 6 177 7 
<< m2 >>
rect 177 6 178 7 
<< m2 >>
rect 178 6 179 7 
<< m2 >>
rect 179 6 180 7 
<< m2 >>
rect 180 6 181 7 
<< m2 >>
rect 181 6 182 7 
<< m2 >>
rect 182 6 183 7 
<< m2 >>
rect 183 6 184 7 
<< m2 >>
rect 184 6 185 7 
<< m2 >>
rect 185 6 186 7 
<< m2 >>
rect 186 6 187 7 
<< m2 >>
rect 187 6 188 7 
<< m2 >>
rect 188 6 189 7 
<< m2 >>
rect 189 6 190 7 
<< m2 >>
rect 190 6 191 7 
<< m2 >>
rect 191 6 192 7 
<< m2 >>
rect 192 6 193 7 
<< m2 >>
rect 193 6 194 7 
<< m2 >>
rect 194 6 195 7 
<< m2 >>
rect 195 6 196 7 
<< m2 >>
rect 196 6 197 7 
<< m2 >>
rect 197 6 198 7 
<< m2 >>
rect 198 6 199 7 
<< m2 >>
rect 199 6 200 7 
<< m2 >>
rect 200 6 201 7 
<< m2 >>
rect 201 6 202 7 
<< m2 >>
rect 202 6 203 7 
<< m2 >>
rect 203 6 204 7 
<< m2 >>
rect 204 6 205 7 
<< m2 >>
rect 205 6 206 7 
<< m2 >>
rect 206 6 207 7 
<< m2 >>
rect 207 6 208 7 
<< m2 >>
rect 208 6 209 7 
<< m2 >>
rect 209 6 210 7 
<< m2 >>
rect 210 6 211 7 
<< m2 >>
rect 211 6 212 7 
<< m2 >>
rect 212 6 213 7 
<< m2 >>
rect 213 6 214 7 
<< m2 >>
rect 214 6 215 7 
<< m2 >>
rect 215 6 216 7 
<< m2 >>
rect 216 6 217 7 
<< m2 >>
rect 217 6 218 7 
<< m2 >>
rect 218 6 219 7 
<< m2 >>
rect 219 6 220 7 
<< m2 >>
rect 220 6 221 7 
<< m2 >>
rect 221 6 222 7 
<< m2 >>
rect 222 6 223 7 
<< m2 >>
rect 223 6 224 7 
<< m2 >>
rect 224 6 225 7 
<< m2 >>
rect 225 6 226 7 
<< m2 >>
rect 226 6 227 7 
<< m2 >>
rect 227 6 228 7 
<< m2 >>
rect 228 6 229 7 
<< m2 >>
rect 229 6 230 7 
<< m2 >>
rect 230 6 231 7 
<< m2 >>
rect 231 6 232 7 
<< m2 >>
rect 232 6 233 7 
<< m2 >>
rect 233 6 234 7 
<< m2 >>
rect 234 6 235 7 
<< m2 >>
rect 235 6 236 7 
<< m2 >>
rect 236 6 237 7 
<< m2 >>
rect 237 6 238 7 
<< m2 >>
rect 238 6 239 7 
<< m2 >>
rect 239 6 240 7 
<< m2 >>
rect 240 6 241 7 
<< m2 >>
rect 241 6 242 7 
<< m2 >>
rect 242 6 243 7 
<< m2 >>
rect 243 6 244 7 
<< m2 >>
rect 244 6 245 7 
<< m2 >>
rect 245 6 246 7 
<< m2 >>
rect 246 6 247 7 
<< m2 >>
rect 247 6 248 7 
<< m2 >>
rect 248 6 249 7 
<< m2 >>
rect 249 6 250 7 
<< m2 >>
rect 250 6 251 7 
<< m2 >>
rect 251 6 252 7 
<< m2 >>
rect 252 6 253 7 
<< m2 >>
rect 253 6 254 7 
<< m2 >>
rect 254 6 255 7 
<< m2 >>
rect 255 6 256 7 
<< m2 >>
rect 256 6 257 7 
<< m2 >>
rect 257 6 258 7 
<< m2 >>
rect 258 6 259 7 
<< m2 >>
rect 259 6 260 7 
<< m2 >>
rect 260 6 261 7 
<< m2 >>
rect 261 6 262 7 
<< m2 >>
rect 262 6 263 7 
<< m2 >>
rect 263 6 264 7 
<< m2 >>
rect 264 6 265 7 
<< m2 >>
rect 265 6 266 7 
<< m2 >>
rect 266 6 267 7 
<< m2 >>
rect 268 6 269 7 
<< m2 >>
rect 270 6 271 7 
<< m2 >>
rect 271 6 272 7 
<< m2 >>
rect 272 6 273 7 
<< m2 >>
rect 273 6 274 7 
<< m2 >>
rect 274 6 275 7 
<< m2 >>
rect 275 6 276 7 
<< m2 >>
rect 276 6 277 7 
<< m2 >>
rect 277 6 278 7 
<< m2 >>
rect 279 6 280 7 
<< m1 >>
rect 343 6 344 7 
<< m1 >>
rect 21 7 22 8 
<< m1 >>
rect 23 7 24 8 
<< m1 >>
rect 46 7 47 8 
<< m1 >>
rect 52 7 53 8 
<< m2 >>
rect 52 7 53 8 
<< m2c >>
rect 52 7 53 8 
<< m1 >>
rect 52 7 53 8 
<< m2 >>
rect 52 7 53 8 
<< m2 >>
rect 62 7 63 8 
<< m1 >>
rect 66 7 67 8 
<< m1 >>
rect 67 7 68 8 
<< m1 >>
rect 68 7 69 8 
<< m1 >>
rect 69 7 70 8 
<< m1 >>
rect 70 7 71 8 
<< m1 >>
rect 71 7 72 8 
<< m1 >>
rect 72 7 73 8 
<< m1 >>
rect 73 7 74 8 
<< m1 >>
rect 74 7 75 8 
<< m1 >>
rect 75 7 76 8 
<< m1 >>
rect 76 7 77 8 
<< m1 >>
rect 77 7 78 8 
<< m1 >>
rect 78 7 79 8 
<< m1 >>
rect 79 7 80 8 
<< m1 >>
rect 80 7 81 8 
<< m1 >>
rect 81 7 82 8 
<< m1 >>
rect 82 7 83 8 
<< m1 >>
rect 83 7 84 8 
<< m1 >>
rect 84 7 85 8 
<< m1 >>
rect 85 7 86 8 
<< m1 >>
rect 86 7 87 8 
<< m1 >>
rect 87 7 88 8 
<< m1 >>
rect 88 7 89 8 
<< m1 >>
rect 89 7 90 8 
<< m1 >>
rect 90 7 91 8 
<< m1 >>
rect 91 7 92 8 
<< m1 >>
rect 92 7 93 8 
<< m1 >>
rect 93 7 94 8 
<< m1 >>
rect 94 7 95 8 
<< m1 >>
rect 95 7 96 8 
<< m1 >>
rect 96 7 97 8 
<< m1 >>
rect 97 7 98 8 
<< m1 >>
rect 98 7 99 8 
<< m1 >>
rect 99 7 100 8 
<< m1 >>
rect 100 7 101 8 
<< m1 >>
rect 101 7 102 8 
<< m1 >>
rect 102 7 103 8 
<< m1 >>
rect 103 7 104 8 
<< m1 >>
rect 104 7 105 8 
<< m1 >>
rect 105 7 106 8 
<< m1 >>
rect 106 7 107 8 
<< m1 >>
rect 107 7 108 8 
<< m1 >>
rect 108 7 109 8 
<< m1 >>
rect 109 7 110 8 
<< m1 >>
rect 110 7 111 8 
<< m1 >>
rect 111 7 112 8 
<< m1 >>
rect 112 7 113 8 
<< m1 >>
rect 113 7 114 8 
<< m1 >>
rect 114 7 115 8 
<< m1 >>
rect 115 7 116 8 
<< m1 >>
rect 116 7 117 8 
<< m1 >>
rect 117 7 118 8 
<< m1 >>
rect 118 7 119 8 
<< m1 >>
rect 119 7 120 8 
<< m1 >>
rect 120 7 121 8 
<< m1 >>
rect 121 7 122 8 
<< m1 >>
rect 122 7 123 8 
<< m1 >>
rect 123 7 124 8 
<< m1 >>
rect 124 7 125 8 
<< m1 >>
rect 125 7 126 8 
<< m1 >>
rect 126 7 127 8 
<< m1 >>
rect 127 7 128 8 
<< m1 >>
rect 128 7 129 8 
<< m1 >>
rect 129 7 130 8 
<< m1 >>
rect 130 7 131 8 
<< m1 >>
rect 131 7 132 8 
<< m1 >>
rect 132 7 133 8 
<< m1 >>
rect 133 7 134 8 
<< m1 >>
rect 134 7 135 8 
<< m1 >>
rect 135 7 136 8 
<< m1 >>
rect 136 7 137 8 
<< m1 >>
rect 137 7 138 8 
<< m1 >>
rect 138 7 139 8 
<< m1 >>
rect 139 7 140 8 
<< m1 >>
rect 140 7 141 8 
<< m1 >>
rect 141 7 142 8 
<< m1 >>
rect 142 7 143 8 
<< m1 >>
rect 143 7 144 8 
<< m1 >>
rect 144 7 145 8 
<< m1 >>
rect 145 7 146 8 
<< m1 >>
rect 146 7 147 8 
<< m1 >>
rect 147 7 148 8 
<< m1 >>
rect 148 7 149 8 
<< m1 >>
rect 149 7 150 8 
<< m1 >>
rect 150 7 151 8 
<< m1 >>
rect 151 7 152 8 
<< m1 >>
rect 152 7 153 8 
<< m1 >>
rect 153 7 154 8 
<< m1 >>
rect 154 7 155 8 
<< m1 >>
rect 155 7 156 8 
<< m1 >>
rect 156 7 157 8 
<< m1 >>
rect 157 7 158 8 
<< m1 >>
rect 158 7 159 8 
<< m1 >>
rect 159 7 160 8 
<< m1 >>
rect 160 7 161 8 
<< m1 >>
rect 161 7 162 8 
<< m1 >>
rect 162 7 163 8 
<< m1 >>
rect 163 7 164 8 
<< m1 >>
rect 164 7 165 8 
<< m1 >>
rect 165 7 166 8 
<< m1 >>
rect 166 7 167 8 
<< m1 >>
rect 167 7 168 8 
<< m1 >>
rect 168 7 169 8 
<< m1 >>
rect 169 7 170 8 
<< m1 >>
rect 170 7 171 8 
<< m1 >>
rect 171 7 172 8 
<< m1 >>
rect 172 7 173 8 
<< m1 >>
rect 173 7 174 8 
<< m1 >>
rect 174 7 175 8 
<< m1 >>
rect 175 7 176 8 
<< m1 >>
rect 176 7 177 8 
<< m1 >>
rect 177 7 178 8 
<< m1 >>
rect 178 7 179 8 
<< m1 >>
rect 179 7 180 8 
<< m1 >>
rect 180 7 181 8 
<< m1 >>
rect 181 7 182 8 
<< m1 >>
rect 182 7 183 8 
<< m1 >>
rect 183 7 184 8 
<< m1 >>
rect 184 7 185 8 
<< m1 >>
rect 185 7 186 8 
<< m1 >>
rect 186 7 187 8 
<< m1 >>
rect 187 7 188 8 
<< m1 >>
rect 188 7 189 8 
<< m1 >>
rect 189 7 190 8 
<< m1 >>
rect 190 7 191 8 
<< m1 >>
rect 191 7 192 8 
<< m1 >>
rect 192 7 193 8 
<< m1 >>
rect 193 7 194 8 
<< m1 >>
rect 194 7 195 8 
<< m1 >>
rect 195 7 196 8 
<< m1 >>
rect 196 7 197 8 
<< m1 >>
rect 197 7 198 8 
<< m1 >>
rect 198 7 199 8 
<< m1 >>
rect 199 7 200 8 
<< m1 >>
rect 200 7 201 8 
<< m1 >>
rect 201 7 202 8 
<< m1 >>
rect 202 7 203 8 
<< m1 >>
rect 203 7 204 8 
<< m1 >>
rect 204 7 205 8 
<< m1 >>
rect 205 7 206 8 
<< m1 >>
rect 206 7 207 8 
<< m1 >>
rect 207 7 208 8 
<< m1 >>
rect 208 7 209 8 
<< m1 >>
rect 209 7 210 8 
<< m1 >>
rect 210 7 211 8 
<< m1 >>
rect 211 7 212 8 
<< m1 >>
rect 212 7 213 8 
<< m1 >>
rect 213 7 214 8 
<< m1 >>
rect 214 7 215 8 
<< m1 >>
rect 215 7 216 8 
<< m1 >>
rect 216 7 217 8 
<< m1 >>
rect 217 7 218 8 
<< m1 >>
rect 218 7 219 8 
<< m1 >>
rect 219 7 220 8 
<< m1 >>
rect 220 7 221 8 
<< m1 >>
rect 221 7 222 8 
<< m1 >>
rect 222 7 223 8 
<< m1 >>
rect 223 7 224 8 
<< m1 >>
rect 224 7 225 8 
<< m1 >>
rect 225 7 226 8 
<< m1 >>
rect 226 7 227 8 
<< m1 >>
rect 227 7 228 8 
<< m1 >>
rect 228 7 229 8 
<< m1 >>
rect 229 7 230 8 
<< m1 >>
rect 230 7 231 8 
<< m1 >>
rect 231 7 232 8 
<< m1 >>
rect 232 7 233 8 
<< m1 >>
rect 233 7 234 8 
<< m1 >>
rect 234 7 235 8 
<< m1 >>
rect 235 7 236 8 
<< m1 >>
rect 236 7 237 8 
<< m1 >>
rect 237 7 238 8 
<< m1 >>
rect 238 7 239 8 
<< m1 >>
rect 239 7 240 8 
<< m1 >>
rect 240 7 241 8 
<< m1 >>
rect 241 7 242 8 
<< m1 >>
rect 242 7 243 8 
<< m1 >>
rect 243 7 244 8 
<< m1 >>
rect 244 7 245 8 
<< m1 >>
rect 245 7 246 8 
<< m1 >>
rect 246 7 247 8 
<< m1 >>
rect 247 7 248 8 
<< m1 >>
rect 248 7 249 8 
<< m1 >>
rect 249 7 250 8 
<< m1 >>
rect 250 7 251 8 
<< m1 >>
rect 251 7 252 8 
<< m1 >>
rect 252 7 253 8 
<< m1 >>
rect 253 7 254 8 
<< m1 >>
rect 254 7 255 8 
<< m1 >>
rect 255 7 256 8 
<< m1 >>
rect 256 7 257 8 
<< m1 >>
rect 257 7 258 8 
<< m1 >>
rect 258 7 259 8 
<< m1 >>
rect 259 7 260 8 
<< m1 >>
rect 260 7 261 8 
<< m1 >>
rect 261 7 262 8 
<< m1 >>
rect 262 7 263 8 
<< m1 >>
rect 263 7 264 8 
<< m1 >>
rect 264 7 265 8 
<< m1 >>
rect 265 7 266 8 
<< m1 >>
rect 266 7 267 8 
<< m2 >>
rect 266 7 267 8 
<< m1 >>
rect 267 7 268 8 
<< m1 >>
rect 268 7 269 8 
<< m2 >>
rect 268 7 269 8 
<< m1 >>
rect 269 7 270 8 
<< m1 >>
rect 270 7 271 8 
<< m1 >>
rect 271 7 272 8 
<< m1 >>
rect 272 7 273 8 
<< m1 >>
rect 273 7 274 8 
<< m1 >>
rect 274 7 275 8 
<< m1 >>
rect 275 7 276 8 
<< m1 >>
rect 276 7 277 8 
<< m1 >>
rect 277 7 278 8 
<< m2 >>
rect 277 7 278 8 
<< m1 >>
rect 278 7 279 8 
<< m1 >>
rect 279 7 280 8 
<< m2 >>
rect 279 7 280 8 
<< m1 >>
rect 280 7 281 8 
<< m1 >>
rect 281 7 282 8 
<< m1 >>
rect 282 7 283 8 
<< m1 >>
rect 283 7 284 8 
<< m1 >>
rect 284 7 285 8 
<< m1 >>
rect 285 7 286 8 
<< m1 >>
rect 286 7 287 8 
<< m1 >>
rect 287 7 288 8 
<< m1 >>
rect 288 7 289 8 
<< m1 >>
rect 289 7 290 8 
<< m1 >>
rect 290 7 291 8 
<< m1 >>
rect 291 7 292 8 
<< m1 >>
rect 292 7 293 8 
<< m1 >>
rect 293 7 294 8 
<< m1 >>
rect 294 7 295 8 
<< m1 >>
rect 295 7 296 8 
<< m1 >>
rect 296 7 297 8 
<< m1 >>
rect 297 7 298 8 
<< m1 >>
rect 298 7 299 8 
<< m1 >>
rect 299 7 300 8 
<< m1 >>
rect 300 7 301 8 
<< m1 >>
rect 301 7 302 8 
<< m1 >>
rect 302 7 303 8 
<< m1 >>
rect 303 7 304 8 
<< m1 >>
rect 304 7 305 8 
<< m1 >>
rect 305 7 306 8 
<< m1 >>
rect 306 7 307 8 
<< m1 >>
rect 307 7 308 8 
<< m1 >>
rect 308 7 309 8 
<< m1 >>
rect 309 7 310 8 
<< m1 >>
rect 310 7 311 8 
<< m1 >>
rect 311 7 312 8 
<< m1 >>
rect 312 7 313 8 
<< m1 >>
rect 313 7 314 8 
<< m1 >>
rect 314 7 315 8 
<< m1 >>
rect 315 7 316 8 
<< m1 >>
rect 316 7 317 8 
<< m1 >>
rect 317 7 318 8 
<< m1 >>
rect 318 7 319 8 
<< m1 >>
rect 319 7 320 8 
<< m1 >>
rect 320 7 321 8 
<< m1 >>
rect 321 7 322 8 
<< m1 >>
rect 322 7 323 8 
<< m1 >>
rect 323 7 324 8 
<< m1 >>
rect 324 7 325 8 
<< m1 >>
rect 325 7 326 8 
<< m1 >>
rect 326 7 327 8 
<< m1 >>
rect 327 7 328 8 
<< m1 >>
rect 328 7 329 8 
<< m1 >>
rect 329 7 330 8 
<< m1 >>
rect 330 7 331 8 
<< m1 >>
rect 331 7 332 8 
<< m1 >>
rect 332 7 333 8 
<< m1 >>
rect 333 7 334 8 
<< m1 >>
rect 334 7 335 8 
<< m1 >>
rect 343 7 344 8 
<< m1 >>
rect 21 8 22 9 
<< m1 >>
rect 23 8 24 9 
<< m1 >>
rect 46 8 47 9 
<< m2 >>
rect 52 8 53 9 
<< m2 >>
rect 62 8 63 9 
<< m2 >>
rect 64 8 65 9 
<< m2 >>
rect 65 8 66 9 
<< m1 >>
rect 66 8 67 9 
<< m2 >>
rect 66 8 67 9 
<< m2c >>
rect 66 8 67 9 
<< m1 >>
rect 66 8 67 9 
<< m2 >>
rect 66 8 67 9 
<< m2 >>
rect 266 8 267 9 
<< m2 >>
rect 268 8 269 9 
<< m2 >>
rect 277 8 278 9 
<< m2 >>
rect 279 8 280 9 
<< m1 >>
rect 334 8 335 9 
<< m1 >>
rect 343 8 344 9 
<< m1 >>
rect 21 9 22 10 
<< m1 >>
rect 23 9 24 10 
<< m1 >>
rect 46 9 47 10 
<< m1 >>
rect 49 9 50 10 
<< m1 >>
rect 50 9 51 10 
<< m1 >>
rect 51 9 52 10 
<< m1 >>
rect 52 9 53 10 
<< m2 >>
rect 52 9 53 10 
<< m1 >>
rect 53 9 54 10 
<< m1 >>
rect 54 9 55 10 
<< m1 >>
rect 55 9 56 10 
<< m1 >>
rect 56 9 57 10 
<< m1 >>
rect 57 9 58 10 
<< m1 >>
rect 58 9 59 10 
<< m1 >>
rect 59 9 60 10 
<< m1 >>
rect 60 9 61 10 
<< m1 >>
rect 61 9 62 10 
<< m1 >>
rect 62 9 63 10 
<< m2 >>
rect 62 9 63 10 
<< m1 >>
rect 63 9 64 10 
<< m1 >>
rect 64 9 65 10 
<< m2 >>
rect 64 9 65 10 
<< m1 >>
rect 266 9 267 10 
<< m2 >>
rect 266 9 267 10 
<< m2c >>
rect 266 9 267 10 
<< m1 >>
rect 266 9 267 10 
<< m2 >>
rect 266 9 267 10 
<< m1 >>
rect 267 9 268 10 
<< m1 >>
rect 268 9 269 10 
<< m2 >>
rect 268 9 269 10 
<< m1 >>
rect 269 9 270 10 
<< m2 >>
rect 269 9 270 10 
<< m1 >>
rect 270 9 271 10 
<< m2 >>
rect 270 9 271 10 
<< m1 >>
rect 271 9 272 10 
<< m2 >>
rect 271 9 272 10 
<< m1 >>
rect 272 9 273 10 
<< m2 >>
rect 272 9 273 10 
<< m1 >>
rect 273 9 274 10 
<< m2 >>
rect 273 9 274 10 
<< m2 >>
rect 274 9 275 10 
<< m1 >>
rect 275 9 276 10 
<< m2 >>
rect 275 9 276 10 
<< m2c >>
rect 275 9 276 10 
<< m1 >>
rect 275 9 276 10 
<< m2 >>
rect 275 9 276 10 
<< m1 >>
rect 277 9 278 10 
<< m2 >>
rect 277 9 278 10 
<< m2c >>
rect 277 9 278 10 
<< m1 >>
rect 277 9 278 10 
<< m2 >>
rect 277 9 278 10 
<< m1 >>
rect 278 9 279 10 
<< m1 >>
rect 279 9 280 10 
<< m2 >>
rect 279 9 280 10 
<< m1 >>
rect 334 9 335 10 
<< m1 >>
rect 343 9 344 10 
<< m1 >>
rect 21 10 22 11 
<< m1 >>
rect 23 10 24 11 
<< m1 >>
rect 46 10 47 11 
<< m1 >>
rect 49 10 50 11 
<< m2 >>
rect 52 10 53 11 
<< m2 >>
rect 62 10 63 11 
<< m1 >>
rect 64 10 65 11 
<< m2 >>
rect 64 10 65 11 
<< m1 >>
rect 273 10 274 11 
<< m1 >>
rect 275 10 276 11 
<< m1 >>
rect 279 10 280 11 
<< m2 >>
rect 279 10 280 11 
<< m1 >>
rect 334 10 335 11 
<< m1 >>
rect 343 10 344 11 
<< m1 >>
rect 21 11 22 12 
<< m1 >>
rect 23 11 24 12 
<< m1 >>
rect 46 11 47 12 
<< m1 >>
rect 49 11 50 12 
<< m1 >>
rect 52 11 53 12 
<< m2 >>
rect 52 11 53 12 
<< m1 >>
rect 62 11 63 12 
<< m2 >>
rect 62 11 63 12 
<< m2c >>
rect 62 11 63 12 
<< m1 >>
rect 62 11 63 12 
<< m2 >>
rect 62 11 63 12 
<< m1 >>
rect 64 11 65 12 
<< m2 >>
rect 64 11 65 12 
<< m1 >>
rect 273 11 274 12 
<< m1 >>
rect 275 11 276 12 
<< m1 >>
rect 279 11 280 12 
<< m2 >>
rect 279 11 280 12 
<< m1 >>
rect 334 11 335 12 
<< m1 >>
rect 343 11 344 12 
<< pdiffusion >>
rect 12 12 13 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< m1 >>
rect 21 12 22 13 
<< m1 >>
rect 23 12 24 13 
<< pdiffusion >>
rect 30 12 31 13 
<< pdiffusion >>
rect 31 12 32 13 
<< pdiffusion >>
rect 32 12 33 13 
<< pdiffusion >>
rect 33 12 34 13 
<< pdiffusion >>
rect 34 12 35 13 
<< pdiffusion >>
rect 35 12 36 13 
<< m1 >>
rect 46 12 47 13 
<< pdiffusion >>
rect 48 12 49 13 
<< m1 >>
rect 49 12 50 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< m1 >>
rect 51 12 52 13 
<< m2 >>
rect 51 12 52 13 
<< m2c >>
rect 51 12 52 13 
<< m1 >>
rect 51 12 52 13 
<< m2 >>
rect 51 12 52 13 
<< pdiffusion >>
rect 51 12 52 13 
<< m1 >>
rect 52 12 53 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< m1 >>
rect 62 12 63 13 
<< m1 >>
rect 64 12 65 13 
<< m2 >>
rect 64 12 65 13 
<< pdiffusion >>
rect 66 12 67 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< pdiffusion >>
rect 84 12 85 13 
<< pdiffusion >>
rect 85 12 86 13 
<< pdiffusion >>
rect 86 12 87 13 
<< pdiffusion >>
rect 87 12 88 13 
<< pdiffusion >>
rect 88 12 89 13 
<< pdiffusion >>
rect 89 12 90 13 
<< pdiffusion >>
rect 102 12 103 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< pdiffusion >>
rect 120 12 121 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< pdiffusion >>
rect 138 12 139 13 
<< pdiffusion >>
rect 139 12 140 13 
<< pdiffusion >>
rect 140 12 141 13 
<< pdiffusion >>
rect 141 12 142 13 
<< pdiffusion >>
rect 142 12 143 13 
<< pdiffusion >>
rect 143 12 144 13 
<< pdiffusion >>
rect 156 12 157 13 
<< pdiffusion >>
rect 157 12 158 13 
<< pdiffusion >>
rect 158 12 159 13 
<< pdiffusion >>
rect 159 12 160 13 
<< pdiffusion >>
rect 160 12 161 13 
<< pdiffusion >>
rect 161 12 162 13 
<< pdiffusion >>
rect 174 12 175 13 
<< pdiffusion >>
rect 175 12 176 13 
<< pdiffusion >>
rect 176 12 177 13 
<< pdiffusion >>
rect 177 12 178 13 
<< pdiffusion >>
rect 178 12 179 13 
<< pdiffusion >>
rect 179 12 180 13 
<< pdiffusion >>
rect 192 12 193 13 
<< pdiffusion >>
rect 193 12 194 13 
<< pdiffusion >>
rect 194 12 195 13 
<< pdiffusion >>
rect 195 12 196 13 
<< pdiffusion >>
rect 196 12 197 13 
<< pdiffusion >>
rect 197 12 198 13 
<< pdiffusion >>
rect 210 12 211 13 
<< pdiffusion >>
rect 211 12 212 13 
<< pdiffusion >>
rect 212 12 213 13 
<< pdiffusion >>
rect 213 12 214 13 
<< pdiffusion >>
rect 214 12 215 13 
<< pdiffusion >>
rect 215 12 216 13 
<< pdiffusion >>
rect 228 12 229 13 
<< pdiffusion >>
rect 229 12 230 13 
<< pdiffusion >>
rect 230 12 231 13 
<< pdiffusion >>
rect 231 12 232 13 
<< pdiffusion >>
rect 232 12 233 13 
<< pdiffusion >>
rect 233 12 234 13 
<< pdiffusion >>
rect 246 12 247 13 
<< pdiffusion >>
rect 247 12 248 13 
<< pdiffusion >>
rect 248 12 249 13 
<< pdiffusion >>
rect 249 12 250 13 
<< pdiffusion >>
rect 250 12 251 13 
<< pdiffusion >>
rect 251 12 252 13 
<< pdiffusion >>
rect 264 12 265 13 
<< pdiffusion >>
rect 265 12 266 13 
<< pdiffusion >>
rect 266 12 267 13 
<< pdiffusion >>
rect 267 12 268 13 
<< pdiffusion >>
rect 268 12 269 13 
<< pdiffusion >>
rect 269 12 270 13 
<< m1 >>
rect 273 12 274 13 
<< m1 >>
rect 275 12 276 13 
<< m1 >>
rect 279 12 280 13 
<< m2 >>
rect 279 12 280 13 
<< pdiffusion >>
rect 282 12 283 13 
<< pdiffusion >>
rect 283 12 284 13 
<< pdiffusion >>
rect 284 12 285 13 
<< pdiffusion >>
rect 285 12 286 13 
<< pdiffusion >>
rect 286 12 287 13 
<< pdiffusion >>
rect 287 12 288 13 
<< pdiffusion >>
rect 300 12 301 13 
<< pdiffusion >>
rect 301 12 302 13 
<< pdiffusion >>
rect 302 12 303 13 
<< pdiffusion >>
rect 303 12 304 13 
<< pdiffusion >>
rect 304 12 305 13 
<< pdiffusion >>
rect 305 12 306 13 
<< pdiffusion >>
rect 318 12 319 13 
<< pdiffusion >>
rect 319 12 320 13 
<< pdiffusion >>
rect 320 12 321 13 
<< pdiffusion >>
rect 321 12 322 13 
<< pdiffusion >>
rect 322 12 323 13 
<< pdiffusion >>
rect 323 12 324 13 
<< m1 >>
rect 334 12 335 13 
<< pdiffusion >>
rect 336 12 337 13 
<< pdiffusion >>
rect 337 12 338 13 
<< pdiffusion >>
rect 338 12 339 13 
<< pdiffusion >>
rect 339 12 340 13 
<< pdiffusion >>
rect 340 12 341 13 
<< pdiffusion >>
rect 341 12 342 13 
<< m1 >>
rect 343 12 344 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< m1 >>
rect 21 13 22 14 
<< m1 >>
rect 23 13 24 14 
<< pdiffusion >>
rect 30 13 31 14 
<< pdiffusion >>
rect 31 13 32 14 
<< pdiffusion >>
rect 32 13 33 14 
<< pdiffusion >>
rect 33 13 34 14 
<< pdiffusion >>
rect 34 13 35 14 
<< pdiffusion >>
rect 35 13 36 14 
<< m1 >>
rect 46 13 47 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< m1 >>
rect 62 13 63 14 
<< m1 >>
rect 64 13 65 14 
<< m2 >>
rect 64 13 65 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< pdiffusion >>
rect 84 13 85 14 
<< pdiffusion >>
rect 85 13 86 14 
<< pdiffusion >>
rect 86 13 87 14 
<< pdiffusion >>
rect 87 13 88 14 
<< pdiffusion >>
rect 88 13 89 14 
<< pdiffusion >>
rect 89 13 90 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< pdiffusion >>
rect 138 13 139 14 
<< pdiffusion >>
rect 139 13 140 14 
<< pdiffusion >>
rect 140 13 141 14 
<< pdiffusion >>
rect 141 13 142 14 
<< pdiffusion >>
rect 142 13 143 14 
<< pdiffusion >>
rect 143 13 144 14 
<< pdiffusion >>
rect 156 13 157 14 
<< pdiffusion >>
rect 157 13 158 14 
<< pdiffusion >>
rect 158 13 159 14 
<< pdiffusion >>
rect 159 13 160 14 
<< pdiffusion >>
rect 160 13 161 14 
<< pdiffusion >>
rect 161 13 162 14 
<< pdiffusion >>
rect 174 13 175 14 
<< pdiffusion >>
rect 175 13 176 14 
<< pdiffusion >>
rect 176 13 177 14 
<< pdiffusion >>
rect 177 13 178 14 
<< pdiffusion >>
rect 178 13 179 14 
<< pdiffusion >>
rect 179 13 180 14 
<< pdiffusion >>
rect 192 13 193 14 
<< pdiffusion >>
rect 193 13 194 14 
<< pdiffusion >>
rect 194 13 195 14 
<< pdiffusion >>
rect 195 13 196 14 
<< pdiffusion >>
rect 196 13 197 14 
<< pdiffusion >>
rect 197 13 198 14 
<< pdiffusion >>
rect 210 13 211 14 
<< pdiffusion >>
rect 211 13 212 14 
<< pdiffusion >>
rect 212 13 213 14 
<< pdiffusion >>
rect 213 13 214 14 
<< pdiffusion >>
rect 214 13 215 14 
<< pdiffusion >>
rect 215 13 216 14 
<< pdiffusion >>
rect 228 13 229 14 
<< pdiffusion >>
rect 229 13 230 14 
<< pdiffusion >>
rect 230 13 231 14 
<< pdiffusion >>
rect 231 13 232 14 
<< pdiffusion >>
rect 232 13 233 14 
<< pdiffusion >>
rect 233 13 234 14 
<< pdiffusion >>
rect 246 13 247 14 
<< pdiffusion >>
rect 247 13 248 14 
<< pdiffusion >>
rect 248 13 249 14 
<< pdiffusion >>
rect 249 13 250 14 
<< pdiffusion >>
rect 250 13 251 14 
<< pdiffusion >>
rect 251 13 252 14 
<< pdiffusion >>
rect 264 13 265 14 
<< pdiffusion >>
rect 265 13 266 14 
<< pdiffusion >>
rect 266 13 267 14 
<< pdiffusion >>
rect 267 13 268 14 
<< pdiffusion >>
rect 268 13 269 14 
<< pdiffusion >>
rect 269 13 270 14 
<< m1 >>
rect 273 13 274 14 
<< m1 >>
rect 275 13 276 14 
<< m1 >>
rect 279 13 280 14 
<< m2 >>
rect 279 13 280 14 
<< pdiffusion >>
rect 282 13 283 14 
<< pdiffusion >>
rect 283 13 284 14 
<< pdiffusion >>
rect 284 13 285 14 
<< pdiffusion >>
rect 285 13 286 14 
<< pdiffusion >>
rect 286 13 287 14 
<< pdiffusion >>
rect 287 13 288 14 
<< pdiffusion >>
rect 300 13 301 14 
<< pdiffusion >>
rect 301 13 302 14 
<< pdiffusion >>
rect 302 13 303 14 
<< pdiffusion >>
rect 303 13 304 14 
<< pdiffusion >>
rect 304 13 305 14 
<< pdiffusion >>
rect 305 13 306 14 
<< pdiffusion >>
rect 318 13 319 14 
<< pdiffusion >>
rect 319 13 320 14 
<< pdiffusion >>
rect 320 13 321 14 
<< pdiffusion >>
rect 321 13 322 14 
<< pdiffusion >>
rect 322 13 323 14 
<< pdiffusion >>
rect 323 13 324 14 
<< m1 >>
rect 334 13 335 14 
<< pdiffusion >>
rect 336 13 337 14 
<< pdiffusion >>
rect 337 13 338 14 
<< pdiffusion >>
rect 338 13 339 14 
<< pdiffusion >>
rect 339 13 340 14 
<< pdiffusion >>
rect 340 13 341 14 
<< pdiffusion >>
rect 341 13 342 14 
<< m1 >>
rect 343 13 344 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< m1 >>
rect 21 14 22 15 
<< m1 >>
rect 23 14 24 15 
<< pdiffusion >>
rect 30 14 31 15 
<< pdiffusion >>
rect 31 14 32 15 
<< pdiffusion >>
rect 32 14 33 15 
<< pdiffusion >>
rect 33 14 34 15 
<< pdiffusion >>
rect 34 14 35 15 
<< pdiffusion >>
rect 35 14 36 15 
<< m1 >>
rect 46 14 47 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< m1 >>
rect 62 14 63 15 
<< m1 >>
rect 64 14 65 15 
<< m2 >>
rect 64 14 65 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< pdiffusion >>
rect 84 14 85 15 
<< pdiffusion >>
rect 85 14 86 15 
<< pdiffusion >>
rect 86 14 87 15 
<< pdiffusion >>
rect 87 14 88 15 
<< pdiffusion >>
rect 88 14 89 15 
<< pdiffusion >>
rect 89 14 90 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< pdiffusion >>
rect 138 14 139 15 
<< pdiffusion >>
rect 139 14 140 15 
<< pdiffusion >>
rect 140 14 141 15 
<< pdiffusion >>
rect 141 14 142 15 
<< pdiffusion >>
rect 142 14 143 15 
<< pdiffusion >>
rect 143 14 144 15 
<< pdiffusion >>
rect 156 14 157 15 
<< pdiffusion >>
rect 157 14 158 15 
<< pdiffusion >>
rect 158 14 159 15 
<< pdiffusion >>
rect 159 14 160 15 
<< pdiffusion >>
rect 160 14 161 15 
<< pdiffusion >>
rect 161 14 162 15 
<< pdiffusion >>
rect 174 14 175 15 
<< pdiffusion >>
rect 175 14 176 15 
<< pdiffusion >>
rect 176 14 177 15 
<< pdiffusion >>
rect 177 14 178 15 
<< pdiffusion >>
rect 178 14 179 15 
<< pdiffusion >>
rect 179 14 180 15 
<< pdiffusion >>
rect 192 14 193 15 
<< pdiffusion >>
rect 193 14 194 15 
<< pdiffusion >>
rect 194 14 195 15 
<< pdiffusion >>
rect 195 14 196 15 
<< pdiffusion >>
rect 196 14 197 15 
<< pdiffusion >>
rect 197 14 198 15 
<< pdiffusion >>
rect 210 14 211 15 
<< pdiffusion >>
rect 211 14 212 15 
<< pdiffusion >>
rect 212 14 213 15 
<< pdiffusion >>
rect 213 14 214 15 
<< pdiffusion >>
rect 214 14 215 15 
<< pdiffusion >>
rect 215 14 216 15 
<< pdiffusion >>
rect 228 14 229 15 
<< pdiffusion >>
rect 229 14 230 15 
<< pdiffusion >>
rect 230 14 231 15 
<< pdiffusion >>
rect 231 14 232 15 
<< pdiffusion >>
rect 232 14 233 15 
<< pdiffusion >>
rect 233 14 234 15 
<< pdiffusion >>
rect 246 14 247 15 
<< pdiffusion >>
rect 247 14 248 15 
<< pdiffusion >>
rect 248 14 249 15 
<< pdiffusion >>
rect 249 14 250 15 
<< pdiffusion >>
rect 250 14 251 15 
<< pdiffusion >>
rect 251 14 252 15 
<< pdiffusion >>
rect 264 14 265 15 
<< pdiffusion >>
rect 265 14 266 15 
<< pdiffusion >>
rect 266 14 267 15 
<< pdiffusion >>
rect 267 14 268 15 
<< pdiffusion >>
rect 268 14 269 15 
<< pdiffusion >>
rect 269 14 270 15 
<< m1 >>
rect 273 14 274 15 
<< m1 >>
rect 275 14 276 15 
<< m1 >>
rect 279 14 280 15 
<< m2 >>
rect 279 14 280 15 
<< pdiffusion >>
rect 282 14 283 15 
<< pdiffusion >>
rect 283 14 284 15 
<< pdiffusion >>
rect 284 14 285 15 
<< pdiffusion >>
rect 285 14 286 15 
<< pdiffusion >>
rect 286 14 287 15 
<< pdiffusion >>
rect 287 14 288 15 
<< pdiffusion >>
rect 300 14 301 15 
<< pdiffusion >>
rect 301 14 302 15 
<< pdiffusion >>
rect 302 14 303 15 
<< pdiffusion >>
rect 303 14 304 15 
<< pdiffusion >>
rect 304 14 305 15 
<< pdiffusion >>
rect 305 14 306 15 
<< pdiffusion >>
rect 318 14 319 15 
<< pdiffusion >>
rect 319 14 320 15 
<< pdiffusion >>
rect 320 14 321 15 
<< pdiffusion >>
rect 321 14 322 15 
<< pdiffusion >>
rect 322 14 323 15 
<< pdiffusion >>
rect 323 14 324 15 
<< m1 >>
rect 334 14 335 15 
<< pdiffusion >>
rect 336 14 337 15 
<< pdiffusion >>
rect 337 14 338 15 
<< pdiffusion >>
rect 338 14 339 15 
<< pdiffusion >>
rect 339 14 340 15 
<< pdiffusion >>
rect 340 14 341 15 
<< pdiffusion >>
rect 341 14 342 15 
<< m1 >>
rect 343 14 344 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< m1 >>
rect 21 15 22 16 
<< m1 >>
rect 23 15 24 16 
<< pdiffusion >>
rect 30 15 31 16 
<< pdiffusion >>
rect 31 15 32 16 
<< pdiffusion >>
rect 32 15 33 16 
<< pdiffusion >>
rect 33 15 34 16 
<< pdiffusion >>
rect 34 15 35 16 
<< pdiffusion >>
rect 35 15 36 16 
<< m1 >>
rect 46 15 47 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< m1 >>
rect 62 15 63 16 
<< m1 >>
rect 64 15 65 16 
<< m2 >>
rect 64 15 65 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< pdiffusion >>
rect 84 15 85 16 
<< pdiffusion >>
rect 85 15 86 16 
<< pdiffusion >>
rect 86 15 87 16 
<< pdiffusion >>
rect 87 15 88 16 
<< pdiffusion >>
rect 88 15 89 16 
<< pdiffusion >>
rect 89 15 90 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< pdiffusion >>
rect 138 15 139 16 
<< pdiffusion >>
rect 139 15 140 16 
<< pdiffusion >>
rect 140 15 141 16 
<< pdiffusion >>
rect 141 15 142 16 
<< pdiffusion >>
rect 142 15 143 16 
<< pdiffusion >>
rect 143 15 144 16 
<< pdiffusion >>
rect 156 15 157 16 
<< pdiffusion >>
rect 157 15 158 16 
<< pdiffusion >>
rect 158 15 159 16 
<< pdiffusion >>
rect 159 15 160 16 
<< pdiffusion >>
rect 160 15 161 16 
<< pdiffusion >>
rect 161 15 162 16 
<< pdiffusion >>
rect 174 15 175 16 
<< pdiffusion >>
rect 175 15 176 16 
<< pdiffusion >>
rect 176 15 177 16 
<< pdiffusion >>
rect 177 15 178 16 
<< pdiffusion >>
rect 178 15 179 16 
<< pdiffusion >>
rect 179 15 180 16 
<< pdiffusion >>
rect 192 15 193 16 
<< pdiffusion >>
rect 193 15 194 16 
<< pdiffusion >>
rect 194 15 195 16 
<< pdiffusion >>
rect 195 15 196 16 
<< pdiffusion >>
rect 196 15 197 16 
<< pdiffusion >>
rect 197 15 198 16 
<< pdiffusion >>
rect 210 15 211 16 
<< pdiffusion >>
rect 211 15 212 16 
<< pdiffusion >>
rect 212 15 213 16 
<< pdiffusion >>
rect 213 15 214 16 
<< pdiffusion >>
rect 214 15 215 16 
<< pdiffusion >>
rect 215 15 216 16 
<< pdiffusion >>
rect 228 15 229 16 
<< pdiffusion >>
rect 229 15 230 16 
<< pdiffusion >>
rect 230 15 231 16 
<< pdiffusion >>
rect 231 15 232 16 
<< pdiffusion >>
rect 232 15 233 16 
<< pdiffusion >>
rect 233 15 234 16 
<< pdiffusion >>
rect 246 15 247 16 
<< pdiffusion >>
rect 247 15 248 16 
<< pdiffusion >>
rect 248 15 249 16 
<< pdiffusion >>
rect 249 15 250 16 
<< pdiffusion >>
rect 250 15 251 16 
<< pdiffusion >>
rect 251 15 252 16 
<< pdiffusion >>
rect 264 15 265 16 
<< pdiffusion >>
rect 265 15 266 16 
<< pdiffusion >>
rect 266 15 267 16 
<< pdiffusion >>
rect 267 15 268 16 
<< pdiffusion >>
rect 268 15 269 16 
<< pdiffusion >>
rect 269 15 270 16 
<< m1 >>
rect 273 15 274 16 
<< m1 >>
rect 275 15 276 16 
<< m1 >>
rect 279 15 280 16 
<< m2 >>
rect 279 15 280 16 
<< pdiffusion >>
rect 282 15 283 16 
<< pdiffusion >>
rect 283 15 284 16 
<< pdiffusion >>
rect 284 15 285 16 
<< pdiffusion >>
rect 285 15 286 16 
<< pdiffusion >>
rect 286 15 287 16 
<< pdiffusion >>
rect 287 15 288 16 
<< pdiffusion >>
rect 300 15 301 16 
<< pdiffusion >>
rect 301 15 302 16 
<< pdiffusion >>
rect 302 15 303 16 
<< pdiffusion >>
rect 303 15 304 16 
<< pdiffusion >>
rect 304 15 305 16 
<< pdiffusion >>
rect 305 15 306 16 
<< pdiffusion >>
rect 318 15 319 16 
<< pdiffusion >>
rect 319 15 320 16 
<< pdiffusion >>
rect 320 15 321 16 
<< pdiffusion >>
rect 321 15 322 16 
<< pdiffusion >>
rect 322 15 323 16 
<< pdiffusion >>
rect 323 15 324 16 
<< m1 >>
rect 334 15 335 16 
<< pdiffusion >>
rect 336 15 337 16 
<< pdiffusion >>
rect 337 15 338 16 
<< pdiffusion >>
rect 338 15 339 16 
<< pdiffusion >>
rect 339 15 340 16 
<< pdiffusion >>
rect 340 15 341 16 
<< pdiffusion >>
rect 341 15 342 16 
<< m1 >>
rect 343 15 344 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< m1 >>
rect 21 16 22 17 
<< m1 >>
rect 23 16 24 17 
<< pdiffusion >>
rect 30 16 31 17 
<< pdiffusion >>
rect 31 16 32 17 
<< pdiffusion >>
rect 32 16 33 17 
<< pdiffusion >>
rect 33 16 34 17 
<< pdiffusion >>
rect 34 16 35 17 
<< pdiffusion >>
rect 35 16 36 17 
<< m1 >>
rect 46 16 47 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< m1 >>
rect 62 16 63 17 
<< m1 >>
rect 64 16 65 17 
<< m2 >>
rect 64 16 65 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< pdiffusion >>
rect 84 16 85 17 
<< pdiffusion >>
rect 85 16 86 17 
<< pdiffusion >>
rect 86 16 87 17 
<< pdiffusion >>
rect 87 16 88 17 
<< pdiffusion >>
rect 88 16 89 17 
<< pdiffusion >>
rect 89 16 90 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< pdiffusion >>
rect 138 16 139 17 
<< pdiffusion >>
rect 139 16 140 17 
<< pdiffusion >>
rect 140 16 141 17 
<< pdiffusion >>
rect 141 16 142 17 
<< pdiffusion >>
rect 142 16 143 17 
<< pdiffusion >>
rect 143 16 144 17 
<< pdiffusion >>
rect 156 16 157 17 
<< pdiffusion >>
rect 157 16 158 17 
<< pdiffusion >>
rect 158 16 159 17 
<< pdiffusion >>
rect 159 16 160 17 
<< pdiffusion >>
rect 160 16 161 17 
<< pdiffusion >>
rect 161 16 162 17 
<< pdiffusion >>
rect 174 16 175 17 
<< pdiffusion >>
rect 175 16 176 17 
<< pdiffusion >>
rect 176 16 177 17 
<< pdiffusion >>
rect 177 16 178 17 
<< pdiffusion >>
rect 178 16 179 17 
<< pdiffusion >>
rect 179 16 180 17 
<< pdiffusion >>
rect 192 16 193 17 
<< pdiffusion >>
rect 193 16 194 17 
<< pdiffusion >>
rect 194 16 195 17 
<< pdiffusion >>
rect 195 16 196 17 
<< pdiffusion >>
rect 196 16 197 17 
<< pdiffusion >>
rect 197 16 198 17 
<< pdiffusion >>
rect 210 16 211 17 
<< pdiffusion >>
rect 211 16 212 17 
<< pdiffusion >>
rect 212 16 213 17 
<< pdiffusion >>
rect 213 16 214 17 
<< pdiffusion >>
rect 214 16 215 17 
<< pdiffusion >>
rect 215 16 216 17 
<< pdiffusion >>
rect 228 16 229 17 
<< pdiffusion >>
rect 229 16 230 17 
<< pdiffusion >>
rect 230 16 231 17 
<< pdiffusion >>
rect 231 16 232 17 
<< pdiffusion >>
rect 232 16 233 17 
<< pdiffusion >>
rect 233 16 234 17 
<< pdiffusion >>
rect 246 16 247 17 
<< pdiffusion >>
rect 247 16 248 17 
<< pdiffusion >>
rect 248 16 249 17 
<< pdiffusion >>
rect 249 16 250 17 
<< pdiffusion >>
rect 250 16 251 17 
<< pdiffusion >>
rect 251 16 252 17 
<< pdiffusion >>
rect 264 16 265 17 
<< pdiffusion >>
rect 265 16 266 17 
<< pdiffusion >>
rect 266 16 267 17 
<< pdiffusion >>
rect 267 16 268 17 
<< pdiffusion >>
rect 268 16 269 17 
<< pdiffusion >>
rect 269 16 270 17 
<< m1 >>
rect 273 16 274 17 
<< m1 >>
rect 275 16 276 17 
<< m1 >>
rect 279 16 280 17 
<< m2 >>
rect 279 16 280 17 
<< pdiffusion >>
rect 282 16 283 17 
<< pdiffusion >>
rect 283 16 284 17 
<< pdiffusion >>
rect 284 16 285 17 
<< pdiffusion >>
rect 285 16 286 17 
<< pdiffusion >>
rect 286 16 287 17 
<< pdiffusion >>
rect 287 16 288 17 
<< pdiffusion >>
rect 300 16 301 17 
<< pdiffusion >>
rect 301 16 302 17 
<< pdiffusion >>
rect 302 16 303 17 
<< pdiffusion >>
rect 303 16 304 17 
<< pdiffusion >>
rect 304 16 305 17 
<< pdiffusion >>
rect 305 16 306 17 
<< pdiffusion >>
rect 318 16 319 17 
<< pdiffusion >>
rect 319 16 320 17 
<< pdiffusion >>
rect 320 16 321 17 
<< pdiffusion >>
rect 321 16 322 17 
<< pdiffusion >>
rect 322 16 323 17 
<< pdiffusion >>
rect 323 16 324 17 
<< m1 >>
rect 334 16 335 17 
<< pdiffusion >>
rect 336 16 337 17 
<< pdiffusion >>
rect 337 16 338 17 
<< pdiffusion >>
rect 338 16 339 17 
<< pdiffusion >>
rect 339 16 340 17 
<< pdiffusion >>
rect 340 16 341 17 
<< pdiffusion >>
rect 341 16 342 17 
<< m1 >>
rect 343 16 344 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< m1 >>
rect 21 17 22 18 
<< m1 >>
rect 23 17 24 18 
<< pdiffusion >>
rect 30 17 31 18 
<< pdiffusion >>
rect 31 17 32 18 
<< pdiffusion >>
rect 32 17 33 18 
<< pdiffusion >>
rect 33 17 34 18 
<< pdiffusion >>
rect 34 17 35 18 
<< pdiffusion >>
rect 35 17 36 18 
<< m1 >>
rect 46 17 47 18 
<< pdiffusion >>
rect 48 17 49 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< m1 >>
rect 62 17 63 18 
<< m1 >>
rect 64 17 65 18 
<< m2 >>
rect 64 17 65 18 
<< pdiffusion >>
rect 66 17 67 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< pdiffusion >>
rect 84 17 85 18 
<< pdiffusion >>
rect 85 17 86 18 
<< pdiffusion >>
rect 86 17 87 18 
<< pdiffusion >>
rect 87 17 88 18 
<< pdiffusion >>
rect 88 17 89 18 
<< pdiffusion >>
rect 89 17 90 18 
<< pdiffusion >>
rect 102 17 103 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< pdiffusion >>
rect 120 17 121 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< pdiffusion >>
rect 138 17 139 18 
<< pdiffusion >>
rect 139 17 140 18 
<< pdiffusion >>
rect 140 17 141 18 
<< pdiffusion >>
rect 141 17 142 18 
<< pdiffusion >>
rect 142 17 143 18 
<< pdiffusion >>
rect 143 17 144 18 
<< pdiffusion >>
rect 156 17 157 18 
<< pdiffusion >>
rect 157 17 158 18 
<< pdiffusion >>
rect 158 17 159 18 
<< pdiffusion >>
rect 159 17 160 18 
<< pdiffusion >>
rect 160 17 161 18 
<< pdiffusion >>
rect 161 17 162 18 
<< pdiffusion >>
rect 174 17 175 18 
<< pdiffusion >>
rect 175 17 176 18 
<< pdiffusion >>
rect 176 17 177 18 
<< pdiffusion >>
rect 177 17 178 18 
<< pdiffusion >>
rect 178 17 179 18 
<< pdiffusion >>
rect 179 17 180 18 
<< pdiffusion >>
rect 192 17 193 18 
<< pdiffusion >>
rect 193 17 194 18 
<< pdiffusion >>
rect 194 17 195 18 
<< pdiffusion >>
rect 195 17 196 18 
<< pdiffusion >>
rect 196 17 197 18 
<< pdiffusion >>
rect 197 17 198 18 
<< pdiffusion >>
rect 210 17 211 18 
<< pdiffusion >>
rect 211 17 212 18 
<< pdiffusion >>
rect 212 17 213 18 
<< pdiffusion >>
rect 213 17 214 18 
<< pdiffusion >>
rect 214 17 215 18 
<< pdiffusion >>
rect 215 17 216 18 
<< pdiffusion >>
rect 228 17 229 18 
<< pdiffusion >>
rect 229 17 230 18 
<< pdiffusion >>
rect 230 17 231 18 
<< pdiffusion >>
rect 231 17 232 18 
<< pdiffusion >>
rect 232 17 233 18 
<< pdiffusion >>
rect 233 17 234 18 
<< pdiffusion >>
rect 246 17 247 18 
<< pdiffusion >>
rect 247 17 248 18 
<< pdiffusion >>
rect 248 17 249 18 
<< pdiffusion >>
rect 249 17 250 18 
<< pdiffusion >>
rect 250 17 251 18 
<< pdiffusion >>
rect 251 17 252 18 
<< pdiffusion >>
rect 264 17 265 18 
<< pdiffusion >>
rect 265 17 266 18 
<< pdiffusion >>
rect 266 17 267 18 
<< pdiffusion >>
rect 267 17 268 18 
<< pdiffusion >>
rect 268 17 269 18 
<< pdiffusion >>
rect 269 17 270 18 
<< m1 >>
rect 273 17 274 18 
<< m1 >>
rect 275 17 276 18 
<< m1 >>
rect 279 17 280 18 
<< m2 >>
rect 279 17 280 18 
<< pdiffusion >>
rect 282 17 283 18 
<< pdiffusion >>
rect 283 17 284 18 
<< pdiffusion >>
rect 284 17 285 18 
<< pdiffusion >>
rect 285 17 286 18 
<< pdiffusion >>
rect 286 17 287 18 
<< pdiffusion >>
rect 287 17 288 18 
<< pdiffusion >>
rect 300 17 301 18 
<< pdiffusion >>
rect 301 17 302 18 
<< pdiffusion >>
rect 302 17 303 18 
<< pdiffusion >>
rect 303 17 304 18 
<< pdiffusion >>
rect 304 17 305 18 
<< pdiffusion >>
rect 305 17 306 18 
<< pdiffusion >>
rect 318 17 319 18 
<< pdiffusion >>
rect 319 17 320 18 
<< pdiffusion >>
rect 320 17 321 18 
<< pdiffusion >>
rect 321 17 322 18 
<< pdiffusion >>
rect 322 17 323 18 
<< pdiffusion >>
rect 323 17 324 18 
<< m1 >>
rect 334 17 335 18 
<< pdiffusion >>
rect 336 17 337 18 
<< pdiffusion >>
rect 337 17 338 18 
<< pdiffusion >>
rect 338 17 339 18 
<< pdiffusion >>
rect 339 17 340 18 
<< m1 >>
rect 340 17 341 18 
<< pdiffusion >>
rect 340 17 341 18 
<< pdiffusion >>
rect 341 17 342 18 
<< m1 >>
rect 343 17 344 18 
<< m1 >>
rect 21 18 22 19 
<< m1 >>
rect 23 18 24 19 
<< m1 >>
rect 46 18 47 19 
<< m1 >>
rect 62 18 63 19 
<< m1 >>
rect 64 18 65 19 
<< m2 >>
rect 64 18 65 19 
<< m1 >>
rect 273 18 274 19 
<< m1 >>
rect 275 18 276 19 
<< m1 >>
rect 279 18 280 19 
<< m2 >>
rect 279 18 280 19 
<< m1 >>
rect 334 18 335 19 
<< m1 >>
rect 340 18 341 19 
<< m1 >>
rect 343 18 344 19 
<< m1 >>
rect 21 19 22 20 
<< m1 >>
rect 23 19 24 20 
<< m1 >>
rect 46 19 47 20 
<< m1 >>
rect 62 19 63 20 
<< m1 >>
rect 64 19 65 20 
<< m2 >>
rect 64 19 65 20 
<< m1 >>
rect 273 19 274 20 
<< m1 >>
rect 275 19 276 20 
<< m1 >>
rect 279 19 280 20 
<< m2 >>
rect 279 19 280 20 
<< m2 >>
rect 280 19 281 20 
<< m1 >>
rect 281 19 282 20 
<< m2 >>
rect 281 19 282 20 
<< m2c >>
rect 281 19 282 20 
<< m1 >>
rect 281 19 282 20 
<< m2 >>
rect 281 19 282 20 
<< m1 >>
rect 334 19 335 20 
<< m1 >>
rect 340 19 341 20 
<< m1 >>
rect 343 19 344 20 
<< m1 >>
rect 21 20 22 21 
<< m1 >>
rect 23 20 24 21 
<< m1 >>
rect 46 20 47 21 
<< m1 >>
rect 62 20 63 21 
<< m1 >>
rect 64 20 65 21 
<< m2 >>
rect 64 20 65 21 
<< m1 >>
rect 273 20 274 21 
<< m1 >>
rect 275 20 276 21 
<< m1 >>
rect 279 20 280 21 
<< m1 >>
rect 281 20 282 21 
<< m1 >>
rect 334 20 335 21 
<< m1 >>
rect 340 20 341 21 
<< m1 >>
rect 343 20 344 21 
<< m1 >>
rect 21 21 22 22 
<< m2 >>
rect 21 21 22 22 
<< m2c >>
rect 21 21 22 22 
<< m1 >>
rect 21 21 22 22 
<< m2 >>
rect 21 21 22 22 
<< m1 >>
rect 23 21 24 22 
<< m2 >>
rect 23 21 24 22 
<< m2c >>
rect 23 21 24 22 
<< m1 >>
rect 23 21 24 22 
<< m2 >>
rect 23 21 24 22 
<< m1 >>
rect 46 21 47 22 
<< m2 >>
rect 46 21 47 22 
<< m2c >>
rect 46 21 47 22 
<< m1 >>
rect 46 21 47 22 
<< m2 >>
rect 46 21 47 22 
<< m1 >>
rect 62 21 63 22 
<< m2 >>
rect 62 21 63 22 
<< m2c >>
rect 62 21 63 22 
<< m1 >>
rect 62 21 63 22 
<< m2 >>
rect 62 21 63 22 
<< m1 >>
rect 64 21 65 22 
<< m2 >>
rect 64 21 65 22 
<< m1 >>
rect 65 21 66 22 
<< m1 >>
rect 66 21 67 22 
<< m2 >>
rect 66 21 67 22 
<< m2c >>
rect 66 21 67 22 
<< m1 >>
rect 66 21 67 22 
<< m2 >>
rect 66 21 67 22 
<< m1 >>
rect 202 21 203 22 
<< m2 >>
rect 202 21 203 22 
<< m2c >>
rect 202 21 203 22 
<< m1 >>
rect 202 21 203 22 
<< m2 >>
rect 202 21 203 22 
<< m1 >>
rect 203 21 204 22 
<< m1 >>
rect 204 21 205 22 
<< m1 >>
rect 205 21 206 22 
<< m1 >>
rect 206 21 207 22 
<< m1 >>
rect 207 21 208 22 
<< m1 >>
rect 208 21 209 22 
<< m1 >>
rect 209 21 210 22 
<< m1 >>
rect 210 21 211 22 
<< m1 >>
rect 266 21 267 22 
<< m2 >>
rect 266 21 267 22 
<< m2c >>
rect 266 21 267 22 
<< m1 >>
rect 266 21 267 22 
<< m2 >>
rect 266 21 267 22 
<< m1 >>
rect 267 21 268 22 
<< m1 >>
rect 268 21 269 22 
<< m1 >>
rect 269 21 270 22 
<< m1 >>
rect 270 21 271 22 
<< m1 >>
rect 271 21 272 22 
<< m2 >>
rect 271 21 272 22 
<< m2c >>
rect 271 21 272 22 
<< m1 >>
rect 271 21 272 22 
<< m2 >>
rect 271 21 272 22 
<< m2 >>
rect 272 21 273 22 
<< m1 >>
rect 273 21 274 22 
<< m2 >>
rect 273 21 274 22 
<< m2 >>
rect 274 21 275 22 
<< m1 >>
rect 275 21 276 22 
<< m2 >>
rect 275 21 276 22 
<< m2 >>
rect 276 21 277 22 
<< m1 >>
rect 277 21 278 22 
<< m2 >>
rect 277 21 278 22 
<< m2c >>
rect 277 21 278 22 
<< m1 >>
rect 277 21 278 22 
<< m2 >>
rect 277 21 278 22 
<< m1 >>
rect 279 21 280 22 
<< m1 >>
rect 281 21 282 22 
<< m1 >>
rect 334 21 335 22 
<< m1 >>
rect 340 21 341 22 
<< m1 >>
rect 343 21 344 22 
<< m2 >>
rect 21 22 22 23 
<< m2 >>
rect 23 22 24 23 
<< m2 >>
rect 46 22 47 23 
<< m2 >>
rect 62 22 63 23 
<< m2 >>
rect 64 22 65 23 
<< m2 >>
rect 66 22 67 23 
<< m2 >>
rect 67 22 68 23 
<< m2 >>
rect 68 22 69 23 
<< m2 >>
rect 69 22 70 23 
<< m2 >>
rect 70 22 71 23 
<< m2 >>
rect 71 22 72 23 
<< m2 >>
rect 72 22 73 23 
<< m2 >>
rect 73 22 74 23 
<< m2 >>
rect 74 22 75 23 
<< m2 >>
rect 75 22 76 23 
<< m2 >>
rect 76 22 77 23 
<< m2 >>
rect 77 22 78 23 
<< m2 >>
rect 78 22 79 23 
<< m2 >>
rect 79 22 80 23 
<< m2 >>
rect 80 22 81 23 
<< m2 >>
rect 81 22 82 23 
<< m2 >>
rect 82 22 83 23 
<< m2 >>
rect 83 22 84 23 
<< m2 >>
rect 84 22 85 23 
<< m2 >>
rect 85 22 86 23 
<< m2 >>
rect 86 22 87 23 
<< m2 >>
rect 87 22 88 23 
<< m2 >>
rect 88 22 89 23 
<< m2 >>
rect 89 22 90 23 
<< m2 >>
rect 90 22 91 23 
<< m2 >>
rect 91 22 92 23 
<< m2 >>
rect 92 22 93 23 
<< m2 >>
rect 93 22 94 23 
<< m2 >>
rect 94 22 95 23 
<< m2 >>
rect 95 22 96 23 
<< m2 >>
rect 96 22 97 23 
<< m2 >>
rect 97 22 98 23 
<< m2 >>
rect 98 22 99 23 
<< m2 >>
rect 99 22 100 23 
<< m2 >>
rect 100 22 101 23 
<< m2 >>
rect 101 22 102 23 
<< m2 >>
rect 102 22 103 23 
<< m2 >>
rect 103 22 104 23 
<< m2 >>
rect 104 22 105 23 
<< m2 >>
rect 105 22 106 23 
<< m2 >>
rect 106 22 107 23 
<< m2 >>
rect 107 22 108 23 
<< m2 >>
rect 108 22 109 23 
<< m2 >>
rect 109 22 110 23 
<< m2 >>
rect 110 22 111 23 
<< m2 >>
rect 111 22 112 23 
<< m2 >>
rect 112 22 113 23 
<< m2 >>
rect 113 22 114 23 
<< m2 >>
rect 114 22 115 23 
<< m2 >>
rect 115 22 116 23 
<< m2 >>
rect 116 22 117 23 
<< m2 >>
rect 117 22 118 23 
<< m2 >>
rect 118 22 119 23 
<< m2 >>
rect 119 22 120 23 
<< m2 >>
rect 120 22 121 23 
<< m2 >>
rect 121 22 122 23 
<< m2 >>
rect 122 22 123 23 
<< m2 >>
rect 123 22 124 23 
<< m2 >>
rect 124 22 125 23 
<< m2 >>
rect 125 22 126 23 
<< m2 >>
rect 126 22 127 23 
<< m2 >>
rect 127 22 128 23 
<< m2 >>
rect 128 22 129 23 
<< m2 >>
rect 129 22 130 23 
<< m2 >>
rect 130 22 131 23 
<< m2 >>
rect 131 22 132 23 
<< m2 >>
rect 132 22 133 23 
<< m2 >>
rect 133 22 134 23 
<< m2 >>
rect 134 22 135 23 
<< m2 >>
rect 135 22 136 23 
<< m2 >>
rect 136 22 137 23 
<< m2 >>
rect 137 22 138 23 
<< m2 >>
rect 138 22 139 23 
<< m2 >>
rect 139 22 140 23 
<< m2 >>
rect 140 22 141 23 
<< m2 >>
rect 141 22 142 23 
<< m2 >>
rect 142 22 143 23 
<< m2 >>
rect 143 22 144 23 
<< m2 >>
rect 144 22 145 23 
<< m2 >>
rect 145 22 146 23 
<< m2 >>
rect 146 22 147 23 
<< m2 >>
rect 147 22 148 23 
<< m2 >>
rect 148 22 149 23 
<< m2 >>
rect 149 22 150 23 
<< m2 >>
rect 150 22 151 23 
<< m2 >>
rect 151 22 152 23 
<< m2 >>
rect 152 22 153 23 
<< m2 >>
rect 153 22 154 23 
<< m2 >>
rect 154 22 155 23 
<< m2 >>
rect 155 22 156 23 
<< m2 >>
rect 156 22 157 23 
<< m2 >>
rect 157 22 158 23 
<< m2 >>
rect 158 22 159 23 
<< m2 >>
rect 159 22 160 23 
<< m2 >>
rect 160 22 161 23 
<< m2 >>
rect 161 22 162 23 
<< m2 >>
rect 162 22 163 23 
<< m2 >>
rect 163 22 164 23 
<< m2 >>
rect 164 22 165 23 
<< m2 >>
rect 165 22 166 23 
<< m2 >>
rect 166 22 167 23 
<< m2 >>
rect 167 22 168 23 
<< m2 >>
rect 168 22 169 23 
<< m2 >>
rect 169 22 170 23 
<< m2 >>
rect 170 22 171 23 
<< m2 >>
rect 171 22 172 23 
<< m2 >>
rect 172 22 173 23 
<< m2 >>
rect 173 22 174 23 
<< m2 >>
rect 174 22 175 23 
<< m2 >>
rect 175 22 176 23 
<< m2 >>
rect 176 22 177 23 
<< m2 >>
rect 177 22 178 23 
<< m2 >>
rect 178 22 179 23 
<< m2 >>
rect 179 22 180 23 
<< m2 >>
rect 180 22 181 23 
<< m2 >>
rect 181 22 182 23 
<< m2 >>
rect 182 22 183 23 
<< m2 >>
rect 183 22 184 23 
<< m2 >>
rect 184 22 185 23 
<< m2 >>
rect 185 22 186 23 
<< m2 >>
rect 186 22 187 23 
<< m2 >>
rect 187 22 188 23 
<< m2 >>
rect 188 22 189 23 
<< m2 >>
rect 189 22 190 23 
<< m2 >>
rect 190 22 191 23 
<< m2 >>
rect 191 22 192 23 
<< m2 >>
rect 192 22 193 23 
<< m2 >>
rect 193 22 194 23 
<< m2 >>
rect 194 22 195 23 
<< m2 >>
rect 195 22 196 23 
<< m2 >>
rect 196 22 197 23 
<< m2 >>
rect 197 22 198 23 
<< m2 >>
rect 198 22 199 23 
<< m2 >>
rect 199 22 200 23 
<< m2 >>
rect 200 22 201 23 
<< m2 >>
rect 201 22 202 23 
<< m2 >>
rect 202 22 203 23 
<< m1 >>
rect 210 22 211 23 
<< m2 >>
rect 266 22 267 23 
<< m1 >>
rect 273 22 274 23 
<< m1 >>
rect 275 22 276 23 
<< m1 >>
rect 277 22 278 23 
<< m1 >>
rect 279 22 280 23 
<< m1 >>
rect 281 22 282 23 
<< m1 >>
rect 334 22 335 23 
<< m1 >>
rect 340 22 341 23 
<< m1 >>
rect 343 22 344 23 
<< m1 >>
rect 19 23 20 24 
<< m1 >>
rect 20 23 21 24 
<< m1 >>
rect 21 23 22 24 
<< m2 >>
rect 21 23 22 24 
<< m1 >>
rect 22 23 23 24 
<< m1 >>
rect 23 23 24 24 
<< m2 >>
rect 23 23 24 24 
<< m1 >>
rect 24 23 25 24 
<< m1 >>
rect 25 23 26 24 
<< m1 >>
rect 26 23 27 24 
<< m1 >>
rect 27 23 28 24 
<< m1 >>
rect 28 23 29 24 
<< m1 >>
rect 29 23 30 24 
<< m1 >>
rect 30 23 31 24 
<< m1 >>
rect 31 23 32 24 
<< m1 >>
rect 32 23 33 24 
<< m1 >>
rect 33 23 34 24 
<< m1 >>
rect 34 23 35 24 
<< m1 >>
rect 35 23 36 24 
<< m1 >>
rect 36 23 37 24 
<< m1 >>
rect 37 23 38 24 
<< m1 >>
rect 38 23 39 24 
<< m1 >>
rect 39 23 40 24 
<< m1 >>
rect 40 23 41 24 
<< m1 >>
rect 41 23 42 24 
<< m1 >>
rect 42 23 43 24 
<< m1 >>
rect 43 23 44 24 
<< m1 >>
rect 44 23 45 24 
<< m1 >>
rect 45 23 46 24 
<< m1 >>
rect 46 23 47 24 
<< m2 >>
rect 46 23 47 24 
<< m1 >>
rect 47 23 48 24 
<< m1 >>
rect 48 23 49 24 
<< m1 >>
rect 49 23 50 24 
<< m1 >>
rect 50 23 51 24 
<< m1 >>
rect 51 23 52 24 
<< m1 >>
rect 52 23 53 24 
<< m1 >>
rect 53 23 54 24 
<< m1 >>
rect 54 23 55 24 
<< m1 >>
rect 55 23 56 24 
<< m1 >>
rect 56 23 57 24 
<< m1 >>
rect 57 23 58 24 
<< m1 >>
rect 58 23 59 24 
<< m1 >>
rect 59 23 60 24 
<< m1 >>
rect 60 23 61 24 
<< m1 >>
rect 61 23 62 24 
<< m1 >>
rect 62 23 63 24 
<< m2 >>
rect 62 23 63 24 
<< m1 >>
rect 63 23 64 24 
<< m1 >>
rect 64 23 65 24 
<< m2 >>
rect 64 23 65 24 
<< m1 >>
rect 65 23 66 24 
<< m1 >>
rect 66 23 67 24 
<< m1 >>
rect 67 23 68 24 
<< m1 >>
rect 68 23 69 24 
<< m1 >>
rect 69 23 70 24 
<< m1 >>
rect 70 23 71 24 
<< m1 >>
rect 71 23 72 24 
<< m1 >>
rect 72 23 73 24 
<< m1 >>
rect 73 23 74 24 
<< m1 >>
rect 74 23 75 24 
<< m1 >>
rect 75 23 76 24 
<< m1 >>
rect 76 23 77 24 
<< m1 >>
rect 77 23 78 24 
<< m1 >>
rect 78 23 79 24 
<< m1 >>
rect 79 23 80 24 
<< m1 >>
rect 80 23 81 24 
<< m1 >>
rect 81 23 82 24 
<< m1 >>
rect 82 23 83 24 
<< m1 >>
rect 83 23 84 24 
<< m1 >>
rect 84 23 85 24 
<< m1 >>
rect 85 23 86 24 
<< m1 >>
rect 86 23 87 24 
<< m1 >>
rect 87 23 88 24 
<< m1 >>
rect 88 23 89 24 
<< m1 >>
rect 89 23 90 24 
<< m1 >>
rect 90 23 91 24 
<< m1 >>
rect 91 23 92 24 
<< m1 >>
rect 92 23 93 24 
<< m1 >>
rect 93 23 94 24 
<< m1 >>
rect 94 23 95 24 
<< m1 >>
rect 95 23 96 24 
<< m1 >>
rect 96 23 97 24 
<< m1 >>
rect 97 23 98 24 
<< m1 >>
rect 98 23 99 24 
<< m1 >>
rect 99 23 100 24 
<< m1 >>
rect 100 23 101 24 
<< m1 >>
rect 101 23 102 24 
<< m1 >>
rect 102 23 103 24 
<< m1 >>
rect 103 23 104 24 
<< m1 >>
rect 104 23 105 24 
<< m1 >>
rect 105 23 106 24 
<< m1 >>
rect 106 23 107 24 
<< m1 >>
rect 107 23 108 24 
<< m1 >>
rect 108 23 109 24 
<< m1 >>
rect 109 23 110 24 
<< m1 >>
rect 110 23 111 24 
<< m1 >>
rect 111 23 112 24 
<< m1 >>
rect 112 23 113 24 
<< m1 >>
rect 113 23 114 24 
<< m1 >>
rect 114 23 115 24 
<< m1 >>
rect 115 23 116 24 
<< m1 >>
rect 116 23 117 24 
<< m1 >>
rect 117 23 118 24 
<< m1 >>
rect 118 23 119 24 
<< m1 >>
rect 119 23 120 24 
<< m1 >>
rect 120 23 121 24 
<< m1 >>
rect 121 23 122 24 
<< m1 >>
rect 122 23 123 24 
<< m1 >>
rect 123 23 124 24 
<< m1 >>
rect 124 23 125 24 
<< m1 >>
rect 125 23 126 24 
<< m1 >>
rect 126 23 127 24 
<< m1 >>
rect 127 23 128 24 
<< m1 >>
rect 128 23 129 24 
<< m1 >>
rect 129 23 130 24 
<< m1 >>
rect 130 23 131 24 
<< m1 >>
rect 131 23 132 24 
<< m1 >>
rect 132 23 133 24 
<< m1 >>
rect 133 23 134 24 
<< m1 >>
rect 134 23 135 24 
<< m1 >>
rect 135 23 136 24 
<< m1 >>
rect 136 23 137 24 
<< m1 >>
rect 137 23 138 24 
<< m1 >>
rect 138 23 139 24 
<< m1 >>
rect 139 23 140 24 
<< m1 >>
rect 140 23 141 24 
<< m1 >>
rect 141 23 142 24 
<< m1 >>
rect 142 23 143 24 
<< m1 >>
rect 143 23 144 24 
<< m1 >>
rect 144 23 145 24 
<< m1 >>
rect 145 23 146 24 
<< m1 >>
rect 146 23 147 24 
<< m1 >>
rect 147 23 148 24 
<< m1 >>
rect 148 23 149 24 
<< m1 >>
rect 149 23 150 24 
<< m1 >>
rect 150 23 151 24 
<< m1 >>
rect 151 23 152 24 
<< m1 >>
rect 152 23 153 24 
<< m1 >>
rect 153 23 154 24 
<< m1 >>
rect 154 23 155 24 
<< m1 >>
rect 155 23 156 24 
<< m1 >>
rect 156 23 157 24 
<< m1 >>
rect 157 23 158 24 
<< m1 >>
rect 158 23 159 24 
<< m1 >>
rect 159 23 160 24 
<< m1 >>
rect 160 23 161 24 
<< m1 >>
rect 161 23 162 24 
<< m1 >>
rect 162 23 163 24 
<< m1 >>
rect 163 23 164 24 
<< m1 >>
rect 164 23 165 24 
<< m1 >>
rect 165 23 166 24 
<< m1 >>
rect 166 23 167 24 
<< m1 >>
rect 167 23 168 24 
<< m1 >>
rect 168 23 169 24 
<< m1 >>
rect 169 23 170 24 
<< m1 >>
rect 170 23 171 24 
<< m1 >>
rect 171 23 172 24 
<< m1 >>
rect 172 23 173 24 
<< m1 >>
rect 173 23 174 24 
<< m1 >>
rect 174 23 175 24 
<< m1 >>
rect 175 23 176 24 
<< m1 >>
rect 176 23 177 24 
<< m1 >>
rect 177 23 178 24 
<< m1 >>
rect 178 23 179 24 
<< m1 >>
rect 179 23 180 24 
<< m1 >>
rect 180 23 181 24 
<< m1 >>
rect 181 23 182 24 
<< m1 >>
rect 182 23 183 24 
<< m1 >>
rect 183 23 184 24 
<< m1 >>
rect 184 23 185 24 
<< m1 >>
rect 185 23 186 24 
<< m1 >>
rect 186 23 187 24 
<< m1 >>
rect 187 23 188 24 
<< m1 >>
rect 188 23 189 24 
<< m1 >>
rect 189 23 190 24 
<< m1 >>
rect 190 23 191 24 
<< m1 >>
rect 191 23 192 24 
<< m1 >>
rect 192 23 193 24 
<< m1 >>
rect 193 23 194 24 
<< m1 >>
rect 194 23 195 24 
<< m1 >>
rect 195 23 196 24 
<< m1 >>
rect 196 23 197 24 
<< m1 >>
rect 197 23 198 24 
<< m1 >>
rect 198 23 199 24 
<< m1 >>
rect 199 23 200 24 
<< m1 >>
rect 200 23 201 24 
<< m1 >>
rect 201 23 202 24 
<< m1 >>
rect 202 23 203 24 
<< m1 >>
rect 203 23 204 24 
<< m1 >>
rect 204 23 205 24 
<< m2 >>
rect 204 23 205 24 
<< m2c >>
rect 204 23 205 24 
<< m1 >>
rect 204 23 205 24 
<< m2 >>
rect 204 23 205 24 
<< m1 >>
rect 210 23 211 24 
<< m1 >>
rect 211 23 212 24 
<< m1 >>
rect 212 23 213 24 
<< m1 >>
rect 213 23 214 24 
<< m1 >>
rect 214 23 215 24 
<< m1 >>
rect 215 23 216 24 
<< m1 >>
rect 216 23 217 24 
<< m1 >>
rect 217 23 218 24 
<< m1 >>
rect 218 23 219 24 
<< m1 >>
rect 219 23 220 24 
<< m1 >>
rect 220 23 221 24 
<< m1 >>
rect 221 23 222 24 
<< m1 >>
rect 222 23 223 24 
<< m1 >>
rect 223 23 224 24 
<< m1 >>
rect 224 23 225 24 
<< m1 >>
rect 225 23 226 24 
<< m1 >>
rect 226 23 227 24 
<< m1 >>
rect 227 23 228 24 
<< m1 >>
rect 228 23 229 24 
<< m1 >>
rect 229 23 230 24 
<< m1 >>
rect 230 23 231 24 
<< m1 >>
rect 231 23 232 24 
<< m1 >>
rect 232 23 233 24 
<< m1 >>
rect 233 23 234 24 
<< m1 >>
rect 234 23 235 24 
<< m1 >>
rect 235 23 236 24 
<< m1 >>
rect 236 23 237 24 
<< m1 >>
rect 237 23 238 24 
<< m1 >>
rect 238 23 239 24 
<< m1 >>
rect 239 23 240 24 
<< m1 >>
rect 240 23 241 24 
<< m1 >>
rect 241 23 242 24 
<< m1 >>
rect 242 23 243 24 
<< m1 >>
rect 243 23 244 24 
<< m1 >>
rect 244 23 245 24 
<< m1 >>
rect 245 23 246 24 
<< m1 >>
rect 246 23 247 24 
<< m1 >>
rect 247 23 248 24 
<< m1 >>
rect 248 23 249 24 
<< m1 >>
rect 249 23 250 24 
<< m1 >>
rect 250 23 251 24 
<< m1 >>
rect 251 23 252 24 
<< m1 >>
rect 252 23 253 24 
<< m1 >>
rect 253 23 254 24 
<< m1 >>
rect 254 23 255 24 
<< m1 >>
rect 255 23 256 24 
<< m1 >>
rect 256 23 257 24 
<< m1 >>
rect 257 23 258 24 
<< m1 >>
rect 258 23 259 24 
<< m1 >>
rect 259 23 260 24 
<< m1 >>
rect 260 23 261 24 
<< m1 >>
rect 261 23 262 24 
<< m1 >>
rect 262 23 263 24 
<< m1 >>
rect 263 23 264 24 
<< m1 >>
rect 264 23 265 24 
<< m1 >>
rect 265 23 266 24 
<< m1 >>
rect 266 23 267 24 
<< m2 >>
rect 266 23 267 24 
<< m1 >>
rect 267 23 268 24 
<< m1 >>
rect 268 23 269 24 
<< m1 >>
rect 269 23 270 24 
<< m1 >>
rect 270 23 271 24 
<< m1 >>
rect 271 23 272 24 
<< m2 >>
rect 271 23 272 24 
<< m2c >>
rect 271 23 272 24 
<< m1 >>
rect 271 23 272 24 
<< m2 >>
rect 271 23 272 24 
<< m1 >>
rect 273 23 274 24 
<< m2 >>
rect 273 23 274 24 
<< m2c >>
rect 273 23 274 24 
<< m1 >>
rect 273 23 274 24 
<< m2 >>
rect 273 23 274 24 
<< m1 >>
rect 275 23 276 24 
<< m2 >>
rect 275 23 276 24 
<< m2c >>
rect 275 23 276 24 
<< m1 >>
rect 275 23 276 24 
<< m2 >>
rect 275 23 276 24 
<< m1 >>
rect 277 23 278 24 
<< m2 >>
rect 277 23 278 24 
<< m2c >>
rect 277 23 278 24 
<< m1 >>
rect 277 23 278 24 
<< m2 >>
rect 277 23 278 24 
<< m1 >>
rect 279 23 280 24 
<< m2 >>
rect 279 23 280 24 
<< m2c >>
rect 279 23 280 24 
<< m1 >>
rect 279 23 280 24 
<< m2 >>
rect 279 23 280 24 
<< m1 >>
rect 281 23 282 24 
<< m2 >>
rect 281 23 282 24 
<< m2c >>
rect 281 23 282 24 
<< m1 >>
rect 281 23 282 24 
<< m2 >>
rect 281 23 282 24 
<< m1 >>
rect 334 23 335 24 
<< m2 >>
rect 334 23 335 24 
<< m2c >>
rect 334 23 335 24 
<< m1 >>
rect 334 23 335 24 
<< m2 >>
rect 334 23 335 24 
<< m1 >>
rect 340 23 341 24 
<< m1 >>
rect 343 23 344 24 
<< m1 >>
rect 19 24 20 25 
<< m2 >>
rect 21 24 22 25 
<< m2 >>
rect 23 24 24 25 
<< m2 >>
rect 46 24 47 25 
<< m2 >>
rect 62 24 63 25 
<< m2 >>
rect 64 24 65 25 
<< m2 >>
rect 204 24 205 25 
<< m2 >>
rect 205 24 206 25 
<< m2 >>
rect 206 24 207 25 
<< m2 >>
rect 207 24 208 25 
<< m2 >>
rect 208 24 209 25 
<< m2 >>
rect 209 24 210 25 
<< m2 >>
rect 210 24 211 25 
<< m2 >>
rect 211 24 212 25 
<< m2 >>
rect 212 24 213 25 
<< m2 >>
rect 213 24 214 25 
<< m2 >>
rect 214 24 215 25 
<< m2 >>
rect 215 24 216 25 
<< m2 >>
rect 216 24 217 25 
<< m2 >>
rect 217 24 218 25 
<< m2 >>
rect 218 24 219 25 
<< m2 >>
rect 219 24 220 25 
<< m2 >>
rect 220 24 221 25 
<< m2 >>
rect 221 24 222 25 
<< m2 >>
rect 222 24 223 25 
<< m2 >>
rect 223 24 224 25 
<< m2 >>
rect 224 24 225 25 
<< m2 >>
rect 225 24 226 25 
<< m2 >>
rect 266 24 267 25 
<< m2 >>
rect 271 24 272 25 
<< m2 >>
rect 273 24 274 25 
<< m2 >>
rect 275 24 276 25 
<< m2 >>
rect 277 24 278 25 
<< m2 >>
rect 279 24 280 25 
<< m2 >>
rect 281 24 282 25 
<< m2 >>
rect 282 24 283 25 
<< m2 >>
rect 283 24 284 25 
<< m2 >>
rect 284 24 285 25 
<< m2 >>
rect 334 24 335 25 
<< m1 >>
rect 340 24 341 25 
<< m1 >>
rect 343 24 344 25 
<< m1 >>
rect 19 25 20 26 
<< m1 >>
rect 21 25 22 26 
<< m2 >>
rect 21 25 22 26 
<< m2c >>
rect 21 25 22 26 
<< m1 >>
rect 21 25 22 26 
<< m2 >>
rect 21 25 22 26 
<< m1 >>
rect 23 25 24 26 
<< m2 >>
rect 23 25 24 26 
<< m2c >>
rect 23 25 24 26 
<< m1 >>
rect 23 25 24 26 
<< m2 >>
rect 23 25 24 26 
<< m1 >>
rect 46 25 47 26 
<< m2 >>
rect 46 25 47 26 
<< m2c >>
rect 46 25 47 26 
<< m1 >>
rect 46 25 47 26 
<< m2 >>
rect 46 25 47 26 
<< m1 >>
rect 62 25 63 26 
<< m2 >>
rect 62 25 63 26 
<< m2c >>
rect 62 25 63 26 
<< m1 >>
rect 62 25 63 26 
<< m2 >>
rect 62 25 63 26 
<< m1 >>
rect 64 25 65 26 
<< m2 >>
rect 64 25 65 26 
<< m2c >>
rect 64 25 65 26 
<< m1 >>
rect 64 25 65 26 
<< m2 >>
rect 64 25 65 26 
<< m1 >>
rect 78 25 79 26 
<< m1 >>
rect 79 25 80 26 
<< m1 >>
rect 80 25 81 26 
<< m2 >>
rect 80 25 81 26 
<< m2c >>
rect 80 25 81 26 
<< m1 >>
rect 80 25 81 26 
<< m2 >>
rect 80 25 81 26 
<< m2 >>
rect 81 25 82 26 
<< m1 >>
rect 82 25 83 26 
<< m2 >>
rect 82 25 83 26 
<< m1 >>
rect 83 25 84 26 
<< m2 >>
rect 83 25 84 26 
<< m1 >>
rect 84 25 85 26 
<< m2 >>
rect 84 25 85 26 
<< m1 >>
rect 85 25 86 26 
<< m2 >>
rect 85 25 86 26 
<< m1 >>
rect 86 25 87 26 
<< m2 >>
rect 86 25 87 26 
<< m1 >>
rect 87 25 88 26 
<< m2 >>
rect 87 25 88 26 
<< m1 >>
rect 88 25 89 26 
<< m2 >>
rect 88 25 89 26 
<< m2 >>
rect 89 25 90 26 
<< m1 >>
rect 90 25 91 26 
<< m2 >>
rect 90 25 91 26 
<< m2c >>
rect 90 25 91 26 
<< m1 >>
rect 90 25 91 26 
<< m2 >>
rect 90 25 91 26 
<< m1 >>
rect 91 25 92 26 
<< m1 >>
rect 92 25 93 26 
<< m2 >>
rect 92 25 93 26 
<< m1 >>
rect 93 25 94 26 
<< m2 >>
rect 93 25 94 26 
<< m1 >>
rect 94 25 95 26 
<< m2 >>
rect 94 25 95 26 
<< m1 >>
rect 95 25 96 26 
<< m2 >>
rect 95 25 96 26 
<< m1 >>
rect 96 25 97 26 
<< m2 >>
rect 96 25 97 26 
<< m1 >>
rect 97 25 98 26 
<< m2 >>
rect 97 25 98 26 
<< m1 >>
rect 98 25 99 26 
<< m2 >>
rect 98 25 99 26 
<< m1 >>
rect 99 25 100 26 
<< m2 >>
rect 99 25 100 26 
<< m1 >>
rect 100 25 101 26 
<< m2 >>
rect 100 25 101 26 
<< m1 >>
rect 101 25 102 26 
<< m2 >>
rect 101 25 102 26 
<< m1 >>
rect 102 25 103 26 
<< m2 >>
rect 102 25 103 26 
<< m1 >>
rect 103 25 104 26 
<< m2 >>
rect 103 25 104 26 
<< m1 >>
rect 104 25 105 26 
<< m2 >>
rect 104 25 105 26 
<< m1 >>
rect 105 25 106 26 
<< m2 >>
rect 105 25 106 26 
<< m1 >>
rect 106 25 107 26 
<< m2 >>
rect 106 25 107 26 
<< m1 >>
rect 107 25 108 26 
<< m2 >>
rect 107 25 108 26 
<< m1 >>
rect 108 25 109 26 
<< m2 >>
rect 108 25 109 26 
<< m1 >>
rect 109 25 110 26 
<< m2 >>
rect 109 25 110 26 
<< m1 >>
rect 110 25 111 26 
<< m2 >>
rect 110 25 111 26 
<< m1 >>
rect 111 25 112 26 
<< m2 >>
rect 111 25 112 26 
<< m1 >>
rect 112 25 113 26 
<< m2 >>
rect 112 25 113 26 
<< m1 >>
rect 113 25 114 26 
<< m2 >>
rect 113 25 114 26 
<< m1 >>
rect 114 25 115 26 
<< m2 >>
rect 114 25 115 26 
<< m1 >>
rect 115 25 116 26 
<< m2 >>
rect 115 25 116 26 
<< m1 >>
rect 116 25 117 26 
<< m2 >>
rect 116 25 117 26 
<< m1 >>
rect 117 25 118 26 
<< m2 >>
rect 117 25 118 26 
<< m1 >>
rect 118 25 119 26 
<< m2 >>
rect 118 25 119 26 
<< m1 >>
rect 119 25 120 26 
<< m2 >>
rect 119 25 120 26 
<< m1 >>
rect 120 25 121 26 
<< m2 >>
rect 120 25 121 26 
<< m1 >>
rect 121 25 122 26 
<< m2 >>
rect 121 25 122 26 
<< m1 >>
rect 122 25 123 26 
<< m2 >>
rect 122 25 123 26 
<< m1 >>
rect 123 25 124 26 
<< m2 >>
rect 123 25 124 26 
<< m1 >>
rect 124 25 125 26 
<< m2 >>
rect 124 25 125 26 
<< m1 >>
rect 125 25 126 26 
<< m2 >>
rect 125 25 126 26 
<< m1 >>
rect 126 25 127 26 
<< m2 >>
rect 126 25 127 26 
<< m1 >>
rect 127 25 128 26 
<< m2 >>
rect 127 25 128 26 
<< m1 >>
rect 128 25 129 26 
<< m2 >>
rect 128 25 129 26 
<< m1 >>
rect 129 25 130 26 
<< m2 >>
rect 129 25 130 26 
<< m1 >>
rect 130 25 131 26 
<< m2 >>
rect 130 25 131 26 
<< m1 >>
rect 131 25 132 26 
<< m2 >>
rect 131 25 132 26 
<< m1 >>
rect 132 25 133 26 
<< m2 >>
rect 132 25 133 26 
<< m1 >>
rect 133 25 134 26 
<< m2 >>
rect 133 25 134 26 
<< m1 >>
rect 134 25 135 26 
<< m2 >>
rect 134 25 135 26 
<< m1 >>
rect 135 25 136 26 
<< m2 >>
rect 135 25 136 26 
<< m1 >>
rect 136 25 137 26 
<< m2 >>
rect 136 25 137 26 
<< m1 >>
rect 137 25 138 26 
<< m2 >>
rect 137 25 138 26 
<< m1 >>
rect 138 25 139 26 
<< m2 >>
rect 138 25 139 26 
<< m1 >>
rect 139 25 140 26 
<< m2 >>
rect 139 25 140 26 
<< m1 >>
rect 140 25 141 26 
<< m2 >>
rect 140 25 141 26 
<< m1 >>
rect 141 25 142 26 
<< m2 >>
rect 141 25 142 26 
<< m1 >>
rect 142 25 143 26 
<< m2 >>
rect 142 25 143 26 
<< m1 >>
rect 143 25 144 26 
<< m2 >>
rect 143 25 144 26 
<< m1 >>
rect 144 25 145 26 
<< m2 >>
rect 144 25 145 26 
<< m1 >>
rect 145 25 146 26 
<< m2 >>
rect 145 25 146 26 
<< m1 >>
rect 146 25 147 26 
<< m2 >>
rect 146 25 147 26 
<< m1 >>
rect 147 25 148 26 
<< m2 >>
rect 147 25 148 26 
<< m1 >>
rect 148 25 149 26 
<< m2 >>
rect 148 25 149 26 
<< m1 >>
rect 149 25 150 26 
<< m2 >>
rect 149 25 150 26 
<< m1 >>
rect 150 25 151 26 
<< m2 >>
rect 150 25 151 26 
<< m1 >>
rect 151 25 152 26 
<< m2 >>
rect 151 25 152 26 
<< m1 >>
rect 152 25 153 26 
<< m2 >>
rect 152 25 153 26 
<< m1 >>
rect 153 25 154 26 
<< m2 >>
rect 153 25 154 26 
<< m1 >>
rect 154 25 155 26 
<< m2 >>
rect 154 25 155 26 
<< m1 >>
rect 155 25 156 26 
<< m2 >>
rect 155 25 156 26 
<< m1 >>
rect 156 25 157 26 
<< m2 >>
rect 156 25 157 26 
<< m1 >>
rect 157 25 158 26 
<< m2 >>
rect 157 25 158 26 
<< m1 >>
rect 158 25 159 26 
<< m2 >>
rect 158 25 159 26 
<< m1 >>
rect 159 25 160 26 
<< m2 >>
rect 159 25 160 26 
<< m1 >>
rect 160 25 161 26 
<< m2 >>
rect 160 25 161 26 
<< m1 >>
rect 161 25 162 26 
<< m2 >>
rect 161 25 162 26 
<< m1 >>
rect 162 25 163 26 
<< m2 >>
rect 162 25 163 26 
<< m1 >>
rect 163 25 164 26 
<< m2 >>
rect 163 25 164 26 
<< m1 >>
rect 164 25 165 26 
<< m2 >>
rect 164 25 165 26 
<< m1 >>
rect 165 25 166 26 
<< m2 >>
rect 165 25 166 26 
<< m1 >>
rect 166 25 167 26 
<< m2 >>
rect 166 25 167 26 
<< m1 >>
rect 167 25 168 26 
<< m2 >>
rect 167 25 168 26 
<< m1 >>
rect 168 25 169 26 
<< m2 >>
rect 168 25 169 26 
<< m1 >>
rect 169 25 170 26 
<< m2 >>
rect 169 25 170 26 
<< m1 >>
rect 170 25 171 26 
<< m2 >>
rect 170 25 171 26 
<< m1 >>
rect 171 25 172 26 
<< m2 >>
rect 171 25 172 26 
<< m1 >>
rect 172 25 173 26 
<< m2 >>
rect 172 25 173 26 
<< m1 >>
rect 173 25 174 26 
<< m2 >>
rect 173 25 174 26 
<< m1 >>
rect 174 25 175 26 
<< m2 >>
rect 174 25 175 26 
<< m1 >>
rect 175 25 176 26 
<< m2 >>
rect 175 25 176 26 
<< m1 >>
rect 176 25 177 26 
<< m2 >>
rect 176 25 177 26 
<< m1 >>
rect 177 25 178 26 
<< m2 >>
rect 177 25 178 26 
<< m1 >>
rect 178 25 179 26 
<< m2 >>
rect 178 25 179 26 
<< m1 >>
rect 179 25 180 26 
<< m2 >>
rect 179 25 180 26 
<< m1 >>
rect 180 25 181 26 
<< m2 >>
rect 180 25 181 26 
<< m1 >>
rect 181 25 182 26 
<< m2 >>
rect 181 25 182 26 
<< m1 >>
rect 182 25 183 26 
<< m2 >>
rect 182 25 183 26 
<< m1 >>
rect 183 25 184 26 
<< m2 >>
rect 183 25 184 26 
<< m1 >>
rect 184 25 185 26 
<< m2 >>
rect 184 25 185 26 
<< m1 >>
rect 185 25 186 26 
<< m2 >>
rect 185 25 186 26 
<< m1 >>
rect 186 25 187 26 
<< m2 >>
rect 186 25 187 26 
<< m1 >>
rect 187 25 188 26 
<< m2 >>
rect 187 25 188 26 
<< m1 >>
rect 188 25 189 26 
<< m2 >>
rect 188 25 189 26 
<< m1 >>
rect 189 25 190 26 
<< m2 >>
rect 189 25 190 26 
<< m1 >>
rect 190 25 191 26 
<< m2 >>
rect 190 25 191 26 
<< m1 >>
rect 191 25 192 26 
<< m2 >>
rect 191 25 192 26 
<< m1 >>
rect 192 25 193 26 
<< m2 >>
rect 192 25 193 26 
<< m1 >>
rect 193 25 194 26 
<< m2 >>
rect 193 25 194 26 
<< m1 >>
rect 194 25 195 26 
<< m2 >>
rect 194 25 195 26 
<< m1 >>
rect 195 25 196 26 
<< m2 >>
rect 195 25 196 26 
<< m1 >>
rect 196 25 197 26 
<< m2 >>
rect 196 25 197 26 
<< m1 >>
rect 197 25 198 26 
<< m2 >>
rect 197 25 198 26 
<< m1 >>
rect 198 25 199 26 
<< m2 >>
rect 198 25 199 26 
<< m2 >>
rect 199 25 200 26 
<< m1 >>
rect 200 25 201 26 
<< m2 >>
rect 200 25 201 26 
<< m1 >>
rect 201 25 202 26 
<< m2 >>
rect 201 25 202 26 
<< m1 >>
rect 202 25 203 26 
<< m2 >>
rect 202 25 203 26 
<< m1 >>
rect 203 25 204 26 
<< m1 >>
rect 204 25 205 26 
<< m1 >>
rect 205 25 206 26 
<< m1 >>
rect 206 25 207 26 
<< m1 >>
rect 207 25 208 26 
<< m1 >>
rect 208 25 209 26 
<< m1 >>
rect 209 25 210 26 
<< m1 >>
rect 210 25 211 26 
<< m1 >>
rect 211 25 212 26 
<< m1 >>
rect 212 25 213 26 
<< m1 >>
rect 213 25 214 26 
<< m1 >>
rect 214 25 215 26 
<< m1 >>
rect 215 25 216 26 
<< m1 >>
rect 216 25 217 26 
<< m1 >>
rect 217 25 218 26 
<< m1 >>
rect 218 25 219 26 
<< m1 >>
rect 219 25 220 26 
<< m1 >>
rect 220 25 221 26 
<< m1 >>
rect 221 25 222 26 
<< m1 >>
rect 222 25 223 26 
<< m1 >>
rect 223 25 224 26 
<< m1 >>
rect 224 25 225 26 
<< m1 >>
rect 225 25 226 26 
<< m2 >>
rect 225 25 226 26 
<< m1 >>
rect 226 25 227 26 
<< m1 >>
rect 227 25 228 26 
<< m1 >>
rect 228 25 229 26 
<< m1 >>
rect 229 25 230 26 
<< m1 >>
rect 230 25 231 26 
<< m1 >>
rect 231 25 232 26 
<< m1 >>
rect 232 25 233 26 
<< m1 >>
rect 233 25 234 26 
<< m1 >>
rect 234 25 235 26 
<< m1 >>
rect 235 25 236 26 
<< m1 >>
rect 236 25 237 26 
<< m1 >>
rect 237 25 238 26 
<< m1 >>
rect 238 25 239 26 
<< m1 >>
rect 239 25 240 26 
<< m1 >>
rect 240 25 241 26 
<< m1 >>
rect 241 25 242 26 
<< m1 >>
rect 242 25 243 26 
<< m1 >>
rect 243 25 244 26 
<< m1 >>
rect 244 25 245 26 
<< m1 >>
rect 245 25 246 26 
<< m1 >>
rect 246 25 247 26 
<< m1 >>
rect 247 25 248 26 
<< m1 >>
rect 248 25 249 26 
<< m1 >>
rect 249 25 250 26 
<< m1 >>
rect 250 25 251 26 
<< m1 >>
rect 251 25 252 26 
<< m1 >>
rect 252 25 253 26 
<< m1 >>
rect 253 25 254 26 
<< m2 >>
rect 253 25 254 26 
<< m1 >>
rect 254 25 255 26 
<< m2 >>
rect 254 25 255 26 
<< m1 >>
rect 255 25 256 26 
<< m2 >>
rect 255 25 256 26 
<< m1 >>
rect 256 25 257 26 
<< m2 >>
rect 256 25 257 26 
<< m1 >>
rect 257 25 258 26 
<< m2 >>
rect 257 25 258 26 
<< m1 >>
rect 258 25 259 26 
<< m2 >>
rect 258 25 259 26 
<< m1 >>
rect 259 25 260 26 
<< m2 >>
rect 259 25 260 26 
<< m1 >>
rect 260 25 261 26 
<< m2 >>
rect 260 25 261 26 
<< m1 >>
rect 261 25 262 26 
<< m2 >>
rect 261 25 262 26 
<< m1 >>
rect 262 25 263 26 
<< m2 >>
rect 262 25 263 26 
<< m1 >>
rect 263 25 264 26 
<< m2 >>
rect 263 25 264 26 
<< m1 >>
rect 264 25 265 26 
<< m2 >>
rect 264 25 265 26 
<< m1 >>
rect 265 25 266 26 
<< m2 >>
rect 265 25 266 26 
<< m1 >>
rect 266 25 267 26 
<< m2 >>
rect 266 25 267 26 
<< m1 >>
rect 267 25 268 26 
<< m1 >>
rect 268 25 269 26 
<< m1 >>
rect 269 25 270 26 
<< m1 >>
rect 270 25 271 26 
<< m1 >>
rect 271 25 272 26 
<< m2 >>
rect 271 25 272 26 
<< m1 >>
rect 272 25 273 26 
<< m1 >>
rect 273 25 274 26 
<< m2 >>
rect 273 25 274 26 
<< m1 >>
rect 274 25 275 26 
<< m1 >>
rect 275 25 276 26 
<< m2 >>
rect 275 25 276 26 
<< m1 >>
rect 276 25 277 26 
<< m1 >>
rect 277 25 278 26 
<< m2 >>
rect 277 25 278 26 
<< m1 >>
rect 278 25 279 26 
<< m1 >>
rect 279 25 280 26 
<< m2 >>
rect 279 25 280 26 
<< m1 >>
rect 280 25 281 26 
<< m1 >>
rect 281 25 282 26 
<< m1 >>
rect 282 25 283 26 
<< m1 >>
rect 283 25 284 26 
<< m1 >>
rect 284 25 285 26 
<< m2 >>
rect 284 25 285 26 
<< m1 >>
rect 285 25 286 26 
<< m1 >>
rect 286 25 287 26 
<< m1 >>
rect 287 25 288 26 
<< m1 >>
rect 288 25 289 26 
<< m1 >>
rect 289 25 290 26 
<< m1 >>
rect 290 25 291 26 
<< m1 >>
rect 291 25 292 26 
<< m1 >>
rect 292 25 293 26 
<< m1 >>
rect 293 25 294 26 
<< m1 >>
rect 294 25 295 26 
<< m1 >>
rect 295 25 296 26 
<< m1 >>
rect 296 25 297 26 
<< m1 >>
rect 297 25 298 26 
<< m1 >>
rect 298 25 299 26 
<< m1 >>
rect 299 25 300 26 
<< m1 >>
rect 300 25 301 26 
<< m1 >>
rect 301 25 302 26 
<< m1 >>
rect 302 25 303 26 
<< m1 >>
rect 303 25 304 26 
<< m1 >>
rect 304 25 305 26 
<< m1 >>
rect 305 25 306 26 
<< m1 >>
rect 306 25 307 26 
<< m1 >>
rect 307 25 308 26 
<< m1 >>
rect 308 25 309 26 
<< m1 >>
rect 309 25 310 26 
<< m1 >>
rect 310 25 311 26 
<< m1 >>
rect 311 25 312 26 
<< m1 >>
rect 312 25 313 26 
<< m1 >>
rect 313 25 314 26 
<< m1 >>
rect 314 25 315 26 
<< m1 >>
rect 315 25 316 26 
<< m1 >>
rect 316 25 317 26 
<< m1 >>
rect 317 25 318 26 
<< m1 >>
rect 318 25 319 26 
<< m1 >>
rect 319 25 320 26 
<< m1 >>
rect 320 25 321 26 
<< m1 >>
rect 321 25 322 26 
<< m1 >>
rect 322 25 323 26 
<< m1 >>
rect 323 25 324 26 
<< m1 >>
rect 324 25 325 26 
<< m1 >>
rect 325 25 326 26 
<< m1 >>
rect 326 25 327 26 
<< m1 >>
rect 327 25 328 26 
<< m1 >>
rect 328 25 329 26 
<< m1 >>
rect 329 25 330 26 
<< m1 >>
rect 330 25 331 26 
<< m1 >>
rect 331 25 332 26 
<< m1 >>
rect 332 25 333 26 
<< m1 >>
rect 333 25 334 26 
<< m1 >>
rect 334 25 335 26 
<< m2 >>
rect 334 25 335 26 
<< m1 >>
rect 335 25 336 26 
<< m1 >>
rect 336 25 337 26 
<< m1 >>
rect 337 25 338 26 
<< m1 >>
rect 338 25 339 26 
<< m1 >>
rect 339 25 340 26 
<< m1 >>
rect 340 25 341 26 
<< m1 >>
rect 343 25 344 26 
<< m1 >>
rect 19 26 20 27 
<< m1 >>
rect 21 26 22 27 
<< m1 >>
rect 23 26 24 27 
<< m1 >>
rect 46 26 47 27 
<< m1 >>
rect 62 26 63 27 
<< m1 >>
rect 64 26 65 27 
<< m1 >>
rect 78 26 79 27 
<< m1 >>
rect 82 26 83 27 
<< m1 >>
rect 88 26 89 27 
<< m2 >>
rect 92 26 93 27 
<< m1 >>
rect 198 26 199 27 
<< m1 >>
rect 200 26 201 27 
<< m2 >>
rect 202 26 203 27 
<< m2 >>
rect 225 26 226 27 
<< m2 >>
rect 253 26 254 27 
<< m2 >>
rect 271 26 272 27 
<< m2 >>
rect 273 26 274 27 
<< m2 >>
rect 275 26 276 27 
<< m2 >>
rect 277 26 278 27 
<< m2 >>
rect 279 26 280 27 
<< m2 >>
rect 284 26 285 27 
<< m2 >>
rect 334 26 335 27 
<< m1 >>
rect 343 26 344 27 
<< m1 >>
rect 19 27 20 28 
<< m1 >>
rect 21 27 22 28 
<< m1 >>
rect 23 27 24 28 
<< m1 >>
rect 31 27 32 28 
<< m1 >>
rect 32 27 33 28 
<< m1 >>
rect 33 27 34 28 
<< m1 >>
rect 34 27 35 28 
<< m1 >>
rect 35 27 36 28 
<< m1 >>
rect 36 27 37 28 
<< m1 >>
rect 37 27 38 28 
<< m1 >>
rect 46 27 47 28 
<< m1 >>
rect 62 27 63 28 
<< m1 >>
rect 64 27 65 28 
<< m1 >>
rect 78 27 79 28 
<< m1 >>
rect 82 27 83 28 
<< m1 >>
rect 88 27 89 28 
<< m1 >>
rect 92 27 93 28 
<< m2 >>
rect 92 27 93 28 
<< m2c >>
rect 92 27 93 28 
<< m1 >>
rect 92 27 93 28 
<< m2 >>
rect 92 27 93 28 
<< m1 >>
rect 198 27 199 28 
<< m1 >>
rect 200 27 201 28 
<< m1 >>
rect 202 27 203 28 
<< m2 >>
rect 202 27 203 28 
<< m2c >>
rect 202 27 203 28 
<< m1 >>
rect 202 27 203 28 
<< m2 >>
rect 202 27 203 28 
<< m1 >>
rect 203 27 204 28 
<< m1 >>
rect 204 27 205 28 
<< m2 >>
rect 225 27 226 28 
<< m1 >>
rect 253 27 254 28 
<< m2 >>
rect 253 27 254 28 
<< m2c >>
rect 253 27 254 28 
<< m1 >>
rect 253 27 254 28 
<< m2 >>
rect 253 27 254 28 
<< m1 >>
rect 271 27 272 28 
<< m2 >>
rect 271 27 272 28 
<< m2c >>
rect 271 27 272 28 
<< m1 >>
rect 271 27 272 28 
<< m2 >>
rect 271 27 272 28 
<< m1 >>
rect 273 27 274 28 
<< m2 >>
rect 273 27 274 28 
<< m2c >>
rect 273 27 274 28 
<< m1 >>
rect 273 27 274 28 
<< m2 >>
rect 273 27 274 28 
<< m1 >>
rect 275 27 276 28 
<< m2 >>
rect 275 27 276 28 
<< m2c >>
rect 275 27 276 28 
<< m1 >>
rect 275 27 276 28 
<< m2 >>
rect 275 27 276 28 
<< m1 >>
rect 277 27 278 28 
<< m2 >>
rect 277 27 278 28 
<< m2c >>
rect 277 27 278 28 
<< m1 >>
rect 277 27 278 28 
<< m2 >>
rect 277 27 278 28 
<< m1 >>
rect 279 27 280 28 
<< m2 >>
rect 279 27 280 28 
<< m2c >>
rect 279 27 280 28 
<< m1 >>
rect 279 27 280 28 
<< m2 >>
rect 279 27 280 28 
<< m1 >>
rect 284 27 285 28 
<< m2 >>
rect 284 27 285 28 
<< m2c >>
rect 284 27 285 28 
<< m1 >>
rect 284 27 285 28 
<< m2 >>
rect 284 27 285 28 
<< m1 >>
rect 285 27 286 28 
<< m1 >>
rect 286 27 287 28 
<< m1 >>
rect 287 27 288 28 
<< m1 >>
rect 288 27 289 28 
<< m1 >>
rect 289 27 290 28 
<< m1 >>
rect 334 27 335 28 
<< m2 >>
rect 334 27 335 28 
<< m2c >>
rect 334 27 335 28 
<< m1 >>
rect 334 27 335 28 
<< m2 >>
rect 334 27 335 28 
<< m1 >>
rect 343 27 344 28 
<< m1 >>
rect 19 28 20 29 
<< m1 >>
rect 21 28 22 29 
<< m1 >>
rect 23 28 24 29 
<< m1 >>
rect 31 28 32 29 
<< m1 >>
rect 37 28 38 29 
<< m1 >>
rect 46 28 47 29 
<< m1 >>
rect 62 28 63 29 
<< m1 >>
rect 64 28 65 29 
<< m1 >>
rect 78 28 79 29 
<< m1 >>
rect 82 28 83 29 
<< m1 >>
rect 88 28 89 29 
<< m1 >>
rect 92 28 93 29 
<< m1 >>
rect 190 28 191 29 
<< m1 >>
rect 191 28 192 29 
<< m1 >>
rect 192 28 193 29 
<< m1 >>
rect 193 28 194 29 
<< m1 >>
rect 198 28 199 29 
<< m2 >>
rect 198 28 199 29 
<< m2c >>
rect 198 28 199 29 
<< m1 >>
rect 198 28 199 29 
<< m2 >>
rect 198 28 199 29 
<< m2 >>
rect 199 28 200 29 
<< m1 >>
rect 200 28 201 29 
<< m2 >>
rect 200 28 201 29 
<< m2 >>
rect 201 28 202 29 
<< m1 >>
rect 204 28 205 29 
<< m2 >>
rect 225 28 226 29 
<< m1 >>
rect 226 28 227 29 
<< m1 >>
rect 227 28 228 29 
<< m1 >>
rect 228 28 229 29 
<< m1 >>
rect 229 28 230 29 
<< m1 >>
rect 253 28 254 29 
<< m1 >>
rect 271 28 272 29 
<< m1 >>
rect 273 28 274 29 
<< m1 >>
rect 275 28 276 29 
<< m1 >>
rect 277 28 278 29 
<< m1 >>
rect 279 28 280 29 
<< m1 >>
rect 289 28 290 29 
<< m1 >>
rect 316 28 317 29 
<< m1 >>
rect 317 28 318 29 
<< m1 >>
rect 318 28 319 29 
<< m1 >>
rect 319 28 320 29 
<< m1 >>
rect 334 28 335 29 
<< m1 >>
rect 343 28 344 29 
<< m1 >>
rect 19 29 20 30 
<< m1 >>
rect 21 29 22 30 
<< m1 >>
rect 23 29 24 30 
<< m1 >>
rect 31 29 32 30 
<< m1 >>
rect 37 29 38 30 
<< m1 >>
rect 46 29 47 30 
<< m1 >>
rect 62 29 63 30 
<< m1 >>
rect 64 29 65 30 
<< m1 >>
rect 78 29 79 30 
<< m1 >>
rect 82 29 83 30 
<< m1 >>
rect 88 29 89 30 
<< m1 >>
rect 92 29 93 30 
<< m1 >>
rect 190 29 191 30 
<< m1 >>
rect 193 29 194 30 
<< m1 >>
rect 200 29 201 30 
<< m2 >>
rect 201 29 202 30 
<< m1 >>
rect 204 29 205 30 
<< m2 >>
rect 225 29 226 30 
<< m1 >>
rect 226 29 227 30 
<< m1 >>
rect 229 29 230 30 
<< m1 >>
rect 253 29 254 30 
<< m1 >>
rect 271 29 272 30 
<< m1 >>
rect 273 29 274 30 
<< m1 >>
rect 275 29 276 30 
<< m1 >>
rect 277 29 278 30 
<< m1 >>
rect 279 29 280 30 
<< m1 >>
rect 289 29 290 30 
<< m1 >>
rect 316 29 317 30 
<< m1 >>
rect 319 29 320 30 
<< m1 >>
rect 334 29 335 30 
<< m1 >>
rect 343 29 344 30 
<< pdiffusion >>
rect 12 30 13 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< pdiffusion >>
rect 15 30 16 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< m1 >>
rect 19 30 20 31 
<< m1 >>
rect 21 30 22 31 
<< m1 >>
rect 23 30 24 31 
<< pdiffusion >>
rect 30 30 31 31 
<< m1 >>
rect 31 30 32 31 
<< pdiffusion >>
rect 31 30 32 31 
<< pdiffusion >>
rect 32 30 33 31 
<< pdiffusion >>
rect 33 30 34 31 
<< pdiffusion >>
rect 34 30 35 31 
<< pdiffusion >>
rect 35 30 36 31 
<< m1 >>
rect 37 30 38 31 
<< m1 >>
rect 46 30 47 31 
<< pdiffusion >>
rect 48 30 49 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 62 30 63 31 
<< m1 >>
rect 64 30 65 31 
<< pdiffusion >>
rect 66 30 67 31 
<< pdiffusion >>
rect 67 30 68 31 
<< pdiffusion >>
rect 68 30 69 31 
<< pdiffusion >>
rect 69 30 70 31 
<< pdiffusion >>
rect 70 30 71 31 
<< pdiffusion >>
rect 71 30 72 31 
<< m1 >>
rect 78 30 79 31 
<< m1 >>
rect 82 30 83 31 
<< pdiffusion >>
rect 84 30 85 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< m1 >>
rect 88 30 89 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< m1 >>
rect 92 30 93 31 
<< pdiffusion >>
rect 102 30 103 31 
<< pdiffusion >>
rect 103 30 104 31 
<< pdiffusion >>
rect 104 30 105 31 
<< pdiffusion >>
rect 105 30 106 31 
<< pdiffusion >>
rect 106 30 107 31 
<< pdiffusion >>
rect 107 30 108 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< pdiffusion >>
rect 138 30 139 31 
<< pdiffusion >>
rect 139 30 140 31 
<< pdiffusion >>
rect 140 30 141 31 
<< pdiffusion >>
rect 141 30 142 31 
<< pdiffusion >>
rect 142 30 143 31 
<< pdiffusion >>
rect 143 30 144 31 
<< pdiffusion >>
rect 156 30 157 31 
<< pdiffusion >>
rect 157 30 158 31 
<< pdiffusion >>
rect 158 30 159 31 
<< pdiffusion >>
rect 159 30 160 31 
<< pdiffusion >>
rect 160 30 161 31 
<< pdiffusion >>
rect 161 30 162 31 
<< pdiffusion >>
rect 174 30 175 31 
<< pdiffusion >>
rect 175 30 176 31 
<< pdiffusion >>
rect 176 30 177 31 
<< pdiffusion >>
rect 177 30 178 31 
<< pdiffusion >>
rect 178 30 179 31 
<< pdiffusion >>
rect 179 30 180 31 
<< m1 >>
rect 190 30 191 31 
<< pdiffusion >>
rect 192 30 193 31 
<< m1 >>
rect 193 30 194 31 
<< pdiffusion >>
rect 193 30 194 31 
<< pdiffusion >>
rect 194 30 195 31 
<< pdiffusion >>
rect 195 30 196 31 
<< pdiffusion >>
rect 196 30 197 31 
<< pdiffusion >>
rect 197 30 198 31 
<< m1 >>
rect 200 30 201 31 
<< m2 >>
rect 201 30 202 31 
<< m1 >>
rect 204 30 205 31 
<< pdiffusion >>
rect 210 30 211 31 
<< pdiffusion >>
rect 211 30 212 31 
<< pdiffusion >>
rect 212 30 213 31 
<< pdiffusion >>
rect 213 30 214 31 
<< pdiffusion >>
rect 214 30 215 31 
<< pdiffusion >>
rect 215 30 216 31 
<< m2 >>
rect 225 30 226 31 
<< m1 >>
rect 226 30 227 31 
<< pdiffusion >>
rect 228 30 229 31 
<< m1 >>
rect 229 30 230 31 
<< pdiffusion >>
rect 229 30 230 31 
<< pdiffusion >>
rect 230 30 231 31 
<< pdiffusion >>
rect 231 30 232 31 
<< pdiffusion >>
rect 232 30 233 31 
<< pdiffusion >>
rect 233 30 234 31 
<< pdiffusion >>
rect 246 30 247 31 
<< pdiffusion >>
rect 247 30 248 31 
<< pdiffusion >>
rect 248 30 249 31 
<< pdiffusion >>
rect 249 30 250 31 
<< pdiffusion >>
rect 250 30 251 31 
<< pdiffusion >>
rect 251 30 252 31 
<< m1 >>
rect 253 30 254 31 
<< pdiffusion >>
rect 264 30 265 31 
<< pdiffusion >>
rect 265 30 266 31 
<< pdiffusion >>
rect 266 30 267 31 
<< pdiffusion >>
rect 267 30 268 31 
<< pdiffusion >>
rect 268 30 269 31 
<< pdiffusion >>
rect 269 30 270 31 
<< m1 >>
rect 271 30 272 31 
<< m1 >>
rect 273 30 274 31 
<< m1 >>
rect 275 30 276 31 
<< m1 >>
rect 277 30 278 31 
<< m1 >>
rect 279 30 280 31 
<< pdiffusion >>
rect 282 30 283 31 
<< pdiffusion >>
rect 283 30 284 31 
<< pdiffusion >>
rect 284 30 285 31 
<< pdiffusion >>
rect 285 30 286 31 
<< pdiffusion >>
rect 286 30 287 31 
<< pdiffusion >>
rect 287 30 288 31 
<< m1 >>
rect 289 30 290 31 
<< pdiffusion >>
rect 300 30 301 31 
<< pdiffusion >>
rect 301 30 302 31 
<< pdiffusion >>
rect 302 30 303 31 
<< pdiffusion >>
rect 303 30 304 31 
<< pdiffusion >>
rect 304 30 305 31 
<< pdiffusion >>
rect 305 30 306 31 
<< m1 >>
rect 316 30 317 31 
<< pdiffusion >>
rect 318 30 319 31 
<< m1 >>
rect 319 30 320 31 
<< pdiffusion >>
rect 319 30 320 31 
<< pdiffusion >>
rect 320 30 321 31 
<< pdiffusion >>
rect 321 30 322 31 
<< pdiffusion >>
rect 322 30 323 31 
<< pdiffusion >>
rect 323 30 324 31 
<< m1 >>
rect 334 30 335 31 
<< pdiffusion >>
rect 336 30 337 31 
<< pdiffusion >>
rect 337 30 338 31 
<< pdiffusion >>
rect 338 30 339 31 
<< pdiffusion >>
rect 339 30 340 31 
<< pdiffusion >>
rect 340 30 341 31 
<< pdiffusion >>
rect 341 30 342 31 
<< m1 >>
rect 343 30 344 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< m1 >>
rect 19 31 20 32 
<< m1 >>
rect 21 31 22 32 
<< m1 >>
rect 23 31 24 32 
<< pdiffusion >>
rect 30 31 31 32 
<< pdiffusion >>
rect 31 31 32 32 
<< pdiffusion >>
rect 32 31 33 32 
<< pdiffusion >>
rect 33 31 34 32 
<< pdiffusion >>
rect 34 31 35 32 
<< pdiffusion >>
rect 35 31 36 32 
<< m1 >>
rect 37 31 38 32 
<< m1 >>
rect 46 31 47 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 62 31 63 32 
<< m1 >>
rect 64 31 65 32 
<< pdiffusion >>
rect 66 31 67 32 
<< pdiffusion >>
rect 67 31 68 32 
<< pdiffusion >>
rect 68 31 69 32 
<< pdiffusion >>
rect 69 31 70 32 
<< pdiffusion >>
rect 70 31 71 32 
<< pdiffusion >>
rect 71 31 72 32 
<< m1 >>
rect 78 31 79 32 
<< m1 >>
rect 82 31 83 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< m1 >>
rect 92 31 93 32 
<< pdiffusion >>
rect 102 31 103 32 
<< pdiffusion >>
rect 103 31 104 32 
<< pdiffusion >>
rect 104 31 105 32 
<< pdiffusion >>
rect 105 31 106 32 
<< pdiffusion >>
rect 106 31 107 32 
<< pdiffusion >>
rect 107 31 108 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< pdiffusion >>
rect 138 31 139 32 
<< pdiffusion >>
rect 139 31 140 32 
<< pdiffusion >>
rect 140 31 141 32 
<< pdiffusion >>
rect 141 31 142 32 
<< pdiffusion >>
rect 142 31 143 32 
<< pdiffusion >>
rect 143 31 144 32 
<< pdiffusion >>
rect 156 31 157 32 
<< pdiffusion >>
rect 157 31 158 32 
<< pdiffusion >>
rect 158 31 159 32 
<< pdiffusion >>
rect 159 31 160 32 
<< pdiffusion >>
rect 160 31 161 32 
<< pdiffusion >>
rect 161 31 162 32 
<< pdiffusion >>
rect 174 31 175 32 
<< pdiffusion >>
rect 175 31 176 32 
<< pdiffusion >>
rect 176 31 177 32 
<< pdiffusion >>
rect 177 31 178 32 
<< pdiffusion >>
rect 178 31 179 32 
<< pdiffusion >>
rect 179 31 180 32 
<< m1 >>
rect 190 31 191 32 
<< pdiffusion >>
rect 192 31 193 32 
<< pdiffusion >>
rect 193 31 194 32 
<< pdiffusion >>
rect 194 31 195 32 
<< pdiffusion >>
rect 195 31 196 32 
<< pdiffusion >>
rect 196 31 197 32 
<< pdiffusion >>
rect 197 31 198 32 
<< m1 >>
rect 200 31 201 32 
<< m2 >>
rect 201 31 202 32 
<< m1 >>
rect 204 31 205 32 
<< pdiffusion >>
rect 210 31 211 32 
<< pdiffusion >>
rect 211 31 212 32 
<< pdiffusion >>
rect 212 31 213 32 
<< pdiffusion >>
rect 213 31 214 32 
<< pdiffusion >>
rect 214 31 215 32 
<< pdiffusion >>
rect 215 31 216 32 
<< m2 >>
rect 225 31 226 32 
<< m1 >>
rect 226 31 227 32 
<< pdiffusion >>
rect 228 31 229 32 
<< pdiffusion >>
rect 229 31 230 32 
<< pdiffusion >>
rect 230 31 231 32 
<< pdiffusion >>
rect 231 31 232 32 
<< pdiffusion >>
rect 232 31 233 32 
<< pdiffusion >>
rect 233 31 234 32 
<< pdiffusion >>
rect 246 31 247 32 
<< pdiffusion >>
rect 247 31 248 32 
<< pdiffusion >>
rect 248 31 249 32 
<< pdiffusion >>
rect 249 31 250 32 
<< pdiffusion >>
rect 250 31 251 32 
<< pdiffusion >>
rect 251 31 252 32 
<< m1 >>
rect 253 31 254 32 
<< pdiffusion >>
rect 264 31 265 32 
<< pdiffusion >>
rect 265 31 266 32 
<< pdiffusion >>
rect 266 31 267 32 
<< pdiffusion >>
rect 267 31 268 32 
<< pdiffusion >>
rect 268 31 269 32 
<< pdiffusion >>
rect 269 31 270 32 
<< m1 >>
rect 271 31 272 32 
<< m1 >>
rect 273 31 274 32 
<< m1 >>
rect 275 31 276 32 
<< m1 >>
rect 277 31 278 32 
<< m1 >>
rect 279 31 280 32 
<< pdiffusion >>
rect 282 31 283 32 
<< pdiffusion >>
rect 283 31 284 32 
<< pdiffusion >>
rect 284 31 285 32 
<< pdiffusion >>
rect 285 31 286 32 
<< pdiffusion >>
rect 286 31 287 32 
<< pdiffusion >>
rect 287 31 288 32 
<< m1 >>
rect 289 31 290 32 
<< pdiffusion >>
rect 300 31 301 32 
<< pdiffusion >>
rect 301 31 302 32 
<< pdiffusion >>
rect 302 31 303 32 
<< pdiffusion >>
rect 303 31 304 32 
<< pdiffusion >>
rect 304 31 305 32 
<< pdiffusion >>
rect 305 31 306 32 
<< m1 >>
rect 316 31 317 32 
<< pdiffusion >>
rect 318 31 319 32 
<< pdiffusion >>
rect 319 31 320 32 
<< pdiffusion >>
rect 320 31 321 32 
<< pdiffusion >>
rect 321 31 322 32 
<< pdiffusion >>
rect 322 31 323 32 
<< pdiffusion >>
rect 323 31 324 32 
<< m1 >>
rect 334 31 335 32 
<< pdiffusion >>
rect 336 31 337 32 
<< pdiffusion >>
rect 337 31 338 32 
<< pdiffusion >>
rect 338 31 339 32 
<< pdiffusion >>
rect 339 31 340 32 
<< pdiffusion >>
rect 340 31 341 32 
<< pdiffusion >>
rect 341 31 342 32 
<< m1 >>
rect 343 31 344 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< m1 >>
rect 19 32 20 33 
<< m1 >>
rect 21 32 22 33 
<< m1 >>
rect 23 32 24 33 
<< pdiffusion >>
rect 30 32 31 33 
<< pdiffusion >>
rect 31 32 32 33 
<< pdiffusion >>
rect 32 32 33 33 
<< pdiffusion >>
rect 33 32 34 33 
<< pdiffusion >>
rect 34 32 35 33 
<< pdiffusion >>
rect 35 32 36 33 
<< m1 >>
rect 37 32 38 33 
<< m1 >>
rect 46 32 47 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 62 32 63 33 
<< m1 >>
rect 64 32 65 33 
<< pdiffusion >>
rect 66 32 67 33 
<< pdiffusion >>
rect 67 32 68 33 
<< pdiffusion >>
rect 68 32 69 33 
<< pdiffusion >>
rect 69 32 70 33 
<< pdiffusion >>
rect 70 32 71 33 
<< pdiffusion >>
rect 71 32 72 33 
<< m1 >>
rect 78 32 79 33 
<< m1 >>
rect 82 32 83 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< m1 >>
rect 92 32 93 33 
<< pdiffusion >>
rect 102 32 103 33 
<< pdiffusion >>
rect 103 32 104 33 
<< pdiffusion >>
rect 104 32 105 33 
<< pdiffusion >>
rect 105 32 106 33 
<< pdiffusion >>
rect 106 32 107 33 
<< pdiffusion >>
rect 107 32 108 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< pdiffusion >>
rect 138 32 139 33 
<< pdiffusion >>
rect 139 32 140 33 
<< pdiffusion >>
rect 140 32 141 33 
<< pdiffusion >>
rect 141 32 142 33 
<< pdiffusion >>
rect 142 32 143 33 
<< pdiffusion >>
rect 143 32 144 33 
<< pdiffusion >>
rect 156 32 157 33 
<< pdiffusion >>
rect 157 32 158 33 
<< pdiffusion >>
rect 158 32 159 33 
<< pdiffusion >>
rect 159 32 160 33 
<< pdiffusion >>
rect 160 32 161 33 
<< pdiffusion >>
rect 161 32 162 33 
<< pdiffusion >>
rect 174 32 175 33 
<< pdiffusion >>
rect 175 32 176 33 
<< pdiffusion >>
rect 176 32 177 33 
<< pdiffusion >>
rect 177 32 178 33 
<< pdiffusion >>
rect 178 32 179 33 
<< pdiffusion >>
rect 179 32 180 33 
<< m1 >>
rect 190 32 191 33 
<< pdiffusion >>
rect 192 32 193 33 
<< pdiffusion >>
rect 193 32 194 33 
<< pdiffusion >>
rect 194 32 195 33 
<< pdiffusion >>
rect 195 32 196 33 
<< pdiffusion >>
rect 196 32 197 33 
<< pdiffusion >>
rect 197 32 198 33 
<< m1 >>
rect 200 32 201 33 
<< m2 >>
rect 201 32 202 33 
<< m1 >>
rect 204 32 205 33 
<< pdiffusion >>
rect 210 32 211 33 
<< pdiffusion >>
rect 211 32 212 33 
<< pdiffusion >>
rect 212 32 213 33 
<< pdiffusion >>
rect 213 32 214 33 
<< pdiffusion >>
rect 214 32 215 33 
<< pdiffusion >>
rect 215 32 216 33 
<< m2 >>
rect 225 32 226 33 
<< m1 >>
rect 226 32 227 33 
<< pdiffusion >>
rect 228 32 229 33 
<< pdiffusion >>
rect 229 32 230 33 
<< pdiffusion >>
rect 230 32 231 33 
<< pdiffusion >>
rect 231 32 232 33 
<< pdiffusion >>
rect 232 32 233 33 
<< pdiffusion >>
rect 233 32 234 33 
<< pdiffusion >>
rect 246 32 247 33 
<< pdiffusion >>
rect 247 32 248 33 
<< pdiffusion >>
rect 248 32 249 33 
<< pdiffusion >>
rect 249 32 250 33 
<< pdiffusion >>
rect 250 32 251 33 
<< pdiffusion >>
rect 251 32 252 33 
<< m1 >>
rect 253 32 254 33 
<< pdiffusion >>
rect 264 32 265 33 
<< pdiffusion >>
rect 265 32 266 33 
<< pdiffusion >>
rect 266 32 267 33 
<< pdiffusion >>
rect 267 32 268 33 
<< pdiffusion >>
rect 268 32 269 33 
<< pdiffusion >>
rect 269 32 270 33 
<< m1 >>
rect 271 32 272 33 
<< m1 >>
rect 273 32 274 33 
<< m1 >>
rect 275 32 276 33 
<< m1 >>
rect 277 32 278 33 
<< m1 >>
rect 279 32 280 33 
<< pdiffusion >>
rect 282 32 283 33 
<< pdiffusion >>
rect 283 32 284 33 
<< pdiffusion >>
rect 284 32 285 33 
<< pdiffusion >>
rect 285 32 286 33 
<< pdiffusion >>
rect 286 32 287 33 
<< pdiffusion >>
rect 287 32 288 33 
<< m1 >>
rect 289 32 290 33 
<< pdiffusion >>
rect 300 32 301 33 
<< pdiffusion >>
rect 301 32 302 33 
<< pdiffusion >>
rect 302 32 303 33 
<< pdiffusion >>
rect 303 32 304 33 
<< pdiffusion >>
rect 304 32 305 33 
<< pdiffusion >>
rect 305 32 306 33 
<< m1 >>
rect 316 32 317 33 
<< pdiffusion >>
rect 318 32 319 33 
<< pdiffusion >>
rect 319 32 320 33 
<< pdiffusion >>
rect 320 32 321 33 
<< pdiffusion >>
rect 321 32 322 33 
<< pdiffusion >>
rect 322 32 323 33 
<< pdiffusion >>
rect 323 32 324 33 
<< m1 >>
rect 334 32 335 33 
<< pdiffusion >>
rect 336 32 337 33 
<< pdiffusion >>
rect 337 32 338 33 
<< pdiffusion >>
rect 338 32 339 33 
<< pdiffusion >>
rect 339 32 340 33 
<< pdiffusion >>
rect 340 32 341 33 
<< pdiffusion >>
rect 341 32 342 33 
<< m1 >>
rect 343 32 344 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< m1 >>
rect 19 33 20 34 
<< m1 >>
rect 21 33 22 34 
<< m1 >>
rect 23 33 24 34 
<< pdiffusion >>
rect 30 33 31 34 
<< pdiffusion >>
rect 31 33 32 34 
<< pdiffusion >>
rect 32 33 33 34 
<< pdiffusion >>
rect 33 33 34 34 
<< pdiffusion >>
rect 34 33 35 34 
<< pdiffusion >>
rect 35 33 36 34 
<< m1 >>
rect 37 33 38 34 
<< m1 >>
rect 46 33 47 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 62 33 63 34 
<< m1 >>
rect 64 33 65 34 
<< pdiffusion >>
rect 66 33 67 34 
<< pdiffusion >>
rect 67 33 68 34 
<< pdiffusion >>
rect 68 33 69 34 
<< pdiffusion >>
rect 69 33 70 34 
<< pdiffusion >>
rect 70 33 71 34 
<< pdiffusion >>
rect 71 33 72 34 
<< m1 >>
rect 78 33 79 34 
<< m1 >>
rect 82 33 83 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< m1 >>
rect 92 33 93 34 
<< pdiffusion >>
rect 102 33 103 34 
<< pdiffusion >>
rect 103 33 104 34 
<< pdiffusion >>
rect 104 33 105 34 
<< pdiffusion >>
rect 105 33 106 34 
<< pdiffusion >>
rect 106 33 107 34 
<< pdiffusion >>
rect 107 33 108 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< pdiffusion >>
rect 138 33 139 34 
<< pdiffusion >>
rect 139 33 140 34 
<< pdiffusion >>
rect 140 33 141 34 
<< pdiffusion >>
rect 141 33 142 34 
<< pdiffusion >>
rect 142 33 143 34 
<< pdiffusion >>
rect 143 33 144 34 
<< pdiffusion >>
rect 156 33 157 34 
<< pdiffusion >>
rect 157 33 158 34 
<< pdiffusion >>
rect 158 33 159 34 
<< pdiffusion >>
rect 159 33 160 34 
<< pdiffusion >>
rect 160 33 161 34 
<< pdiffusion >>
rect 161 33 162 34 
<< pdiffusion >>
rect 174 33 175 34 
<< pdiffusion >>
rect 175 33 176 34 
<< pdiffusion >>
rect 176 33 177 34 
<< pdiffusion >>
rect 177 33 178 34 
<< pdiffusion >>
rect 178 33 179 34 
<< pdiffusion >>
rect 179 33 180 34 
<< m1 >>
rect 190 33 191 34 
<< pdiffusion >>
rect 192 33 193 34 
<< pdiffusion >>
rect 193 33 194 34 
<< pdiffusion >>
rect 194 33 195 34 
<< pdiffusion >>
rect 195 33 196 34 
<< pdiffusion >>
rect 196 33 197 34 
<< pdiffusion >>
rect 197 33 198 34 
<< m1 >>
rect 200 33 201 34 
<< m2 >>
rect 201 33 202 34 
<< m1 >>
rect 204 33 205 34 
<< pdiffusion >>
rect 210 33 211 34 
<< pdiffusion >>
rect 211 33 212 34 
<< pdiffusion >>
rect 212 33 213 34 
<< pdiffusion >>
rect 213 33 214 34 
<< pdiffusion >>
rect 214 33 215 34 
<< pdiffusion >>
rect 215 33 216 34 
<< m2 >>
rect 225 33 226 34 
<< m1 >>
rect 226 33 227 34 
<< pdiffusion >>
rect 228 33 229 34 
<< pdiffusion >>
rect 229 33 230 34 
<< pdiffusion >>
rect 230 33 231 34 
<< pdiffusion >>
rect 231 33 232 34 
<< pdiffusion >>
rect 232 33 233 34 
<< pdiffusion >>
rect 233 33 234 34 
<< pdiffusion >>
rect 246 33 247 34 
<< pdiffusion >>
rect 247 33 248 34 
<< pdiffusion >>
rect 248 33 249 34 
<< pdiffusion >>
rect 249 33 250 34 
<< pdiffusion >>
rect 250 33 251 34 
<< pdiffusion >>
rect 251 33 252 34 
<< m1 >>
rect 253 33 254 34 
<< pdiffusion >>
rect 264 33 265 34 
<< pdiffusion >>
rect 265 33 266 34 
<< pdiffusion >>
rect 266 33 267 34 
<< pdiffusion >>
rect 267 33 268 34 
<< pdiffusion >>
rect 268 33 269 34 
<< pdiffusion >>
rect 269 33 270 34 
<< m1 >>
rect 271 33 272 34 
<< m1 >>
rect 273 33 274 34 
<< m1 >>
rect 275 33 276 34 
<< m1 >>
rect 277 33 278 34 
<< m1 >>
rect 279 33 280 34 
<< pdiffusion >>
rect 282 33 283 34 
<< pdiffusion >>
rect 283 33 284 34 
<< pdiffusion >>
rect 284 33 285 34 
<< pdiffusion >>
rect 285 33 286 34 
<< pdiffusion >>
rect 286 33 287 34 
<< pdiffusion >>
rect 287 33 288 34 
<< m1 >>
rect 289 33 290 34 
<< pdiffusion >>
rect 300 33 301 34 
<< pdiffusion >>
rect 301 33 302 34 
<< pdiffusion >>
rect 302 33 303 34 
<< pdiffusion >>
rect 303 33 304 34 
<< pdiffusion >>
rect 304 33 305 34 
<< pdiffusion >>
rect 305 33 306 34 
<< m1 >>
rect 316 33 317 34 
<< pdiffusion >>
rect 318 33 319 34 
<< pdiffusion >>
rect 319 33 320 34 
<< pdiffusion >>
rect 320 33 321 34 
<< pdiffusion >>
rect 321 33 322 34 
<< pdiffusion >>
rect 322 33 323 34 
<< pdiffusion >>
rect 323 33 324 34 
<< m1 >>
rect 334 33 335 34 
<< pdiffusion >>
rect 336 33 337 34 
<< pdiffusion >>
rect 337 33 338 34 
<< pdiffusion >>
rect 338 33 339 34 
<< pdiffusion >>
rect 339 33 340 34 
<< pdiffusion >>
rect 340 33 341 34 
<< pdiffusion >>
rect 341 33 342 34 
<< m1 >>
rect 343 33 344 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< m1 >>
rect 19 34 20 35 
<< m1 >>
rect 21 34 22 35 
<< m1 >>
rect 23 34 24 35 
<< pdiffusion >>
rect 30 34 31 35 
<< pdiffusion >>
rect 31 34 32 35 
<< pdiffusion >>
rect 32 34 33 35 
<< pdiffusion >>
rect 33 34 34 35 
<< pdiffusion >>
rect 34 34 35 35 
<< pdiffusion >>
rect 35 34 36 35 
<< m1 >>
rect 37 34 38 35 
<< m1 >>
rect 46 34 47 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 62 34 63 35 
<< m1 >>
rect 64 34 65 35 
<< pdiffusion >>
rect 66 34 67 35 
<< pdiffusion >>
rect 67 34 68 35 
<< pdiffusion >>
rect 68 34 69 35 
<< pdiffusion >>
rect 69 34 70 35 
<< pdiffusion >>
rect 70 34 71 35 
<< pdiffusion >>
rect 71 34 72 35 
<< m1 >>
rect 78 34 79 35 
<< m1 >>
rect 82 34 83 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< m1 >>
rect 92 34 93 35 
<< pdiffusion >>
rect 102 34 103 35 
<< pdiffusion >>
rect 103 34 104 35 
<< pdiffusion >>
rect 104 34 105 35 
<< pdiffusion >>
rect 105 34 106 35 
<< pdiffusion >>
rect 106 34 107 35 
<< pdiffusion >>
rect 107 34 108 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< pdiffusion >>
rect 138 34 139 35 
<< pdiffusion >>
rect 139 34 140 35 
<< pdiffusion >>
rect 140 34 141 35 
<< pdiffusion >>
rect 141 34 142 35 
<< pdiffusion >>
rect 142 34 143 35 
<< pdiffusion >>
rect 143 34 144 35 
<< pdiffusion >>
rect 156 34 157 35 
<< pdiffusion >>
rect 157 34 158 35 
<< pdiffusion >>
rect 158 34 159 35 
<< pdiffusion >>
rect 159 34 160 35 
<< pdiffusion >>
rect 160 34 161 35 
<< pdiffusion >>
rect 161 34 162 35 
<< pdiffusion >>
rect 174 34 175 35 
<< pdiffusion >>
rect 175 34 176 35 
<< pdiffusion >>
rect 176 34 177 35 
<< pdiffusion >>
rect 177 34 178 35 
<< pdiffusion >>
rect 178 34 179 35 
<< pdiffusion >>
rect 179 34 180 35 
<< m1 >>
rect 190 34 191 35 
<< pdiffusion >>
rect 192 34 193 35 
<< pdiffusion >>
rect 193 34 194 35 
<< pdiffusion >>
rect 194 34 195 35 
<< pdiffusion >>
rect 195 34 196 35 
<< pdiffusion >>
rect 196 34 197 35 
<< pdiffusion >>
rect 197 34 198 35 
<< m1 >>
rect 200 34 201 35 
<< m2 >>
rect 201 34 202 35 
<< m1 >>
rect 204 34 205 35 
<< pdiffusion >>
rect 210 34 211 35 
<< pdiffusion >>
rect 211 34 212 35 
<< pdiffusion >>
rect 212 34 213 35 
<< pdiffusion >>
rect 213 34 214 35 
<< pdiffusion >>
rect 214 34 215 35 
<< pdiffusion >>
rect 215 34 216 35 
<< m2 >>
rect 225 34 226 35 
<< m1 >>
rect 226 34 227 35 
<< pdiffusion >>
rect 228 34 229 35 
<< pdiffusion >>
rect 229 34 230 35 
<< pdiffusion >>
rect 230 34 231 35 
<< pdiffusion >>
rect 231 34 232 35 
<< pdiffusion >>
rect 232 34 233 35 
<< pdiffusion >>
rect 233 34 234 35 
<< pdiffusion >>
rect 246 34 247 35 
<< pdiffusion >>
rect 247 34 248 35 
<< pdiffusion >>
rect 248 34 249 35 
<< pdiffusion >>
rect 249 34 250 35 
<< pdiffusion >>
rect 250 34 251 35 
<< pdiffusion >>
rect 251 34 252 35 
<< m1 >>
rect 253 34 254 35 
<< pdiffusion >>
rect 264 34 265 35 
<< pdiffusion >>
rect 265 34 266 35 
<< pdiffusion >>
rect 266 34 267 35 
<< pdiffusion >>
rect 267 34 268 35 
<< pdiffusion >>
rect 268 34 269 35 
<< pdiffusion >>
rect 269 34 270 35 
<< m1 >>
rect 271 34 272 35 
<< m1 >>
rect 273 34 274 35 
<< m1 >>
rect 275 34 276 35 
<< m1 >>
rect 277 34 278 35 
<< m1 >>
rect 279 34 280 35 
<< pdiffusion >>
rect 282 34 283 35 
<< pdiffusion >>
rect 283 34 284 35 
<< pdiffusion >>
rect 284 34 285 35 
<< pdiffusion >>
rect 285 34 286 35 
<< pdiffusion >>
rect 286 34 287 35 
<< pdiffusion >>
rect 287 34 288 35 
<< m1 >>
rect 289 34 290 35 
<< pdiffusion >>
rect 300 34 301 35 
<< pdiffusion >>
rect 301 34 302 35 
<< pdiffusion >>
rect 302 34 303 35 
<< pdiffusion >>
rect 303 34 304 35 
<< pdiffusion >>
rect 304 34 305 35 
<< pdiffusion >>
rect 305 34 306 35 
<< m1 >>
rect 316 34 317 35 
<< pdiffusion >>
rect 318 34 319 35 
<< pdiffusion >>
rect 319 34 320 35 
<< pdiffusion >>
rect 320 34 321 35 
<< pdiffusion >>
rect 321 34 322 35 
<< pdiffusion >>
rect 322 34 323 35 
<< pdiffusion >>
rect 323 34 324 35 
<< m1 >>
rect 334 34 335 35 
<< pdiffusion >>
rect 336 34 337 35 
<< pdiffusion >>
rect 337 34 338 35 
<< pdiffusion >>
rect 338 34 339 35 
<< pdiffusion >>
rect 339 34 340 35 
<< pdiffusion >>
rect 340 34 341 35 
<< pdiffusion >>
rect 341 34 342 35 
<< m1 >>
rect 343 34 344 35 
<< pdiffusion >>
rect 12 35 13 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< m1 >>
rect 19 35 20 36 
<< m1 >>
rect 21 35 22 36 
<< m1 >>
rect 23 35 24 36 
<< pdiffusion >>
rect 30 35 31 36 
<< pdiffusion >>
rect 31 35 32 36 
<< pdiffusion >>
rect 32 35 33 36 
<< pdiffusion >>
rect 33 35 34 36 
<< pdiffusion >>
rect 34 35 35 36 
<< pdiffusion >>
rect 35 35 36 36 
<< m1 >>
rect 37 35 38 36 
<< m1 >>
rect 46 35 47 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 62 35 63 36 
<< m1 >>
rect 64 35 65 36 
<< pdiffusion >>
rect 66 35 67 36 
<< pdiffusion >>
rect 67 35 68 36 
<< pdiffusion >>
rect 68 35 69 36 
<< pdiffusion >>
rect 69 35 70 36 
<< pdiffusion >>
rect 70 35 71 36 
<< pdiffusion >>
rect 71 35 72 36 
<< m1 >>
rect 78 35 79 36 
<< m1 >>
rect 82 35 83 36 
<< pdiffusion >>
rect 84 35 85 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< m1 >>
rect 92 35 93 36 
<< pdiffusion >>
rect 102 35 103 36 
<< pdiffusion >>
rect 103 35 104 36 
<< pdiffusion >>
rect 104 35 105 36 
<< pdiffusion >>
rect 105 35 106 36 
<< pdiffusion >>
rect 106 35 107 36 
<< pdiffusion >>
rect 107 35 108 36 
<< pdiffusion >>
rect 120 35 121 36 
<< m1 >>
rect 121 35 122 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< pdiffusion >>
rect 138 35 139 36 
<< pdiffusion >>
rect 139 35 140 36 
<< pdiffusion >>
rect 140 35 141 36 
<< pdiffusion >>
rect 141 35 142 36 
<< pdiffusion >>
rect 142 35 143 36 
<< pdiffusion >>
rect 143 35 144 36 
<< pdiffusion >>
rect 156 35 157 36 
<< pdiffusion >>
rect 157 35 158 36 
<< pdiffusion >>
rect 158 35 159 36 
<< pdiffusion >>
rect 159 35 160 36 
<< pdiffusion >>
rect 160 35 161 36 
<< pdiffusion >>
rect 161 35 162 36 
<< pdiffusion >>
rect 174 35 175 36 
<< pdiffusion >>
rect 175 35 176 36 
<< pdiffusion >>
rect 176 35 177 36 
<< pdiffusion >>
rect 177 35 178 36 
<< pdiffusion >>
rect 178 35 179 36 
<< pdiffusion >>
rect 179 35 180 36 
<< m1 >>
rect 190 35 191 36 
<< pdiffusion >>
rect 192 35 193 36 
<< pdiffusion >>
rect 193 35 194 36 
<< pdiffusion >>
rect 194 35 195 36 
<< pdiffusion >>
rect 195 35 196 36 
<< pdiffusion >>
rect 196 35 197 36 
<< pdiffusion >>
rect 197 35 198 36 
<< m1 >>
rect 200 35 201 36 
<< m2 >>
rect 201 35 202 36 
<< m1 >>
rect 204 35 205 36 
<< pdiffusion >>
rect 210 35 211 36 
<< pdiffusion >>
rect 211 35 212 36 
<< pdiffusion >>
rect 212 35 213 36 
<< pdiffusion >>
rect 213 35 214 36 
<< pdiffusion >>
rect 214 35 215 36 
<< pdiffusion >>
rect 215 35 216 36 
<< m2 >>
rect 225 35 226 36 
<< m1 >>
rect 226 35 227 36 
<< pdiffusion >>
rect 228 35 229 36 
<< pdiffusion >>
rect 229 35 230 36 
<< pdiffusion >>
rect 230 35 231 36 
<< pdiffusion >>
rect 231 35 232 36 
<< pdiffusion >>
rect 232 35 233 36 
<< pdiffusion >>
rect 233 35 234 36 
<< pdiffusion >>
rect 246 35 247 36 
<< m1 >>
rect 247 35 248 36 
<< pdiffusion >>
rect 247 35 248 36 
<< pdiffusion >>
rect 248 35 249 36 
<< pdiffusion >>
rect 249 35 250 36 
<< pdiffusion >>
rect 250 35 251 36 
<< pdiffusion >>
rect 251 35 252 36 
<< m1 >>
rect 253 35 254 36 
<< pdiffusion >>
rect 264 35 265 36 
<< m1 >>
rect 265 35 266 36 
<< pdiffusion >>
rect 265 35 266 36 
<< pdiffusion >>
rect 266 35 267 36 
<< pdiffusion >>
rect 267 35 268 36 
<< pdiffusion >>
rect 268 35 269 36 
<< pdiffusion >>
rect 269 35 270 36 
<< m1 >>
rect 271 35 272 36 
<< m1 >>
rect 273 35 274 36 
<< m1 >>
rect 275 35 276 36 
<< m1 >>
rect 277 35 278 36 
<< m1 >>
rect 279 35 280 36 
<< pdiffusion >>
rect 282 35 283 36 
<< pdiffusion >>
rect 283 35 284 36 
<< pdiffusion >>
rect 284 35 285 36 
<< pdiffusion >>
rect 285 35 286 36 
<< pdiffusion >>
rect 286 35 287 36 
<< pdiffusion >>
rect 287 35 288 36 
<< m1 >>
rect 289 35 290 36 
<< pdiffusion >>
rect 300 35 301 36 
<< pdiffusion >>
rect 301 35 302 36 
<< pdiffusion >>
rect 302 35 303 36 
<< pdiffusion >>
rect 303 35 304 36 
<< m1 >>
rect 304 35 305 36 
<< pdiffusion >>
rect 304 35 305 36 
<< pdiffusion >>
rect 305 35 306 36 
<< m1 >>
rect 316 35 317 36 
<< pdiffusion >>
rect 318 35 319 36 
<< pdiffusion >>
rect 319 35 320 36 
<< pdiffusion >>
rect 320 35 321 36 
<< pdiffusion >>
rect 321 35 322 36 
<< pdiffusion >>
rect 322 35 323 36 
<< pdiffusion >>
rect 323 35 324 36 
<< m1 >>
rect 334 35 335 36 
<< pdiffusion >>
rect 336 35 337 36 
<< m1 >>
rect 337 35 338 36 
<< pdiffusion >>
rect 337 35 338 36 
<< pdiffusion >>
rect 338 35 339 36 
<< pdiffusion >>
rect 339 35 340 36 
<< m1 >>
rect 340 35 341 36 
<< pdiffusion >>
rect 340 35 341 36 
<< pdiffusion >>
rect 341 35 342 36 
<< m1 >>
rect 343 35 344 36 
<< m1 >>
rect 19 36 20 37 
<< m1 >>
rect 21 36 22 37 
<< m1 >>
rect 23 36 24 37 
<< m1 >>
rect 37 36 38 37 
<< m1 >>
rect 46 36 47 37 
<< m1 >>
rect 62 36 63 37 
<< m1 >>
rect 64 36 65 37 
<< m1 >>
rect 78 36 79 37 
<< m1 >>
rect 82 36 83 37 
<< m1 >>
rect 92 36 93 37 
<< m1 >>
rect 121 36 122 37 
<< m1 >>
rect 190 36 191 37 
<< m1 >>
rect 200 36 201 37 
<< m2 >>
rect 201 36 202 37 
<< m1 >>
rect 204 36 205 37 
<< m2 >>
rect 225 36 226 37 
<< m1 >>
rect 226 36 227 37 
<< m1 >>
rect 247 36 248 37 
<< m1 >>
rect 253 36 254 37 
<< m1 >>
rect 265 36 266 37 
<< m1 >>
rect 271 36 272 37 
<< m1 >>
rect 273 36 274 37 
<< m1 >>
rect 275 36 276 37 
<< m1 >>
rect 277 36 278 37 
<< m1 >>
rect 279 36 280 37 
<< m1 >>
rect 289 36 290 37 
<< m1 >>
rect 304 36 305 37 
<< m1 >>
rect 316 36 317 37 
<< m2 >>
rect 316 36 317 37 
<< m2c >>
rect 316 36 317 37 
<< m1 >>
rect 316 36 317 37 
<< m2 >>
rect 316 36 317 37 
<< m1 >>
rect 334 36 335 37 
<< m1 >>
rect 337 36 338 37 
<< m1 >>
rect 340 36 341 37 
<< m1 >>
rect 343 36 344 37 
<< m1 >>
rect 19 37 20 38 
<< m1 >>
rect 21 37 22 38 
<< m1 >>
rect 23 37 24 38 
<< m1 >>
rect 37 37 38 38 
<< m1 >>
rect 46 37 47 38 
<< m1 >>
rect 62 37 63 38 
<< m1 >>
rect 64 37 65 38 
<< m1 >>
rect 78 37 79 38 
<< m1 >>
rect 82 37 83 38 
<< m1 >>
rect 92 37 93 38 
<< m1 >>
rect 121 37 122 38 
<< m1 >>
rect 190 37 191 38 
<< m1 >>
rect 200 37 201 38 
<< m2 >>
rect 201 37 202 38 
<< m1 >>
rect 204 37 205 38 
<< m2 >>
rect 204 37 205 38 
<< m2c >>
rect 204 37 205 38 
<< m1 >>
rect 204 37 205 38 
<< m2 >>
rect 204 37 205 38 
<< m2 >>
rect 225 37 226 38 
<< m1 >>
rect 226 37 227 38 
<< m2 >>
rect 226 37 227 38 
<< m2 >>
rect 227 37 228 38 
<< m1 >>
rect 228 37 229 38 
<< m2 >>
rect 228 37 229 38 
<< m2c >>
rect 228 37 229 38 
<< m1 >>
rect 228 37 229 38 
<< m2 >>
rect 228 37 229 38 
<< m1 >>
rect 247 37 248 38 
<< m1 >>
rect 253 37 254 38 
<< m1 >>
rect 265 37 266 38 
<< m1 >>
rect 271 37 272 38 
<< m1 >>
rect 273 37 274 38 
<< m1 >>
rect 275 37 276 38 
<< m1 >>
rect 277 37 278 38 
<< m1 >>
rect 279 37 280 38 
<< m1 >>
rect 289 37 290 38 
<< m1 >>
rect 304 37 305 38 
<< m2 >>
rect 316 37 317 38 
<< m1 >>
rect 334 37 335 38 
<< m1 >>
rect 337 37 338 38 
<< m1 >>
rect 340 37 341 38 
<< m1 >>
rect 343 37 344 38 
<< m1 >>
rect 19 38 20 39 
<< m1 >>
rect 21 38 22 39 
<< m1 >>
rect 23 38 24 39 
<< m1 >>
rect 37 38 38 39 
<< m1 >>
rect 46 38 47 39 
<< m1 >>
rect 62 38 63 39 
<< m2 >>
rect 62 38 63 39 
<< m2c >>
rect 62 38 63 39 
<< m1 >>
rect 62 38 63 39 
<< m2 >>
rect 62 38 63 39 
<< m1 >>
rect 64 38 65 39 
<< m2 >>
rect 64 38 65 39 
<< m2c >>
rect 64 38 65 39 
<< m1 >>
rect 64 38 65 39 
<< m2 >>
rect 64 38 65 39 
<< m1 >>
rect 78 38 79 39 
<< m1 >>
rect 82 38 83 39 
<< m1 >>
rect 92 38 93 39 
<< m1 >>
rect 121 38 122 39 
<< m1 >>
rect 122 38 123 39 
<< m1 >>
rect 123 38 124 39 
<< m1 >>
rect 124 38 125 39 
<< m1 >>
rect 125 38 126 39 
<< m1 >>
rect 126 38 127 39 
<< m1 >>
rect 127 38 128 39 
<< m1 >>
rect 190 38 191 39 
<< m1 >>
rect 200 38 201 39 
<< m2 >>
rect 201 38 202 39 
<< m2 >>
rect 204 38 205 39 
<< m1 >>
rect 226 38 227 39 
<< m1 >>
rect 228 38 229 39 
<< m1 >>
rect 247 38 248 39 
<< m1 >>
rect 248 38 249 39 
<< m1 >>
rect 249 38 250 39 
<< m1 >>
rect 250 38 251 39 
<< m1 >>
rect 251 38 252 39 
<< m1 >>
rect 252 38 253 39 
<< m1 >>
rect 253 38 254 39 
<< m1 >>
rect 265 38 266 39 
<< m1 >>
rect 271 38 272 39 
<< m2 >>
rect 271 38 272 39 
<< m2c >>
rect 271 38 272 39 
<< m1 >>
rect 271 38 272 39 
<< m2 >>
rect 271 38 272 39 
<< m1 >>
rect 273 38 274 39 
<< m2 >>
rect 273 38 274 39 
<< m2c >>
rect 273 38 274 39 
<< m1 >>
rect 273 38 274 39 
<< m2 >>
rect 273 38 274 39 
<< m1 >>
rect 275 38 276 39 
<< m2 >>
rect 275 38 276 39 
<< m2c >>
rect 275 38 276 39 
<< m1 >>
rect 275 38 276 39 
<< m2 >>
rect 275 38 276 39 
<< m1 >>
rect 277 38 278 39 
<< m2 >>
rect 277 38 278 39 
<< m2c >>
rect 277 38 278 39 
<< m1 >>
rect 277 38 278 39 
<< m2 >>
rect 277 38 278 39 
<< m1 >>
rect 279 38 280 39 
<< m2 >>
rect 279 38 280 39 
<< m2c >>
rect 279 38 280 39 
<< m1 >>
rect 279 38 280 39 
<< m2 >>
rect 279 38 280 39 
<< m1 >>
rect 289 38 290 39 
<< m2 >>
rect 289 38 290 39 
<< m2c >>
rect 289 38 290 39 
<< m1 >>
rect 289 38 290 39 
<< m2 >>
rect 289 38 290 39 
<< m1 >>
rect 304 38 305 39 
<< m1 >>
rect 305 38 306 39 
<< m1 >>
rect 306 38 307 39 
<< m1 >>
rect 307 38 308 39 
<< m1 >>
rect 308 38 309 39 
<< m1 >>
rect 309 38 310 39 
<< m1 >>
rect 310 38 311 39 
<< m1 >>
rect 311 38 312 39 
<< m1 >>
rect 312 38 313 39 
<< m1 >>
rect 313 38 314 39 
<< m1 >>
rect 314 38 315 39 
<< m1 >>
rect 315 38 316 39 
<< m1 >>
rect 316 38 317 39 
<< m2 >>
rect 316 38 317 39 
<< m1 >>
rect 317 38 318 39 
<< m1 >>
rect 318 38 319 39 
<< m2 >>
rect 318 38 319 39 
<< m2c >>
rect 318 38 319 39 
<< m1 >>
rect 318 38 319 39 
<< m2 >>
rect 318 38 319 39 
<< m1 >>
rect 334 38 335 39 
<< m2 >>
rect 334 38 335 39 
<< m2c >>
rect 334 38 335 39 
<< m1 >>
rect 334 38 335 39 
<< m2 >>
rect 334 38 335 39 
<< m1 >>
rect 337 38 338 39 
<< m1 >>
rect 338 38 339 39 
<< m2 >>
rect 338 38 339 39 
<< m2c >>
rect 338 38 339 39 
<< m1 >>
rect 338 38 339 39 
<< m2 >>
rect 338 38 339 39 
<< m2 >>
rect 339 38 340 39 
<< m1 >>
rect 340 38 341 39 
<< m2 >>
rect 340 38 341 39 
<< m2 >>
rect 341 38 342 39 
<< m2 >>
rect 342 38 343 39 
<< m1 >>
rect 343 38 344 39 
<< m2 >>
rect 343 38 344 39 
<< m1 >>
rect 19 39 20 40 
<< m1 >>
rect 21 39 22 40 
<< m1 >>
rect 23 39 24 40 
<< m1 >>
rect 37 39 38 40 
<< m1 >>
rect 46 39 47 40 
<< m2 >>
rect 62 39 63 40 
<< m2 >>
rect 64 39 65 40 
<< m1 >>
rect 78 39 79 40 
<< m1 >>
rect 82 39 83 40 
<< m1 >>
rect 92 39 93 40 
<< m1 >>
rect 127 39 128 40 
<< m1 >>
rect 190 39 191 40 
<< m1 >>
rect 200 39 201 40 
<< m2 >>
rect 201 39 202 40 
<< m1 >>
rect 202 39 203 40 
<< m2 >>
rect 202 39 203 40 
<< m2c >>
rect 202 39 203 40 
<< m1 >>
rect 202 39 203 40 
<< m2 >>
rect 202 39 203 40 
<< m1 >>
rect 203 39 204 40 
<< m1 >>
rect 204 39 205 40 
<< m2 >>
rect 204 39 205 40 
<< m1 >>
rect 205 39 206 40 
<< m1 >>
rect 206 39 207 40 
<< m1 >>
rect 207 39 208 40 
<< m1 >>
rect 208 39 209 40 
<< m1 >>
rect 209 39 210 40 
<< m1 >>
rect 210 39 211 40 
<< m2 >>
rect 210 39 211 40 
<< m2c >>
rect 210 39 211 40 
<< m1 >>
rect 210 39 211 40 
<< m2 >>
rect 210 39 211 40 
<< m1 >>
rect 226 39 227 40 
<< m2 >>
rect 226 39 227 40 
<< m2c >>
rect 226 39 227 40 
<< m1 >>
rect 226 39 227 40 
<< m2 >>
rect 226 39 227 40 
<< m1 >>
rect 228 39 229 40 
<< m2 >>
rect 228 39 229 40 
<< m2c >>
rect 228 39 229 40 
<< m1 >>
rect 228 39 229 40 
<< m2 >>
rect 228 39 229 40 
<< m1 >>
rect 265 39 266 40 
<< m2 >>
rect 271 39 272 40 
<< m2 >>
rect 273 39 274 40 
<< m2 >>
rect 275 39 276 40 
<< m2 >>
rect 277 39 278 40 
<< m2 >>
rect 279 39 280 40 
<< m2 >>
rect 289 39 290 40 
<< m2 >>
rect 316 39 317 40 
<< m2 >>
rect 318 39 319 40 
<< m2 >>
rect 334 39 335 40 
<< m1 >>
rect 340 39 341 40 
<< m1 >>
rect 343 39 344 40 
<< m2 >>
rect 343 39 344 40 
<< m1 >>
rect 19 40 20 41 
<< m1 >>
rect 21 40 22 41 
<< m1 >>
rect 23 40 24 41 
<< m1 >>
rect 37 40 38 41 
<< m1 >>
rect 46 40 47 41 
<< m1 >>
rect 55 40 56 41 
<< m1 >>
rect 56 40 57 41 
<< m1 >>
rect 57 40 58 41 
<< m1 >>
rect 58 40 59 41 
<< m1 >>
rect 59 40 60 41 
<< m1 >>
rect 60 40 61 41 
<< m1 >>
rect 61 40 62 41 
<< m1 >>
rect 62 40 63 41 
<< m2 >>
rect 62 40 63 41 
<< m1 >>
rect 63 40 64 41 
<< m1 >>
rect 64 40 65 41 
<< m2 >>
rect 64 40 65 41 
<< m1 >>
rect 65 40 66 41 
<< m1 >>
rect 66 40 67 41 
<< m1 >>
rect 67 40 68 41 
<< m1 >>
rect 68 40 69 41 
<< m1 >>
rect 69 40 70 41 
<< m1 >>
rect 70 40 71 41 
<< m1 >>
rect 71 40 72 41 
<< m1 >>
rect 72 40 73 41 
<< m1 >>
rect 73 40 74 41 
<< m1 >>
rect 74 40 75 41 
<< m1 >>
rect 75 40 76 41 
<< m1 >>
rect 76 40 77 41 
<< m2 >>
rect 76 40 77 41 
<< m2c >>
rect 76 40 77 41 
<< m1 >>
rect 76 40 77 41 
<< m2 >>
rect 76 40 77 41 
<< m2 >>
rect 77 40 78 41 
<< m1 >>
rect 78 40 79 41 
<< m2 >>
rect 78 40 79 41 
<< m2 >>
rect 79 40 80 41 
<< m1 >>
rect 80 40 81 41 
<< m2 >>
rect 80 40 81 41 
<< m2c >>
rect 80 40 81 41 
<< m1 >>
rect 80 40 81 41 
<< m2 >>
rect 80 40 81 41 
<< m2 >>
rect 81 40 82 41 
<< m1 >>
rect 82 40 83 41 
<< m2 >>
rect 82 40 83 41 
<< m2 >>
rect 83 40 84 41 
<< m1 >>
rect 84 40 85 41 
<< m2 >>
rect 84 40 85 41 
<< m2c >>
rect 84 40 85 41 
<< m1 >>
rect 84 40 85 41 
<< m2 >>
rect 84 40 85 41 
<< m1 >>
rect 85 40 86 41 
<< m1 >>
rect 86 40 87 41 
<< m1 >>
rect 87 40 88 41 
<< m1 >>
rect 88 40 89 41 
<< m1 >>
rect 89 40 90 41 
<< m1 >>
rect 90 40 91 41 
<< m1 >>
rect 91 40 92 41 
<< m1 >>
rect 92 40 93 41 
<< m1 >>
rect 127 40 128 41 
<< m1 >>
rect 190 40 191 41 
<< m1 >>
rect 191 40 192 41 
<< m1 >>
rect 192 40 193 41 
<< m1 >>
rect 193 40 194 41 
<< m1 >>
rect 200 40 201 41 
<< m2 >>
rect 204 40 205 41 
<< m2 >>
rect 210 40 211 41 
<< m2 >>
rect 226 40 227 41 
<< m2 >>
rect 228 40 229 41 
<< m2 >>
rect 229 40 230 41 
<< m2 >>
rect 230 40 231 41 
<< m2 >>
rect 231 40 232 41 
<< m2 >>
rect 232 40 233 41 
<< m2 >>
rect 233 40 234 41 
<< m2 >>
rect 234 40 235 41 
<< m2 >>
rect 235 40 236 41 
<< m2 >>
rect 236 40 237 41 
<< m2 >>
rect 237 40 238 41 
<< m2 >>
rect 238 40 239 41 
<< m2 >>
rect 239 40 240 41 
<< m2 >>
rect 240 40 241 41 
<< m2 >>
rect 241 40 242 41 
<< m2 >>
rect 242 40 243 41 
<< m2 >>
rect 243 40 244 41 
<< m2 >>
rect 244 40 245 41 
<< m2 >>
rect 245 40 246 41 
<< m2 >>
rect 246 40 247 41 
<< m2 >>
rect 247 40 248 41 
<< m2 >>
rect 248 40 249 41 
<< m2 >>
rect 249 40 250 41 
<< m2 >>
rect 250 40 251 41 
<< m2 >>
rect 251 40 252 41 
<< m2 >>
rect 252 40 253 41 
<< m2 >>
rect 253 40 254 41 
<< m2 >>
rect 254 40 255 41 
<< m2 >>
rect 255 40 256 41 
<< m2 >>
rect 256 40 257 41 
<< m2 >>
rect 257 40 258 41 
<< m2 >>
rect 258 40 259 41 
<< m2 >>
rect 259 40 260 41 
<< m2 >>
rect 260 40 261 41 
<< m2 >>
rect 261 40 262 41 
<< m2 >>
rect 262 40 263 41 
<< m2 >>
rect 263 40 264 41 
<< m2 >>
rect 264 40 265 41 
<< m1 >>
rect 265 40 266 41 
<< m2 >>
rect 265 40 266 41 
<< m2 >>
rect 266 40 267 41 
<< m1 >>
rect 267 40 268 41 
<< m2 >>
rect 267 40 268 41 
<< m2c >>
rect 267 40 268 41 
<< m1 >>
rect 267 40 268 41 
<< m2 >>
rect 267 40 268 41 
<< m1 >>
rect 268 40 269 41 
<< m1 >>
rect 269 40 270 41 
<< m1 >>
rect 270 40 271 41 
<< m1 >>
rect 271 40 272 41 
<< m2 >>
rect 271 40 272 41 
<< m1 >>
rect 272 40 273 41 
<< m1 >>
rect 273 40 274 41 
<< m2 >>
rect 273 40 274 41 
<< m1 >>
rect 274 40 275 41 
<< m1 >>
rect 275 40 276 41 
<< m2 >>
rect 275 40 276 41 
<< m1 >>
rect 276 40 277 41 
<< m1 >>
rect 277 40 278 41 
<< m2 >>
rect 277 40 278 41 
<< m1 >>
rect 278 40 279 41 
<< m1 >>
rect 279 40 280 41 
<< m2 >>
rect 279 40 280 41 
<< m1 >>
rect 280 40 281 41 
<< m1 >>
rect 281 40 282 41 
<< m1 >>
rect 282 40 283 41 
<< m1 >>
rect 283 40 284 41 
<< m1 >>
rect 284 40 285 41 
<< m1 >>
rect 285 40 286 41 
<< m1 >>
rect 286 40 287 41 
<< m1 >>
rect 287 40 288 41 
<< m1 >>
rect 288 40 289 41 
<< m1 >>
rect 289 40 290 41 
<< m2 >>
rect 289 40 290 41 
<< m1 >>
rect 290 40 291 41 
<< m1 >>
rect 291 40 292 41 
<< m1 >>
rect 292 40 293 41 
<< m1 >>
rect 293 40 294 41 
<< m1 >>
rect 294 40 295 41 
<< m1 >>
rect 295 40 296 41 
<< m1 >>
rect 296 40 297 41 
<< m1 >>
rect 297 40 298 41 
<< m1 >>
rect 298 40 299 41 
<< m1 >>
rect 299 40 300 41 
<< m1 >>
rect 300 40 301 41 
<< m1 >>
rect 301 40 302 41 
<< m1 >>
rect 302 40 303 41 
<< m1 >>
rect 303 40 304 41 
<< m1 >>
rect 304 40 305 41 
<< m1 >>
rect 305 40 306 41 
<< m1 >>
rect 306 40 307 41 
<< m1 >>
rect 307 40 308 41 
<< m1 >>
rect 308 40 309 41 
<< m1 >>
rect 309 40 310 41 
<< m1 >>
rect 310 40 311 41 
<< m1 >>
rect 311 40 312 41 
<< m1 >>
rect 312 40 313 41 
<< m1 >>
rect 313 40 314 41 
<< m1 >>
rect 314 40 315 41 
<< m1 >>
rect 315 40 316 41 
<< m1 >>
rect 316 40 317 41 
<< m2 >>
rect 316 40 317 41 
<< m1 >>
rect 317 40 318 41 
<< m1 >>
rect 318 40 319 41 
<< m2 >>
rect 318 40 319 41 
<< m1 >>
rect 319 40 320 41 
<< m1 >>
rect 334 40 335 41 
<< m2 >>
rect 334 40 335 41 
<< m1 >>
rect 335 40 336 41 
<< m1 >>
rect 336 40 337 41 
<< m1 >>
rect 337 40 338 41 
<< m1 >>
rect 338 40 339 41 
<< m1 >>
rect 339 40 340 41 
<< m1 >>
rect 340 40 341 41 
<< m1 >>
rect 343 40 344 41 
<< m2 >>
rect 343 40 344 41 
<< m1 >>
rect 19 41 20 42 
<< m1 >>
rect 21 41 22 42 
<< m1 >>
rect 23 41 24 42 
<< m1 >>
rect 37 41 38 42 
<< m1 >>
rect 46 41 47 42 
<< m1 >>
rect 55 41 56 42 
<< m2 >>
rect 62 41 63 42 
<< m2 >>
rect 64 41 65 42 
<< m1 >>
rect 78 41 79 42 
<< m1 >>
rect 82 41 83 42 
<< m1 >>
rect 127 41 128 42 
<< m2 >>
rect 189 41 190 42 
<< m2 >>
rect 190 41 191 42 
<< m2 >>
rect 191 41 192 42 
<< m2 >>
rect 192 41 193 42 
<< m1 >>
rect 193 41 194 42 
<< m2 >>
rect 193 41 194 42 
<< m2 >>
rect 194 41 195 42 
<< m1 >>
rect 195 41 196 42 
<< m2 >>
rect 195 41 196 42 
<< m2c >>
rect 195 41 196 42 
<< m1 >>
rect 195 41 196 42 
<< m2 >>
rect 195 41 196 42 
<< m1 >>
rect 196 41 197 42 
<< m1 >>
rect 197 41 198 42 
<< m1 >>
rect 198 41 199 42 
<< m2 >>
rect 198 41 199 42 
<< m2c >>
rect 198 41 199 42 
<< m1 >>
rect 198 41 199 42 
<< m2 >>
rect 198 41 199 42 
<< m2 >>
rect 199 41 200 42 
<< m1 >>
rect 200 41 201 42 
<< m2 >>
rect 200 41 201 42 
<< m2 >>
rect 201 41 202 42 
<< m1 >>
rect 202 41 203 42 
<< m2 >>
rect 202 41 203 42 
<< m2c >>
rect 202 41 203 42 
<< m1 >>
rect 202 41 203 42 
<< m2 >>
rect 202 41 203 42 
<< m1 >>
rect 203 41 204 42 
<< m1 >>
rect 204 41 205 42 
<< m2 >>
rect 204 41 205 42 
<< m1 >>
rect 205 41 206 42 
<< m1 >>
rect 206 41 207 42 
<< m1 >>
rect 207 41 208 42 
<< m1 >>
rect 208 41 209 42 
<< m1 >>
rect 209 41 210 42 
<< m1 >>
rect 210 41 211 42 
<< m2 >>
rect 210 41 211 42 
<< m1 >>
rect 211 41 212 42 
<< m1 >>
rect 212 41 213 42 
<< m1 >>
rect 213 41 214 42 
<< m1 >>
rect 214 41 215 42 
<< m1 >>
rect 215 41 216 42 
<< m1 >>
rect 216 41 217 42 
<< m1 >>
rect 217 41 218 42 
<< m1 >>
rect 218 41 219 42 
<< m1 >>
rect 219 41 220 42 
<< m1 >>
rect 220 41 221 42 
<< m1 >>
rect 221 41 222 42 
<< m1 >>
rect 222 41 223 42 
<< m1 >>
rect 223 41 224 42 
<< m1 >>
rect 224 41 225 42 
<< m1 >>
rect 225 41 226 42 
<< m1 >>
rect 226 41 227 42 
<< m2 >>
rect 226 41 227 42 
<< m1 >>
rect 227 41 228 42 
<< m1 >>
rect 228 41 229 42 
<< m1 >>
rect 229 41 230 42 
<< m1 >>
rect 230 41 231 42 
<< m1 >>
rect 231 41 232 42 
<< m1 >>
rect 232 41 233 42 
<< m1 >>
rect 233 41 234 42 
<< m1 >>
rect 234 41 235 42 
<< m1 >>
rect 235 41 236 42 
<< m1 >>
rect 236 41 237 42 
<< m1 >>
rect 237 41 238 42 
<< m1 >>
rect 238 41 239 42 
<< m1 >>
rect 239 41 240 42 
<< m1 >>
rect 240 41 241 42 
<< m1 >>
rect 241 41 242 42 
<< m1 >>
rect 242 41 243 42 
<< m1 >>
rect 243 41 244 42 
<< m1 >>
rect 244 41 245 42 
<< m1 >>
rect 245 41 246 42 
<< m1 >>
rect 246 41 247 42 
<< m1 >>
rect 247 41 248 42 
<< m1 >>
rect 248 41 249 42 
<< m1 >>
rect 249 41 250 42 
<< m1 >>
rect 250 41 251 42 
<< m1 >>
rect 251 41 252 42 
<< m1 >>
rect 252 41 253 42 
<< m1 >>
rect 253 41 254 42 
<< m1 >>
rect 254 41 255 42 
<< m1 >>
rect 255 41 256 42 
<< m1 >>
rect 256 41 257 42 
<< m1 >>
rect 257 41 258 42 
<< m1 >>
rect 258 41 259 42 
<< m1 >>
rect 259 41 260 42 
<< m1 >>
rect 260 41 261 42 
<< m1 >>
rect 261 41 262 42 
<< m1 >>
rect 262 41 263 42 
<< m1 >>
rect 263 41 264 42 
<< m1 >>
rect 264 41 265 42 
<< m1 >>
rect 265 41 266 42 
<< m2 >>
rect 271 41 272 42 
<< m2 >>
rect 273 41 274 42 
<< m2 >>
rect 275 41 276 42 
<< m2 >>
rect 277 41 278 42 
<< m2 >>
rect 279 41 280 42 
<< m2 >>
rect 289 41 290 42 
<< m2 >>
rect 316 41 317 42 
<< m2 >>
rect 318 41 319 42 
<< m1 >>
rect 319 41 320 42 
<< m1 >>
rect 334 41 335 42 
<< m2 >>
rect 334 41 335 42 
<< m1 >>
rect 343 41 344 42 
<< m2 >>
rect 343 41 344 42 
<< m1 >>
rect 19 42 20 43 
<< m1 >>
rect 21 42 22 43 
<< m1 >>
rect 23 42 24 43 
<< m1 >>
rect 37 42 38 43 
<< m1 >>
rect 46 42 47 43 
<< m1 >>
rect 55 42 56 43 
<< m1 >>
rect 60 42 61 43 
<< m1 >>
rect 61 42 62 43 
<< m1 >>
rect 62 42 63 43 
<< m2 >>
rect 62 42 63 43 
<< m1 >>
rect 63 42 64 43 
<< m1 >>
rect 64 42 65 43 
<< m2 >>
rect 64 42 65 43 
<< m2c >>
rect 64 42 65 43 
<< m1 >>
rect 64 42 65 43 
<< m2 >>
rect 64 42 65 43 
<< m1 >>
rect 78 42 79 43 
<< m2 >>
rect 78 42 79 43 
<< m2c >>
rect 78 42 79 43 
<< m1 >>
rect 78 42 79 43 
<< m2 >>
rect 78 42 79 43 
<< m1 >>
rect 82 42 83 43 
<< m1 >>
rect 127 42 128 43 
<< m2 >>
rect 189 42 190 43 
<< m1 >>
rect 193 42 194 43 
<< m1 >>
rect 200 42 201 43 
<< m2 >>
rect 204 42 205 43 
<< m2 >>
rect 210 42 211 43 
<< m2 >>
rect 211 42 212 43 
<< m2 >>
rect 212 42 213 43 
<< m2 >>
rect 213 42 214 43 
<< m2 >>
rect 214 42 215 43 
<< m2 >>
rect 215 42 216 43 
<< m2 >>
rect 216 42 217 43 
<< m2 >>
rect 217 42 218 43 
<< m2 >>
rect 218 42 219 43 
<< m2 >>
rect 219 42 220 43 
<< m2 >>
rect 220 42 221 43 
<< m2 >>
rect 226 42 227 43 
<< m1 >>
rect 271 42 272 43 
<< m2 >>
rect 271 42 272 43 
<< m2c >>
rect 271 42 272 43 
<< m1 >>
rect 271 42 272 43 
<< m2 >>
rect 271 42 272 43 
<< m1 >>
rect 273 42 274 43 
<< m2 >>
rect 273 42 274 43 
<< m2c >>
rect 273 42 274 43 
<< m1 >>
rect 273 42 274 43 
<< m2 >>
rect 273 42 274 43 
<< m1 >>
rect 275 42 276 43 
<< m2 >>
rect 275 42 276 43 
<< m2c >>
rect 275 42 276 43 
<< m1 >>
rect 275 42 276 43 
<< m2 >>
rect 275 42 276 43 
<< m1 >>
rect 277 42 278 43 
<< m2 >>
rect 277 42 278 43 
<< m2c >>
rect 277 42 278 43 
<< m1 >>
rect 277 42 278 43 
<< m2 >>
rect 277 42 278 43 
<< m1 >>
rect 279 42 280 43 
<< m2 >>
rect 279 42 280 43 
<< m2c >>
rect 279 42 280 43 
<< m1 >>
rect 279 42 280 43 
<< m2 >>
rect 279 42 280 43 
<< m1 >>
rect 280 42 281 43 
<< m1 >>
rect 289 42 290 43 
<< m2 >>
rect 289 42 290 43 
<< m2c >>
rect 289 42 290 43 
<< m1 >>
rect 289 42 290 43 
<< m2 >>
rect 289 42 290 43 
<< m1 >>
rect 316 42 317 43 
<< m2 >>
rect 316 42 317 43 
<< m2c >>
rect 316 42 317 43 
<< m1 >>
rect 316 42 317 43 
<< m2 >>
rect 316 42 317 43 
<< m2 >>
rect 318 42 319 43 
<< m1 >>
rect 319 42 320 43 
<< m1 >>
rect 334 42 335 43 
<< m2 >>
rect 334 42 335 43 
<< m1 >>
rect 337 42 338 43 
<< m1 >>
rect 338 42 339 43 
<< m1 >>
rect 339 42 340 43 
<< m1 >>
rect 340 42 341 43 
<< m1 >>
rect 341 42 342 43 
<< m1 >>
rect 342 42 343 43 
<< m1 >>
rect 343 42 344 43 
<< m2 >>
rect 343 42 344 43 
<< m1 >>
rect 19 43 20 44 
<< m1 >>
rect 21 43 22 44 
<< m1 >>
rect 23 43 24 44 
<< m1 >>
rect 37 43 38 44 
<< m1 >>
rect 46 43 47 44 
<< m1 >>
rect 55 43 56 44 
<< m1 >>
rect 60 43 61 44 
<< m2 >>
rect 62 43 63 44 
<< m1 >>
rect 66 43 67 44 
<< m2 >>
rect 66 43 67 44 
<< m1 >>
rect 67 43 68 44 
<< m2 >>
rect 67 43 68 44 
<< m1 >>
rect 68 43 69 44 
<< m2 >>
rect 68 43 69 44 
<< m1 >>
rect 69 43 70 44 
<< m2 >>
rect 69 43 70 44 
<< m1 >>
rect 70 43 71 44 
<< m2 >>
rect 70 43 71 44 
<< m1 >>
rect 71 43 72 44 
<< m2 >>
rect 71 43 72 44 
<< m2 >>
rect 72 43 73 44 
<< m2 >>
rect 73 43 74 44 
<< m2 >>
rect 74 43 75 44 
<< m2 >>
rect 75 43 76 44 
<< m2 >>
rect 78 43 79 44 
<< m2 >>
rect 81 43 82 44 
<< m1 >>
rect 82 43 83 44 
<< m2 >>
rect 82 43 83 44 
<< m2 >>
rect 83 43 84 44 
<< m1 >>
rect 84 43 85 44 
<< m2 >>
rect 84 43 85 44 
<< m1 >>
rect 85 43 86 44 
<< m2 >>
rect 85 43 86 44 
<< m1 >>
rect 86 43 87 44 
<< m2 >>
rect 86 43 87 44 
<< m1 >>
rect 87 43 88 44 
<< m2 >>
rect 87 43 88 44 
<< m1 >>
rect 88 43 89 44 
<< m1 >>
rect 89 43 90 44 
<< m1 >>
rect 90 43 91 44 
<< m1 >>
rect 91 43 92 44 
<< m1 >>
rect 92 43 93 44 
<< m1 >>
rect 93 43 94 44 
<< m1 >>
rect 94 43 95 44 
<< m1 >>
rect 95 43 96 44 
<< m1 >>
rect 96 43 97 44 
<< m1 >>
rect 97 43 98 44 
<< m1 >>
rect 98 43 99 44 
<< m1 >>
rect 99 43 100 44 
<< m1 >>
rect 100 43 101 44 
<< m1 >>
rect 101 43 102 44 
<< m1 >>
rect 102 43 103 44 
<< m1 >>
rect 103 43 104 44 
<< m1 >>
rect 104 43 105 44 
<< m1 >>
rect 105 43 106 44 
<< m1 >>
rect 106 43 107 44 
<< m1 >>
rect 107 43 108 44 
<< m1 >>
rect 108 43 109 44 
<< m1 >>
rect 109 43 110 44 
<< m1 >>
rect 110 43 111 44 
<< m1 >>
rect 111 43 112 44 
<< m1 >>
rect 112 43 113 44 
<< m1 >>
rect 113 43 114 44 
<< m1 >>
rect 114 43 115 44 
<< m1 >>
rect 115 43 116 44 
<< m1 >>
rect 116 43 117 44 
<< m1 >>
rect 117 43 118 44 
<< m1 >>
rect 118 43 119 44 
<< m1 >>
rect 119 43 120 44 
<< m1 >>
rect 120 43 121 44 
<< m1 >>
rect 121 43 122 44 
<< m1 >>
rect 122 43 123 44 
<< m1 >>
rect 123 43 124 44 
<< m1 >>
rect 124 43 125 44 
<< m1 >>
rect 125 43 126 44 
<< m2 >>
rect 125 43 126 44 
<< m2c >>
rect 125 43 126 44 
<< m1 >>
rect 125 43 126 44 
<< m2 >>
rect 125 43 126 44 
<< m2 >>
rect 126 43 127 44 
<< m1 >>
rect 127 43 128 44 
<< m2 >>
rect 127 43 128 44 
<< m2 >>
rect 128 43 129 44 
<< m1 >>
rect 129 43 130 44 
<< m2 >>
rect 129 43 130 44 
<< m2c >>
rect 129 43 130 44 
<< m1 >>
rect 129 43 130 44 
<< m2 >>
rect 129 43 130 44 
<< m1 >>
rect 130 43 131 44 
<< m1 >>
rect 131 43 132 44 
<< m1 >>
rect 132 43 133 44 
<< m1 >>
rect 133 43 134 44 
<< m1 >>
rect 134 43 135 44 
<< m1 >>
rect 135 43 136 44 
<< m1 >>
rect 136 43 137 44 
<< m1 >>
rect 137 43 138 44 
<< m2 >>
rect 137 43 138 44 
<< m2c >>
rect 137 43 138 44 
<< m1 >>
rect 137 43 138 44 
<< m2 >>
rect 137 43 138 44 
<< m2 >>
rect 138 43 139 44 
<< m1 >>
rect 139 43 140 44 
<< m2 >>
rect 139 43 140 44 
<< m1 >>
rect 140 43 141 44 
<< m2 >>
rect 140 43 141 44 
<< m1 >>
rect 141 43 142 44 
<< m2 >>
rect 141 43 142 44 
<< m1 >>
rect 142 43 143 44 
<< m2 >>
rect 142 43 143 44 
<< m1 >>
rect 143 43 144 44 
<< m2 >>
rect 143 43 144 44 
<< m1 >>
rect 144 43 145 44 
<< m2 >>
rect 144 43 145 44 
<< m1 >>
rect 145 43 146 44 
<< m2 >>
rect 145 43 146 44 
<< m1 >>
rect 146 43 147 44 
<< m2 >>
rect 146 43 147 44 
<< m1 >>
rect 147 43 148 44 
<< m2 >>
rect 147 43 148 44 
<< m1 >>
rect 148 43 149 44 
<< m2 >>
rect 148 43 149 44 
<< m1 >>
rect 149 43 150 44 
<< m2 >>
rect 149 43 150 44 
<< m1 >>
rect 150 43 151 44 
<< m2 >>
rect 150 43 151 44 
<< m1 >>
rect 151 43 152 44 
<< m2 >>
rect 151 43 152 44 
<< m1 >>
rect 152 43 153 44 
<< m2 >>
rect 152 43 153 44 
<< m1 >>
rect 153 43 154 44 
<< m2 >>
rect 153 43 154 44 
<< m1 >>
rect 154 43 155 44 
<< m2 >>
rect 154 43 155 44 
<< m1 >>
rect 155 43 156 44 
<< m2 >>
rect 155 43 156 44 
<< m1 >>
rect 156 43 157 44 
<< m2 >>
rect 156 43 157 44 
<< m1 >>
rect 157 43 158 44 
<< m2 >>
rect 157 43 158 44 
<< m1 >>
rect 158 43 159 44 
<< m2 >>
rect 158 43 159 44 
<< m1 >>
rect 159 43 160 44 
<< m2 >>
rect 159 43 160 44 
<< m1 >>
rect 160 43 161 44 
<< m2 >>
rect 160 43 161 44 
<< m1 >>
rect 161 43 162 44 
<< m2 >>
rect 161 43 162 44 
<< m1 >>
rect 162 43 163 44 
<< m2 >>
rect 162 43 163 44 
<< m1 >>
rect 163 43 164 44 
<< m2 >>
rect 163 43 164 44 
<< m1 >>
rect 164 43 165 44 
<< m2 >>
rect 164 43 165 44 
<< m1 >>
rect 165 43 166 44 
<< m2 >>
rect 165 43 166 44 
<< m1 >>
rect 166 43 167 44 
<< m2 >>
rect 166 43 167 44 
<< m1 >>
rect 167 43 168 44 
<< m2 >>
rect 167 43 168 44 
<< m1 >>
rect 168 43 169 44 
<< m2 >>
rect 168 43 169 44 
<< m1 >>
rect 169 43 170 44 
<< m2 >>
rect 169 43 170 44 
<< m1 >>
rect 170 43 171 44 
<< m2 >>
rect 170 43 171 44 
<< m1 >>
rect 171 43 172 44 
<< m2 >>
rect 171 43 172 44 
<< m1 >>
rect 172 43 173 44 
<< m2 >>
rect 172 43 173 44 
<< m1 >>
rect 173 43 174 44 
<< m2 >>
rect 173 43 174 44 
<< m1 >>
rect 174 43 175 44 
<< m2 >>
rect 174 43 175 44 
<< m1 >>
rect 175 43 176 44 
<< m2 >>
rect 175 43 176 44 
<< m1 >>
rect 176 43 177 44 
<< m2 >>
rect 176 43 177 44 
<< m1 >>
rect 177 43 178 44 
<< m2 >>
rect 177 43 178 44 
<< m1 >>
rect 178 43 179 44 
<< m2 >>
rect 178 43 179 44 
<< m1 >>
rect 179 43 180 44 
<< m2 >>
rect 179 43 180 44 
<< m1 >>
rect 180 43 181 44 
<< m2 >>
rect 180 43 181 44 
<< m1 >>
rect 181 43 182 44 
<< m2 >>
rect 181 43 182 44 
<< m1 >>
rect 182 43 183 44 
<< m2 >>
rect 182 43 183 44 
<< m1 >>
rect 183 43 184 44 
<< m2 >>
rect 183 43 184 44 
<< m1 >>
rect 184 43 185 44 
<< m2 >>
rect 184 43 185 44 
<< m1 >>
rect 185 43 186 44 
<< m2 >>
rect 185 43 186 44 
<< m1 >>
rect 186 43 187 44 
<< m2 >>
rect 186 43 187 44 
<< m1 >>
rect 187 43 188 44 
<< m2 >>
rect 187 43 188 44 
<< m1 >>
rect 188 43 189 44 
<< m2 >>
rect 188 43 189 44 
<< m1 >>
rect 189 43 190 44 
<< m2 >>
rect 189 43 190 44 
<< m1 >>
rect 190 43 191 44 
<< m1 >>
rect 191 43 192 44 
<< m2 >>
rect 191 43 192 44 
<< m2c >>
rect 191 43 192 44 
<< m1 >>
rect 191 43 192 44 
<< m2 >>
rect 191 43 192 44 
<< m2 >>
rect 192 43 193 44 
<< m1 >>
rect 193 43 194 44 
<< m2 >>
rect 193 43 194 44 
<< m2 >>
rect 194 43 195 44 
<< m1 >>
rect 200 43 201 44 
<< m1 >>
rect 204 43 205 44 
<< m2 >>
rect 204 43 205 44 
<< m2c >>
rect 204 43 205 44 
<< m1 >>
rect 204 43 205 44 
<< m2 >>
rect 204 43 205 44 
<< m1 >>
rect 220 43 221 44 
<< m2 >>
rect 220 43 221 44 
<< m2c >>
rect 220 43 221 44 
<< m1 >>
rect 220 43 221 44 
<< m2 >>
rect 220 43 221 44 
<< m1 >>
rect 226 43 227 44 
<< m2 >>
rect 226 43 227 44 
<< m2c >>
rect 226 43 227 44 
<< m1 >>
rect 226 43 227 44 
<< m2 >>
rect 226 43 227 44 
<< m1 >>
rect 271 43 272 44 
<< m1 >>
rect 273 43 274 44 
<< m1 >>
rect 275 43 276 44 
<< m1 >>
rect 277 43 278 44 
<< m1 >>
rect 280 43 281 44 
<< m1 >>
rect 289 43 290 44 
<< m1 >>
rect 316 43 317 44 
<< m2 >>
rect 318 43 319 44 
<< m1 >>
rect 319 43 320 44 
<< m2 >>
rect 319 43 320 44 
<< m2 >>
rect 320 43 321 44 
<< m1 >>
rect 334 43 335 44 
<< m2 >>
rect 334 43 335 44 
<< m1 >>
rect 337 43 338 44 
<< m2 >>
rect 343 43 344 44 
<< m1 >>
rect 19 44 20 45 
<< m1 >>
rect 21 44 22 45 
<< m1 >>
rect 23 44 24 45 
<< m1 >>
rect 37 44 38 45 
<< m1 >>
rect 46 44 47 45 
<< m1 >>
rect 55 44 56 45 
<< m1 >>
rect 60 44 61 45 
<< m1 >>
rect 62 44 63 45 
<< m2 >>
rect 62 44 63 45 
<< m2c >>
rect 62 44 63 45 
<< m1 >>
rect 62 44 63 45 
<< m2 >>
rect 62 44 63 45 
<< m1 >>
rect 63 44 64 45 
<< m1 >>
rect 64 44 65 45 
<< m1 >>
rect 65 44 66 45 
<< m1 >>
rect 66 44 67 45 
<< m2 >>
rect 66 44 67 45 
<< m1 >>
rect 71 44 72 45 
<< m1 >>
rect 73 44 74 45 
<< m1 >>
rect 74 44 75 45 
<< m1 >>
rect 75 44 76 45 
<< m2 >>
rect 75 44 76 45 
<< m1 >>
rect 76 44 77 45 
<< m1 >>
rect 77 44 78 45 
<< m1 >>
rect 78 44 79 45 
<< m2 >>
rect 78 44 79 45 
<< m1 >>
rect 79 44 80 45 
<< m1 >>
rect 80 44 81 45 
<< m2 >>
rect 80 44 81 45 
<< m2c >>
rect 80 44 81 45 
<< m1 >>
rect 80 44 81 45 
<< m2 >>
rect 80 44 81 45 
<< m2 >>
rect 81 44 82 45 
<< m1 >>
rect 82 44 83 45 
<< m1 >>
rect 84 44 85 45 
<< m2 >>
rect 87 44 88 45 
<< m1 >>
rect 127 44 128 45 
<< m1 >>
rect 139 44 140 45 
<< m1 >>
rect 193 44 194 45 
<< m2 >>
rect 194 44 195 45 
<< m1 >>
rect 200 44 201 45 
<< m1 >>
rect 204 44 205 45 
<< m1 >>
rect 220 44 221 45 
<< m1 >>
rect 226 44 227 45 
<< m1 >>
rect 271 44 272 45 
<< m1 >>
rect 273 44 274 45 
<< m2 >>
rect 274 44 275 45 
<< m1 >>
rect 275 44 276 45 
<< m2 >>
rect 275 44 276 45 
<< m2c >>
rect 275 44 276 45 
<< m1 >>
rect 275 44 276 45 
<< m2 >>
rect 275 44 276 45 
<< m1 >>
rect 277 44 278 45 
<< m1 >>
rect 280 44 281 45 
<< m1 >>
rect 289 44 290 45 
<< m1 >>
rect 316 44 317 45 
<< m1 >>
rect 319 44 320 45 
<< m2 >>
rect 320 44 321 45 
<< m1 >>
rect 334 44 335 45 
<< m2 >>
rect 334 44 335 45 
<< m1 >>
rect 337 44 338 45 
<< m1 >>
rect 343 44 344 45 
<< m2 >>
rect 343 44 344 45 
<< m2c >>
rect 343 44 344 45 
<< m1 >>
rect 343 44 344 45 
<< m2 >>
rect 343 44 344 45 
<< m1 >>
rect 19 45 20 46 
<< m1 >>
rect 21 45 22 46 
<< m1 >>
rect 23 45 24 46 
<< m1 >>
rect 37 45 38 46 
<< m1 >>
rect 46 45 47 46 
<< m1 >>
rect 55 45 56 46 
<< m1 >>
rect 60 45 61 46 
<< m2 >>
rect 66 45 67 46 
<< m1 >>
rect 71 45 72 46 
<< m1 >>
rect 73 45 74 46 
<< m2 >>
rect 75 45 76 46 
<< m2 >>
rect 78 45 79 46 
<< m1 >>
rect 82 45 83 46 
<< m1 >>
rect 84 45 85 46 
<< m2 >>
rect 87 45 88 46 
<< m2 >>
rect 88 45 89 46 
<< m2 >>
rect 89 45 90 46 
<< m2 >>
rect 90 45 91 46 
<< m2 >>
rect 91 45 92 46 
<< m2 >>
rect 92 45 93 46 
<< m1 >>
rect 93 45 94 46 
<< m2 >>
rect 93 45 94 46 
<< m2c >>
rect 93 45 94 46 
<< m1 >>
rect 93 45 94 46 
<< m2 >>
rect 93 45 94 46 
<< m1 >>
rect 94 45 95 46 
<< m1 >>
rect 95 45 96 46 
<< m1 >>
rect 96 45 97 46 
<< m1 >>
rect 97 45 98 46 
<< m1 >>
rect 127 45 128 46 
<< m1 >>
rect 139 45 140 46 
<< m1 >>
rect 193 45 194 46 
<< m2 >>
rect 194 45 195 46 
<< m1 >>
rect 195 45 196 46 
<< m2 >>
rect 195 45 196 46 
<< m2c >>
rect 195 45 196 46 
<< m1 >>
rect 195 45 196 46 
<< m2 >>
rect 195 45 196 46 
<< m1 >>
rect 196 45 197 46 
<< m1 >>
rect 197 45 198 46 
<< m1 >>
rect 198 45 199 46 
<< m1 >>
rect 200 45 201 46 
<< m1 >>
rect 204 45 205 46 
<< m1 >>
rect 220 45 221 46 
<< m1 >>
rect 226 45 227 46 
<< m1 >>
rect 271 45 272 46 
<< m1 >>
rect 273 45 274 46 
<< m2 >>
rect 274 45 275 46 
<< m1 >>
rect 277 45 278 46 
<< m1 >>
rect 280 45 281 46 
<< m1 >>
rect 289 45 290 46 
<< m1 >>
rect 316 45 317 46 
<< m1 >>
rect 319 45 320 46 
<< m2 >>
rect 320 45 321 46 
<< m1 >>
rect 321 45 322 46 
<< m2 >>
rect 321 45 322 46 
<< m2c >>
rect 321 45 322 46 
<< m1 >>
rect 321 45 322 46 
<< m2 >>
rect 321 45 322 46 
<< m1 >>
rect 322 45 323 46 
<< m1 >>
rect 323 45 324 46 
<< m1 >>
rect 324 45 325 46 
<< m1 >>
rect 325 45 326 46 
<< m1 >>
rect 326 45 327 46 
<< m1 >>
rect 327 45 328 46 
<< m1 >>
rect 334 45 335 46 
<< m2 >>
rect 334 45 335 46 
<< m1 >>
rect 337 45 338 46 
<< m1 >>
rect 343 45 344 46 
<< m1 >>
rect 19 46 20 47 
<< m1 >>
rect 21 46 22 47 
<< m1 >>
rect 23 46 24 47 
<< m1 >>
rect 37 46 38 47 
<< m1 >>
rect 46 46 47 47 
<< m1 >>
rect 55 46 56 47 
<< m2 >>
rect 56 46 57 47 
<< m1 >>
rect 57 46 58 47 
<< m2 >>
rect 57 46 58 47 
<< m1 >>
rect 58 46 59 47 
<< m2 >>
rect 58 46 59 47 
<< m2c >>
rect 58 46 59 47 
<< m1 >>
rect 58 46 59 47 
<< m2 >>
rect 58 46 59 47 
<< m2 >>
rect 59 46 60 47 
<< m1 >>
rect 60 46 61 47 
<< m2 >>
rect 60 46 61 47 
<< m2 >>
rect 61 46 62 47 
<< m1 >>
rect 62 46 63 47 
<< m2 >>
rect 62 46 63 47 
<< m2c >>
rect 62 46 63 47 
<< m1 >>
rect 62 46 63 47 
<< m2 >>
rect 62 46 63 47 
<< m1 >>
rect 63 46 64 47 
<< m1 >>
rect 64 46 65 47 
<< m1 >>
rect 65 46 66 47 
<< m1 >>
rect 66 46 67 47 
<< m2 >>
rect 66 46 67 47 
<< m2c >>
rect 66 46 67 47 
<< m1 >>
rect 66 46 67 47 
<< m2 >>
rect 66 46 67 47 
<< m1 >>
rect 71 46 72 47 
<< m2 >>
rect 71 46 72 47 
<< m2c >>
rect 71 46 72 47 
<< m1 >>
rect 71 46 72 47 
<< m2 >>
rect 71 46 72 47 
<< m2 >>
rect 72 46 73 47 
<< m1 >>
rect 73 46 74 47 
<< m2 >>
rect 73 46 74 47 
<< m1 >>
rect 75 46 76 47 
<< m2 >>
rect 75 46 76 47 
<< m2c >>
rect 75 46 76 47 
<< m1 >>
rect 75 46 76 47 
<< m2 >>
rect 75 46 76 47 
<< m1 >>
rect 78 46 79 47 
<< m2 >>
rect 78 46 79 47 
<< m2c >>
rect 78 46 79 47 
<< m1 >>
rect 78 46 79 47 
<< m2 >>
rect 78 46 79 47 
<< m2 >>
rect 81 46 82 47 
<< m1 >>
rect 82 46 83 47 
<< m2 >>
rect 82 46 83 47 
<< m2 >>
rect 83 46 84 47 
<< m1 >>
rect 84 46 85 47 
<< m2 >>
rect 84 46 85 47 
<< m2c >>
rect 84 46 85 47 
<< m1 >>
rect 84 46 85 47 
<< m2 >>
rect 84 46 85 47 
<< m1 >>
rect 88 46 89 47 
<< m1 >>
rect 89 46 90 47 
<< m1 >>
rect 90 46 91 47 
<< m1 >>
rect 91 46 92 47 
<< m1 >>
rect 97 46 98 47 
<< m1 >>
rect 127 46 128 47 
<< m1 >>
rect 139 46 140 47 
<< m1 >>
rect 193 46 194 47 
<< m1 >>
rect 198 46 199 47 
<< m2 >>
rect 198 46 199 47 
<< m2c >>
rect 198 46 199 47 
<< m1 >>
rect 198 46 199 47 
<< m2 >>
rect 198 46 199 47 
<< m2 >>
rect 199 46 200 47 
<< m1 >>
rect 200 46 201 47 
<< m2 >>
rect 200 46 201 47 
<< m2 >>
rect 201 46 202 47 
<< m1 >>
rect 204 46 205 47 
<< m1 >>
rect 220 46 221 47 
<< m1 >>
rect 226 46 227 47 
<< m1 >>
rect 250 46 251 47 
<< m1 >>
rect 251 46 252 47 
<< m1 >>
rect 252 46 253 47 
<< m1 >>
rect 253 46 254 47 
<< m1 >>
rect 254 46 255 47 
<< m1 >>
rect 255 46 256 47 
<< m1 >>
rect 256 46 257 47 
<< m1 >>
rect 257 46 258 47 
<< m1 >>
rect 258 46 259 47 
<< m1 >>
rect 259 46 260 47 
<< m1 >>
rect 260 46 261 47 
<< m1 >>
rect 261 46 262 47 
<< m1 >>
rect 262 46 263 47 
<< m1 >>
rect 271 46 272 47 
<< m1 >>
rect 273 46 274 47 
<< m2 >>
rect 274 46 275 47 
<< m1 >>
rect 277 46 278 47 
<< m1 >>
rect 280 46 281 47 
<< m1 >>
rect 289 46 290 47 
<< m1 >>
rect 304 46 305 47 
<< m1 >>
rect 305 46 306 47 
<< m1 >>
rect 306 46 307 47 
<< m1 >>
rect 307 46 308 47 
<< m1 >>
rect 316 46 317 47 
<< m1 >>
rect 319 46 320 47 
<< m1 >>
rect 327 46 328 47 
<< m1 >>
rect 334 46 335 47 
<< m2 >>
rect 334 46 335 47 
<< m1 >>
rect 337 46 338 47 
<< m1 >>
rect 343 46 344 47 
<< m1 >>
rect 19 47 20 48 
<< m1 >>
rect 21 47 22 48 
<< m1 >>
rect 23 47 24 48 
<< m1 >>
rect 37 47 38 48 
<< m1 >>
rect 46 47 47 48 
<< m1 >>
rect 55 47 56 48 
<< m2 >>
rect 56 47 57 48 
<< m1 >>
rect 60 47 61 48 
<< m1 >>
rect 73 47 74 48 
<< m2 >>
rect 73 47 74 48 
<< m1 >>
rect 75 47 76 48 
<< m1 >>
rect 78 47 79 48 
<< m2 >>
rect 81 47 82 48 
<< m1 >>
rect 82 47 83 48 
<< m1 >>
rect 88 47 89 48 
<< m1 >>
rect 91 47 92 48 
<< m1 >>
rect 97 47 98 48 
<< m1 >>
rect 127 47 128 48 
<< m1 >>
rect 139 47 140 48 
<< m1 >>
rect 193 47 194 48 
<< m1 >>
rect 200 47 201 48 
<< m2 >>
rect 201 47 202 48 
<< m1 >>
rect 204 47 205 48 
<< m1 >>
rect 220 47 221 48 
<< m1 >>
rect 226 47 227 48 
<< m1 >>
rect 250 47 251 48 
<< m1 >>
rect 262 47 263 48 
<< m1 >>
rect 271 47 272 48 
<< m1 >>
rect 273 47 274 48 
<< m2 >>
rect 274 47 275 48 
<< m1 >>
rect 277 47 278 48 
<< m1 >>
rect 280 47 281 48 
<< m1 >>
rect 289 47 290 48 
<< m1 >>
rect 304 47 305 48 
<< m1 >>
rect 307 47 308 48 
<< m1 >>
rect 316 47 317 48 
<< m1 >>
rect 319 47 320 48 
<< m1 >>
rect 327 47 328 48 
<< m1 >>
rect 334 47 335 48 
<< m2 >>
rect 334 47 335 48 
<< m1 >>
rect 337 47 338 48 
<< m1 >>
rect 343 47 344 48 
<< pdiffusion >>
rect 12 48 13 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< m1 >>
rect 19 48 20 49 
<< m1 >>
rect 21 48 22 49 
<< m1 >>
rect 23 48 24 49 
<< pdiffusion >>
rect 30 48 31 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< m1 >>
rect 37 48 38 49 
<< m1 >>
rect 46 48 47 49 
<< pdiffusion >>
rect 48 48 49 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 55 48 56 49 
<< m2 >>
rect 56 48 57 49 
<< m1 >>
rect 60 48 61 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< m1 >>
rect 73 48 74 49 
<< m2 >>
rect 73 48 74 49 
<< m1 >>
rect 75 48 76 49 
<< m1 >>
rect 78 48 79 49 
<< m2 >>
rect 81 48 82 49 
<< m1 >>
rect 82 48 83 49 
<< pdiffusion >>
rect 84 48 85 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< m1 >>
rect 88 48 89 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< m1 >>
rect 97 48 98 49 
<< pdiffusion >>
rect 102 48 103 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< pdiffusion >>
rect 120 48 121 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< m1 >>
rect 127 48 128 49 
<< pdiffusion >>
rect 138 48 139 49 
<< m1 >>
rect 139 48 140 49 
<< pdiffusion >>
rect 139 48 140 49 
<< pdiffusion >>
rect 140 48 141 49 
<< pdiffusion >>
rect 141 48 142 49 
<< pdiffusion >>
rect 142 48 143 49 
<< pdiffusion >>
rect 143 48 144 49 
<< pdiffusion >>
rect 156 48 157 49 
<< pdiffusion >>
rect 157 48 158 49 
<< pdiffusion >>
rect 158 48 159 49 
<< pdiffusion >>
rect 159 48 160 49 
<< pdiffusion >>
rect 160 48 161 49 
<< pdiffusion >>
rect 161 48 162 49 
<< pdiffusion >>
rect 174 48 175 49 
<< pdiffusion >>
rect 175 48 176 49 
<< pdiffusion >>
rect 176 48 177 49 
<< pdiffusion >>
rect 177 48 178 49 
<< pdiffusion >>
rect 178 48 179 49 
<< pdiffusion >>
rect 179 48 180 49 
<< pdiffusion >>
rect 192 48 193 49 
<< m1 >>
rect 193 48 194 49 
<< pdiffusion >>
rect 193 48 194 49 
<< pdiffusion >>
rect 194 48 195 49 
<< pdiffusion >>
rect 195 48 196 49 
<< pdiffusion >>
rect 196 48 197 49 
<< pdiffusion >>
rect 197 48 198 49 
<< m1 >>
rect 200 48 201 49 
<< m2 >>
rect 201 48 202 49 
<< m1 >>
rect 204 48 205 49 
<< pdiffusion >>
rect 210 48 211 49 
<< pdiffusion >>
rect 211 48 212 49 
<< pdiffusion >>
rect 212 48 213 49 
<< pdiffusion >>
rect 213 48 214 49 
<< pdiffusion >>
rect 214 48 215 49 
<< pdiffusion >>
rect 215 48 216 49 
<< m1 >>
rect 220 48 221 49 
<< m1 >>
rect 226 48 227 49 
<< pdiffusion >>
rect 228 48 229 49 
<< pdiffusion >>
rect 229 48 230 49 
<< pdiffusion >>
rect 230 48 231 49 
<< pdiffusion >>
rect 231 48 232 49 
<< pdiffusion >>
rect 232 48 233 49 
<< pdiffusion >>
rect 233 48 234 49 
<< pdiffusion >>
rect 246 48 247 49 
<< pdiffusion >>
rect 247 48 248 49 
<< pdiffusion >>
rect 248 48 249 49 
<< pdiffusion >>
rect 249 48 250 49 
<< m1 >>
rect 250 48 251 49 
<< pdiffusion >>
rect 250 48 251 49 
<< pdiffusion >>
rect 251 48 252 49 
<< m1 >>
rect 262 48 263 49 
<< pdiffusion >>
rect 264 48 265 49 
<< pdiffusion >>
rect 265 48 266 49 
<< pdiffusion >>
rect 266 48 267 49 
<< pdiffusion >>
rect 267 48 268 49 
<< pdiffusion >>
rect 268 48 269 49 
<< pdiffusion >>
rect 269 48 270 49 
<< m1 >>
rect 271 48 272 49 
<< m1 >>
rect 273 48 274 49 
<< m2 >>
rect 274 48 275 49 
<< m1 >>
rect 277 48 278 49 
<< m1 >>
rect 280 48 281 49 
<< pdiffusion >>
rect 282 48 283 49 
<< pdiffusion >>
rect 283 48 284 49 
<< pdiffusion >>
rect 284 48 285 49 
<< pdiffusion >>
rect 285 48 286 49 
<< pdiffusion >>
rect 286 48 287 49 
<< pdiffusion >>
rect 287 48 288 49 
<< m1 >>
rect 289 48 290 49 
<< pdiffusion >>
rect 300 48 301 49 
<< pdiffusion >>
rect 301 48 302 49 
<< pdiffusion >>
rect 302 48 303 49 
<< pdiffusion >>
rect 303 48 304 49 
<< m1 >>
rect 304 48 305 49 
<< pdiffusion >>
rect 304 48 305 49 
<< pdiffusion >>
rect 305 48 306 49 
<< m1 >>
rect 307 48 308 49 
<< m1 >>
rect 316 48 317 49 
<< pdiffusion >>
rect 318 48 319 49 
<< m1 >>
rect 319 48 320 49 
<< pdiffusion >>
rect 319 48 320 49 
<< pdiffusion >>
rect 320 48 321 49 
<< pdiffusion >>
rect 321 48 322 49 
<< pdiffusion >>
rect 322 48 323 49 
<< pdiffusion >>
rect 323 48 324 49 
<< m1 >>
rect 327 48 328 49 
<< m1 >>
rect 334 48 335 49 
<< m2 >>
rect 334 48 335 49 
<< pdiffusion >>
rect 336 48 337 49 
<< m1 >>
rect 337 48 338 49 
<< pdiffusion >>
rect 337 48 338 49 
<< pdiffusion >>
rect 338 48 339 49 
<< pdiffusion >>
rect 339 48 340 49 
<< pdiffusion >>
rect 340 48 341 49 
<< pdiffusion >>
rect 341 48 342 49 
<< m1 >>
rect 343 48 344 49 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< m1 >>
rect 19 49 20 50 
<< m1 >>
rect 21 49 22 50 
<< m1 >>
rect 23 49 24 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< m1 >>
rect 37 49 38 50 
<< m1 >>
rect 46 49 47 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 55 49 56 50 
<< m2 >>
rect 56 49 57 50 
<< m1 >>
rect 60 49 61 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< m1 >>
rect 73 49 74 50 
<< m2 >>
rect 73 49 74 50 
<< m1 >>
rect 75 49 76 50 
<< m1 >>
rect 78 49 79 50 
<< m2 >>
rect 81 49 82 50 
<< m1 >>
rect 82 49 83 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< m1 >>
rect 97 49 98 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< m1 >>
rect 127 49 128 50 
<< pdiffusion >>
rect 138 49 139 50 
<< pdiffusion >>
rect 139 49 140 50 
<< pdiffusion >>
rect 140 49 141 50 
<< pdiffusion >>
rect 141 49 142 50 
<< pdiffusion >>
rect 142 49 143 50 
<< pdiffusion >>
rect 143 49 144 50 
<< pdiffusion >>
rect 156 49 157 50 
<< pdiffusion >>
rect 157 49 158 50 
<< pdiffusion >>
rect 158 49 159 50 
<< pdiffusion >>
rect 159 49 160 50 
<< pdiffusion >>
rect 160 49 161 50 
<< pdiffusion >>
rect 161 49 162 50 
<< pdiffusion >>
rect 174 49 175 50 
<< pdiffusion >>
rect 175 49 176 50 
<< pdiffusion >>
rect 176 49 177 50 
<< pdiffusion >>
rect 177 49 178 50 
<< pdiffusion >>
rect 178 49 179 50 
<< pdiffusion >>
rect 179 49 180 50 
<< pdiffusion >>
rect 192 49 193 50 
<< pdiffusion >>
rect 193 49 194 50 
<< pdiffusion >>
rect 194 49 195 50 
<< pdiffusion >>
rect 195 49 196 50 
<< pdiffusion >>
rect 196 49 197 50 
<< pdiffusion >>
rect 197 49 198 50 
<< m1 >>
rect 200 49 201 50 
<< m2 >>
rect 201 49 202 50 
<< m1 >>
rect 204 49 205 50 
<< pdiffusion >>
rect 210 49 211 50 
<< pdiffusion >>
rect 211 49 212 50 
<< pdiffusion >>
rect 212 49 213 50 
<< pdiffusion >>
rect 213 49 214 50 
<< pdiffusion >>
rect 214 49 215 50 
<< pdiffusion >>
rect 215 49 216 50 
<< m1 >>
rect 220 49 221 50 
<< m1 >>
rect 226 49 227 50 
<< pdiffusion >>
rect 228 49 229 50 
<< pdiffusion >>
rect 229 49 230 50 
<< pdiffusion >>
rect 230 49 231 50 
<< pdiffusion >>
rect 231 49 232 50 
<< pdiffusion >>
rect 232 49 233 50 
<< pdiffusion >>
rect 233 49 234 50 
<< pdiffusion >>
rect 246 49 247 50 
<< pdiffusion >>
rect 247 49 248 50 
<< pdiffusion >>
rect 248 49 249 50 
<< pdiffusion >>
rect 249 49 250 50 
<< pdiffusion >>
rect 250 49 251 50 
<< pdiffusion >>
rect 251 49 252 50 
<< m1 >>
rect 262 49 263 50 
<< pdiffusion >>
rect 264 49 265 50 
<< pdiffusion >>
rect 265 49 266 50 
<< pdiffusion >>
rect 266 49 267 50 
<< pdiffusion >>
rect 267 49 268 50 
<< pdiffusion >>
rect 268 49 269 50 
<< pdiffusion >>
rect 269 49 270 50 
<< m1 >>
rect 271 49 272 50 
<< m1 >>
rect 273 49 274 50 
<< m2 >>
rect 274 49 275 50 
<< m1 >>
rect 277 49 278 50 
<< m1 >>
rect 280 49 281 50 
<< pdiffusion >>
rect 282 49 283 50 
<< pdiffusion >>
rect 283 49 284 50 
<< pdiffusion >>
rect 284 49 285 50 
<< pdiffusion >>
rect 285 49 286 50 
<< pdiffusion >>
rect 286 49 287 50 
<< pdiffusion >>
rect 287 49 288 50 
<< m1 >>
rect 289 49 290 50 
<< pdiffusion >>
rect 300 49 301 50 
<< pdiffusion >>
rect 301 49 302 50 
<< pdiffusion >>
rect 302 49 303 50 
<< pdiffusion >>
rect 303 49 304 50 
<< pdiffusion >>
rect 304 49 305 50 
<< pdiffusion >>
rect 305 49 306 50 
<< m1 >>
rect 307 49 308 50 
<< m1 >>
rect 316 49 317 50 
<< pdiffusion >>
rect 318 49 319 50 
<< pdiffusion >>
rect 319 49 320 50 
<< pdiffusion >>
rect 320 49 321 50 
<< pdiffusion >>
rect 321 49 322 50 
<< pdiffusion >>
rect 322 49 323 50 
<< pdiffusion >>
rect 323 49 324 50 
<< m1 >>
rect 327 49 328 50 
<< m1 >>
rect 334 49 335 50 
<< m2 >>
rect 334 49 335 50 
<< pdiffusion >>
rect 336 49 337 50 
<< pdiffusion >>
rect 337 49 338 50 
<< pdiffusion >>
rect 338 49 339 50 
<< pdiffusion >>
rect 339 49 340 50 
<< pdiffusion >>
rect 340 49 341 50 
<< pdiffusion >>
rect 341 49 342 50 
<< m1 >>
rect 343 49 344 50 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< m1 >>
rect 19 50 20 51 
<< m1 >>
rect 21 50 22 51 
<< m1 >>
rect 23 50 24 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< m1 >>
rect 37 50 38 51 
<< m1 >>
rect 46 50 47 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 55 50 56 51 
<< m2 >>
rect 56 50 57 51 
<< m1 >>
rect 60 50 61 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< m1 >>
rect 73 50 74 51 
<< m2 >>
rect 73 50 74 51 
<< m1 >>
rect 75 50 76 51 
<< m1 >>
rect 78 50 79 51 
<< m2 >>
rect 81 50 82 51 
<< m1 >>
rect 82 50 83 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< m1 >>
rect 97 50 98 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< m1 >>
rect 127 50 128 51 
<< pdiffusion >>
rect 138 50 139 51 
<< pdiffusion >>
rect 139 50 140 51 
<< pdiffusion >>
rect 140 50 141 51 
<< pdiffusion >>
rect 141 50 142 51 
<< pdiffusion >>
rect 142 50 143 51 
<< pdiffusion >>
rect 143 50 144 51 
<< pdiffusion >>
rect 156 50 157 51 
<< pdiffusion >>
rect 157 50 158 51 
<< pdiffusion >>
rect 158 50 159 51 
<< pdiffusion >>
rect 159 50 160 51 
<< pdiffusion >>
rect 160 50 161 51 
<< pdiffusion >>
rect 161 50 162 51 
<< pdiffusion >>
rect 174 50 175 51 
<< pdiffusion >>
rect 175 50 176 51 
<< pdiffusion >>
rect 176 50 177 51 
<< pdiffusion >>
rect 177 50 178 51 
<< pdiffusion >>
rect 178 50 179 51 
<< pdiffusion >>
rect 179 50 180 51 
<< pdiffusion >>
rect 192 50 193 51 
<< pdiffusion >>
rect 193 50 194 51 
<< pdiffusion >>
rect 194 50 195 51 
<< pdiffusion >>
rect 195 50 196 51 
<< pdiffusion >>
rect 196 50 197 51 
<< pdiffusion >>
rect 197 50 198 51 
<< m1 >>
rect 200 50 201 51 
<< m2 >>
rect 201 50 202 51 
<< m1 >>
rect 204 50 205 51 
<< pdiffusion >>
rect 210 50 211 51 
<< pdiffusion >>
rect 211 50 212 51 
<< pdiffusion >>
rect 212 50 213 51 
<< pdiffusion >>
rect 213 50 214 51 
<< pdiffusion >>
rect 214 50 215 51 
<< pdiffusion >>
rect 215 50 216 51 
<< m1 >>
rect 220 50 221 51 
<< m1 >>
rect 226 50 227 51 
<< pdiffusion >>
rect 228 50 229 51 
<< pdiffusion >>
rect 229 50 230 51 
<< pdiffusion >>
rect 230 50 231 51 
<< pdiffusion >>
rect 231 50 232 51 
<< pdiffusion >>
rect 232 50 233 51 
<< pdiffusion >>
rect 233 50 234 51 
<< pdiffusion >>
rect 246 50 247 51 
<< pdiffusion >>
rect 247 50 248 51 
<< pdiffusion >>
rect 248 50 249 51 
<< pdiffusion >>
rect 249 50 250 51 
<< pdiffusion >>
rect 250 50 251 51 
<< pdiffusion >>
rect 251 50 252 51 
<< m1 >>
rect 262 50 263 51 
<< pdiffusion >>
rect 264 50 265 51 
<< pdiffusion >>
rect 265 50 266 51 
<< pdiffusion >>
rect 266 50 267 51 
<< pdiffusion >>
rect 267 50 268 51 
<< pdiffusion >>
rect 268 50 269 51 
<< pdiffusion >>
rect 269 50 270 51 
<< m1 >>
rect 271 50 272 51 
<< m1 >>
rect 273 50 274 51 
<< m2 >>
rect 274 50 275 51 
<< m1 >>
rect 277 50 278 51 
<< m1 >>
rect 280 50 281 51 
<< pdiffusion >>
rect 282 50 283 51 
<< pdiffusion >>
rect 283 50 284 51 
<< pdiffusion >>
rect 284 50 285 51 
<< pdiffusion >>
rect 285 50 286 51 
<< pdiffusion >>
rect 286 50 287 51 
<< pdiffusion >>
rect 287 50 288 51 
<< m1 >>
rect 289 50 290 51 
<< pdiffusion >>
rect 300 50 301 51 
<< pdiffusion >>
rect 301 50 302 51 
<< pdiffusion >>
rect 302 50 303 51 
<< pdiffusion >>
rect 303 50 304 51 
<< pdiffusion >>
rect 304 50 305 51 
<< pdiffusion >>
rect 305 50 306 51 
<< m1 >>
rect 307 50 308 51 
<< m1 >>
rect 316 50 317 51 
<< pdiffusion >>
rect 318 50 319 51 
<< pdiffusion >>
rect 319 50 320 51 
<< pdiffusion >>
rect 320 50 321 51 
<< pdiffusion >>
rect 321 50 322 51 
<< pdiffusion >>
rect 322 50 323 51 
<< pdiffusion >>
rect 323 50 324 51 
<< m1 >>
rect 327 50 328 51 
<< m1 >>
rect 334 50 335 51 
<< m2 >>
rect 334 50 335 51 
<< pdiffusion >>
rect 336 50 337 51 
<< pdiffusion >>
rect 337 50 338 51 
<< pdiffusion >>
rect 338 50 339 51 
<< pdiffusion >>
rect 339 50 340 51 
<< pdiffusion >>
rect 340 50 341 51 
<< pdiffusion >>
rect 341 50 342 51 
<< m1 >>
rect 343 50 344 51 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< m1 >>
rect 19 51 20 52 
<< m1 >>
rect 21 51 22 52 
<< m1 >>
rect 23 51 24 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< m1 >>
rect 37 51 38 52 
<< m1 >>
rect 46 51 47 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 55 51 56 52 
<< m2 >>
rect 56 51 57 52 
<< m1 >>
rect 60 51 61 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< m1 >>
rect 73 51 74 52 
<< m2 >>
rect 73 51 74 52 
<< m1 >>
rect 75 51 76 52 
<< m1 >>
rect 78 51 79 52 
<< m2 >>
rect 81 51 82 52 
<< m1 >>
rect 82 51 83 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< m1 >>
rect 97 51 98 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< m1 >>
rect 127 51 128 52 
<< pdiffusion >>
rect 138 51 139 52 
<< pdiffusion >>
rect 139 51 140 52 
<< pdiffusion >>
rect 140 51 141 52 
<< pdiffusion >>
rect 141 51 142 52 
<< pdiffusion >>
rect 142 51 143 52 
<< pdiffusion >>
rect 143 51 144 52 
<< pdiffusion >>
rect 156 51 157 52 
<< pdiffusion >>
rect 157 51 158 52 
<< pdiffusion >>
rect 158 51 159 52 
<< pdiffusion >>
rect 159 51 160 52 
<< pdiffusion >>
rect 160 51 161 52 
<< pdiffusion >>
rect 161 51 162 52 
<< pdiffusion >>
rect 174 51 175 52 
<< pdiffusion >>
rect 175 51 176 52 
<< pdiffusion >>
rect 176 51 177 52 
<< pdiffusion >>
rect 177 51 178 52 
<< pdiffusion >>
rect 178 51 179 52 
<< pdiffusion >>
rect 179 51 180 52 
<< pdiffusion >>
rect 192 51 193 52 
<< pdiffusion >>
rect 193 51 194 52 
<< pdiffusion >>
rect 194 51 195 52 
<< pdiffusion >>
rect 195 51 196 52 
<< pdiffusion >>
rect 196 51 197 52 
<< pdiffusion >>
rect 197 51 198 52 
<< m1 >>
rect 200 51 201 52 
<< m2 >>
rect 201 51 202 52 
<< m1 >>
rect 204 51 205 52 
<< m2 >>
rect 204 51 205 52 
<< m2c >>
rect 204 51 205 52 
<< m1 >>
rect 204 51 205 52 
<< m2 >>
rect 204 51 205 52 
<< pdiffusion >>
rect 210 51 211 52 
<< pdiffusion >>
rect 211 51 212 52 
<< pdiffusion >>
rect 212 51 213 52 
<< pdiffusion >>
rect 213 51 214 52 
<< pdiffusion >>
rect 214 51 215 52 
<< pdiffusion >>
rect 215 51 216 52 
<< m1 >>
rect 220 51 221 52 
<< m1 >>
rect 226 51 227 52 
<< pdiffusion >>
rect 228 51 229 52 
<< pdiffusion >>
rect 229 51 230 52 
<< pdiffusion >>
rect 230 51 231 52 
<< pdiffusion >>
rect 231 51 232 52 
<< pdiffusion >>
rect 232 51 233 52 
<< pdiffusion >>
rect 233 51 234 52 
<< pdiffusion >>
rect 246 51 247 52 
<< pdiffusion >>
rect 247 51 248 52 
<< pdiffusion >>
rect 248 51 249 52 
<< pdiffusion >>
rect 249 51 250 52 
<< pdiffusion >>
rect 250 51 251 52 
<< pdiffusion >>
rect 251 51 252 52 
<< m1 >>
rect 262 51 263 52 
<< pdiffusion >>
rect 264 51 265 52 
<< pdiffusion >>
rect 265 51 266 52 
<< pdiffusion >>
rect 266 51 267 52 
<< pdiffusion >>
rect 267 51 268 52 
<< pdiffusion >>
rect 268 51 269 52 
<< pdiffusion >>
rect 269 51 270 52 
<< m1 >>
rect 271 51 272 52 
<< m1 >>
rect 273 51 274 52 
<< m2 >>
rect 274 51 275 52 
<< m1 >>
rect 277 51 278 52 
<< m1 >>
rect 280 51 281 52 
<< pdiffusion >>
rect 282 51 283 52 
<< pdiffusion >>
rect 283 51 284 52 
<< pdiffusion >>
rect 284 51 285 52 
<< pdiffusion >>
rect 285 51 286 52 
<< pdiffusion >>
rect 286 51 287 52 
<< pdiffusion >>
rect 287 51 288 52 
<< m1 >>
rect 289 51 290 52 
<< pdiffusion >>
rect 300 51 301 52 
<< pdiffusion >>
rect 301 51 302 52 
<< pdiffusion >>
rect 302 51 303 52 
<< pdiffusion >>
rect 303 51 304 52 
<< pdiffusion >>
rect 304 51 305 52 
<< pdiffusion >>
rect 305 51 306 52 
<< m1 >>
rect 307 51 308 52 
<< m1 >>
rect 316 51 317 52 
<< pdiffusion >>
rect 318 51 319 52 
<< pdiffusion >>
rect 319 51 320 52 
<< pdiffusion >>
rect 320 51 321 52 
<< pdiffusion >>
rect 321 51 322 52 
<< pdiffusion >>
rect 322 51 323 52 
<< pdiffusion >>
rect 323 51 324 52 
<< m1 >>
rect 327 51 328 52 
<< m1 >>
rect 334 51 335 52 
<< m2 >>
rect 334 51 335 52 
<< pdiffusion >>
rect 336 51 337 52 
<< pdiffusion >>
rect 337 51 338 52 
<< pdiffusion >>
rect 338 51 339 52 
<< pdiffusion >>
rect 339 51 340 52 
<< pdiffusion >>
rect 340 51 341 52 
<< pdiffusion >>
rect 341 51 342 52 
<< m1 >>
rect 343 51 344 52 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< m1 >>
rect 19 52 20 53 
<< m1 >>
rect 21 52 22 53 
<< m1 >>
rect 23 52 24 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< m1 >>
rect 37 52 38 53 
<< m1 >>
rect 46 52 47 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 55 52 56 53 
<< m2 >>
rect 56 52 57 53 
<< m1 >>
rect 60 52 61 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< m1 >>
rect 73 52 74 53 
<< m2 >>
rect 73 52 74 53 
<< m1 >>
rect 75 52 76 53 
<< m1 >>
rect 78 52 79 53 
<< m2 >>
rect 81 52 82 53 
<< m1 >>
rect 82 52 83 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< m1 >>
rect 97 52 98 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< m1 >>
rect 127 52 128 53 
<< pdiffusion >>
rect 138 52 139 53 
<< pdiffusion >>
rect 139 52 140 53 
<< pdiffusion >>
rect 140 52 141 53 
<< pdiffusion >>
rect 141 52 142 53 
<< pdiffusion >>
rect 142 52 143 53 
<< pdiffusion >>
rect 143 52 144 53 
<< pdiffusion >>
rect 156 52 157 53 
<< pdiffusion >>
rect 157 52 158 53 
<< pdiffusion >>
rect 158 52 159 53 
<< pdiffusion >>
rect 159 52 160 53 
<< pdiffusion >>
rect 160 52 161 53 
<< pdiffusion >>
rect 161 52 162 53 
<< pdiffusion >>
rect 174 52 175 53 
<< pdiffusion >>
rect 175 52 176 53 
<< pdiffusion >>
rect 176 52 177 53 
<< pdiffusion >>
rect 177 52 178 53 
<< pdiffusion >>
rect 178 52 179 53 
<< pdiffusion >>
rect 179 52 180 53 
<< pdiffusion >>
rect 192 52 193 53 
<< pdiffusion >>
rect 193 52 194 53 
<< pdiffusion >>
rect 194 52 195 53 
<< pdiffusion >>
rect 195 52 196 53 
<< pdiffusion >>
rect 196 52 197 53 
<< pdiffusion >>
rect 197 52 198 53 
<< m1 >>
rect 200 52 201 53 
<< m2 >>
rect 201 52 202 53 
<< m2 >>
rect 204 52 205 53 
<< pdiffusion >>
rect 210 52 211 53 
<< pdiffusion >>
rect 211 52 212 53 
<< pdiffusion >>
rect 212 52 213 53 
<< pdiffusion >>
rect 213 52 214 53 
<< pdiffusion >>
rect 214 52 215 53 
<< pdiffusion >>
rect 215 52 216 53 
<< m1 >>
rect 220 52 221 53 
<< m1 >>
rect 226 52 227 53 
<< pdiffusion >>
rect 228 52 229 53 
<< pdiffusion >>
rect 229 52 230 53 
<< pdiffusion >>
rect 230 52 231 53 
<< pdiffusion >>
rect 231 52 232 53 
<< pdiffusion >>
rect 232 52 233 53 
<< pdiffusion >>
rect 233 52 234 53 
<< pdiffusion >>
rect 246 52 247 53 
<< pdiffusion >>
rect 247 52 248 53 
<< pdiffusion >>
rect 248 52 249 53 
<< pdiffusion >>
rect 249 52 250 53 
<< pdiffusion >>
rect 250 52 251 53 
<< pdiffusion >>
rect 251 52 252 53 
<< m1 >>
rect 262 52 263 53 
<< pdiffusion >>
rect 264 52 265 53 
<< pdiffusion >>
rect 265 52 266 53 
<< pdiffusion >>
rect 266 52 267 53 
<< pdiffusion >>
rect 267 52 268 53 
<< pdiffusion >>
rect 268 52 269 53 
<< pdiffusion >>
rect 269 52 270 53 
<< m1 >>
rect 271 52 272 53 
<< m1 >>
rect 273 52 274 53 
<< m2 >>
rect 274 52 275 53 
<< m1 >>
rect 277 52 278 53 
<< m1 >>
rect 280 52 281 53 
<< pdiffusion >>
rect 282 52 283 53 
<< pdiffusion >>
rect 283 52 284 53 
<< pdiffusion >>
rect 284 52 285 53 
<< pdiffusion >>
rect 285 52 286 53 
<< pdiffusion >>
rect 286 52 287 53 
<< pdiffusion >>
rect 287 52 288 53 
<< m1 >>
rect 289 52 290 53 
<< pdiffusion >>
rect 300 52 301 53 
<< pdiffusion >>
rect 301 52 302 53 
<< pdiffusion >>
rect 302 52 303 53 
<< pdiffusion >>
rect 303 52 304 53 
<< pdiffusion >>
rect 304 52 305 53 
<< pdiffusion >>
rect 305 52 306 53 
<< m1 >>
rect 307 52 308 53 
<< m1 >>
rect 316 52 317 53 
<< pdiffusion >>
rect 318 52 319 53 
<< pdiffusion >>
rect 319 52 320 53 
<< pdiffusion >>
rect 320 52 321 53 
<< pdiffusion >>
rect 321 52 322 53 
<< pdiffusion >>
rect 322 52 323 53 
<< pdiffusion >>
rect 323 52 324 53 
<< m1 >>
rect 327 52 328 53 
<< m1 >>
rect 334 52 335 53 
<< m2 >>
rect 334 52 335 53 
<< pdiffusion >>
rect 336 52 337 53 
<< pdiffusion >>
rect 337 52 338 53 
<< pdiffusion >>
rect 338 52 339 53 
<< pdiffusion >>
rect 339 52 340 53 
<< pdiffusion >>
rect 340 52 341 53 
<< pdiffusion >>
rect 341 52 342 53 
<< m1 >>
rect 343 52 344 53 
<< pdiffusion >>
rect 12 53 13 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< m1 >>
rect 19 53 20 54 
<< m1 >>
rect 21 53 22 54 
<< m1 >>
rect 23 53 24 54 
<< pdiffusion >>
rect 30 53 31 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< m1 >>
rect 37 53 38 54 
<< m1 >>
rect 46 53 47 54 
<< pdiffusion >>
rect 48 53 49 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 55 53 56 54 
<< m2 >>
rect 56 53 57 54 
<< m1 >>
rect 60 53 61 54 
<< pdiffusion >>
rect 66 53 67 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< m1 >>
rect 73 53 74 54 
<< m2 >>
rect 73 53 74 54 
<< m1 >>
rect 75 53 76 54 
<< m1 >>
rect 78 53 79 54 
<< m2 >>
rect 81 53 82 54 
<< m1 >>
rect 82 53 83 54 
<< pdiffusion >>
rect 84 53 85 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< m1 >>
rect 97 53 98 54 
<< pdiffusion >>
rect 102 53 103 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< pdiffusion >>
rect 120 53 121 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< m1 >>
rect 127 53 128 54 
<< pdiffusion >>
rect 138 53 139 54 
<< pdiffusion >>
rect 139 53 140 54 
<< pdiffusion >>
rect 140 53 141 54 
<< pdiffusion >>
rect 141 53 142 54 
<< pdiffusion >>
rect 142 53 143 54 
<< pdiffusion >>
rect 143 53 144 54 
<< pdiffusion >>
rect 156 53 157 54 
<< pdiffusion >>
rect 157 53 158 54 
<< pdiffusion >>
rect 158 53 159 54 
<< pdiffusion >>
rect 159 53 160 54 
<< pdiffusion >>
rect 160 53 161 54 
<< pdiffusion >>
rect 161 53 162 54 
<< pdiffusion >>
rect 174 53 175 54 
<< pdiffusion >>
rect 175 53 176 54 
<< pdiffusion >>
rect 176 53 177 54 
<< pdiffusion >>
rect 177 53 178 54 
<< pdiffusion >>
rect 178 53 179 54 
<< pdiffusion >>
rect 179 53 180 54 
<< pdiffusion >>
rect 192 53 193 54 
<< pdiffusion >>
rect 193 53 194 54 
<< pdiffusion >>
rect 194 53 195 54 
<< pdiffusion >>
rect 195 53 196 54 
<< pdiffusion >>
rect 196 53 197 54 
<< pdiffusion >>
rect 197 53 198 54 
<< m1 >>
rect 200 53 201 54 
<< m2 >>
rect 201 53 202 54 
<< m1 >>
rect 202 53 203 54 
<< m2 >>
rect 202 53 203 54 
<< m2c >>
rect 202 53 203 54 
<< m1 >>
rect 202 53 203 54 
<< m2 >>
rect 202 53 203 54 
<< m1 >>
rect 203 53 204 54 
<< m1 >>
rect 204 53 205 54 
<< m2 >>
rect 204 53 205 54 
<< m1 >>
rect 205 53 206 54 
<< m1 >>
rect 206 53 207 54 
<< m1 >>
rect 207 53 208 54 
<< m1 >>
rect 208 53 209 54 
<< pdiffusion >>
rect 210 53 211 54 
<< m1 >>
rect 211 53 212 54 
<< pdiffusion >>
rect 211 53 212 54 
<< pdiffusion >>
rect 212 53 213 54 
<< pdiffusion >>
rect 213 53 214 54 
<< pdiffusion >>
rect 214 53 215 54 
<< pdiffusion >>
rect 215 53 216 54 
<< m1 >>
rect 220 53 221 54 
<< m1 >>
rect 226 53 227 54 
<< pdiffusion >>
rect 228 53 229 54 
<< pdiffusion >>
rect 229 53 230 54 
<< pdiffusion >>
rect 230 53 231 54 
<< pdiffusion >>
rect 231 53 232 54 
<< pdiffusion >>
rect 232 53 233 54 
<< pdiffusion >>
rect 233 53 234 54 
<< pdiffusion >>
rect 246 53 247 54 
<< pdiffusion >>
rect 247 53 248 54 
<< pdiffusion >>
rect 248 53 249 54 
<< pdiffusion >>
rect 249 53 250 54 
<< pdiffusion >>
rect 250 53 251 54 
<< pdiffusion >>
rect 251 53 252 54 
<< m1 >>
rect 262 53 263 54 
<< pdiffusion >>
rect 264 53 265 54 
<< m1 >>
rect 265 53 266 54 
<< pdiffusion >>
rect 265 53 266 54 
<< pdiffusion >>
rect 266 53 267 54 
<< pdiffusion >>
rect 267 53 268 54 
<< pdiffusion >>
rect 268 53 269 54 
<< pdiffusion >>
rect 269 53 270 54 
<< m1 >>
rect 271 53 272 54 
<< m1 >>
rect 273 53 274 54 
<< m2 >>
rect 274 53 275 54 
<< m1 >>
rect 277 53 278 54 
<< m1 >>
rect 280 53 281 54 
<< pdiffusion >>
rect 282 53 283 54 
<< pdiffusion >>
rect 283 53 284 54 
<< pdiffusion >>
rect 284 53 285 54 
<< pdiffusion >>
rect 285 53 286 54 
<< m1 >>
rect 286 53 287 54 
<< pdiffusion >>
rect 286 53 287 54 
<< pdiffusion >>
rect 287 53 288 54 
<< m1 >>
rect 289 53 290 54 
<< pdiffusion >>
rect 300 53 301 54 
<< pdiffusion >>
rect 301 53 302 54 
<< pdiffusion >>
rect 302 53 303 54 
<< pdiffusion >>
rect 303 53 304 54 
<< pdiffusion >>
rect 304 53 305 54 
<< pdiffusion >>
rect 305 53 306 54 
<< m1 >>
rect 307 53 308 54 
<< m1 >>
rect 316 53 317 54 
<< pdiffusion >>
rect 318 53 319 54 
<< pdiffusion >>
rect 319 53 320 54 
<< pdiffusion >>
rect 320 53 321 54 
<< pdiffusion >>
rect 321 53 322 54 
<< pdiffusion >>
rect 322 53 323 54 
<< pdiffusion >>
rect 323 53 324 54 
<< m1 >>
rect 327 53 328 54 
<< m1 >>
rect 334 53 335 54 
<< m2 >>
rect 334 53 335 54 
<< pdiffusion >>
rect 336 53 337 54 
<< pdiffusion >>
rect 337 53 338 54 
<< pdiffusion >>
rect 338 53 339 54 
<< pdiffusion >>
rect 339 53 340 54 
<< pdiffusion >>
rect 340 53 341 54 
<< pdiffusion >>
rect 341 53 342 54 
<< m1 >>
rect 343 53 344 54 
<< m1 >>
rect 19 54 20 55 
<< m1 >>
rect 21 54 22 55 
<< m1 >>
rect 23 54 24 55 
<< m1 >>
rect 37 54 38 55 
<< m1 >>
rect 46 54 47 55 
<< m1 >>
rect 55 54 56 55 
<< m2 >>
rect 56 54 57 55 
<< m1 >>
rect 60 54 61 55 
<< m1 >>
rect 73 54 74 55 
<< m2 >>
rect 73 54 74 55 
<< m1 >>
rect 75 54 76 55 
<< m1 >>
rect 78 54 79 55 
<< m2 >>
rect 81 54 82 55 
<< m1 >>
rect 82 54 83 55 
<< m1 >>
rect 91 54 92 55 
<< m1 >>
rect 97 54 98 55 
<< m1 >>
rect 127 54 128 55 
<< m1 >>
rect 200 54 201 55 
<< m2 >>
rect 204 54 205 55 
<< m1 >>
rect 208 54 209 55 
<< m1 >>
rect 211 54 212 55 
<< m1 >>
rect 220 54 221 55 
<< m1 >>
rect 226 54 227 55 
<< m1 >>
rect 262 54 263 55 
<< m1 >>
rect 265 54 266 55 
<< m1 >>
rect 271 54 272 55 
<< m1 >>
rect 273 54 274 55 
<< m2 >>
rect 274 54 275 55 
<< m1 >>
rect 277 54 278 55 
<< m1 >>
rect 280 54 281 55 
<< m1 >>
rect 286 54 287 55 
<< m1 >>
rect 289 54 290 55 
<< m1 >>
rect 307 54 308 55 
<< m1 >>
rect 316 54 317 55 
<< m1 >>
rect 327 54 328 55 
<< m1 >>
rect 334 54 335 55 
<< m2 >>
rect 334 54 335 55 
<< m1 >>
rect 343 54 344 55 
<< m1 >>
rect 19 55 20 56 
<< m1 >>
rect 21 55 22 56 
<< m1 >>
rect 23 55 24 56 
<< m1 >>
rect 37 55 38 56 
<< m1 >>
rect 46 55 47 56 
<< m1 >>
rect 53 55 54 56 
<< m2 >>
rect 53 55 54 56 
<< m2c >>
rect 53 55 54 56 
<< m1 >>
rect 53 55 54 56 
<< m2 >>
rect 53 55 54 56 
<< m2 >>
rect 54 55 55 56 
<< m1 >>
rect 55 55 56 56 
<< m2 >>
rect 55 55 56 56 
<< m2 >>
rect 56 55 57 56 
<< m1 >>
rect 60 55 61 56 
<< m1 >>
rect 71 55 72 56 
<< m2 >>
rect 71 55 72 56 
<< m2c >>
rect 71 55 72 56 
<< m1 >>
rect 71 55 72 56 
<< m2 >>
rect 71 55 72 56 
<< m1 >>
rect 72 55 73 56 
<< m1 >>
rect 73 55 74 56 
<< m2 >>
rect 73 55 74 56 
<< m1 >>
rect 75 55 76 56 
<< m2 >>
rect 75 55 76 56 
<< m2c >>
rect 75 55 76 56 
<< m1 >>
rect 75 55 76 56 
<< m2 >>
rect 75 55 76 56 
<< m1 >>
rect 78 55 79 56 
<< m2 >>
rect 78 55 79 56 
<< m2c >>
rect 78 55 79 56 
<< m1 >>
rect 78 55 79 56 
<< m2 >>
rect 78 55 79 56 
<< m2 >>
rect 81 55 82 56 
<< m1 >>
rect 82 55 83 56 
<< m1 >>
rect 91 55 92 56 
<< m1 >>
rect 97 55 98 56 
<< m1 >>
rect 127 55 128 56 
<< m1 >>
rect 200 55 201 56 
<< m2 >>
rect 200 55 201 56 
<< m2c >>
rect 200 55 201 56 
<< m1 >>
rect 200 55 201 56 
<< m2 >>
rect 200 55 201 56 
<< m1 >>
rect 204 55 205 56 
<< m2 >>
rect 204 55 205 56 
<< m2c >>
rect 204 55 205 56 
<< m1 >>
rect 204 55 205 56 
<< m2 >>
rect 204 55 205 56 
<< m1 >>
rect 208 55 209 56 
<< m1 >>
rect 209 55 210 56 
<< m2 >>
rect 209 55 210 56 
<< m2c >>
rect 209 55 210 56 
<< m1 >>
rect 209 55 210 56 
<< m2 >>
rect 209 55 210 56 
<< m2 >>
rect 210 55 211 56 
<< m1 >>
rect 211 55 212 56 
<< m1 >>
rect 220 55 221 56 
<< m1 >>
rect 226 55 227 56 
<< m1 >>
rect 262 55 263 56 
<< m1 >>
rect 265 55 266 56 
<< m1 >>
rect 271 55 272 56 
<< m1 >>
rect 273 55 274 56 
<< m2 >>
rect 274 55 275 56 
<< m1 >>
rect 277 55 278 56 
<< m1 >>
rect 280 55 281 56 
<< m1 >>
rect 286 55 287 56 
<< m1 >>
rect 287 55 288 56 
<< m1 >>
rect 288 55 289 56 
<< m1 >>
rect 289 55 290 56 
<< m1 >>
rect 307 55 308 56 
<< m1 >>
rect 316 55 317 56 
<< m1 >>
rect 327 55 328 56 
<< m1 >>
rect 334 55 335 56 
<< m2 >>
rect 334 55 335 56 
<< m1 >>
rect 343 55 344 56 
<< m1 >>
rect 19 56 20 57 
<< m1 >>
rect 21 56 22 57 
<< m1 >>
rect 23 56 24 57 
<< m1 >>
rect 37 56 38 57 
<< m1 >>
rect 46 56 47 57 
<< m1 >>
rect 53 56 54 57 
<< m1 >>
rect 55 56 56 57 
<< m1 >>
rect 60 56 61 57 
<< m2 >>
rect 71 56 72 57 
<< m2 >>
rect 73 56 74 57 
<< m2 >>
rect 75 56 76 57 
<< m2 >>
rect 78 56 79 57 
<< m2 >>
rect 81 56 82 57 
<< m1 >>
rect 82 56 83 57 
<< m2 >>
rect 90 56 91 57 
<< m1 >>
rect 91 56 92 57 
<< m2 >>
rect 91 56 92 57 
<< m2 >>
rect 92 56 93 57 
<< m1 >>
rect 93 56 94 57 
<< m2 >>
rect 93 56 94 57 
<< m2c >>
rect 93 56 94 57 
<< m1 >>
rect 93 56 94 57 
<< m2 >>
rect 93 56 94 57 
<< m1 >>
rect 94 56 95 57 
<< m1 >>
rect 95 56 96 57 
<< m2 >>
rect 95 56 96 57 
<< m2c >>
rect 95 56 96 57 
<< m1 >>
rect 95 56 96 57 
<< m2 >>
rect 95 56 96 57 
<< m1 >>
rect 97 56 98 57 
<< m2 >>
rect 97 56 98 57 
<< m2c >>
rect 97 56 98 57 
<< m1 >>
rect 97 56 98 57 
<< m2 >>
rect 97 56 98 57 
<< m1 >>
rect 127 56 128 57 
<< m2 >>
rect 200 56 201 57 
<< m2 >>
rect 204 56 205 57 
<< m2 >>
rect 210 56 211 57 
<< m1 >>
rect 211 56 212 57 
<< m1 >>
rect 220 56 221 57 
<< m2 >>
rect 220 56 221 57 
<< m2c >>
rect 220 56 221 57 
<< m1 >>
rect 220 56 221 57 
<< m2 >>
rect 220 56 221 57 
<< m1 >>
rect 226 56 227 57 
<< m2 >>
rect 226 56 227 57 
<< m2c >>
rect 226 56 227 57 
<< m1 >>
rect 226 56 227 57 
<< m2 >>
rect 226 56 227 57 
<< m1 >>
rect 262 56 263 57 
<< m1 >>
rect 265 56 266 57 
<< m1 >>
rect 271 56 272 57 
<< m1 >>
rect 273 56 274 57 
<< m2 >>
rect 274 56 275 57 
<< m1 >>
rect 277 56 278 57 
<< m1 >>
rect 280 56 281 57 
<< m1 >>
rect 307 56 308 57 
<< m1 >>
rect 316 56 317 57 
<< m1 >>
rect 327 56 328 57 
<< m1 >>
rect 334 56 335 57 
<< m2 >>
rect 334 56 335 57 
<< m1 >>
rect 343 56 344 57 
<< m1 >>
rect 19 57 20 58 
<< m1 >>
rect 21 57 22 58 
<< m1 >>
rect 23 57 24 58 
<< m1 >>
rect 35 57 36 58 
<< m2 >>
rect 35 57 36 58 
<< m2c >>
rect 35 57 36 58 
<< m1 >>
rect 35 57 36 58 
<< m2 >>
rect 35 57 36 58 
<< m2 >>
rect 36 57 37 58 
<< m1 >>
rect 37 57 38 58 
<< m2 >>
rect 37 57 38 58 
<< m2 >>
rect 38 57 39 58 
<< m1 >>
rect 39 57 40 58 
<< m2 >>
rect 39 57 40 58 
<< m2c >>
rect 39 57 40 58 
<< m1 >>
rect 39 57 40 58 
<< m2 >>
rect 39 57 40 58 
<< m1 >>
rect 40 57 41 58 
<< m1 >>
rect 41 57 42 58 
<< m1 >>
rect 42 57 43 58 
<< m1 >>
rect 43 57 44 58 
<< m1 >>
rect 44 57 45 58 
<< m2 >>
rect 44 57 45 58 
<< m2c >>
rect 44 57 45 58 
<< m1 >>
rect 44 57 45 58 
<< m2 >>
rect 44 57 45 58 
<< m2 >>
rect 45 57 46 58 
<< m1 >>
rect 46 57 47 58 
<< m2 >>
rect 46 57 47 58 
<< m2 >>
rect 47 57 48 58 
<< m1 >>
rect 48 57 49 58 
<< m2 >>
rect 48 57 49 58 
<< m2c >>
rect 48 57 49 58 
<< m1 >>
rect 48 57 49 58 
<< m2 >>
rect 48 57 49 58 
<< m1 >>
rect 53 57 54 58 
<< m1 >>
rect 55 57 56 58 
<< m1 >>
rect 60 57 61 58 
<< m1 >>
rect 68 57 69 58 
<< m1 >>
rect 69 57 70 58 
<< m1 >>
rect 70 57 71 58 
<< m1 >>
rect 71 57 72 58 
<< m2 >>
rect 71 57 72 58 
<< m1 >>
rect 72 57 73 58 
<< m1 >>
rect 73 57 74 58 
<< m2 >>
rect 73 57 74 58 
<< m1 >>
rect 74 57 75 58 
<< m1 >>
rect 75 57 76 58 
<< m2 >>
rect 75 57 76 58 
<< m1 >>
rect 76 57 77 58 
<< m1 >>
rect 77 57 78 58 
<< m1 >>
rect 78 57 79 58 
<< m2 >>
rect 78 57 79 58 
<< m1 >>
rect 79 57 80 58 
<< m1 >>
rect 80 57 81 58 
<< m2 >>
rect 80 57 81 58 
<< m2c >>
rect 80 57 81 58 
<< m1 >>
rect 80 57 81 58 
<< m2 >>
rect 80 57 81 58 
<< m2 >>
rect 81 57 82 58 
<< m1 >>
rect 82 57 83 58 
<< m2 >>
rect 90 57 91 58 
<< m1 >>
rect 91 57 92 58 
<< m2 >>
rect 95 57 96 58 
<< m2 >>
rect 97 57 98 58 
<< m1 >>
rect 127 57 128 58 
<< m2 >>
rect 197 57 198 58 
<< m1 >>
rect 198 57 199 58 
<< m2 >>
rect 198 57 199 58 
<< m2c >>
rect 198 57 199 58 
<< m1 >>
rect 198 57 199 58 
<< m2 >>
rect 198 57 199 58 
<< m1 >>
rect 199 57 200 58 
<< m1 >>
rect 200 57 201 58 
<< m2 >>
rect 200 57 201 58 
<< m1 >>
rect 201 57 202 58 
<< m1 >>
rect 202 57 203 58 
<< m1 >>
rect 203 57 204 58 
<< m1 >>
rect 204 57 205 58 
<< m2 >>
rect 204 57 205 58 
<< m1 >>
rect 205 57 206 58 
<< m1 >>
rect 206 57 207 58 
<< m1 >>
rect 207 57 208 58 
<< m1 >>
rect 208 57 209 58 
<< m1 >>
rect 209 57 210 58 
<< m1 >>
rect 210 57 211 58 
<< m2 >>
rect 210 57 211 58 
<< m1 >>
rect 211 57 212 58 
<< m2 >>
rect 220 57 221 58 
<< m2 >>
rect 226 57 227 58 
<< m1 >>
rect 262 57 263 58 
<< m1 >>
rect 265 57 266 58 
<< m1 >>
rect 271 57 272 58 
<< m1 >>
rect 273 57 274 58 
<< m2 >>
rect 274 57 275 58 
<< m1 >>
rect 277 57 278 58 
<< m1 >>
rect 280 57 281 58 
<< m1 >>
rect 307 57 308 58 
<< m1 >>
rect 316 57 317 58 
<< m1 >>
rect 327 57 328 58 
<< m1 >>
rect 334 57 335 58 
<< m2 >>
rect 334 57 335 58 
<< m1 >>
rect 343 57 344 58 
<< m1 >>
rect 19 58 20 59 
<< m1 >>
rect 21 58 22 59 
<< m1 >>
rect 23 58 24 59 
<< m1 >>
rect 35 58 36 59 
<< m1 >>
rect 37 58 38 59 
<< m1 >>
rect 46 58 47 59 
<< m1 >>
rect 48 58 49 59 
<< m1 >>
rect 49 58 50 59 
<< m1 >>
rect 50 58 51 59 
<< m1 >>
rect 51 58 52 59 
<< m1 >>
rect 52 58 53 59 
<< m1 >>
rect 53 58 54 59 
<< m1 >>
rect 55 58 56 59 
<< m1 >>
rect 60 58 61 59 
<< m2 >>
rect 64 58 65 59 
<< m2 >>
rect 65 58 66 59 
<< m2 >>
rect 66 58 67 59 
<< m2 >>
rect 67 58 68 59 
<< m1 >>
rect 68 58 69 59 
<< m2 >>
rect 68 58 69 59 
<< m2 >>
rect 69 58 70 59 
<< m2 >>
rect 70 58 71 59 
<< m2 >>
rect 71 58 72 59 
<< m2 >>
rect 73 58 74 59 
<< m2 >>
rect 75 58 76 59 
<< m2 >>
rect 78 58 79 59 
<< m1 >>
rect 82 58 83 59 
<< m2 >>
rect 90 58 91 59 
<< m1 >>
rect 91 58 92 59 
<< m2 >>
rect 92 58 93 59 
<< m1 >>
rect 93 58 94 59 
<< m2 >>
rect 93 58 94 59 
<< m2c >>
rect 93 58 94 59 
<< m1 >>
rect 93 58 94 59 
<< m2 >>
rect 93 58 94 59 
<< m1 >>
rect 94 58 95 59 
<< m1 >>
rect 95 58 96 59 
<< m2 >>
rect 95 58 96 59 
<< m1 >>
rect 96 58 97 59 
<< m1 >>
rect 97 58 98 59 
<< m2 >>
rect 97 58 98 59 
<< m1 >>
rect 98 58 99 59 
<< m1 >>
rect 99 58 100 59 
<< m1 >>
rect 100 58 101 59 
<< m1 >>
rect 101 58 102 59 
<< m1 >>
rect 102 58 103 59 
<< m1 >>
rect 103 58 104 59 
<< m1 >>
rect 104 58 105 59 
<< m1 >>
rect 105 58 106 59 
<< m1 >>
rect 106 58 107 59 
<< m1 >>
rect 107 58 108 59 
<< m1 >>
rect 108 58 109 59 
<< m1 >>
rect 109 58 110 59 
<< m1 >>
rect 110 58 111 59 
<< m1 >>
rect 111 58 112 59 
<< m1 >>
rect 112 58 113 59 
<< m1 >>
rect 113 58 114 59 
<< m1 >>
rect 114 58 115 59 
<< m1 >>
rect 115 58 116 59 
<< m1 >>
rect 116 58 117 59 
<< m1 >>
rect 117 58 118 59 
<< m1 >>
rect 118 58 119 59 
<< m1 >>
rect 119 58 120 59 
<< m1 >>
rect 120 58 121 59 
<< m1 >>
rect 121 58 122 59 
<< m1 >>
rect 122 58 123 59 
<< m1 >>
rect 123 58 124 59 
<< m1 >>
rect 124 58 125 59 
<< m1 >>
rect 125 58 126 59 
<< m2 >>
rect 125 58 126 59 
<< m2c >>
rect 125 58 126 59 
<< m1 >>
rect 125 58 126 59 
<< m2 >>
rect 125 58 126 59 
<< m2 >>
rect 126 58 127 59 
<< m1 >>
rect 127 58 128 59 
<< m2 >>
rect 127 58 128 59 
<< m1 >>
rect 128 58 129 59 
<< m2 >>
rect 128 58 129 59 
<< m1 >>
rect 129 58 130 59 
<< m2 >>
rect 129 58 130 59 
<< m1 >>
rect 130 58 131 59 
<< m2 >>
rect 130 58 131 59 
<< m1 >>
rect 131 58 132 59 
<< m2 >>
rect 131 58 132 59 
<< m1 >>
rect 132 58 133 59 
<< m2 >>
rect 132 58 133 59 
<< m1 >>
rect 133 58 134 59 
<< m2 >>
rect 133 58 134 59 
<< m1 >>
rect 134 58 135 59 
<< m2 >>
rect 134 58 135 59 
<< m1 >>
rect 135 58 136 59 
<< m2 >>
rect 135 58 136 59 
<< m1 >>
rect 136 58 137 59 
<< m2 >>
rect 136 58 137 59 
<< m1 >>
rect 137 58 138 59 
<< m2 >>
rect 137 58 138 59 
<< m1 >>
rect 138 58 139 59 
<< m2 >>
rect 138 58 139 59 
<< m1 >>
rect 139 58 140 59 
<< m2 >>
rect 139 58 140 59 
<< m1 >>
rect 140 58 141 59 
<< m2 >>
rect 140 58 141 59 
<< m1 >>
rect 141 58 142 59 
<< m2 >>
rect 141 58 142 59 
<< m1 >>
rect 142 58 143 59 
<< m2 >>
rect 142 58 143 59 
<< m1 >>
rect 143 58 144 59 
<< m2 >>
rect 143 58 144 59 
<< m1 >>
rect 144 58 145 59 
<< m2 >>
rect 144 58 145 59 
<< m1 >>
rect 145 58 146 59 
<< m2 >>
rect 145 58 146 59 
<< m1 >>
rect 146 58 147 59 
<< m2 >>
rect 146 58 147 59 
<< m1 >>
rect 147 58 148 59 
<< m2 >>
rect 147 58 148 59 
<< m1 >>
rect 148 58 149 59 
<< m2 >>
rect 148 58 149 59 
<< m1 >>
rect 149 58 150 59 
<< m2 >>
rect 149 58 150 59 
<< m1 >>
rect 150 58 151 59 
<< m2 >>
rect 150 58 151 59 
<< m1 >>
rect 151 58 152 59 
<< m2 >>
rect 151 58 152 59 
<< m1 >>
rect 152 58 153 59 
<< m2 >>
rect 152 58 153 59 
<< m1 >>
rect 153 58 154 59 
<< m2 >>
rect 153 58 154 59 
<< m1 >>
rect 154 58 155 59 
<< m2 >>
rect 154 58 155 59 
<< m1 >>
rect 155 58 156 59 
<< m2 >>
rect 155 58 156 59 
<< m1 >>
rect 156 58 157 59 
<< m2 >>
rect 156 58 157 59 
<< m1 >>
rect 157 58 158 59 
<< m2 >>
rect 157 58 158 59 
<< m1 >>
rect 158 58 159 59 
<< m2 >>
rect 158 58 159 59 
<< m1 >>
rect 159 58 160 59 
<< m2 >>
rect 159 58 160 59 
<< m1 >>
rect 160 58 161 59 
<< m2 >>
rect 160 58 161 59 
<< m1 >>
rect 161 58 162 59 
<< m2 >>
rect 161 58 162 59 
<< m1 >>
rect 162 58 163 59 
<< m2 >>
rect 162 58 163 59 
<< m1 >>
rect 163 58 164 59 
<< m2 >>
rect 163 58 164 59 
<< m1 >>
rect 164 58 165 59 
<< m2 >>
rect 164 58 165 59 
<< m1 >>
rect 165 58 166 59 
<< m2 >>
rect 165 58 166 59 
<< m1 >>
rect 166 58 167 59 
<< m2 >>
rect 166 58 167 59 
<< m1 >>
rect 167 58 168 59 
<< m2 >>
rect 167 58 168 59 
<< m1 >>
rect 168 58 169 59 
<< m2 >>
rect 168 58 169 59 
<< m1 >>
rect 169 58 170 59 
<< m2 >>
rect 169 58 170 59 
<< m1 >>
rect 170 58 171 59 
<< m2 >>
rect 170 58 171 59 
<< m1 >>
rect 171 58 172 59 
<< m2 >>
rect 171 58 172 59 
<< m1 >>
rect 172 58 173 59 
<< m2 >>
rect 172 58 173 59 
<< m1 >>
rect 173 58 174 59 
<< m2 >>
rect 173 58 174 59 
<< m1 >>
rect 174 58 175 59 
<< m2 >>
rect 174 58 175 59 
<< m1 >>
rect 175 58 176 59 
<< m2 >>
rect 175 58 176 59 
<< m1 >>
rect 176 58 177 59 
<< m2 >>
rect 176 58 177 59 
<< m1 >>
rect 177 58 178 59 
<< m2 >>
rect 177 58 178 59 
<< m1 >>
rect 178 58 179 59 
<< m2 >>
rect 178 58 179 59 
<< m1 >>
rect 179 58 180 59 
<< m2 >>
rect 179 58 180 59 
<< m1 >>
rect 180 58 181 59 
<< m2 >>
rect 180 58 181 59 
<< m1 >>
rect 181 58 182 59 
<< m2 >>
rect 181 58 182 59 
<< m1 >>
rect 182 58 183 59 
<< m2 >>
rect 182 58 183 59 
<< m1 >>
rect 183 58 184 59 
<< m2 >>
rect 183 58 184 59 
<< m1 >>
rect 184 58 185 59 
<< m2 >>
rect 184 58 185 59 
<< m1 >>
rect 185 58 186 59 
<< m2 >>
rect 185 58 186 59 
<< m1 >>
rect 186 58 187 59 
<< m2 >>
rect 186 58 187 59 
<< m1 >>
rect 187 58 188 59 
<< m2 >>
rect 187 58 188 59 
<< m1 >>
rect 188 58 189 59 
<< m2 >>
rect 188 58 189 59 
<< m1 >>
rect 189 58 190 59 
<< m2 >>
rect 189 58 190 59 
<< m1 >>
rect 190 58 191 59 
<< m2 >>
rect 190 58 191 59 
<< m1 >>
rect 191 58 192 59 
<< m2 >>
rect 191 58 192 59 
<< m1 >>
rect 192 58 193 59 
<< m2 >>
rect 192 58 193 59 
<< m1 >>
rect 193 58 194 59 
<< m2 >>
rect 193 58 194 59 
<< m1 >>
rect 194 58 195 59 
<< m2 >>
rect 194 58 195 59 
<< m1 >>
rect 195 58 196 59 
<< m2 >>
rect 195 58 196 59 
<< m1 >>
rect 196 58 197 59 
<< m2 >>
rect 196 58 197 59 
<< m2 >>
rect 197 58 198 59 
<< m2 >>
rect 200 58 201 59 
<< m2 >>
rect 204 58 205 59 
<< m2 >>
rect 210 58 211 59 
<< m2 >>
rect 211 58 212 59 
<< m2 >>
rect 212 58 213 59 
<< m1 >>
rect 213 58 214 59 
<< m2 >>
rect 213 58 214 59 
<< m2c >>
rect 213 58 214 59 
<< m1 >>
rect 213 58 214 59 
<< m2 >>
rect 213 58 214 59 
<< m1 >>
rect 214 58 215 59 
<< m1 >>
rect 215 58 216 59 
<< m1 >>
rect 216 58 217 59 
<< m1 >>
rect 217 58 218 59 
<< m1 >>
rect 218 58 219 59 
<< m1 >>
rect 219 58 220 59 
<< m1 >>
rect 220 58 221 59 
<< m2 >>
rect 220 58 221 59 
<< m1 >>
rect 221 58 222 59 
<< m1 >>
rect 222 58 223 59 
<< m1 >>
rect 223 58 224 59 
<< m1 >>
rect 224 58 225 59 
<< m1 >>
rect 225 58 226 59 
<< m1 >>
rect 226 58 227 59 
<< m2 >>
rect 226 58 227 59 
<< m1 >>
rect 227 58 228 59 
<< m1 >>
rect 228 58 229 59 
<< m1 >>
rect 229 58 230 59 
<< m1 >>
rect 230 58 231 59 
<< m1 >>
rect 231 58 232 59 
<< m1 >>
rect 232 58 233 59 
<< m1 >>
rect 233 58 234 59 
<< m1 >>
rect 234 58 235 59 
<< m1 >>
rect 235 58 236 59 
<< m1 >>
rect 236 58 237 59 
<< m1 >>
rect 237 58 238 59 
<< m1 >>
rect 238 58 239 59 
<< m1 >>
rect 239 58 240 59 
<< m1 >>
rect 240 58 241 59 
<< m1 >>
rect 241 58 242 59 
<< m1 >>
rect 242 58 243 59 
<< m1 >>
rect 243 58 244 59 
<< m1 >>
rect 244 58 245 59 
<< m1 >>
rect 245 58 246 59 
<< m1 >>
rect 246 58 247 59 
<< m1 >>
rect 247 58 248 59 
<< m1 >>
rect 248 58 249 59 
<< m1 >>
rect 249 58 250 59 
<< m1 >>
rect 250 58 251 59 
<< m1 >>
rect 251 58 252 59 
<< m1 >>
rect 252 58 253 59 
<< m1 >>
rect 253 58 254 59 
<< m1 >>
rect 254 58 255 59 
<< m1 >>
rect 255 58 256 59 
<< m1 >>
rect 256 58 257 59 
<< m1 >>
rect 257 58 258 59 
<< m1 >>
rect 258 58 259 59 
<< m1 >>
rect 259 58 260 59 
<< m1 >>
rect 260 58 261 59 
<< m1 >>
rect 262 58 263 59 
<< m1 >>
rect 265 58 266 59 
<< m1 >>
rect 271 58 272 59 
<< m1 >>
rect 273 58 274 59 
<< m2 >>
rect 274 58 275 59 
<< m1 >>
rect 277 58 278 59 
<< m1 >>
rect 280 58 281 59 
<< m1 >>
rect 307 58 308 59 
<< m1 >>
rect 316 58 317 59 
<< m1 >>
rect 327 58 328 59 
<< m1 >>
rect 334 58 335 59 
<< m2 >>
rect 334 58 335 59 
<< m1 >>
rect 343 58 344 59 
<< m1 >>
rect 19 59 20 60 
<< m2 >>
rect 19 59 20 60 
<< m2c >>
rect 19 59 20 60 
<< m1 >>
rect 19 59 20 60 
<< m2 >>
rect 19 59 20 60 
<< m1 >>
rect 21 59 22 60 
<< m2 >>
rect 21 59 22 60 
<< m2c >>
rect 21 59 22 60 
<< m1 >>
rect 21 59 22 60 
<< m2 >>
rect 21 59 22 60 
<< m1 >>
rect 23 59 24 60 
<< m2 >>
rect 23 59 24 60 
<< m2c >>
rect 23 59 24 60 
<< m1 >>
rect 23 59 24 60 
<< m2 >>
rect 23 59 24 60 
<< m1 >>
rect 35 59 36 60 
<< m2 >>
rect 35 59 36 60 
<< m2c >>
rect 35 59 36 60 
<< m1 >>
rect 35 59 36 60 
<< m2 >>
rect 35 59 36 60 
<< m1 >>
rect 37 59 38 60 
<< m2 >>
rect 37 59 38 60 
<< m2c >>
rect 37 59 38 60 
<< m1 >>
rect 37 59 38 60 
<< m2 >>
rect 37 59 38 60 
<< m1 >>
rect 46 59 47 60 
<< m2 >>
rect 46 59 47 60 
<< m2c >>
rect 46 59 47 60 
<< m1 >>
rect 46 59 47 60 
<< m2 >>
rect 46 59 47 60 
<< m1 >>
rect 55 59 56 60 
<< m2 >>
rect 55 59 56 60 
<< m2c >>
rect 55 59 56 60 
<< m1 >>
rect 55 59 56 60 
<< m2 >>
rect 55 59 56 60 
<< m1 >>
rect 60 59 61 60 
<< m2 >>
rect 60 59 61 60 
<< m2c >>
rect 60 59 61 60 
<< m1 >>
rect 60 59 61 60 
<< m2 >>
rect 60 59 61 60 
<< m1 >>
rect 62 59 63 60 
<< m2 >>
rect 62 59 63 60 
<< m2c >>
rect 62 59 63 60 
<< m1 >>
rect 62 59 63 60 
<< m2 >>
rect 62 59 63 60 
<< m1 >>
rect 63 59 64 60 
<< m1 >>
rect 64 59 65 60 
<< m2 >>
rect 64 59 65 60 
<< m1 >>
rect 65 59 66 60 
<< m1 >>
rect 66 59 67 60 
<< m1 >>
rect 67 59 68 60 
<< m1 >>
rect 68 59 69 60 
<< m1 >>
rect 73 59 74 60 
<< m2 >>
rect 73 59 74 60 
<< m2c >>
rect 73 59 74 60 
<< m1 >>
rect 73 59 74 60 
<< m2 >>
rect 73 59 74 60 
<< m1 >>
rect 75 59 76 60 
<< m2 >>
rect 75 59 76 60 
<< m2c >>
rect 75 59 76 60 
<< m1 >>
rect 75 59 76 60 
<< m2 >>
rect 75 59 76 60 
<< m1 >>
rect 78 59 79 60 
<< m2 >>
rect 78 59 79 60 
<< m2c >>
rect 78 59 79 60 
<< m1 >>
rect 78 59 79 60 
<< m2 >>
rect 78 59 79 60 
<< m1 >>
rect 82 59 83 60 
<< m2 >>
rect 82 59 83 60 
<< m2c >>
rect 82 59 83 60 
<< m1 >>
rect 82 59 83 60 
<< m2 >>
rect 82 59 83 60 
<< m2 >>
rect 90 59 91 60 
<< m1 >>
rect 91 59 92 60 
<< m2 >>
rect 92 59 93 60 
<< m2 >>
rect 95 59 96 60 
<< m2 >>
rect 97 59 98 60 
<< m1 >>
rect 196 59 197 60 
<< m1 >>
rect 200 59 201 60 
<< m2 >>
rect 200 59 201 60 
<< m2c >>
rect 200 59 201 60 
<< m1 >>
rect 200 59 201 60 
<< m2 >>
rect 200 59 201 60 
<< m1 >>
rect 204 59 205 60 
<< m2 >>
rect 204 59 205 60 
<< m2c >>
rect 204 59 205 60 
<< m1 >>
rect 204 59 205 60 
<< m2 >>
rect 204 59 205 60 
<< m2 >>
rect 220 59 221 60 
<< m2 >>
rect 226 59 227 60 
<< m1 >>
rect 260 59 261 60 
<< m1 >>
rect 262 59 263 60 
<< m1 >>
rect 265 59 266 60 
<< m1 >>
rect 271 59 272 60 
<< m1 >>
rect 273 59 274 60 
<< m2 >>
rect 274 59 275 60 
<< m1 >>
rect 277 59 278 60 
<< m1 >>
rect 280 59 281 60 
<< m1 >>
rect 307 59 308 60 
<< m1 >>
rect 316 59 317 60 
<< m1 >>
rect 327 59 328 60 
<< m1 >>
rect 334 59 335 60 
<< m2 >>
rect 334 59 335 60 
<< m1 >>
rect 343 59 344 60 
<< m2 >>
rect 19 60 20 61 
<< m2 >>
rect 21 60 22 61 
<< m2 >>
rect 23 60 24 61 
<< m2 >>
rect 30 60 31 61 
<< m2 >>
rect 31 60 32 61 
<< m2 >>
rect 32 60 33 61 
<< m2 >>
rect 33 60 34 61 
<< m2 >>
rect 34 60 35 61 
<< m2 >>
rect 35 60 36 61 
<< m2 >>
rect 37 60 38 61 
<< m2 >>
rect 46 60 47 61 
<< m2 >>
rect 55 60 56 61 
<< m2 >>
rect 60 60 61 61 
<< m2 >>
rect 62 60 63 61 
<< m2 >>
rect 64 60 65 61 
<< m2 >>
rect 73 60 74 61 
<< m2 >>
rect 75 60 76 61 
<< m2 >>
rect 78 60 79 61 
<< m2 >>
rect 82 60 83 61 
<< m2 >>
rect 90 60 91 61 
<< m1 >>
rect 91 60 92 61 
<< m2 >>
rect 92 60 93 61 
<< m1 >>
rect 95 60 96 61 
<< m2 >>
rect 95 60 96 61 
<< m2c >>
rect 95 60 96 61 
<< m1 >>
rect 95 60 96 61 
<< m2 >>
rect 95 60 96 61 
<< m1 >>
rect 96 60 97 61 
<< m1 >>
rect 97 60 98 61 
<< m2 >>
rect 97 60 98 61 
<< m1 >>
rect 98 60 99 61 
<< m2 >>
rect 98 60 99 61 
<< m1 >>
rect 99 60 100 61 
<< m2 >>
rect 99 60 100 61 
<< m1 >>
rect 100 60 101 61 
<< m2 >>
rect 100 60 101 61 
<< m1 >>
rect 101 60 102 61 
<< m2 >>
rect 101 60 102 61 
<< m1 >>
rect 102 60 103 61 
<< m2 >>
rect 102 60 103 61 
<< m1 >>
rect 103 60 104 61 
<< m2 >>
rect 103 60 104 61 
<< m1 >>
rect 104 60 105 61 
<< m2 >>
rect 104 60 105 61 
<< m1 >>
rect 105 60 106 61 
<< m2 >>
rect 105 60 106 61 
<< m1 >>
rect 106 60 107 61 
<< m2 >>
rect 106 60 107 61 
<< m1 >>
rect 107 60 108 61 
<< m2 >>
rect 107 60 108 61 
<< m1 >>
rect 108 60 109 61 
<< m2 >>
rect 108 60 109 61 
<< m1 >>
rect 109 60 110 61 
<< m2 >>
rect 109 60 110 61 
<< m1 >>
rect 110 60 111 61 
<< m2 >>
rect 110 60 111 61 
<< m1 >>
rect 111 60 112 61 
<< m2 >>
rect 111 60 112 61 
<< m1 >>
rect 112 60 113 61 
<< m2 >>
rect 112 60 113 61 
<< m1 >>
rect 113 60 114 61 
<< m2 >>
rect 113 60 114 61 
<< m1 >>
rect 114 60 115 61 
<< m2 >>
rect 114 60 115 61 
<< m1 >>
rect 115 60 116 61 
<< m2 >>
rect 115 60 116 61 
<< m1 >>
rect 116 60 117 61 
<< m2 >>
rect 116 60 117 61 
<< m1 >>
rect 117 60 118 61 
<< m2 >>
rect 117 60 118 61 
<< m1 >>
rect 118 60 119 61 
<< m2 >>
rect 118 60 119 61 
<< m1 >>
rect 119 60 120 61 
<< m2 >>
rect 119 60 120 61 
<< m1 >>
rect 120 60 121 61 
<< m2 >>
rect 120 60 121 61 
<< m1 >>
rect 121 60 122 61 
<< m2 >>
rect 121 60 122 61 
<< m1 >>
rect 122 60 123 61 
<< m2 >>
rect 122 60 123 61 
<< m1 >>
rect 123 60 124 61 
<< m2 >>
rect 123 60 124 61 
<< m1 >>
rect 124 60 125 61 
<< m2 >>
rect 124 60 125 61 
<< m2 >>
rect 125 60 126 61 
<< m1 >>
rect 126 60 127 61 
<< m2 >>
rect 126 60 127 61 
<< m2c >>
rect 126 60 127 61 
<< m1 >>
rect 126 60 127 61 
<< m2 >>
rect 126 60 127 61 
<< m1 >>
rect 127 60 128 61 
<< m1 >>
rect 128 60 129 61 
<< m1 >>
rect 129 60 130 61 
<< m1 >>
rect 130 60 131 61 
<< m1 >>
rect 131 60 132 61 
<< m1 >>
rect 132 60 133 61 
<< m1 >>
rect 133 60 134 61 
<< m1 >>
rect 134 60 135 61 
<< m1 >>
rect 135 60 136 61 
<< m1 >>
rect 136 60 137 61 
<< m1 >>
rect 137 60 138 61 
<< m1 >>
rect 138 60 139 61 
<< m1 >>
rect 139 60 140 61 
<< m1 >>
rect 140 60 141 61 
<< m1 >>
rect 141 60 142 61 
<< m1 >>
rect 142 60 143 61 
<< m1 >>
rect 143 60 144 61 
<< m1 >>
rect 144 60 145 61 
<< m1 >>
rect 145 60 146 61 
<< m1 >>
rect 146 60 147 61 
<< m1 >>
rect 147 60 148 61 
<< m1 >>
rect 148 60 149 61 
<< m1 >>
rect 149 60 150 61 
<< m1 >>
rect 150 60 151 61 
<< m1 >>
rect 151 60 152 61 
<< m1 >>
rect 152 60 153 61 
<< m1 >>
rect 153 60 154 61 
<< m1 >>
rect 154 60 155 61 
<< m1 >>
rect 155 60 156 61 
<< m1 >>
rect 156 60 157 61 
<< m1 >>
rect 157 60 158 61 
<< m1 >>
rect 158 60 159 61 
<< m1 >>
rect 159 60 160 61 
<< m1 >>
rect 160 60 161 61 
<< m1 >>
rect 161 60 162 61 
<< m1 >>
rect 162 60 163 61 
<< m1 >>
rect 163 60 164 61 
<< m1 >>
rect 164 60 165 61 
<< m1 >>
rect 165 60 166 61 
<< m1 >>
rect 166 60 167 61 
<< m1 >>
rect 167 60 168 61 
<< m1 >>
rect 168 60 169 61 
<< m1 >>
rect 169 60 170 61 
<< m1 >>
rect 170 60 171 61 
<< m1 >>
rect 171 60 172 61 
<< m1 >>
rect 172 60 173 61 
<< m1 >>
rect 173 60 174 61 
<< m1 >>
rect 174 60 175 61 
<< m1 >>
rect 175 60 176 61 
<< m1 >>
rect 176 60 177 61 
<< m1 >>
rect 177 60 178 61 
<< m1 >>
rect 178 60 179 61 
<< m1 >>
rect 179 60 180 61 
<< m1 >>
rect 180 60 181 61 
<< m1 >>
rect 181 60 182 61 
<< m1 >>
rect 182 60 183 61 
<< m1 >>
rect 183 60 184 61 
<< m1 >>
rect 184 60 185 61 
<< m1 >>
rect 185 60 186 61 
<< m1 >>
rect 186 60 187 61 
<< m1 >>
rect 187 60 188 61 
<< m1 >>
rect 188 60 189 61 
<< m1 >>
rect 189 60 190 61 
<< m1 >>
rect 190 60 191 61 
<< m1 >>
rect 191 60 192 61 
<< m1 >>
rect 192 60 193 61 
<< m1 >>
rect 193 60 194 61 
<< m1 >>
rect 194 60 195 61 
<< m2 >>
rect 194 60 195 61 
<< m2c >>
rect 194 60 195 61 
<< m1 >>
rect 194 60 195 61 
<< m2 >>
rect 194 60 195 61 
<< m2 >>
rect 195 60 196 61 
<< m1 >>
rect 196 60 197 61 
<< m2 >>
rect 196 60 197 61 
<< m2 >>
rect 197 60 198 61 
<< m1 >>
rect 198 60 199 61 
<< m2 >>
rect 198 60 199 61 
<< m2c >>
rect 198 60 199 61 
<< m1 >>
rect 198 60 199 61 
<< m2 >>
rect 198 60 199 61 
<< m1 >>
rect 200 60 201 61 
<< m2 >>
rect 204 60 205 61 
<< m2 >>
rect 205 60 206 61 
<< m2 >>
rect 206 60 207 61 
<< m2 >>
rect 207 60 208 61 
<< m2 >>
rect 208 60 209 61 
<< m2 >>
rect 209 60 210 61 
<< m2 >>
rect 210 60 211 61 
<< m2 >>
rect 211 60 212 61 
<< m2 >>
rect 212 60 213 61 
<< m2 >>
rect 220 60 221 61 
<< m1 >>
rect 224 60 225 61 
<< m1 >>
rect 225 60 226 61 
<< m1 >>
rect 226 60 227 61 
<< m2 >>
rect 226 60 227 61 
<< m2c >>
rect 226 60 227 61 
<< m1 >>
rect 226 60 227 61 
<< m2 >>
rect 226 60 227 61 
<< m1 >>
rect 260 60 261 61 
<< m1 >>
rect 262 60 263 61 
<< m1 >>
rect 265 60 266 61 
<< m1 >>
rect 271 60 272 61 
<< m1 >>
rect 273 60 274 61 
<< m2 >>
rect 274 60 275 61 
<< m1 >>
rect 277 60 278 61 
<< m1 >>
rect 280 60 281 61 
<< m1 >>
rect 307 60 308 61 
<< m1 >>
rect 316 60 317 61 
<< m1 >>
rect 327 60 328 61 
<< m1 >>
rect 334 60 335 61 
<< m2 >>
rect 334 60 335 61 
<< m1 >>
rect 343 60 344 61 
<< m1 >>
rect 19 61 20 62 
<< m2 >>
rect 19 61 20 62 
<< m1 >>
rect 20 61 21 62 
<< m1 >>
rect 21 61 22 62 
<< m2 >>
rect 21 61 22 62 
<< m1 >>
rect 22 61 23 62 
<< m1 >>
rect 23 61 24 62 
<< m2 >>
rect 23 61 24 62 
<< m1 >>
rect 24 61 25 62 
<< m1 >>
rect 25 61 26 62 
<< m1 >>
rect 26 61 27 62 
<< m1 >>
rect 27 61 28 62 
<< m1 >>
rect 28 61 29 62 
<< m1 >>
rect 29 61 30 62 
<< m1 >>
rect 30 61 31 62 
<< m2 >>
rect 30 61 31 62 
<< m1 >>
rect 31 61 32 62 
<< m1 >>
rect 32 61 33 62 
<< m1 >>
rect 33 61 34 62 
<< m1 >>
rect 34 61 35 62 
<< m1 >>
rect 35 61 36 62 
<< m1 >>
rect 36 61 37 62 
<< m1 >>
rect 37 61 38 62 
<< m2 >>
rect 37 61 38 62 
<< m1 >>
rect 38 61 39 62 
<< m1 >>
rect 39 61 40 62 
<< m1 >>
rect 40 61 41 62 
<< m1 >>
rect 41 61 42 62 
<< m1 >>
rect 42 61 43 62 
<< m1 >>
rect 43 61 44 62 
<< m1 >>
rect 44 61 45 62 
<< m1 >>
rect 45 61 46 62 
<< m1 >>
rect 46 61 47 62 
<< m2 >>
rect 46 61 47 62 
<< m1 >>
rect 47 61 48 62 
<< m1 >>
rect 48 61 49 62 
<< m1 >>
rect 49 61 50 62 
<< m1 >>
rect 50 61 51 62 
<< m1 >>
rect 51 61 52 62 
<< m1 >>
rect 52 61 53 62 
<< m1 >>
rect 53 61 54 62 
<< m1 >>
rect 54 61 55 62 
<< m1 >>
rect 55 61 56 62 
<< m2 >>
rect 55 61 56 62 
<< m1 >>
rect 56 61 57 62 
<< m1 >>
rect 57 61 58 62 
<< m1 >>
rect 58 61 59 62 
<< m1 >>
rect 59 61 60 62 
<< m1 >>
rect 60 61 61 62 
<< m2 >>
rect 60 61 61 62 
<< m1 >>
rect 61 61 62 62 
<< m1 >>
rect 62 61 63 62 
<< m2 >>
rect 62 61 63 62 
<< m1 >>
rect 63 61 64 62 
<< m1 >>
rect 64 61 65 62 
<< m2 >>
rect 64 61 65 62 
<< m1 >>
rect 65 61 66 62 
<< m1 >>
rect 66 61 67 62 
<< m1 >>
rect 67 61 68 62 
<< m1 >>
rect 68 61 69 62 
<< m1 >>
rect 69 61 70 62 
<< m1 >>
rect 70 61 71 62 
<< m1 >>
rect 71 61 72 62 
<< m1 >>
rect 72 61 73 62 
<< m1 >>
rect 73 61 74 62 
<< m2 >>
rect 73 61 74 62 
<< m1 >>
rect 74 61 75 62 
<< m1 >>
rect 75 61 76 62 
<< m2 >>
rect 75 61 76 62 
<< m1 >>
rect 76 61 77 62 
<< m1 >>
rect 77 61 78 62 
<< m1 >>
rect 78 61 79 62 
<< m2 >>
rect 78 61 79 62 
<< m1 >>
rect 79 61 80 62 
<< m1 >>
rect 80 61 81 62 
<< m1 >>
rect 81 61 82 62 
<< m1 >>
rect 82 61 83 62 
<< m2 >>
rect 82 61 83 62 
<< m1 >>
rect 83 61 84 62 
<< m1 >>
rect 84 61 85 62 
<< m1 >>
rect 85 61 86 62 
<< m1 >>
rect 86 61 87 62 
<< m1 >>
rect 87 61 88 62 
<< m1 >>
rect 88 61 89 62 
<< m1 >>
rect 89 61 90 62 
<< m2 >>
rect 89 61 90 62 
<< m2c >>
rect 89 61 90 62 
<< m1 >>
rect 89 61 90 62 
<< m2 >>
rect 89 61 90 62 
<< m2 >>
rect 90 61 91 62 
<< m1 >>
rect 91 61 92 62 
<< m2 >>
rect 92 61 93 62 
<< m1 >>
rect 124 61 125 62 
<< m2 >>
rect 154 61 155 62 
<< m2 >>
rect 155 61 156 62 
<< m2 >>
rect 156 61 157 62 
<< m2 >>
rect 157 61 158 62 
<< m2 >>
rect 158 61 159 62 
<< m1 >>
rect 196 61 197 62 
<< m1 >>
rect 198 61 199 62 
<< m2 >>
rect 198 61 199 62 
<< m2 >>
rect 199 61 200 62 
<< m1 >>
rect 200 61 201 62 
<< m2 >>
rect 200 61 201 62 
<< m2 >>
rect 201 61 202 62 
<< m1 >>
rect 202 61 203 62 
<< m2 >>
rect 202 61 203 62 
<< m2c >>
rect 202 61 203 62 
<< m1 >>
rect 202 61 203 62 
<< m2 >>
rect 202 61 203 62 
<< m1 >>
rect 203 61 204 62 
<< m1 >>
rect 204 61 205 62 
<< m1 >>
rect 205 61 206 62 
<< m1 >>
rect 206 61 207 62 
<< m1 >>
rect 207 61 208 62 
<< m1 >>
rect 208 61 209 62 
<< m1 >>
rect 209 61 210 62 
<< m1 >>
rect 210 61 211 62 
<< m1 >>
rect 211 61 212 62 
<< m1 >>
rect 212 61 213 62 
<< m2 >>
rect 212 61 213 62 
<< m1 >>
rect 213 61 214 62 
<< m1 >>
rect 214 61 215 62 
<< m1 >>
rect 215 61 216 62 
<< m1 >>
rect 216 61 217 62 
<< m1 >>
rect 217 61 218 62 
<< m1 >>
rect 218 61 219 62 
<< m1 >>
rect 219 61 220 62 
<< m1 >>
rect 220 61 221 62 
<< m2 >>
rect 220 61 221 62 
<< m1 >>
rect 221 61 222 62 
<< m1 >>
rect 222 61 223 62 
<< m2 >>
rect 222 61 223 62 
<< m2c >>
rect 222 61 223 62 
<< m1 >>
rect 222 61 223 62 
<< m2 >>
rect 222 61 223 62 
<< m2 >>
rect 223 61 224 62 
<< m1 >>
rect 224 61 225 62 
<< m1 >>
rect 229 61 230 62 
<< m1 >>
rect 230 61 231 62 
<< m1 >>
rect 231 61 232 62 
<< m1 >>
rect 232 61 233 62 
<< m1 >>
rect 233 61 234 62 
<< m1 >>
rect 234 61 235 62 
<< m1 >>
rect 235 61 236 62 
<< m1 >>
rect 236 61 237 62 
<< m1 >>
rect 237 61 238 62 
<< m1 >>
rect 238 61 239 62 
<< m1 >>
rect 239 61 240 62 
<< m1 >>
rect 240 61 241 62 
<< m1 >>
rect 241 61 242 62 
<< m1 >>
rect 242 61 243 62 
<< m1 >>
rect 243 61 244 62 
<< m1 >>
rect 244 61 245 62 
<< m1 >>
rect 245 61 246 62 
<< m1 >>
rect 246 61 247 62 
<< m1 >>
rect 247 61 248 62 
<< m1 >>
rect 248 61 249 62 
<< m1 >>
rect 249 61 250 62 
<< m1 >>
rect 250 61 251 62 
<< m1 >>
rect 251 61 252 62 
<< m1 >>
rect 252 61 253 62 
<< m1 >>
rect 253 61 254 62 
<< m1 >>
rect 260 61 261 62 
<< m1 >>
rect 262 61 263 62 
<< m1 >>
rect 264 61 265 62 
<< m1 >>
rect 265 61 266 62 
<< m1 >>
rect 271 61 272 62 
<< m1 >>
rect 273 61 274 62 
<< m2 >>
rect 274 61 275 62 
<< m1 >>
rect 277 61 278 62 
<< m1 >>
rect 280 61 281 62 
<< m1 >>
rect 307 61 308 62 
<< m1 >>
rect 316 61 317 62 
<< m1 >>
rect 327 61 328 62 
<< m1 >>
rect 334 61 335 62 
<< m2 >>
rect 334 61 335 62 
<< m1 >>
rect 343 61 344 62 
<< m1 >>
rect 19 62 20 63 
<< m2 >>
rect 19 62 20 63 
<< m2 >>
rect 21 62 22 63 
<< m2 >>
rect 23 62 24 63 
<< m2 >>
rect 30 62 31 63 
<< m2 >>
rect 37 62 38 63 
<< m2 >>
rect 46 62 47 63 
<< m2 >>
rect 55 62 56 63 
<< m2 >>
rect 60 62 61 63 
<< m2 >>
rect 62 62 63 63 
<< m2 >>
rect 64 62 65 63 
<< m2 >>
rect 73 62 74 63 
<< m2 >>
rect 75 62 76 63 
<< m2 >>
rect 78 62 79 63 
<< m2 >>
rect 82 62 83 63 
<< m1 >>
rect 91 62 92 63 
<< m2 >>
rect 92 62 93 63 
<< m1 >>
rect 124 62 125 63 
<< m1 >>
rect 154 62 155 63 
<< m2 >>
rect 154 62 155 63 
<< m2c >>
rect 154 62 155 63 
<< m1 >>
rect 154 62 155 63 
<< m2 >>
rect 154 62 155 63 
<< m1 >>
rect 158 62 159 63 
<< m2 >>
rect 158 62 159 63 
<< m2c >>
rect 158 62 159 63 
<< m1 >>
rect 158 62 159 63 
<< m2 >>
rect 158 62 159 63 
<< m1 >>
rect 159 62 160 63 
<< m1 >>
rect 160 62 161 63 
<< m1 >>
rect 161 62 162 63 
<< m1 >>
rect 162 62 163 63 
<< m1 >>
rect 163 62 164 63 
<< m1 >>
rect 164 62 165 63 
<< m1 >>
rect 165 62 166 63 
<< m1 >>
rect 166 62 167 63 
<< m1 >>
rect 167 62 168 63 
<< m1 >>
rect 168 62 169 63 
<< m1 >>
rect 169 62 170 63 
<< m1 >>
rect 170 62 171 63 
<< m1 >>
rect 171 62 172 63 
<< m2 >>
rect 171 62 172 63 
<< m2c >>
rect 171 62 172 63 
<< m1 >>
rect 171 62 172 63 
<< m2 >>
rect 171 62 172 63 
<< m1 >>
rect 196 62 197 63 
<< m1 >>
rect 200 62 201 63 
<< m2 >>
rect 212 62 213 63 
<< m2 >>
rect 220 62 221 63 
<< m2 >>
rect 223 62 224 63 
<< m1 >>
rect 224 62 225 63 
<< m2 >>
rect 224 62 225 63 
<< m2 >>
rect 225 62 226 63 
<< m1 >>
rect 226 62 227 63 
<< m2 >>
rect 226 62 227 63 
<< m2c >>
rect 226 62 227 63 
<< m1 >>
rect 226 62 227 63 
<< m2 >>
rect 226 62 227 63 
<< m1 >>
rect 229 62 230 63 
<< m1 >>
rect 253 62 254 63 
<< m1 >>
rect 260 62 261 63 
<< m1 >>
rect 262 62 263 63 
<< m1 >>
rect 264 62 265 63 
<< m1 >>
rect 271 62 272 63 
<< m1 >>
rect 273 62 274 63 
<< m2 >>
rect 274 62 275 63 
<< m1 >>
rect 277 62 278 63 
<< m1 >>
rect 280 62 281 63 
<< m1 >>
rect 307 62 308 63 
<< m1 >>
rect 316 62 317 63 
<< m1 >>
rect 327 62 328 63 
<< m1 >>
rect 334 62 335 63 
<< m2 >>
rect 334 62 335 63 
<< m1 >>
rect 343 62 344 63 
<< m1 >>
rect 19 63 20 64 
<< m2 >>
rect 19 63 20 64 
<< m1 >>
rect 21 63 22 64 
<< m2 >>
rect 21 63 22 64 
<< m2c >>
rect 21 63 22 64 
<< m1 >>
rect 21 63 22 64 
<< m2 >>
rect 21 63 22 64 
<< m1 >>
rect 23 63 24 64 
<< m2 >>
rect 23 63 24 64 
<< m2c >>
rect 23 63 24 64 
<< m1 >>
rect 23 63 24 64 
<< m2 >>
rect 23 63 24 64 
<< m1 >>
rect 28 63 29 64 
<< m1 >>
rect 29 63 30 64 
<< m1 >>
rect 30 63 31 64 
<< m2 >>
rect 30 63 31 64 
<< m2c >>
rect 30 63 31 64 
<< m1 >>
rect 30 63 31 64 
<< m2 >>
rect 30 63 31 64 
<< m1 >>
rect 37 63 38 64 
<< m2 >>
rect 37 63 38 64 
<< m2c >>
rect 37 63 38 64 
<< m1 >>
rect 37 63 38 64 
<< m2 >>
rect 37 63 38 64 
<< m1 >>
rect 46 63 47 64 
<< m2 >>
rect 46 63 47 64 
<< m2c >>
rect 46 63 47 64 
<< m1 >>
rect 46 63 47 64 
<< m2 >>
rect 46 63 47 64 
<< m1 >>
rect 55 63 56 64 
<< m2 >>
rect 55 63 56 64 
<< m2c >>
rect 55 63 56 64 
<< m1 >>
rect 55 63 56 64 
<< m2 >>
rect 55 63 56 64 
<< m1 >>
rect 60 63 61 64 
<< m2 >>
rect 60 63 61 64 
<< m2c >>
rect 60 63 61 64 
<< m1 >>
rect 60 63 61 64 
<< m2 >>
rect 60 63 61 64 
<< m1 >>
rect 62 63 63 64 
<< m2 >>
rect 62 63 63 64 
<< m2c >>
rect 62 63 63 64 
<< m1 >>
rect 62 63 63 64 
<< m2 >>
rect 62 63 63 64 
<< m1 >>
rect 64 63 65 64 
<< m2 >>
rect 64 63 65 64 
<< m2c >>
rect 64 63 65 64 
<< m1 >>
rect 64 63 65 64 
<< m2 >>
rect 64 63 65 64 
<< m1 >>
rect 73 63 74 64 
<< m2 >>
rect 73 63 74 64 
<< m2c >>
rect 73 63 74 64 
<< m1 >>
rect 73 63 74 64 
<< m2 >>
rect 73 63 74 64 
<< m1 >>
rect 75 63 76 64 
<< m2 >>
rect 75 63 76 64 
<< m2c >>
rect 75 63 76 64 
<< m1 >>
rect 75 63 76 64 
<< m2 >>
rect 75 63 76 64 
<< m1 >>
rect 78 63 79 64 
<< m2 >>
rect 78 63 79 64 
<< m2c >>
rect 78 63 79 64 
<< m1 >>
rect 78 63 79 64 
<< m2 >>
rect 78 63 79 64 
<< m1 >>
rect 82 63 83 64 
<< m2 >>
rect 82 63 83 64 
<< m2c >>
rect 82 63 83 64 
<< m1 >>
rect 82 63 83 64 
<< m2 >>
rect 82 63 83 64 
<< m1 >>
rect 91 63 92 64 
<< m2 >>
rect 92 63 93 64 
<< m1 >>
rect 103 63 104 64 
<< m1 >>
rect 104 63 105 64 
<< m1 >>
rect 105 63 106 64 
<< m1 >>
rect 106 63 107 64 
<< m1 >>
rect 107 63 108 64 
<< m1 >>
rect 108 63 109 64 
<< m1 >>
rect 109 63 110 64 
<< m1 >>
rect 110 63 111 64 
<< m1 >>
rect 111 63 112 64 
<< m1 >>
rect 112 63 113 64 
<< m1 >>
rect 113 63 114 64 
<< m1 >>
rect 114 63 115 64 
<< m1 >>
rect 115 63 116 64 
<< m1 >>
rect 116 63 117 64 
<< m1 >>
rect 117 63 118 64 
<< m1 >>
rect 118 63 119 64 
<< m1 >>
rect 124 63 125 64 
<< m1 >>
rect 154 63 155 64 
<< m2 >>
rect 171 63 172 64 
<< m1 >>
rect 196 63 197 64 
<< m1 >>
rect 200 63 201 64 
<< m1 >>
rect 212 63 213 64 
<< m2 >>
rect 212 63 213 64 
<< m2c >>
rect 212 63 213 64 
<< m1 >>
rect 212 63 213 64 
<< m2 >>
rect 212 63 213 64 
<< m1 >>
rect 213 63 214 64 
<< m1 >>
rect 214 63 215 64 
<< m1 >>
rect 215 63 216 64 
<< m1 >>
rect 216 63 217 64 
<< m1 >>
rect 217 63 218 64 
<< m1 >>
rect 220 63 221 64 
<< m2 >>
rect 220 63 221 64 
<< m2c >>
rect 220 63 221 64 
<< m1 >>
rect 220 63 221 64 
<< m2 >>
rect 220 63 221 64 
<< m1 >>
rect 224 63 225 64 
<< m1 >>
rect 226 63 227 64 
<< m1 >>
rect 229 63 230 64 
<< m1 >>
rect 253 63 254 64 
<< m1 >>
rect 260 63 261 64 
<< m1 >>
rect 262 63 263 64 
<< m1 >>
rect 264 63 265 64 
<< m1 >>
rect 271 63 272 64 
<< m1 >>
rect 273 63 274 64 
<< m2 >>
rect 274 63 275 64 
<< m1 >>
rect 277 63 278 64 
<< m1 >>
rect 280 63 281 64 
<< m1 >>
rect 283 63 284 64 
<< m1 >>
rect 284 63 285 64 
<< m1 >>
rect 285 63 286 64 
<< m1 >>
rect 286 63 287 64 
<< m1 >>
rect 287 63 288 64 
<< m1 >>
rect 288 63 289 64 
<< m1 >>
rect 289 63 290 64 
<< m1 >>
rect 307 63 308 64 
<< m1 >>
rect 316 63 317 64 
<< m1 >>
rect 327 63 328 64 
<< m1 >>
rect 334 63 335 64 
<< m2 >>
rect 334 63 335 64 
<< m1 >>
rect 343 63 344 64 
<< m1 >>
rect 10 64 11 65 
<< m1 >>
rect 11 64 12 65 
<< m1 >>
rect 12 64 13 65 
<< m1 >>
rect 13 64 14 65 
<< m1 >>
rect 19 64 20 65 
<< m2 >>
rect 19 64 20 65 
<< m1 >>
rect 21 64 22 65 
<< m1 >>
rect 23 64 24 65 
<< m1 >>
rect 28 64 29 65 
<< m1 >>
rect 37 64 38 65 
<< m1 >>
rect 46 64 47 65 
<< m1 >>
rect 55 64 56 65 
<< m1 >>
rect 60 64 61 65 
<< m1 >>
rect 62 64 63 65 
<< m1 >>
rect 64 64 65 65 
<< m1 >>
rect 73 64 74 65 
<< m1 >>
rect 75 64 76 65 
<< m1 >>
rect 78 64 79 65 
<< m1 >>
rect 82 64 83 65 
<< m1 >>
rect 91 64 92 65 
<< m2 >>
rect 92 64 93 65 
<< m1 >>
rect 103 64 104 65 
<< m1 >>
rect 118 64 119 65 
<< m1 >>
rect 124 64 125 65 
<< m1 >>
rect 136 64 137 65 
<< m1 >>
rect 137 64 138 65 
<< m1 >>
rect 138 64 139 65 
<< m1 >>
rect 139 64 140 65 
<< m1 >>
rect 142 64 143 65 
<< m1 >>
rect 143 64 144 65 
<< m1 >>
rect 144 64 145 65 
<< m1 >>
rect 145 64 146 65 
<< m1 >>
rect 154 64 155 65 
<< m2 >>
rect 171 64 172 65 
<< m1 >>
rect 172 64 173 65 
<< m1 >>
rect 173 64 174 65 
<< m1 >>
rect 174 64 175 65 
<< m1 >>
rect 175 64 176 65 
<< m1 >>
rect 196 64 197 65 
<< m1 >>
rect 200 64 201 65 
<< m1 >>
rect 217 64 218 65 
<< m1 >>
rect 220 64 221 65 
<< m1 >>
rect 224 64 225 65 
<< m1 >>
rect 226 64 227 65 
<< m1 >>
rect 229 64 230 65 
<< m1 >>
rect 253 64 254 65 
<< m2 >>
rect 259 64 260 65 
<< m1 >>
rect 260 64 261 65 
<< m2 >>
rect 260 64 261 65 
<< m2 >>
rect 261 64 262 65 
<< m1 >>
rect 262 64 263 65 
<< m2 >>
rect 262 64 263 65 
<< m2 >>
rect 263 64 264 65 
<< m1 >>
rect 264 64 265 65 
<< m2 >>
rect 264 64 265 65 
<< m2c >>
rect 264 64 265 65 
<< m1 >>
rect 264 64 265 65 
<< m2 >>
rect 264 64 265 65 
<< m1 >>
rect 271 64 272 65 
<< m1 >>
rect 273 64 274 65 
<< m2 >>
rect 274 64 275 65 
<< m1 >>
rect 277 64 278 65 
<< m1 >>
rect 280 64 281 65 
<< m1 >>
rect 283 64 284 65 
<< m1 >>
rect 289 64 290 65 
<< m1 >>
rect 307 64 308 65 
<< m1 >>
rect 316 64 317 65 
<< m1 >>
rect 322 64 323 65 
<< m1 >>
rect 323 64 324 65 
<< m1 >>
rect 324 64 325 65 
<< m1 >>
rect 325 64 326 65 
<< m2 >>
rect 325 64 326 65 
<< m2c >>
rect 325 64 326 65 
<< m1 >>
rect 325 64 326 65 
<< m2 >>
rect 325 64 326 65 
<< m2 >>
rect 326 64 327 65 
<< m1 >>
rect 327 64 328 65 
<< m2 >>
rect 327 64 328 65 
<< m2 >>
rect 328 64 329 65 
<< m1 >>
rect 329 64 330 65 
<< m2 >>
rect 329 64 330 65 
<< m2c >>
rect 329 64 330 65 
<< m1 >>
rect 329 64 330 65 
<< m2 >>
rect 329 64 330 65 
<< m1 >>
rect 334 64 335 65 
<< m2 >>
rect 334 64 335 65 
<< m1 >>
rect 343 64 344 65 
<< m1 >>
rect 10 65 11 66 
<< m1 >>
rect 13 65 14 66 
<< m1 >>
rect 19 65 20 66 
<< m2 >>
rect 19 65 20 66 
<< m1 >>
rect 21 65 22 66 
<< m1 >>
rect 23 65 24 66 
<< m1 >>
rect 28 65 29 66 
<< m1 >>
rect 37 65 38 66 
<< m1 >>
rect 46 65 47 66 
<< m1 >>
rect 55 65 56 66 
<< m2 >>
rect 56 65 57 66 
<< m1 >>
rect 57 65 58 66 
<< m2 >>
rect 57 65 58 66 
<< m2c >>
rect 57 65 58 66 
<< m1 >>
rect 57 65 58 66 
<< m2 >>
rect 57 65 58 66 
<< m1 >>
rect 58 65 59 66 
<< m1 >>
rect 59 65 60 66 
<< m1 >>
rect 60 65 61 66 
<< m1 >>
rect 62 65 63 66 
<< m1 >>
rect 64 65 65 66 
<< m1 >>
rect 73 65 74 66 
<< m1 >>
rect 75 65 76 66 
<< m1 >>
rect 78 65 79 66 
<< m1 >>
rect 82 65 83 66 
<< m1 >>
rect 91 65 92 66 
<< m2 >>
rect 92 65 93 66 
<< m1 >>
rect 103 65 104 66 
<< m1 >>
rect 118 65 119 66 
<< m1 >>
rect 124 65 125 66 
<< m1 >>
rect 136 65 137 66 
<< m1 >>
rect 139 65 140 66 
<< m1 >>
rect 142 65 143 66 
<< m1 >>
rect 145 65 146 66 
<< m1 >>
rect 154 65 155 66 
<< m2 >>
rect 171 65 172 66 
<< m1 >>
rect 172 65 173 66 
<< m1 >>
rect 175 65 176 66 
<< m1 >>
rect 196 65 197 66 
<< m1 >>
rect 200 65 201 66 
<< m1 >>
rect 217 65 218 66 
<< m1 >>
rect 218 65 219 66 
<< m2 >>
rect 218 65 219 66 
<< m2c >>
rect 218 65 219 66 
<< m1 >>
rect 218 65 219 66 
<< m2 >>
rect 218 65 219 66 
<< m2 >>
rect 219 65 220 66 
<< m1 >>
rect 220 65 221 66 
<< m2 >>
rect 220 65 221 66 
<< m2 >>
rect 221 65 222 66 
<< m1 >>
rect 222 65 223 66 
<< m2 >>
rect 222 65 223 66 
<< m2c >>
rect 222 65 223 66 
<< m1 >>
rect 222 65 223 66 
<< m2 >>
rect 222 65 223 66 
<< m2 >>
rect 223 65 224 66 
<< m1 >>
rect 224 65 225 66 
<< m1 >>
rect 226 65 227 66 
<< m1 >>
rect 229 65 230 66 
<< m1 >>
rect 253 65 254 66 
<< m2 >>
rect 259 65 260 66 
<< m1 >>
rect 260 65 261 66 
<< m1 >>
rect 262 65 263 66 
<< m1 >>
rect 271 65 272 66 
<< m1 >>
rect 273 65 274 66 
<< m2 >>
rect 274 65 275 66 
<< m1 >>
rect 277 65 278 66 
<< m1 >>
rect 280 65 281 66 
<< m1 >>
rect 283 65 284 66 
<< m1 >>
rect 289 65 290 66 
<< m1 >>
rect 307 65 308 66 
<< m1 >>
rect 316 65 317 66 
<< m1 >>
rect 322 65 323 66 
<< m1 >>
rect 327 65 328 66 
<< m1 >>
rect 329 65 330 66 
<< m1 >>
rect 334 65 335 66 
<< m2 >>
rect 334 65 335 66 
<< m1 >>
rect 343 65 344 66 
<< m1 >>
rect 10 66 11 67 
<< pdiffusion >>
rect 12 66 13 67 
<< m1 >>
rect 13 66 14 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< m1 >>
rect 19 66 20 67 
<< m2 >>
rect 19 66 20 67 
<< m1 >>
rect 21 66 22 67 
<< m1 >>
rect 23 66 24 67 
<< m1 >>
rect 28 66 29 67 
<< pdiffusion >>
rect 30 66 31 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< m1 >>
rect 37 66 38 67 
<< m1 >>
rect 46 66 47 67 
<< pdiffusion >>
rect 48 66 49 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 55 66 56 67 
<< m2 >>
rect 56 66 57 67 
<< m1 >>
rect 62 66 63 67 
<< m1 >>
rect 64 66 65 67 
<< pdiffusion >>
rect 66 66 67 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< m1 >>
rect 73 66 74 67 
<< m1 >>
rect 75 66 76 67 
<< m1 >>
rect 78 66 79 67 
<< m1 >>
rect 82 66 83 67 
<< pdiffusion >>
rect 84 66 85 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< m1 >>
rect 91 66 92 67 
<< m2 >>
rect 92 66 93 67 
<< pdiffusion >>
rect 102 66 103 67 
<< m1 >>
rect 103 66 104 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< m1 >>
rect 118 66 119 67 
<< pdiffusion >>
rect 120 66 121 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< m1 >>
rect 124 66 125 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< m1 >>
rect 136 66 137 67 
<< pdiffusion >>
rect 138 66 139 67 
<< m1 >>
rect 139 66 140 67 
<< pdiffusion >>
rect 139 66 140 67 
<< pdiffusion >>
rect 140 66 141 67 
<< pdiffusion >>
rect 141 66 142 67 
<< m1 >>
rect 142 66 143 67 
<< pdiffusion >>
rect 142 66 143 67 
<< pdiffusion >>
rect 143 66 144 67 
<< m1 >>
rect 145 66 146 67 
<< m1 >>
rect 154 66 155 67 
<< pdiffusion >>
rect 156 66 157 67 
<< pdiffusion >>
rect 157 66 158 67 
<< pdiffusion >>
rect 158 66 159 67 
<< pdiffusion >>
rect 159 66 160 67 
<< pdiffusion >>
rect 160 66 161 67 
<< pdiffusion >>
rect 161 66 162 67 
<< m2 >>
rect 171 66 172 67 
<< m1 >>
rect 172 66 173 67 
<< pdiffusion >>
rect 174 66 175 67 
<< m1 >>
rect 175 66 176 67 
<< pdiffusion >>
rect 175 66 176 67 
<< pdiffusion >>
rect 176 66 177 67 
<< pdiffusion >>
rect 177 66 178 67 
<< pdiffusion >>
rect 178 66 179 67 
<< pdiffusion >>
rect 179 66 180 67 
<< pdiffusion >>
rect 192 66 193 67 
<< pdiffusion >>
rect 193 66 194 67 
<< pdiffusion >>
rect 194 66 195 67 
<< pdiffusion >>
rect 195 66 196 67 
<< m1 >>
rect 196 66 197 67 
<< pdiffusion >>
rect 196 66 197 67 
<< pdiffusion >>
rect 197 66 198 67 
<< m1 >>
rect 200 66 201 67 
<< pdiffusion >>
rect 210 66 211 67 
<< pdiffusion >>
rect 211 66 212 67 
<< pdiffusion >>
rect 212 66 213 67 
<< pdiffusion >>
rect 213 66 214 67 
<< pdiffusion >>
rect 214 66 215 67 
<< pdiffusion >>
rect 215 66 216 67 
<< m1 >>
rect 220 66 221 67 
<< m2 >>
rect 223 66 224 67 
<< m1 >>
rect 224 66 225 67 
<< m1 >>
rect 226 66 227 67 
<< pdiffusion >>
rect 228 66 229 67 
<< m1 >>
rect 229 66 230 67 
<< pdiffusion >>
rect 229 66 230 67 
<< pdiffusion >>
rect 230 66 231 67 
<< pdiffusion >>
rect 231 66 232 67 
<< pdiffusion >>
rect 232 66 233 67 
<< pdiffusion >>
rect 233 66 234 67 
<< pdiffusion >>
rect 246 66 247 67 
<< pdiffusion >>
rect 247 66 248 67 
<< pdiffusion >>
rect 248 66 249 67 
<< pdiffusion >>
rect 249 66 250 67 
<< pdiffusion >>
rect 250 66 251 67 
<< pdiffusion >>
rect 251 66 252 67 
<< m1 >>
rect 253 66 254 67 
<< m2 >>
rect 259 66 260 67 
<< m1 >>
rect 260 66 261 67 
<< m1 >>
rect 262 66 263 67 
<< pdiffusion >>
rect 264 66 265 67 
<< pdiffusion >>
rect 265 66 266 67 
<< pdiffusion >>
rect 266 66 267 67 
<< pdiffusion >>
rect 267 66 268 67 
<< pdiffusion >>
rect 268 66 269 67 
<< pdiffusion >>
rect 269 66 270 67 
<< m1 >>
rect 271 66 272 67 
<< m1 >>
rect 273 66 274 67 
<< m2 >>
rect 274 66 275 67 
<< m1 >>
rect 277 66 278 67 
<< m1 >>
rect 280 66 281 67 
<< pdiffusion >>
rect 282 66 283 67 
<< m1 >>
rect 283 66 284 67 
<< pdiffusion >>
rect 283 66 284 67 
<< pdiffusion >>
rect 284 66 285 67 
<< pdiffusion >>
rect 285 66 286 67 
<< pdiffusion >>
rect 286 66 287 67 
<< pdiffusion >>
rect 287 66 288 67 
<< m1 >>
rect 289 66 290 67 
<< pdiffusion >>
rect 300 66 301 67 
<< pdiffusion >>
rect 301 66 302 67 
<< pdiffusion >>
rect 302 66 303 67 
<< pdiffusion >>
rect 303 66 304 67 
<< pdiffusion >>
rect 304 66 305 67 
<< pdiffusion >>
rect 305 66 306 67 
<< m1 >>
rect 307 66 308 67 
<< m1 >>
rect 316 66 317 67 
<< pdiffusion >>
rect 318 66 319 67 
<< pdiffusion >>
rect 319 66 320 67 
<< pdiffusion >>
rect 320 66 321 67 
<< pdiffusion >>
rect 321 66 322 67 
<< m1 >>
rect 322 66 323 67 
<< pdiffusion >>
rect 322 66 323 67 
<< pdiffusion >>
rect 323 66 324 67 
<< m1 >>
rect 327 66 328 67 
<< m1 >>
rect 329 66 330 67 
<< m1 >>
rect 334 66 335 67 
<< m2 >>
rect 334 66 335 67 
<< pdiffusion >>
rect 336 66 337 67 
<< pdiffusion >>
rect 337 66 338 67 
<< pdiffusion >>
rect 338 66 339 67 
<< pdiffusion >>
rect 339 66 340 67 
<< pdiffusion >>
rect 340 66 341 67 
<< pdiffusion >>
rect 341 66 342 67 
<< m1 >>
rect 343 66 344 67 
<< m1 >>
rect 10 67 11 68 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< m1 >>
rect 19 67 20 68 
<< m2 >>
rect 19 67 20 68 
<< m1 >>
rect 21 67 22 68 
<< m1 >>
rect 23 67 24 68 
<< m1 >>
rect 28 67 29 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< m1 >>
rect 37 67 38 68 
<< m1 >>
rect 46 67 47 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 55 67 56 68 
<< m2 >>
rect 56 67 57 68 
<< m1 >>
rect 62 67 63 68 
<< m1 >>
rect 64 67 65 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< m1 >>
rect 73 67 74 68 
<< m1 >>
rect 75 67 76 68 
<< m1 >>
rect 78 67 79 68 
<< m1 >>
rect 82 67 83 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< m1 >>
rect 91 67 92 68 
<< m2 >>
rect 92 67 93 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< m1 >>
rect 118 67 119 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< m1 >>
rect 136 67 137 68 
<< pdiffusion >>
rect 138 67 139 68 
<< pdiffusion >>
rect 139 67 140 68 
<< pdiffusion >>
rect 140 67 141 68 
<< pdiffusion >>
rect 141 67 142 68 
<< pdiffusion >>
rect 142 67 143 68 
<< pdiffusion >>
rect 143 67 144 68 
<< m1 >>
rect 145 67 146 68 
<< m1 >>
rect 154 67 155 68 
<< pdiffusion >>
rect 156 67 157 68 
<< pdiffusion >>
rect 157 67 158 68 
<< pdiffusion >>
rect 158 67 159 68 
<< pdiffusion >>
rect 159 67 160 68 
<< pdiffusion >>
rect 160 67 161 68 
<< pdiffusion >>
rect 161 67 162 68 
<< m2 >>
rect 171 67 172 68 
<< m1 >>
rect 172 67 173 68 
<< pdiffusion >>
rect 174 67 175 68 
<< pdiffusion >>
rect 175 67 176 68 
<< pdiffusion >>
rect 176 67 177 68 
<< pdiffusion >>
rect 177 67 178 68 
<< pdiffusion >>
rect 178 67 179 68 
<< pdiffusion >>
rect 179 67 180 68 
<< pdiffusion >>
rect 192 67 193 68 
<< pdiffusion >>
rect 193 67 194 68 
<< pdiffusion >>
rect 194 67 195 68 
<< pdiffusion >>
rect 195 67 196 68 
<< pdiffusion >>
rect 196 67 197 68 
<< pdiffusion >>
rect 197 67 198 68 
<< m1 >>
rect 200 67 201 68 
<< pdiffusion >>
rect 210 67 211 68 
<< pdiffusion >>
rect 211 67 212 68 
<< pdiffusion >>
rect 212 67 213 68 
<< pdiffusion >>
rect 213 67 214 68 
<< pdiffusion >>
rect 214 67 215 68 
<< pdiffusion >>
rect 215 67 216 68 
<< m1 >>
rect 220 67 221 68 
<< m2 >>
rect 223 67 224 68 
<< m1 >>
rect 224 67 225 68 
<< m1 >>
rect 226 67 227 68 
<< pdiffusion >>
rect 228 67 229 68 
<< pdiffusion >>
rect 229 67 230 68 
<< pdiffusion >>
rect 230 67 231 68 
<< pdiffusion >>
rect 231 67 232 68 
<< pdiffusion >>
rect 232 67 233 68 
<< pdiffusion >>
rect 233 67 234 68 
<< pdiffusion >>
rect 246 67 247 68 
<< pdiffusion >>
rect 247 67 248 68 
<< pdiffusion >>
rect 248 67 249 68 
<< pdiffusion >>
rect 249 67 250 68 
<< pdiffusion >>
rect 250 67 251 68 
<< pdiffusion >>
rect 251 67 252 68 
<< m1 >>
rect 253 67 254 68 
<< m2 >>
rect 259 67 260 68 
<< m1 >>
rect 260 67 261 68 
<< m1 >>
rect 262 67 263 68 
<< pdiffusion >>
rect 264 67 265 68 
<< pdiffusion >>
rect 265 67 266 68 
<< pdiffusion >>
rect 266 67 267 68 
<< pdiffusion >>
rect 267 67 268 68 
<< pdiffusion >>
rect 268 67 269 68 
<< pdiffusion >>
rect 269 67 270 68 
<< m1 >>
rect 271 67 272 68 
<< m1 >>
rect 273 67 274 68 
<< m2 >>
rect 274 67 275 68 
<< m1 >>
rect 277 67 278 68 
<< m1 >>
rect 280 67 281 68 
<< pdiffusion >>
rect 282 67 283 68 
<< pdiffusion >>
rect 283 67 284 68 
<< pdiffusion >>
rect 284 67 285 68 
<< pdiffusion >>
rect 285 67 286 68 
<< pdiffusion >>
rect 286 67 287 68 
<< pdiffusion >>
rect 287 67 288 68 
<< m1 >>
rect 289 67 290 68 
<< pdiffusion >>
rect 300 67 301 68 
<< pdiffusion >>
rect 301 67 302 68 
<< pdiffusion >>
rect 302 67 303 68 
<< pdiffusion >>
rect 303 67 304 68 
<< pdiffusion >>
rect 304 67 305 68 
<< pdiffusion >>
rect 305 67 306 68 
<< m1 >>
rect 307 67 308 68 
<< m1 >>
rect 316 67 317 68 
<< pdiffusion >>
rect 318 67 319 68 
<< pdiffusion >>
rect 319 67 320 68 
<< pdiffusion >>
rect 320 67 321 68 
<< pdiffusion >>
rect 321 67 322 68 
<< pdiffusion >>
rect 322 67 323 68 
<< pdiffusion >>
rect 323 67 324 68 
<< m1 >>
rect 327 67 328 68 
<< m1 >>
rect 329 67 330 68 
<< m1 >>
rect 334 67 335 68 
<< m2 >>
rect 334 67 335 68 
<< pdiffusion >>
rect 336 67 337 68 
<< pdiffusion >>
rect 337 67 338 68 
<< pdiffusion >>
rect 338 67 339 68 
<< pdiffusion >>
rect 339 67 340 68 
<< pdiffusion >>
rect 340 67 341 68 
<< pdiffusion >>
rect 341 67 342 68 
<< m1 >>
rect 343 67 344 68 
<< m1 >>
rect 10 68 11 69 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< m1 >>
rect 19 68 20 69 
<< m2 >>
rect 19 68 20 69 
<< m1 >>
rect 21 68 22 69 
<< m1 >>
rect 23 68 24 69 
<< m1 >>
rect 28 68 29 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< m1 >>
rect 37 68 38 69 
<< m1 >>
rect 46 68 47 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 55 68 56 69 
<< m2 >>
rect 56 68 57 69 
<< m1 >>
rect 62 68 63 69 
<< m1 >>
rect 64 68 65 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< m1 >>
rect 73 68 74 69 
<< m1 >>
rect 75 68 76 69 
<< m1 >>
rect 78 68 79 69 
<< m1 >>
rect 82 68 83 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< m1 >>
rect 91 68 92 69 
<< m2 >>
rect 92 68 93 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< m1 >>
rect 118 68 119 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< m1 >>
rect 136 68 137 69 
<< pdiffusion >>
rect 138 68 139 69 
<< pdiffusion >>
rect 139 68 140 69 
<< pdiffusion >>
rect 140 68 141 69 
<< pdiffusion >>
rect 141 68 142 69 
<< pdiffusion >>
rect 142 68 143 69 
<< pdiffusion >>
rect 143 68 144 69 
<< m1 >>
rect 145 68 146 69 
<< m1 >>
rect 154 68 155 69 
<< pdiffusion >>
rect 156 68 157 69 
<< pdiffusion >>
rect 157 68 158 69 
<< pdiffusion >>
rect 158 68 159 69 
<< pdiffusion >>
rect 159 68 160 69 
<< pdiffusion >>
rect 160 68 161 69 
<< pdiffusion >>
rect 161 68 162 69 
<< m2 >>
rect 171 68 172 69 
<< m1 >>
rect 172 68 173 69 
<< pdiffusion >>
rect 174 68 175 69 
<< pdiffusion >>
rect 175 68 176 69 
<< pdiffusion >>
rect 176 68 177 69 
<< pdiffusion >>
rect 177 68 178 69 
<< pdiffusion >>
rect 178 68 179 69 
<< pdiffusion >>
rect 179 68 180 69 
<< pdiffusion >>
rect 192 68 193 69 
<< pdiffusion >>
rect 193 68 194 69 
<< pdiffusion >>
rect 194 68 195 69 
<< pdiffusion >>
rect 195 68 196 69 
<< pdiffusion >>
rect 196 68 197 69 
<< pdiffusion >>
rect 197 68 198 69 
<< m1 >>
rect 200 68 201 69 
<< pdiffusion >>
rect 210 68 211 69 
<< pdiffusion >>
rect 211 68 212 69 
<< pdiffusion >>
rect 212 68 213 69 
<< pdiffusion >>
rect 213 68 214 69 
<< pdiffusion >>
rect 214 68 215 69 
<< pdiffusion >>
rect 215 68 216 69 
<< m1 >>
rect 220 68 221 69 
<< m2 >>
rect 223 68 224 69 
<< m1 >>
rect 224 68 225 69 
<< m1 >>
rect 226 68 227 69 
<< pdiffusion >>
rect 228 68 229 69 
<< pdiffusion >>
rect 229 68 230 69 
<< pdiffusion >>
rect 230 68 231 69 
<< pdiffusion >>
rect 231 68 232 69 
<< pdiffusion >>
rect 232 68 233 69 
<< pdiffusion >>
rect 233 68 234 69 
<< pdiffusion >>
rect 246 68 247 69 
<< pdiffusion >>
rect 247 68 248 69 
<< pdiffusion >>
rect 248 68 249 69 
<< pdiffusion >>
rect 249 68 250 69 
<< pdiffusion >>
rect 250 68 251 69 
<< pdiffusion >>
rect 251 68 252 69 
<< m1 >>
rect 253 68 254 69 
<< m2 >>
rect 259 68 260 69 
<< m1 >>
rect 260 68 261 69 
<< m1 >>
rect 262 68 263 69 
<< pdiffusion >>
rect 264 68 265 69 
<< pdiffusion >>
rect 265 68 266 69 
<< pdiffusion >>
rect 266 68 267 69 
<< pdiffusion >>
rect 267 68 268 69 
<< pdiffusion >>
rect 268 68 269 69 
<< pdiffusion >>
rect 269 68 270 69 
<< m1 >>
rect 271 68 272 69 
<< m1 >>
rect 273 68 274 69 
<< m2 >>
rect 274 68 275 69 
<< m1 >>
rect 277 68 278 69 
<< m1 >>
rect 280 68 281 69 
<< pdiffusion >>
rect 282 68 283 69 
<< pdiffusion >>
rect 283 68 284 69 
<< pdiffusion >>
rect 284 68 285 69 
<< pdiffusion >>
rect 285 68 286 69 
<< pdiffusion >>
rect 286 68 287 69 
<< pdiffusion >>
rect 287 68 288 69 
<< m1 >>
rect 289 68 290 69 
<< pdiffusion >>
rect 300 68 301 69 
<< pdiffusion >>
rect 301 68 302 69 
<< pdiffusion >>
rect 302 68 303 69 
<< pdiffusion >>
rect 303 68 304 69 
<< pdiffusion >>
rect 304 68 305 69 
<< pdiffusion >>
rect 305 68 306 69 
<< m1 >>
rect 307 68 308 69 
<< m1 >>
rect 316 68 317 69 
<< pdiffusion >>
rect 318 68 319 69 
<< pdiffusion >>
rect 319 68 320 69 
<< pdiffusion >>
rect 320 68 321 69 
<< pdiffusion >>
rect 321 68 322 69 
<< pdiffusion >>
rect 322 68 323 69 
<< pdiffusion >>
rect 323 68 324 69 
<< m1 >>
rect 327 68 328 69 
<< m1 >>
rect 329 68 330 69 
<< m1 >>
rect 334 68 335 69 
<< m2 >>
rect 334 68 335 69 
<< pdiffusion >>
rect 336 68 337 69 
<< pdiffusion >>
rect 337 68 338 69 
<< pdiffusion >>
rect 338 68 339 69 
<< pdiffusion >>
rect 339 68 340 69 
<< pdiffusion >>
rect 340 68 341 69 
<< pdiffusion >>
rect 341 68 342 69 
<< m1 >>
rect 343 68 344 69 
<< m1 >>
rect 10 69 11 70 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< m1 >>
rect 19 69 20 70 
<< m2 >>
rect 19 69 20 70 
<< m1 >>
rect 21 69 22 70 
<< m1 >>
rect 23 69 24 70 
<< m1 >>
rect 28 69 29 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< m1 >>
rect 37 69 38 70 
<< m1 >>
rect 46 69 47 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 55 69 56 70 
<< m2 >>
rect 56 69 57 70 
<< m1 >>
rect 62 69 63 70 
<< m1 >>
rect 64 69 65 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< m1 >>
rect 73 69 74 70 
<< m1 >>
rect 75 69 76 70 
<< m1 >>
rect 78 69 79 70 
<< m1 >>
rect 82 69 83 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< m1 >>
rect 91 69 92 70 
<< m2 >>
rect 92 69 93 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< m1 >>
rect 118 69 119 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< m1 >>
rect 136 69 137 70 
<< pdiffusion >>
rect 138 69 139 70 
<< pdiffusion >>
rect 139 69 140 70 
<< pdiffusion >>
rect 140 69 141 70 
<< pdiffusion >>
rect 141 69 142 70 
<< pdiffusion >>
rect 142 69 143 70 
<< pdiffusion >>
rect 143 69 144 70 
<< m1 >>
rect 145 69 146 70 
<< m1 >>
rect 154 69 155 70 
<< pdiffusion >>
rect 156 69 157 70 
<< pdiffusion >>
rect 157 69 158 70 
<< pdiffusion >>
rect 158 69 159 70 
<< pdiffusion >>
rect 159 69 160 70 
<< pdiffusion >>
rect 160 69 161 70 
<< pdiffusion >>
rect 161 69 162 70 
<< m2 >>
rect 171 69 172 70 
<< m1 >>
rect 172 69 173 70 
<< pdiffusion >>
rect 174 69 175 70 
<< pdiffusion >>
rect 175 69 176 70 
<< pdiffusion >>
rect 176 69 177 70 
<< pdiffusion >>
rect 177 69 178 70 
<< pdiffusion >>
rect 178 69 179 70 
<< pdiffusion >>
rect 179 69 180 70 
<< pdiffusion >>
rect 192 69 193 70 
<< pdiffusion >>
rect 193 69 194 70 
<< pdiffusion >>
rect 194 69 195 70 
<< pdiffusion >>
rect 195 69 196 70 
<< pdiffusion >>
rect 196 69 197 70 
<< pdiffusion >>
rect 197 69 198 70 
<< m1 >>
rect 200 69 201 70 
<< pdiffusion >>
rect 210 69 211 70 
<< pdiffusion >>
rect 211 69 212 70 
<< pdiffusion >>
rect 212 69 213 70 
<< pdiffusion >>
rect 213 69 214 70 
<< pdiffusion >>
rect 214 69 215 70 
<< pdiffusion >>
rect 215 69 216 70 
<< m1 >>
rect 220 69 221 70 
<< m2 >>
rect 223 69 224 70 
<< m1 >>
rect 224 69 225 70 
<< m1 >>
rect 226 69 227 70 
<< pdiffusion >>
rect 228 69 229 70 
<< pdiffusion >>
rect 229 69 230 70 
<< pdiffusion >>
rect 230 69 231 70 
<< pdiffusion >>
rect 231 69 232 70 
<< pdiffusion >>
rect 232 69 233 70 
<< pdiffusion >>
rect 233 69 234 70 
<< pdiffusion >>
rect 246 69 247 70 
<< pdiffusion >>
rect 247 69 248 70 
<< pdiffusion >>
rect 248 69 249 70 
<< pdiffusion >>
rect 249 69 250 70 
<< pdiffusion >>
rect 250 69 251 70 
<< pdiffusion >>
rect 251 69 252 70 
<< m1 >>
rect 253 69 254 70 
<< m2 >>
rect 259 69 260 70 
<< m1 >>
rect 260 69 261 70 
<< m1 >>
rect 262 69 263 70 
<< pdiffusion >>
rect 264 69 265 70 
<< pdiffusion >>
rect 265 69 266 70 
<< pdiffusion >>
rect 266 69 267 70 
<< pdiffusion >>
rect 267 69 268 70 
<< pdiffusion >>
rect 268 69 269 70 
<< pdiffusion >>
rect 269 69 270 70 
<< m1 >>
rect 271 69 272 70 
<< m1 >>
rect 273 69 274 70 
<< m2 >>
rect 274 69 275 70 
<< m1 >>
rect 277 69 278 70 
<< m1 >>
rect 280 69 281 70 
<< pdiffusion >>
rect 282 69 283 70 
<< pdiffusion >>
rect 283 69 284 70 
<< pdiffusion >>
rect 284 69 285 70 
<< pdiffusion >>
rect 285 69 286 70 
<< pdiffusion >>
rect 286 69 287 70 
<< pdiffusion >>
rect 287 69 288 70 
<< m1 >>
rect 289 69 290 70 
<< pdiffusion >>
rect 300 69 301 70 
<< pdiffusion >>
rect 301 69 302 70 
<< pdiffusion >>
rect 302 69 303 70 
<< pdiffusion >>
rect 303 69 304 70 
<< pdiffusion >>
rect 304 69 305 70 
<< pdiffusion >>
rect 305 69 306 70 
<< m1 >>
rect 307 69 308 70 
<< m1 >>
rect 316 69 317 70 
<< pdiffusion >>
rect 318 69 319 70 
<< pdiffusion >>
rect 319 69 320 70 
<< pdiffusion >>
rect 320 69 321 70 
<< pdiffusion >>
rect 321 69 322 70 
<< pdiffusion >>
rect 322 69 323 70 
<< pdiffusion >>
rect 323 69 324 70 
<< m1 >>
rect 327 69 328 70 
<< m1 >>
rect 329 69 330 70 
<< m1 >>
rect 334 69 335 70 
<< m2 >>
rect 334 69 335 70 
<< pdiffusion >>
rect 336 69 337 70 
<< pdiffusion >>
rect 337 69 338 70 
<< pdiffusion >>
rect 338 69 339 70 
<< pdiffusion >>
rect 339 69 340 70 
<< pdiffusion >>
rect 340 69 341 70 
<< pdiffusion >>
rect 341 69 342 70 
<< m1 >>
rect 343 69 344 70 
<< m1 >>
rect 10 70 11 71 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< m1 >>
rect 19 70 20 71 
<< m2 >>
rect 19 70 20 71 
<< m1 >>
rect 21 70 22 71 
<< m1 >>
rect 23 70 24 71 
<< m1 >>
rect 28 70 29 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< m1 >>
rect 37 70 38 71 
<< m1 >>
rect 46 70 47 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 55 70 56 71 
<< m2 >>
rect 56 70 57 71 
<< m1 >>
rect 62 70 63 71 
<< m1 >>
rect 64 70 65 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< m1 >>
rect 73 70 74 71 
<< m1 >>
rect 75 70 76 71 
<< m1 >>
rect 78 70 79 71 
<< m1 >>
rect 82 70 83 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< m1 >>
rect 91 70 92 71 
<< m2 >>
rect 92 70 93 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< m1 >>
rect 118 70 119 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< m1 >>
rect 136 70 137 71 
<< pdiffusion >>
rect 138 70 139 71 
<< pdiffusion >>
rect 139 70 140 71 
<< pdiffusion >>
rect 140 70 141 71 
<< pdiffusion >>
rect 141 70 142 71 
<< pdiffusion >>
rect 142 70 143 71 
<< pdiffusion >>
rect 143 70 144 71 
<< m1 >>
rect 145 70 146 71 
<< m1 >>
rect 154 70 155 71 
<< pdiffusion >>
rect 156 70 157 71 
<< pdiffusion >>
rect 157 70 158 71 
<< pdiffusion >>
rect 158 70 159 71 
<< pdiffusion >>
rect 159 70 160 71 
<< pdiffusion >>
rect 160 70 161 71 
<< pdiffusion >>
rect 161 70 162 71 
<< m2 >>
rect 171 70 172 71 
<< m1 >>
rect 172 70 173 71 
<< pdiffusion >>
rect 174 70 175 71 
<< pdiffusion >>
rect 175 70 176 71 
<< pdiffusion >>
rect 176 70 177 71 
<< pdiffusion >>
rect 177 70 178 71 
<< pdiffusion >>
rect 178 70 179 71 
<< pdiffusion >>
rect 179 70 180 71 
<< pdiffusion >>
rect 192 70 193 71 
<< pdiffusion >>
rect 193 70 194 71 
<< pdiffusion >>
rect 194 70 195 71 
<< pdiffusion >>
rect 195 70 196 71 
<< pdiffusion >>
rect 196 70 197 71 
<< pdiffusion >>
rect 197 70 198 71 
<< m1 >>
rect 200 70 201 71 
<< pdiffusion >>
rect 210 70 211 71 
<< pdiffusion >>
rect 211 70 212 71 
<< pdiffusion >>
rect 212 70 213 71 
<< pdiffusion >>
rect 213 70 214 71 
<< pdiffusion >>
rect 214 70 215 71 
<< pdiffusion >>
rect 215 70 216 71 
<< m1 >>
rect 220 70 221 71 
<< m2 >>
rect 223 70 224 71 
<< m1 >>
rect 224 70 225 71 
<< m1 >>
rect 226 70 227 71 
<< pdiffusion >>
rect 228 70 229 71 
<< pdiffusion >>
rect 229 70 230 71 
<< pdiffusion >>
rect 230 70 231 71 
<< pdiffusion >>
rect 231 70 232 71 
<< pdiffusion >>
rect 232 70 233 71 
<< pdiffusion >>
rect 233 70 234 71 
<< pdiffusion >>
rect 246 70 247 71 
<< pdiffusion >>
rect 247 70 248 71 
<< pdiffusion >>
rect 248 70 249 71 
<< pdiffusion >>
rect 249 70 250 71 
<< pdiffusion >>
rect 250 70 251 71 
<< pdiffusion >>
rect 251 70 252 71 
<< m1 >>
rect 253 70 254 71 
<< m2 >>
rect 259 70 260 71 
<< m1 >>
rect 260 70 261 71 
<< m1 >>
rect 262 70 263 71 
<< pdiffusion >>
rect 264 70 265 71 
<< pdiffusion >>
rect 265 70 266 71 
<< pdiffusion >>
rect 266 70 267 71 
<< pdiffusion >>
rect 267 70 268 71 
<< pdiffusion >>
rect 268 70 269 71 
<< pdiffusion >>
rect 269 70 270 71 
<< m1 >>
rect 271 70 272 71 
<< m1 >>
rect 273 70 274 71 
<< m2 >>
rect 274 70 275 71 
<< m1 >>
rect 277 70 278 71 
<< m1 >>
rect 280 70 281 71 
<< pdiffusion >>
rect 282 70 283 71 
<< pdiffusion >>
rect 283 70 284 71 
<< pdiffusion >>
rect 284 70 285 71 
<< pdiffusion >>
rect 285 70 286 71 
<< pdiffusion >>
rect 286 70 287 71 
<< pdiffusion >>
rect 287 70 288 71 
<< m1 >>
rect 289 70 290 71 
<< pdiffusion >>
rect 300 70 301 71 
<< pdiffusion >>
rect 301 70 302 71 
<< pdiffusion >>
rect 302 70 303 71 
<< pdiffusion >>
rect 303 70 304 71 
<< pdiffusion >>
rect 304 70 305 71 
<< pdiffusion >>
rect 305 70 306 71 
<< m1 >>
rect 307 70 308 71 
<< m1 >>
rect 316 70 317 71 
<< pdiffusion >>
rect 318 70 319 71 
<< pdiffusion >>
rect 319 70 320 71 
<< pdiffusion >>
rect 320 70 321 71 
<< pdiffusion >>
rect 321 70 322 71 
<< pdiffusion >>
rect 322 70 323 71 
<< pdiffusion >>
rect 323 70 324 71 
<< m1 >>
rect 327 70 328 71 
<< m1 >>
rect 329 70 330 71 
<< m1 >>
rect 334 70 335 71 
<< m2 >>
rect 334 70 335 71 
<< pdiffusion >>
rect 336 70 337 71 
<< pdiffusion >>
rect 337 70 338 71 
<< pdiffusion >>
rect 338 70 339 71 
<< pdiffusion >>
rect 339 70 340 71 
<< pdiffusion >>
rect 340 70 341 71 
<< pdiffusion >>
rect 341 70 342 71 
<< m1 >>
rect 343 70 344 71 
<< m1 >>
rect 10 71 11 72 
<< pdiffusion >>
rect 12 71 13 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< m1 >>
rect 19 71 20 72 
<< m2 >>
rect 19 71 20 72 
<< m1 >>
rect 21 71 22 72 
<< m1 >>
rect 23 71 24 72 
<< m1 >>
rect 28 71 29 72 
<< pdiffusion >>
rect 30 71 31 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< m1 >>
rect 37 71 38 72 
<< m1 >>
rect 46 71 47 72 
<< pdiffusion >>
rect 48 71 49 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 55 71 56 72 
<< m2 >>
rect 56 71 57 72 
<< m1 >>
rect 62 71 63 72 
<< m1 >>
rect 64 71 65 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< m1 >>
rect 70 71 71 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< m1 >>
rect 73 71 74 72 
<< m1 >>
rect 75 71 76 72 
<< m1 >>
rect 78 71 79 72 
<< m1 >>
rect 82 71 83 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< m1 >>
rect 91 71 92 72 
<< m2 >>
rect 92 71 93 72 
<< pdiffusion >>
rect 102 71 103 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< m1 >>
rect 118 71 119 72 
<< pdiffusion >>
rect 120 71 121 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< m1 >>
rect 136 71 137 72 
<< pdiffusion >>
rect 138 71 139 72 
<< pdiffusion >>
rect 139 71 140 72 
<< pdiffusion >>
rect 140 71 141 72 
<< pdiffusion >>
rect 141 71 142 72 
<< pdiffusion >>
rect 142 71 143 72 
<< pdiffusion >>
rect 143 71 144 72 
<< m1 >>
rect 145 71 146 72 
<< m1 >>
rect 154 71 155 72 
<< pdiffusion >>
rect 156 71 157 72 
<< pdiffusion >>
rect 157 71 158 72 
<< pdiffusion >>
rect 158 71 159 72 
<< pdiffusion >>
rect 159 71 160 72 
<< m1 >>
rect 160 71 161 72 
<< pdiffusion >>
rect 160 71 161 72 
<< pdiffusion >>
rect 161 71 162 72 
<< m2 >>
rect 171 71 172 72 
<< m1 >>
rect 172 71 173 72 
<< pdiffusion >>
rect 174 71 175 72 
<< pdiffusion >>
rect 175 71 176 72 
<< pdiffusion >>
rect 176 71 177 72 
<< pdiffusion >>
rect 177 71 178 72 
<< pdiffusion >>
rect 178 71 179 72 
<< pdiffusion >>
rect 179 71 180 72 
<< pdiffusion >>
rect 192 71 193 72 
<< pdiffusion >>
rect 193 71 194 72 
<< pdiffusion >>
rect 194 71 195 72 
<< pdiffusion >>
rect 195 71 196 72 
<< pdiffusion >>
rect 196 71 197 72 
<< pdiffusion >>
rect 197 71 198 72 
<< m1 >>
rect 200 71 201 72 
<< pdiffusion >>
rect 210 71 211 72 
<< pdiffusion >>
rect 211 71 212 72 
<< pdiffusion >>
rect 212 71 213 72 
<< pdiffusion >>
rect 213 71 214 72 
<< pdiffusion >>
rect 214 71 215 72 
<< pdiffusion >>
rect 215 71 216 72 
<< m1 >>
rect 220 71 221 72 
<< m2 >>
rect 223 71 224 72 
<< m1 >>
rect 224 71 225 72 
<< m1 >>
rect 226 71 227 72 
<< pdiffusion >>
rect 228 71 229 72 
<< pdiffusion >>
rect 229 71 230 72 
<< pdiffusion >>
rect 230 71 231 72 
<< pdiffusion >>
rect 231 71 232 72 
<< pdiffusion >>
rect 232 71 233 72 
<< pdiffusion >>
rect 233 71 234 72 
<< pdiffusion >>
rect 246 71 247 72 
<< pdiffusion >>
rect 247 71 248 72 
<< pdiffusion >>
rect 248 71 249 72 
<< pdiffusion >>
rect 249 71 250 72 
<< pdiffusion >>
rect 250 71 251 72 
<< pdiffusion >>
rect 251 71 252 72 
<< m1 >>
rect 253 71 254 72 
<< m2 >>
rect 259 71 260 72 
<< m1 >>
rect 260 71 261 72 
<< m1 >>
rect 262 71 263 72 
<< pdiffusion >>
rect 264 71 265 72 
<< pdiffusion >>
rect 265 71 266 72 
<< pdiffusion >>
rect 266 71 267 72 
<< pdiffusion >>
rect 267 71 268 72 
<< pdiffusion >>
rect 268 71 269 72 
<< pdiffusion >>
rect 269 71 270 72 
<< m1 >>
rect 271 71 272 72 
<< m1 >>
rect 273 71 274 72 
<< m2 >>
rect 274 71 275 72 
<< m1 >>
rect 277 71 278 72 
<< m1 >>
rect 280 71 281 72 
<< pdiffusion >>
rect 282 71 283 72 
<< pdiffusion >>
rect 283 71 284 72 
<< pdiffusion >>
rect 284 71 285 72 
<< pdiffusion >>
rect 285 71 286 72 
<< pdiffusion >>
rect 286 71 287 72 
<< pdiffusion >>
rect 287 71 288 72 
<< m1 >>
rect 289 71 290 72 
<< pdiffusion >>
rect 300 71 301 72 
<< pdiffusion >>
rect 301 71 302 72 
<< pdiffusion >>
rect 302 71 303 72 
<< pdiffusion >>
rect 303 71 304 72 
<< m1 >>
rect 304 71 305 72 
<< pdiffusion >>
rect 304 71 305 72 
<< pdiffusion >>
rect 305 71 306 72 
<< m1 >>
rect 307 71 308 72 
<< m1 >>
rect 316 71 317 72 
<< pdiffusion >>
rect 318 71 319 72 
<< pdiffusion >>
rect 319 71 320 72 
<< pdiffusion >>
rect 320 71 321 72 
<< pdiffusion >>
rect 321 71 322 72 
<< pdiffusion >>
rect 322 71 323 72 
<< pdiffusion >>
rect 323 71 324 72 
<< m1 >>
rect 327 71 328 72 
<< m1 >>
rect 329 71 330 72 
<< m1 >>
rect 334 71 335 72 
<< m2 >>
rect 334 71 335 72 
<< pdiffusion >>
rect 336 71 337 72 
<< pdiffusion >>
rect 337 71 338 72 
<< pdiffusion >>
rect 338 71 339 72 
<< pdiffusion >>
rect 339 71 340 72 
<< pdiffusion >>
rect 340 71 341 72 
<< pdiffusion >>
rect 341 71 342 72 
<< m1 >>
rect 343 71 344 72 
<< m1 >>
rect 10 72 11 73 
<< m1 >>
rect 19 72 20 73 
<< m2 >>
rect 19 72 20 73 
<< m1 >>
rect 21 72 22 73 
<< m1 >>
rect 23 72 24 73 
<< m1 >>
rect 28 72 29 73 
<< m1 >>
rect 37 72 38 73 
<< m1 >>
rect 46 72 47 73 
<< m1 >>
rect 55 72 56 73 
<< m2 >>
rect 56 72 57 73 
<< m1 >>
rect 62 72 63 73 
<< m1 >>
rect 64 72 65 73 
<< m1 >>
rect 70 72 71 73 
<< m1 >>
rect 73 72 74 73 
<< m1 >>
rect 75 72 76 73 
<< m1 >>
rect 78 72 79 73 
<< m1 >>
rect 82 72 83 73 
<< m1 >>
rect 91 72 92 73 
<< m2 >>
rect 92 72 93 73 
<< m1 >>
rect 118 72 119 73 
<< m1 >>
rect 136 72 137 73 
<< m1 >>
rect 145 72 146 73 
<< m1 >>
rect 154 72 155 73 
<< m1 >>
rect 160 72 161 73 
<< m2 >>
rect 171 72 172 73 
<< m1 >>
rect 172 72 173 73 
<< m1 >>
rect 200 72 201 73 
<< m1 >>
rect 220 72 221 73 
<< m2 >>
rect 223 72 224 73 
<< m1 >>
rect 224 72 225 73 
<< m1 >>
rect 226 72 227 73 
<< m1 >>
rect 253 72 254 73 
<< m2 >>
rect 253 72 254 73 
<< m2c >>
rect 253 72 254 73 
<< m1 >>
rect 253 72 254 73 
<< m2 >>
rect 253 72 254 73 
<< m2 >>
rect 259 72 260 73 
<< m1 >>
rect 260 72 261 73 
<< m1 >>
rect 262 72 263 73 
<< m1 >>
rect 271 72 272 73 
<< m1 >>
rect 273 72 274 73 
<< m2 >>
rect 274 72 275 73 
<< m1 >>
rect 277 72 278 73 
<< m1 >>
rect 280 72 281 73 
<< m1 >>
rect 289 72 290 73 
<< m1 >>
rect 304 72 305 73 
<< m1 >>
rect 307 72 308 73 
<< m1 >>
rect 316 72 317 73 
<< m1 >>
rect 327 72 328 73 
<< m2 >>
rect 327 72 328 73 
<< m2c >>
rect 327 72 328 73 
<< m1 >>
rect 327 72 328 73 
<< m2 >>
rect 327 72 328 73 
<< m1 >>
rect 329 72 330 73 
<< m2 >>
rect 329 72 330 73 
<< m2c >>
rect 329 72 330 73 
<< m1 >>
rect 329 72 330 73 
<< m2 >>
rect 329 72 330 73 
<< m1 >>
rect 334 72 335 73 
<< m2 >>
rect 334 72 335 73 
<< m1 >>
rect 343 72 344 73 
<< m1 >>
rect 10 73 11 74 
<< m1 >>
rect 19 73 20 74 
<< m2 >>
rect 19 73 20 74 
<< m1 >>
rect 21 73 22 74 
<< m1 >>
rect 23 73 24 74 
<< m1 >>
rect 28 73 29 74 
<< m1 >>
rect 37 73 38 74 
<< m1 >>
rect 46 73 47 74 
<< m1 >>
rect 55 73 56 74 
<< m2 >>
rect 56 73 57 74 
<< m1 >>
rect 62 73 63 74 
<< m1 >>
rect 64 73 65 74 
<< m1 >>
rect 70 73 71 74 
<< m1 >>
rect 71 73 72 74 
<< m1 >>
rect 72 73 73 74 
<< m1 >>
rect 73 73 74 74 
<< m1 >>
rect 75 73 76 74 
<< m1 >>
rect 78 73 79 74 
<< m1 >>
rect 82 73 83 74 
<< m1 >>
rect 91 73 92 74 
<< m2 >>
rect 92 73 93 74 
<< m1 >>
rect 118 73 119 74 
<< m1 >>
rect 136 73 137 74 
<< m1 >>
rect 145 73 146 74 
<< m1 >>
rect 154 73 155 74 
<< m1 >>
rect 160 73 161 74 
<< m2 >>
rect 171 73 172 74 
<< m1 >>
rect 172 73 173 74 
<< m2 >>
rect 172 73 173 74 
<< m2 >>
rect 173 73 174 74 
<< m1 >>
rect 174 73 175 74 
<< m2 >>
rect 174 73 175 74 
<< m2c >>
rect 174 73 175 74 
<< m1 >>
rect 174 73 175 74 
<< m2 >>
rect 174 73 175 74 
<< m1 >>
rect 200 73 201 74 
<< m1 >>
rect 220 73 221 74 
<< m2 >>
rect 223 73 224 74 
<< m1 >>
rect 224 73 225 74 
<< m1 >>
rect 226 73 227 74 
<< m2 >>
rect 253 73 254 74 
<< m2 >>
rect 259 73 260 74 
<< m1 >>
rect 260 73 261 74 
<< m1 >>
rect 262 73 263 74 
<< m1 >>
rect 271 73 272 74 
<< m1 >>
rect 273 73 274 74 
<< m2 >>
rect 274 73 275 74 
<< m1 >>
rect 277 73 278 74 
<< m1 >>
rect 280 73 281 74 
<< m1 >>
rect 289 73 290 74 
<< m1 >>
rect 304 73 305 74 
<< m1 >>
rect 305 73 306 74 
<< m1 >>
rect 306 73 307 74 
<< m1 >>
rect 307 73 308 74 
<< m1 >>
rect 316 73 317 74 
<< m2 >>
rect 327 73 328 74 
<< m2 >>
rect 329 73 330 74 
<< m1 >>
rect 334 73 335 74 
<< m2 >>
rect 334 73 335 74 
<< m1 >>
rect 343 73 344 74 
<< m1 >>
rect 10 74 11 75 
<< m1 >>
rect 19 74 20 75 
<< m2 >>
rect 19 74 20 75 
<< m1 >>
rect 21 74 22 75 
<< m1 >>
rect 23 74 24 75 
<< m1 >>
rect 28 74 29 75 
<< m1 >>
rect 37 74 38 75 
<< m1 >>
rect 46 74 47 75 
<< m1 >>
rect 55 74 56 75 
<< m2 >>
rect 56 74 57 75 
<< m1 >>
rect 62 74 63 75 
<< m1 >>
rect 64 74 65 75 
<< m2 >>
rect 71 74 72 75 
<< m2 >>
rect 72 74 73 75 
<< m2 >>
rect 73 74 74 75 
<< m2 >>
rect 74 74 75 75 
<< m1 >>
rect 75 74 76 75 
<< m2 >>
rect 75 74 76 75 
<< m2c >>
rect 75 74 76 75 
<< m1 >>
rect 75 74 76 75 
<< m2 >>
rect 75 74 76 75 
<< m1 >>
rect 78 74 79 75 
<< m1 >>
rect 82 74 83 75 
<< m1 >>
rect 91 74 92 75 
<< m2 >>
rect 92 74 93 75 
<< m1 >>
rect 118 74 119 75 
<< m1 >>
rect 136 74 137 75 
<< m1 >>
rect 145 74 146 75 
<< m1 >>
rect 154 74 155 75 
<< m1 >>
rect 160 74 161 75 
<< m1 >>
rect 172 74 173 75 
<< m1 >>
rect 174 74 175 75 
<< m1 >>
rect 200 74 201 75 
<< m1 >>
rect 220 74 221 75 
<< m2 >>
rect 223 74 224 75 
<< m1 >>
rect 224 74 225 75 
<< m1 >>
rect 226 74 227 75 
<< m1 >>
rect 248 74 249 75 
<< m2 >>
rect 248 74 249 75 
<< m2c >>
rect 248 74 249 75 
<< m1 >>
rect 248 74 249 75 
<< m2 >>
rect 248 74 249 75 
<< m1 >>
rect 249 74 250 75 
<< m1 >>
rect 250 74 251 75 
<< m1 >>
rect 251 74 252 75 
<< m1 >>
rect 252 74 253 75 
<< m1 >>
rect 253 74 254 75 
<< m2 >>
rect 253 74 254 75 
<< m1 >>
rect 254 74 255 75 
<< m1 >>
rect 255 74 256 75 
<< m1 >>
rect 256 74 257 75 
<< m1 >>
rect 257 74 258 75 
<< m1 >>
rect 258 74 259 75 
<< m2 >>
rect 258 74 259 75 
<< m2c >>
rect 258 74 259 75 
<< m1 >>
rect 258 74 259 75 
<< m2 >>
rect 258 74 259 75 
<< m2 >>
rect 259 74 260 75 
<< m1 >>
rect 260 74 261 75 
<< m1 >>
rect 262 74 263 75 
<< m1 >>
rect 271 74 272 75 
<< m1 >>
rect 273 74 274 75 
<< m2 >>
rect 274 74 275 75 
<< m1 >>
rect 277 74 278 75 
<< m1 >>
rect 280 74 281 75 
<< m1 >>
rect 289 74 290 75 
<< m1 >>
rect 316 74 317 75 
<< m2 >>
rect 316 74 317 75 
<< m2c >>
rect 316 74 317 75 
<< m1 >>
rect 316 74 317 75 
<< m2 >>
rect 316 74 317 75 
<< m1 >>
rect 322 74 323 75 
<< m1 >>
rect 323 74 324 75 
<< m1 >>
rect 324 74 325 75 
<< m1 >>
rect 325 74 326 75 
<< m1 >>
rect 326 74 327 75 
<< m1 >>
rect 327 74 328 75 
<< m2 >>
rect 327 74 328 75 
<< m1 >>
rect 328 74 329 75 
<< m1 >>
rect 329 74 330 75 
<< m2 >>
rect 329 74 330 75 
<< m1 >>
rect 330 74 331 75 
<< m1 >>
rect 331 74 332 75 
<< m1 >>
rect 332 74 333 75 
<< m1 >>
rect 333 74 334 75 
<< m1 >>
rect 334 74 335 75 
<< m2 >>
rect 334 74 335 75 
<< m1 >>
rect 343 74 344 75 
<< m1 >>
rect 10 75 11 76 
<< m1 >>
rect 19 75 20 76 
<< m2 >>
rect 19 75 20 76 
<< m1 >>
rect 21 75 22 76 
<< m1 >>
rect 23 75 24 76 
<< m1 >>
rect 28 75 29 76 
<< m1 >>
rect 37 75 38 76 
<< m1 >>
rect 46 75 47 76 
<< m1 >>
rect 55 75 56 76 
<< m2 >>
rect 56 75 57 76 
<< m1 >>
rect 62 75 63 76 
<< m1 >>
rect 64 75 65 76 
<< m2 >>
rect 71 75 72 76 
<< m1 >>
rect 78 75 79 76 
<< m1 >>
rect 82 75 83 76 
<< m1 >>
rect 91 75 92 76 
<< m2 >>
rect 92 75 93 76 
<< m1 >>
rect 118 75 119 76 
<< m1 >>
rect 136 75 137 76 
<< m1 >>
rect 145 75 146 76 
<< m2 >>
rect 145 75 146 76 
<< m2c >>
rect 145 75 146 76 
<< m1 >>
rect 145 75 146 76 
<< m2 >>
rect 145 75 146 76 
<< m1 >>
rect 154 75 155 76 
<< m1 >>
rect 155 75 156 76 
<< m1 >>
rect 156 75 157 76 
<< m2 >>
rect 156 75 157 76 
<< m2c >>
rect 156 75 157 76 
<< m1 >>
rect 156 75 157 76 
<< m2 >>
rect 156 75 157 76 
<< m1 >>
rect 160 75 161 76 
<< m2 >>
rect 160 75 161 76 
<< m2c >>
rect 160 75 161 76 
<< m1 >>
rect 160 75 161 76 
<< m2 >>
rect 160 75 161 76 
<< m1 >>
rect 172 75 173 76 
<< m1 >>
rect 174 75 175 76 
<< m1 >>
rect 200 75 201 76 
<< m1 >>
rect 220 75 221 76 
<< m2 >>
rect 223 75 224 76 
<< m1 >>
rect 224 75 225 76 
<< m1 >>
rect 226 75 227 76 
<< m2 >>
rect 248 75 249 76 
<< m2 >>
rect 253 75 254 76 
<< m1 >>
rect 260 75 261 76 
<< m1 >>
rect 262 75 263 76 
<< m1 >>
rect 271 75 272 76 
<< m1 >>
rect 273 75 274 76 
<< m2 >>
rect 274 75 275 76 
<< m1 >>
rect 277 75 278 76 
<< m1 >>
rect 280 75 281 76 
<< m1 >>
rect 289 75 290 76 
<< m2 >>
rect 316 75 317 76 
<< m1 >>
rect 322 75 323 76 
<< m2 >>
rect 327 75 328 76 
<< m2 >>
rect 329 75 330 76 
<< m2 >>
rect 334 75 335 76 
<< m1 >>
rect 343 75 344 76 
<< m1 >>
rect 10 76 11 77 
<< m1 >>
rect 19 76 20 77 
<< m2 >>
rect 19 76 20 77 
<< m1 >>
rect 21 76 22 77 
<< m1 >>
rect 23 76 24 77 
<< m1 >>
rect 28 76 29 77 
<< m1 >>
rect 37 76 38 77 
<< m1 >>
rect 46 76 47 77 
<< m1 >>
rect 55 76 56 77 
<< m2 >>
rect 56 76 57 77 
<< m1 >>
rect 57 76 58 77 
<< m1 >>
rect 58 76 59 77 
<< m1 >>
rect 59 76 60 77 
<< m1 >>
rect 60 76 61 77 
<< m2 >>
rect 60 76 61 77 
<< m2c >>
rect 60 76 61 77 
<< m1 >>
rect 60 76 61 77 
<< m2 >>
rect 60 76 61 77 
<< m2 >>
rect 61 76 62 77 
<< m1 >>
rect 62 76 63 77 
<< m2 >>
rect 62 76 63 77 
<< m2 >>
rect 63 76 64 77 
<< m1 >>
rect 64 76 65 77 
<< m2 >>
rect 64 76 65 77 
<< m2 >>
rect 65 76 66 77 
<< m1 >>
rect 66 76 67 77 
<< m2 >>
rect 66 76 67 77 
<< m2c >>
rect 66 76 67 77 
<< m1 >>
rect 66 76 67 77 
<< m2 >>
rect 66 76 67 77 
<< m1 >>
rect 67 76 68 77 
<< m1 >>
rect 68 76 69 77 
<< m1 >>
rect 69 76 70 77 
<< m1 >>
rect 70 76 71 77 
<< m1 >>
rect 71 76 72 77 
<< m2 >>
rect 71 76 72 77 
<< m1 >>
rect 72 76 73 77 
<< m1 >>
rect 73 76 74 77 
<< m2 >>
rect 73 76 74 77 
<< m2c >>
rect 73 76 74 77 
<< m1 >>
rect 73 76 74 77 
<< m2 >>
rect 73 76 74 77 
<< m1 >>
rect 78 76 79 77 
<< m1 >>
rect 82 76 83 77 
<< m1 >>
rect 91 76 92 77 
<< m2 >>
rect 92 76 93 77 
<< m1 >>
rect 118 76 119 77 
<< m1 >>
rect 136 76 137 77 
<< m2 >>
rect 145 76 146 77 
<< m2 >>
rect 156 76 157 77 
<< m2 >>
rect 160 76 161 77 
<< m1 >>
rect 172 76 173 77 
<< m1 >>
rect 174 76 175 77 
<< m1 >>
rect 175 76 176 77 
<< m1 >>
rect 176 76 177 77 
<< m1 >>
rect 177 76 178 77 
<< m1 >>
rect 178 76 179 77 
<< m1 >>
rect 179 76 180 77 
<< m1 >>
rect 180 76 181 77 
<< m1 >>
rect 181 76 182 77 
<< m1 >>
rect 182 76 183 77 
<< m1 >>
rect 183 76 184 77 
<< m1 >>
rect 184 76 185 77 
<< m1 >>
rect 185 76 186 77 
<< m1 >>
rect 186 76 187 77 
<< m1 >>
rect 187 76 188 77 
<< m1 >>
rect 188 76 189 77 
<< m1 >>
rect 189 76 190 77 
<< m1 >>
rect 190 76 191 77 
<< m1 >>
rect 191 76 192 77 
<< m1 >>
rect 192 76 193 77 
<< m1 >>
rect 193 76 194 77 
<< m1 >>
rect 194 76 195 77 
<< m1 >>
rect 195 76 196 77 
<< m1 >>
rect 196 76 197 77 
<< m1 >>
rect 197 76 198 77 
<< m1 >>
rect 198 76 199 77 
<< m2 >>
rect 198 76 199 77 
<< m2c >>
rect 198 76 199 77 
<< m1 >>
rect 198 76 199 77 
<< m2 >>
rect 198 76 199 77 
<< m2 >>
rect 199 76 200 77 
<< m1 >>
rect 200 76 201 77 
<< m2 >>
rect 200 76 201 77 
<< m2 >>
rect 201 76 202 77 
<< m1 >>
rect 202 76 203 77 
<< m2 >>
rect 202 76 203 77 
<< m2c >>
rect 202 76 203 77 
<< m1 >>
rect 202 76 203 77 
<< m2 >>
rect 202 76 203 77 
<< m1 >>
rect 203 76 204 77 
<< m1 >>
rect 220 76 221 77 
<< m2 >>
rect 223 76 224 77 
<< m1 >>
rect 224 76 225 77 
<< m1 >>
rect 226 76 227 77 
<< m1 >>
rect 227 76 228 77 
<< m1 >>
rect 228 76 229 77 
<< m1 >>
rect 229 76 230 77 
<< m1 >>
rect 230 76 231 77 
<< m1 >>
rect 231 76 232 77 
<< m1 >>
rect 232 76 233 77 
<< m1 >>
rect 233 76 234 77 
<< m1 >>
rect 234 76 235 77 
<< m1 >>
rect 235 76 236 77 
<< m1 >>
rect 236 76 237 77 
<< m1 >>
rect 237 76 238 77 
<< m1 >>
rect 238 76 239 77 
<< m1 >>
rect 239 76 240 77 
<< m1 >>
rect 240 76 241 77 
<< m1 >>
rect 241 76 242 77 
<< m1 >>
rect 242 76 243 77 
<< m1 >>
rect 243 76 244 77 
<< m1 >>
rect 244 76 245 77 
<< m1 >>
rect 245 76 246 77 
<< m1 >>
rect 246 76 247 77 
<< m1 >>
rect 247 76 248 77 
<< m1 >>
rect 248 76 249 77 
<< m2 >>
rect 248 76 249 77 
<< m1 >>
rect 249 76 250 77 
<< m1 >>
rect 250 76 251 77 
<< m1 >>
rect 251 76 252 77 
<< m1 >>
rect 252 76 253 77 
<< m1 >>
rect 253 76 254 77 
<< m2 >>
rect 253 76 254 77 
<< m1 >>
rect 254 76 255 77 
<< m1 >>
rect 255 76 256 77 
<< m1 >>
rect 256 76 257 77 
<< m1 >>
rect 257 76 258 77 
<< m1 >>
rect 258 76 259 77 
<< m2 >>
rect 258 76 259 77 
<< m2c >>
rect 258 76 259 77 
<< m1 >>
rect 258 76 259 77 
<< m2 >>
rect 258 76 259 77 
<< m2 >>
rect 259 76 260 77 
<< m1 >>
rect 260 76 261 77 
<< m2 >>
rect 260 76 261 77 
<< m2 >>
rect 261 76 262 77 
<< m1 >>
rect 262 76 263 77 
<< m2 >>
rect 262 76 263 77 
<< m2 >>
rect 263 76 264 77 
<< m1 >>
rect 264 76 265 77 
<< m2 >>
rect 264 76 265 77 
<< m2c >>
rect 264 76 265 77 
<< m1 >>
rect 264 76 265 77 
<< m2 >>
rect 264 76 265 77 
<< m1 >>
rect 265 76 266 77 
<< m1 >>
rect 266 76 267 77 
<< m1 >>
rect 267 76 268 77 
<< m1 >>
rect 268 76 269 77 
<< m1 >>
rect 271 76 272 77 
<< m1 >>
rect 273 76 274 77 
<< m2 >>
rect 274 76 275 77 
<< m1 >>
rect 277 76 278 77 
<< m1 >>
rect 280 76 281 77 
<< m1 >>
rect 289 76 290 77 
<< m1 >>
rect 290 76 291 77 
<< m1 >>
rect 291 76 292 77 
<< m1 >>
rect 292 76 293 77 
<< m1 >>
rect 293 76 294 77 
<< m1 >>
rect 294 76 295 77 
<< m1 >>
rect 295 76 296 77 
<< m1 >>
rect 296 76 297 77 
<< m1 >>
rect 297 76 298 77 
<< m1 >>
rect 298 76 299 77 
<< m1 >>
rect 299 76 300 77 
<< m1 >>
rect 300 76 301 77 
<< m1 >>
rect 301 76 302 77 
<< m1 >>
rect 302 76 303 77 
<< m1 >>
rect 303 76 304 77 
<< m1 >>
rect 304 76 305 77 
<< m1 >>
rect 305 76 306 77 
<< m1 >>
rect 306 76 307 77 
<< m1 >>
rect 307 76 308 77 
<< m1 >>
rect 308 76 309 77 
<< m1 >>
rect 309 76 310 77 
<< m1 >>
rect 310 76 311 77 
<< m1 >>
rect 311 76 312 77 
<< m1 >>
rect 312 76 313 77 
<< m1 >>
rect 313 76 314 77 
<< m1 >>
rect 314 76 315 77 
<< m1 >>
rect 315 76 316 77 
<< m1 >>
rect 316 76 317 77 
<< m2 >>
rect 316 76 317 77 
<< m1 >>
rect 317 76 318 77 
<< m1 >>
rect 318 76 319 77 
<< m1 >>
rect 319 76 320 77 
<< m1 >>
rect 320 76 321 77 
<< m2 >>
rect 320 76 321 77 
<< m2c >>
rect 320 76 321 77 
<< m1 >>
rect 320 76 321 77 
<< m2 >>
rect 320 76 321 77 
<< m2 >>
rect 321 76 322 77 
<< m1 >>
rect 322 76 323 77 
<< m2 >>
rect 322 76 323 77 
<< m2 >>
rect 323 76 324 77 
<< m1 >>
rect 324 76 325 77 
<< m2 >>
rect 324 76 325 77 
<< m2c >>
rect 324 76 325 77 
<< m1 >>
rect 324 76 325 77 
<< m2 >>
rect 324 76 325 77 
<< m1 >>
rect 327 76 328 77 
<< m2 >>
rect 327 76 328 77 
<< m2c >>
rect 327 76 328 77 
<< m1 >>
rect 327 76 328 77 
<< m2 >>
rect 327 76 328 77 
<< m1 >>
rect 329 76 330 77 
<< m2 >>
rect 329 76 330 77 
<< m2c >>
rect 329 76 330 77 
<< m1 >>
rect 329 76 330 77 
<< m2 >>
rect 329 76 330 77 
<< m1 >>
rect 330 76 331 77 
<< m1 >>
rect 331 76 332 77 
<< m1 >>
rect 334 76 335 77 
<< m2 >>
rect 334 76 335 77 
<< m2c >>
rect 334 76 335 77 
<< m1 >>
rect 334 76 335 77 
<< m2 >>
rect 334 76 335 77 
<< m1 >>
rect 343 76 344 77 
<< m1 >>
rect 10 77 11 78 
<< m1 >>
rect 19 77 20 78 
<< m2 >>
rect 19 77 20 78 
<< m1 >>
rect 21 77 22 78 
<< m1 >>
rect 23 77 24 78 
<< m1 >>
rect 28 77 29 78 
<< m1 >>
rect 37 77 38 78 
<< m1 >>
rect 46 77 47 78 
<< m1 >>
rect 55 77 56 78 
<< m2 >>
rect 56 77 57 78 
<< m1 >>
rect 57 77 58 78 
<< m1 >>
rect 62 77 63 78 
<< m1 >>
rect 64 77 65 78 
<< m2 >>
rect 71 77 72 78 
<< m2 >>
rect 73 77 74 78 
<< m1 >>
rect 78 77 79 78 
<< m1 >>
rect 82 77 83 78 
<< m1 >>
rect 91 77 92 78 
<< m2 >>
rect 92 77 93 78 
<< m1 >>
rect 115 77 116 78 
<< m1 >>
rect 116 77 117 78 
<< m2 >>
rect 116 77 117 78 
<< m2c >>
rect 116 77 117 78 
<< m1 >>
rect 116 77 117 78 
<< m2 >>
rect 116 77 117 78 
<< m2 >>
rect 117 77 118 78 
<< m1 >>
rect 118 77 119 78 
<< m2 >>
rect 118 77 119 78 
<< m2 >>
rect 119 77 120 78 
<< m1 >>
rect 120 77 121 78 
<< m2 >>
rect 120 77 121 78 
<< m2c >>
rect 120 77 121 78 
<< m1 >>
rect 120 77 121 78 
<< m2 >>
rect 120 77 121 78 
<< m1 >>
rect 121 77 122 78 
<< m1 >>
rect 122 77 123 78 
<< m1 >>
rect 123 77 124 78 
<< m1 >>
rect 124 77 125 78 
<< m1 >>
rect 125 77 126 78 
<< m1 >>
rect 126 77 127 78 
<< m1 >>
rect 127 77 128 78 
<< m1 >>
rect 128 77 129 78 
<< m1 >>
rect 129 77 130 78 
<< m1 >>
rect 130 77 131 78 
<< m1 >>
rect 131 77 132 78 
<< m1 >>
rect 132 77 133 78 
<< m1 >>
rect 133 77 134 78 
<< m1 >>
rect 134 77 135 78 
<< m2 >>
rect 134 77 135 78 
<< m2c >>
rect 134 77 135 78 
<< m1 >>
rect 134 77 135 78 
<< m2 >>
rect 134 77 135 78 
<< m2 >>
rect 135 77 136 78 
<< m1 >>
rect 136 77 137 78 
<< m2 >>
rect 136 77 137 78 
<< m2 >>
rect 137 77 138 78 
<< m1 >>
rect 138 77 139 78 
<< m2 >>
rect 138 77 139 78 
<< m2c >>
rect 138 77 139 78 
<< m1 >>
rect 138 77 139 78 
<< m2 >>
rect 138 77 139 78 
<< m1 >>
rect 139 77 140 78 
<< m1 >>
rect 140 77 141 78 
<< m1 >>
rect 141 77 142 78 
<< m1 >>
rect 142 77 143 78 
<< m1 >>
rect 143 77 144 78 
<< m1 >>
rect 144 77 145 78 
<< m1 >>
rect 145 77 146 78 
<< m2 >>
rect 145 77 146 78 
<< m1 >>
rect 146 77 147 78 
<< m1 >>
rect 147 77 148 78 
<< m1 >>
rect 148 77 149 78 
<< m1 >>
rect 149 77 150 78 
<< m1 >>
rect 150 77 151 78 
<< m1 >>
rect 151 77 152 78 
<< m1 >>
rect 152 77 153 78 
<< m1 >>
rect 153 77 154 78 
<< m1 >>
rect 154 77 155 78 
<< m1 >>
rect 155 77 156 78 
<< m1 >>
rect 156 77 157 78 
<< m2 >>
rect 156 77 157 78 
<< m1 >>
rect 157 77 158 78 
<< m1 >>
rect 158 77 159 78 
<< m1 >>
rect 159 77 160 78 
<< m1 >>
rect 160 77 161 78 
<< m2 >>
rect 160 77 161 78 
<< m1 >>
rect 161 77 162 78 
<< m1 >>
rect 162 77 163 78 
<< m1 >>
rect 163 77 164 78 
<< m1 >>
rect 164 77 165 78 
<< m1 >>
rect 165 77 166 78 
<< m1 >>
rect 166 77 167 78 
<< m1 >>
rect 167 77 168 78 
<< m1 >>
rect 168 77 169 78 
<< m2 >>
rect 168 77 169 78 
<< m2c >>
rect 168 77 169 78 
<< m1 >>
rect 168 77 169 78 
<< m2 >>
rect 168 77 169 78 
<< m1 >>
rect 172 77 173 78 
<< m1 >>
rect 200 77 201 78 
<< m1 >>
rect 203 77 204 78 
<< m1 >>
rect 220 77 221 78 
<< m2 >>
rect 223 77 224 78 
<< m1 >>
rect 224 77 225 78 
<< m2 >>
rect 236 77 237 78 
<< m2 >>
rect 237 77 238 78 
<< m2 >>
rect 238 77 239 78 
<< m2 >>
rect 239 77 240 78 
<< m2 >>
rect 240 77 241 78 
<< m2 >>
rect 241 77 242 78 
<< m2 >>
rect 242 77 243 78 
<< m2 >>
rect 243 77 244 78 
<< m2 >>
rect 244 77 245 78 
<< m2 >>
rect 245 77 246 78 
<< m2 >>
rect 246 77 247 78 
<< m2 >>
rect 247 77 248 78 
<< m2 >>
rect 248 77 249 78 
<< m2 >>
rect 253 77 254 78 
<< m1 >>
rect 260 77 261 78 
<< m1 >>
rect 262 77 263 78 
<< m1 >>
rect 268 77 269 78 
<< m1 >>
rect 271 77 272 78 
<< m1 >>
rect 273 77 274 78 
<< m2 >>
rect 274 77 275 78 
<< m1 >>
rect 277 77 278 78 
<< m1 >>
rect 280 77 281 78 
<< m2 >>
rect 316 77 317 78 
<< m1 >>
rect 322 77 323 78 
<< m1 >>
rect 324 77 325 78 
<< m1 >>
rect 327 77 328 78 
<< m1 >>
rect 331 77 332 78 
<< m1 >>
rect 334 77 335 78 
<< m1 >>
rect 343 77 344 78 
<< m1 >>
rect 10 78 11 79 
<< m1 >>
rect 19 78 20 79 
<< m2 >>
rect 19 78 20 79 
<< m1 >>
rect 21 78 22 79 
<< m1 >>
rect 23 78 24 79 
<< m1 >>
rect 28 78 29 79 
<< m1 >>
rect 37 78 38 79 
<< m1 >>
rect 46 78 47 79 
<< m1 >>
rect 55 78 56 79 
<< m2 >>
rect 56 78 57 79 
<< m1 >>
rect 57 78 58 79 
<< m1 >>
rect 59 78 60 79 
<< m1 >>
rect 60 78 61 79 
<< m2 >>
rect 60 78 61 79 
<< m2c >>
rect 60 78 61 79 
<< m1 >>
rect 60 78 61 79 
<< m2 >>
rect 60 78 61 79 
<< m2 >>
rect 61 78 62 79 
<< m1 >>
rect 62 78 63 79 
<< m2 >>
rect 62 78 63 79 
<< m2 >>
rect 63 78 64 79 
<< m1 >>
rect 64 78 65 79 
<< m2 >>
rect 64 78 65 79 
<< m2 >>
rect 65 78 66 79 
<< m1 >>
rect 66 78 67 79 
<< m2 >>
rect 66 78 67 79 
<< m2c >>
rect 66 78 67 79 
<< m1 >>
rect 66 78 67 79 
<< m2 >>
rect 66 78 67 79 
<< m1 >>
rect 67 78 68 79 
<< m1 >>
rect 68 78 69 79 
<< m1 >>
rect 69 78 70 79 
<< m1 >>
rect 70 78 71 79 
<< m1 >>
rect 71 78 72 79 
<< m2 >>
rect 71 78 72 79 
<< m1 >>
rect 72 78 73 79 
<< m1 >>
rect 73 78 74 79 
<< m2 >>
rect 73 78 74 79 
<< m1 >>
rect 74 78 75 79 
<< m1 >>
rect 75 78 76 79 
<< m1 >>
rect 76 78 77 79 
<< m2 >>
rect 76 78 77 79 
<< m2c >>
rect 76 78 77 79 
<< m1 >>
rect 76 78 77 79 
<< m2 >>
rect 76 78 77 79 
<< m2 >>
rect 77 78 78 79 
<< m1 >>
rect 78 78 79 79 
<< m2 >>
rect 78 78 79 79 
<< m2 >>
rect 79 78 80 79 
<< m1 >>
rect 80 78 81 79 
<< m2 >>
rect 80 78 81 79 
<< m2c >>
rect 80 78 81 79 
<< m1 >>
rect 80 78 81 79 
<< m2 >>
rect 80 78 81 79 
<< m2 >>
rect 81 78 82 79 
<< m1 >>
rect 82 78 83 79 
<< m1 >>
rect 91 78 92 79 
<< m2 >>
rect 92 78 93 79 
<< m1 >>
rect 115 78 116 79 
<< m1 >>
rect 118 78 119 79 
<< m1 >>
rect 136 78 137 79 
<< m2 >>
rect 145 78 146 79 
<< m2 >>
rect 156 78 157 79 
<< m2 >>
rect 160 78 161 79 
<< m2 >>
rect 168 78 169 79 
<< m1 >>
rect 172 78 173 79 
<< m1 >>
rect 200 78 201 79 
<< m1 >>
rect 203 78 204 79 
<< m1 >>
rect 220 78 221 79 
<< m2 >>
rect 223 78 224 79 
<< m1 >>
rect 224 78 225 79 
<< m2 >>
rect 224 78 225 79 
<< m2 >>
rect 225 78 226 79 
<< m2 >>
rect 226 78 227 79 
<< m2 >>
rect 227 78 228 79 
<< m2 >>
rect 228 78 229 79 
<< m2 >>
rect 229 78 230 79 
<< m2 >>
rect 230 78 231 79 
<< m2 >>
rect 231 78 232 79 
<< m2 >>
rect 232 78 233 79 
<< m2 >>
rect 233 78 234 79 
<< m1 >>
rect 234 78 235 79 
<< m2 >>
rect 234 78 235 79 
<< m2c >>
rect 234 78 235 79 
<< m1 >>
rect 234 78 235 79 
<< m2 >>
rect 234 78 235 79 
<< m1 >>
rect 235 78 236 79 
<< m1 >>
rect 236 78 237 79 
<< m2 >>
rect 236 78 237 79 
<< m1 >>
rect 237 78 238 79 
<< m2 >>
rect 253 78 254 79 
<< m1 >>
rect 254 78 255 79 
<< m1 >>
rect 255 78 256 79 
<< m1 >>
rect 256 78 257 79 
<< m1 >>
rect 257 78 258 79 
<< m1 >>
rect 258 78 259 79 
<< m2 >>
rect 258 78 259 79 
<< m2c >>
rect 258 78 259 79 
<< m1 >>
rect 258 78 259 79 
<< m2 >>
rect 258 78 259 79 
<< m2 >>
rect 259 78 260 79 
<< m1 >>
rect 260 78 261 79 
<< m2 >>
rect 260 78 261 79 
<< m2 >>
rect 261 78 262 79 
<< m1 >>
rect 262 78 263 79 
<< m2 >>
rect 262 78 263 79 
<< m2 >>
rect 263 78 264 79 
<< m1 >>
rect 264 78 265 79 
<< m2 >>
rect 264 78 265 79 
<< m2c >>
rect 264 78 265 79 
<< m1 >>
rect 264 78 265 79 
<< m2 >>
rect 264 78 265 79 
<< m1 >>
rect 265 78 266 79 
<< m1 >>
rect 266 78 267 79 
<< m2 >>
rect 266 78 267 79 
<< m2c >>
rect 266 78 267 79 
<< m1 >>
rect 266 78 267 79 
<< m2 >>
rect 266 78 267 79 
<< m2 >>
rect 267 78 268 79 
<< m1 >>
rect 268 78 269 79 
<< m2 >>
rect 268 78 269 79 
<< m2 >>
rect 269 78 270 79 
<< m2 >>
rect 270 78 271 79 
<< m1 >>
rect 271 78 272 79 
<< m2 >>
rect 271 78 272 79 
<< m2 >>
rect 272 78 273 79 
<< m1 >>
rect 273 78 274 79 
<< m2 >>
rect 273 78 274 79 
<< m2 >>
rect 274 78 275 79 
<< m1 >>
rect 277 78 278 79 
<< m1 >>
rect 280 78 281 79 
<< m1 >>
rect 316 78 317 79 
<< m2 >>
rect 316 78 317 79 
<< m2c >>
rect 316 78 317 79 
<< m1 >>
rect 316 78 317 79 
<< m2 >>
rect 316 78 317 79 
<< m1 >>
rect 322 78 323 79 
<< m1 >>
rect 324 78 325 79 
<< m1 >>
rect 325 78 326 79 
<< m2 >>
rect 325 78 326 79 
<< m2c >>
rect 325 78 326 79 
<< m1 >>
rect 325 78 326 79 
<< m2 >>
rect 325 78 326 79 
<< m2 >>
rect 326 78 327 79 
<< m1 >>
rect 327 78 328 79 
<< m2 >>
rect 327 78 328 79 
<< m2 >>
rect 328 78 329 79 
<< m1 >>
rect 329 78 330 79 
<< m2 >>
rect 329 78 330 79 
<< m2c >>
rect 329 78 330 79 
<< m1 >>
rect 329 78 330 79 
<< m2 >>
rect 329 78 330 79 
<< m1 >>
rect 331 78 332 79 
<< m1 >>
rect 334 78 335 79 
<< m1 >>
rect 343 78 344 79 
<< m1 >>
rect 10 79 11 80 
<< m1 >>
rect 19 79 20 80 
<< m2 >>
rect 19 79 20 80 
<< m1 >>
rect 21 79 22 80 
<< m1 >>
rect 23 79 24 80 
<< m1 >>
rect 28 79 29 80 
<< m1 >>
rect 37 79 38 80 
<< m1 >>
rect 46 79 47 80 
<< m1 >>
rect 55 79 56 80 
<< m2 >>
rect 56 79 57 80 
<< m1 >>
rect 57 79 58 80 
<< m1 >>
rect 59 79 60 80 
<< m1 >>
rect 62 79 63 80 
<< m1 >>
rect 64 79 65 80 
<< m2 >>
rect 71 79 72 80 
<< m2 >>
rect 73 79 74 80 
<< m1 >>
rect 78 79 79 80 
<< m2 >>
rect 81 79 82 80 
<< m1 >>
rect 82 79 83 80 
<< m1 >>
rect 91 79 92 80 
<< m2 >>
rect 92 79 93 80 
<< m1 >>
rect 115 79 116 80 
<< m2 >>
rect 117 79 118 80 
<< m1 >>
rect 118 79 119 80 
<< m2 >>
rect 118 79 119 80 
<< m1 >>
rect 119 79 120 80 
<< m2 >>
rect 119 79 120 80 
<< m1 >>
rect 120 79 121 80 
<< m2 >>
rect 120 79 121 80 
<< m1 >>
rect 121 79 122 80 
<< m2 >>
rect 121 79 122 80 
<< m1 >>
rect 122 79 123 80 
<< m2 >>
rect 122 79 123 80 
<< m1 >>
rect 123 79 124 80 
<< m2 >>
rect 123 79 124 80 
<< m1 >>
rect 124 79 125 80 
<< m2 >>
rect 124 79 125 80 
<< m1 >>
rect 125 79 126 80 
<< m2 >>
rect 125 79 126 80 
<< m1 >>
rect 126 79 127 80 
<< m2 >>
rect 126 79 127 80 
<< m1 >>
rect 127 79 128 80 
<< m2 >>
rect 127 79 128 80 
<< m1 >>
rect 128 79 129 80 
<< m2 >>
rect 128 79 129 80 
<< m1 >>
rect 129 79 130 80 
<< m2 >>
rect 129 79 130 80 
<< m1 >>
rect 130 79 131 80 
<< m2 >>
rect 130 79 131 80 
<< m1 >>
rect 131 79 132 80 
<< m2 >>
rect 131 79 132 80 
<< m1 >>
rect 132 79 133 80 
<< m2 >>
rect 132 79 133 80 
<< m1 >>
rect 133 79 134 80 
<< m2 >>
rect 133 79 134 80 
<< m1 >>
rect 134 79 135 80 
<< m2 >>
rect 134 79 135 80 
<< m2 >>
rect 135 79 136 80 
<< m1 >>
rect 136 79 137 80 
<< m2 >>
rect 136 79 137 80 
<< m2 >>
rect 137 79 138 80 
<< m1 >>
rect 138 79 139 80 
<< m2 >>
rect 138 79 139 80 
<< m1 >>
rect 139 79 140 80 
<< m2 >>
rect 139 79 140 80 
<< m1 >>
rect 140 79 141 80 
<< m2 >>
rect 140 79 141 80 
<< m1 >>
rect 141 79 142 80 
<< m1 >>
rect 142 79 143 80 
<< m1 >>
rect 143 79 144 80 
<< m1 >>
rect 144 79 145 80 
<< m1 >>
rect 145 79 146 80 
<< m2 >>
rect 145 79 146 80 
<< m1 >>
rect 146 79 147 80 
<< m1 >>
rect 147 79 148 80 
<< m1 >>
rect 148 79 149 80 
<< m1 >>
rect 149 79 150 80 
<< m1 >>
rect 150 79 151 80 
<< m1 >>
rect 151 79 152 80 
<< m1 >>
rect 152 79 153 80 
<< m1 >>
rect 153 79 154 80 
<< m1 >>
rect 154 79 155 80 
<< m1 >>
rect 155 79 156 80 
<< m1 >>
rect 156 79 157 80 
<< m2 >>
rect 156 79 157 80 
<< m1 >>
rect 157 79 158 80 
<< m1 >>
rect 158 79 159 80 
<< m1 >>
rect 159 79 160 80 
<< m1 >>
rect 160 79 161 80 
<< m2 >>
rect 160 79 161 80 
<< m1 >>
rect 161 79 162 80 
<< m1 >>
rect 162 79 163 80 
<< m1 >>
rect 163 79 164 80 
<< m1 >>
rect 164 79 165 80 
<< m1 >>
rect 165 79 166 80 
<< m1 >>
rect 166 79 167 80 
<< m1 >>
rect 167 79 168 80 
<< m1 >>
rect 168 79 169 80 
<< m2 >>
rect 168 79 169 80 
<< m1 >>
rect 169 79 170 80 
<< m1 >>
rect 170 79 171 80 
<< m2 >>
rect 170 79 171 80 
<< m2c >>
rect 170 79 171 80 
<< m1 >>
rect 170 79 171 80 
<< m2 >>
rect 170 79 171 80 
<< m2 >>
rect 171 79 172 80 
<< m1 >>
rect 172 79 173 80 
<< m2 >>
rect 172 79 173 80 
<< m2 >>
rect 173 79 174 80 
<< m1 >>
rect 174 79 175 80 
<< m2 >>
rect 174 79 175 80 
<< m2c >>
rect 174 79 175 80 
<< m1 >>
rect 174 79 175 80 
<< m2 >>
rect 174 79 175 80 
<< m1 >>
rect 175 79 176 80 
<< m1 >>
rect 176 79 177 80 
<< m1 >>
rect 177 79 178 80 
<< m1 >>
rect 178 79 179 80 
<< m1 >>
rect 179 79 180 80 
<< m1 >>
rect 180 79 181 80 
<< m1 >>
rect 181 79 182 80 
<< m1 >>
rect 182 79 183 80 
<< m1 >>
rect 183 79 184 80 
<< m1 >>
rect 184 79 185 80 
<< m1 >>
rect 185 79 186 80 
<< m1 >>
rect 186 79 187 80 
<< m1 >>
rect 187 79 188 80 
<< m1 >>
rect 188 79 189 80 
<< m1 >>
rect 189 79 190 80 
<< m1 >>
rect 190 79 191 80 
<< m1 >>
rect 191 79 192 80 
<< m1 >>
rect 192 79 193 80 
<< m1 >>
rect 193 79 194 80 
<< m1 >>
rect 194 79 195 80 
<< m1 >>
rect 195 79 196 80 
<< m1 >>
rect 196 79 197 80 
<< m1 >>
rect 197 79 198 80 
<< m1 >>
rect 198 79 199 80 
<< m2 >>
rect 198 79 199 80 
<< m2c >>
rect 198 79 199 80 
<< m1 >>
rect 198 79 199 80 
<< m2 >>
rect 198 79 199 80 
<< m2 >>
rect 199 79 200 80 
<< m1 >>
rect 200 79 201 80 
<< m2 >>
rect 200 79 201 80 
<< m2 >>
rect 201 79 202 80 
<< m1 >>
rect 203 79 204 80 
<< m1 >>
rect 220 79 221 80 
<< m1 >>
rect 224 79 225 80 
<< m1 >>
rect 226 79 227 80 
<< m1 >>
rect 227 79 228 80 
<< m1 >>
rect 228 79 229 80 
<< m1 >>
rect 229 79 230 80 
<< m1 >>
rect 230 79 231 80 
<< m1 >>
rect 231 79 232 80 
<< m1 >>
rect 232 79 233 80 
<< m2 >>
rect 236 79 237 80 
<< m1 >>
rect 237 79 238 80 
<< m2 >>
rect 253 79 254 80 
<< m1 >>
rect 254 79 255 80 
<< m1 >>
rect 260 79 261 80 
<< m1 >>
rect 262 79 263 80 
<< m1 >>
rect 268 79 269 80 
<< m1 >>
rect 271 79 272 80 
<< m1 >>
rect 273 79 274 80 
<< m1 >>
rect 277 79 278 80 
<< m1 >>
rect 280 79 281 80 
<< m1 >>
rect 316 79 317 80 
<< m1 >>
rect 322 79 323 80 
<< m1 >>
rect 327 79 328 80 
<< m1 >>
rect 329 79 330 80 
<< m1 >>
rect 331 79 332 80 
<< m1 >>
rect 334 79 335 80 
<< m1 >>
rect 343 79 344 80 
<< m1 >>
rect 10 80 11 81 
<< m1 >>
rect 19 80 20 81 
<< m2 >>
rect 19 80 20 81 
<< m1 >>
rect 21 80 22 81 
<< m1 >>
rect 23 80 24 81 
<< m1 >>
rect 28 80 29 81 
<< m1 >>
rect 37 80 38 81 
<< m1 >>
rect 46 80 47 81 
<< m1 >>
rect 55 80 56 81 
<< m2 >>
rect 56 80 57 81 
<< m1 >>
rect 57 80 58 81 
<< m1 >>
rect 59 80 60 81 
<< m2 >>
rect 61 80 62 81 
<< m1 >>
rect 62 80 63 81 
<< m2 >>
rect 62 80 63 81 
<< m2 >>
rect 63 80 64 81 
<< m1 >>
rect 64 80 65 81 
<< m2 >>
rect 64 80 65 81 
<< m2c >>
rect 64 80 65 81 
<< m1 >>
rect 64 80 65 81 
<< m2 >>
rect 64 80 65 81 
<< m1 >>
rect 71 80 72 81 
<< m2 >>
rect 71 80 72 81 
<< m2c >>
rect 71 80 72 81 
<< m1 >>
rect 71 80 72 81 
<< m2 >>
rect 71 80 72 81 
<< m1 >>
rect 73 80 74 81 
<< m2 >>
rect 73 80 74 81 
<< m2c >>
rect 73 80 74 81 
<< m1 >>
rect 73 80 74 81 
<< m2 >>
rect 73 80 74 81 
<< m1 >>
rect 78 80 79 81 
<< m2 >>
rect 81 80 82 81 
<< m1 >>
rect 82 80 83 81 
<< m1 >>
rect 91 80 92 81 
<< m2 >>
rect 92 80 93 81 
<< m1 >>
rect 115 80 116 81 
<< m2 >>
rect 117 80 118 81 
<< m1 >>
rect 134 80 135 81 
<< m1 >>
rect 136 80 137 81 
<< m1 >>
rect 138 80 139 81 
<< m2 >>
rect 140 80 141 81 
<< m2 >>
rect 145 80 146 81 
<< m2 >>
rect 156 80 157 81 
<< m2 >>
rect 157 80 158 81 
<< m2 >>
rect 160 80 161 81 
<< m2 >>
rect 168 80 169 81 
<< m1 >>
rect 172 80 173 81 
<< m1 >>
rect 200 80 201 81 
<< m2 >>
rect 201 80 202 81 
<< m1 >>
rect 203 80 204 81 
<< m1 >>
rect 220 80 221 81 
<< m1 >>
rect 224 80 225 81 
<< m1 >>
rect 226 80 227 81 
<< m1 >>
rect 232 80 233 81 
<< m2 >>
rect 236 80 237 81 
<< m1 >>
rect 237 80 238 81 
<< m2 >>
rect 253 80 254 81 
<< m1 >>
rect 254 80 255 81 
<< m1 >>
rect 260 80 261 81 
<< m1 >>
rect 262 80 263 81 
<< m1 >>
rect 268 80 269 81 
<< m1 >>
rect 271 80 272 81 
<< m1 >>
rect 273 80 274 81 
<< m1 >>
rect 277 80 278 81 
<< m1 >>
rect 280 80 281 81 
<< m1 >>
rect 316 80 317 81 
<< m1 >>
rect 322 80 323 81 
<< m1 >>
rect 325 80 326 81 
<< m2 >>
rect 325 80 326 81 
<< m2c >>
rect 325 80 326 81 
<< m1 >>
rect 325 80 326 81 
<< m2 >>
rect 325 80 326 81 
<< m2 >>
rect 326 80 327 81 
<< m1 >>
rect 327 80 328 81 
<< m2 >>
rect 327 80 328 81 
<< m2 >>
rect 328 80 329 81 
<< m1 >>
rect 329 80 330 81 
<< m2 >>
rect 329 80 330 81 
<< m2 >>
rect 330 80 331 81 
<< m1 >>
rect 331 80 332 81 
<< m2 >>
rect 331 80 332 81 
<< m2c >>
rect 331 80 332 81 
<< m1 >>
rect 331 80 332 81 
<< m2 >>
rect 331 80 332 81 
<< m1 >>
rect 334 80 335 81 
<< m2 >>
rect 334 80 335 81 
<< m2c >>
rect 334 80 335 81 
<< m1 >>
rect 334 80 335 81 
<< m2 >>
rect 334 80 335 81 
<< m1 >>
rect 343 80 344 81 
<< m1 >>
rect 10 81 11 82 
<< m1 >>
rect 19 81 20 82 
<< m2 >>
rect 19 81 20 82 
<< m1 >>
rect 21 81 22 82 
<< m1 >>
rect 23 81 24 82 
<< m1 >>
rect 28 81 29 82 
<< m1 >>
rect 37 81 38 82 
<< m1 >>
rect 46 81 47 82 
<< m1 >>
rect 55 81 56 82 
<< m2 >>
rect 56 81 57 82 
<< m1 >>
rect 57 81 58 82 
<< m1 >>
rect 59 81 60 82 
<< m2 >>
rect 61 81 62 82 
<< m1 >>
rect 62 81 63 82 
<< m1 >>
rect 71 81 72 82 
<< m1 >>
rect 73 81 74 82 
<< m1 >>
rect 78 81 79 82 
<< m2 >>
rect 81 81 82 82 
<< m1 >>
rect 82 81 83 82 
<< m1 >>
rect 91 81 92 82 
<< m2 >>
rect 92 81 93 82 
<< m1 >>
rect 115 81 116 82 
<< m1 >>
rect 117 81 118 82 
<< m2 >>
rect 117 81 118 82 
<< m2c >>
rect 117 81 118 82 
<< m1 >>
rect 117 81 118 82 
<< m2 >>
rect 117 81 118 82 
<< m1 >>
rect 134 81 135 82 
<< m1 >>
rect 136 81 137 82 
<< m1 >>
rect 138 81 139 82 
<< m1 >>
rect 140 81 141 82 
<< m2 >>
rect 140 81 141 82 
<< m2c >>
rect 140 81 141 82 
<< m1 >>
rect 140 81 141 82 
<< m2 >>
rect 140 81 141 82 
<< m1 >>
rect 141 81 142 82 
<< m1 >>
rect 142 81 143 82 
<< m1 >>
rect 143 81 144 82 
<< m1 >>
rect 144 81 145 82 
<< m1 >>
rect 145 81 146 82 
<< m2 >>
rect 145 81 146 82 
<< m1 >>
rect 146 81 147 82 
<< m2 >>
rect 146 81 147 82 
<< m1 >>
rect 147 81 148 82 
<< m2 >>
rect 147 81 148 82 
<< m2 >>
rect 148 81 149 82 
<< m1 >>
rect 149 81 150 82 
<< m2 >>
rect 149 81 150 82 
<< m2c >>
rect 149 81 150 82 
<< m1 >>
rect 149 81 150 82 
<< m2 >>
rect 149 81 150 82 
<< m1 >>
rect 157 81 158 82 
<< m2 >>
rect 157 81 158 82 
<< m2c >>
rect 157 81 158 82 
<< m1 >>
rect 157 81 158 82 
<< m2 >>
rect 157 81 158 82 
<< m1 >>
rect 160 81 161 82 
<< m2 >>
rect 160 81 161 82 
<< m2c >>
rect 160 81 161 82 
<< m1 >>
rect 160 81 161 82 
<< m2 >>
rect 160 81 161 82 
<< m1 >>
rect 161 81 162 82 
<< m1 >>
rect 162 81 163 82 
<< m1 >>
rect 163 81 164 82 
<< m1 >>
rect 168 81 169 82 
<< m2 >>
rect 168 81 169 82 
<< m2c >>
rect 168 81 169 82 
<< m1 >>
rect 168 81 169 82 
<< m2 >>
rect 168 81 169 82 
<< m1 >>
rect 172 81 173 82 
<< m1 >>
rect 200 81 201 82 
<< m2 >>
rect 201 81 202 82 
<< m1 >>
rect 203 81 204 82 
<< m1 >>
rect 220 81 221 82 
<< m1 >>
rect 224 81 225 82 
<< m1 >>
rect 226 81 227 82 
<< m2 >>
rect 231 81 232 82 
<< m1 >>
rect 232 81 233 82 
<< m2 >>
rect 232 81 233 82 
<< m2 >>
rect 233 81 234 82 
<< m1 >>
rect 234 81 235 82 
<< m2 >>
rect 234 81 235 82 
<< m2c >>
rect 234 81 235 82 
<< m1 >>
rect 234 81 235 82 
<< m2 >>
rect 234 81 235 82 
<< m1 >>
rect 235 81 236 82 
<< m2 >>
rect 236 81 237 82 
<< m1 >>
rect 237 81 238 82 
<< m2 >>
rect 253 81 254 82 
<< m1 >>
rect 254 81 255 82 
<< m1 >>
rect 260 81 261 82 
<< m1 >>
rect 262 81 263 82 
<< m1 >>
rect 268 81 269 82 
<< m1 >>
rect 271 81 272 82 
<< m1 >>
rect 273 81 274 82 
<< m1 >>
rect 277 81 278 82 
<< m1 >>
rect 280 81 281 82 
<< m1 >>
rect 316 81 317 82 
<< m1 >>
rect 322 81 323 82 
<< m1 >>
rect 325 81 326 82 
<< m1 >>
rect 327 81 328 82 
<< m1 >>
rect 329 81 330 82 
<< m2 >>
rect 334 81 335 82 
<< m1 >>
rect 343 81 344 82 
<< m1 >>
rect 10 82 11 83 
<< m1 >>
rect 19 82 20 83 
<< m2 >>
rect 19 82 20 83 
<< m1 >>
rect 21 82 22 83 
<< m1 >>
rect 23 82 24 83 
<< m1 >>
rect 28 82 29 83 
<< m1 >>
rect 37 82 38 83 
<< m1 >>
rect 46 82 47 83 
<< m1 >>
rect 55 82 56 83 
<< m2 >>
rect 56 82 57 83 
<< m1 >>
rect 57 82 58 83 
<< m1 >>
rect 59 82 60 83 
<< m2 >>
rect 61 82 62 83 
<< m1 >>
rect 62 82 63 83 
<< m1 >>
rect 64 82 65 83 
<< m1 >>
rect 65 82 66 83 
<< m1 >>
rect 66 82 67 83 
<< m1 >>
rect 67 82 68 83 
<< m1 >>
rect 71 82 72 83 
<< m2 >>
rect 71 82 72 83 
<< m2c >>
rect 71 82 72 83 
<< m1 >>
rect 71 82 72 83 
<< m2 >>
rect 71 82 72 83 
<< m2 >>
rect 72 82 73 83 
<< m1 >>
rect 73 82 74 83 
<< m2 >>
rect 73 82 74 83 
<< m1 >>
rect 78 82 79 83 
<< m2 >>
rect 81 82 82 83 
<< m1 >>
rect 82 82 83 83 
<< m1 >>
rect 91 82 92 83 
<< m2 >>
rect 92 82 93 83 
<< m1 >>
rect 115 82 116 83 
<< m1 >>
rect 117 82 118 83 
<< m1 >>
rect 124 82 125 83 
<< m1 >>
rect 125 82 126 83 
<< m1 >>
rect 126 82 127 83 
<< m1 >>
rect 127 82 128 83 
<< m2 >>
rect 127 82 128 83 
<< m1 >>
rect 128 82 129 83 
<< m2 >>
rect 128 82 129 83 
<< m1 >>
rect 129 82 130 83 
<< m2 >>
rect 129 82 130 83 
<< m1 >>
rect 130 82 131 83 
<< m2 >>
rect 130 82 131 83 
<< m1 >>
rect 131 82 132 83 
<< m2 >>
rect 131 82 132 83 
<< m1 >>
rect 132 82 133 83 
<< m2 >>
rect 132 82 133 83 
<< m2 >>
rect 133 82 134 83 
<< m1 >>
rect 134 82 135 83 
<< m2 >>
rect 134 82 135 83 
<< m2 >>
rect 135 82 136 83 
<< m1 >>
rect 136 82 137 83 
<< m2 >>
rect 136 82 137 83 
<< m2 >>
rect 137 82 138 83 
<< m1 >>
rect 138 82 139 83 
<< m2 >>
rect 138 82 139 83 
<< m2c >>
rect 138 82 139 83 
<< m1 >>
rect 138 82 139 83 
<< m2 >>
rect 138 82 139 83 
<< m1 >>
rect 147 82 148 83 
<< m1 >>
rect 149 82 150 83 
<< m1 >>
rect 157 82 158 83 
<< m1 >>
rect 163 82 164 83 
<< m1 >>
rect 168 82 169 83 
<< m1 >>
rect 172 82 173 83 
<< m1 >>
rect 200 82 201 83 
<< m2 >>
rect 201 82 202 83 
<< m1 >>
rect 203 82 204 83 
<< m1 >>
rect 220 82 221 83 
<< m1 >>
rect 224 82 225 83 
<< m1 >>
rect 226 82 227 83 
<< m1 >>
rect 229 82 230 83 
<< m1 >>
rect 230 82 231 83 
<< m2 >>
rect 230 82 231 83 
<< m2c >>
rect 230 82 231 83 
<< m1 >>
rect 230 82 231 83 
<< m2 >>
rect 230 82 231 83 
<< m2 >>
rect 231 82 232 83 
<< m1 >>
rect 232 82 233 83 
<< m1 >>
rect 235 82 236 83 
<< m2 >>
rect 236 82 237 83 
<< m1 >>
rect 237 82 238 83 
<< m2 >>
rect 253 82 254 83 
<< m1 >>
rect 254 82 255 83 
<< m1 >>
rect 260 82 261 83 
<< m1 >>
rect 262 82 263 83 
<< m1 >>
rect 268 82 269 83 
<< m1 >>
rect 271 82 272 83 
<< m1 >>
rect 273 82 274 83 
<< m1 >>
rect 277 82 278 83 
<< m1 >>
rect 280 82 281 83 
<< m1 >>
rect 316 82 317 83 
<< m1 >>
rect 322 82 323 83 
<< m1 >>
rect 325 82 326 83 
<< m1 >>
rect 327 82 328 83 
<< m1 >>
rect 329 82 330 83 
<< m1 >>
rect 334 82 335 83 
<< m2 >>
rect 334 82 335 83 
<< m1 >>
rect 335 82 336 83 
<< m1 >>
rect 336 82 337 83 
<< m1 >>
rect 337 82 338 83 
<< m1 >>
rect 343 82 344 83 
<< m1 >>
rect 10 83 11 84 
<< m1 >>
rect 19 83 20 84 
<< m2 >>
rect 19 83 20 84 
<< m1 >>
rect 21 83 22 84 
<< m1 >>
rect 23 83 24 84 
<< m1 >>
rect 28 83 29 84 
<< m1 >>
rect 37 83 38 84 
<< m1 >>
rect 46 83 47 84 
<< m1 >>
rect 55 83 56 84 
<< m2 >>
rect 56 83 57 84 
<< m1 >>
rect 57 83 58 84 
<< m1 >>
rect 59 83 60 84 
<< m2 >>
rect 61 83 62 84 
<< m1 >>
rect 62 83 63 84 
<< m1 >>
rect 64 83 65 84 
<< m1 >>
rect 67 83 68 84 
<< m1 >>
rect 73 83 74 84 
<< m2 >>
rect 73 83 74 84 
<< m1 >>
rect 78 83 79 84 
<< m2 >>
rect 81 83 82 84 
<< m1 >>
rect 82 83 83 84 
<< m1 >>
rect 91 83 92 84 
<< m2 >>
rect 92 83 93 84 
<< m1 >>
rect 115 83 116 84 
<< m1 >>
rect 117 83 118 84 
<< m1 >>
rect 124 83 125 84 
<< m2 >>
rect 127 83 128 84 
<< m1 >>
rect 132 83 133 84 
<< m1 >>
rect 134 83 135 84 
<< m1 >>
rect 136 83 137 84 
<< m1 >>
rect 147 83 148 84 
<< m1 >>
rect 149 83 150 84 
<< m1 >>
rect 157 83 158 84 
<< m1 >>
rect 163 83 164 84 
<< m1 >>
rect 164 83 165 84 
<< m1 >>
rect 165 83 166 84 
<< m1 >>
rect 166 83 167 84 
<< m2 >>
rect 166 83 167 84 
<< m2c >>
rect 166 83 167 84 
<< m1 >>
rect 166 83 167 84 
<< m2 >>
rect 166 83 167 84 
<< m2 >>
rect 167 83 168 84 
<< m1 >>
rect 168 83 169 84 
<< m1 >>
rect 172 83 173 84 
<< m1 >>
rect 200 83 201 84 
<< m2 >>
rect 201 83 202 84 
<< m1 >>
rect 203 83 204 84 
<< m1 >>
rect 220 83 221 84 
<< m1 >>
rect 224 83 225 84 
<< m1 >>
rect 226 83 227 84 
<< m1 >>
rect 229 83 230 84 
<< m1 >>
rect 232 83 233 84 
<< m1 >>
rect 235 83 236 84 
<< m2 >>
rect 236 83 237 84 
<< m1 >>
rect 237 83 238 84 
<< m2 >>
rect 253 83 254 84 
<< m1 >>
rect 254 83 255 84 
<< m1 >>
rect 260 83 261 84 
<< m1 >>
rect 262 83 263 84 
<< m1 >>
rect 268 83 269 84 
<< m1 >>
rect 271 83 272 84 
<< m1 >>
rect 273 83 274 84 
<< m1 >>
rect 277 83 278 84 
<< m1 >>
rect 280 83 281 84 
<< m1 >>
rect 316 83 317 84 
<< m1 >>
rect 322 83 323 84 
<< m1 >>
rect 325 83 326 84 
<< m1 >>
rect 327 83 328 84 
<< m1 >>
rect 329 83 330 84 
<< m1 >>
rect 334 83 335 84 
<< m2 >>
rect 334 83 335 84 
<< m1 >>
rect 337 83 338 84 
<< m1 >>
rect 343 83 344 84 
<< m1 >>
rect 10 84 11 85 
<< pdiffusion >>
rect 12 84 13 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< m1 >>
rect 19 84 20 85 
<< m2 >>
rect 19 84 20 85 
<< m1 >>
rect 21 84 22 85 
<< m1 >>
rect 23 84 24 85 
<< m1 >>
rect 28 84 29 85 
<< m1 >>
rect 37 84 38 85 
<< m1 >>
rect 46 84 47 85 
<< pdiffusion >>
rect 48 84 49 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< m1 >>
rect 55 84 56 85 
<< m2 >>
rect 56 84 57 85 
<< m1 >>
rect 57 84 58 85 
<< m1 >>
rect 59 84 60 85 
<< m2 >>
rect 61 84 62 85 
<< m1 >>
rect 62 84 63 85 
<< m1 >>
rect 64 84 65 85 
<< pdiffusion >>
rect 66 84 67 85 
<< m1 >>
rect 67 84 68 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< m1 >>
rect 73 84 74 85 
<< m2 >>
rect 73 84 74 85 
<< m1 >>
rect 78 84 79 85 
<< m2 >>
rect 81 84 82 85 
<< m1 >>
rect 82 84 83 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 91 84 92 85 
<< m2 >>
rect 92 84 93 85 
<< pdiffusion >>
rect 102 84 103 85 
<< pdiffusion >>
rect 103 84 104 85 
<< pdiffusion >>
rect 104 84 105 85 
<< pdiffusion >>
rect 105 84 106 85 
<< pdiffusion >>
rect 106 84 107 85 
<< pdiffusion >>
rect 107 84 108 85 
<< m1 >>
rect 115 84 116 85 
<< m1 >>
rect 117 84 118 85 
<< pdiffusion >>
rect 120 84 121 85 
<< pdiffusion >>
rect 121 84 122 85 
<< pdiffusion >>
rect 122 84 123 85 
<< pdiffusion >>
rect 123 84 124 85 
<< m1 >>
rect 124 84 125 85 
<< pdiffusion >>
rect 124 84 125 85 
<< pdiffusion >>
rect 125 84 126 85 
<< m1 >>
rect 127 84 128 85 
<< m2 >>
rect 127 84 128 85 
<< m2c >>
rect 127 84 128 85 
<< m1 >>
rect 127 84 128 85 
<< m2 >>
rect 127 84 128 85 
<< m1 >>
rect 132 84 133 85 
<< m1 >>
rect 134 84 135 85 
<< m1 >>
rect 136 84 137 85 
<< pdiffusion >>
rect 138 84 139 85 
<< pdiffusion >>
rect 139 84 140 85 
<< pdiffusion >>
rect 140 84 141 85 
<< pdiffusion >>
rect 141 84 142 85 
<< pdiffusion >>
rect 142 84 143 85 
<< pdiffusion >>
rect 143 84 144 85 
<< m1 >>
rect 147 84 148 85 
<< m1 >>
rect 149 84 150 85 
<< pdiffusion >>
rect 156 84 157 85 
<< m1 >>
rect 157 84 158 85 
<< pdiffusion >>
rect 157 84 158 85 
<< pdiffusion >>
rect 158 84 159 85 
<< pdiffusion >>
rect 159 84 160 85 
<< pdiffusion >>
rect 160 84 161 85 
<< pdiffusion >>
rect 161 84 162 85 
<< m2 >>
rect 167 84 168 85 
<< m1 >>
rect 168 84 169 85 
<< m1 >>
rect 172 84 173 85 
<< pdiffusion >>
rect 174 84 175 85 
<< pdiffusion >>
rect 175 84 176 85 
<< pdiffusion >>
rect 176 84 177 85 
<< pdiffusion >>
rect 177 84 178 85 
<< pdiffusion >>
rect 178 84 179 85 
<< pdiffusion >>
rect 179 84 180 85 
<< pdiffusion >>
rect 192 84 193 85 
<< pdiffusion >>
rect 193 84 194 85 
<< pdiffusion >>
rect 194 84 195 85 
<< pdiffusion >>
rect 195 84 196 85 
<< pdiffusion >>
rect 196 84 197 85 
<< pdiffusion >>
rect 197 84 198 85 
<< m1 >>
rect 200 84 201 85 
<< m2 >>
rect 201 84 202 85 
<< m1 >>
rect 203 84 204 85 
<< pdiffusion >>
rect 210 84 211 85 
<< pdiffusion >>
rect 211 84 212 85 
<< pdiffusion >>
rect 212 84 213 85 
<< pdiffusion >>
rect 213 84 214 85 
<< pdiffusion >>
rect 214 84 215 85 
<< pdiffusion >>
rect 215 84 216 85 
<< m1 >>
rect 220 84 221 85 
<< m1 >>
rect 224 84 225 85 
<< m1 >>
rect 226 84 227 85 
<< pdiffusion >>
rect 228 84 229 85 
<< m1 >>
rect 229 84 230 85 
<< pdiffusion >>
rect 229 84 230 85 
<< pdiffusion >>
rect 230 84 231 85 
<< pdiffusion >>
rect 231 84 232 85 
<< m1 >>
rect 232 84 233 85 
<< pdiffusion >>
rect 232 84 233 85 
<< pdiffusion >>
rect 233 84 234 85 
<< m1 >>
rect 235 84 236 85 
<< m2 >>
rect 236 84 237 85 
<< m1 >>
rect 237 84 238 85 
<< pdiffusion >>
rect 246 84 247 85 
<< pdiffusion >>
rect 247 84 248 85 
<< pdiffusion >>
rect 248 84 249 85 
<< pdiffusion >>
rect 249 84 250 85 
<< pdiffusion >>
rect 250 84 251 85 
<< pdiffusion >>
rect 251 84 252 85 
<< m2 >>
rect 253 84 254 85 
<< m1 >>
rect 254 84 255 85 
<< m1 >>
rect 260 84 261 85 
<< m1 >>
rect 262 84 263 85 
<< pdiffusion >>
rect 264 84 265 85 
<< pdiffusion >>
rect 265 84 266 85 
<< pdiffusion >>
rect 266 84 267 85 
<< pdiffusion >>
rect 267 84 268 85 
<< m1 >>
rect 268 84 269 85 
<< pdiffusion >>
rect 268 84 269 85 
<< pdiffusion >>
rect 269 84 270 85 
<< m1 >>
rect 271 84 272 85 
<< m1 >>
rect 273 84 274 85 
<< m1 >>
rect 277 84 278 85 
<< m1 >>
rect 280 84 281 85 
<< pdiffusion >>
rect 282 84 283 85 
<< pdiffusion >>
rect 283 84 284 85 
<< pdiffusion >>
rect 284 84 285 85 
<< pdiffusion >>
rect 285 84 286 85 
<< pdiffusion >>
rect 286 84 287 85 
<< pdiffusion >>
rect 287 84 288 85 
<< pdiffusion >>
rect 300 84 301 85 
<< pdiffusion >>
rect 301 84 302 85 
<< pdiffusion >>
rect 302 84 303 85 
<< pdiffusion >>
rect 303 84 304 85 
<< pdiffusion >>
rect 304 84 305 85 
<< pdiffusion >>
rect 305 84 306 85 
<< m1 >>
rect 316 84 317 85 
<< pdiffusion >>
rect 318 84 319 85 
<< pdiffusion >>
rect 319 84 320 85 
<< pdiffusion >>
rect 320 84 321 85 
<< pdiffusion >>
rect 321 84 322 85 
<< m1 >>
rect 322 84 323 85 
<< pdiffusion >>
rect 322 84 323 85 
<< pdiffusion >>
rect 323 84 324 85 
<< m1 >>
rect 325 84 326 85 
<< m1 >>
rect 327 84 328 85 
<< m1 >>
rect 329 84 330 85 
<< m1 >>
rect 334 84 335 85 
<< m2 >>
rect 334 84 335 85 
<< pdiffusion >>
rect 336 84 337 85 
<< m1 >>
rect 337 84 338 85 
<< pdiffusion >>
rect 337 84 338 85 
<< pdiffusion >>
rect 338 84 339 85 
<< pdiffusion >>
rect 339 84 340 85 
<< pdiffusion >>
rect 340 84 341 85 
<< pdiffusion >>
rect 341 84 342 85 
<< m1 >>
rect 343 84 344 85 
<< m1 >>
rect 10 85 11 86 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< m1 >>
rect 19 85 20 86 
<< m2 >>
rect 19 85 20 86 
<< m1 >>
rect 21 85 22 86 
<< m1 >>
rect 23 85 24 86 
<< m1 >>
rect 28 85 29 86 
<< m1 >>
rect 37 85 38 86 
<< m1 >>
rect 46 85 47 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< m1 >>
rect 55 85 56 86 
<< m2 >>
rect 56 85 57 86 
<< m1 >>
rect 57 85 58 86 
<< m1 >>
rect 59 85 60 86 
<< m2 >>
rect 61 85 62 86 
<< m1 >>
rect 62 85 63 86 
<< m1 >>
rect 64 85 65 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< m1 >>
rect 73 85 74 86 
<< m2 >>
rect 73 85 74 86 
<< m1 >>
rect 78 85 79 86 
<< m2 >>
rect 81 85 82 86 
<< m1 >>
rect 82 85 83 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 91 85 92 86 
<< m2 >>
rect 92 85 93 86 
<< pdiffusion >>
rect 102 85 103 86 
<< pdiffusion >>
rect 103 85 104 86 
<< pdiffusion >>
rect 104 85 105 86 
<< pdiffusion >>
rect 105 85 106 86 
<< pdiffusion >>
rect 106 85 107 86 
<< pdiffusion >>
rect 107 85 108 86 
<< m1 >>
rect 115 85 116 86 
<< m1 >>
rect 117 85 118 86 
<< pdiffusion >>
rect 120 85 121 86 
<< pdiffusion >>
rect 121 85 122 86 
<< pdiffusion >>
rect 122 85 123 86 
<< pdiffusion >>
rect 123 85 124 86 
<< pdiffusion >>
rect 124 85 125 86 
<< pdiffusion >>
rect 125 85 126 86 
<< m1 >>
rect 127 85 128 86 
<< m1 >>
rect 132 85 133 86 
<< m1 >>
rect 134 85 135 86 
<< m1 >>
rect 136 85 137 86 
<< pdiffusion >>
rect 138 85 139 86 
<< pdiffusion >>
rect 139 85 140 86 
<< pdiffusion >>
rect 140 85 141 86 
<< pdiffusion >>
rect 141 85 142 86 
<< pdiffusion >>
rect 142 85 143 86 
<< pdiffusion >>
rect 143 85 144 86 
<< m1 >>
rect 147 85 148 86 
<< m1 >>
rect 149 85 150 86 
<< pdiffusion >>
rect 156 85 157 86 
<< pdiffusion >>
rect 157 85 158 86 
<< pdiffusion >>
rect 158 85 159 86 
<< pdiffusion >>
rect 159 85 160 86 
<< pdiffusion >>
rect 160 85 161 86 
<< pdiffusion >>
rect 161 85 162 86 
<< m2 >>
rect 167 85 168 86 
<< m1 >>
rect 168 85 169 86 
<< m1 >>
rect 172 85 173 86 
<< pdiffusion >>
rect 174 85 175 86 
<< pdiffusion >>
rect 175 85 176 86 
<< pdiffusion >>
rect 176 85 177 86 
<< pdiffusion >>
rect 177 85 178 86 
<< pdiffusion >>
rect 178 85 179 86 
<< pdiffusion >>
rect 179 85 180 86 
<< pdiffusion >>
rect 192 85 193 86 
<< pdiffusion >>
rect 193 85 194 86 
<< pdiffusion >>
rect 194 85 195 86 
<< pdiffusion >>
rect 195 85 196 86 
<< pdiffusion >>
rect 196 85 197 86 
<< pdiffusion >>
rect 197 85 198 86 
<< m1 >>
rect 200 85 201 86 
<< m2 >>
rect 201 85 202 86 
<< m1 >>
rect 203 85 204 86 
<< pdiffusion >>
rect 210 85 211 86 
<< pdiffusion >>
rect 211 85 212 86 
<< pdiffusion >>
rect 212 85 213 86 
<< pdiffusion >>
rect 213 85 214 86 
<< pdiffusion >>
rect 214 85 215 86 
<< pdiffusion >>
rect 215 85 216 86 
<< m1 >>
rect 220 85 221 86 
<< m1 >>
rect 224 85 225 86 
<< m1 >>
rect 226 85 227 86 
<< pdiffusion >>
rect 228 85 229 86 
<< pdiffusion >>
rect 229 85 230 86 
<< pdiffusion >>
rect 230 85 231 86 
<< pdiffusion >>
rect 231 85 232 86 
<< pdiffusion >>
rect 232 85 233 86 
<< pdiffusion >>
rect 233 85 234 86 
<< m1 >>
rect 235 85 236 86 
<< m2 >>
rect 236 85 237 86 
<< m1 >>
rect 237 85 238 86 
<< pdiffusion >>
rect 246 85 247 86 
<< pdiffusion >>
rect 247 85 248 86 
<< pdiffusion >>
rect 248 85 249 86 
<< pdiffusion >>
rect 249 85 250 86 
<< pdiffusion >>
rect 250 85 251 86 
<< pdiffusion >>
rect 251 85 252 86 
<< m2 >>
rect 253 85 254 86 
<< m1 >>
rect 254 85 255 86 
<< m1 >>
rect 260 85 261 86 
<< m1 >>
rect 262 85 263 86 
<< pdiffusion >>
rect 264 85 265 86 
<< pdiffusion >>
rect 265 85 266 86 
<< pdiffusion >>
rect 266 85 267 86 
<< pdiffusion >>
rect 267 85 268 86 
<< pdiffusion >>
rect 268 85 269 86 
<< pdiffusion >>
rect 269 85 270 86 
<< m1 >>
rect 271 85 272 86 
<< m1 >>
rect 273 85 274 86 
<< m1 >>
rect 277 85 278 86 
<< m1 >>
rect 280 85 281 86 
<< pdiffusion >>
rect 282 85 283 86 
<< pdiffusion >>
rect 283 85 284 86 
<< pdiffusion >>
rect 284 85 285 86 
<< pdiffusion >>
rect 285 85 286 86 
<< pdiffusion >>
rect 286 85 287 86 
<< pdiffusion >>
rect 287 85 288 86 
<< pdiffusion >>
rect 300 85 301 86 
<< pdiffusion >>
rect 301 85 302 86 
<< pdiffusion >>
rect 302 85 303 86 
<< pdiffusion >>
rect 303 85 304 86 
<< pdiffusion >>
rect 304 85 305 86 
<< pdiffusion >>
rect 305 85 306 86 
<< m1 >>
rect 316 85 317 86 
<< pdiffusion >>
rect 318 85 319 86 
<< pdiffusion >>
rect 319 85 320 86 
<< pdiffusion >>
rect 320 85 321 86 
<< pdiffusion >>
rect 321 85 322 86 
<< pdiffusion >>
rect 322 85 323 86 
<< pdiffusion >>
rect 323 85 324 86 
<< m1 >>
rect 325 85 326 86 
<< m1 >>
rect 327 85 328 86 
<< m1 >>
rect 329 85 330 86 
<< m1 >>
rect 334 85 335 86 
<< m2 >>
rect 334 85 335 86 
<< pdiffusion >>
rect 336 85 337 86 
<< pdiffusion >>
rect 337 85 338 86 
<< pdiffusion >>
rect 338 85 339 86 
<< pdiffusion >>
rect 339 85 340 86 
<< pdiffusion >>
rect 340 85 341 86 
<< pdiffusion >>
rect 341 85 342 86 
<< m1 >>
rect 343 85 344 86 
<< m1 >>
rect 10 86 11 87 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< m1 >>
rect 19 86 20 87 
<< m2 >>
rect 19 86 20 87 
<< m1 >>
rect 21 86 22 87 
<< m1 >>
rect 23 86 24 87 
<< m1 >>
rect 28 86 29 87 
<< m1 >>
rect 37 86 38 87 
<< m1 >>
rect 46 86 47 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< m1 >>
rect 55 86 56 87 
<< m2 >>
rect 56 86 57 87 
<< m1 >>
rect 57 86 58 87 
<< m1 >>
rect 59 86 60 87 
<< m2 >>
rect 61 86 62 87 
<< m1 >>
rect 62 86 63 87 
<< m1 >>
rect 64 86 65 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< m1 >>
rect 73 86 74 87 
<< m2 >>
rect 73 86 74 87 
<< m1 >>
rect 78 86 79 87 
<< m2 >>
rect 81 86 82 87 
<< m1 >>
rect 82 86 83 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 91 86 92 87 
<< m2 >>
rect 92 86 93 87 
<< pdiffusion >>
rect 102 86 103 87 
<< pdiffusion >>
rect 103 86 104 87 
<< pdiffusion >>
rect 104 86 105 87 
<< pdiffusion >>
rect 105 86 106 87 
<< pdiffusion >>
rect 106 86 107 87 
<< pdiffusion >>
rect 107 86 108 87 
<< m1 >>
rect 115 86 116 87 
<< m1 >>
rect 117 86 118 87 
<< pdiffusion >>
rect 120 86 121 87 
<< pdiffusion >>
rect 121 86 122 87 
<< pdiffusion >>
rect 122 86 123 87 
<< pdiffusion >>
rect 123 86 124 87 
<< pdiffusion >>
rect 124 86 125 87 
<< pdiffusion >>
rect 125 86 126 87 
<< m1 >>
rect 127 86 128 87 
<< m1 >>
rect 132 86 133 87 
<< m1 >>
rect 134 86 135 87 
<< m1 >>
rect 136 86 137 87 
<< pdiffusion >>
rect 138 86 139 87 
<< pdiffusion >>
rect 139 86 140 87 
<< pdiffusion >>
rect 140 86 141 87 
<< pdiffusion >>
rect 141 86 142 87 
<< pdiffusion >>
rect 142 86 143 87 
<< pdiffusion >>
rect 143 86 144 87 
<< m1 >>
rect 147 86 148 87 
<< m1 >>
rect 149 86 150 87 
<< pdiffusion >>
rect 156 86 157 87 
<< pdiffusion >>
rect 157 86 158 87 
<< pdiffusion >>
rect 158 86 159 87 
<< pdiffusion >>
rect 159 86 160 87 
<< pdiffusion >>
rect 160 86 161 87 
<< pdiffusion >>
rect 161 86 162 87 
<< m2 >>
rect 167 86 168 87 
<< m1 >>
rect 168 86 169 87 
<< m1 >>
rect 172 86 173 87 
<< pdiffusion >>
rect 174 86 175 87 
<< pdiffusion >>
rect 175 86 176 87 
<< pdiffusion >>
rect 176 86 177 87 
<< pdiffusion >>
rect 177 86 178 87 
<< pdiffusion >>
rect 178 86 179 87 
<< pdiffusion >>
rect 179 86 180 87 
<< pdiffusion >>
rect 192 86 193 87 
<< pdiffusion >>
rect 193 86 194 87 
<< pdiffusion >>
rect 194 86 195 87 
<< pdiffusion >>
rect 195 86 196 87 
<< pdiffusion >>
rect 196 86 197 87 
<< pdiffusion >>
rect 197 86 198 87 
<< m1 >>
rect 200 86 201 87 
<< m2 >>
rect 201 86 202 87 
<< m1 >>
rect 203 86 204 87 
<< pdiffusion >>
rect 210 86 211 87 
<< pdiffusion >>
rect 211 86 212 87 
<< pdiffusion >>
rect 212 86 213 87 
<< pdiffusion >>
rect 213 86 214 87 
<< pdiffusion >>
rect 214 86 215 87 
<< pdiffusion >>
rect 215 86 216 87 
<< m1 >>
rect 220 86 221 87 
<< m1 >>
rect 224 86 225 87 
<< m1 >>
rect 226 86 227 87 
<< pdiffusion >>
rect 228 86 229 87 
<< pdiffusion >>
rect 229 86 230 87 
<< pdiffusion >>
rect 230 86 231 87 
<< pdiffusion >>
rect 231 86 232 87 
<< pdiffusion >>
rect 232 86 233 87 
<< pdiffusion >>
rect 233 86 234 87 
<< m1 >>
rect 235 86 236 87 
<< m2 >>
rect 236 86 237 87 
<< m1 >>
rect 237 86 238 87 
<< pdiffusion >>
rect 246 86 247 87 
<< pdiffusion >>
rect 247 86 248 87 
<< pdiffusion >>
rect 248 86 249 87 
<< pdiffusion >>
rect 249 86 250 87 
<< pdiffusion >>
rect 250 86 251 87 
<< pdiffusion >>
rect 251 86 252 87 
<< m2 >>
rect 253 86 254 87 
<< m1 >>
rect 254 86 255 87 
<< m1 >>
rect 260 86 261 87 
<< m1 >>
rect 262 86 263 87 
<< pdiffusion >>
rect 264 86 265 87 
<< pdiffusion >>
rect 265 86 266 87 
<< pdiffusion >>
rect 266 86 267 87 
<< pdiffusion >>
rect 267 86 268 87 
<< pdiffusion >>
rect 268 86 269 87 
<< pdiffusion >>
rect 269 86 270 87 
<< m1 >>
rect 271 86 272 87 
<< m1 >>
rect 273 86 274 87 
<< m1 >>
rect 277 86 278 87 
<< m1 >>
rect 280 86 281 87 
<< pdiffusion >>
rect 282 86 283 87 
<< pdiffusion >>
rect 283 86 284 87 
<< pdiffusion >>
rect 284 86 285 87 
<< pdiffusion >>
rect 285 86 286 87 
<< pdiffusion >>
rect 286 86 287 87 
<< pdiffusion >>
rect 287 86 288 87 
<< pdiffusion >>
rect 300 86 301 87 
<< pdiffusion >>
rect 301 86 302 87 
<< pdiffusion >>
rect 302 86 303 87 
<< pdiffusion >>
rect 303 86 304 87 
<< pdiffusion >>
rect 304 86 305 87 
<< pdiffusion >>
rect 305 86 306 87 
<< m1 >>
rect 316 86 317 87 
<< pdiffusion >>
rect 318 86 319 87 
<< pdiffusion >>
rect 319 86 320 87 
<< pdiffusion >>
rect 320 86 321 87 
<< pdiffusion >>
rect 321 86 322 87 
<< pdiffusion >>
rect 322 86 323 87 
<< pdiffusion >>
rect 323 86 324 87 
<< m1 >>
rect 325 86 326 87 
<< m1 >>
rect 327 86 328 87 
<< m1 >>
rect 329 86 330 87 
<< m1 >>
rect 334 86 335 87 
<< m2 >>
rect 334 86 335 87 
<< pdiffusion >>
rect 336 86 337 87 
<< pdiffusion >>
rect 337 86 338 87 
<< pdiffusion >>
rect 338 86 339 87 
<< pdiffusion >>
rect 339 86 340 87 
<< pdiffusion >>
rect 340 86 341 87 
<< pdiffusion >>
rect 341 86 342 87 
<< m1 >>
rect 343 86 344 87 
<< m1 >>
rect 10 87 11 88 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< m1 >>
rect 19 87 20 88 
<< m2 >>
rect 19 87 20 88 
<< m1 >>
rect 21 87 22 88 
<< m1 >>
rect 23 87 24 88 
<< m1 >>
rect 28 87 29 88 
<< m1 >>
rect 37 87 38 88 
<< m1 >>
rect 46 87 47 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< m1 >>
rect 55 87 56 88 
<< m2 >>
rect 56 87 57 88 
<< m1 >>
rect 57 87 58 88 
<< m1 >>
rect 59 87 60 88 
<< m2 >>
rect 61 87 62 88 
<< m1 >>
rect 62 87 63 88 
<< m1 >>
rect 64 87 65 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< m1 >>
rect 73 87 74 88 
<< m2 >>
rect 73 87 74 88 
<< m1 >>
rect 78 87 79 88 
<< m2 >>
rect 81 87 82 88 
<< m1 >>
rect 82 87 83 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 91 87 92 88 
<< m2 >>
rect 92 87 93 88 
<< pdiffusion >>
rect 102 87 103 88 
<< pdiffusion >>
rect 103 87 104 88 
<< pdiffusion >>
rect 104 87 105 88 
<< pdiffusion >>
rect 105 87 106 88 
<< pdiffusion >>
rect 106 87 107 88 
<< pdiffusion >>
rect 107 87 108 88 
<< m1 >>
rect 115 87 116 88 
<< m1 >>
rect 117 87 118 88 
<< pdiffusion >>
rect 120 87 121 88 
<< pdiffusion >>
rect 121 87 122 88 
<< pdiffusion >>
rect 122 87 123 88 
<< pdiffusion >>
rect 123 87 124 88 
<< pdiffusion >>
rect 124 87 125 88 
<< pdiffusion >>
rect 125 87 126 88 
<< m1 >>
rect 127 87 128 88 
<< m1 >>
rect 132 87 133 88 
<< m1 >>
rect 134 87 135 88 
<< m1 >>
rect 136 87 137 88 
<< pdiffusion >>
rect 138 87 139 88 
<< pdiffusion >>
rect 139 87 140 88 
<< pdiffusion >>
rect 140 87 141 88 
<< pdiffusion >>
rect 141 87 142 88 
<< pdiffusion >>
rect 142 87 143 88 
<< pdiffusion >>
rect 143 87 144 88 
<< m1 >>
rect 147 87 148 88 
<< m1 >>
rect 149 87 150 88 
<< pdiffusion >>
rect 156 87 157 88 
<< pdiffusion >>
rect 157 87 158 88 
<< pdiffusion >>
rect 158 87 159 88 
<< pdiffusion >>
rect 159 87 160 88 
<< pdiffusion >>
rect 160 87 161 88 
<< pdiffusion >>
rect 161 87 162 88 
<< m2 >>
rect 167 87 168 88 
<< m1 >>
rect 168 87 169 88 
<< m1 >>
rect 172 87 173 88 
<< pdiffusion >>
rect 174 87 175 88 
<< pdiffusion >>
rect 175 87 176 88 
<< pdiffusion >>
rect 176 87 177 88 
<< pdiffusion >>
rect 177 87 178 88 
<< pdiffusion >>
rect 178 87 179 88 
<< pdiffusion >>
rect 179 87 180 88 
<< pdiffusion >>
rect 192 87 193 88 
<< pdiffusion >>
rect 193 87 194 88 
<< pdiffusion >>
rect 194 87 195 88 
<< pdiffusion >>
rect 195 87 196 88 
<< pdiffusion >>
rect 196 87 197 88 
<< pdiffusion >>
rect 197 87 198 88 
<< m1 >>
rect 200 87 201 88 
<< m2 >>
rect 201 87 202 88 
<< m1 >>
rect 203 87 204 88 
<< pdiffusion >>
rect 210 87 211 88 
<< pdiffusion >>
rect 211 87 212 88 
<< pdiffusion >>
rect 212 87 213 88 
<< pdiffusion >>
rect 213 87 214 88 
<< pdiffusion >>
rect 214 87 215 88 
<< pdiffusion >>
rect 215 87 216 88 
<< m1 >>
rect 220 87 221 88 
<< m1 >>
rect 224 87 225 88 
<< m1 >>
rect 226 87 227 88 
<< pdiffusion >>
rect 228 87 229 88 
<< pdiffusion >>
rect 229 87 230 88 
<< pdiffusion >>
rect 230 87 231 88 
<< pdiffusion >>
rect 231 87 232 88 
<< pdiffusion >>
rect 232 87 233 88 
<< pdiffusion >>
rect 233 87 234 88 
<< m1 >>
rect 235 87 236 88 
<< m2 >>
rect 236 87 237 88 
<< m1 >>
rect 237 87 238 88 
<< pdiffusion >>
rect 246 87 247 88 
<< pdiffusion >>
rect 247 87 248 88 
<< pdiffusion >>
rect 248 87 249 88 
<< pdiffusion >>
rect 249 87 250 88 
<< pdiffusion >>
rect 250 87 251 88 
<< pdiffusion >>
rect 251 87 252 88 
<< m2 >>
rect 253 87 254 88 
<< m1 >>
rect 254 87 255 88 
<< m1 >>
rect 260 87 261 88 
<< m1 >>
rect 262 87 263 88 
<< pdiffusion >>
rect 264 87 265 88 
<< pdiffusion >>
rect 265 87 266 88 
<< pdiffusion >>
rect 266 87 267 88 
<< pdiffusion >>
rect 267 87 268 88 
<< pdiffusion >>
rect 268 87 269 88 
<< pdiffusion >>
rect 269 87 270 88 
<< m1 >>
rect 271 87 272 88 
<< m1 >>
rect 273 87 274 88 
<< m1 >>
rect 277 87 278 88 
<< m1 >>
rect 280 87 281 88 
<< pdiffusion >>
rect 282 87 283 88 
<< pdiffusion >>
rect 283 87 284 88 
<< pdiffusion >>
rect 284 87 285 88 
<< pdiffusion >>
rect 285 87 286 88 
<< pdiffusion >>
rect 286 87 287 88 
<< pdiffusion >>
rect 287 87 288 88 
<< pdiffusion >>
rect 300 87 301 88 
<< pdiffusion >>
rect 301 87 302 88 
<< pdiffusion >>
rect 302 87 303 88 
<< pdiffusion >>
rect 303 87 304 88 
<< pdiffusion >>
rect 304 87 305 88 
<< pdiffusion >>
rect 305 87 306 88 
<< m1 >>
rect 316 87 317 88 
<< pdiffusion >>
rect 318 87 319 88 
<< pdiffusion >>
rect 319 87 320 88 
<< pdiffusion >>
rect 320 87 321 88 
<< pdiffusion >>
rect 321 87 322 88 
<< pdiffusion >>
rect 322 87 323 88 
<< pdiffusion >>
rect 323 87 324 88 
<< m1 >>
rect 325 87 326 88 
<< m1 >>
rect 327 87 328 88 
<< m1 >>
rect 329 87 330 88 
<< m1 >>
rect 334 87 335 88 
<< m2 >>
rect 334 87 335 88 
<< pdiffusion >>
rect 336 87 337 88 
<< pdiffusion >>
rect 337 87 338 88 
<< pdiffusion >>
rect 338 87 339 88 
<< pdiffusion >>
rect 339 87 340 88 
<< pdiffusion >>
rect 340 87 341 88 
<< pdiffusion >>
rect 341 87 342 88 
<< m1 >>
rect 343 87 344 88 
<< m1 >>
rect 10 88 11 89 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< m1 >>
rect 19 88 20 89 
<< m2 >>
rect 19 88 20 89 
<< m1 >>
rect 21 88 22 89 
<< m1 >>
rect 23 88 24 89 
<< m1 >>
rect 28 88 29 89 
<< m1 >>
rect 37 88 38 89 
<< m1 >>
rect 46 88 47 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< m1 >>
rect 55 88 56 89 
<< m2 >>
rect 56 88 57 89 
<< m1 >>
rect 57 88 58 89 
<< m1 >>
rect 59 88 60 89 
<< m2 >>
rect 61 88 62 89 
<< m1 >>
rect 62 88 63 89 
<< m1 >>
rect 64 88 65 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< m1 >>
rect 73 88 74 89 
<< m2 >>
rect 73 88 74 89 
<< m1 >>
rect 78 88 79 89 
<< m2 >>
rect 81 88 82 89 
<< m1 >>
rect 82 88 83 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 91 88 92 89 
<< m2 >>
rect 92 88 93 89 
<< pdiffusion >>
rect 102 88 103 89 
<< pdiffusion >>
rect 103 88 104 89 
<< pdiffusion >>
rect 104 88 105 89 
<< pdiffusion >>
rect 105 88 106 89 
<< pdiffusion >>
rect 106 88 107 89 
<< pdiffusion >>
rect 107 88 108 89 
<< m1 >>
rect 115 88 116 89 
<< m1 >>
rect 117 88 118 89 
<< pdiffusion >>
rect 120 88 121 89 
<< pdiffusion >>
rect 121 88 122 89 
<< pdiffusion >>
rect 122 88 123 89 
<< pdiffusion >>
rect 123 88 124 89 
<< pdiffusion >>
rect 124 88 125 89 
<< pdiffusion >>
rect 125 88 126 89 
<< m1 >>
rect 127 88 128 89 
<< m1 >>
rect 132 88 133 89 
<< m1 >>
rect 134 88 135 89 
<< m1 >>
rect 136 88 137 89 
<< pdiffusion >>
rect 138 88 139 89 
<< pdiffusion >>
rect 139 88 140 89 
<< pdiffusion >>
rect 140 88 141 89 
<< pdiffusion >>
rect 141 88 142 89 
<< pdiffusion >>
rect 142 88 143 89 
<< pdiffusion >>
rect 143 88 144 89 
<< m1 >>
rect 147 88 148 89 
<< m1 >>
rect 149 88 150 89 
<< pdiffusion >>
rect 156 88 157 89 
<< pdiffusion >>
rect 157 88 158 89 
<< pdiffusion >>
rect 158 88 159 89 
<< pdiffusion >>
rect 159 88 160 89 
<< pdiffusion >>
rect 160 88 161 89 
<< pdiffusion >>
rect 161 88 162 89 
<< m2 >>
rect 167 88 168 89 
<< m1 >>
rect 168 88 169 89 
<< m1 >>
rect 172 88 173 89 
<< pdiffusion >>
rect 174 88 175 89 
<< pdiffusion >>
rect 175 88 176 89 
<< pdiffusion >>
rect 176 88 177 89 
<< pdiffusion >>
rect 177 88 178 89 
<< pdiffusion >>
rect 178 88 179 89 
<< pdiffusion >>
rect 179 88 180 89 
<< pdiffusion >>
rect 192 88 193 89 
<< pdiffusion >>
rect 193 88 194 89 
<< pdiffusion >>
rect 194 88 195 89 
<< pdiffusion >>
rect 195 88 196 89 
<< pdiffusion >>
rect 196 88 197 89 
<< pdiffusion >>
rect 197 88 198 89 
<< m1 >>
rect 200 88 201 89 
<< m2 >>
rect 201 88 202 89 
<< m1 >>
rect 203 88 204 89 
<< pdiffusion >>
rect 210 88 211 89 
<< pdiffusion >>
rect 211 88 212 89 
<< pdiffusion >>
rect 212 88 213 89 
<< pdiffusion >>
rect 213 88 214 89 
<< pdiffusion >>
rect 214 88 215 89 
<< pdiffusion >>
rect 215 88 216 89 
<< m1 >>
rect 220 88 221 89 
<< m1 >>
rect 224 88 225 89 
<< m1 >>
rect 226 88 227 89 
<< pdiffusion >>
rect 228 88 229 89 
<< pdiffusion >>
rect 229 88 230 89 
<< pdiffusion >>
rect 230 88 231 89 
<< pdiffusion >>
rect 231 88 232 89 
<< pdiffusion >>
rect 232 88 233 89 
<< pdiffusion >>
rect 233 88 234 89 
<< m1 >>
rect 235 88 236 89 
<< m2 >>
rect 236 88 237 89 
<< m1 >>
rect 237 88 238 89 
<< pdiffusion >>
rect 246 88 247 89 
<< pdiffusion >>
rect 247 88 248 89 
<< pdiffusion >>
rect 248 88 249 89 
<< pdiffusion >>
rect 249 88 250 89 
<< pdiffusion >>
rect 250 88 251 89 
<< pdiffusion >>
rect 251 88 252 89 
<< m2 >>
rect 253 88 254 89 
<< m1 >>
rect 254 88 255 89 
<< m1 >>
rect 260 88 261 89 
<< m1 >>
rect 262 88 263 89 
<< pdiffusion >>
rect 264 88 265 89 
<< pdiffusion >>
rect 265 88 266 89 
<< pdiffusion >>
rect 266 88 267 89 
<< pdiffusion >>
rect 267 88 268 89 
<< pdiffusion >>
rect 268 88 269 89 
<< pdiffusion >>
rect 269 88 270 89 
<< m1 >>
rect 271 88 272 89 
<< m1 >>
rect 273 88 274 89 
<< m1 >>
rect 277 88 278 89 
<< m1 >>
rect 280 88 281 89 
<< pdiffusion >>
rect 282 88 283 89 
<< pdiffusion >>
rect 283 88 284 89 
<< pdiffusion >>
rect 284 88 285 89 
<< pdiffusion >>
rect 285 88 286 89 
<< pdiffusion >>
rect 286 88 287 89 
<< pdiffusion >>
rect 287 88 288 89 
<< pdiffusion >>
rect 300 88 301 89 
<< pdiffusion >>
rect 301 88 302 89 
<< pdiffusion >>
rect 302 88 303 89 
<< pdiffusion >>
rect 303 88 304 89 
<< pdiffusion >>
rect 304 88 305 89 
<< pdiffusion >>
rect 305 88 306 89 
<< m1 >>
rect 316 88 317 89 
<< pdiffusion >>
rect 318 88 319 89 
<< pdiffusion >>
rect 319 88 320 89 
<< pdiffusion >>
rect 320 88 321 89 
<< pdiffusion >>
rect 321 88 322 89 
<< pdiffusion >>
rect 322 88 323 89 
<< pdiffusion >>
rect 323 88 324 89 
<< m1 >>
rect 325 88 326 89 
<< m1 >>
rect 327 88 328 89 
<< m1 >>
rect 329 88 330 89 
<< m1 >>
rect 334 88 335 89 
<< m2 >>
rect 334 88 335 89 
<< pdiffusion >>
rect 336 88 337 89 
<< pdiffusion >>
rect 337 88 338 89 
<< pdiffusion >>
rect 338 88 339 89 
<< pdiffusion >>
rect 339 88 340 89 
<< pdiffusion >>
rect 340 88 341 89 
<< pdiffusion >>
rect 341 88 342 89 
<< m1 >>
rect 343 88 344 89 
<< m1 >>
rect 10 89 11 90 
<< pdiffusion >>
rect 12 89 13 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< m1 >>
rect 19 89 20 90 
<< m2 >>
rect 19 89 20 90 
<< m1 >>
rect 21 89 22 90 
<< m1 >>
rect 23 89 24 90 
<< m1 >>
rect 28 89 29 90 
<< m1 >>
rect 37 89 38 90 
<< m1 >>
rect 46 89 47 90 
<< pdiffusion >>
rect 48 89 49 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< m1 >>
rect 55 89 56 90 
<< m2 >>
rect 56 89 57 90 
<< m1 >>
rect 57 89 58 90 
<< m1 >>
rect 59 89 60 90 
<< m2 >>
rect 61 89 62 90 
<< m1 >>
rect 62 89 63 90 
<< m1 >>
rect 64 89 65 90 
<< pdiffusion >>
rect 66 89 67 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< m1 >>
rect 73 89 74 90 
<< m2 >>
rect 73 89 74 90 
<< m1 >>
rect 78 89 79 90 
<< m2 >>
rect 81 89 82 90 
<< m1 >>
rect 82 89 83 90 
<< pdiffusion >>
rect 84 89 85 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 91 89 92 90 
<< m2 >>
rect 92 89 93 90 
<< pdiffusion >>
rect 102 89 103 90 
<< pdiffusion >>
rect 103 89 104 90 
<< pdiffusion >>
rect 104 89 105 90 
<< pdiffusion >>
rect 105 89 106 90 
<< pdiffusion >>
rect 106 89 107 90 
<< pdiffusion >>
rect 107 89 108 90 
<< m1 >>
rect 115 89 116 90 
<< m1 >>
rect 117 89 118 90 
<< pdiffusion >>
rect 120 89 121 90 
<< pdiffusion >>
rect 121 89 122 90 
<< pdiffusion >>
rect 122 89 123 90 
<< pdiffusion >>
rect 123 89 124 90 
<< m1 >>
rect 124 89 125 90 
<< pdiffusion >>
rect 124 89 125 90 
<< pdiffusion >>
rect 125 89 126 90 
<< m1 >>
rect 127 89 128 90 
<< m1 >>
rect 132 89 133 90 
<< m1 >>
rect 134 89 135 90 
<< m1 >>
rect 136 89 137 90 
<< pdiffusion >>
rect 138 89 139 90 
<< pdiffusion >>
rect 139 89 140 90 
<< pdiffusion >>
rect 140 89 141 90 
<< pdiffusion >>
rect 141 89 142 90 
<< pdiffusion >>
rect 142 89 143 90 
<< pdiffusion >>
rect 143 89 144 90 
<< m1 >>
rect 147 89 148 90 
<< m1 >>
rect 149 89 150 90 
<< pdiffusion >>
rect 156 89 157 90 
<< m1 >>
rect 157 89 158 90 
<< pdiffusion >>
rect 157 89 158 90 
<< pdiffusion >>
rect 158 89 159 90 
<< pdiffusion >>
rect 159 89 160 90 
<< pdiffusion >>
rect 160 89 161 90 
<< pdiffusion >>
rect 161 89 162 90 
<< m2 >>
rect 167 89 168 90 
<< m1 >>
rect 168 89 169 90 
<< m1 >>
rect 172 89 173 90 
<< pdiffusion >>
rect 174 89 175 90 
<< pdiffusion >>
rect 175 89 176 90 
<< pdiffusion >>
rect 176 89 177 90 
<< pdiffusion >>
rect 177 89 178 90 
<< pdiffusion >>
rect 178 89 179 90 
<< pdiffusion >>
rect 179 89 180 90 
<< pdiffusion >>
rect 192 89 193 90 
<< pdiffusion >>
rect 193 89 194 90 
<< pdiffusion >>
rect 194 89 195 90 
<< pdiffusion >>
rect 195 89 196 90 
<< pdiffusion >>
rect 196 89 197 90 
<< pdiffusion >>
rect 197 89 198 90 
<< m1 >>
rect 200 89 201 90 
<< m2 >>
rect 201 89 202 90 
<< m1 >>
rect 203 89 204 90 
<< pdiffusion >>
rect 210 89 211 90 
<< pdiffusion >>
rect 211 89 212 90 
<< pdiffusion >>
rect 212 89 213 90 
<< pdiffusion >>
rect 213 89 214 90 
<< pdiffusion >>
rect 214 89 215 90 
<< pdiffusion >>
rect 215 89 216 90 
<< m1 >>
rect 220 89 221 90 
<< m1 >>
rect 224 89 225 90 
<< m1 >>
rect 226 89 227 90 
<< pdiffusion >>
rect 228 89 229 90 
<< pdiffusion >>
rect 229 89 230 90 
<< pdiffusion >>
rect 230 89 231 90 
<< pdiffusion >>
rect 231 89 232 90 
<< pdiffusion >>
rect 232 89 233 90 
<< pdiffusion >>
rect 233 89 234 90 
<< m1 >>
rect 235 89 236 90 
<< m2 >>
rect 236 89 237 90 
<< m1 >>
rect 237 89 238 90 
<< pdiffusion >>
rect 246 89 247 90 
<< pdiffusion >>
rect 247 89 248 90 
<< pdiffusion >>
rect 248 89 249 90 
<< pdiffusion >>
rect 249 89 250 90 
<< pdiffusion >>
rect 250 89 251 90 
<< pdiffusion >>
rect 251 89 252 90 
<< m2 >>
rect 253 89 254 90 
<< m1 >>
rect 254 89 255 90 
<< m1 >>
rect 260 89 261 90 
<< m1 >>
rect 262 89 263 90 
<< pdiffusion >>
rect 264 89 265 90 
<< pdiffusion >>
rect 265 89 266 90 
<< pdiffusion >>
rect 266 89 267 90 
<< pdiffusion >>
rect 267 89 268 90 
<< pdiffusion >>
rect 268 89 269 90 
<< pdiffusion >>
rect 269 89 270 90 
<< m1 >>
rect 271 89 272 90 
<< m1 >>
rect 273 89 274 90 
<< m1 >>
rect 277 89 278 90 
<< m1 >>
rect 280 89 281 90 
<< pdiffusion >>
rect 282 89 283 90 
<< pdiffusion >>
rect 283 89 284 90 
<< pdiffusion >>
rect 284 89 285 90 
<< pdiffusion >>
rect 285 89 286 90 
<< pdiffusion >>
rect 286 89 287 90 
<< pdiffusion >>
rect 287 89 288 90 
<< pdiffusion >>
rect 300 89 301 90 
<< pdiffusion >>
rect 301 89 302 90 
<< pdiffusion >>
rect 302 89 303 90 
<< pdiffusion >>
rect 303 89 304 90 
<< pdiffusion >>
rect 304 89 305 90 
<< pdiffusion >>
rect 305 89 306 90 
<< m1 >>
rect 316 89 317 90 
<< pdiffusion >>
rect 318 89 319 90 
<< pdiffusion >>
rect 319 89 320 90 
<< pdiffusion >>
rect 320 89 321 90 
<< pdiffusion >>
rect 321 89 322 90 
<< m1 >>
rect 322 89 323 90 
<< pdiffusion >>
rect 322 89 323 90 
<< pdiffusion >>
rect 323 89 324 90 
<< m1 >>
rect 325 89 326 90 
<< m1 >>
rect 327 89 328 90 
<< m1 >>
rect 329 89 330 90 
<< m1 >>
rect 334 89 335 90 
<< m2 >>
rect 334 89 335 90 
<< pdiffusion >>
rect 336 89 337 90 
<< m1 >>
rect 337 89 338 90 
<< pdiffusion >>
rect 337 89 338 90 
<< pdiffusion >>
rect 338 89 339 90 
<< pdiffusion >>
rect 339 89 340 90 
<< m1 >>
rect 340 89 341 90 
<< pdiffusion >>
rect 340 89 341 90 
<< pdiffusion >>
rect 341 89 342 90 
<< m1 >>
rect 343 89 344 90 
<< m1 >>
rect 10 90 11 91 
<< m1 >>
rect 19 90 20 91 
<< m2 >>
rect 19 90 20 91 
<< m1 >>
rect 21 90 22 91 
<< m1 >>
rect 23 90 24 91 
<< m1 >>
rect 28 90 29 91 
<< m1 >>
rect 37 90 38 91 
<< m1 >>
rect 46 90 47 91 
<< m1 >>
rect 55 90 56 91 
<< m2 >>
rect 56 90 57 91 
<< m1 >>
rect 57 90 58 91 
<< m1 >>
rect 59 90 60 91 
<< m2 >>
rect 61 90 62 91 
<< m1 >>
rect 62 90 63 91 
<< m1 >>
rect 64 90 65 91 
<< m1 >>
rect 73 90 74 91 
<< m2 >>
rect 73 90 74 91 
<< m1 >>
rect 78 90 79 91 
<< m2 >>
rect 81 90 82 91 
<< m1 >>
rect 82 90 83 91 
<< m1 >>
rect 91 90 92 91 
<< m2 >>
rect 92 90 93 91 
<< m1 >>
rect 115 90 116 91 
<< m1 >>
rect 117 90 118 91 
<< m1 >>
rect 124 90 125 91 
<< m1 >>
rect 127 90 128 91 
<< m1 >>
rect 132 90 133 91 
<< m1 >>
rect 134 90 135 91 
<< m1 >>
rect 136 90 137 91 
<< m1 >>
rect 147 90 148 91 
<< m1 >>
rect 149 90 150 91 
<< m1 >>
rect 157 90 158 91 
<< m2 >>
rect 167 90 168 91 
<< m1 >>
rect 168 90 169 91 
<< m1 >>
rect 172 90 173 91 
<< m1 >>
rect 200 90 201 91 
<< m2 >>
rect 201 90 202 91 
<< m1 >>
rect 203 90 204 91 
<< m1 >>
rect 220 90 221 91 
<< m1 >>
rect 224 90 225 91 
<< m1 >>
rect 226 90 227 91 
<< m1 >>
rect 235 90 236 91 
<< m2 >>
rect 236 90 237 91 
<< m1 >>
rect 237 90 238 91 
<< m2 >>
rect 253 90 254 91 
<< m1 >>
rect 254 90 255 91 
<< m1 >>
rect 260 90 261 91 
<< m1 >>
rect 262 90 263 91 
<< m1 >>
rect 271 90 272 91 
<< m1 >>
rect 273 90 274 91 
<< m1 >>
rect 277 90 278 91 
<< m1 >>
rect 280 90 281 91 
<< m1 >>
rect 316 90 317 91 
<< m1 >>
rect 322 90 323 91 
<< m1 >>
rect 325 90 326 91 
<< m1 >>
rect 327 90 328 91 
<< m1 >>
rect 329 90 330 91 
<< m1 >>
rect 334 90 335 91 
<< m2 >>
rect 334 90 335 91 
<< m1 >>
rect 337 90 338 91 
<< m1 >>
rect 340 90 341 91 
<< m1 >>
rect 343 90 344 91 
<< m1 >>
rect 10 91 11 92 
<< m1 >>
rect 19 91 20 92 
<< m2 >>
rect 19 91 20 92 
<< m1 >>
rect 21 91 22 92 
<< m1 >>
rect 23 91 24 92 
<< m1 >>
rect 28 91 29 92 
<< m1 >>
rect 37 91 38 92 
<< m1 >>
rect 46 91 47 92 
<< m1 >>
rect 53 91 54 92 
<< m2 >>
rect 53 91 54 92 
<< m2c >>
rect 53 91 54 92 
<< m1 >>
rect 53 91 54 92 
<< m2 >>
rect 53 91 54 92 
<< m2 >>
rect 54 91 55 92 
<< m1 >>
rect 55 91 56 92 
<< m2 >>
rect 55 91 56 92 
<< m2 >>
rect 56 91 57 92 
<< m1 >>
rect 57 91 58 92 
<< m1 >>
rect 59 91 60 92 
<< m2 >>
rect 61 91 62 92 
<< m1 >>
rect 62 91 63 92 
<< m1 >>
rect 64 91 65 92 
<< m1 >>
rect 73 91 74 92 
<< m2 >>
rect 73 91 74 92 
<< m1 >>
rect 78 91 79 92 
<< m2 >>
rect 81 91 82 92 
<< m1 >>
rect 82 91 83 92 
<< m1 >>
rect 91 91 92 92 
<< m2 >>
rect 92 91 93 92 
<< m1 >>
rect 115 91 116 92 
<< m1 >>
rect 117 91 118 92 
<< m1 >>
rect 124 91 125 92 
<< m1 >>
rect 127 91 128 92 
<< m1 >>
rect 132 91 133 92 
<< m1 >>
rect 134 91 135 92 
<< m1 >>
rect 136 91 137 92 
<< m1 >>
rect 147 91 148 92 
<< m1 >>
rect 149 91 150 92 
<< m1 >>
rect 150 91 151 92 
<< m1 >>
rect 151 91 152 92 
<< m1 >>
rect 152 91 153 92 
<< m1 >>
rect 153 91 154 92 
<< m1 >>
rect 154 91 155 92 
<< m1 >>
rect 155 91 156 92 
<< m2 >>
rect 155 91 156 92 
<< m2c >>
rect 155 91 156 92 
<< m1 >>
rect 155 91 156 92 
<< m2 >>
rect 155 91 156 92 
<< m2 >>
rect 156 91 157 92 
<< m1 >>
rect 157 91 158 92 
<< m2 >>
rect 167 91 168 92 
<< m1 >>
rect 168 91 169 92 
<< m1 >>
rect 172 91 173 92 
<< m1 >>
rect 200 91 201 92 
<< m2 >>
rect 201 91 202 92 
<< m1 >>
rect 203 91 204 92 
<< m1 >>
rect 220 91 221 92 
<< m1 >>
rect 224 91 225 92 
<< m1 >>
rect 226 91 227 92 
<< m1 >>
rect 235 91 236 92 
<< m2 >>
rect 236 91 237 92 
<< m1 >>
rect 237 91 238 92 
<< m2 >>
rect 253 91 254 92 
<< m1 >>
rect 254 91 255 92 
<< m1 >>
rect 260 91 261 92 
<< m1 >>
rect 262 91 263 92 
<< m1 >>
rect 271 91 272 92 
<< m1 >>
rect 273 91 274 92 
<< m1 >>
rect 277 91 278 92 
<< m1 >>
rect 280 91 281 92 
<< m1 >>
rect 316 91 317 92 
<< m1 >>
rect 322 91 323 92 
<< m1 >>
rect 325 91 326 92 
<< m1 >>
rect 327 91 328 92 
<< m1 >>
rect 329 91 330 92 
<< m1 >>
rect 334 91 335 92 
<< m2 >>
rect 334 91 335 92 
<< m2 >>
rect 335 91 336 92 
<< m1 >>
rect 336 91 337 92 
<< m2 >>
rect 336 91 337 92 
<< m2c >>
rect 336 91 337 92 
<< m1 >>
rect 336 91 337 92 
<< m2 >>
rect 336 91 337 92 
<< m1 >>
rect 337 91 338 92 
<< m1 >>
rect 340 91 341 92 
<< m1 >>
rect 341 91 342 92 
<< m1 >>
rect 342 91 343 92 
<< m1 >>
rect 343 91 344 92 
<< m1 >>
rect 10 92 11 93 
<< m1 >>
rect 19 92 20 93 
<< m2 >>
rect 19 92 20 93 
<< m1 >>
rect 21 92 22 93 
<< m1 >>
rect 23 92 24 93 
<< m1 >>
rect 28 92 29 93 
<< m1 >>
rect 37 92 38 93 
<< m1 >>
rect 46 92 47 93 
<< m1 >>
rect 53 92 54 93 
<< m1 >>
rect 55 92 56 93 
<< m1 >>
rect 57 92 58 93 
<< m1 >>
rect 59 92 60 93 
<< m2 >>
rect 61 92 62 93 
<< m1 >>
rect 62 92 63 93 
<< m1 >>
rect 64 92 65 93 
<< m1 >>
rect 73 92 74 93 
<< m2 >>
rect 73 92 74 93 
<< m1 >>
rect 78 92 79 93 
<< m2 >>
rect 81 92 82 93 
<< m1 >>
rect 82 92 83 93 
<< m1 >>
rect 91 92 92 93 
<< m2 >>
rect 92 92 93 93 
<< m1 >>
rect 115 92 116 93 
<< m1 >>
rect 117 92 118 93 
<< m1 >>
rect 124 92 125 93 
<< m1 >>
rect 127 92 128 93 
<< m1 >>
rect 132 92 133 93 
<< m1 >>
rect 134 92 135 93 
<< m1 >>
rect 136 92 137 93 
<< m1 >>
rect 147 92 148 93 
<< m2 >>
rect 156 92 157 93 
<< m1 >>
rect 157 92 158 93 
<< m2 >>
rect 167 92 168 93 
<< m1 >>
rect 168 92 169 93 
<< m1 >>
rect 172 92 173 93 
<< m1 >>
rect 200 92 201 93 
<< m2 >>
rect 201 92 202 93 
<< m1 >>
rect 203 92 204 93 
<< m2 >>
rect 219 92 220 93 
<< m1 >>
rect 220 92 221 93 
<< m2 >>
rect 220 92 221 93 
<< m2 >>
rect 221 92 222 93 
<< m1 >>
rect 222 92 223 93 
<< m2 >>
rect 222 92 223 93 
<< m2c >>
rect 222 92 223 93 
<< m1 >>
rect 222 92 223 93 
<< m2 >>
rect 222 92 223 93 
<< m2 >>
rect 223 92 224 93 
<< m1 >>
rect 224 92 225 93 
<< m2 >>
rect 224 92 225 93 
<< m2 >>
rect 225 92 226 93 
<< m1 >>
rect 226 92 227 93 
<< m2 >>
rect 226 92 227 93 
<< m2 >>
rect 227 92 228 93 
<< m1 >>
rect 228 92 229 93 
<< m2 >>
rect 228 92 229 93 
<< m2c >>
rect 228 92 229 93 
<< m1 >>
rect 228 92 229 93 
<< m2 >>
rect 228 92 229 93 
<< m1 >>
rect 235 92 236 93 
<< m2 >>
rect 236 92 237 93 
<< m1 >>
rect 237 92 238 93 
<< m1 >>
rect 252 92 253 93 
<< m2 >>
rect 252 92 253 93 
<< m2c >>
rect 252 92 253 93 
<< m1 >>
rect 252 92 253 93 
<< m2 >>
rect 252 92 253 93 
<< m2 >>
rect 253 92 254 93 
<< m1 >>
rect 254 92 255 93 
<< m1 >>
rect 260 92 261 93 
<< m1 >>
rect 262 92 263 93 
<< m1 >>
rect 271 92 272 93 
<< m2 >>
rect 271 92 272 93 
<< m2c >>
rect 271 92 272 93 
<< m1 >>
rect 271 92 272 93 
<< m2 >>
rect 271 92 272 93 
<< m1 >>
rect 273 92 274 93 
<< m2 >>
rect 273 92 274 93 
<< m2c >>
rect 273 92 274 93 
<< m1 >>
rect 273 92 274 93 
<< m2 >>
rect 273 92 274 93 
<< m1 >>
rect 277 92 278 93 
<< m2 >>
rect 277 92 278 93 
<< m2c >>
rect 277 92 278 93 
<< m1 >>
rect 277 92 278 93 
<< m2 >>
rect 277 92 278 93 
<< m1 >>
rect 280 92 281 93 
<< m2 >>
rect 280 92 281 93 
<< m2c >>
rect 280 92 281 93 
<< m1 >>
rect 280 92 281 93 
<< m2 >>
rect 280 92 281 93 
<< m1 >>
rect 316 92 317 93 
<< m2 >>
rect 316 92 317 93 
<< m2c >>
rect 316 92 317 93 
<< m1 >>
rect 316 92 317 93 
<< m2 >>
rect 316 92 317 93 
<< m1 >>
rect 320 92 321 93 
<< m2 >>
rect 320 92 321 93 
<< m2c >>
rect 320 92 321 93 
<< m1 >>
rect 320 92 321 93 
<< m2 >>
rect 320 92 321 93 
<< m1 >>
rect 321 92 322 93 
<< m1 >>
rect 322 92 323 93 
<< m1 >>
rect 325 92 326 93 
<< m2 >>
rect 325 92 326 93 
<< m2c >>
rect 325 92 326 93 
<< m1 >>
rect 325 92 326 93 
<< m2 >>
rect 325 92 326 93 
<< m1 >>
rect 327 92 328 93 
<< m2 >>
rect 327 92 328 93 
<< m2c >>
rect 327 92 328 93 
<< m1 >>
rect 327 92 328 93 
<< m2 >>
rect 327 92 328 93 
<< m1 >>
rect 329 92 330 93 
<< m2 >>
rect 329 92 330 93 
<< m2c >>
rect 329 92 330 93 
<< m1 >>
rect 329 92 330 93 
<< m2 >>
rect 329 92 330 93 
<< m1 >>
rect 334 92 335 93 
<< m1 >>
rect 10 93 11 94 
<< m1 >>
rect 19 93 20 94 
<< m2 >>
rect 19 93 20 94 
<< m1 >>
rect 21 93 22 94 
<< m1 >>
rect 23 93 24 94 
<< m1 >>
rect 28 93 29 94 
<< m1 >>
rect 37 93 38 94 
<< m1 >>
rect 46 93 47 94 
<< m1 >>
rect 53 93 54 94 
<< m1 >>
rect 55 93 56 94 
<< m2 >>
rect 56 93 57 94 
<< m1 >>
rect 57 93 58 94 
<< m2 >>
rect 57 93 58 94 
<< m2c >>
rect 57 93 58 94 
<< m1 >>
rect 57 93 58 94 
<< m2 >>
rect 57 93 58 94 
<< m1 >>
rect 59 93 60 94 
<< m2 >>
rect 61 93 62 94 
<< m1 >>
rect 62 93 63 94 
<< m1 >>
rect 64 93 65 94 
<< m1 >>
rect 73 93 74 94 
<< m2 >>
rect 73 93 74 94 
<< m1 >>
rect 78 93 79 94 
<< m2 >>
rect 81 93 82 94 
<< m1 >>
rect 82 93 83 94 
<< m1 >>
rect 91 93 92 94 
<< m2 >>
rect 92 93 93 94 
<< m1 >>
rect 115 93 116 94 
<< m2 >>
rect 115 93 116 94 
<< m2c >>
rect 115 93 116 94 
<< m1 >>
rect 115 93 116 94 
<< m2 >>
rect 115 93 116 94 
<< m1 >>
rect 117 93 118 94 
<< m1 >>
rect 124 93 125 94 
<< m1 >>
rect 127 93 128 94 
<< m1 >>
rect 132 93 133 94 
<< m1 >>
rect 134 93 135 94 
<< m2 >>
rect 134 93 135 94 
<< m2c >>
rect 134 93 135 94 
<< m1 >>
rect 134 93 135 94 
<< m2 >>
rect 134 93 135 94 
<< m2 >>
rect 135 93 136 94 
<< m1 >>
rect 136 93 137 94 
<< m2 >>
rect 136 93 137 94 
<< m2 >>
rect 137 93 138 94 
<< m1 >>
rect 138 93 139 94 
<< m2 >>
rect 138 93 139 94 
<< m2c >>
rect 138 93 139 94 
<< m1 >>
rect 138 93 139 94 
<< m2 >>
rect 138 93 139 94 
<< m1 >>
rect 147 93 148 94 
<< m2 >>
rect 156 93 157 94 
<< m1 >>
rect 157 93 158 94 
<< m2 >>
rect 167 93 168 94 
<< m1 >>
rect 168 93 169 94 
<< m1 >>
rect 169 93 170 94 
<< m1 >>
rect 170 93 171 94 
<< m2 >>
rect 170 93 171 94 
<< m2c >>
rect 170 93 171 94 
<< m1 >>
rect 170 93 171 94 
<< m2 >>
rect 170 93 171 94 
<< m2 >>
rect 171 93 172 94 
<< m1 >>
rect 172 93 173 94 
<< m2 >>
rect 172 93 173 94 
<< m2 >>
rect 173 93 174 94 
<< m1 >>
rect 174 93 175 94 
<< m2 >>
rect 174 93 175 94 
<< m2c >>
rect 174 93 175 94 
<< m1 >>
rect 174 93 175 94 
<< m2 >>
rect 174 93 175 94 
<< m1 >>
rect 200 93 201 94 
<< m2 >>
rect 201 93 202 94 
<< m1 >>
rect 203 93 204 94 
<< m2 >>
rect 219 93 220 94 
<< m1 >>
rect 220 93 221 94 
<< m1 >>
rect 224 93 225 94 
<< m1 >>
rect 226 93 227 94 
<< m1 >>
rect 228 93 229 94 
<< m1 >>
rect 235 93 236 94 
<< m2 >>
rect 236 93 237 94 
<< m1 >>
rect 237 93 238 94 
<< m1 >>
rect 252 93 253 94 
<< m1 >>
rect 254 93 255 94 
<< m1 >>
rect 260 93 261 94 
<< m1 >>
rect 262 93 263 94 
<< m2 >>
rect 271 93 272 94 
<< m2 >>
rect 273 93 274 94 
<< m2 >>
rect 277 93 278 94 
<< m2 >>
rect 278 93 279 94 
<< m2 >>
rect 280 93 281 94 
<< m2 >>
rect 316 93 317 94 
<< m2 >>
rect 320 93 321 94 
<< m2 >>
rect 325 93 326 94 
<< m2 >>
rect 327 93 328 94 
<< m2 >>
rect 329 93 330 94 
<< m1 >>
rect 334 93 335 94 
<< m1 >>
rect 10 94 11 95 
<< m1 >>
rect 19 94 20 95 
<< m2 >>
rect 19 94 20 95 
<< m1 >>
rect 21 94 22 95 
<< m1 >>
rect 23 94 24 95 
<< m1 >>
rect 28 94 29 95 
<< m1 >>
rect 37 94 38 95 
<< m1 >>
rect 46 94 47 95 
<< m1 >>
rect 48 94 49 95 
<< m1 >>
rect 49 94 50 95 
<< m1 >>
rect 50 94 51 95 
<< m1 >>
rect 51 94 52 95 
<< m1 >>
rect 52 94 53 95 
<< m1 >>
rect 53 94 54 95 
<< m1 >>
rect 55 94 56 95 
<< m2 >>
rect 56 94 57 95 
<< m1 >>
rect 59 94 60 95 
<< m2 >>
rect 61 94 62 95 
<< m1 >>
rect 62 94 63 95 
<< m1 >>
rect 64 94 65 95 
<< m1 >>
rect 73 94 74 95 
<< m2 >>
rect 73 94 74 95 
<< m1 >>
rect 78 94 79 95 
<< m2 >>
rect 81 94 82 95 
<< m1 >>
rect 82 94 83 95 
<< m1 >>
rect 91 94 92 95 
<< m2 >>
rect 92 94 93 95 
<< m2 >>
rect 115 94 116 95 
<< m1 >>
rect 117 94 118 95 
<< m1 >>
rect 124 94 125 95 
<< m1 >>
rect 127 94 128 95 
<< m1 >>
rect 132 94 133 95 
<< m1 >>
rect 136 94 137 95 
<< m1 >>
rect 138 94 139 95 
<< m1 >>
rect 147 94 148 95 
<< m2 >>
rect 156 94 157 95 
<< m1 >>
rect 157 94 158 95 
<< m2 >>
rect 157 94 158 95 
<< m2 >>
rect 158 94 159 95 
<< m2 >>
rect 159 94 160 95 
<< m2 >>
rect 160 94 161 95 
<< m2 >>
rect 161 94 162 95 
<< m2 >>
rect 162 94 163 95 
<< m2 >>
rect 163 94 164 95 
<< m2 >>
rect 167 94 168 95 
<< m1 >>
rect 172 94 173 95 
<< m1 >>
rect 174 94 175 95 
<< m1 >>
rect 200 94 201 95 
<< m2 >>
rect 201 94 202 95 
<< m1 >>
rect 203 94 204 95 
<< m2 >>
rect 219 94 220 95 
<< m1 >>
rect 220 94 221 95 
<< m1 >>
rect 221 94 222 95 
<< m1 >>
rect 222 94 223 95 
<< m2 >>
rect 222 94 223 95 
<< m2c >>
rect 222 94 223 95 
<< m1 >>
rect 222 94 223 95 
<< m2 >>
rect 222 94 223 95 
<< m2 >>
rect 223 94 224 95 
<< m1 >>
rect 224 94 225 95 
<< m2 >>
rect 224 94 225 95 
<< m2 >>
rect 225 94 226 95 
<< m1 >>
rect 226 94 227 95 
<< m2 >>
rect 226 94 227 95 
<< m1 >>
rect 228 94 229 95 
<< m1 >>
rect 229 94 230 95 
<< m1 >>
rect 230 94 231 95 
<< m1 >>
rect 231 94 232 95 
<< m1 >>
rect 232 94 233 95 
<< m1 >>
rect 233 94 234 95 
<< m2 >>
rect 233 94 234 95 
<< m2c >>
rect 233 94 234 95 
<< m1 >>
rect 233 94 234 95 
<< m2 >>
rect 233 94 234 95 
<< m2 >>
rect 234 94 235 95 
<< m1 >>
rect 235 94 236 95 
<< m2 >>
rect 235 94 236 95 
<< m2 >>
rect 236 94 237 95 
<< m1 >>
rect 237 94 238 95 
<< m1 >>
rect 252 94 253 95 
<< m2 >>
rect 252 94 253 95 
<< m2c >>
rect 252 94 253 95 
<< m1 >>
rect 252 94 253 95 
<< m2 >>
rect 252 94 253 95 
<< m1 >>
rect 254 94 255 95 
<< m2 >>
rect 254 94 255 95 
<< m2c >>
rect 254 94 255 95 
<< m1 >>
rect 254 94 255 95 
<< m2 >>
rect 254 94 255 95 
<< m1 >>
rect 258 94 259 95 
<< m2 >>
rect 258 94 259 95 
<< m2c >>
rect 258 94 259 95 
<< m1 >>
rect 258 94 259 95 
<< m2 >>
rect 258 94 259 95 
<< m2 >>
rect 259 94 260 95 
<< m1 >>
rect 260 94 261 95 
<< m2 >>
rect 260 94 261 95 
<< m2 >>
rect 261 94 262 95 
<< m1 >>
rect 262 94 263 95 
<< m2 >>
rect 262 94 263 95 
<< m2 >>
rect 263 94 264 95 
<< m1 >>
rect 264 94 265 95 
<< m2 >>
rect 264 94 265 95 
<< m2c >>
rect 264 94 265 95 
<< m1 >>
rect 264 94 265 95 
<< m2 >>
rect 264 94 265 95 
<< m1 >>
rect 265 94 266 95 
<< m1 >>
rect 266 94 267 95 
<< m1 >>
rect 267 94 268 95 
<< m1 >>
rect 268 94 269 95 
<< m1 >>
rect 269 94 270 95 
<< m1 >>
rect 270 94 271 95 
<< m1 >>
rect 271 94 272 95 
<< m2 >>
rect 271 94 272 95 
<< m1 >>
rect 272 94 273 95 
<< m1 >>
rect 273 94 274 95 
<< m2 >>
rect 273 94 274 95 
<< m1 >>
rect 274 94 275 95 
<< m1 >>
rect 275 94 276 95 
<< m1 >>
rect 276 94 277 95 
<< m1 >>
rect 277 94 278 95 
<< m1 >>
rect 278 94 279 95 
<< m2 >>
rect 278 94 279 95 
<< m1 >>
rect 279 94 280 95 
<< m1 >>
rect 280 94 281 95 
<< m2 >>
rect 280 94 281 95 
<< m1 >>
rect 281 94 282 95 
<< m1 >>
rect 282 94 283 95 
<< m2 >>
rect 282 94 283 95 
<< m1 >>
rect 283 94 284 95 
<< m2 >>
rect 283 94 284 95 
<< m1 >>
rect 284 94 285 95 
<< m2 >>
rect 284 94 285 95 
<< m1 >>
rect 285 94 286 95 
<< m2 >>
rect 285 94 286 95 
<< m1 >>
rect 286 94 287 95 
<< m2 >>
rect 286 94 287 95 
<< m1 >>
rect 287 94 288 95 
<< m2 >>
rect 287 94 288 95 
<< m1 >>
rect 288 94 289 95 
<< m2 >>
rect 288 94 289 95 
<< m1 >>
rect 289 94 290 95 
<< m2 >>
rect 289 94 290 95 
<< m1 >>
rect 290 94 291 95 
<< m2 >>
rect 290 94 291 95 
<< m1 >>
rect 291 94 292 95 
<< m2 >>
rect 291 94 292 95 
<< m1 >>
rect 292 94 293 95 
<< m2 >>
rect 292 94 293 95 
<< m1 >>
rect 293 94 294 95 
<< m2 >>
rect 293 94 294 95 
<< m1 >>
rect 294 94 295 95 
<< m2 >>
rect 294 94 295 95 
<< m1 >>
rect 295 94 296 95 
<< m2 >>
rect 295 94 296 95 
<< m1 >>
rect 296 94 297 95 
<< m2 >>
rect 296 94 297 95 
<< m1 >>
rect 297 94 298 95 
<< m2 >>
rect 297 94 298 95 
<< m1 >>
rect 298 94 299 95 
<< m2 >>
rect 298 94 299 95 
<< m1 >>
rect 299 94 300 95 
<< m2 >>
rect 299 94 300 95 
<< m1 >>
rect 300 94 301 95 
<< m2 >>
rect 300 94 301 95 
<< m1 >>
rect 301 94 302 95 
<< m2 >>
rect 301 94 302 95 
<< m1 >>
rect 302 94 303 95 
<< m2 >>
rect 302 94 303 95 
<< m1 >>
rect 303 94 304 95 
<< m2 >>
rect 303 94 304 95 
<< m1 >>
rect 304 94 305 95 
<< m2 >>
rect 304 94 305 95 
<< m1 >>
rect 305 94 306 95 
<< m2 >>
rect 305 94 306 95 
<< m1 >>
rect 306 94 307 95 
<< m2 >>
rect 306 94 307 95 
<< m1 >>
rect 307 94 308 95 
<< m2 >>
rect 307 94 308 95 
<< m1 >>
rect 308 94 309 95 
<< m2 >>
rect 308 94 309 95 
<< m1 >>
rect 309 94 310 95 
<< m2 >>
rect 309 94 310 95 
<< m1 >>
rect 310 94 311 95 
<< m2 >>
rect 310 94 311 95 
<< m1 >>
rect 311 94 312 95 
<< m2 >>
rect 311 94 312 95 
<< m1 >>
rect 312 94 313 95 
<< m2 >>
rect 312 94 313 95 
<< m1 >>
rect 313 94 314 95 
<< m2 >>
rect 313 94 314 95 
<< m1 >>
rect 314 94 315 95 
<< m2 >>
rect 314 94 315 95 
<< m1 >>
rect 315 94 316 95 
<< m2 >>
rect 315 94 316 95 
<< m1 >>
rect 316 94 317 95 
<< m2 >>
rect 316 94 317 95 
<< m1 >>
rect 317 94 318 95 
<< m1 >>
rect 318 94 319 95 
<< m1 >>
rect 319 94 320 95 
<< m1 >>
rect 320 94 321 95 
<< m2 >>
rect 320 94 321 95 
<< m1 >>
rect 321 94 322 95 
<< m1 >>
rect 322 94 323 95 
<< m1 >>
rect 323 94 324 95 
<< m1 >>
rect 324 94 325 95 
<< m1 >>
rect 325 94 326 95 
<< m2 >>
rect 325 94 326 95 
<< m1 >>
rect 326 94 327 95 
<< m1 >>
rect 327 94 328 95 
<< m2 >>
rect 327 94 328 95 
<< m1 >>
rect 328 94 329 95 
<< m1 >>
rect 329 94 330 95 
<< m2 >>
rect 329 94 330 95 
<< m1 >>
rect 330 94 331 95 
<< m1 >>
rect 331 94 332 95 
<< m1 >>
rect 332 94 333 95 
<< m1 >>
rect 333 94 334 95 
<< m1 >>
rect 334 94 335 95 
<< m1 >>
rect 10 95 11 96 
<< m1 >>
rect 19 95 20 96 
<< m2 >>
rect 19 95 20 96 
<< m1 >>
rect 21 95 22 96 
<< m1 >>
rect 23 95 24 96 
<< m1 >>
rect 28 95 29 96 
<< m1 >>
rect 37 95 38 96 
<< m1 >>
rect 46 95 47 96 
<< m1 >>
rect 48 95 49 96 
<< m1 >>
rect 55 95 56 96 
<< m2 >>
rect 56 95 57 96 
<< m1 >>
rect 59 95 60 96 
<< m2 >>
rect 61 95 62 96 
<< m1 >>
rect 62 95 63 96 
<< m1 >>
rect 64 95 65 96 
<< m1 >>
rect 73 95 74 96 
<< m2 >>
rect 73 95 74 96 
<< m1 >>
rect 78 95 79 96 
<< m2 >>
rect 81 95 82 96 
<< m1 >>
rect 82 95 83 96 
<< m1 >>
rect 91 95 92 96 
<< m2 >>
rect 92 95 93 96 
<< m1 >>
rect 109 95 110 96 
<< m2 >>
rect 109 95 110 96 
<< m2c >>
rect 109 95 110 96 
<< m1 >>
rect 109 95 110 96 
<< m2 >>
rect 109 95 110 96 
<< m1 >>
rect 110 95 111 96 
<< m1 >>
rect 111 95 112 96 
<< m1 >>
rect 112 95 113 96 
<< m1 >>
rect 113 95 114 96 
<< m1 >>
rect 114 95 115 96 
<< m1 >>
rect 115 95 116 96 
<< m2 >>
rect 115 95 116 96 
<< m1 >>
rect 116 95 117 96 
<< m1 >>
rect 117 95 118 96 
<< m1 >>
rect 124 95 125 96 
<< m1 >>
rect 127 95 128 96 
<< m1 >>
rect 132 95 133 96 
<< m1 >>
rect 136 95 137 96 
<< m2 >>
rect 136 95 137 96 
<< m2c >>
rect 136 95 137 96 
<< m1 >>
rect 136 95 137 96 
<< m2 >>
rect 136 95 137 96 
<< m1 >>
rect 138 95 139 96 
<< m1 >>
rect 139 95 140 96 
<< m1 >>
rect 140 95 141 96 
<< m1 >>
rect 141 95 142 96 
<< m1 >>
rect 142 95 143 96 
<< m1 >>
rect 143 95 144 96 
<< m1 >>
rect 144 95 145 96 
<< m1 >>
rect 145 95 146 96 
<< m2 >>
rect 145 95 146 96 
<< m2c >>
rect 145 95 146 96 
<< m1 >>
rect 145 95 146 96 
<< m2 >>
rect 145 95 146 96 
<< m1 >>
rect 147 95 148 96 
<< m2 >>
rect 147 95 148 96 
<< m2c >>
rect 147 95 148 96 
<< m1 >>
rect 147 95 148 96 
<< m2 >>
rect 147 95 148 96 
<< m1 >>
rect 157 95 158 96 
<< m1 >>
rect 158 95 159 96 
<< m1 >>
rect 159 95 160 96 
<< m1 >>
rect 160 95 161 96 
<< m1 >>
rect 161 95 162 96 
<< m1 >>
rect 162 95 163 96 
<< m1 >>
rect 163 95 164 96 
<< m2 >>
rect 163 95 164 96 
<< m1 >>
rect 164 95 165 96 
<< m1 >>
rect 165 95 166 96 
<< m1 >>
rect 166 95 167 96 
<< m1 >>
rect 167 95 168 96 
<< m2 >>
rect 167 95 168 96 
<< m1 >>
rect 168 95 169 96 
<< m1 >>
rect 169 95 170 96 
<< m1 >>
rect 170 95 171 96 
<< m2 >>
rect 170 95 171 96 
<< m2c >>
rect 170 95 171 96 
<< m1 >>
rect 170 95 171 96 
<< m2 >>
rect 170 95 171 96 
<< m1 >>
rect 172 95 173 96 
<< m2 >>
rect 172 95 173 96 
<< m2c >>
rect 172 95 173 96 
<< m1 >>
rect 172 95 173 96 
<< m2 >>
rect 172 95 173 96 
<< m1 >>
rect 174 95 175 96 
<< m1 >>
rect 175 95 176 96 
<< m1 >>
rect 176 95 177 96 
<< m1 >>
rect 177 95 178 96 
<< m1 >>
rect 178 95 179 96 
<< m2 >>
rect 178 95 179 96 
<< m2c >>
rect 178 95 179 96 
<< m1 >>
rect 178 95 179 96 
<< m2 >>
rect 178 95 179 96 
<< m1 >>
rect 199 95 200 96 
<< m2 >>
rect 199 95 200 96 
<< m2c >>
rect 199 95 200 96 
<< m1 >>
rect 199 95 200 96 
<< m2 >>
rect 199 95 200 96 
<< m1 >>
rect 200 95 201 96 
<< m2 >>
rect 201 95 202 96 
<< m1 >>
rect 203 95 204 96 
<< m2 >>
rect 203 95 204 96 
<< m2c >>
rect 203 95 204 96 
<< m1 >>
rect 203 95 204 96 
<< m2 >>
rect 203 95 204 96 
<< m2 >>
rect 219 95 220 96 
<< m1 >>
rect 224 95 225 96 
<< m1 >>
rect 226 95 227 96 
<< m2 >>
rect 226 95 227 96 
<< m1 >>
rect 235 95 236 96 
<< m1 >>
rect 237 95 238 96 
<< m2 >>
rect 252 95 253 96 
<< m2 >>
rect 254 95 255 96 
<< m1 >>
rect 258 95 259 96 
<< m1 >>
rect 260 95 261 96 
<< m1 >>
rect 262 95 263 96 
<< m2 >>
rect 271 95 272 96 
<< m2 >>
rect 273 95 274 96 
<< m2 >>
rect 278 95 279 96 
<< m2 >>
rect 280 95 281 96 
<< m2 >>
rect 282 95 283 96 
<< m2 >>
rect 316 95 317 96 
<< m2 >>
rect 317 95 318 96 
<< m2 >>
rect 318 95 319 96 
<< m2 >>
rect 319 95 320 96 
<< m2 >>
rect 320 95 321 96 
<< m2 >>
rect 325 95 326 96 
<< m2 >>
rect 327 95 328 96 
<< m2 >>
rect 329 95 330 96 
<< m1 >>
rect 10 96 11 97 
<< m1 >>
rect 19 96 20 97 
<< m2 >>
rect 19 96 20 97 
<< m1 >>
rect 21 96 22 97 
<< m1 >>
rect 23 96 24 97 
<< m1 >>
rect 28 96 29 97 
<< m1 >>
rect 37 96 38 97 
<< m1 >>
rect 46 96 47 97 
<< m2 >>
rect 46 96 47 97 
<< m2c >>
rect 46 96 47 97 
<< m1 >>
rect 46 96 47 97 
<< m2 >>
rect 46 96 47 97 
<< m2 >>
rect 47 96 48 97 
<< m1 >>
rect 48 96 49 97 
<< m2 >>
rect 48 96 49 97 
<< m2 >>
rect 49 96 50 97 
<< m1 >>
rect 50 96 51 97 
<< m2 >>
rect 50 96 51 97 
<< m2c >>
rect 50 96 51 97 
<< m1 >>
rect 50 96 51 97 
<< m2 >>
rect 50 96 51 97 
<< m1 >>
rect 55 96 56 97 
<< m2 >>
rect 56 96 57 97 
<< m1 >>
rect 59 96 60 97 
<< m2 >>
rect 61 96 62 97 
<< m1 >>
rect 62 96 63 97 
<< m1 >>
rect 64 96 65 97 
<< m1 >>
rect 73 96 74 97 
<< m2 >>
rect 73 96 74 97 
<< m1 >>
rect 78 96 79 97 
<< m2 >>
rect 81 96 82 97 
<< m1 >>
rect 82 96 83 97 
<< m1 >>
rect 91 96 92 97 
<< m2 >>
rect 92 96 93 97 
<< m2 >>
rect 109 96 110 97 
<< m2 >>
rect 115 96 116 97 
<< m1 >>
rect 124 96 125 97 
<< m1 >>
rect 127 96 128 97 
<< m1 >>
rect 132 96 133 97 
<< m2 >>
rect 136 96 137 97 
<< m2 >>
rect 145 96 146 97 
<< m2 >>
rect 147 96 148 97 
<< m2 >>
rect 163 96 164 97 
<< m2 >>
rect 167 96 168 97 
<< m2 >>
rect 170 96 171 97 
<< m2 >>
rect 172 96 173 97 
<< m2 >>
rect 178 96 179 97 
<< m2 >>
rect 199 96 200 97 
<< m2 >>
rect 201 96 202 97 
<< m2 >>
rect 203 96 204 97 
<< m2 >>
rect 210 96 211 97 
<< m2 >>
rect 211 96 212 97 
<< m2 >>
rect 212 96 213 97 
<< m2 >>
rect 213 96 214 97 
<< m2 >>
rect 214 96 215 97 
<< m2 >>
rect 215 96 216 97 
<< m1 >>
rect 216 96 217 97 
<< m2 >>
rect 216 96 217 97 
<< m2c >>
rect 216 96 217 97 
<< m1 >>
rect 216 96 217 97 
<< m2 >>
rect 216 96 217 97 
<< m1 >>
rect 217 96 218 97 
<< m1 >>
rect 218 96 219 97 
<< m1 >>
rect 219 96 220 97 
<< m2 >>
rect 219 96 220 97 
<< m1 >>
rect 220 96 221 97 
<< m1 >>
rect 221 96 222 97 
<< m1 >>
rect 222 96 223 97 
<< m1 >>
rect 223 96 224 97 
<< m1 >>
rect 224 96 225 97 
<< m1 >>
rect 226 96 227 97 
<< m2 >>
rect 226 96 227 97 
<< m1 >>
rect 235 96 236 97 
<< m1 >>
rect 237 96 238 97 
<< m1 >>
rect 238 96 239 97 
<< m1 >>
rect 239 96 240 97 
<< m1 >>
rect 240 96 241 97 
<< m1 >>
rect 241 96 242 97 
<< m1 >>
rect 242 96 243 97 
<< m1 >>
rect 243 96 244 97 
<< m1 >>
rect 244 96 245 97 
<< m1 >>
rect 245 96 246 97 
<< m1 >>
rect 246 96 247 97 
<< m1 >>
rect 247 96 248 97 
<< m1 >>
rect 248 96 249 97 
<< m1 >>
rect 249 96 250 97 
<< m1 >>
rect 250 96 251 97 
<< m1 >>
rect 251 96 252 97 
<< m1 >>
rect 252 96 253 97 
<< m2 >>
rect 252 96 253 97 
<< m1 >>
rect 253 96 254 97 
<< m1 >>
rect 254 96 255 97 
<< m2 >>
rect 254 96 255 97 
<< m1 >>
rect 255 96 256 97 
<< m1 >>
rect 256 96 257 97 
<< m2 >>
rect 256 96 257 97 
<< m2c >>
rect 256 96 257 97 
<< m1 >>
rect 256 96 257 97 
<< m2 >>
rect 256 96 257 97 
<< m2 >>
rect 257 96 258 97 
<< m1 >>
rect 258 96 259 97 
<< m2 >>
rect 258 96 259 97 
<< m2 >>
rect 259 96 260 97 
<< m1 >>
rect 260 96 261 97 
<< m2 >>
rect 260 96 261 97 
<< m2 >>
rect 261 96 262 97 
<< m1 >>
rect 262 96 263 97 
<< m2 >>
rect 262 96 263 97 
<< m2 >>
rect 263 96 264 97 
<< m1 >>
rect 264 96 265 97 
<< m2 >>
rect 264 96 265 97 
<< m2c >>
rect 264 96 265 97 
<< m1 >>
rect 264 96 265 97 
<< m2 >>
rect 264 96 265 97 
<< m1 >>
rect 265 96 266 97 
<< m1 >>
rect 266 96 267 97 
<< m1 >>
rect 267 96 268 97 
<< m1 >>
rect 268 96 269 97 
<< m1 >>
rect 269 96 270 97 
<< m1 >>
rect 270 96 271 97 
<< m1 >>
rect 271 96 272 97 
<< m2 >>
rect 271 96 272 97 
<< m1 >>
rect 272 96 273 97 
<< m1 >>
rect 273 96 274 97 
<< m2 >>
rect 273 96 274 97 
<< m1 >>
rect 274 96 275 97 
<< m2 >>
rect 274 96 275 97 
<< m2 >>
rect 275 96 276 97 
<< m1 >>
rect 276 96 277 97 
<< m2 >>
rect 276 96 277 97 
<< m2c >>
rect 276 96 277 97 
<< m1 >>
rect 276 96 277 97 
<< m2 >>
rect 276 96 277 97 
<< m1 >>
rect 278 96 279 97 
<< m2 >>
rect 278 96 279 97 
<< m2c >>
rect 278 96 279 97 
<< m1 >>
rect 278 96 279 97 
<< m2 >>
rect 278 96 279 97 
<< m1 >>
rect 280 96 281 97 
<< m2 >>
rect 280 96 281 97 
<< m2c >>
rect 280 96 281 97 
<< m1 >>
rect 280 96 281 97 
<< m2 >>
rect 280 96 281 97 
<< m1 >>
rect 281 96 282 97 
<< m1 >>
rect 282 96 283 97 
<< m2 >>
rect 282 96 283 97 
<< m1 >>
rect 283 96 284 97 
<< m1 >>
rect 284 96 285 97 
<< m1 >>
rect 285 96 286 97 
<< m1 >>
rect 286 96 287 97 
<< m1 >>
rect 287 96 288 97 
<< m1 >>
rect 288 96 289 97 
<< m1 >>
rect 289 96 290 97 
<< m1 >>
rect 290 96 291 97 
<< m1 >>
rect 291 96 292 97 
<< m1 >>
rect 292 96 293 97 
<< m1 >>
rect 293 96 294 97 
<< m1 >>
rect 294 96 295 97 
<< m1 >>
rect 295 96 296 97 
<< m1 >>
rect 296 96 297 97 
<< m2 >>
rect 296 96 297 97 
<< m1 >>
rect 297 96 298 97 
<< m2 >>
rect 297 96 298 97 
<< m1 >>
rect 298 96 299 97 
<< m2 >>
rect 298 96 299 97 
<< m1 >>
rect 299 96 300 97 
<< m2 >>
rect 299 96 300 97 
<< m1 >>
rect 300 96 301 97 
<< m2 >>
rect 300 96 301 97 
<< m1 >>
rect 301 96 302 97 
<< m2 >>
rect 301 96 302 97 
<< m1 >>
rect 302 96 303 97 
<< m2 >>
rect 302 96 303 97 
<< m1 >>
rect 303 96 304 97 
<< m2 >>
rect 303 96 304 97 
<< m1 >>
rect 304 96 305 97 
<< m2 >>
rect 304 96 305 97 
<< m1 >>
rect 305 96 306 97 
<< m2 >>
rect 305 96 306 97 
<< m1 >>
rect 306 96 307 97 
<< m2 >>
rect 306 96 307 97 
<< m1 >>
rect 307 96 308 97 
<< m2 >>
rect 307 96 308 97 
<< m2 >>
rect 308 96 309 97 
<< m1 >>
rect 309 96 310 97 
<< m2 >>
rect 309 96 310 97 
<< m2c >>
rect 309 96 310 97 
<< m1 >>
rect 309 96 310 97 
<< m2 >>
rect 309 96 310 97 
<< m1 >>
rect 310 96 311 97 
<< m1 >>
rect 311 96 312 97 
<< m2 >>
rect 311 96 312 97 
<< m2c >>
rect 311 96 312 97 
<< m1 >>
rect 311 96 312 97 
<< m2 >>
rect 311 96 312 97 
<< m1 >>
rect 316 96 317 97 
<< m2 >>
rect 316 96 317 97 
<< m2c >>
rect 316 96 317 97 
<< m1 >>
rect 316 96 317 97 
<< m2 >>
rect 316 96 317 97 
<< m1 >>
rect 318 96 319 97 
<< m1 >>
rect 319 96 320 97 
<< m1 >>
rect 320 96 321 97 
<< m1 >>
rect 321 96 322 97 
<< m1 >>
rect 322 96 323 97 
<< m1 >>
rect 323 96 324 97 
<< m1 >>
rect 324 96 325 97 
<< m1 >>
rect 325 96 326 97 
<< m2 >>
rect 325 96 326 97 
<< m2c >>
rect 325 96 326 97 
<< m1 >>
rect 325 96 326 97 
<< m2 >>
rect 325 96 326 97 
<< m1 >>
rect 327 96 328 97 
<< m2 >>
rect 327 96 328 97 
<< m2c >>
rect 327 96 328 97 
<< m1 >>
rect 327 96 328 97 
<< m2 >>
rect 327 96 328 97 
<< m1 >>
rect 329 96 330 97 
<< m2 >>
rect 329 96 330 97 
<< m2c >>
rect 329 96 330 97 
<< m1 >>
rect 329 96 330 97 
<< m2 >>
rect 329 96 330 97 
<< m1 >>
rect 10 97 11 98 
<< m1 >>
rect 19 97 20 98 
<< m2 >>
rect 19 97 20 98 
<< m1 >>
rect 21 97 22 98 
<< m1 >>
rect 23 97 24 98 
<< m1 >>
rect 28 97 29 98 
<< m1 >>
rect 37 97 38 98 
<< m2 >>
rect 37 97 38 98 
<< m2c >>
rect 37 97 38 98 
<< m1 >>
rect 37 97 38 98 
<< m2 >>
rect 37 97 38 98 
<< m1 >>
rect 48 97 49 98 
<< m1 >>
rect 50 97 51 98 
<< m1 >>
rect 55 97 56 98 
<< m2 >>
rect 56 97 57 98 
<< m1 >>
rect 59 97 60 98 
<< m2 >>
rect 61 97 62 98 
<< m1 >>
rect 62 97 63 98 
<< m1 >>
rect 64 97 65 98 
<< m1 >>
rect 73 97 74 98 
<< m2 >>
rect 73 97 74 98 
<< m1 >>
rect 78 97 79 98 
<< m2 >>
rect 81 97 82 98 
<< m1 >>
rect 82 97 83 98 
<< m1 >>
rect 91 97 92 98 
<< m2 >>
rect 92 97 93 98 
<< m1 >>
rect 109 97 110 98 
<< m2 >>
rect 109 97 110 98 
<< m1 >>
rect 110 97 111 98 
<< m1 >>
rect 111 97 112 98 
<< m1 >>
rect 112 97 113 98 
<< m1 >>
rect 113 97 114 98 
<< m1 >>
rect 114 97 115 98 
<< m1 >>
rect 115 97 116 98 
<< m2 >>
rect 115 97 116 98 
<< m1 >>
rect 116 97 117 98 
<< m1 >>
rect 117 97 118 98 
<< m1 >>
rect 118 97 119 98 
<< m1 >>
rect 119 97 120 98 
<< m1 >>
rect 120 97 121 98 
<< m1 >>
rect 121 97 122 98 
<< m1 >>
rect 122 97 123 98 
<< m2 >>
rect 122 97 123 98 
<< m2c >>
rect 122 97 123 98 
<< m1 >>
rect 122 97 123 98 
<< m2 >>
rect 122 97 123 98 
<< m2 >>
rect 123 97 124 98 
<< m1 >>
rect 124 97 125 98 
<< m2 >>
rect 124 97 125 98 
<< m2 >>
rect 125 97 126 98 
<< m1 >>
rect 126 97 127 98 
<< m2 >>
rect 126 97 127 98 
<< m2c >>
rect 126 97 127 98 
<< m1 >>
rect 126 97 127 98 
<< m2 >>
rect 126 97 127 98 
<< m1 >>
rect 127 97 128 98 
<< m1 >>
rect 132 97 133 98 
<< m1 >>
rect 136 97 137 98 
<< m2 >>
rect 136 97 137 98 
<< m1 >>
rect 137 97 138 98 
<< m1 >>
rect 138 97 139 98 
<< m1 >>
rect 139 97 140 98 
<< m1 >>
rect 140 97 141 98 
<< m1 >>
rect 141 97 142 98 
<< m1 >>
rect 142 97 143 98 
<< m1 >>
rect 143 97 144 98 
<< m1 >>
rect 144 97 145 98 
<< m1 >>
rect 145 97 146 98 
<< m2 >>
rect 145 97 146 98 
<< m1 >>
rect 146 97 147 98 
<< m1 >>
rect 147 97 148 98 
<< m2 >>
rect 147 97 148 98 
<< m1 >>
rect 148 97 149 98 
<< m1 >>
rect 149 97 150 98 
<< m1 >>
rect 150 97 151 98 
<< m1 >>
rect 151 97 152 98 
<< m1 >>
rect 152 97 153 98 
<< m1 >>
rect 153 97 154 98 
<< m1 >>
rect 154 97 155 98 
<< m1 >>
rect 155 97 156 98 
<< m1 >>
rect 156 97 157 98 
<< m1 >>
rect 157 97 158 98 
<< m1 >>
rect 158 97 159 98 
<< m1 >>
rect 159 97 160 98 
<< m1 >>
rect 160 97 161 98 
<< m1 >>
rect 161 97 162 98 
<< m1 >>
rect 162 97 163 98 
<< m1 >>
rect 163 97 164 98 
<< m2 >>
rect 163 97 164 98 
<< m1 >>
rect 164 97 165 98 
<< m1 >>
rect 165 97 166 98 
<< m1 >>
rect 166 97 167 98 
<< m1 >>
rect 167 97 168 98 
<< m2 >>
rect 167 97 168 98 
<< m1 >>
rect 168 97 169 98 
<< m1 >>
rect 169 97 170 98 
<< m1 >>
rect 170 97 171 98 
<< m2 >>
rect 170 97 171 98 
<< m1 >>
rect 171 97 172 98 
<< m1 >>
rect 172 97 173 98 
<< m2 >>
rect 172 97 173 98 
<< m1 >>
rect 173 97 174 98 
<< m1 >>
rect 174 97 175 98 
<< m1 >>
rect 175 97 176 98 
<< m1 >>
rect 176 97 177 98 
<< m1 >>
rect 177 97 178 98 
<< m1 >>
rect 178 97 179 98 
<< m2 >>
rect 178 97 179 98 
<< m1 >>
rect 179 97 180 98 
<< m1 >>
rect 180 97 181 98 
<< m1 >>
rect 181 97 182 98 
<< m1 >>
rect 182 97 183 98 
<< m1 >>
rect 183 97 184 98 
<< m1 >>
rect 184 97 185 98 
<< m1 >>
rect 185 97 186 98 
<< m1 >>
rect 186 97 187 98 
<< m1 >>
rect 187 97 188 98 
<< m1 >>
rect 188 97 189 98 
<< m1 >>
rect 189 97 190 98 
<< m1 >>
rect 190 97 191 98 
<< m1 >>
rect 191 97 192 98 
<< m1 >>
rect 192 97 193 98 
<< m1 >>
rect 193 97 194 98 
<< m1 >>
rect 194 97 195 98 
<< m1 >>
rect 195 97 196 98 
<< m1 >>
rect 196 97 197 98 
<< m1 >>
rect 197 97 198 98 
<< m1 >>
rect 198 97 199 98 
<< m1 >>
rect 199 97 200 98 
<< m2 >>
rect 199 97 200 98 
<< m1 >>
rect 200 97 201 98 
<< m1 >>
rect 201 97 202 98 
<< m2 >>
rect 201 97 202 98 
<< m1 >>
rect 202 97 203 98 
<< m1 >>
rect 203 97 204 98 
<< m2 >>
rect 203 97 204 98 
<< m1 >>
rect 204 97 205 98 
<< m1 >>
rect 205 97 206 98 
<< m1 >>
rect 206 97 207 98 
<< m1 >>
rect 207 97 208 98 
<< m1 >>
rect 208 97 209 98 
<< m1 >>
rect 209 97 210 98 
<< m1 >>
rect 210 97 211 98 
<< m2 >>
rect 210 97 211 98 
<< m1 >>
rect 211 97 212 98 
<< m1 >>
rect 212 97 213 98 
<< m1 >>
rect 213 97 214 98 
<< m1 >>
rect 214 97 215 98 
<< m2 >>
rect 218 97 219 98 
<< m2 >>
rect 219 97 220 98 
<< m1 >>
rect 226 97 227 98 
<< m2 >>
rect 226 97 227 98 
<< m1 >>
rect 235 97 236 98 
<< m2 >>
rect 252 97 253 98 
<< m2 >>
rect 254 97 255 98 
<< m1 >>
rect 258 97 259 98 
<< m1 >>
rect 260 97 261 98 
<< m1 >>
rect 262 97 263 98 
<< m2 >>
rect 271 97 272 98 
<< m1 >>
rect 274 97 275 98 
<< m1 >>
rect 276 97 277 98 
<< m1 >>
rect 278 97 279 98 
<< m2 >>
rect 282 97 283 98 
<< m2 >>
rect 296 97 297 98 
<< m1 >>
rect 307 97 308 98 
<< m2 >>
rect 311 97 312 98 
<< m1 >>
rect 316 97 317 98 
<< m1 >>
rect 318 97 319 98 
<< m1 >>
rect 327 97 328 98 
<< m1 >>
rect 329 97 330 98 
<< m1 >>
rect 10 98 11 99 
<< m1 >>
rect 19 98 20 99 
<< m2 >>
rect 19 98 20 99 
<< m1 >>
rect 21 98 22 99 
<< m1 >>
rect 23 98 24 99 
<< m1 >>
rect 28 98 29 99 
<< m2 >>
rect 37 98 38 99 
<< m2 >>
rect 46 98 47 99 
<< m2 >>
rect 47 98 48 99 
<< m1 >>
rect 48 98 49 99 
<< m2 >>
rect 48 98 49 99 
<< m2c >>
rect 48 98 49 99 
<< m1 >>
rect 48 98 49 99 
<< m2 >>
rect 48 98 49 99 
<< m1 >>
rect 50 98 51 99 
<< m1 >>
rect 55 98 56 99 
<< m2 >>
rect 56 98 57 99 
<< m1 >>
rect 59 98 60 99 
<< m2 >>
rect 61 98 62 99 
<< m1 >>
rect 62 98 63 99 
<< m1 >>
rect 64 98 65 99 
<< m1 >>
rect 73 98 74 99 
<< m2 >>
rect 73 98 74 99 
<< m1 >>
rect 78 98 79 99 
<< m2 >>
rect 81 98 82 99 
<< m1 >>
rect 82 98 83 99 
<< m1 >>
rect 91 98 92 99 
<< m2 >>
rect 92 98 93 99 
<< m1 >>
rect 109 98 110 99 
<< m2 >>
rect 109 98 110 99 
<< m2 >>
rect 115 98 116 99 
<< m1 >>
rect 124 98 125 99 
<< m1 >>
rect 132 98 133 99 
<< m1 >>
rect 136 98 137 99 
<< m2 >>
rect 136 98 137 99 
<< m2 >>
rect 145 98 146 99 
<< m2 >>
rect 147 98 148 99 
<< m2 >>
rect 163 98 164 99 
<< m2 >>
rect 167 98 168 99 
<< m2 >>
rect 170 98 171 99 
<< m2 >>
rect 172 98 173 99 
<< m2 >>
rect 178 98 179 99 
<< m2 >>
rect 199 98 200 99 
<< m2 >>
rect 201 98 202 99 
<< m2 >>
rect 203 98 204 99 
<< m2 >>
rect 210 98 211 99 
<< m1 >>
rect 214 98 215 99 
<< m1 >>
rect 218 98 219 99 
<< m2 >>
rect 218 98 219 99 
<< m2c >>
rect 218 98 219 99 
<< m1 >>
rect 218 98 219 99 
<< m2 >>
rect 218 98 219 99 
<< m1 >>
rect 226 98 227 99 
<< m2 >>
rect 226 98 227 99 
<< m1 >>
rect 235 98 236 99 
<< m1 >>
rect 252 98 253 99 
<< m2 >>
rect 252 98 253 99 
<< m2c >>
rect 252 98 253 99 
<< m1 >>
rect 252 98 253 99 
<< m2 >>
rect 252 98 253 99 
<< m1 >>
rect 254 98 255 99 
<< m2 >>
rect 254 98 255 99 
<< m2c >>
rect 254 98 255 99 
<< m1 >>
rect 254 98 255 99 
<< m2 >>
rect 254 98 255 99 
<< m1 >>
rect 258 98 259 99 
<< m1 >>
rect 260 98 261 99 
<< m1 >>
rect 262 98 263 99 
<< m1 >>
rect 271 98 272 99 
<< m2 >>
rect 271 98 272 99 
<< m2c >>
rect 271 98 272 99 
<< m1 >>
rect 271 98 272 99 
<< m2 >>
rect 271 98 272 99 
<< m1 >>
rect 274 98 275 99 
<< m1 >>
rect 276 98 277 99 
<< m1 >>
rect 278 98 279 99 
<< m2 >>
rect 279 98 280 99 
<< m1 >>
rect 280 98 281 99 
<< m2 >>
rect 280 98 281 99 
<< m2c >>
rect 280 98 281 99 
<< m1 >>
rect 280 98 281 99 
<< m2 >>
rect 280 98 281 99 
<< m1 >>
rect 281 98 282 99 
<< m1 >>
rect 282 98 283 99 
<< m2 >>
rect 282 98 283 99 
<< m2c >>
rect 282 98 283 99 
<< m1 >>
rect 282 98 283 99 
<< m2 >>
rect 282 98 283 99 
<< m1 >>
rect 296 98 297 99 
<< m2 >>
rect 296 98 297 99 
<< m2c >>
rect 296 98 297 99 
<< m1 >>
rect 296 98 297 99 
<< m2 >>
rect 296 98 297 99 
<< m1 >>
rect 307 98 308 99 
<< m2 >>
rect 308 98 309 99 
<< m1 >>
rect 309 98 310 99 
<< m2 >>
rect 309 98 310 99 
<< m2c >>
rect 309 98 310 99 
<< m1 >>
rect 309 98 310 99 
<< m2 >>
rect 309 98 310 99 
<< m1 >>
rect 310 98 311 99 
<< m1 >>
rect 311 98 312 99 
<< m2 >>
rect 311 98 312 99 
<< m1 >>
rect 312 98 313 99 
<< m1 >>
rect 313 98 314 99 
<< m1 >>
rect 314 98 315 99 
<< m2 >>
rect 314 98 315 99 
<< m2c >>
rect 314 98 315 99 
<< m1 >>
rect 314 98 315 99 
<< m2 >>
rect 314 98 315 99 
<< m2 >>
rect 315 98 316 99 
<< m1 >>
rect 316 98 317 99 
<< m2 >>
rect 316 98 317 99 
<< m2 >>
rect 317 98 318 99 
<< m1 >>
rect 318 98 319 99 
<< m2 >>
rect 318 98 319 99 
<< m2c >>
rect 318 98 319 99 
<< m1 >>
rect 318 98 319 99 
<< m2 >>
rect 318 98 319 99 
<< m1 >>
rect 327 98 328 99 
<< m1 >>
rect 329 98 330 99 
<< m1 >>
rect 10 99 11 100 
<< m1 >>
rect 19 99 20 100 
<< m2 >>
rect 19 99 20 100 
<< m1 >>
rect 21 99 22 100 
<< m1 >>
rect 23 99 24 100 
<< m1 >>
rect 28 99 29 100 
<< m1 >>
rect 31 99 32 100 
<< m1 >>
rect 32 99 33 100 
<< m1 >>
rect 33 99 34 100 
<< m1 >>
rect 34 99 35 100 
<< m1 >>
rect 35 99 36 100 
<< m1 >>
rect 36 99 37 100 
<< m1 >>
rect 37 99 38 100 
<< m2 >>
rect 37 99 38 100 
<< m1 >>
rect 38 99 39 100 
<< m1 >>
rect 39 99 40 100 
<< m1 >>
rect 40 99 41 100 
<< m1 >>
rect 41 99 42 100 
<< m1 >>
rect 42 99 43 100 
<< m1 >>
rect 43 99 44 100 
<< m1 >>
rect 44 99 45 100 
<< m1 >>
rect 45 99 46 100 
<< m1 >>
rect 46 99 47 100 
<< m2 >>
rect 46 99 47 100 
<< m1 >>
rect 50 99 51 100 
<< m1 >>
rect 55 99 56 100 
<< m2 >>
rect 56 99 57 100 
<< m1 >>
rect 59 99 60 100 
<< m2 >>
rect 61 99 62 100 
<< m1 >>
rect 62 99 63 100 
<< m1 >>
rect 64 99 65 100 
<< m1 >>
rect 73 99 74 100 
<< m2 >>
rect 73 99 74 100 
<< m1 >>
rect 78 99 79 100 
<< m2 >>
rect 81 99 82 100 
<< m1 >>
rect 82 99 83 100 
<< m1 >>
rect 91 99 92 100 
<< m2 >>
rect 92 99 93 100 
<< m1 >>
rect 109 99 110 100 
<< m2 >>
rect 109 99 110 100 
<< m1 >>
rect 115 99 116 100 
<< m2 >>
rect 115 99 116 100 
<< m2c >>
rect 115 99 116 100 
<< m1 >>
rect 115 99 116 100 
<< m2 >>
rect 115 99 116 100 
<< m1 >>
rect 124 99 125 100 
<< m1 >>
rect 125 99 126 100 
<< m1 >>
rect 126 99 127 100 
<< m1 >>
rect 127 99 128 100 
<< m1 >>
rect 128 99 129 100 
<< m1 >>
rect 129 99 130 100 
<< m1 >>
rect 130 99 131 100 
<< m1 >>
rect 132 99 133 100 
<< m1 >>
rect 136 99 137 100 
<< m2 >>
rect 136 99 137 100 
<< m2 >>
rect 145 99 146 100 
<< m1 >>
rect 147 99 148 100 
<< m2 >>
rect 147 99 148 100 
<< m2c >>
rect 147 99 148 100 
<< m1 >>
rect 147 99 148 100 
<< m2 >>
rect 147 99 148 100 
<< m2 >>
rect 163 99 164 100 
<< m2 >>
rect 167 99 168 100 
<< m2 >>
rect 170 99 171 100 
<< m2 >>
rect 172 99 173 100 
<< m1 >>
rect 178 99 179 100 
<< m2 >>
rect 178 99 179 100 
<< m2c >>
rect 178 99 179 100 
<< m1 >>
rect 178 99 179 100 
<< m2 >>
rect 178 99 179 100 
<< m1 >>
rect 199 99 200 100 
<< m2 >>
rect 199 99 200 100 
<< m2c >>
rect 199 99 200 100 
<< m1 >>
rect 199 99 200 100 
<< m2 >>
rect 199 99 200 100 
<< m1 >>
rect 201 99 202 100 
<< m2 >>
rect 201 99 202 100 
<< m2c >>
rect 201 99 202 100 
<< m1 >>
rect 201 99 202 100 
<< m2 >>
rect 201 99 202 100 
<< m1 >>
rect 203 99 204 100 
<< m2 >>
rect 203 99 204 100 
<< m2c >>
rect 203 99 204 100 
<< m1 >>
rect 203 99 204 100 
<< m2 >>
rect 203 99 204 100 
<< m1 >>
rect 204 99 205 100 
<< m1 >>
rect 205 99 206 100 
<< m2 >>
rect 205 99 206 100 
<< m2c >>
rect 205 99 206 100 
<< m1 >>
rect 205 99 206 100 
<< m2 >>
rect 205 99 206 100 
<< m1 >>
rect 208 99 209 100 
<< m1 >>
rect 209 99 210 100 
<< m1 >>
rect 210 99 211 100 
<< m2 >>
rect 210 99 211 100 
<< m2c >>
rect 210 99 211 100 
<< m1 >>
rect 210 99 211 100 
<< m2 >>
rect 210 99 211 100 
<< m1 >>
rect 214 99 215 100 
<< m1 >>
rect 218 99 219 100 
<< m1 >>
rect 226 99 227 100 
<< m2 >>
rect 226 99 227 100 
<< m1 >>
rect 235 99 236 100 
<< m1 >>
rect 252 99 253 100 
<< m1 >>
rect 254 99 255 100 
<< m1 >>
rect 258 99 259 100 
<< m1 >>
rect 260 99 261 100 
<< m1 >>
rect 262 99 263 100 
<< m1 >>
rect 271 99 272 100 
<< m1 >>
rect 274 99 275 100 
<< m1 >>
rect 276 99 277 100 
<< m1 >>
rect 278 99 279 100 
<< m2 >>
rect 279 99 280 100 
<< m1 >>
rect 296 99 297 100 
<< m1 >>
rect 307 99 308 100 
<< m2 >>
rect 308 99 309 100 
<< m2 >>
rect 311 99 312 100 
<< m1 >>
rect 316 99 317 100 
<< m1 >>
rect 327 99 328 100 
<< m1 >>
rect 329 99 330 100 
<< m1 >>
rect 10 100 11 101 
<< m1 >>
rect 19 100 20 101 
<< m2 >>
rect 19 100 20 101 
<< m1 >>
rect 21 100 22 101 
<< m1 >>
rect 23 100 24 101 
<< m1 >>
rect 28 100 29 101 
<< m1 >>
rect 31 100 32 101 
<< m2 >>
rect 37 100 38 101 
<< m1 >>
rect 46 100 47 101 
<< m2 >>
rect 46 100 47 101 
<< m1 >>
rect 49 100 50 101 
<< m1 >>
rect 50 100 51 101 
<< m1 >>
rect 55 100 56 101 
<< m2 >>
rect 56 100 57 101 
<< m1 >>
rect 59 100 60 101 
<< m2 >>
rect 61 100 62 101 
<< m1 >>
rect 62 100 63 101 
<< m1 >>
rect 64 100 65 101 
<< m1 >>
rect 73 100 74 101 
<< m2 >>
rect 73 100 74 101 
<< m1 >>
rect 78 100 79 101 
<< m2 >>
rect 81 100 82 101 
<< m1 >>
rect 82 100 83 101 
<< m1 >>
rect 91 100 92 101 
<< m2 >>
rect 92 100 93 101 
<< m1 >>
rect 109 100 110 101 
<< m2 >>
rect 109 100 110 101 
<< m1 >>
rect 115 100 116 101 
<< m1 >>
rect 130 100 131 101 
<< m1 >>
rect 132 100 133 101 
<< m1 >>
rect 136 100 137 101 
<< m2 >>
rect 136 100 137 101 
<< m1 >>
rect 142 100 143 101 
<< m1 >>
rect 143 100 144 101 
<< m1 >>
rect 144 100 145 101 
<< m1 >>
rect 145 100 146 101 
<< m2 >>
rect 145 100 146 101 
<< m1 >>
rect 147 100 148 101 
<< m1 >>
rect 163 100 164 101 
<< m2 >>
rect 163 100 164 101 
<< m1 >>
rect 164 100 165 101 
<< m1 >>
rect 165 100 166 101 
<< m1 >>
rect 166 100 167 101 
<< m1 >>
rect 167 100 168 101 
<< m2 >>
rect 167 100 168 101 
<< m1 >>
rect 168 100 169 101 
<< m1 >>
rect 169 100 170 101 
<< m1 >>
rect 170 100 171 101 
<< m2 >>
rect 170 100 171 101 
<< m1 >>
rect 171 100 172 101 
<< m1 >>
rect 172 100 173 101 
<< m2 >>
rect 172 100 173 101 
<< m1 >>
rect 173 100 174 101 
<< m1 >>
rect 174 100 175 101 
<< m1 >>
rect 175 100 176 101 
<< m1 >>
rect 178 100 179 101 
<< m1 >>
rect 190 100 191 101 
<< m1 >>
rect 191 100 192 101 
<< m1 >>
rect 192 100 193 101 
<< m1 >>
rect 193 100 194 101 
<< m1 >>
rect 199 100 200 101 
<< m1 >>
rect 201 100 202 101 
<< m2 >>
rect 205 100 206 101 
<< m1 >>
rect 208 100 209 101 
<< m1 >>
rect 214 100 215 101 
<< m1 >>
rect 218 100 219 101 
<< m1 >>
rect 226 100 227 101 
<< m2 >>
rect 226 100 227 101 
<< m1 >>
rect 232 100 233 101 
<< m1 >>
rect 233 100 234 101 
<< m2 >>
rect 233 100 234 101 
<< m2c >>
rect 233 100 234 101 
<< m1 >>
rect 233 100 234 101 
<< m2 >>
rect 233 100 234 101 
<< m2 >>
rect 234 100 235 101 
<< m1 >>
rect 235 100 236 101 
<< m2 >>
rect 235 100 236 101 
<< m2 >>
rect 236 100 237 101 
<< m1 >>
rect 252 100 253 101 
<< m2 >>
rect 252 100 253 101 
<< m2c >>
rect 252 100 253 101 
<< m1 >>
rect 252 100 253 101 
<< m2 >>
rect 252 100 253 101 
<< m2 >>
rect 253 100 254 101 
<< m1 >>
rect 254 100 255 101 
<< m2 >>
rect 254 100 255 101 
<< m2 >>
rect 255 100 256 101 
<< m1 >>
rect 258 100 259 101 
<< m1 >>
rect 260 100 261 101 
<< m1 >>
rect 262 100 263 101 
<< m1 >>
rect 271 100 272 101 
<< m1 >>
rect 274 100 275 101 
<< m1 >>
rect 276 100 277 101 
<< m1 >>
rect 278 100 279 101 
<< m2 >>
rect 279 100 280 101 
<< m1 >>
rect 296 100 297 101 
<< m1 >>
rect 307 100 308 101 
<< m2 >>
rect 308 100 309 101 
<< m1 >>
rect 311 100 312 101 
<< m2 >>
rect 311 100 312 101 
<< m2c >>
rect 311 100 312 101 
<< m1 >>
rect 311 100 312 101 
<< m2 >>
rect 311 100 312 101 
<< m1 >>
rect 312 100 313 101 
<< m1 >>
rect 313 100 314 101 
<< m1 >>
rect 314 100 315 101 
<< m2 >>
rect 314 100 315 101 
<< m2c >>
rect 314 100 315 101 
<< m1 >>
rect 314 100 315 101 
<< m2 >>
rect 314 100 315 101 
<< m2 >>
rect 315 100 316 101 
<< m1 >>
rect 316 100 317 101 
<< m1 >>
rect 327 100 328 101 
<< m1 >>
rect 329 100 330 101 
<< m1 >>
rect 10 101 11 102 
<< m1 >>
rect 19 101 20 102 
<< m2 >>
rect 19 101 20 102 
<< m1 >>
rect 21 101 22 102 
<< m1 >>
rect 23 101 24 102 
<< m1 >>
rect 28 101 29 102 
<< m1 >>
rect 31 101 32 102 
<< m1 >>
rect 37 101 38 102 
<< m2 >>
rect 37 101 38 102 
<< m2c >>
rect 37 101 38 102 
<< m1 >>
rect 37 101 38 102 
<< m2 >>
rect 37 101 38 102 
<< m1 >>
rect 44 101 45 102 
<< m2 >>
rect 44 101 45 102 
<< m2c >>
rect 44 101 45 102 
<< m1 >>
rect 44 101 45 102 
<< m2 >>
rect 44 101 45 102 
<< m2 >>
rect 45 101 46 102 
<< m1 >>
rect 46 101 47 102 
<< m2 >>
rect 46 101 47 102 
<< m1 >>
rect 49 101 50 102 
<< m1 >>
rect 55 101 56 102 
<< m2 >>
rect 56 101 57 102 
<< m1 >>
rect 59 101 60 102 
<< m2 >>
rect 61 101 62 102 
<< m1 >>
rect 62 101 63 102 
<< m1 >>
rect 64 101 65 102 
<< m1 >>
rect 73 101 74 102 
<< m2 >>
rect 73 101 74 102 
<< m1 >>
rect 78 101 79 102 
<< m2 >>
rect 81 101 82 102 
<< m1 >>
rect 82 101 83 102 
<< m1 >>
rect 91 101 92 102 
<< m2 >>
rect 92 101 93 102 
<< m1 >>
rect 109 101 110 102 
<< m2 >>
rect 109 101 110 102 
<< m1 >>
rect 115 101 116 102 
<< m1 >>
rect 130 101 131 102 
<< m1 >>
rect 132 101 133 102 
<< m1 >>
rect 136 101 137 102 
<< m2 >>
rect 136 101 137 102 
<< m1 >>
rect 142 101 143 102 
<< m1 >>
rect 145 101 146 102 
<< m2 >>
rect 145 101 146 102 
<< m1 >>
rect 147 101 148 102 
<< m1 >>
rect 163 101 164 102 
<< m2 >>
rect 163 101 164 102 
<< m2 >>
rect 167 101 168 102 
<< m2 >>
rect 170 101 171 102 
<< m2 >>
rect 172 101 173 102 
<< m1 >>
rect 175 101 176 102 
<< m1 >>
rect 178 101 179 102 
<< m1 >>
rect 190 101 191 102 
<< m1 >>
rect 193 101 194 102 
<< m1 >>
rect 199 101 200 102 
<< m1 >>
rect 201 101 202 102 
<< m2 >>
rect 202 101 203 102 
<< m1 >>
rect 203 101 204 102 
<< m2 >>
rect 203 101 204 102 
<< m2c >>
rect 203 101 204 102 
<< m1 >>
rect 203 101 204 102 
<< m2 >>
rect 203 101 204 102 
<< m1 >>
rect 204 101 205 102 
<< m1 >>
rect 205 101 206 102 
<< m2 >>
rect 205 101 206 102 
<< m1 >>
rect 206 101 207 102 
<< m1 >>
rect 207 101 208 102 
<< m1 >>
rect 208 101 209 102 
<< m1 >>
rect 214 101 215 102 
<< m1 >>
rect 218 101 219 102 
<< m1 >>
rect 226 101 227 102 
<< m2 >>
rect 226 101 227 102 
<< m1 >>
rect 232 101 233 102 
<< m1 >>
rect 235 101 236 102 
<< m2 >>
rect 236 101 237 102 
<< m1 >>
rect 254 101 255 102 
<< m2 >>
rect 255 101 256 102 
<< m1 >>
rect 258 101 259 102 
<< m1 >>
rect 260 101 261 102 
<< m1 >>
rect 262 101 263 102 
<< m1 >>
rect 271 101 272 102 
<< m1 >>
rect 274 101 275 102 
<< m1 >>
rect 276 101 277 102 
<< m1 >>
rect 278 101 279 102 
<< m2 >>
rect 279 101 280 102 
<< m1 >>
rect 296 101 297 102 
<< m1 >>
rect 307 101 308 102 
<< m2 >>
rect 308 101 309 102 
<< m2 >>
rect 315 101 316 102 
<< m1 >>
rect 316 101 317 102 
<< m1 >>
rect 327 101 328 102 
<< m1 >>
rect 329 101 330 102 
<< m1 >>
rect 10 102 11 103 
<< pdiffusion >>
rect 12 102 13 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< m1 >>
rect 19 102 20 103 
<< m2 >>
rect 19 102 20 103 
<< m1 >>
rect 21 102 22 103 
<< m1 >>
rect 23 102 24 103 
<< m1 >>
rect 28 102 29 103 
<< pdiffusion >>
rect 30 102 31 103 
<< m1 >>
rect 31 102 32 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< pdiffusion >>
rect 33 102 34 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< m1 >>
rect 37 102 38 103 
<< m1 >>
rect 44 102 45 103 
<< m1 >>
rect 46 102 47 103 
<< pdiffusion >>
rect 48 102 49 103 
<< m1 >>
rect 49 102 50 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m1 >>
rect 55 102 56 103 
<< m2 >>
rect 56 102 57 103 
<< m1 >>
rect 59 102 60 103 
<< m2 >>
rect 61 102 62 103 
<< m1 >>
rect 62 102 63 103 
<< m1 >>
rect 64 102 65 103 
<< pdiffusion >>
rect 66 102 67 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< m1 >>
rect 73 102 74 103 
<< m2 >>
rect 73 102 74 103 
<< m1 >>
rect 78 102 79 103 
<< m2 >>
rect 81 102 82 103 
<< m1 >>
rect 82 102 83 103 
<< pdiffusion >>
rect 84 102 85 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< m1 >>
rect 91 102 92 103 
<< m2 >>
rect 92 102 93 103 
<< pdiffusion >>
rect 102 102 103 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< m1 >>
rect 109 102 110 103 
<< m2 >>
rect 109 102 110 103 
<< m1 >>
rect 115 102 116 103 
<< pdiffusion >>
rect 120 102 121 103 
<< pdiffusion >>
rect 121 102 122 103 
<< pdiffusion >>
rect 122 102 123 103 
<< pdiffusion >>
rect 123 102 124 103 
<< pdiffusion >>
rect 124 102 125 103 
<< pdiffusion >>
rect 125 102 126 103 
<< m1 >>
rect 130 102 131 103 
<< m1 >>
rect 132 102 133 103 
<< m1 >>
rect 136 102 137 103 
<< m2 >>
rect 136 102 137 103 
<< pdiffusion >>
rect 138 102 139 103 
<< pdiffusion >>
rect 139 102 140 103 
<< pdiffusion >>
rect 140 102 141 103 
<< pdiffusion >>
rect 141 102 142 103 
<< m1 >>
rect 142 102 143 103 
<< pdiffusion >>
rect 142 102 143 103 
<< pdiffusion >>
rect 143 102 144 103 
<< m1 >>
rect 145 102 146 103 
<< m2 >>
rect 145 102 146 103 
<< m1 >>
rect 147 102 148 103 
<< pdiffusion >>
rect 156 102 157 103 
<< pdiffusion >>
rect 157 102 158 103 
<< pdiffusion >>
rect 158 102 159 103 
<< pdiffusion >>
rect 159 102 160 103 
<< pdiffusion >>
rect 160 102 161 103 
<< pdiffusion >>
rect 161 102 162 103 
<< m1 >>
rect 163 102 164 103 
<< m2 >>
rect 163 102 164 103 
<< m2 >>
rect 164 102 165 103 
<< m1 >>
rect 165 102 166 103 
<< m2 >>
rect 165 102 166 103 
<< m2c >>
rect 165 102 166 103 
<< m1 >>
rect 165 102 166 103 
<< m2 >>
rect 165 102 166 103 
<< m1 >>
rect 166 102 167 103 
<< m1 >>
rect 167 102 168 103 
<< m2 >>
rect 167 102 168 103 
<< m1 >>
rect 170 102 171 103 
<< m2 >>
rect 170 102 171 103 
<< m2c >>
rect 170 102 171 103 
<< m1 >>
rect 170 102 171 103 
<< m2 >>
rect 170 102 171 103 
<< m1 >>
rect 172 102 173 103 
<< m2 >>
rect 172 102 173 103 
<< m2c >>
rect 172 102 173 103 
<< m1 >>
rect 172 102 173 103 
<< m2 >>
rect 172 102 173 103 
<< pdiffusion >>
rect 174 102 175 103 
<< m1 >>
rect 175 102 176 103 
<< pdiffusion >>
rect 175 102 176 103 
<< pdiffusion >>
rect 176 102 177 103 
<< pdiffusion >>
rect 177 102 178 103 
<< m1 >>
rect 178 102 179 103 
<< pdiffusion >>
rect 178 102 179 103 
<< pdiffusion >>
rect 179 102 180 103 
<< m1 >>
rect 190 102 191 103 
<< pdiffusion >>
rect 192 102 193 103 
<< m1 >>
rect 193 102 194 103 
<< pdiffusion >>
rect 193 102 194 103 
<< pdiffusion >>
rect 194 102 195 103 
<< pdiffusion >>
rect 195 102 196 103 
<< pdiffusion >>
rect 196 102 197 103 
<< pdiffusion >>
rect 197 102 198 103 
<< m1 >>
rect 199 102 200 103 
<< m1 >>
rect 201 102 202 103 
<< m2 >>
rect 202 102 203 103 
<< m2 >>
rect 205 102 206 103 
<< pdiffusion >>
rect 210 102 211 103 
<< pdiffusion >>
rect 211 102 212 103 
<< pdiffusion >>
rect 212 102 213 103 
<< pdiffusion >>
rect 213 102 214 103 
<< m1 >>
rect 214 102 215 103 
<< pdiffusion >>
rect 214 102 215 103 
<< pdiffusion >>
rect 215 102 216 103 
<< m1 >>
rect 218 102 219 103 
<< m1 >>
rect 226 102 227 103 
<< m2 >>
rect 226 102 227 103 
<< pdiffusion >>
rect 228 102 229 103 
<< pdiffusion >>
rect 229 102 230 103 
<< pdiffusion >>
rect 230 102 231 103 
<< pdiffusion >>
rect 231 102 232 103 
<< m1 >>
rect 232 102 233 103 
<< pdiffusion >>
rect 232 102 233 103 
<< pdiffusion >>
rect 233 102 234 103 
<< m1 >>
rect 235 102 236 103 
<< m2 >>
rect 236 102 237 103 
<< pdiffusion >>
rect 246 102 247 103 
<< pdiffusion >>
rect 247 102 248 103 
<< pdiffusion >>
rect 248 102 249 103 
<< pdiffusion >>
rect 249 102 250 103 
<< pdiffusion >>
rect 250 102 251 103 
<< pdiffusion >>
rect 251 102 252 103 
<< m1 >>
rect 254 102 255 103 
<< m2 >>
rect 255 102 256 103 
<< m1 >>
rect 258 102 259 103 
<< m1 >>
rect 260 102 261 103 
<< m1 >>
rect 262 102 263 103 
<< pdiffusion >>
rect 264 102 265 103 
<< pdiffusion >>
rect 265 102 266 103 
<< pdiffusion >>
rect 266 102 267 103 
<< pdiffusion >>
rect 267 102 268 103 
<< pdiffusion >>
rect 268 102 269 103 
<< pdiffusion >>
rect 269 102 270 103 
<< m1 >>
rect 271 102 272 103 
<< m1 >>
rect 274 102 275 103 
<< m1 >>
rect 276 102 277 103 
<< m1 >>
rect 278 102 279 103 
<< m2 >>
rect 279 102 280 103 
<< pdiffusion >>
rect 282 102 283 103 
<< pdiffusion >>
rect 283 102 284 103 
<< pdiffusion >>
rect 284 102 285 103 
<< pdiffusion >>
rect 285 102 286 103 
<< pdiffusion >>
rect 286 102 287 103 
<< pdiffusion >>
rect 287 102 288 103 
<< m1 >>
rect 296 102 297 103 
<< pdiffusion >>
rect 300 102 301 103 
<< pdiffusion >>
rect 301 102 302 103 
<< pdiffusion >>
rect 302 102 303 103 
<< pdiffusion >>
rect 303 102 304 103 
<< pdiffusion >>
rect 304 102 305 103 
<< pdiffusion >>
rect 305 102 306 103 
<< m1 >>
rect 307 102 308 103 
<< m2 >>
rect 308 102 309 103 
<< m2 >>
rect 315 102 316 103 
<< m1 >>
rect 316 102 317 103 
<< pdiffusion >>
rect 318 102 319 103 
<< pdiffusion >>
rect 319 102 320 103 
<< pdiffusion >>
rect 320 102 321 103 
<< pdiffusion >>
rect 321 102 322 103 
<< pdiffusion >>
rect 322 102 323 103 
<< pdiffusion >>
rect 323 102 324 103 
<< m1 >>
rect 327 102 328 103 
<< m1 >>
rect 329 102 330 103 
<< pdiffusion >>
rect 336 102 337 103 
<< pdiffusion >>
rect 337 102 338 103 
<< pdiffusion >>
rect 338 102 339 103 
<< pdiffusion >>
rect 339 102 340 103 
<< pdiffusion >>
rect 340 102 341 103 
<< pdiffusion >>
rect 341 102 342 103 
<< m1 >>
rect 10 103 11 104 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< m1 >>
rect 19 103 20 104 
<< m2 >>
rect 19 103 20 104 
<< m1 >>
rect 21 103 22 104 
<< m1 >>
rect 23 103 24 104 
<< m1 >>
rect 28 103 29 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< m1 >>
rect 37 103 38 104 
<< m1 >>
rect 44 103 45 104 
<< m1 >>
rect 46 103 47 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m1 >>
rect 55 103 56 104 
<< m2 >>
rect 56 103 57 104 
<< m1 >>
rect 59 103 60 104 
<< m2 >>
rect 61 103 62 104 
<< m1 >>
rect 62 103 63 104 
<< m1 >>
rect 64 103 65 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< m1 >>
rect 73 103 74 104 
<< m2 >>
rect 73 103 74 104 
<< m1 >>
rect 78 103 79 104 
<< m2 >>
rect 81 103 82 104 
<< m1 >>
rect 82 103 83 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< m1 >>
rect 91 103 92 104 
<< m2 >>
rect 92 103 93 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< m1 >>
rect 109 103 110 104 
<< m2 >>
rect 109 103 110 104 
<< m1 >>
rect 115 103 116 104 
<< pdiffusion >>
rect 120 103 121 104 
<< pdiffusion >>
rect 121 103 122 104 
<< pdiffusion >>
rect 122 103 123 104 
<< pdiffusion >>
rect 123 103 124 104 
<< pdiffusion >>
rect 124 103 125 104 
<< pdiffusion >>
rect 125 103 126 104 
<< m1 >>
rect 130 103 131 104 
<< m1 >>
rect 132 103 133 104 
<< m1 >>
rect 136 103 137 104 
<< m2 >>
rect 136 103 137 104 
<< pdiffusion >>
rect 138 103 139 104 
<< pdiffusion >>
rect 139 103 140 104 
<< pdiffusion >>
rect 140 103 141 104 
<< pdiffusion >>
rect 141 103 142 104 
<< pdiffusion >>
rect 142 103 143 104 
<< pdiffusion >>
rect 143 103 144 104 
<< m1 >>
rect 145 103 146 104 
<< m2 >>
rect 145 103 146 104 
<< m1 >>
rect 147 103 148 104 
<< pdiffusion >>
rect 156 103 157 104 
<< pdiffusion >>
rect 157 103 158 104 
<< pdiffusion >>
rect 158 103 159 104 
<< pdiffusion >>
rect 159 103 160 104 
<< pdiffusion >>
rect 160 103 161 104 
<< pdiffusion >>
rect 161 103 162 104 
<< m1 >>
rect 163 103 164 104 
<< m1 >>
rect 167 103 168 104 
<< m2 >>
rect 167 103 168 104 
<< m1 >>
rect 170 103 171 104 
<< m1 >>
rect 172 103 173 104 
<< pdiffusion >>
rect 174 103 175 104 
<< pdiffusion >>
rect 175 103 176 104 
<< pdiffusion >>
rect 176 103 177 104 
<< pdiffusion >>
rect 177 103 178 104 
<< pdiffusion >>
rect 178 103 179 104 
<< pdiffusion >>
rect 179 103 180 104 
<< m1 >>
rect 190 103 191 104 
<< pdiffusion >>
rect 192 103 193 104 
<< pdiffusion >>
rect 193 103 194 104 
<< pdiffusion >>
rect 194 103 195 104 
<< pdiffusion >>
rect 195 103 196 104 
<< pdiffusion >>
rect 196 103 197 104 
<< pdiffusion >>
rect 197 103 198 104 
<< m1 >>
rect 199 103 200 104 
<< m1 >>
rect 201 103 202 104 
<< m2 >>
rect 202 103 203 104 
<< m1 >>
rect 205 103 206 104 
<< m2 >>
rect 205 103 206 104 
<< m2c >>
rect 205 103 206 104 
<< m1 >>
rect 205 103 206 104 
<< m2 >>
rect 205 103 206 104 
<< pdiffusion >>
rect 210 103 211 104 
<< pdiffusion >>
rect 211 103 212 104 
<< pdiffusion >>
rect 212 103 213 104 
<< pdiffusion >>
rect 213 103 214 104 
<< pdiffusion >>
rect 214 103 215 104 
<< pdiffusion >>
rect 215 103 216 104 
<< m1 >>
rect 218 103 219 104 
<< m1 >>
rect 226 103 227 104 
<< m2 >>
rect 226 103 227 104 
<< pdiffusion >>
rect 228 103 229 104 
<< pdiffusion >>
rect 229 103 230 104 
<< pdiffusion >>
rect 230 103 231 104 
<< pdiffusion >>
rect 231 103 232 104 
<< pdiffusion >>
rect 232 103 233 104 
<< pdiffusion >>
rect 233 103 234 104 
<< m1 >>
rect 235 103 236 104 
<< m2 >>
rect 236 103 237 104 
<< pdiffusion >>
rect 246 103 247 104 
<< pdiffusion >>
rect 247 103 248 104 
<< pdiffusion >>
rect 248 103 249 104 
<< pdiffusion >>
rect 249 103 250 104 
<< pdiffusion >>
rect 250 103 251 104 
<< pdiffusion >>
rect 251 103 252 104 
<< m1 >>
rect 254 103 255 104 
<< m2 >>
rect 255 103 256 104 
<< m1 >>
rect 258 103 259 104 
<< m1 >>
rect 260 103 261 104 
<< m1 >>
rect 262 103 263 104 
<< pdiffusion >>
rect 264 103 265 104 
<< pdiffusion >>
rect 265 103 266 104 
<< pdiffusion >>
rect 266 103 267 104 
<< pdiffusion >>
rect 267 103 268 104 
<< pdiffusion >>
rect 268 103 269 104 
<< pdiffusion >>
rect 269 103 270 104 
<< m1 >>
rect 271 103 272 104 
<< m1 >>
rect 274 103 275 104 
<< m1 >>
rect 276 103 277 104 
<< m1 >>
rect 278 103 279 104 
<< m2 >>
rect 279 103 280 104 
<< pdiffusion >>
rect 282 103 283 104 
<< pdiffusion >>
rect 283 103 284 104 
<< pdiffusion >>
rect 284 103 285 104 
<< pdiffusion >>
rect 285 103 286 104 
<< pdiffusion >>
rect 286 103 287 104 
<< pdiffusion >>
rect 287 103 288 104 
<< m1 >>
rect 296 103 297 104 
<< pdiffusion >>
rect 300 103 301 104 
<< pdiffusion >>
rect 301 103 302 104 
<< pdiffusion >>
rect 302 103 303 104 
<< pdiffusion >>
rect 303 103 304 104 
<< pdiffusion >>
rect 304 103 305 104 
<< pdiffusion >>
rect 305 103 306 104 
<< m1 >>
rect 307 103 308 104 
<< m2 >>
rect 308 103 309 104 
<< m2 >>
rect 315 103 316 104 
<< m1 >>
rect 316 103 317 104 
<< pdiffusion >>
rect 318 103 319 104 
<< pdiffusion >>
rect 319 103 320 104 
<< pdiffusion >>
rect 320 103 321 104 
<< pdiffusion >>
rect 321 103 322 104 
<< pdiffusion >>
rect 322 103 323 104 
<< pdiffusion >>
rect 323 103 324 104 
<< m1 >>
rect 327 103 328 104 
<< m1 >>
rect 329 103 330 104 
<< pdiffusion >>
rect 336 103 337 104 
<< pdiffusion >>
rect 337 103 338 104 
<< pdiffusion >>
rect 338 103 339 104 
<< pdiffusion >>
rect 339 103 340 104 
<< pdiffusion >>
rect 340 103 341 104 
<< pdiffusion >>
rect 341 103 342 104 
<< m1 >>
rect 10 104 11 105 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< m1 >>
rect 19 104 20 105 
<< m2 >>
rect 19 104 20 105 
<< m1 >>
rect 21 104 22 105 
<< m1 >>
rect 23 104 24 105 
<< m1 >>
rect 28 104 29 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< m1 >>
rect 37 104 38 105 
<< m1 >>
rect 44 104 45 105 
<< m1 >>
rect 46 104 47 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m1 >>
rect 55 104 56 105 
<< m2 >>
rect 56 104 57 105 
<< m1 >>
rect 59 104 60 105 
<< m2 >>
rect 61 104 62 105 
<< m1 >>
rect 62 104 63 105 
<< m1 >>
rect 64 104 65 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< m1 >>
rect 73 104 74 105 
<< m2 >>
rect 73 104 74 105 
<< m1 >>
rect 78 104 79 105 
<< m2 >>
rect 81 104 82 105 
<< m1 >>
rect 82 104 83 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< m1 >>
rect 91 104 92 105 
<< m2 >>
rect 92 104 93 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< m1 >>
rect 109 104 110 105 
<< m2 >>
rect 109 104 110 105 
<< m1 >>
rect 115 104 116 105 
<< pdiffusion >>
rect 120 104 121 105 
<< pdiffusion >>
rect 121 104 122 105 
<< pdiffusion >>
rect 122 104 123 105 
<< pdiffusion >>
rect 123 104 124 105 
<< pdiffusion >>
rect 124 104 125 105 
<< pdiffusion >>
rect 125 104 126 105 
<< m1 >>
rect 130 104 131 105 
<< m1 >>
rect 132 104 133 105 
<< m1 >>
rect 136 104 137 105 
<< m2 >>
rect 136 104 137 105 
<< pdiffusion >>
rect 138 104 139 105 
<< pdiffusion >>
rect 139 104 140 105 
<< pdiffusion >>
rect 140 104 141 105 
<< pdiffusion >>
rect 141 104 142 105 
<< pdiffusion >>
rect 142 104 143 105 
<< pdiffusion >>
rect 143 104 144 105 
<< m1 >>
rect 145 104 146 105 
<< m2 >>
rect 145 104 146 105 
<< m1 >>
rect 147 104 148 105 
<< pdiffusion >>
rect 156 104 157 105 
<< pdiffusion >>
rect 157 104 158 105 
<< pdiffusion >>
rect 158 104 159 105 
<< pdiffusion >>
rect 159 104 160 105 
<< pdiffusion >>
rect 160 104 161 105 
<< pdiffusion >>
rect 161 104 162 105 
<< m1 >>
rect 163 104 164 105 
<< m1 >>
rect 167 104 168 105 
<< m2 >>
rect 167 104 168 105 
<< m2 >>
rect 168 104 169 105 
<< m2 >>
rect 169 104 170 105 
<< m1 >>
rect 170 104 171 105 
<< m1 >>
rect 172 104 173 105 
<< pdiffusion >>
rect 174 104 175 105 
<< pdiffusion >>
rect 175 104 176 105 
<< pdiffusion >>
rect 176 104 177 105 
<< pdiffusion >>
rect 177 104 178 105 
<< pdiffusion >>
rect 178 104 179 105 
<< pdiffusion >>
rect 179 104 180 105 
<< m1 >>
rect 190 104 191 105 
<< pdiffusion >>
rect 192 104 193 105 
<< pdiffusion >>
rect 193 104 194 105 
<< pdiffusion >>
rect 194 104 195 105 
<< pdiffusion >>
rect 195 104 196 105 
<< pdiffusion >>
rect 196 104 197 105 
<< pdiffusion >>
rect 197 104 198 105 
<< m1 >>
rect 199 104 200 105 
<< m1 >>
rect 201 104 202 105 
<< m2 >>
rect 202 104 203 105 
<< m1 >>
rect 205 104 206 105 
<< pdiffusion >>
rect 210 104 211 105 
<< pdiffusion >>
rect 211 104 212 105 
<< pdiffusion >>
rect 212 104 213 105 
<< pdiffusion >>
rect 213 104 214 105 
<< pdiffusion >>
rect 214 104 215 105 
<< pdiffusion >>
rect 215 104 216 105 
<< m1 >>
rect 218 104 219 105 
<< m1 >>
rect 226 104 227 105 
<< m2 >>
rect 226 104 227 105 
<< pdiffusion >>
rect 228 104 229 105 
<< pdiffusion >>
rect 229 104 230 105 
<< pdiffusion >>
rect 230 104 231 105 
<< pdiffusion >>
rect 231 104 232 105 
<< pdiffusion >>
rect 232 104 233 105 
<< pdiffusion >>
rect 233 104 234 105 
<< m1 >>
rect 235 104 236 105 
<< m2 >>
rect 236 104 237 105 
<< pdiffusion >>
rect 246 104 247 105 
<< pdiffusion >>
rect 247 104 248 105 
<< pdiffusion >>
rect 248 104 249 105 
<< pdiffusion >>
rect 249 104 250 105 
<< pdiffusion >>
rect 250 104 251 105 
<< pdiffusion >>
rect 251 104 252 105 
<< m1 >>
rect 254 104 255 105 
<< m2 >>
rect 255 104 256 105 
<< m1 >>
rect 258 104 259 105 
<< m1 >>
rect 260 104 261 105 
<< m1 >>
rect 262 104 263 105 
<< pdiffusion >>
rect 264 104 265 105 
<< pdiffusion >>
rect 265 104 266 105 
<< pdiffusion >>
rect 266 104 267 105 
<< pdiffusion >>
rect 267 104 268 105 
<< pdiffusion >>
rect 268 104 269 105 
<< pdiffusion >>
rect 269 104 270 105 
<< m1 >>
rect 271 104 272 105 
<< m1 >>
rect 274 104 275 105 
<< m1 >>
rect 276 104 277 105 
<< m1 >>
rect 278 104 279 105 
<< m2 >>
rect 279 104 280 105 
<< pdiffusion >>
rect 282 104 283 105 
<< pdiffusion >>
rect 283 104 284 105 
<< pdiffusion >>
rect 284 104 285 105 
<< pdiffusion >>
rect 285 104 286 105 
<< pdiffusion >>
rect 286 104 287 105 
<< pdiffusion >>
rect 287 104 288 105 
<< m1 >>
rect 296 104 297 105 
<< pdiffusion >>
rect 300 104 301 105 
<< pdiffusion >>
rect 301 104 302 105 
<< pdiffusion >>
rect 302 104 303 105 
<< pdiffusion >>
rect 303 104 304 105 
<< pdiffusion >>
rect 304 104 305 105 
<< pdiffusion >>
rect 305 104 306 105 
<< m1 >>
rect 307 104 308 105 
<< m2 >>
rect 308 104 309 105 
<< m2 >>
rect 315 104 316 105 
<< m1 >>
rect 316 104 317 105 
<< pdiffusion >>
rect 318 104 319 105 
<< pdiffusion >>
rect 319 104 320 105 
<< pdiffusion >>
rect 320 104 321 105 
<< pdiffusion >>
rect 321 104 322 105 
<< pdiffusion >>
rect 322 104 323 105 
<< pdiffusion >>
rect 323 104 324 105 
<< m1 >>
rect 327 104 328 105 
<< m1 >>
rect 329 104 330 105 
<< pdiffusion >>
rect 336 104 337 105 
<< pdiffusion >>
rect 337 104 338 105 
<< pdiffusion >>
rect 338 104 339 105 
<< pdiffusion >>
rect 339 104 340 105 
<< pdiffusion >>
rect 340 104 341 105 
<< pdiffusion >>
rect 341 104 342 105 
<< m1 >>
rect 10 105 11 106 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< m1 >>
rect 19 105 20 106 
<< m2 >>
rect 19 105 20 106 
<< m1 >>
rect 21 105 22 106 
<< m1 >>
rect 23 105 24 106 
<< m1 >>
rect 28 105 29 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< m1 >>
rect 37 105 38 106 
<< m1 >>
rect 44 105 45 106 
<< m1 >>
rect 46 105 47 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m1 >>
rect 55 105 56 106 
<< m2 >>
rect 56 105 57 106 
<< m1 >>
rect 59 105 60 106 
<< m2 >>
rect 61 105 62 106 
<< m1 >>
rect 62 105 63 106 
<< m1 >>
rect 64 105 65 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< m1 >>
rect 73 105 74 106 
<< m2 >>
rect 73 105 74 106 
<< m1 >>
rect 78 105 79 106 
<< m2 >>
rect 81 105 82 106 
<< m1 >>
rect 82 105 83 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< m1 >>
rect 91 105 92 106 
<< m2 >>
rect 92 105 93 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< m1 >>
rect 109 105 110 106 
<< m2 >>
rect 109 105 110 106 
<< m1 >>
rect 115 105 116 106 
<< pdiffusion >>
rect 120 105 121 106 
<< pdiffusion >>
rect 121 105 122 106 
<< pdiffusion >>
rect 122 105 123 106 
<< pdiffusion >>
rect 123 105 124 106 
<< pdiffusion >>
rect 124 105 125 106 
<< pdiffusion >>
rect 125 105 126 106 
<< m1 >>
rect 130 105 131 106 
<< m1 >>
rect 132 105 133 106 
<< m1 >>
rect 136 105 137 106 
<< m2 >>
rect 136 105 137 106 
<< pdiffusion >>
rect 138 105 139 106 
<< pdiffusion >>
rect 139 105 140 106 
<< pdiffusion >>
rect 140 105 141 106 
<< pdiffusion >>
rect 141 105 142 106 
<< pdiffusion >>
rect 142 105 143 106 
<< pdiffusion >>
rect 143 105 144 106 
<< m1 >>
rect 145 105 146 106 
<< m2 >>
rect 145 105 146 106 
<< m1 >>
rect 147 105 148 106 
<< pdiffusion >>
rect 156 105 157 106 
<< pdiffusion >>
rect 157 105 158 106 
<< pdiffusion >>
rect 158 105 159 106 
<< pdiffusion >>
rect 159 105 160 106 
<< pdiffusion >>
rect 160 105 161 106 
<< pdiffusion >>
rect 161 105 162 106 
<< m1 >>
rect 163 105 164 106 
<< m1 >>
rect 167 105 168 106 
<< m2 >>
rect 169 105 170 106 
<< m1 >>
rect 170 105 171 106 
<< m1 >>
rect 172 105 173 106 
<< pdiffusion >>
rect 174 105 175 106 
<< pdiffusion >>
rect 175 105 176 106 
<< pdiffusion >>
rect 176 105 177 106 
<< pdiffusion >>
rect 177 105 178 106 
<< pdiffusion >>
rect 178 105 179 106 
<< pdiffusion >>
rect 179 105 180 106 
<< m1 >>
rect 190 105 191 106 
<< pdiffusion >>
rect 192 105 193 106 
<< pdiffusion >>
rect 193 105 194 106 
<< pdiffusion >>
rect 194 105 195 106 
<< pdiffusion >>
rect 195 105 196 106 
<< pdiffusion >>
rect 196 105 197 106 
<< pdiffusion >>
rect 197 105 198 106 
<< m1 >>
rect 199 105 200 106 
<< m1 >>
rect 201 105 202 106 
<< m2 >>
rect 202 105 203 106 
<< m1 >>
rect 205 105 206 106 
<< pdiffusion >>
rect 210 105 211 106 
<< pdiffusion >>
rect 211 105 212 106 
<< pdiffusion >>
rect 212 105 213 106 
<< pdiffusion >>
rect 213 105 214 106 
<< pdiffusion >>
rect 214 105 215 106 
<< pdiffusion >>
rect 215 105 216 106 
<< m1 >>
rect 218 105 219 106 
<< m1 >>
rect 226 105 227 106 
<< m2 >>
rect 226 105 227 106 
<< pdiffusion >>
rect 228 105 229 106 
<< pdiffusion >>
rect 229 105 230 106 
<< pdiffusion >>
rect 230 105 231 106 
<< pdiffusion >>
rect 231 105 232 106 
<< pdiffusion >>
rect 232 105 233 106 
<< pdiffusion >>
rect 233 105 234 106 
<< m1 >>
rect 235 105 236 106 
<< m2 >>
rect 236 105 237 106 
<< m1 >>
rect 237 105 238 106 
<< m2 >>
rect 237 105 238 106 
<< m2c >>
rect 237 105 238 106 
<< m1 >>
rect 237 105 238 106 
<< m2 >>
rect 237 105 238 106 
<< m1 >>
rect 238 105 239 106 
<< m1 >>
rect 239 105 240 106 
<< m1 >>
rect 240 105 241 106 
<< m1 >>
rect 241 105 242 106 
<< m1 >>
rect 242 105 243 106 
<< m1 >>
rect 243 105 244 106 
<< m1 >>
rect 244 105 245 106 
<< pdiffusion >>
rect 246 105 247 106 
<< pdiffusion >>
rect 247 105 248 106 
<< pdiffusion >>
rect 248 105 249 106 
<< pdiffusion >>
rect 249 105 250 106 
<< pdiffusion >>
rect 250 105 251 106 
<< pdiffusion >>
rect 251 105 252 106 
<< m1 >>
rect 254 105 255 106 
<< m2 >>
rect 255 105 256 106 
<< m1 >>
rect 258 105 259 106 
<< m1 >>
rect 260 105 261 106 
<< m1 >>
rect 262 105 263 106 
<< pdiffusion >>
rect 264 105 265 106 
<< pdiffusion >>
rect 265 105 266 106 
<< pdiffusion >>
rect 266 105 267 106 
<< pdiffusion >>
rect 267 105 268 106 
<< pdiffusion >>
rect 268 105 269 106 
<< pdiffusion >>
rect 269 105 270 106 
<< m1 >>
rect 271 105 272 106 
<< m1 >>
rect 274 105 275 106 
<< m1 >>
rect 276 105 277 106 
<< m1 >>
rect 278 105 279 106 
<< m2 >>
rect 279 105 280 106 
<< pdiffusion >>
rect 282 105 283 106 
<< pdiffusion >>
rect 283 105 284 106 
<< pdiffusion >>
rect 284 105 285 106 
<< pdiffusion >>
rect 285 105 286 106 
<< pdiffusion >>
rect 286 105 287 106 
<< pdiffusion >>
rect 287 105 288 106 
<< m1 >>
rect 296 105 297 106 
<< pdiffusion >>
rect 300 105 301 106 
<< pdiffusion >>
rect 301 105 302 106 
<< pdiffusion >>
rect 302 105 303 106 
<< pdiffusion >>
rect 303 105 304 106 
<< pdiffusion >>
rect 304 105 305 106 
<< pdiffusion >>
rect 305 105 306 106 
<< m1 >>
rect 307 105 308 106 
<< m2 >>
rect 308 105 309 106 
<< m2 >>
rect 315 105 316 106 
<< m1 >>
rect 316 105 317 106 
<< pdiffusion >>
rect 318 105 319 106 
<< pdiffusion >>
rect 319 105 320 106 
<< pdiffusion >>
rect 320 105 321 106 
<< pdiffusion >>
rect 321 105 322 106 
<< pdiffusion >>
rect 322 105 323 106 
<< pdiffusion >>
rect 323 105 324 106 
<< m1 >>
rect 327 105 328 106 
<< m1 >>
rect 329 105 330 106 
<< pdiffusion >>
rect 336 105 337 106 
<< pdiffusion >>
rect 337 105 338 106 
<< pdiffusion >>
rect 338 105 339 106 
<< pdiffusion >>
rect 339 105 340 106 
<< pdiffusion >>
rect 340 105 341 106 
<< pdiffusion >>
rect 341 105 342 106 
<< m1 >>
rect 10 106 11 107 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< m1 >>
rect 19 106 20 107 
<< m2 >>
rect 19 106 20 107 
<< m1 >>
rect 21 106 22 107 
<< m1 >>
rect 23 106 24 107 
<< m1 >>
rect 28 106 29 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< m1 >>
rect 37 106 38 107 
<< m1 >>
rect 44 106 45 107 
<< m1 >>
rect 46 106 47 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m1 >>
rect 55 106 56 107 
<< m2 >>
rect 56 106 57 107 
<< m1 >>
rect 59 106 60 107 
<< m2 >>
rect 61 106 62 107 
<< m1 >>
rect 62 106 63 107 
<< m1 >>
rect 64 106 65 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< m1 >>
rect 73 106 74 107 
<< m2 >>
rect 73 106 74 107 
<< m1 >>
rect 78 106 79 107 
<< m2 >>
rect 81 106 82 107 
<< m1 >>
rect 82 106 83 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< m1 >>
rect 91 106 92 107 
<< m2 >>
rect 92 106 93 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< m1 >>
rect 109 106 110 107 
<< m2 >>
rect 109 106 110 107 
<< m1 >>
rect 115 106 116 107 
<< pdiffusion >>
rect 120 106 121 107 
<< pdiffusion >>
rect 121 106 122 107 
<< pdiffusion >>
rect 122 106 123 107 
<< pdiffusion >>
rect 123 106 124 107 
<< pdiffusion >>
rect 124 106 125 107 
<< pdiffusion >>
rect 125 106 126 107 
<< m1 >>
rect 130 106 131 107 
<< m1 >>
rect 132 106 133 107 
<< m1 >>
rect 136 106 137 107 
<< m2 >>
rect 136 106 137 107 
<< pdiffusion >>
rect 138 106 139 107 
<< pdiffusion >>
rect 139 106 140 107 
<< pdiffusion >>
rect 140 106 141 107 
<< pdiffusion >>
rect 141 106 142 107 
<< pdiffusion >>
rect 142 106 143 107 
<< pdiffusion >>
rect 143 106 144 107 
<< m1 >>
rect 145 106 146 107 
<< m2 >>
rect 145 106 146 107 
<< m1 >>
rect 147 106 148 107 
<< pdiffusion >>
rect 156 106 157 107 
<< pdiffusion >>
rect 157 106 158 107 
<< pdiffusion >>
rect 158 106 159 107 
<< pdiffusion >>
rect 159 106 160 107 
<< pdiffusion >>
rect 160 106 161 107 
<< pdiffusion >>
rect 161 106 162 107 
<< m1 >>
rect 163 106 164 107 
<< m1 >>
rect 167 106 168 107 
<< m2 >>
rect 169 106 170 107 
<< m1 >>
rect 170 106 171 107 
<< m1 >>
rect 172 106 173 107 
<< pdiffusion >>
rect 174 106 175 107 
<< pdiffusion >>
rect 175 106 176 107 
<< pdiffusion >>
rect 176 106 177 107 
<< pdiffusion >>
rect 177 106 178 107 
<< pdiffusion >>
rect 178 106 179 107 
<< pdiffusion >>
rect 179 106 180 107 
<< m1 >>
rect 190 106 191 107 
<< pdiffusion >>
rect 192 106 193 107 
<< pdiffusion >>
rect 193 106 194 107 
<< pdiffusion >>
rect 194 106 195 107 
<< pdiffusion >>
rect 195 106 196 107 
<< pdiffusion >>
rect 196 106 197 107 
<< pdiffusion >>
rect 197 106 198 107 
<< m1 >>
rect 199 106 200 107 
<< m1 >>
rect 201 106 202 107 
<< m2 >>
rect 202 106 203 107 
<< m1 >>
rect 205 106 206 107 
<< pdiffusion >>
rect 210 106 211 107 
<< pdiffusion >>
rect 211 106 212 107 
<< pdiffusion >>
rect 212 106 213 107 
<< pdiffusion >>
rect 213 106 214 107 
<< pdiffusion >>
rect 214 106 215 107 
<< pdiffusion >>
rect 215 106 216 107 
<< m1 >>
rect 218 106 219 107 
<< m1 >>
rect 226 106 227 107 
<< m2 >>
rect 226 106 227 107 
<< pdiffusion >>
rect 228 106 229 107 
<< pdiffusion >>
rect 229 106 230 107 
<< pdiffusion >>
rect 230 106 231 107 
<< pdiffusion >>
rect 231 106 232 107 
<< pdiffusion >>
rect 232 106 233 107 
<< pdiffusion >>
rect 233 106 234 107 
<< m1 >>
rect 235 106 236 107 
<< m1 >>
rect 244 106 245 107 
<< pdiffusion >>
rect 246 106 247 107 
<< pdiffusion >>
rect 247 106 248 107 
<< pdiffusion >>
rect 248 106 249 107 
<< pdiffusion >>
rect 249 106 250 107 
<< pdiffusion >>
rect 250 106 251 107 
<< pdiffusion >>
rect 251 106 252 107 
<< m1 >>
rect 254 106 255 107 
<< m2 >>
rect 255 106 256 107 
<< m1 >>
rect 258 106 259 107 
<< m1 >>
rect 260 106 261 107 
<< m1 >>
rect 262 106 263 107 
<< pdiffusion >>
rect 264 106 265 107 
<< pdiffusion >>
rect 265 106 266 107 
<< pdiffusion >>
rect 266 106 267 107 
<< pdiffusion >>
rect 267 106 268 107 
<< pdiffusion >>
rect 268 106 269 107 
<< pdiffusion >>
rect 269 106 270 107 
<< m1 >>
rect 271 106 272 107 
<< m1 >>
rect 274 106 275 107 
<< m1 >>
rect 276 106 277 107 
<< m1 >>
rect 278 106 279 107 
<< m2 >>
rect 279 106 280 107 
<< pdiffusion >>
rect 282 106 283 107 
<< pdiffusion >>
rect 283 106 284 107 
<< pdiffusion >>
rect 284 106 285 107 
<< pdiffusion >>
rect 285 106 286 107 
<< pdiffusion >>
rect 286 106 287 107 
<< pdiffusion >>
rect 287 106 288 107 
<< m1 >>
rect 296 106 297 107 
<< pdiffusion >>
rect 300 106 301 107 
<< pdiffusion >>
rect 301 106 302 107 
<< pdiffusion >>
rect 302 106 303 107 
<< pdiffusion >>
rect 303 106 304 107 
<< pdiffusion >>
rect 304 106 305 107 
<< pdiffusion >>
rect 305 106 306 107 
<< m1 >>
rect 307 106 308 107 
<< m2 >>
rect 308 106 309 107 
<< m2 >>
rect 315 106 316 107 
<< m1 >>
rect 316 106 317 107 
<< pdiffusion >>
rect 318 106 319 107 
<< pdiffusion >>
rect 319 106 320 107 
<< pdiffusion >>
rect 320 106 321 107 
<< pdiffusion >>
rect 321 106 322 107 
<< pdiffusion >>
rect 322 106 323 107 
<< pdiffusion >>
rect 323 106 324 107 
<< m1 >>
rect 327 106 328 107 
<< m1 >>
rect 329 106 330 107 
<< pdiffusion >>
rect 336 106 337 107 
<< pdiffusion >>
rect 337 106 338 107 
<< pdiffusion >>
rect 338 106 339 107 
<< pdiffusion >>
rect 339 106 340 107 
<< pdiffusion >>
rect 340 106 341 107 
<< pdiffusion >>
rect 341 106 342 107 
<< m1 >>
rect 10 107 11 108 
<< pdiffusion >>
rect 12 107 13 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< m1 >>
rect 19 107 20 108 
<< m2 >>
rect 19 107 20 108 
<< m1 >>
rect 21 107 22 108 
<< m1 >>
rect 23 107 24 108 
<< m1 >>
rect 28 107 29 108 
<< pdiffusion >>
rect 30 107 31 108 
<< m1 >>
rect 31 107 32 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< m1 >>
rect 37 107 38 108 
<< m1 >>
rect 44 107 45 108 
<< m1 >>
rect 46 107 47 108 
<< pdiffusion >>
rect 48 107 49 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< m1 >>
rect 52 107 53 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m1 >>
rect 55 107 56 108 
<< m2 >>
rect 56 107 57 108 
<< m1 >>
rect 59 107 60 108 
<< m2 >>
rect 61 107 62 108 
<< m1 >>
rect 62 107 63 108 
<< m1 >>
rect 64 107 65 108 
<< pdiffusion >>
rect 66 107 67 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< m1 >>
rect 70 107 71 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< m1 >>
rect 73 107 74 108 
<< m2 >>
rect 73 107 74 108 
<< m1 >>
rect 78 107 79 108 
<< m2 >>
rect 81 107 82 108 
<< m1 >>
rect 82 107 83 108 
<< pdiffusion >>
rect 84 107 85 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< m1 >>
rect 91 107 92 108 
<< m2 >>
rect 92 107 93 108 
<< pdiffusion >>
rect 102 107 103 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< m1 >>
rect 109 107 110 108 
<< m2 >>
rect 109 107 110 108 
<< m1 >>
rect 115 107 116 108 
<< pdiffusion >>
rect 120 107 121 108 
<< pdiffusion >>
rect 121 107 122 108 
<< pdiffusion >>
rect 122 107 123 108 
<< pdiffusion >>
rect 123 107 124 108 
<< pdiffusion >>
rect 124 107 125 108 
<< pdiffusion >>
rect 125 107 126 108 
<< m1 >>
rect 130 107 131 108 
<< m1 >>
rect 132 107 133 108 
<< m1 >>
rect 136 107 137 108 
<< m2 >>
rect 136 107 137 108 
<< pdiffusion >>
rect 138 107 139 108 
<< pdiffusion >>
rect 139 107 140 108 
<< pdiffusion >>
rect 140 107 141 108 
<< pdiffusion >>
rect 141 107 142 108 
<< pdiffusion >>
rect 142 107 143 108 
<< pdiffusion >>
rect 143 107 144 108 
<< m1 >>
rect 145 107 146 108 
<< m2 >>
rect 145 107 146 108 
<< m1 >>
rect 147 107 148 108 
<< pdiffusion >>
rect 156 107 157 108 
<< pdiffusion >>
rect 157 107 158 108 
<< pdiffusion >>
rect 158 107 159 108 
<< pdiffusion >>
rect 159 107 160 108 
<< pdiffusion >>
rect 160 107 161 108 
<< pdiffusion >>
rect 161 107 162 108 
<< m1 >>
rect 163 107 164 108 
<< m1 >>
rect 167 107 168 108 
<< m2 >>
rect 169 107 170 108 
<< m1 >>
rect 170 107 171 108 
<< m1 >>
rect 172 107 173 108 
<< pdiffusion >>
rect 174 107 175 108 
<< pdiffusion >>
rect 175 107 176 108 
<< pdiffusion >>
rect 176 107 177 108 
<< pdiffusion >>
rect 177 107 178 108 
<< pdiffusion >>
rect 178 107 179 108 
<< pdiffusion >>
rect 179 107 180 108 
<< m1 >>
rect 190 107 191 108 
<< pdiffusion >>
rect 192 107 193 108 
<< pdiffusion >>
rect 193 107 194 108 
<< pdiffusion >>
rect 194 107 195 108 
<< pdiffusion >>
rect 195 107 196 108 
<< pdiffusion >>
rect 196 107 197 108 
<< pdiffusion >>
rect 197 107 198 108 
<< m1 >>
rect 199 107 200 108 
<< m1 >>
rect 201 107 202 108 
<< m2 >>
rect 202 107 203 108 
<< m1 >>
rect 205 107 206 108 
<< pdiffusion >>
rect 210 107 211 108 
<< pdiffusion >>
rect 211 107 212 108 
<< pdiffusion >>
rect 212 107 213 108 
<< pdiffusion >>
rect 213 107 214 108 
<< m1 >>
rect 214 107 215 108 
<< pdiffusion >>
rect 214 107 215 108 
<< pdiffusion >>
rect 215 107 216 108 
<< m1 >>
rect 218 107 219 108 
<< m1 >>
rect 226 107 227 108 
<< m2 >>
rect 226 107 227 108 
<< pdiffusion >>
rect 228 107 229 108 
<< pdiffusion >>
rect 229 107 230 108 
<< pdiffusion >>
rect 230 107 231 108 
<< pdiffusion >>
rect 231 107 232 108 
<< m1 >>
rect 232 107 233 108 
<< pdiffusion >>
rect 232 107 233 108 
<< pdiffusion >>
rect 233 107 234 108 
<< m1 >>
rect 235 107 236 108 
<< m2 >>
rect 235 107 236 108 
<< m2c >>
rect 235 107 236 108 
<< m1 >>
rect 235 107 236 108 
<< m2 >>
rect 235 107 236 108 
<< m1 >>
rect 244 107 245 108 
<< pdiffusion >>
rect 246 107 247 108 
<< pdiffusion >>
rect 247 107 248 108 
<< pdiffusion >>
rect 248 107 249 108 
<< pdiffusion >>
rect 249 107 250 108 
<< m1 >>
rect 250 107 251 108 
<< pdiffusion >>
rect 250 107 251 108 
<< pdiffusion >>
rect 251 107 252 108 
<< m1 >>
rect 254 107 255 108 
<< m2 >>
rect 255 107 256 108 
<< m1 >>
rect 258 107 259 108 
<< m1 >>
rect 260 107 261 108 
<< m1 >>
rect 262 107 263 108 
<< pdiffusion >>
rect 264 107 265 108 
<< pdiffusion >>
rect 265 107 266 108 
<< pdiffusion >>
rect 266 107 267 108 
<< pdiffusion >>
rect 267 107 268 108 
<< pdiffusion >>
rect 268 107 269 108 
<< pdiffusion >>
rect 269 107 270 108 
<< m1 >>
rect 271 107 272 108 
<< m1 >>
rect 274 107 275 108 
<< m1 >>
rect 276 107 277 108 
<< m1 >>
rect 278 107 279 108 
<< m2 >>
rect 279 107 280 108 
<< pdiffusion >>
rect 282 107 283 108 
<< pdiffusion >>
rect 283 107 284 108 
<< pdiffusion >>
rect 284 107 285 108 
<< pdiffusion >>
rect 285 107 286 108 
<< pdiffusion >>
rect 286 107 287 108 
<< pdiffusion >>
rect 287 107 288 108 
<< m1 >>
rect 296 107 297 108 
<< pdiffusion >>
rect 300 107 301 108 
<< pdiffusion >>
rect 301 107 302 108 
<< pdiffusion >>
rect 302 107 303 108 
<< pdiffusion >>
rect 303 107 304 108 
<< pdiffusion >>
rect 304 107 305 108 
<< pdiffusion >>
rect 305 107 306 108 
<< m1 >>
rect 307 107 308 108 
<< m2 >>
rect 308 107 309 108 
<< m2 >>
rect 315 107 316 108 
<< m1 >>
rect 316 107 317 108 
<< pdiffusion >>
rect 318 107 319 108 
<< pdiffusion >>
rect 319 107 320 108 
<< pdiffusion >>
rect 320 107 321 108 
<< pdiffusion >>
rect 321 107 322 108 
<< pdiffusion >>
rect 322 107 323 108 
<< pdiffusion >>
rect 323 107 324 108 
<< m1 >>
rect 327 107 328 108 
<< m1 >>
rect 329 107 330 108 
<< pdiffusion >>
rect 336 107 337 108 
<< pdiffusion >>
rect 337 107 338 108 
<< pdiffusion >>
rect 338 107 339 108 
<< pdiffusion >>
rect 339 107 340 108 
<< pdiffusion >>
rect 340 107 341 108 
<< pdiffusion >>
rect 341 107 342 108 
<< m1 >>
rect 10 108 11 109 
<< m1 >>
rect 19 108 20 109 
<< m2 >>
rect 19 108 20 109 
<< m1 >>
rect 21 108 22 109 
<< m1 >>
rect 23 108 24 109 
<< m1 >>
rect 28 108 29 109 
<< m1 >>
rect 31 108 32 109 
<< m1 >>
rect 37 108 38 109 
<< m1 >>
rect 44 108 45 109 
<< m1 >>
rect 46 108 47 109 
<< m1 >>
rect 52 108 53 109 
<< m1 >>
rect 55 108 56 109 
<< m2 >>
rect 56 108 57 109 
<< m1 >>
rect 59 108 60 109 
<< m2 >>
rect 61 108 62 109 
<< m1 >>
rect 62 108 63 109 
<< m1 >>
rect 64 108 65 109 
<< m1 >>
rect 70 108 71 109 
<< m1 >>
rect 73 108 74 109 
<< m2 >>
rect 73 108 74 109 
<< m1 >>
rect 78 108 79 109 
<< m2 >>
rect 81 108 82 109 
<< m1 >>
rect 82 108 83 109 
<< m1 >>
rect 91 108 92 109 
<< m2 >>
rect 92 108 93 109 
<< m1 >>
rect 109 108 110 109 
<< m2 >>
rect 109 108 110 109 
<< m1 >>
rect 115 108 116 109 
<< m1 >>
rect 130 108 131 109 
<< m1 >>
rect 132 108 133 109 
<< m1 >>
rect 136 108 137 109 
<< m2 >>
rect 136 108 137 109 
<< m1 >>
rect 145 108 146 109 
<< m2 >>
rect 145 108 146 109 
<< m1 >>
rect 147 108 148 109 
<< m1 >>
rect 163 108 164 109 
<< m1 >>
rect 167 108 168 109 
<< m2 >>
rect 169 108 170 109 
<< m1 >>
rect 170 108 171 109 
<< m1 >>
rect 172 108 173 109 
<< m1 >>
rect 190 108 191 109 
<< m1 >>
rect 199 108 200 109 
<< m1 >>
rect 201 108 202 109 
<< m2 >>
rect 202 108 203 109 
<< m1 >>
rect 205 108 206 109 
<< m1 >>
rect 214 108 215 109 
<< m1 >>
rect 218 108 219 109 
<< m1 >>
rect 226 108 227 109 
<< m2 >>
rect 226 108 227 109 
<< m1 >>
rect 232 108 233 109 
<< m2 >>
rect 235 108 236 109 
<< m1 >>
rect 244 108 245 109 
<< m1 >>
rect 250 108 251 109 
<< m1 >>
rect 254 108 255 109 
<< m2 >>
rect 255 108 256 109 
<< m1 >>
rect 258 108 259 109 
<< m1 >>
rect 260 108 261 109 
<< m1 >>
rect 262 108 263 109 
<< m1 >>
rect 271 108 272 109 
<< m1 >>
rect 274 108 275 109 
<< m1 >>
rect 276 108 277 109 
<< m1 >>
rect 278 108 279 109 
<< m2 >>
rect 279 108 280 109 
<< m1 >>
rect 296 108 297 109 
<< m1 >>
rect 307 108 308 109 
<< m2 >>
rect 308 108 309 109 
<< m2 >>
rect 315 108 316 109 
<< m1 >>
rect 316 108 317 109 
<< m1 >>
rect 327 108 328 109 
<< m1 >>
rect 329 108 330 109 
<< m1 >>
rect 10 109 11 110 
<< m1 >>
rect 19 109 20 110 
<< m2 >>
rect 19 109 20 110 
<< m1 >>
rect 21 109 22 110 
<< m1 >>
rect 23 109 24 110 
<< m1 >>
rect 28 109 29 110 
<< m1 >>
rect 31 109 32 110 
<< m1 >>
rect 37 109 38 110 
<< m1 >>
rect 44 109 45 110 
<< m1 >>
rect 46 109 47 110 
<< m1 >>
rect 52 109 53 110 
<< m1 >>
rect 55 109 56 110 
<< m2 >>
rect 56 109 57 110 
<< m1 >>
rect 59 109 60 110 
<< m2 >>
rect 61 109 62 110 
<< m1 >>
rect 62 109 63 110 
<< m1 >>
rect 64 109 65 110 
<< m1 >>
rect 70 109 71 110 
<< m1 >>
rect 71 109 72 110 
<< m2 >>
rect 71 109 72 110 
<< m2c >>
rect 71 109 72 110 
<< m1 >>
rect 71 109 72 110 
<< m2 >>
rect 71 109 72 110 
<< m2 >>
rect 72 109 73 110 
<< m1 >>
rect 73 109 74 110 
<< m2 >>
rect 73 109 74 110 
<< m1 >>
rect 78 109 79 110 
<< m2 >>
rect 81 109 82 110 
<< m1 >>
rect 82 109 83 110 
<< m1 >>
rect 91 109 92 110 
<< m2 >>
rect 92 109 93 110 
<< m1 >>
rect 109 109 110 110 
<< m2 >>
rect 109 109 110 110 
<< m1 >>
rect 115 109 116 110 
<< m1 >>
rect 130 109 131 110 
<< m1 >>
rect 132 109 133 110 
<< m1 >>
rect 136 109 137 110 
<< m2 >>
rect 136 109 137 110 
<< m1 >>
rect 145 109 146 110 
<< m2 >>
rect 145 109 146 110 
<< m1 >>
rect 147 109 148 110 
<< m1 >>
rect 163 109 164 110 
<< m1 >>
rect 167 109 168 110 
<< m2 >>
rect 169 109 170 110 
<< m1 >>
rect 170 109 171 110 
<< m1 >>
rect 172 109 173 110 
<< m1 >>
rect 190 109 191 110 
<< m1 >>
rect 199 109 200 110 
<< m1 >>
rect 201 109 202 110 
<< m2 >>
rect 202 109 203 110 
<< m1 >>
rect 205 109 206 110 
<< m1 >>
rect 214 109 215 110 
<< m1 >>
rect 215 109 216 110 
<< m1 >>
rect 216 109 217 110 
<< m1 >>
rect 217 109 218 110 
<< m1 >>
rect 218 109 219 110 
<< m1 >>
rect 226 109 227 110 
<< m2 >>
rect 226 109 227 110 
<< m1 >>
rect 232 109 233 110 
<< m1 >>
rect 233 109 234 110 
<< m1 >>
rect 234 109 235 110 
<< m1 >>
rect 235 109 236 110 
<< m2 >>
rect 235 109 236 110 
<< m1 >>
rect 244 109 245 110 
<< m1 >>
rect 250 109 251 110 
<< m1 >>
rect 251 109 252 110 
<< m1 >>
rect 252 109 253 110 
<< m1 >>
rect 253 109 254 110 
<< m1 >>
rect 254 109 255 110 
<< m2 >>
rect 255 109 256 110 
<< m1 >>
rect 258 109 259 110 
<< m1 >>
rect 260 109 261 110 
<< m1 >>
rect 262 109 263 110 
<< m1 >>
rect 269 109 270 110 
<< m2 >>
rect 269 109 270 110 
<< m2c >>
rect 269 109 270 110 
<< m1 >>
rect 269 109 270 110 
<< m2 >>
rect 269 109 270 110 
<< m2 >>
rect 270 109 271 110 
<< m1 >>
rect 271 109 272 110 
<< m2 >>
rect 271 109 272 110 
<< m2 >>
rect 272 109 273 110 
<< m2 >>
rect 273 109 274 110 
<< m1 >>
rect 274 109 275 110 
<< m2 >>
rect 274 109 275 110 
<< m2 >>
rect 275 109 276 110 
<< m1 >>
rect 276 109 277 110 
<< m2 >>
rect 276 109 277 110 
<< m2 >>
rect 277 109 278 110 
<< m1 >>
rect 278 109 279 110 
<< m2 >>
rect 278 109 279 110 
<< m2 >>
rect 279 109 280 110 
<< m1 >>
rect 296 109 297 110 
<< m1 >>
rect 307 109 308 110 
<< m2 >>
rect 308 109 309 110 
<< m2 >>
rect 315 109 316 110 
<< m1 >>
rect 316 109 317 110 
<< m2 >>
rect 316 109 317 110 
<< m2 >>
rect 317 109 318 110 
<< m1 >>
rect 318 109 319 110 
<< m2 >>
rect 318 109 319 110 
<< m2c >>
rect 318 109 319 110 
<< m1 >>
rect 318 109 319 110 
<< m2 >>
rect 318 109 319 110 
<< m1 >>
rect 327 109 328 110 
<< m1 >>
rect 329 109 330 110 
<< m1 >>
rect 10 110 11 111 
<< m1 >>
rect 19 110 20 111 
<< m2 >>
rect 19 110 20 111 
<< m1 >>
rect 21 110 22 111 
<< m1 >>
rect 23 110 24 111 
<< m2 >>
rect 27 110 28 111 
<< m1 >>
rect 28 110 29 111 
<< m2 >>
rect 28 110 29 111 
<< m2 >>
rect 29 110 30 111 
<< m1 >>
rect 30 110 31 111 
<< m2 >>
rect 30 110 31 111 
<< m2c >>
rect 30 110 31 111 
<< m1 >>
rect 30 110 31 111 
<< m2 >>
rect 30 110 31 111 
<< m1 >>
rect 31 110 32 111 
<< m1 >>
rect 37 110 38 111 
<< m2 >>
rect 37 110 38 111 
<< m2c >>
rect 37 110 38 111 
<< m1 >>
rect 37 110 38 111 
<< m2 >>
rect 37 110 38 111 
<< m1 >>
rect 44 110 45 111 
<< m1 >>
rect 46 110 47 111 
<< m1 >>
rect 50 110 51 111 
<< m2 >>
rect 50 110 51 111 
<< m2c >>
rect 50 110 51 111 
<< m1 >>
rect 50 110 51 111 
<< m2 >>
rect 50 110 51 111 
<< m2 >>
rect 51 110 52 111 
<< m1 >>
rect 52 110 53 111 
<< m2 >>
rect 52 110 53 111 
<< m2 >>
rect 53 110 54 111 
<< m2 >>
rect 54 110 55 111 
<< m1 >>
rect 55 110 56 111 
<< m2 >>
rect 55 110 56 111 
<< m2 >>
rect 56 110 57 111 
<< m1 >>
rect 59 110 60 111 
<< m2 >>
rect 61 110 62 111 
<< m1 >>
rect 62 110 63 111 
<< m1 >>
rect 64 110 65 111 
<< m1 >>
rect 73 110 74 111 
<< m1 >>
rect 78 110 79 111 
<< m2 >>
rect 81 110 82 111 
<< m1 >>
rect 82 110 83 111 
<< m1 >>
rect 91 110 92 111 
<< m2 >>
rect 92 110 93 111 
<< m1 >>
rect 109 110 110 111 
<< m2 >>
rect 109 110 110 111 
<< m1 >>
rect 115 110 116 111 
<< m1 >>
rect 130 110 131 111 
<< m1 >>
rect 132 110 133 111 
<< m1 >>
rect 136 110 137 111 
<< m2 >>
rect 136 110 137 111 
<< m1 >>
rect 145 110 146 111 
<< m2 >>
rect 145 110 146 111 
<< m1 >>
rect 147 110 148 111 
<< m1 >>
rect 163 110 164 111 
<< m1 >>
rect 167 110 168 111 
<< m2 >>
rect 169 110 170 111 
<< m1 >>
rect 170 110 171 111 
<< m1 >>
rect 172 110 173 111 
<< m1 >>
rect 190 110 191 111 
<< m1 >>
rect 199 110 200 111 
<< m1 >>
rect 201 110 202 111 
<< m2 >>
rect 202 110 203 111 
<< m1 >>
rect 205 110 206 111 
<< m1 >>
rect 226 110 227 111 
<< m2 >>
rect 226 110 227 111 
<< m1 >>
rect 235 110 236 111 
<< m2 >>
rect 235 110 236 111 
<< m1 >>
rect 244 110 245 111 
<< m2 >>
rect 255 110 256 111 
<< m1 >>
rect 256 110 257 111 
<< m2 >>
rect 256 110 257 111 
<< m2c >>
rect 256 110 257 111 
<< m1 >>
rect 256 110 257 111 
<< m2 >>
rect 256 110 257 111 
<< m1 >>
rect 258 110 259 111 
<< m1 >>
rect 260 110 261 111 
<< m1 >>
rect 262 110 263 111 
<< m1 >>
rect 269 110 270 111 
<< m1 >>
rect 271 110 272 111 
<< m1 >>
rect 274 110 275 111 
<< m1 >>
rect 276 110 277 111 
<< m1 >>
rect 278 110 279 111 
<< m1 >>
rect 296 110 297 111 
<< m1 >>
rect 307 110 308 111 
<< m2 >>
rect 308 110 309 111 
<< m1 >>
rect 316 110 317 111 
<< m1 >>
rect 318 110 319 111 
<< m1 >>
rect 327 110 328 111 
<< m1 >>
rect 329 110 330 111 
<< m1 >>
rect 10 111 11 112 
<< m1 >>
rect 19 111 20 112 
<< m2 >>
rect 19 111 20 112 
<< m1 >>
rect 21 111 22 112 
<< m1 >>
rect 23 111 24 112 
<< m2 >>
rect 27 111 28 112 
<< m1 >>
rect 28 111 29 112 
<< m2 >>
rect 37 111 38 112 
<< m1 >>
rect 44 111 45 112 
<< m1 >>
rect 46 111 47 112 
<< m1 >>
rect 50 111 51 112 
<< m1 >>
rect 52 111 53 112 
<< m1 >>
rect 55 111 56 112 
<< m1 >>
rect 59 111 60 112 
<< m2 >>
rect 61 111 62 112 
<< m1 >>
rect 62 111 63 112 
<< m1 >>
rect 64 111 65 112 
<< m1 >>
rect 73 111 74 112 
<< m1 >>
rect 78 111 79 112 
<< m2 >>
rect 81 111 82 112 
<< m1 >>
rect 82 111 83 112 
<< m1 >>
rect 91 111 92 112 
<< m2 >>
rect 92 111 93 112 
<< m1 >>
rect 109 111 110 112 
<< m2 >>
rect 109 111 110 112 
<< m1 >>
rect 115 111 116 112 
<< m1 >>
rect 130 111 131 112 
<< m1 >>
rect 132 111 133 112 
<< m1 >>
rect 136 111 137 112 
<< m2 >>
rect 136 111 137 112 
<< m1 >>
rect 145 111 146 112 
<< m2 >>
rect 145 111 146 112 
<< m1 >>
rect 147 111 148 112 
<< m1 >>
rect 163 111 164 112 
<< m1 >>
rect 167 111 168 112 
<< m2 >>
rect 169 111 170 112 
<< m1 >>
rect 170 111 171 112 
<< m1 >>
rect 172 111 173 112 
<< m1 >>
rect 190 111 191 112 
<< m1 >>
rect 199 111 200 112 
<< m1 >>
rect 201 111 202 112 
<< m2 >>
rect 202 111 203 112 
<< m1 >>
rect 205 111 206 112 
<< m1 >>
rect 226 111 227 112 
<< m2 >>
rect 226 111 227 112 
<< m1 >>
rect 235 111 236 112 
<< m2 >>
rect 235 111 236 112 
<< m1 >>
rect 244 111 245 112 
<< m1 >>
rect 256 111 257 112 
<< m1 >>
rect 258 111 259 112 
<< m1 >>
rect 260 111 261 112 
<< m1 >>
rect 262 111 263 112 
<< m1 >>
rect 269 111 270 112 
<< m1 >>
rect 271 111 272 112 
<< m1 >>
rect 274 111 275 112 
<< m1 >>
rect 276 111 277 112 
<< m1 >>
rect 278 111 279 112 
<< m1 >>
rect 296 111 297 112 
<< m1 >>
rect 307 111 308 112 
<< m2 >>
rect 308 111 309 112 
<< m1 >>
rect 316 111 317 112 
<< m1 >>
rect 318 111 319 112 
<< m1 >>
rect 327 111 328 112 
<< m1 >>
rect 329 111 330 112 
<< m1 >>
rect 10 112 11 113 
<< m1 >>
rect 19 112 20 113 
<< m2 >>
rect 19 112 20 113 
<< m1 >>
rect 21 112 22 113 
<< m1 >>
rect 23 112 24 113 
<< m2 >>
rect 27 112 28 113 
<< m1 >>
rect 28 112 29 113 
<< m1 >>
rect 31 112 32 113 
<< m1 >>
rect 32 112 33 113 
<< m1 >>
rect 33 112 34 113 
<< m1 >>
rect 34 112 35 113 
<< m1 >>
rect 35 112 36 113 
<< m1 >>
rect 36 112 37 113 
<< m1 >>
rect 37 112 38 113 
<< m2 >>
rect 37 112 38 113 
<< m1 >>
rect 38 112 39 113 
<< m1 >>
rect 39 112 40 113 
<< m1 >>
rect 40 112 41 113 
<< m1 >>
rect 41 112 42 113 
<< m1 >>
rect 42 112 43 113 
<< m1 >>
rect 43 112 44 113 
<< m1 >>
rect 44 112 45 113 
<< m1 >>
rect 46 112 47 113 
<< m2 >>
rect 47 112 48 113 
<< m1 >>
rect 48 112 49 113 
<< m2 >>
rect 48 112 49 113 
<< m2c >>
rect 48 112 49 113 
<< m1 >>
rect 48 112 49 113 
<< m2 >>
rect 48 112 49 113 
<< m1 >>
rect 49 112 50 113 
<< m1 >>
rect 50 112 51 113 
<< m1 >>
rect 52 112 53 113 
<< m1 >>
rect 55 112 56 113 
<< m1 >>
rect 59 112 60 113 
<< m2 >>
rect 61 112 62 113 
<< m1 >>
rect 62 112 63 113 
<< m1 >>
rect 64 112 65 113 
<< m1 >>
rect 73 112 74 113 
<< m1 >>
rect 78 112 79 113 
<< m2 >>
rect 81 112 82 113 
<< m1 >>
rect 82 112 83 113 
<< m1 >>
rect 91 112 92 113 
<< m2 >>
rect 92 112 93 113 
<< m1 >>
rect 109 112 110 113 
<< m2 >>
rect 109 112 110 113 
<< m1 >>
rect 115 112 116 113 
<< m1 >>
rect 130 112 131 113 
<< m1 >>
rect 132 112 133 113 
<< m1 >>
rect 136 112 137 113 
<< m2 >>
rect 136 112 137 113 
<< m1 >>
rect 145 112 146 113 
<< m2 >>
rect 145 112 146 113 
<< m1 >>
rect 147 112 148 113 
<< m1 >>
rect 163 112 164 113 
<< m1 >>
rect 167 112 168 113 
<< m2 >>
rect 169 112 170 113 
<< m1 >>
rect 170 112 171 113 
<< m1 >>
rect 172 112 173 113 
<< m1 >>
rect 175 112 176 113 
<< m1 >>
rect 176 112 177 113 
<< m1 >>
rect 177 112 178 113 
<< m1 >>
rect 178 112 179 113 
<< m1 >>
rect 179 112 180 113 
<< m1 >>
rect 180 112 181 113 
<< m1 >>
rect 181 112 182 113 
<< m1 >>
rect 182 112 183 113 
<< m1 >>
rect 183 112 184 113 
<< m1 >>
rect 184 112 185 113 
<< m1 >>
rect 185 112 186 113 
<< m1 >>
rect 186 112 187 113 
<< m1 >>
rect 187 112 188 113 
<< m1 >>
rect 188 112 189 113 
<< m1 >>
rect 189 112 190 113 
<< m1 >>
rect 190 112 191 113 
<< m1 >>
rect 199 112 200 113 
<< m1 >>
rect 201 112 202 113 
<< m2 >>
rect 202 112 203 113 
<< m1 >>
rect 205 112 206 113 
<< m1 >>
rect 226 112 227 113 
<< m2 >>
rect 226 112 227 113 
<< m1 >>
rect 235 112 236 113 
<< m2 >>
rect 235 112 236 113 
<< m1 >>
rect 244 112 245 113 
<< m1 >>
rect 256 112 257 113 
<< m2 >>
rect 256 112 257 113 
<< m2c >>
rect 256 112 257 113 
<< m1 >>
rect 256 112 257 113 
<< m2 >>
rect 256 112 257 113 
<< m2 >>
rect 257 112 258 113 
<< m1 >>
rect 258 112 259 113 
<< m2 >>
rect 258 112 259 113 
<< m2 >>
rect 259 112 260 113 
<< m1 >>
rect 260 112 261 113 
<< m2 >>
rect 260 112 261 113 
<< m2 >>
rect 261 112 262 113 
<< m1 >>
rect 262 112 263 113 
<< m2 >>
rect 262 112 263 113 
<< m2 >>
rect 263 112 264 113 
<< m1 >>
rect 264 112 265 113 
<< m2 >>
rect 264 112 265 113 
<< m2c >>
rect 264 112 265 113 
<< m1 >>
rect 264 112 265 113 
<< m2 >>
rect 264 112 265 113 
<< m1 >>
rect 265 112 266 113 
<< m1 >>
rect 266 112 267 113 
<< m1 >>
rect 267 112 268 113 
<< m1 >>
rect 268 112 269 113 
<< m1 >>
rect 269 112 270 113 
<< m1 >>
rect 271 112 272 113 
<< m1 >>
rect 274 112 275 113 
<< m1 >>
rect 276 112 277 113 
<< m1 >>
rect 278 112 279 113 
<< m1 >>
rect 296 112 297 113 
<< m1 >>
rect 307 112 308 113 
<< m2 >>
rect 308 112 309 113 
<< m1 >>
rect 316 112 317 113 
<< m1 >>
rect 318 112 319 113 
<< m1 >>
rect 319 112 320 113 
<< m1 >>
rect 320 112 321 113 
<< m1 >>
rect 321 112 322 113 
<< m1 >>
rect 322 112 323 113 
<< m1 >>
rect 323 112 324 113 
<< m1 >>
rect 324 112 325 113 
<< m1 >>
rect 325 112 326 113 
<< m2 >>
rect 325 112 326 113 
<< m2c >>
rect 325 112 326 113 
<< m1 >>
rect 325 112 326 113 
<< m2 >>
rect 325 112 326 113 
<< m2 >>
rect 326 112 327 113 
<< m1 >>
rect 327 112 328 113 
<< m2 >>
rect 327 112 328 113 
<< m2 >>
rect 328 112 329 113 
<< m1 >>
rect 329 112 330 113 
<< m2 >>
rect 329 112 330 113 
<< m2 >>
rect 330 112 331 113 
<< m1 >>
rect 331 112 332 113 
<< m2 >>
rect 331 112 332 113 
<< m2c >>
rect 331 112 332 113 
<< m1 >>
rect 331 112 332 113 
<< m2 >>
rect 331 112 332 113 
<< m1 >>
rect 10 113 11 114 
<< m1 >>
rect 19 113 20 114 
<< m2 >>
rect 19 113 20 114 
<< m1 >>
rect 21 113 22 114 
<< m1 >>
rect 23 113 24 114 
<< m2 >>
rect 27 113 28 114 
<< m1 >>
rect 28 113 29 114 
<< m1 >>
rect 31 113 32 114 
<< m2 >>
rect 37 113 38 114 
<< m1 >>
rect 46 113 47 114 
<< m2 >>
rect 47 113 48 114 
<< m1 >>
rect 52 113 53 114 
<< m1 >>
rect 55 113 56 114 
<< m1 >>
rect 59 113 60 114 
<< m2 >>
rect 61 113 62 114 
<< m1 >>
rect 62 113 63 114 
<< m1 >>
rect 64 113 65 114 
<< m1 >>
rect 73 113 74 114 
<< m1 >>
rect 78 113 79 114 
<< m2 >>
rect 81 113 82 114 
<< m1 >>
rect 82 113 83 114 
<< m1 >>
rect 91 113 92 114 
<< m2 >>
rect 92 113 93 114 
<< m1 >>
rect 109 113 110 114 
<< m2 >>
rect 109 113 110 114 
<< m1 >>
rect 115 113 116 114 
<< m1 >>
rect 130 113 131 114 
<< m1 >>
rect 132 113 133 114 
<< m1 >>
rect 136 113 137 114 
<< m2 >>
rect 136 113 137 114 
<< m1 >>
rect 145 113 146 114 
<< m2 >>
rect 145 113 146 114 
<< m1 >>
rect 147 113 148 114 
<< m1 >>
rect 163 113 164 114 
<< m1 >>
rect 167 113 168 114 
<< m2 >>
rect 169 113 170 114 
<< m1 >>
rect 170 113 171 114 
<< m1 >>
rect 172 113 173 114 
<< m1 >>
rect 175 113 176 114 
<< m1 >>
rect 199 113 200 114 
<< m1 >>
rect 201 113 202 114 
<< m2 >>
rect 202 113 203 114 
<< m1 >>
rect 205 113 206 114 
<< m1 >>
rect 226 113 227 114 
<< m2 >>
rect 226 113 227 114 
<< m1 >>
rect 235 113 236 114 
<< m2 >>
rect 235 113 236 114 
<< m1 >>
rect 244 113 245 114 
<< m1 >>
rect 258 113 259 114 
<< m1 >>
rect 260 113 261 114 
<< m1 >>
rect 262 113 263 114 
<< m1 >>
rect 271 113 272 114 
<< m1 >>
rect 274 113 275 114 
<< m1 >>
rect 276 113 277 114 
<< m1 >>
rect 278 113 279 114 
<< m1 >>
rect 296 113 297 114 
<< m2 >>
rect 296 113 297 114 
<< m2c >>
rect 296 113 297 114 
<< m1 >>
rect 296 113 297 114 
<< m2 >>
rect 296 113 297 114 
<< m1 >>
rect 307 113 308 114 
<< m2 >>
rect 308 113 309 114 
<< m1 >>
rect 316 113 317 114 
<< m1 >>
rect 327 113 328 114 
<< m1 >>
rect 329 113 330 114 
<< m1 >>
rect 331 113 332 114 
<< m1 >>
rect 10 114 11 115 
<< m1 >>
rect 19 114 20 115 
<< m2 >>
rect 19 114 20 115 
<< m1 >>
rect 21 114 22 115 
<< m1 >>
rect 23 114 24 115 
<< m2 >>
rect 27 114 28 115 
<< m1 >>
rect 28 114 29 115 
<< m1 >>
rect 31 114 32 115 
<< m1 >>
rect 37 114 38 115 
<< m2 >>
rect 37 114 38 115 
<< m2c >>
rect 37 114 38 115 
<< m1 >>
rect 37 114 38 115 
<< m2 >>
rect 37 114 38 115 
<< m1 >>
rect 42 114 43 115 
<< m1 >>
rect 43 114 44 115 
<< m1 >>
rect 44 114 45 115 
<< m2 >>
rect 44 114 45 115 
<< m2c >>
rect 44 114 45 115 
<< m1 >>
rect 44 114 45 115 
<< m2 >>
rect 44 114 45 115 
<< m2 >>
rect 45 114 46 115 
<< m1 >>
rect 46 114 47 115 
<< m2 >>
rect 46 114 47 115 
<< m2 >>
rect 47 114 48 115 
<< m1 >>
rect 52 114 53 115 
<< m1 >>
rect 55 114 56 115 
<< m1 >>
rect 59 114 60 115 
<< m2 >>
rect 61 114 62 115 
<< m1 >>
rect 62 114 63 115 
<< m1 >>
rect 64 114 65 115 
<< m1 >>
rect 73 114 74 115 
<< m1 >>
rect 78 114 79 115 
<< m2 >>
rect 81 114 82 115 
<< m1 >>
rect 82 114 83 115 
<< m1 >>
rect 91 114 92 115 
<< m2 >>
rect 92 114 93 115 
<< m1 >>
rect 109 114 110 115 
<< m2 >>
rect 109 114 110 115 
<< m1 >>
rect 115 114 116 115 
<< m1 >>
rect 130 114 131 115 
<< m1 >>
rect 132 114 133 115 
<< m1 >>
rect 136 114 137 115 
<< m2 >>
rect 136 114 137 115 
<< m1 >>
rect 145 114 146 115 
<< m2 >>
rect 145 114 146 115 
<< m1 >>
rect 147 114 148 115 
<< m1 >>
rect 163 114 164 115 
<< m1 >>
rect 167 114 168 115 
<< m2 >>
rect 167 114 168 115 
<< m2c >>
rect 167 114 168 115 
<< m1 >>
rect 167 114 168 115 
<< m2 >>
rect 167 114 168 115 
<< m2 >>
rect 169 114 170 115 
<< m1 >>
rect 170 114 171 115 
<< m2 >>
rect 170 114 171 115 
<< m2 >>
rect 171 114 172 115 
<< m1 >>
rect 172 114 173 115 
<< m2 >>
rect 172 114 173 115 
<< m2 >>
rect 173 114 174 115 
<< m2 >>
rect 174 114 175 115 
<< m1 >>
rect 175 114 176 115 
<< m2 >>
rect 175 114 176 115 
<< m2 >>
rect 176 114 177 115 
<< m1 >>
rect 177 114 178 115 
<< m2 >>
rect 177 114 178 115 
<< m2c >>
rect 177 114 178 115 
<< m1 >>
rect 177 114 178 115 
<< m2 >>
rect 177 114 178 115 
<< m1 >>
rect 178 114 179 115 
<< m1 >>
rect 179 114 180 115 
<< m1 >>
rect 180 114 181 115 
<< m1 >>
rect 181 114 182 115 
<< m1 >>
rect 199 114 200 115 
<< m1 >>
rect 201 114 202 115 
<< m2 >>
rect 202 114 203 115 
<< m1 >>
rect 205 114 206 115 
<< m1 >>
rect 226 114 227 115 
<< m2 >>
rect 226 114 227 115 
<< m1 >>
rect 235 114 236 115 
<< m2 >>
rect 235 114 236 115 
<< m1 >>
rect 244 114 245 115 
<< m1 >>
rect 258 114 259 115 
<< m1 >>
rect 260 114 261 115 
<< m1 >>
rect 262 114 263 115 
<< m1 >>
rect 271 114 272 115 
<< m1 >>
rect 274 114 275 115 
<< m1 >>
rect 276 114 277 115 
<< m1 >>
rect 278 114 279 115 
<< m2 >>
rect 296 114 297 115 
<< m2 >>
rect 300 114 301 115 
<< m2 >>
rect 301 114 302 115 
<< m2 >>
rect 302 114 303 115 
<< m2 >>
rect 303 114 304 115 
<< m2 >>
rect 304 114 305 115 
<< m2 >>
rect 305 114 306 115 
<< m2 >>
rect 306 114 307 115 
<< m1 >>
rect 307 114 308 115 
<< m2 >>
rect 307 114 308 115 
<< m2 >>
rect 308 114 309 115 
<< m1 >>
rect 316 114 317 115 
<< m1 >>
rect 327 114 328 115 
<< m1 >>
rect 329 114 330 115 
<< m1 >>
rect 331 114 332 115 
<< m1 >>
rect 10 115 11 116 
<< m1 >>
rect 19 115 20 116 
<< m2 >>
rect 19 115 20 116 
<< m1 >>
rect 21 115 22 116 
<< m1 >>
rect 23 115 24 116 
<< m2 >>
rect 27 115 28 116 
<< m1 >>
rect 28 115 29 116 
<< m1 >>
rect 31 115 32 116 
<< m1 >>
rect 37 115 38 116 
<< m1 >>
rect 42 115 43 116 
<< m1 >>
rect 46 115 47 116 
<< m1 >>
rect 52 115 53 116 
<< m1 >>
rect 55 115 56 116 
<< m1 >>
rect 59 115 60 116 
<< m2 >>
rect 61 115 62 116 
<< m1 >>
rect 62 115 63 116 
<< m1 >>
rect 64 115 65 116 
<< m1 >>
rect 73 115 74 116 
<< m1 >>
rect 78 115 79 116 
<< m2 >>
rect 81 115 82 116 
<< m1 >>
rect 82 115 83 116 
<< m1 >>
rect 91 115 92 116 
<< m2 >>
rect 92 115 93 116 
<< m1 >>
rect 109 115 110 116 
<< m2 >>
rect 109 115 110 116 
<< m1 >>
rect 115 115 116 116 
<< m1 >>
rect 130 115 131 116 
<< m1 >>
rect 132 115 133 116 
<< m1 >>
rect 136 115 137 116 
<< m2 >>
rect 136 115 137 116 
<< m1 >>
rect 145 115 146 116 
<< m2 >>
rect 145 115 146 116 
<< m1 >>
rect 147 115 148 116 
<< m1 >>
rect 154 115 155 116 
<< m1 >>
rect 155 115 156 116 
<< m1 >>
rect 156 115 157 116 
<< m1 >>
rect 157 115 158 116 
<< m1 >>
rect 158 115 159 116 
<< m1 >>
rect 159 115 160 116 
<< m1 >>
rect 160 115 161 116 
<< m1 >>
rect 161 115 162 116 
<< m1 >>
rect 163 115 164 116 
<< m2 >>
rect 167 115 168 116 
<< m1 >>
rect 170 115 171 116 
<< m1 >>
rect 172 115 173 116 
<< m1 >>
rect 175 115 176 116 
<< m1 >>
rect 181 115 182 116 
<< m1 >>
rect 199 115 200 116 
<< m1 >>
rect 201 115 202 116 
<< m2 >>
rect 202 115 203 116 
<< m1 >>
rect 205 115 206 116 
<< m1 >>
rect 226 115 227 116 
<< m2 >>
rect 226 115 227 116 
<< m1 >>
rect 235 115 236 116 
<< m2 >>
rect 235 115 236 116 
<< m1 >>
rect 244 115 245 116 
<< m1 >>
rect 253 115 254 116 
<< m1 >>
rect 254 115 255 116 
<< m1 >>
rect 255 115 256 116 
<< m1 >>
rect 256 115 257 116 
<< m2 >>
rect 256 115 257 116 
<< m2c >>
rect 256 115 257 116 
<< m1 >>
rect 256 115 257 116 
<< m2 >>
rect 256 115 257 116 
<< m2 >>
rect 257 115 258 116 
<< m1 >>
rect 258 115 259 116 
<< m2 >>
rect 258 115 259 116 
<< m2 >>
rect 259 115 260 116 
<< m1 >>
rect 260 115 261 116 
<< m2 >>
rect 260 115 261 116 
<< m2 >>
rect 261 115 262 116 
<< m1 >>
rect 262 115 263 116 
<< m2 >>
rect 262 115 263 116 
<< m2 >>
rect 263 115 264 116 
<< m1 >>
rect 264 115 265 116 
<< m2 >>
rect 264 115 265 116 
<< m1 >>
rect 265 115 266 116 
<< m2 >>
rect 265 115 266 116 
<< m1 >>
rect 266 115 267 116 
<< m2 >>
rect 266 115 267 116 
<< m1 >>
rect 267 115 268 116 
<< m2 >>
rect 267 115 268 116 
<< m1 >>
rect 268 115 269 116 
<< m2 >>
rect 268 115 269 116 
<< m1 >>
rect 269 115 270 116 
<< m2 >>
rect 269 115 270 116 
<< m1 >>
rect 270 115 271 116 
<< m2 >>
rect 270 115 271 116 
<< m1 >>
rect 271 115 272 116 
<< m2 >>
rect 271 115 272 116 
<< m2 >>
rect 272 115 273 116 
<< m2 >>
rect 273 115 274 116 
<< m1 >>
rect 274 115 275 116 
<< m2 >>
rect 274 115 275 116 
<< m2 >>
rect 275 115 276 116 
<< m1 >>
rect 276 115 277 116 
<< m2 >>
rect 276 115 277 116 
<< m2 >>
rect 277 115 278 116 
<< m1 >>
rect 278 115 279 116 
<< m2 >>
rect 278 115 279 116 
<< m2 >>
rect 279 115 280 116 
<< m1 >>
rect 280 115 281 116 
<< m2 >>
rect 280 115 281 116 
<< m2c >>
rect 280 115 281 116 
<< m1 >>
rect 280 115 281 116 
<< m2 >>
rect 280 115 281 116 
<< m1 >>
rect 281 115 282 116 
<< m1 >>
rect 282 115 283 116 
<< m2 >>
rect 282 115 283 116 
<< m1 >>
rect 283 115 284 116 
<< m2 >>
rect 283 115 284 116 
<< m1 >>
rect 284 115 285 116 
<< m2 >>
rect 284 115 285 116 
<< m1 >>
rect 285 115 286 116 
<< m1 >>
rect 286 115 287 116 
<< m1 >>
rect 287 115 288 116 
<< m1 >>
rect 288 115 289 116 
<< m1 >>
rect 289 115 290 116 
<< m1 >>
rect 290 115 291 116 
<< m1 >>
rect 291 115 292 116 
<< m1 >>
rect 292 115 293 116 
<< m1 >>
rect 293 115 294 116 
<< m1 >>
rect 294 115 295 116 
<< m1 >>
rect 295 115 296 116 
<< m1 >>
rect 296 115 297 116 
<< m2 >>
rect 296 115 297 116 
<< m1 >>
rect 297 115 298 116 
<< m1 >>
rect 298 115 299 116 
<< m1 >>
rect 299 115 300 116 
<< m1 >>
rect 300 115 301 116 
<< m2 >>
rect 300 115 301 116 
<< m1 >>
rect 301 115 302 116 
<< m1 >>
rect 302 115 303 116 
<< m1 >>
rect 303 115 304 116 
<< m1 >>
rect 304 115 305 116 
<< m1 >>
rect 305 115 306 116 
<< m1 >>
rect 307 115 308 116 
<< m1 >>
rect 316 115 317 116 
<< m1 >>
rect 327 115 328 116 
<< m1 >>
rect 329 115 330 116 
<< m1 >>
rect 331 115 332 116 
<< m1 >>
rect 10 116 11 117 
<< m1 >>
rect 19 116 20 117 
<< m2 >>
rect 19 116 20 117 
<< m1 >>
rect 21 116 22 117 
<< m1 >>
rect 23 116 24 117 
<< m2 >>
rect 27 116 28 117 
<< m1 >>
rect 28 116 29 117 
<< m1 >>
rect 31 116 32 117 
<< m1 >>
rect 37 116 38 117 
<< m1 >>
rect 42 116 43 117 
<< m1 >>
rect 46 116 47 117 
<< m1 >>
rect 52 116 53 117 
<< m1 >>
rect 55 116 56 117 
<< m1 >>
rect 59 116 60 117 
<< m2 >>
rect 61 116 62 117 
<< m1 >>
rect 62 116 63 117 
<< m1 >>
rect 64 116 65 117 
<< m1 >>
rect 73 116 74 117 
<< m1 >>
rect 78 116 79 117 
<< m2 >>
rect 81 116 82 117 
<< m1 >>
rect 82 116 83 117 
<< m1 >>
rect 91 116 92 117 
<< m2 >>
rect 92 116 93 117 
<< m1 >>
rect 109 116 110 117 
<< m2 >>
rect 109 116 110 117 
<< m1 >>
rect 115 116 116 117 
<< m1 >>
rect 130 116 131 117 
<< m1 >>
rect 132 116 133 117 
<< m1 >>
rect 136 116 137 117 
<< m2 >>
rect 136 116 137 117 
<< m1 >>
rect 145 116 146 117 
<< m2 >>
rect 145 116 146 117 
<< m1 >>
rect 147 116 148 117 
<< m1 >>
rect 154 116 155 117 
<< m1 >>
rect 161 116 162 117 
<< m2 >>
rect 161 116 162 117 
<< m2c >>
rect 161 116 162 117 
<< m1 >>
rect 161 116 162 117 
<< m2 >>
rect 161 116 162 117 
<< m2 >>
rect 162 116 163 117 
<< m1 >>
rect 163 116 164 117 
<< m2 >>
rect 163 116 164 117 
<< m2 >>
rect 164 116 165 117 
<< m1 >>
rect 165 116 166 117 
<< m2 >>
rect 165 116 166 117 
<< m2c >>
rect 165 116 166 117 
<< m1 >>
rect 165 116 166 117 
<< m2 >>
rect 165 116 166 117 
<< m1 >>
rect 166 116 167 117 
<< m1 >>
rect 167 116 168 117 
<< m2 >>
rect 167 116 168 117 
<< m1 >>
rect 168 116 169 117 
<< m1 >>
rect 170 116 171 117 
<< m1 >>
rect 172 116 173 117 
<< m1 >>
rect 175 116 176 117 
<< m1 >>
rect 181 116 182 117 
<< m1 >>
rect 199 116 200 117 
<< m1 >>
rect 201 116 202 117 
<< m2 >>
rect 202 116 203 117 
<< m1 >>
rect 205 116 206 117 
<< m1 >>
rect 226 116 227 117 
<< m2 >>
rect 226 116 227 117 
<< m1 >>
rect 235 116 236 117 
<< m2 >>
rect 235 116 236 117 
<< m1 >>
rect 244 116 245 117 
<< m1 >>
rect 253 116 254 117 
<< m1 >>
rect 258 116 259 117 
<< m1 >>
rect 260 116 261 117 
<< m1 >>
rect 262 116 263 117 
<< m1 >>
rect 264 116 265 117 
<< m1 >>
rect 274 116 275 117 
<< m1 >>
rect 276 116 277 117 
<< m1 >>
rect 278 116 279 117 
<< m2 >>
rect 282 116 283 117 
<< m2 >>
rect 284 116 285 117 
<< m2 >>
rect 296 116 297 117 
<< m2 >>
rect 300 116 301 117 
<< m1 >>
rect 305 116 306 117 
<< m1 >>
rect 307 116 308 117 
<< m1 >>
rect 316 116 317 117 
<< m1 >>
rect 327 116 328 117 
<< m1 >>
rect 329 116 330 117 
<< m1 >>
rect 331 116 332 117 
<< m1 >>
rect 10 117 11 118 
<< m1 >>
rect 19 117 20 118 
<< m2 >>
rect 19 117 20 118 
<< m1 >>
rect 21 117 22 118 
<< m1 >>
rect 23 117 24 118 
<< m2 >>
rect 27 117 28 118 
<< m1 >>
rect 28 117 29 118 
<< m1 >>
rect 31 117 32 118 
<< m1 >>
rect 37 117 38 118 
<< m1 >>
rect 42 117 43 118 
<< m1 >>
rect 46 117 47 118 
<< m1 >>
rect 52 117 53 118 
<< m1 >>
rect 53 117 54 118 
<< m1 >>
rect 55 117 56 118 
<< m1 >>
rect 59 117 60 118 
<< m2 >>
rect 61 117 62 118 
<< m1 >>
rect 62 117 63 118 
<< m1 >>
rect 64 117 65 118 
<< m1 >>
rect 73 117 74 118 
<< m1 >>
rect 78 117 79 118 
<< m2 >>
rect 81 117 82 118 
<< m1 >>
rect 82 117 83 118 
<< m1 >>
rect 91 117 92 118 
<< m2 >>
rect 92 117 93 118 
<< m1 >>
rect 109 117 110 118 
<< m2 >>
rect 109 117 110 118 
<< m1 >>
rect 115 117 116 118 
<< m1 >>
rect 130 117 131 118 
<< m1 >>
rect 132 117 133 118 
<< m1 >>
rect 136 117 137 118 
<< m2 >>
rect 136 117 137 118 
<< m1 >>
rect 145 117 146 118 
<< m2 >>
rect 145 117 146 118 
<< m1 >>
rect 147 117 148 118 
<< m1 >>
rect 154 117 155 118 
<< m1 >>
rect 163 117 164 118 
<< m2 >>
rect 167 117 168 118 
<< m1 >>
rect 168 117 169 118 
<< m1 >>
rect 170 117 171 118 
<< m1 >>
rect 172 117 173 118 
<< m1 >>
rect 175 117 176 118 
<< m1 >>
rect 181 117 182 118 
<< m1 >>
rect 199 117 200 118 
<< m1 >>
rect 201 117 202 118 
<< m2 >>
rect 202 117 203 118 
<< m1 >>
rect 205 117 206 118 
<< m1 >>
rect 226 117 227 118 
<< m2 >>
rect 226 117 227 118 
<< m1 >>
rect 235 117 236 118 
<< m2 >>
rect 235 117 236 118 
<< m1 >>
rect 244 117 245 118 
<< m1 >>
rect 253 117 254 118 
<< m1 >>
rect 258 117 259 118 
<< m1 >>
rect 260 117 261 118 
<< m1 >>
rect 262 117 263 118 
<< m1 >>
rect 264 117 265 118 
<< m1 >>
rect 274 117 275 118 
<< m1 >>
rect 276 117 277 118 
<< m1 >>
rect 278 117 279 118 
<< m1 >>
rect 282 117 283 118 
<< m2 >>
rect 282 117 283 118 
<< m2c >>
rect 282 117 283 118 
<< m1 >>
rect 282 117 283 118 
<< m2 >>
rect 282 117 283 118 
<< m1 >>
rect 284 117 285 118 
<< m2 >>
rect 284 117 285 118 
<< m2c >>
rect 284 117 285 118 
<< m1 >>
rect 284 117 285 118 
<< m2 >>
rect 284 117 285 118 
<< m1 >>
rect 285 117 286 118 
<< m1 >>
rect 286 117 287 118 
<< m1 >>
rect 287 117 288 118 
<< m1 >>
rect 288 117 289 118 
<< m1 >>
rect 289 117 290 118 
<< m1 >>
rect 296 117 297 118 
<< m2 >>
rect 296 117 297 118 
<< m2c >>
rect 296 117 297 118 
<< m1 >>
rect 296 117 297 118 
<< m2 >>
rect 296 117 297 118 
<< m1 >>
rect 298 117 299 118 
<< m1 >>
rect 299 117 300 118 
<< m1 >>
rect 300 117 301 118 
<< m2 >>
rect 300 117 301 118 
<< m2c >>
rect 300 117 301 118 
<< m1 >>
rect 300 117 301 118 
<< m2 >>
rect 300 117 301 118 
<< m1 >>
rect 305 117 306 118 
<< m1 >>
rect 307 117 308 118 
<< m1 >>
rect 316 117 317 118 
<< m1 >>
rect 327 117 328 118 
<< m1 >>
rect 329 117 330 118 
<< m1 >>
rect 331 117 332 118 
<< m1 >>
rect 10 118 11 119 
<< m1 >>
rect 19 118 20 119 
<< m2 >>
rect 19 118 20 119 
<< m1 >>
rect 21 118 22 119 
<< m1 >>
rect 23 118 24 119 
<< m2 >>
rect 27 118 28 119 
<< m1 >>
rect 28 118 29 119 
<< m1 >>
rect 31 118 32 119 
<< m1 >>
rect 37 118 38 119 
<< m1 >>
rect 42 118 43 119 
<< m1 >>
rect 46 118 47 119 
<< m1 >>
rect 53 118 54 119 
<< m2 >>
rect 53 118 54 119 
<< m2c >>
rect 53 118 54 119 
<< m1 >>
rect 53 118 54 119 
<< m2 >>
rect 53 118 54 119 
<< m2 >>
rect 54 118 55 119 
<< m1 >>
rect 55 118 56 119 
<< m2 >>
rect 55 118 56 119 
<< m2 >>
rect 56 118 57 119 
<< m1 >>
rect 59 118 60 119 
<< m2 >>
rect 61 118 62 119 
<< m1 >>
rect 62 118 63 119 
<< m1 >>
rect 64 118 65 119 
<< m1 >>
rect 73 118 74 119 
<< m1 >>
rect 78 118 79 119 
<< m2 >>
rect 81 118 82 119 
<< m1 >>
rect 82 118 83 119 
<< m1 >>
rect 91 118 92 119 
<< m2 >>
rect 92 118 93 119 
<< m1 >>
rect 106 118 107 119 
<< m1 >>
rect 107 118 108 119 
<< m2 >>
rect 107 118 108 119 
<< m2c >>
rect 107 118 108 119 
<< m1 >>
rect 107 118 108 119 
<< m2 >>
rect 107 118 108 119 
<< m2 >>
rect 108 118 109 119 
<< m1 >>
rect 109 118 110 119 
<< m2 >>
rect 109 118 110 119 
<< m1 >>
rect 115 118 116 119 
<< m1 >>
rect 130 118 131 119 
<< m1 >>
rect 132 118 133 119 
<< m1 >>
rect 136 118 137 119 
<< m2 >>
rect 136 118 137 119 
<< m1 >>
rect 145 118 146 119 
<< m2 >>
rect 145 118 146 119 
<< m1 >>
rect 147 118 148 119 
<< m1 >>
rect 154 118 155 119 
<< m1 >>
rect 160 118 161 119 
<< m1 >>
rect 161 118 162 119 
<< m2 >>
rect 161 118 162 119 
<< m2c >>
rect 161 118 162 119 
<< m1 >>
rect 161 118 162 119 
<< m2 >>
rect 161 118 162 119 
<< m2 >>
rect 162 118 163 119 
<< m1 >>
rect 163 118 164 119 
<< m2 >>
rect 163 118 164 119 
<< m2 >>
rect 164 118 165 119 
<< m2 >>
rect 167 118 168 119 
<< m1 >>
rect 168 118 169 119 
<< m1 >>
rect 170 118 171 119 
<< m1 >>
rect 172 118 173 119 
<< m1 >>
rect 175 118 176 119 
<< m1 >>
rect 181 118 182 119 
<< m1 >>
rect 199 118 200 119 
<< m1 >>
rect 201 118 202 119 
<< m2 >>
rect 202 118 203 119 
<< m1 >>
rect 205 118 206 119 
<< m1 >>
rect 226 118 227 119 
<< m2 >>
rect 226 118 227 119 
<< m1 >>
rect 235 118 236 119 
<< m2 >>
rect 235 118 236 119 
<< m1 >>
rect 244 118 245 119 
<< m1 >>
rect 253 118 254 119 
<< m2 >>
rect 257 118 258 119 
<< m1 >>
rect 258 118 259 119 
<< m2 >>
rect 258 118 259 119 
<< m2 >>
rect 259 118 260 119 
<< m1 >>
rect 260 118 261 119 
<< m2 >>
rect 260 118 261 119 
<< m2 >>
rect 261 118 262 119 
<< m1 >>
rect 262 118 263 119 
<< m2 >>
rect 262 118 263 119 
<< m2 >>
rect 263 118 264 119 
<< m1 >>
rect 264 118 265 119 
<< m2 >>
rect 264 118 265 119 
<< m2c >>
rect 264 118 265 119 
<< m1 >>
rect 264 118 265 119 
<< m2 >>
rect 264 118 265 119 
<< m1 >>
rect 274 118 275 119 
<< m1 >>
rect 276 118 277 119 
<< m1 >>
rect 278 118 279 119 
<< m1 >>
rect 280 118 281 119 
<< m1 >>
rect 281 118 282 119 
<< m1 >>
rect 282 118 283 119 
<< m1 >>
rect 289 118 290 119 
<< m1 >>
rect 296 118 297 119 
<< m1 >>
rect 298 118 299 119 
<< m1 >>
rect 305 118 306 119 
<< m2 >>
rect 305 118 306 119 
<< m2c >>
rect 305 118 306 119 
<< m1 >>
rect 305 118 306 119 
<< m2 >>
rect 305 118 306 119 
<< m2 >>
rect 306 118 307 119 
<< m1 >>
rect 307 118 308 119 
<< m2 >>
rect 307 118 308 119 
<< m2 >>
rect 308 118 309 119 
<< m1 >>
rect 316 118 317 119 
<< m1 >>
rect 327 118 328 119 
<< m1 >>
rect 329 118 330 119 
<< m1 >>
rect 331 118 332 119 
<< m1 >>
rect 340 118 341 119 
<< m1 >>
rect 341 118 342 119 
<< m1 >>
rect 342 118 343 119 
<< m1 >>
rect 343 118 344 119 
<< m1 >>
rect 344 118 345 119 
<< m1 >>
rect 345 118 346 119 
<< m1 >>
rect 10 119 11 120 
<< m1 >>
rect 19 119 20 120 
<< m2 >>
rect 19 119 20 120 
<< m1 >>
rect 21 119 22 120 
<< m1 >>
rect 23 119 24 120 
<< m2 >>
rect 27 119 28 120 
<< m1 >>
rect 28 119 29 120 
<< m1 >>
rect 31 119 32 120 
<< m1 >>
rect 37 119 38 120 
<< m1 >>
rect 42 119 43 120 
<< m1 >>
rect 46 119 47 120 
<< m1 >>
rect 55 119 56 120 
<< m2 >>
rect 56 119 57 120 
<< m1 >>
rect 59 119 60 120 
<< m2 >>
rect 61 119 62 120 
<< m1 >>
rect 62 119 63 120 
<< m1 >>
rect 64 119 65 120 
<< m1 >>
rect 73 119 74 120 
<< m1 >>
rect 78 119 79 120 
<< m2 >>
rect 81 119 82 120 
<< m1 >>
rect 82 119 83 120 
<< m1 >>
rect 91 119 92 120 
<< m2 >>
rect 92 119 93 120 
<< m1 >>
rect 106 119 107 120 
<< m1 >>
rect 109 119 110 120 
<< m1 >>
rect 115 119 116 120 
<< m1 >>
rect 130 119 131 120 
<< m1 >>
rect 132 119 133 120 
<< m1 >>
rect 136 119 137 120 
<< m2 >>
rect 136 119 137 120 
<< m1 >>
rect 145 119 146 120 
<< m2 >>
rect 145 119 146 120 
<< m1 >>
rect 147 119 148 120 
<< m1 >>
rect 154 119 155 120 
<< m1 >>
rect 160 119 161 120 
<< m1 >>
rect 163 119 164 120 
<< m2 >>
rect 164 119 165 120 
<< m2 >>
rect 167 119 168 120 
<< m1 >>
rect 168 119 169 120 
<< m1 >>
rect 170 119 171 120 
<< m1 >>
rect 172 119 173 120 
<< m1 >>
rect 175 119 176 120 
<< m1 >>
rect 181 119 182 120 
<< m1 >>
rect 199 119 200 120 
<< m1 >>
rect 201 119 202 120 
<< m2 >>
rect 202 119 203 120 
<< m1 >>
rect 205 119 206 120 
<< m1 >>
rect 226 119 227 120 
<< m2 >>
rect 226 119 227 120 
<< m1 >>
rect 235 119 236 120 
<< m2 >>
rect 235 119 236 120 
<< m1 >>
rect 244 119 245 120 
<< m1 >>
rect 253 119 254 120 
<< m2 >>
rect 257 119 258 120 
<< m1 >>
rect 258 119 259 120 
<< m1 >>
rect 260 119 261 120 
<< m1 >>
rect 262 119 263 120 
<< m1 >>
rect 274 119 275 120 
<< m1 >>
rect 276 119 277 120 
<< m1 >>
rect 278 119 279 120 
<< m1 >>
rect 280 119 281 120 
<< m1 >>
rect 289 119 290 120 
<< m1 >>
rect 296 119 297 120 
<< m1 >>
rect 298 119 299 120 
<< m1 >>
rect 307 119 308 120 
<< m2 >>
rect 308 119 309 120 
<< m1 >>
rect 316 119 317 120 
<< m1 >>
rect 327 119 328 120 
<< m1 >>
rect 329 119 330 120 
<< m1 >>
rect 331 119 332 120 
<< m1 >>
rect 340 119 341 120 
<< m1 >>
rect 345 119 346 120 
<< m1 >>
rect 10 120 11 121 
<< pdiffusion >>
rect 12 120 13 121 
<< pdiffusion >>
rect 13 120 14 121 
<< pdiffusion >>
rect 14 120 15 121 
<< pdiffusion >>
rect 15 120 16 121 
<< pdiffusion >>
rect 16 120 17 121 
<< pdiffusion >>
rect 17 120 18 121 
<< m1 >>
rect 19 120 20 121 
<< m2 >>
rect 19 120 20 121 
<< m1 >>
rect 21 120 22 121 
<< m1 >>
rect 23 120 24 121 
<< m2 >>
rect 27 120 28 121 
<< m1 >>
rect 28 120 29 121 
<< pdiffusion >>
rect 30 120 31 121 
<< m1 >>
rect 31 120 32 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< m1 >>
rect 37 120 38 121 
<< m1 >>
rect 42 120 43 121 
<< m1 >>
rect 46 120 47 121 
<< pdiffusion >>
rect 48 120 49 121 
<< pdiffusion >>
rect 49 120 50 121 
<< pdiffusion >>
rect 50 120 51 121 
<< pdiffusion >>
rect 51 120 52 121 
<< pdiffusion >>
rect 52 120 53 121 
<< pdiffusion >>
rect 53 120 54 121 
<< m1 >>
rect 55 120 56 121 
<< m2 >>
rect 56 120 57 121 
<< m1 >>
rect 59 120 60 121 
<< m2 >>
rect 61 120 62 121 
<< m1 >>
rect 62 120 63 121 
<< m1 >>
rect 64 120 65 121 
<< pdiffusion >>
rect 66 120 67 121 
<< pdiffusion >>
rect 67 120 68 121 
<< pdiffusion >>
rect 68 120 69 121 
<< pdiffusion >>
rect 69 120 70 121 
<< pdiffusion >>
rect 70 120 71 121 
<< pdiffusion >>
rect 71 120 72 121 
<< m1 >>
rect 73 120 74 121 
<< m1 >>
rect 78 120 79 121 
<< m2 >>
rect 81 120 82 121 
<< m1 >>
rect 82 120 83 121 
<< pdiffusion >>
rect 84 120 85 121 
<< pdiffusion >>
rect 85 120 86 121 
<< pdiffusion >>
rect 86 120 87 121 
<< pdiffusion >>
rect 87 120 88 121 
<< pdiffusion >>
rect 88 120 89 121 
<< pdiffusion >>
rect 89 120 90 121 
<< m1 >>
rect 91 120 92 121 
<< m2 >>
rect 92 120 93 121 
<< pdiffusion >>
rect 102 120 103 121 
<< pdiffusion >>
rect 103 120 104 121 
<< pdiffusion >>
rect 104 120 105 121 
<< pdiffusion >>
rect 105 120 106 121 
<< m1 >>
rect 106 120 107 121 
<< pdiffusion >>
rect 106 120 107 121 
<< pdiffusion >>
rect 107 120 108 121 
<< m1 >>
rect 109 120 110 121 
<< m2 >>
rect 110 120 111 121 
<< m1 >>
rect 111 120 112 121 
<< m2 >>
rect 111 120 112 121 
<< m2c >>
rect 111 120 112 121 
<< m1 >>
rect 111 120 112 121 
<< m2 >>
rect 111 120 112 121 
<< m1 >>
rect 112 120 113 121 
<< m1 >>
rect 113 120 114 121 
<< m1 >>
rect 114 120 115 121 
<< m1 >>
rect 115 120 116 121 
<< pdiffusion >>
rect 120 120 121 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< m1 >>
rect 130 120 131 121 
<< m1 >>
rect 132 120 133 121 
<< m1 >>
rect 136 120 137 121 
<< m2 >>
rect 136 120 137 121 
<< pdiffusion >>
rect 138 120 139 121 
<< pdiffusion >>
rect 139 120 140 121 
<< pdiffusion >>
rect 140 120 141 121 
<< pdiffusion >>
rect 141 120 142 121 
<< pdiffusion >>
rect 142 120 143 121 
<< pdiffusion >>
rect 143 120 144 121 
<< m1 >>
rect 145 120 146 121 
<< m2 >>
rect 145 120 146 121 
<< m1 >>
rect 147 120 148 121 
<< m1 >>
rect 154 120 155 121 
<< pdiffusion >>
rect 156 120 157 121 
<< pdiffusion >>
rect 157 120 158 121 
<< pdiffusion >>
rect 158 120 159 121 
<< pdiffusion >>
rect 159 120 160 121 
<< m1 >>
rect 160 120 161 121 
<< pdiffusion >>
rect 160 120 161 121 
<< pdiffusion >>
rect 161 120 162 121 
<< m1 >>
rect 163 120 164 121 
<< m2 >>
rect 164 120 165 121 
<< m2 >>
rect 167 120 168 121 
<< m1 >>
rect 168 120 169 121 
<< m1 >>
rect 170 120 171 121 
<< m1 >>
rect 172 120 173 121 
<< pdiffusion >>
rect 174 120 175 121 
<< m1 >>
rect 175 120 176 121 
<< pdiffusion >>
rect 175 120 176 121 
<< pdiffusion >>
rect 176 120 177 121 
<< pdiffusion >>
rect 177 120 178 121 
<< pdiffusion >>
rect 178 120 179 121 
<< pdiffusion >>
rect 179 120 180 121 
<< m1 >>
rect 181 120 182 121 
<< pdiffusion >>
rect 192 120 193 121 
<< pdiffusion >>
rect 193 120 194 121 
<< pdiffusion >>
rect 194 120 195 121 
<< pdiffusion >>
rect 195 120 196 121 
<< pdiffusion >>
rect 196 120 197 121 
<< pdiffusion >>
rect 197 120 198 121 
<< m1 >>
rect 199 120 200 121 
<< m1 >>
rect 201 120 202 121 
<< m2 >>
rect 202 120 203 121 
<< m1 >>
rect 205 120 206 121 
<< pdiffusion >>
rect 210 120 211 121 
<< pdiffusion >>
rect 211 120 212 121 
<< pdiffusion >>
rect 212 120 213 121 
<< pdiffusion >>
rect 213 120 214 121 
<< pdiffusion >>
rect 214 120 215 121 
<< pdiffusion >>
rect 215 120 216 121 
<< m1 >>
rect 226 120 227 121 
<< m2 >>
rect 226 120 227 121 
<< pdiffusion >>
rect 228 120 229 121 
<< pdiffusion >>
rect 229 120 230 121 
<< pdiffusion >>
rect 230 120 231 121 
<< pdiffusion >>
rect 231 120 232 121 
<< pdiffusion >>
rect 232 120 233 121 
<< pdiffusion >>
rect 233 120 234 121 
<< m1 >>
rect 235 120 236 121 
<< m2 >>
rect 235 120 236 121 
<< m1 >>
rect 244 120 245 121 
<< pdiffusion >>
rect 246 120 247 121 
<< pdiffusion >>
rect 247 120 248 121 
<< pdiffusion >>
rect 248 120 249 121 
<< pdiffusion >>
rect 249 120 250 121 
<< pdiffusion >>
rect 250 120 251 121 
<< pdiffusion >>
rect 251 120 252 121 
<< m1 >>
rect 253 120 254 121 
<< m2 >>
rect 257 120 258 121 
<< m1 >>
rect 258 120 259 121 
<< m1 >>
rect 260 120 261 121 
<< m1 >>
rect 262 120 263 121 
<< pdiffusion >>
rect 264 120 265 121 
<< pdiffusion >>
rect 265 120 266 121 
<< pdiffusion >>
rect 266 120 267 121 
<< pdiffusion >>
rect 267 120 268 121 
<< pdiffusion >>
rect 268 120 269 121 
<< pdiffusion >>
rect 269 120 270 121 
<< m1 >>
rect 274 120 275 121 
<< m1 >>
rect 276 120 277 121 
<< m1 >>
rect 278 120 279 121 
<< m1 >>
rect 280 120 281 121 
<< pdiffusion >>
rect 282 120 283 121 
<< pdiffusion >>
rect 283 120 284 121 
<< pdiffusion >>
rect 284 120 285 121 
<< pdiffusion >>
rect 285 120 286 121 
<< pdiffusion >>
rect 286 120 287 121 
<< pdiffusion >>
rect 287 120 288 121 
<< m1 >>
rect 289 120 290 121 
<< m1 >>
rect 296 120 297 121 
<< m1 >>
rect 298 120 299 121 
<< pdiffusion >>
rect 300 120 301 121 
<< pdiffusion >>
rect 301 120 302 121 
<< pdiffusion >>
rect 302 120 303 121 
<< pdiffusion >>
rect 303 120 304 121 
<< pdiffusion >>
rect 304 120 305 121 
<< pdiffusion >>
rect 305 120 306 121 
<< m1 >>
rect 307 120 308 121 
<< m2 >>
rect 308 120 309 121 
<< m1 >>
rect 316 120 317 121 
<< pdiffusion >>
rect 318 120 319 121 
<< pdiffusion >>
rect 319 120 320 121 
<< pdiffusion >>
rect 320 120 321 121 
<< pdiffusion >>
rect 321 120 322 121 
<< pdiffusion >>
rect 322 120 323 121 
<< pdiffusion >>
rect 323 120 324 121 
<< m1 >>
rect 327 120 328 121 
<< m1 >>
rect 329 120 330 121 
<< m1 >>
rect 331 120 332 121 
<< pdiffusion >>
rect 336 120 337 121 
<< pdiffusion >>
rect 337 120 338 121 
<< pdiffusion >>
rect 338 120 339 121 
<< pdiffusion >>
rect 339 120 340 121 
<< m1 >>
rect 340 120 341 121 
<< pdiffusion >>
rect 340 120 341 121 
<< pdiffusion >>
rect 341 120 342 121 
<< m1 >>
rect 345 120 346 121 
<< m1 >>
rect 10 121 11 122 
<< pdiffusion >>
rect 12 121 13 122 
<< pdiffusion >>
rect 13 121 14 122 
<< pdiffusion >>
rect 14 121 15 122 
<< pdiffusion >>
rect 15 121 16 122 
<< pdiffusion >>
rect 16 121 17 122 
<< pdiffusion >>
rect 17 121 18 122 
<< m1 >>
rect 19 121 20 122 
<< m2 >>
rect 19 121 20 122 
<< m1 >>
rect 21 121 22 122 
<< m1 >>
rect 23 121 24 122 
<< m2 >>
rect 27 121 28 122 
<< m1 >>
rect 28 121 29 122 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< m1 >>
rect 37 121 38 122 
<< m1 >>
rect 42 121 43 122 
<< m1 >>
rect 46 121 47 122 
<< pdiffusion >>
rect 48 121 49 122 
<< pdiffusion >>
rect 49 121 50 122 
<< pdiffusion >>
rect 50 121 51 122 
<< pdiffusion >>
rect 51 121 52 122 
<< pdiffusion >>
rect 52 121 53 122 
<< pdiffusion >>
rect 53 121 54 122 
<< m1 >>
rect 55 121 56 122 
<< m2 >>
rect 56 121 57 122 
<< m1 >>
rect 59 121 60 122 
<< m2 >>
rect 61 121 62 122 
<< m1 >>
rect 62 121 63 122 
<< m1 >>
rect 64 121 65 122 
<< pdiffusion >>
rect 66 121 67 122 
<< pdiffusion >>
rect 67 121 68 122 
<< pdiffusion >>
rect 68 121 69 122 
<< pdiffusion >>
rect 69 121 70 122 
<< pdiffusion >>
rect 70 121 71 122 
<< pdiffusion >>
rect 71 121 72 122 
<< m1 >>
rect 73 121 74 122 
<< m1 >>
rect 78 121 79 122 
<< m2 >>
rect 81 121 82 122 
<< m1 >>
rect 82 121 83 122 
<< pdiffusion >>
rect 84 121 85 122 
<< pdiffusion >>
rect 85 121 86 122 
<< pdiffusion >>
rect 86 121 87 122 
<< pdiffusion >>
rect 87 121 88 122 
<< pdiffusion >>
rect 88 121 89 122 
<< pdiffusion >>
rect 89 121 90 122 
<< m1 >>
rect 91 121 92 122 
<< m2 >>
rect 92 121 93 122 
<< pdiffusion >>
rect 102 121 103 122 
<< pdiffusion >>
rect 103 121 104 122 
<< pdiffusion >>
rect 104 121 105 122 
<< pdiffusion >>
rect 105 121 106 122 
<< pdiffusion >>
rect 106 121 107 122 
<< pdiffusion >>
rect 107 121 108 122 
<< m1 >>
rect 109 121 110 122 
<< m2 >>
rect 110 121 111 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< m1 >>
rect 130 121 131 122 
<< m1 >>
rect 132 121 133 122 
<< m1 >>
rect 136 121 137 122 
<< m2 >>
rect 136 121 137 122 
<< pdiffusion >>
rect 138 121 139 122 
<< pdiffusion >>
rect 139 121 140 122 
<< pdiffusion >>
rect 140 121 141 122 
<< pdiffusion >>
rect 141 121 142 122 
<< pdiffusion >>
rect 142 121 143 122 
<< pdiffusion >>
rect 143 121 144 122 
<< m1 >>
rect 145 121 146 122 
<< m2 >>
rect 145 121 146 122 
<< m1 >>
rect 147 121 148 122 
<< m1 >>
rect 154 121 155 122 
<< pdiffusion >>
rect 156 121 157 122 
<< pdiffusion >>
rect 157 121 158 122 
<< pdiffusion >>
rect 158 121 159 122 
<< pdiffusion >>
rect 159 121 160 122 
<< pdiffusion >>
rect 160 121 161 122 
<< pdiffusion >>
rect 161 121 162 122 
<< m1 >>
rect 163 121 164 122 
<< m2 >>
rect 164 121 165 122 
<< m2 >>
rect 167 121 168 122 
<< m1 >>
rect 168 121 169 122 
<< m1 >>
rect 170 121 171 122 
<< m1 >>
rect 172 121 173 122 
<< pdiffusion >>
rect 174 121 175 122 
<< pdiffusion >>
rect 175 121 176 122 
<< pdiffusion >>
rect 176 121 177 122 
<< pdiffusion >>
rect 177 121 178 122 
<< pdiffusion >>
rect 178 121 179 122 
<< pdiffusion >>
rect 179 121 180 122 
<< m1 >>
rect 181 121 182 122 
<< pdiffusion >>
rect 192 121 193 122 
<< pdiffusion >>
rect 193 121 194 122 
<< pdiffusion >>
rect 194 121 195 122 
<< pdiffusion >>
rect 195 121 196 122 
<< pdiffusion >>
rect 196 121 197 122 
<< pdiffusion >>
rect 197 121 198 122 
<< m1 >>
rect 199 121 200 122 
<< m1 >>
rect 201 121 202 122 
<< m2 >>
rect 202 121 203 122 
<< m1 >>
rect 205 121 206 122 
<< pdiffusion >>
rect 210 121 211 122 
<< pdiffusion >>
rect 211 121 212 122 
<< pdiffusion >>
rect 212 121 213 122 
<< pdiffusion >>
rect 213 121 214 122 
<< pdiffusion >>
rect 214 121 215 122 
<< pdiffusion >>
rect 215 121 216 122 
<< m1 >>
rect 226 121 227 122 
<< m2 >>
rect 226 121 227 122 
<< pdiffusion >>
rect 228 121 229 122 
<< pdiffusion >>
rect 229 121 230 122 
<< pdiffusion >>
rect 230 121 231 122 
<< pdiffusion >>
rect 231 121 232 122 
<< pdiffusion >>
rect 232 121 233 122 
<< pdiffusion >>
rect 233 121 234 122 
<< m1 >>
rect 235 121 236 122 
<< m2 >>
rect 235 121 236 122 
<< m1 >>
rect 244 121 245 122 
<< pdiffusion >>
rect 246 121 247 122 
<< pdiffusion >>
rect 247 121 248 122 
<< pdiffusion >>
rect 248 121 249 122 
<< pdiffusion >>
rect 249 121 250 122 
<< pdiffusion >>
rect 250 121 251 122 
<< pdiffusion >>
rect 251 121 252 122 
<< m1 >>
rect 253 121 254 122 
<< m2 >>
rect 257 121 258 122 
<< m1 >>
rect 258 121 259 122 
<< m1 >>
rect 260 121 261 122 
<< m1 >>
rect 262 121 263 122 
<< pdiffusion >>
rect 264 121 265 122 
<< pdiffusion >>
rect 265 121 266 122 
<< pdiffusion >>
rect 266 121 267 122 
<< pdiffusion >>
rect 267 121 268 122 
<< pdiffusion >>
rect 268 121 269 122 
<< pdiffusion >>
rect 269 121 270 122 
<< m1 >>
rect 274 121 275 122 
<< m1 >>
rect 276 121 277 122 
<< m1 >>
rect 278 121 279 122 
<< m1 >>
rect 280 121 281 122 
<< pdiffusion >>
rect 282 121 283 122 
<< pdiffusion >>
rect 283 121 284 122 
<< pdiffusion >>
rect 284 121 285 122 
<< pdiffusion >>
rect 285 121 286 122 
<< pdiffusion >>
rect 286 121 287 122 
<< pdiffusion >>
rect 287 121 288 122 
<< m1 >>
rect 289 121 290 122 
<< m1 >>
rect 296 121 297 122 
<< m1 >>
rect 298 121 299 122 
<< pdiffusion >>
rect 300 121 301 122 
<< pdiffusion >>
rect 301 121 302 122 
<< pdiffusion >>
rect 302 121 303 122 
<< pdiffusion >>
rect 303 121 304 122 
<< pdiffusion >>
rect 304 121 305 122 
<< pdiffusion >>
rect 305 121 306 122 
<< m1 >>
rect 307 121 308 122 
<< m2 >>
rect 308 121 309 122 
<< m1 >>
rect 316 121 317 122 
<< pdiffusion >>
rect 318 121 319 122 
<< pdiffusion >>
rect 319 121 320 122 
<< pdiffusion >>
rect 320 121 321 122 
<< pdiffusion >>
rect 321 121 322 122 
<< pdiffusion >>
rect 322 121 323 122 
<< pdiffusion >>
rect 323 121 324 122 
<< m1 >>
rect 327 121 328 122 
<< m1 >>
rect 329 121 330 122 
<< m1 >>
rect 331 121 332 122 
<< pdiffusion >>
rect 336 121 337 122 
<< pdiffusion >>
rect 337 121 338 122 
<< pdiffusion >>
rect 338 121 339 122 
<< pdiffusion >>
rect 339 121 340 122 
<< pdiffusion >>
rect 340 121 341 122 
<< pdiffusion >>
rect 341 121 342 122 
<< m1 >>
rect 345 121 346 122 
<< m1 >>
rect 10 122 11 123 
<< pdiffusion >>
rect 12 122 13 123 
<< pdiffusion >>
rect 13 122 14 123 
<< pdiffusion >>
rect 14 122 15 123 
<< pdiffusion >>
rect 15 122 16 123 
<< pdiffusion >>
rect 16 122 17 123 
<< pdiffusion >>
rect 17 122 18 123 
<< m1 >>
rect 19 122 20 123 
<< m2 >>
rect 19 122 20 123 
<< m1 >>
rect 21 122 22 123 
<< m1 >>
rect 23 122 24 123 
<< m2 >>
rect 27 122 28 123 
<< m1 >>
rect 28 122 29 123 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< m1 >>
rect 37 122 38 123 
<< m1 >>
rect 42 122 43 123 
<< m1 >>
rect 46 122 47 123 
<< pdiffusion >>
rect 48 122 49 123 
<< pdiffusion >>
rect 49 122 50 123 
<< pdiffusion >>
rect 50 122 51 123 
<< pdiffusion >>
rect 51 122 52 123 
<< pdiffusion >>
rect 52 122 53 123 
<< pdiffusion >>
rect 53 122 54 123 
<< m1 >>
rect 55 122 56 123 
<< m2 >>
rect 56 122 57 123 
<< m1 >>
rect 59 122 60 123 
<< m2 >>
rect 61 122 62 123 
<< m1 >>
rect 62 122 63 123 
<< m1 >>
rect 64 122 65 123 
<< pdiffusion >>
rect 66 122 67 123 
<< pdiffusion >>
rect 67 122 68 123 
<< pdiffusion >>
rect 68 122 69 123 
<< pdiffusion >>
rect 69 122 70 123 
<< pdiffusion >>
rect 70 122 71 123 
<< pdiffusion >>
rect 71 122 72 123 
<< m1 >>
rect 73 122 74 123 
<< m1 >>
rect 78 122 79 123 
<< m2 >>
rect 81 122 82 123 
<< m1 >>
rect 82 122 83 123 
<< pdiffusion >>
rect 84 122 85 123 
<< pdiffusion >>
rect 85 122 86 123 
<< pdiffusion >>
rect 86 122 87 123 
<< pdiffusion >>
rect 87 122 88 123 
<< pdiffusion >>
rect 88 122 89 123 
<< pdiffusion >>
rect 89 122 90 123 
<< m1 >>
rect 91 122 92 123 
<< m2 >>
rect 92 122 93 123 
<< pdiffusion >>
rect 102 122 103 123 
<< pdiffusion >>
rect 103 122 104 123 
<< pdiffusion >>
rect 104 122 105 123 
<< pdiffusion >>
rect 105 122 106 123 
<< pdiffusion >>
rect 106 122 107 123 
<< pdiffusion >>
rect 107 122 108 123 
<< m1 >>
rect 109 122 110 123 
<< m2 >>
rect 110 122 111 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< m1 >>
rect 130 122 131 123 
<< m1 >>
rect 132 122 133 123 
<< m1 >>
rect 136 122 137 123 
<< m2 >>
rect 136 122 137 123 
<< pdiffusion >>
rect 138 122 139 123 
<< pdiffusion >>
rect 139 122 140 123 
<< pdiffusion >>
rect 140 122 141 123 
<< pdiffusion >>
rect 141 122 142 123 
<< pdiffusion >>
rect 142 122 143 123 
<< pdiffusion >>
rect 143 122 144 123 
<< m1 >>
rect 145 122 146 123 
<< m2 >>
rect 145 122 146 123 
<< m1 >>
rect 147 122 148 123 
<< m1 >>
rect 154 122 155 123 
<< pdiffusion >>
rect 156 122 157 123 
<< pdiffusion >>
rect 157 122 158 123 
<< pdiffusion >>
rect 158 122 159 123 
<< pdiffusion >>
rect 159 122 160 123 
<< pdiffusion >>
rect 160 122 161 123 
<< pdiffusion >>
rect 161 122 162 123 
<< m1 >>
rect 163 122 164 123 
<< m2 >>
rect 164 122 165 123 
<< m2 >>
rect 167 122 168 123 
<< m1 >>
rect 168 122 169 123 
<< m1 >>
rect 170 122 171 123 
<< m1 >>
rect 172 122 173 123 
<< pdiffusion >>
rect 174 122 175 123 
<< pdiffusion >>
rect 175 122 176 123 
<< pdiffusion >>
rect 176 122 177 123 
<< pdiffusion >>
rect 177 122 178 123 
<< pdiffusion >>
rect 178 122 179 123 
<< pdiffusion >>
rect 179 122 180 123 
<< m1 >>
rect 181 122 182 123 
<< pdiffusion >>
rect 192 122 193 123 
<< pdiffusion >>
rect 193 122 194 123 
<< pdiffusion >>
rect 194 122 195 123 
<< pdiffusion >>
rect 195 122 196 123 
<< pdiffusion >>
rect 196 122 197 123 
<< pdiffusion >>
rect 197 122 198 123 
<< m1 >>
rect 199 122 200 123 
<< m1 >>
rect 201 122 202 123 
<< m2 >>
rect 202 122 203 123 
<< m1 >>
rect 205 122 206 123 
<< pdiffusion >>
rect 210 122 211 123 
<< pdiffusion >>
rect 211 122 212 123 
<< pdiffusion >>
rect 212 122 213 123 
<< pdiffusion >>
rect 213 122 214 123 
<< pdiffusion >>
rect 214 122 215 123 
<< pdiffusion >>
rect 215 122 216 123 
<< m1 >>
rect 226 122 227 123 
<< m2 >>
rect 226 122 227 123 
<< pdiffusion >>
rect 228 122 229 123 
<< pdiffusion >>
rect 229 122 230 123 
<< pdiffusion >>
rect 230 122 231 123 
<< pdiffusion >>
rect 231 122 232 123 
<< pdiffusion >>
rect 232 122 233 123 
<< pdiffusion >>
rect 233 122 234 123 
<< m1 >>
rect 235 122 236 123 
<< m2 >>
rect 235 122 236 123 
<< m1 >>
rect 244 122 245 123 
<< pdiffusion >>
rect 246 122 247 123 
<< pdiffusion >>
rect 247 122 248 123 
<< pdiffusion >>
rect 248 122 249 123 
<< pdiffusion >>
rect 249 122 250 123 
<< pdiffusion >>
rect 250 122 251 123 
<< pdiffusion >>
rect 251 122 252 123 
<< m1 >>
rect 253 122 254 123 
<< m2 >>
rect 257 122 258 123 
<< m1 >>
rect 258 122 259 123 
<< m1 >>
rect 260 122 261 123 
<< m1 >>
rect 262 122 263 123 
<< pdiffusion >>
rect 264 122 265 123 
<< pdiffusion >>
rect 265 122 266 123 
<< pdiffusion >>
rect 266 122 267 123 
<< pdiffusion >>
rect 267 122 268 123 
<< pdiffusion >>
rect 268 122 269 123 
<< pdiffusion >>
rect 269 122 270 123 
<< m1 >>
rect 274 122 275 123 
<< m1 >>
rect 276 122 277 123 
<< m1 >>
rect 278 122 279 123 
<< m1 >>
rect 280 122 281 123 
<< pdiffusion >>
rect 282 122 283 123 
<< pdiffusion >>
rect 283 122 284 123 
<< pdiffusion >>
rect 284 122 285 123 
<< pdiffusion >>
rect 285 122 286 123 
<< pdiffusion >>
rect 286 122 287 123 
<< pdiffusion >>
rect 287 122 288 123 
<< m1 >>
rect 289 122 290 123 
<< m1 >>
rect 296 122 297 123 
<< m1 >>
rect 298 122 299 123 
<< pdiffusion >>
rect 300 122 301 123 
<< pdiffusion >>
rect 301 122 302 123 
<< pdiffusion >>
rect 302 122 303 123 
<< pdiffusion >>
rect 303 122 304 123 
<< pdiffusion >>
rect 304 122 305 123 
<< pdiffusion >>
rect 305 122 306 123 
<< m1 >>
rect 307 122 308 123 
<< m2 >>
rect 308 122 309 123 
<< m1 >>
rect 316 122 317 123 
<< pdiffusion >>
rect 318 122 319 123 
<< pdiffusion >>
rect 319 122 320 123 
<< pdiffusion >>
rect 320 122 321 123 
<< pdiffusion >>
rect 321 122 322 123 
<< pdiffusion >>
rect 322 122 323 123 
<< pdiffusion >>
rect 323 122 324 123 
<< m1 >>
rect 327 122 328 123 
<< m1 >>
rect 329 122 330 123 
<< m1 >>
rect 331 122 332 123 
<< pdiffusion >>
rect 336 122 337 123 
<< pdiffusion >>
rect 337 122 338 123 
<< pdiffusion >>
rect 338 122 339 123 
<< pdiffusion >>
rect 339 122 340 123 
<< pdiffusion >>
rect 340 122 341 123 
<< pdiffusion >>
rect 341 122 342 123 
<< m1 >>
rect 345 122 346 123 
<< m1 >>
rect 10 123 11 124 
<< pdiffusion >>
rect 12 123 13 124 
<< pdiffusion >>
rect 13 123 14 124 
<< pdiffusion >>
rect 14 123 15 124 
<< pdiffusion >>
rect 15 123 16 124 
<< pdiffusion >>
rect 16 123 17 124 
<< pdiffusion >>
rect 17 123 18 124 
<< m1 >>
rect 19 123 20 124 
<< m2 >>
rect 19 123 20 124 
<< m1 >>
rect 21 123 22 124 
<< m1 >>
rect 23 123 24 124 
<< m2 >>
rect 27 123 28 124 
<< m1 >>
rect 28 123 29 124 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< m1 >>
rect 37 123 38 124 
<< m1 >>
rect 42 123 43 124 
<< m1 >>
rect 46 123 47 124 
<< pdiffusion >>
rect 48 123 49 124 
<< pdiffusion >>
rect 49 123 50 124 
<< pdiffusion >>
rect 50 123 51 124 
<< pdiffusion >>
rect 51 123 52 124 
<< pdiffusion >>
rect 52 123 53 124 
<< pdiffusion >>
rect 53 123 54 124 
<< m1 >>
rect 55 123 56 124 
<< m2 >>
rect 56 123 57 124 
<< m1 >>
rect 59 123 60 124 
<< m2 >>
rect 61 123 62 124 
<< m1 >>
rect 62 123 63 124 
<< m1 >>
rect 64 123 65 124 
<< pdiffusion >>
rect 66 123 67 124 
<< pdiffusion >>
rect 67 123 68 124 
<< pdiffusion >>
rect 68 123 69 124 
<< pdiffusion >>
rect 69 123 70 124 
<< pdiffusion >>
rect 70 123 71 124 
<< pdiffusion >>
rect 71 123 72 124 
<< m1 >>
rect 73 123 74 124 
<< m1 >>
rect 78 123 79 124 
<< m2 >>
rect 81 123 82 124 
<< m1 >>
rect 82 123 83 124 
<< pdiffusion >>
rect 84 123 85 124 
<< pdiffusion >>
rect 85 123 86 124 
<< pdiffusion >>
rect 86 123 87 124 
<< pdiffusion >>
rect 87 123 88 124 
<< pdiffusion >>
rect 88 123 89 124 
<< pdiffusion >>
rect 89 123 90 124 
<< m1 >>
rect 91 123 92 124 
<< m2 >>
rect 92 123 93 124 
<< pdiffusion >>
rect 102 123 103 124 
<< pdiffusion >>
rect 103 123 104 124 
<< pdiffusion >>
rect 104 123 105 124 
<< pdiffusion >>
rect 105 123 106 124 
<< pdiffusion >>
rect 106 123 107 124 
<< pdiffusion >>
rect 107 123 108 124 
<< m1 >>
rect 109 123 110 124 
<< m2 >>
rect 110 123 111 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< m1 >>
rect 130 123 131 124 
<< m1 >>
rect 132 123 133 124 
<< m1 >>
rect 136 123 137 124 
<< m2 >>
rect 136 123 137 124 
<< pdiffusion >>
rect 138 123 139 124 
<< pdiffusion >>
rect 139 123 140 124 
<< pdiffusion >>
rect 140 123 141 124 
<< pdiffusion >>
rect 141 123 142 124 
<< pdiffusion >>
rect 142 123 143 124 
<< pdiffusion >>
rect 143 123 144 124 
<< m1 >>
rect 145 123 146 124 
<< m2 >>
rect 145 123 146 124 
<< m1 >>
rect 147 123 148 124 
<< m1 >>
rect 154 123 155 124 
<< pdiffusion >>
rect 156 123 157 124 
<< pdiffusion >>
rect 157 123 158 124 
<< pdiffusion >>
rect 158 123 159 124 
<< pdiffusion >>
rect 159 123 160 124 
<< pdiffusion >>
rect 160 123 161 124 
<< pdiffusion >>
rect 161 123 162 124 
<< m1 >>
rect 163 123 164 124 
<< m2 >>
rect 164 123 165 124 
<< m2 >>
rect 167 123 168 124 
<< m1 >>
rect 168 123 169 124 
<< m1 >>
rect 170 123 171 124 
<< m1 >>
rect 172 123 173 124 
<< pdiffusion >>
rect 174 123 175 124 
<< pdiffusion >>
rect 175 123 176 124 
<< pdiffusion >>
rect 176 123 177 124 
<< pdiffusion >>
rect 177 123 178 124 
<< pdiffusion >>
rect 178 123 179 124 
<< pdiffusion >>
rect 179 123 180 124 
<< m1 >>
rect 181 123 182 124 
<< pdiffusion >>
rect 192 123 193 124 
<< pdiffusion >>
rect 193 123 194 124 
<< pdiffusion >>
rect 194 123 195 124 
<< pdiffusion >>
rect 195 123 196 124 
<< pdiffusion >>
rect 196 123 197 124 
<< pdiffusion >>
rect 197 123 198 124 
<< m1 >>
rect 199 123 200 124 
<< m1 >>
rect 201 123 202 124 
<< m2 >>
rect 202 123 203 124 
<< m1 >>
rect 205 123 206 124 
<< pdiffusion >>
rect 210 123 211 124 
<< pdiffusion >>
rect 211 123 212 124 
<< pdiffusion >>
rect 212 123 213 124 
<< pdiffusion >>
rect 213 123 214 124 
<< pdiffusion >>
rect 214 123 215 124 
<< pdiffusion >>
rect 215 123 216 124 
<< m1 >>
rect 226 123 227 124 
<< m2 >>
rect 226 123 227 124 
<< pdiffusion >>
rect 228 123 229 124 
<< pdiffusion >>
rect 229 123 230 124 
<< pdiffusion >>
rect 230 123 231 124 
<< pdiffusion >>
rect 231 123 232 124 
<< pdiffusion >>
rect 232 123 233 124 
<< pdiffusion >>
rect 233 123 234 124 
<< m1 >>
rect 235 123 236 124 
<< m2 >>
rect 235 123 236 124 
<< m1 >>
rect 244 123 245 124 
<< pdiffusion >>
rect 246 123 247 124 
<< pdiffusion >>
rect 247 123 248 124 
<< pdiffusion >>
rect 248 123 249 124 
<< pdiffusion >>
rect 249 123 250 124 
<< pdiffusion >>
rect 250 123 251 124 
<< pdiffusion >>
rect 251 123 252 124 
<< m1 >>
rect 253 123 254 124 
<< m2 >>
rect 257 123 258 124 
<< m1 >>
rect 258 123 259 124 
<< m1 >>
rect 260 123 261 124 
<< m1 >>
rect 262 123 263 124 
<< pdiffusion >>
rect 264 123 265 124 
<< pdiffusion >>
rect 265 123 266 124 
<< pdiffusion >>
rect 266 123 267 124 
<< pdiffusion >>
rect 267 123 268 124 
<< pdiffusion >>
rect 268 123 269 124 
<< pdiffusion >>
rect 269 123 270 124 
<< m1 >>
rect 274 123 275 124 
<< m1 >>
rect 276 123 277 124 
<< m1 >>
rect 278 123 279 124 
<< m1 >>
rect 280 123 281 124 
<< pdiffusion >>
rect 282 123 283 124 
<< pdiffusion >>
rect 283 123 284 124 
<< pdiffusion >>
rect 284 123 285 124 
<< pdiffusion >>
rect 285 123 286 124 
<< pdiffusion >>
rect 286 123 287 124 
<< pdiffusion >>
rect 287 123 288 124 
<< m1 >>
rect 289 123 290 124 
<< m1 >>
rect 296 123 297 124 
<< m1 >>
rect 298 123 299 124 
<< pdiffusion >>
rect 300 123 301 124 
<< pdiffusion >>
rect 301 123 302 124 
<< pdiffusion >>
rect 302 123 303 124 
<< pdiffusion >>
rect 303 123 304 124 
<< pdiffusion >>
rect 304 123 305 124 
<< pdiffusion >>
rect 305 123 306 124 
<< m1 >>
rect 307 123 308 124 
<< m2 >>
rect 308 123 309 124 
<< m1 >>
rect 316 123 317 124 
<< pdiffusion >>
rect 318 123 319 124 
<< pdiffusion >>
rect 319 123 320 124 
<< pdiffusion >>
rect 320 123 321 124 
<< pdiffusion >>
rect 321 123 322 124 
<< pdiffusion >>
rect 322 123 323 124 
<< pdiffusion >>
rect 323 123 324 124 
<< m1 >>
rect 327 123 328 124 
<< m1 >>
rect 329 123 330 124 
<< m1 >>
rect 331 123 332 124 
<< pdiffusion >>
rect 336 123 337 124 
<< pdiffusion >>
rect 337 123 338 124 
<< pdiffusion >>
rect 338 123 339 124 
<< pdiffusion >>
rect 339 123 340 124 
<< pdiffusion >>
rect 340 123 341 124 
<< pdiffusion >>
rect 341 123 342 124 
<< m1 >>
rect 345 123 346 124 
<< m1 >>
rect 10 124 11 125 
<< pdiffusion >>
rect 12 124 13 125 
<< pdiffusion >>
rect 13 124 14 125 
<< pdiffusion >>
rect 14 124 15 125 
<< pdiffusion >>
rect 15 124 16 125 
<< pdiffusion >>
rect 16 124 17 125 
<< pdiffusion >>
rect 17 124 18 125 
<< m1 >>
rect 19 124 20 125 
<< m2 >>
rect 19 124 20 125 
<< m1 >>
rect 21 124 22 125 
<< m1 >>
rect 23 124 24 125 
<< m2 >>
rect 27 124 28 125 
<< m1 >>
rect 28 124 29 125 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< m1 >>
rect 37 124 38 125 
<< m1 >>
rect 42 124 43 125 
<< m1 >>
rect 46 124 47 125 
<< pdiffusion >>
rect 48 124 49 125 
<< pdiffusion >>
rect 49 124 50 125 
<< pdiffusion >>
rect 50 124 51 125 
<< pdiffusion >>
rect 51 124 52 125 
<< pdiffusion >>
rect 52 124 53 125 
<< pdiffusion >>
rect 53 124 54 125 
<< m1 >>
rect 55 124 56 125 
<< m2 >>
rect 56 124 57 125 
<< m1 >>
rect 59 124 60 125 
<< m2 >>
rect 61 124 62 125 
<< m1 >>
rect 62 124 63 125 
<< m1 >>
rect 64 124 65 125 
<< pdiffusion >>
rect 66 124 67 125 
<< pdiffusion >>
rect 67 124 68 125 
<< pdiffusion >>
rect 68 124 69 125 
<< pdiffusion >>
rect 69 124 70 125 
<< pdiffusion >>
rect 70 124 71 125 
<< pdiffusion >>
rect 71 124 72 125 
<< m1 >>
rect 73 124 74 125 
<< m1 >>
rect 78 124 79 125 
<< m2 >>
rect 81 124 82 125 
<< m1 >>
rect 82 124 83 125 
<< pdiffusion >>
rect 84 124 85 125 
<< pdiffusion >>
rect 85 124 86 125 
<< pdiffusion >>
rect 86 124 87 125 
<< pdiffusion >>
rect 87 124 88 125 
<< pdiffusion >>
rect 88 124 89 125 
<< pdiffusion >>
rect 89 124 90 125 
<< m1 >>
rect 91 124 92 125 
<< m2 >>
rect 92 124 93 125 
<< pdiffusion >>
rect 102 124 103 125 
<< pdiffusion >>
rect 103 124 104 125 
<< pdiffusion >>
rect 104 124 105 125 
<< pdiffusion >>
rect 105 124 106 125 
<< pdiffusion >>
rect 106 124 107 125 
<< pdiffusion >>
rect 107 124 108 125 
<< m1 >>
rect 109 124 110 125 
<< m2 >>
rect 110 124 111 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< m1 >>
rect 130 124 131 125 
<< m1 >>
rect 132 124 133 125 
<< m1 >>
rect 136 124 137 125 
<< m2 >>
rect 136 124 137 125 
<< pdiffusion >>
rect 138 124 139 125 
<< pdiffusion >>
rect 139 124 140 125 
<< pdiffusion >>
rect 140 124 141 125 
<< pdiffusion >>
rect 141 124 142 125 
<< pdiffusion >>
rect 142 124 143 125 
<< pdiffusion >>
rect 143 124 144 125 
<< m1 >>
rect 145 124 146 125 
<< m2 >>
rect 145 124 146 125 
<< m1 >>
rect 147 124 148 125 
<< m1 >>
rect 154 124 155 125 
<< pdiffusion >>
rect 156 124 157 125 
<< pdiffusion >>
rect 157 124 158 125 
<< pdiffusion >>
rect 158 124 159 125 
<< pdiffusion >>
rect 159 124 160 125 
<< pdiffusion >>
rect 160 124 161 125 
<< pdiffusion >>
rect 161 124 162 125 
<< m1 >>
rect 163 124 164 125 
<< m2 >>
rect 164 124 165 125 
<< m2 >>
rect 167 124 168 125 
<< m1 >>
rect 168 124 169 125 
<< m1 >>
rect 170 124 171 125 
<< m1 >>
rect 172 124 173 125 
<< pdiffusion >>
rect 174 124 175 125 
<< pdiffusion >>
rect 175 124 176 125 
<< pdiffusion >>
rect 176 124 177 125 
<< pdiffusion >>
rect 177 124 178 125 
<< pdiffusion >>
rect 178 124 179 125 
<< pdiffusion >>
rect 179 124 180 125 
<< m1 >>
rect 181 124 182 125 
<< pdiffusion >>
rect 192 124 193 125 
<< pdiffusion >>
rect 193 124 194 125 
<< pdiffusion >>
rect 194 124 195 125 
<< pdiffusion >>
rect 195 124 196 125 
<< pdiffusion >>
rect 196 124 197 125 
<< pdiffusion >>
rect 197 124 198 125 
<< m1 >>
rect 199 124 200 125 
<< m1 >>
rect 201 124 202 125 
<< m2 >>
rect 202 124 203 125 
<< m1 >>
rect 205 124 206 125 
<< pdiffusion >>
rect 210 124 211 125 
<< pdiffusion >>
rect 211 124 212 125 
<< pdiffusion >>
rect 212 124 213 125 
<< pdiffusion >>
rect 213 124 214 125 
<< pdiffusion >>
rect 214 124 215 125 
<< pdiffusion >>
rect 215 124 216 125 
<< m1 >>
rect 226 124 227 125 
<< m2 >>
rect 226 124 227 125 
<< pdiffusion >>
rect 228 124 229 125 
<< pdiffusion >>
rect 229 124 230 125 
<< pdiffusion >>
rect 230 124 231 125 
<< pdiffusion >>
rect 231 124 232 125 
<< pdiffusion >>
rect 232 124 233 125 
<< pdiffusion >>
rect 233 124 234 125 
<< m1 >>
rect 235 124 236 125 
<< m2 >>
rect 235 124 236 125 
<< m1 >>
rect 244 124 245 125 
<< pdiffusion >>
rect 246 124 247 125 
<< pdiffusion >>
rect 247 124 248 125 
<< pdiffusion >>
rect 248 124 249 125 
<< pdiffusion >>
rect 249 124 250 125 
<< pdiffusion >>
rect 250 124 251 125 
<< pdiffusion >>
rect 251 124 252 125 
<< m1 >>
rect 253 124 254 125 
<< m2 >>
rect 257 124 258 125 
<< m1 >>
rect 258 124 259 125 
<< m1 >>
rect 260 124 261 125 
<< m1 >>
rect 262 124 263 125 
<< pdiffusion >>
rect 264 124 265 125 
<< pdiffusion >>
rect 265 124 266 125 
<< pdiffusion >>
rect 266 124 267 125 
<< pdiffusion >>
rect 267 124 268 125 
<< pdiffusion >>
rect 268 124 269 125 
<< pdiffusion >>
rect 269 124 270 125 
<< m1 >>
rect 274 124 275 125 
<< m1 >>
rect 276 124 277 125 
<< m1 >>
rect 278 124 279 125 
<< m1 >>
rect 280 124 281 125 
<< pdiffusion >>
rect 282 124 283 125 
<< pdiffusion >>
rect 283 124 284 125 
<< pdiffusion >>
rect 284 124 285 125 
<< pdiffusion >>
rect 285 124 286 125 
<< pdiffusion >>
rect 286 124 287 125 
<< pdiffusion >>
rect 287 124 288 125 
<< m1 >>
rect 289 124 290 125 
<< m1 >>
rect 296 124 297 125 
<< m1 >>
rect 298 124 299 125 
<< pdiffusion >>
rect 300 124 301 125 
<< pdiffusion >>
rect 301 124 302 125 
<< pdiffusion >>
rect 302 124 303 125 
<< pdiffusion >>
rect 303 124 304 125 
<< pdiffusion >>
rect 304 124 305 125 
<< pdiffusion >>
rect 305 124 306 125 
<< m1 >>
rect 307 124 308 125 
<< m2 >>
rect 308 124 309 125 
<< m1 >>
rect 316 124 317 125 
<< pdiffusion >>
rect 318 124 319 125 
<< pdiffusion >>
rect 319 124 320 125 
<< pdiffusion >>
rect 320 124 321 125 
<< pdiffusion >>
rect 321 124 322 125 
<< pdiffusion >>
rect 322 124 323 125 
<< pdiffusion >>
rect 323 124 324 125 
<< m1 >>
rect 327 124 328 125 
<< m1 >>
rect 329 124 330 125 
<< m1 >>
rect 331 124 332 125 
<< pdiffusion >>
rect 336 124 337 125 
<< pdiffusion >>
rect 337 124 338 125 
<< pdiffusion >>
rect 338 124 339 125 
<< pdiffusion >>
rect 339 124 340 125 
<< pdiffusion >>
rect 340 124 341 125 
<< pdiffusion >>
rect 341 124 342 125 
<< m1 >>
rect 345 124 346 125 
<< m1 >>
rect 10 125 11 126 
<< pdiffusion >>
rect 12 125 13 126 
<< pdiffusion >>
rect 13 125 14 126 
<< pdiffusion >>
rect 14 125 15 126 
<< pdiffusion >>
rect 15 125 16 126 
<< pdiffusion >>
rect 16 125 17 126 
<< pdiffusion >>
rect 17 125 18 126 
<< m1 >>
rect 19 125 20 126 
<< m2 >>
rect 19 125 20 126 
<< m1 >>
rect 21 125 22 126 
<< m1 >>
rect 23 125 24 126 
<< m2 >>
rect 27 125 28 126 
<< m1 >>
rect 28 125 29 126 
<< pdiffusion >>
rect 30 125 31 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< m1 >>
rect 37 125 38 126 
<< m1 >>
rect 42 125 43 126 
<< m1 >>
rect 46 125 47 126 
<< pdiffusion >>
rect 48 125 49 126 
<< m1 >>
rect 49 125 50 126 
<< pdiffusion >>
rect 49 125 50 126 
<< pdiffusion >>
rect 50 125 51 126 
<< pdiffusion >>
rect 51 125 52 126 
<< pdiffusion >>
rect 52 125 53 126 
<< pdiffusion >>
rect 53 125 54 126 
<< m1 >>
rect 55 125 56 126 
<< m2 >>
rect 56 125 57 126 
<< m1 >>
rect 59 125 60 126 
<< m2 >>
rect 61 125 62 126 
<< m1 >>
rect 62 125 63 126 
<< m1 >>
rect 64 125 65 126 
<< pdiffusion >>
rect 66 125 67 126 
<< pdiffusion >>
rect 67 125 68 126 
<< pdiffusion >>
rect 68 125 69 126 
<< pdiffusion >>
rect 69 125 70 126 
<< pdiffusion >>
rect 70 125 71 126 
<< pdiffusion >>
rect 71 125 72 126 
<< m1 >>
rect 73 125 74 126 
<< m1 >>
rect 78 125 79 126 
<< m2 >>
rect 81 125 82 126 
<< m1 >>
rect 82 125 83 126 
<< pdiffusion >>
rect 84 125 85 126 
<< pdiffusion >>
rect 85 125 86 126 
<< pdiffusion >>
rect 86 125 87 126 
<< pdiffusion >>
rect 87 125 88 126 
<< pdiffusion >>
rect 88 125 89 126 
<< pdiffusion >>
rect 89 125 90 126 
<< m1 >>
rect 91 125 92 126 
<< m2 >>
rect 92 125 93 126 
<< pdiffusion >>
rect 102 125 103 126 
<< pdiffusion >>
rect 103 125 104 126 
<< pdiffusion >>
rect 104 125 105 126 
<< pdiffusion >>
rect 105 125 106 126 
<< pdiffusion >>
rect 106 125 107 126 
<< pdiffusion >>
rect 107 125 108 126 
<< m1 >>
rect 109 125 110 126 
<< m2 >>
rect 110 125 111 126 
<< pdiffusion >>
rect 120 125 121 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< m1 >>
rect 130 125 131 126 
<< m1 >>
rect 132 125 133 126 
<< m1 >>
rect 136 125 137 126 
<< m2 >>
rect 136 125 137 126 
<< pdiffusion >>
rect 138 125 139 126 
<< pdiffusion >>
rect 139 125 140 126 
<< pdiffusion >>
rect 140 125 141 126 
<< pdiffusion >>
rect 141 125 142 126 
<< pdiffusion >>
rect 142 125 143 126 
<< pdiffusion >>
rect 143 125 144 126 
<< m1 >>
rect 145 125 146 126 
<< m2 >>
rect 145 125 146 126 
<< m1 >>
rect 147 125 148 126 
<< m1 >>
rect 154 125 155 126 
<< pdiffusion >>
rect 156 125 157 126 
<< pdiffusion >>
rect 157 125 158 126 
<< pdiffusion >>
rect 158 125 159 126 
<< pdiffusion >>
rect 159 125 160 126 
<< pdiffusion >>
rect 160 125 161 126 
<< pdiffusion >>
rect 161 125 162 126 
<< m1 >>
rect 163 125 164 126 
<< m2 >>
rect 164 125 165 126 
<< m2 >>
rect 167 125 168 126 
<< m1 >>
rect 168 125 169 126 
<< m1 >>
rect 170 125 171 126 
<< m1 >>
rect 172 125 173 126 
<< pdiffusion >>
rect 174 125 175 126 
<< pdiffusion >>
rect 175 125 176 126 
<< pdiffusion >>
rect 176 125 177 126 
<< pdiffusion >>
rect 177 125 178 126 
<< pdiffusion >>
rect 178 125 179 126 
<< pdiffusion >>
rect 179 125 180 126 
<< m1 >>
rect 181 125 182 126 
<< pdiffusion >>
rect 192 125 193 126 
<< m1 >>
rect 193 125 194 126 
<< pdiffusion >>
rect 193 125 194 126 
<< pdiffusion >>
rect 194 125 195 126 
<< pdiffusion >>
rect 195 125 196 126 
<< pdiffusion >>
rect 196 125 197 126 
<< pdiffusion >>
rect 197 125 198 126 
<< m1 >>
rect 199 125 200 126 
<< m1 >>
rect 201 125 202 126 
<< m2 >>
rect 202 125 203 126 
<< m1 >>
rect 205 125 206 126 
<< pdiffusion >>
rect 210 125 211 126 
<< m1 >>
rect 211 125 212 126 
<< pdiffusion >>
rect 211 125 212 126 
<< pdiffusion >>
rect 212 125 213 126 
<< pdiffusion >>
rect 213 125 214 126 
<< pdiffusion >>
rect 214 125 215 126 
<< pdiffusion >>
rect 215 125 216 126 
<< m1 >>
rect 226 125 227 126 
<< m2 >>
rect 226 125 227 126 
<< pdiffusion >>
rect 228 125 229 126 
<< pdiffusion >>
rect 229 125 230 126 
<< pdiffusion >>
rect 230 125 231 126 
<< pdiffusion >>
rect 231 125 232 126 
<< pdiffusion >>
rect 232 125 233 126 
<< pdiffusion >>
rect 233 125 234 126 
<< m1 >>
rect 235 125 236 126 
<< m2 >>
rect 235 125 236 126 
<< m1 >>
rect 244 125 245 126 
<< pdiffusion >>
rect 246 125 247 126 
<< m1 >>
rect 247 125 248 126 
<< pdiffusion >>
rect 247 125 248 126 
<< pdiffusion >>
rect 248 125 249 126 
<< pdiffusion >>
rect 249 125 250 126 
<< pdiffusion >>
rect 250 125 251 126 
<< pdiffusion >>
rect 251 125 252 126 
<< m1 >>
rect 253 125 254 126 
<< m2 >>
rect 257 125 258 126 
<< m1 >>
rect 258 125 259 126 
<< m1 >>
rect 260 125 261 126 
<< m1 >>
rect 262 125 263 126 
<< pdiffusion >>
rect 264 125 265 126 
<< pdiffusion >>
rect 265 125 266 126 
<< pdiffusion >>
rect 266 125 267 126 
<< pdiffusion >>
rect 267 125 268 126 
<< m1 >>
rect 268 125 269 126 
<< pdiffusion >>
rect 268 125 269 126 
<< pdiffusion >>
rect 269 125 270 126 
<< m1 >>
rect 274 125 275 126 
<< m1 >>
rect 276 125 277 126 
<< m1 >>
rect 278 125 279 126 
<< m1 >>
rect 280 125 281 126 
<< pdiffusion >>
rect 282 125 283 126 
<< m1 >>
rect 283 125 284 126 
<< pdiffusion >>
rect 283 125 284 126 
<< pdiffusion >>
rect 284 125 285 126 
<< pdiffusion >>
rect 285 125 286 126 
<< m1 >>
rect 286 125 287 126 
<< pdiffusion >>
rect 286 125 287 126 
<< pdiffusion >>
rect 287 125 288 126 
<< m1 >>
rect 289 125 290 126 
<< m1 >>
rect 296 125 297 126 
<< m1 >>
rect 298 125 299 126 
<< pdiffusion >>
rect 300 125 301 126 
<< pdiffusion >>
rect 301 125 302 126 
<< pdiffusion >>
rect 302 125 303 126 
<< pdiffusion >>
rect 303 125 304 126 
<< pdiffusion >>
rect 304 125 305 126 
<< pdiffusion >>
rect 305 125 306 126 
<< m1 >>
rect 307 125 308 126 
<< m2 >>
rect 308 125 309 126 
<< m1 >>
rect 316 125 317 126 
<< pdiffusion >>
rect 318 125 319 126 
<< m1 >>
rect 319 125 320 126 
<< pdiffusion >>
rect 319 125 320 126 
<< pdiffusion >>
rect 320 125 321 126 
<< pdiffusion >>
rect 321 125 322 126 
<< m1 >>
rect 322 125 323 126 
<< pdiffusion >>
rect 322 125 323 126 
<< pdiffusion >>
rect 323 125 324 126 
<< m1 >>
rect 327 125 328 126 
<< m1 >>
rect 329 125 330 126 
<< m1 >>
rect 331 125 332 126 
<< pdiffusion >>
rect 336 125 337 126 
<< pdiffusion >>
rect 337 125 338 126 
<< pdiffusion >>
rect 338 125 339 126 
<< pdiffusion >>
rect 339 125 340 126 
<< pdiffusion >>
rect 340 125 341 126 
<< pdiffusion >>
rect 341 125 342 126 
<< m1 >>
rect 345 125 346 126 
<< m1 >>
rect 10 126 11 127 
<< m1 >>
rect 19 126 20 127 
<< m2 >>
rect 19 126 20 127 
<< m1 >>
rect 21 126 22 127 
<< m1 >>
rect 23 126 24 127 
<< m2 >>
rect 27 126 28 127 
<< m1 >>
rect 28 126 29 127 
<< m1 >>
rect 37 126 38 127 
<< m1 >>
rect 42 126 43 127 
<< m1 >>
rect 46 126 47 127 
<< m1 >>
rect 49 126 50 127 
<< m1 >>
rect 55 126 56 127 
<< m2 >>
rect 56 126 57 127 
<< m1 >>
rect 59 126 60 127 
<< m2 >>
rect 61 126 62 127 
<< m1 >>
rect 62 126 63 127 
<< m1 >>
rect 64 126 65 127 
<< m1 >>
rect 73 126 74 127 
<< m1 >>
rect 78 126 79 127 
<< m2 >>
rect 81 126 82 127 
<< m1 >>
rect 82 126 83 127 
<< m1 >>
rect 91 126 92 127 
<< m2 >>
rect 92 126 93 127 
<< m1 >>
rect 109 126 110 127 
<< m2 >>
rect 110 126 111 127 
<< m1 >>
rect 130 126 131 127 
<< m1 >>
rect 132 126 133 127 
<< m1 >>
rect 136 126 137 127 
<< m2 >>
rect 136 126 137 127 
<< m1 >>
rect 145 126 146 127 
<< m2 >>
rect 145 126 146 127 
<< m1 >>
rect 147 126 148 127 
<< m1 >>
rect 154 126 155 127 
<< m1 >>
rect 163 126 164 127 
<< m2 >>
rect 164 126 165 127 
<< m2 >>
rect 167 126 168 127 
<< m1 >>
rect 168 126 169 127 
<< m1 >>
rect 170 126 171 127 
<< m1 >>
rect 172 126 173 127 
<< m1 >>
rect 181 126 182 127 
<< m1 >>
rect 193 126 194 127 
<< m1 >>
rect 199 126 200 127 
<< m1 >>
rect 201 126 202 127 
<< m2 >>
rect 202 126 203 127 
<< m1 >>
rect 205 126 206 127 
<< m1 >>
rect 211 126 212 127 
<< m1 >>
rect 226 126 227 127 
<< m2 >>
rect 226 126 227 127 
<< m1 >>
rect 235 126 236 127 
<< m2 >>
rect 235 126 236 127 
<< m1 >>
rect 244 126 245 127 
<< m1 >>
rect 247 126 248 127 
<< m1 >>
rect 253 126 254 127 
<< m2 >>
rect 253 126 254 127 
<< m2c >>
rect 253 126 254 127 
<< m1 >>
rect 253 126 254 127 
<< m2 >>
rect 253 126 254 127 
<< m2 >>
rect 257 126 258 127 
<< m1 >>
rect 258 126 259 127 
<< m1 >>
rect 260 126 261 127 
<< m1 >>
rect 262 126 263 127 
<< m1 >>
rect 268 126 269 127 
<< m1 >>
rect 274 126 275 127 
<< m1 >>
rect 276 126 277 127 
<< m1 >>
rect 278 126 279 127 
<< m1 >>
rect 280 126 281 127 
<< m1 >>
rect 283 126 284 127 
<< m1 >>
rect 286 126 287 127 
<< m1 >>
rect 289 126 290 127 
<< m1 >>
rect 296 126 297 127 
<< m1 >>
rect 298 126 299 127 
<< m1 >>
rect 307 126 308 127 
<< m2 >>
rect 308 126 309 127 
<< m1 >>
rect 316 126 317 127 
<< m1 >>
rect 319 126 320 127 
<< m1 >>
rect 322 126 323 127 
<< m1 >>
rect 327 126 328 127 
<< m1 >>
rect 329 126 330 127 
<< m1 >>
rect 331 126 332 127 
<< m1 >>
rect 345 126 346 127 
<< m1 >>
rect 10 127 11 128 
<< m1 >>
rect 19 127 20 128 
<< m2 >>
rect 19 127 20 128 
<< m1 >>
rect 21 127 22 128 
<< m1 >>
rect 23 127 24 128 
<< m2 >>
rect 27 127 28 128 
<< m1 >>
rect 28 127 29 128 
<< m1 >>
rect 37 127 38 128 
<< m1 >>
rect 42 127 43 128 
<< m1 >>
rect 46 127 47 128 
<< m1 >>
rect 49 127 50 128 
<< m1 >>
rect 55 127 56 128 
<< m2 >>
rect 56 127 57 128 
<< m1 >>
rect 59 127 60 128 
<< m2 >>
rect 59 127 60 128 
<< m2c >>
rect 59 127 60 128 
<< m1 >>
rect 59 127 60 128 
<< m2 >>
rect 59 127 60 128 
<< m2 >>
rect 61 127 62 128 
<< m1 >>
rect 62 127 63 128 
<< m1 >>
rect 64 127 65 128 
<< m1 >>
rect 73 127 74 128 
<< m1 >>
rect 78 127 79 128 
<< m2 >>
rect 81 127 82 128 
<< m1 >>
rect 82 127 83 128 
<< m2 >>
rect 82 127 83 128 
<< m2 >>
rect 83 127 84 128 
<< m1 >>
rect 84 127 85 128 
<< m2 >>
rect 84 127 85 128 
<< m2c >>
rect 84 127 85 128 
<< m1 >>
rect 84 127 85 128 
<< m2 >>
rect 84 127 85 128 
<< m1 >>
rect 91 127 92 128 
<< m2 >>
rect 92 127 93 128 
<< m1 >>
rect 107 127 108 128 
<< m2 >>
rect 107 127 108 128 
<< m2c >>
rect 107 127 108 128 
<< m1 >>
rect 107 127 108 128 
<< m2 >>
rect 107 127 108 128 
<< m2 >>
rect 108 127 109 128 
<< m1 >>
rect 109 127 110 128 
<< m2 >>
rect 109 127 110 128 
<< m2 >>
rect 110 127 111 128 
<< m1 >>
rect 130 127 131 128 
<< m1 >>
rect 132 127 133 128 
<< m1 >>
rect 136 127 137 128 
<< m2 >>
rect 136 127 137 128 
<< m1 >>
rect 145 127 146 128 
<< m2 >>
rect 145 127 146 128 
<< m1 >>
rect 147 127 148 128 
<< m1 >>
rect 154 127 155 128 
<< m1 >>
rect 163 127 164 128 
<< m2 >>
rect 164 127 165 128 
<< m2 >>
rect 167 127 168 128 
<< m1 >>
rect 168 127 169 128 
<< m2 >>
rect 168 127 169 128 
<< m2 >>
rect 169 127 170 128 
<< m1 >>
rect 170 127 171 128 
<< m2 >>
rect 170 127 171 128 
<< m2 >>
rect 171 127 172 128 
<< m1 >>
rect 172 127 173 128 
<< m2 >>
rect 172 127 173 128 
<< m2 >>
rect 173 127 174 128 
<< m1 >>
rect 174 127 175 128 
<< m2 >>
rect 174 127 175 128 
<< m2c >>
rect 174 127 175 128 
<< m1 >>
rect 174 127 175 128 
<< m2 >>
rect 174 127 175 128 
<< m1 >>
rect 181 127 182 128 
<< m1 >>
rect 193 127 194 128 
<< m1 >>
rect 197 127 198 128 
<< m2 >>
rect 197 127 198 128 
<< m2c >>
rect 197 127 198 128 
<< m1 >>
rect 197 127 198 128 
<< m2 >>
rect 197 127 198 128 
<< m2 >>
rect 198 127 199 128 
<< m1 >>
rect 199 127 200 128 
<< m2 >>
rect 199 127 200 128 
<< m2 >>
rect 200 127 201 128 
<< m1 >>
rect 201 127 202 128 
<< m2 >>
rect 201 127 202 128 
<< m2 >>
rect 202 127 203 128 
<< m1 >>
rect 205 127 206 128 
<< m2 >>
rect 205 127 206 128 
<< m2c >>
rect 205 127 206 128 
<< m1 >>
rect 205 127 206 128 
<< m2 >>
rect 205 127 206 128 
<< m1 >>
rect 211 127 212 128 
<< m1 >>
rect 226 127 227 128 
<< m2 >>
rect 226 127 227 128 
<< m1 >>
rect 235 127 236 128 
<< m2 >>
rect 235 127 236 128 
<< m1 >>
rect 244 127 245 128 
<< m1 >>
rect 247 127 248 128 
<< m2 >>
rect 251 127 252 128 
<< m2 >>
rect 252 127 253 128 
<< m2 >>
rect 253 127 254 128 
<< m2 >>
rect 257 127 258 128 
<< m1 >>
rect 258 127 259 128 
<< m1 >>
rect 260 127 261 128 
<< m1 >>
rect 262 127 263 128 
<< m1 >>
rect 268 127 269 128 
<< m1 >>
rect 274 127 275 128 
<< m1 >>
rect 276 127 277 128 
<< m1 >>
rect 278 127 279 128 
<< m1 >>
rect 280 127 281 128 
<< m1 >>
rect 283 127 284 128 
<< m1 >>
rect 286 127 287 128 
<< m1 >>
rect 289 127 290 128 
<< m1 >>
rect 296 127 297 128 
<< m1 >>
rect 298 127 299 128 
<< m1 >>
rect 307 127 308 128 
<< m2 >>
rect 308 127 309 128 
<< m1 >>
rect 316 127 317 128 
<< m1 >>
rect 317 127 318 128 
<< m1 >>
rect 318 127 319 128 
<< m1 >>
rect 319 127 320 128 
<< m1 >>
rect 322 127 323 128 
<< m1 >>
rect 323 127 324 128 
<< m1 >>
rect 324 127 325 128 
<< m1 >>
rect 325 127 326 128 
<< m1 >>
rect 327 127 328 128 
<< m1 >>
rect 329 127 330 128 
<< m1 >>
rect 331 127 332 128 
<< m1 >>
rect 345 127 346 128 
<< m1 >>
rect 10 128 11 129 
<< m1 >>
rect 19 128 20 129 
<< m2 >>
rect 19 128 20 129 
<< m1 >>
rect 21 128 22 129 
<< m1 >>
rect 23 128 24 129 
<< m2 >>
rect 27 128 28 129 
<< m1 >>
rect 28 128 29 129 
<< m1 >>
rect 37 128 38 129 
<< m1 >>
rect 42 128 43 129 
<< m1 >>
rect 46 128 47 129 
<< m1 >>
rect 49 128 50 129 
<< m1 >>
rect 50 128 51 129 
<< m1 >>
rect 51 128 52 129 
<< m1 >>
rect 52 128 53 129 
<< m1 >>
rect 53 128 54 129 
<< m1 >>
rect 54 128 55 129 
<< m1 >>
rect 55 128 56 129 
<< m2 >>
rect 56 128 57 129 
<< m2 >>
rect 59 128 60 129 
<< m2 >>
rect 61 128 62 129 
<< m1 >>
rect 62 128 63 129 
<< m1 >>
rect 64 128 65 129 
<< m1 >>
rect 73 128 74 129 
<< m1 >>
rect 78 128 79 129 
<< m1 >>
rect 82 128 83 129 
<< m1 >>
rect 84 128 85 129 
<< m1 >>
rect 91 128 92 129 
<< m2 >>
rect 92 128 93 129 
<< m1 >>
rect 106 128 107 129 
<< m1 >>
rect 107 128 108 129 
<< m1 >>
rect 109 128 110 129 
<< m1 >>
rect 130 128 131 129 
<< m1 >>
rect 132 128 133 129 
<< m1 >>
rect 136 128 137 129 
<< m2 >>
rect 136 128 137 129 
<< m1 >>
rect 145 128 146 129 
<< m2 >>
rect 145 128 146 129 
<< m1 >>
rect 147 128 148 129 
<< m1 >>
rect 154 128 155 129 
<< m1 >>
rect 163 128 164 129 
<< m2 >>
rect 164 128 165 129 
<< m1 >>
rect 168 128 169 129 
<< m1 >>
rect 170 128 171 129 
<< m1 >>
rect 172 128 173 129 
<< m1 >>
rect 174 128 175 129 
<< m1 >>
rect 181 128 182 129 
<< m1 >>
rect 193 128 194 129 
<< m1 >>
rect 194 128 195 129 
<< m1 >>
rect 195 128 196 129 
<< m1 >>
rect 196 128 197 129 
<< m1 >>
rect 197 128 198 129 
<< m1 >>
rect 199 128 200 129 
<< m1 >>
rect 201 128 202 129 
<< m2 >>
rect 205 128 206 129 
<< m1 >>
rect 211 128 212 129 
<< m1 >>
rect 226 128 227 129 
<< m2 >>
rect 226 128 227 129 
<< m1 >>
rect 235 128 236 129 
<< m2 >>
rect 235 128 236 129 
<< m1 >>
rect 244 128 245 129 
<< m1 >>
rect 247 128 248 129 
<< m1 >>
rect 248 128 249 129 
<< m1 >>
rect 249 128 250 129 
<< m1 >>
rect 250 128 251 129 
<< m1 >>
rect 251 128 252 129 
<< m2 >>
rect 251 128 252 129 
<< m1 >>
rect 252 128 253 129 
<< m1 >>
rect 253 128 254 129 
<< m1 >>
rect 254 128 255 129 
<< m1 >>
rect 255 128 256 129 
<< m2 >>
rect 255 128 256 129 
<< m1 >>
rect 256 128 257 129 
<< m2 >>
rect 256 128 257 129 
<< m1 >>
rect 257 128 258 129 
<< m2 >>
rect 257 128 258 129 
<< m1 >>
rect 258 128 259 129 
<< m1 >>
rect 260 128 261 129 
<< m1 >>
rect 262 128 263 129 
<< m1 >>
rect 268 128 269 129 
<< m1 >>
rect 274 128 275 129 
<< m1 >>
rect 276 128 277 129 
<< m1 >>
rect 278 128 279 129 
<< m1 >>
rect 280 128 281 129 
<< m1 >>
rect 283 128 284 129 
<< m1 >>
rect 286 128 287 129 
<< m1 >>
rect 289 128 290 129 
<< m1 >>
rect 296 128 297 129 
<< m1 >>
rect 298 128 299 129 
<< m1 >>
rect 307 128 308 129 
<< m2 >>
rect 308 128 309 129 
<< m1 >>
rect 325 128 326 129 
<< m1 >>
rect 327 128 328 129 
<< m1 >>
rect 329 128 330 129 
<< m1 >>
rect 331 128 332 129 
<< m1 >>
rect 345 128 346 129 
<< m1 >>
rect 10 129 11 130 
<< m1 >>
rect 19 129 20 130 
<< m2 >>
rect 19 129 20 130 
<< m1 >>
rect 21 129 22 130 
<< m1 >>
rect 23 129 24 130 
<< m2 >>
rect 27 129 28 130 
<< m1 >>
rect 28 129 29 130 
<< m1 >>
rect 37 129 38 130 
<< m1 >>
rect 42 129 43 130 
<< m1 >>
rect 46 129 47 130 
<< m2 >>
rect 56 129 57 130 
<< m1 >>
rect 57 129 58 130 
<< m2 >>
rect 57 129 58 130 
<< m2c >>
rect 57 129 58 130 
<< m1 >>
rect 57 129 58 130 
<< m2 >>
rect 57 129 58 130 
<< m1 >>
rect 58 129 59 130 
<< m2 >>
rect 59 129 60 130 
<< m2 >>
rect 61 129 62 130 
<< m1 >>
rect 62 129 63 130 
<< m1 >>
rect 64 129 65 130 
<< m1 >>
rect 73 129 74 130 
<< m1 >>
rect 78 129 79 130 
<< m1 >>
rect 82 129 83 130 
<< m1 >>
rect 84 129 85 130 
<< m1 >>
rect 91 129 92 130 
<< m2 >>
rect 92 129 93 130 
<< m1 >>
rect 106 129 107 130 
<< m1 >>
rect 109 129 110 130 
<< m1 >>
rect 130 129 131 130 
<< m1 >>
rect 132 129 133 130 
<< m1 >>
rect 136 129 137 130 
<< m2 >>
rect 136 129 137 130 
<< m1 >>
rect 145 129 146 130 
<< m2 >>
rect 145 129 146 130 
<< m1 >>
rect 147 129 148 130 
<< m1 >>
rect 154 129 155 130 
<< m1 >>
rect 163 129 164 130 
<< m2 >>
rect 164 129 165 130 
<< m1 >>
rect 168 129 169 130 
<< m1 >>
rect 170 129 171 130 
<< m1 >>
rect 172 129 173 130 
<< m1 >>
rect 174 129 175 130 
<< m1 >>
rect 181 129 182 130 
<< m1 >>
rect 199 129 200 130 
<< m1 >>
rect 201 129 202 130 
<< m2 >>
rect 202 129 203 130 
<< m1 >>
rect 203 129 204 130 
<< m2 >>
rect 203 129 204 130 
<< m2c >>
rect 203 129 204 130 
<< m1 >>
rect 203 129 204 130 
<< m2 >>
rect 203 129 204 130 
<< m1 >>
rect 204 129 205 130 
<< m1 >>
rect 205 129 206 130 
<< m2 >>
rect 205 129 206 130 
<< m1 >>
rect 206 129 207 130 
<< m1 >>
rect 207 129 208 130 
<< m1 >>
rect 208 129 209 130 
<< m1 >>
rect 209 129 210 130 
<< m1 >>
rect 210 129 211 130 
<< m1 >>
rect 211 129 212 130 
<< m1 >>
rect 226 129 227 130 
<< m2 >>
rect 226 129 227 130 
<< m1 >>
rect 235 129 236 130 
<< m2 >>
rect 235 129 236 130 
<< m1 >>
rect 244 129 245 130 
<< m2 >>
rect 251 129 252 130 
<< m2 >>
rect 255 129 256 130 
<< m2 >>
rect 258 129 259 130 
<< m2 >>
rect 259 129 260 130 
<< m1 >>
rect 260 129 261 130 
<< m2 >>
rect 260 129 261 130 
<< m2 >>
rect 261 129 262 130 
<< m1 >>
rect 262 129 263 130 
<< m2 >>
rect 262 129 263 130 
<< m2 >>
rect 263 129 264 130 
<< m1 >>
rect 264 129 265 130 
<< m2 >>
rect 264 129 265 130 
<< m2c >>
rect 264 129 265 130 
<< m1 >>
rect 264 129 265 130 
<< m2 >>
rect 264 129 265 130 
<< m1 >>
rect 266 129 267 130 
<< m2 >>
rect 266 129 267 130 
<< m2c >>
rect 266 129 267 130 
<< m1 >>
rect 266 129 267 130 
<< m2 >>
rect 266 129 267 130 
<< m1 >>
rect 267 129 268 130 
<< m1 >>
rect 268 129 269 130 
<< m2 >>
rect 268 129 269 130 
<< m2 >>
rect 269 129 270 130 
<< m1 >>
rect 270 129 271 130 
<< m2 >>
rect 270 129 271 130 
<< m2c >>
rect 270 129 271 130 
<< m1 >>
rect 270 129 271 130 
<< m2 >>
rect 270 129 271 130 
<< m1 >>
rect 271 129 272 130 
<< m1 >>
rect 272 129 273 130 
<< m2 >>
rect 272 129 273 130 
<< m2c >>
rect 272 129 273 130 
<< m1 >>
rect 272 129 273 130 
<< m2 >>
rect 272 129 273 130 
<< m2 >>
rect 273 129 274 130 
<< m1 >>
rect 274 129 275 130 
<< m2 >>
rect 274 129 275 130 
<< m2 >>
rect 275 129 276 130 
<< m1 >>
rect 276 129 277 130 
<< m2 >>
rect 276 129 277 130 
<< m2 >>
rect 277 129 278 130 
<< m1 >>
rect 278 129 279 130 
<< m2 >>
rect 278 129 279 130 
<< m2 >>
rect 279 129 280 130 
<< m1 >>
rect 280 129 281 130 
<< m2 >>
rect 280 129 281 130 
<< m2c >>
rect 280 129 281 130 
<< m1 >>
rect 280 129 281 130 
<< m2 >>
rect 280 129 281 130 
<< m1 >>
rect 283 129 284 130 
<< m1 >>
rect 286 129 287 130 
<< m1 >>
rect 289 129 290 130 
<< m1 >>
rect 296 129 297 130 
<< m1 >>
rect 298 129 299 130 
<< m1 >>
rect 307 129 308 130 
<< m2 >>
rect 308 129 309 130 
<< m1 >>
rect 325 129 326 130 
<< m1 >>
rect 327 129 328 130 
<< m1 >>
rect 329 129 330 130 
<< m1 >>
rect 331 129 332 130 
<< m1 >>
rect 345 129 346 130 
<< m1 >>
rect 10 130 11 131 
<< m1 >>
rect 19 130 20 131 
<< m2 >>
rect 19 130 20 131 
<< m1 >>
rect 21 130 22 131 
<< m1 >>
rect 23 130 24 131 
<< m2 >>
rect 27 130 28 131 
<< m1 >>
rect 28 130 29 131 
<< m1 >>
rect 37 130 38 131 
<< m1 >>
rect 42 130 43 131 
<< m1 >>
rect 46 130 47 131 
<< m1 >>
rect 58 130 59 131 
<< m2 >>
rect 59 130 60 131 
<< m2 >>
rect 61 130 62 131 
<< m1 >>
rect 62 130 63 131 
<< m1 >>
rect 64 130 65 131 
<< m1 >>
rect 73 130 74 131 
<< m1 >>
rect 78 130 79 131 
<< m1 >>
rect 82 130 83 131 
<< m1 >>
rect 84 130 85 131 
<< m1 >>
rect 85 130 86 131 
<< m1 >>
rect 91 130 92 131 
<< m2 >>
rect 92 130 93 131 
<< m1 >>
rect 106 130 107 131 
<< m1 >>
rect 109 130 110 131 
<< m1 >>
rect 130 130 131 131 
<< m1 >>
rect 132 130 133 131 
<< m1 >>
rect 136 130 137 131 
<< m2 >>
rect 136 130 137 131 
<< m1 >>
rect 145 130 146 131 
<< m2 >>
rect 145 130 146 131 
<< m1 >>
rect 147 130 148 131 
<< m1 >>
rect 154 130 155 131 
<< m1 >>
rect 163 130 164 131 
<< m2 >>
rect 164 130 165 131 
<< m1 >>
rect 168 130 169 131 
<< m1 >>
rect 170 130 171 131 
<< m1 >>
rect 172 130 173 131 
<< m1 >>
rect 174 130 175 131 
<< m1 >>
rect 175 130 176 131 
<< m1 >>
rect 176 130 177 131 
<< m1 >>
rect 181 130 182 131 
<< m1 >>
rect 182 130 183 131 
<< m1 >>
rect 183 130 184 131 
<< m1 >>
rect 184 130 185 131 
<< m1 >>
rect 185 130 186 131 
<< m1 >>
rect 186 130 187 131 
<< m1 >>
rect 187 130 188 131 
<< m1 >>
rect 188 130 189 131 
<< m1 >>
rect 189 130 190 131 
<< m1 >>
rect 190 130 191 131 
<< m1 >>
rect 191 130 192 131 
<< m1 >>
rect 192 130 193 131 
<< m2 >>
rect 192 130 193 131 
<< m2c >>
rect 192 130 193 131 
<< m1 >>
rect 192 130 193 131 
<< m2 >>
rect 192 130 193 131 
<< m1 >>
rect 197 130 198 131 
<< m2 >>
rect 197 130 198 131 
<< m2c >>
rect 197 130 198 131 
<< m1 >>
rect 197 130 198 131 
<< m2 >>
rect 197 130 198 131 
<< m2 >>
rect 198 130 199 131 
<< m1 >>
rect 199 130 200 131 
<< m2 >>
rect 199 130 200 131 
<< m2 >>
rect 200 130 201 131 
<< m1 >>
rect 201 130 202 131 
<< m2 >>
rect 201 130 202 131 
<< m2 >>
rect 202 130 203 131 
<< m2 >>
rect 205 130 206 131 
<< m1 >>
rect 226 130 227 131 
<< m2 >>
rect 226 130 227 131 
<< m1 >>
rect 235 130 236 131 
<< m2 >>
rect 235 130 236 131 
<< m1 >>
rect 244 130 245 131 
<< m2 >>
rect 251 130 252 131 
<< m1 >>
rect 255 130 256 131 
<< m2 >>
rect 255 130 256 131 
<< m1 >>
rect 258 130 259 131 
<< m2 >>
rect 258 130 259 131 
<< m1 >>
rect 260 130 261 131 
<< m1 >>
rect 262 130 263 131 
<< m2 >>
rect 264 130 265 131 
<< m2 >>
rect 265 130 266 131 
<< m2 >>
rect 266 130 267 131 
<< m2 >>
rect 268 130 269 131 
<< m1 >>
rect 274 130 275 131 
<< m1 >>
rect 276 130 277 131 
<< m1 >>
rect 278 130 279 131 
<< m1 >>
rect 283 130 284 131 
<< m1 >>
rect 286 130 287 131 
<< m1 >>
rect 289 130 290 131 
<< m1 >>
rect 296 130 297 131 
<< m1 >>
rect 298 130 299 131 
<< m1 >>
rect 307 130 308 131 
<< m2 >>
rect 308 130 309 131 
<< m1 >>
rect 325 130 326 131 
<< m1 >>
rect 327 130 328 131 
<< m1 >>
rect 329 130 330 131 
<< m1 >>
rect 331 130 332 131 
<< m1 >>
rect 332 130 333 131 
<< m1 >>
rect 333 130 334 131 
<< m1 >>
rect 334 130 335 131 
<< m1 >>
rect 335 130 336 131 
<< m1 >>
rect 336 130 337 131 
<< m1 >>
rect 337 130 338 131 
<< m1 >>
rect 338 130 339 131 
<< m1 >>
rect 345 130 346 131 
<< m1 >>
rect 10 131 11 132 
<< m1 >>
rect 19 131 20 132 
<< m2 >>
rect 19 131 20 132 
<< m1 >>
rect 21 131 22 132 
<< m1 >>
rect 23 131 24 132 
<< m2 >>
rect 27 131 28 132 
<< m1 >>
rect 28 131 29 132 
<< m1 >>
rect 37 131 38 132 
<< m1 >>
rect 42 131 43 132 
<< m1 >>
rect 46 131 47 132 
<< m1 >>
rect 58 131 59 132 
<< m2 >>
rect 59 131 60 132 
<< m2 >>
rect 61 131 62 132 
<< m1 >>
rect 62 131 63 132 
<< m1 >>
rect 64 131 65 132 
<< m1 >>
rect 73 131 74 132 
<< m1 >>
rect 78 131 79 132 
<< m1 >>
rect 82 131 83 132 
<< m1 >>
rect 85 131 86 132 
<< m1 >>
rect 91 131 92 132 
<< m2 >>
rect 92 131 93 132 
<< m1 >>
rect 106 131 107 132 
<< m1 >>
rect 109 131 110 132 
<< m1 >>
rect 130 131 131 132 
<< m1 >>
rect 132 131 133 132 
<< m1 >>
rect 136 131 137 132 
<< m2 >>
rect 136 131 137 132 
<< m1 >>
rect 145 131 146 132 
<< m2 >>
rect 145 131 146 132 
<< m1 >>
rect 147 131 148 132 
<< m1 >>
rect 154 131 155 132 
<< m1 >>
rect 163 131 164 132 
<< m2 >>
rect 164 131 165 132 
<< m1 >>
rect 168 131 169 132 
<< m1 >>
rect 170 131 171 132 
<< m1 >>
rect 172 131 173 132 
<< m1 >>
rect 176 131 177 132 
<< m2 >>
rect 176 131 177 132 
<< m2c >>
rect 176 131 177 132 
<< m1 >>
rect 176 131 177 132 
<< m2 >>
rect 176 131 177 132 
<< m2 >>
rect 192 131 193 132 
<< m1 >>
rect 197 131 198 132 
<< m1 >>
rect 199 131 200 132 
<< m1 >>
rect 201 131 202 132 
<< m1 >>
rect 205 131 206 132 
<< m2 >>
rect 205 131 206 132 
<< m2c >>
rect 205 131 206 132 
<< m1 >>
rect 205 131 206 132 
<< m2 >>
rect 205 131 206 132 
<< m1 >>
rect 226 131 227 132 
<< m2 >>
rect 226 131 227 132 
<< m1 >>
rect 235 131 236 132 
<< m2 >>
rect 235 131 236 132 
<< m1 >>
rect 244 131 245 132 
<< m1 >>
rect 245 131 246 132 
<< m1 >>
rect 246 131 247 132 
<< m1 >>
rect 247 131 248 132 
<< m1 >>
rect 248 131 249 132 
<< m1 >>
rect 249 131 250 132 
<< m1 >>
rect 250 131 251 132 
<< m1 >>
rect 251 131 252 132 
<< m2 >>
rect 251 131 252 132 
<< m1 >>
rect 252 131 253 132 
<< m1 >>
rect 253 131 254 132 
<< m2 >>
rect 253 131 254 132 
<< m2c >>
rect 253 131 254 132 
<< m1 >>
rect 253 131 254 132 
<< m2 >>
rect 253 131 254 132 
<< m1 >>
rect 255 131 256 132 
<< m2 >>
rect 255 131 256 132 
<< m2c >>
rect 255 131 256 132 
<< m1 >>
rect 255 131 256 132 
<< m2 >>
rect 255 131 256 132 
<< m1 >>
rect 258 131 259 132 
<< m2 >>
rect 258 131 259 132 
<< m2c >>
rect 258 131 259 132 
<< m1 >>
rect 258 131 259 132 
<< m2 >>
rect 258 131 259 132 
<< m1 >>
rect 260 131 261 132 
<< m2 >>
rect 260 131 261 132 
<< m2c >>
rect 260 131 261 132 
<< m1 >>
rect 260 131 261 132 
<< m2 >>
rect 260 131 261 132 
<< m2 >>
rect 261 131 262 132 
<< m1 >>
rect 262 131 263 132 
<< m2 >>
rect 262 131 263 132 
<< m1 >>
rect 263 131 264 132 
<< m1 >>
rect 264 131 265 132 
<< m1 >>
rect 265 131 266 132 
<< m1 >>
rect 266 131 267 132 
<< m1 >>
rect 267 131 268 132 
<< m1 >>
rect 268 131 269 132 
<< m2 >>
rect 268 131 269 132 
<< m1 >>
rect 269 131 270 132 
<< m1 >>
rect 270 131 271 132 
<< m1 >>
rect 271 131 272 132 
<< m1 >>
rect 272 131 273 132 
<< m2 >>
rect 272 131 273 132 
<< m2c >>
rect 272 131 273 132 
<< m1 >>
rect 272 131 273 132 
<< m2 >>
rect 272 131 273 132 
<< m1 >>
rect 274 131 275 132 
<< m2 >>
rect 274 131 275 132 
<< m2c >>
rect 274 131 275 132 
<< m1 >>
rect 274 131 275 132 
<< m2 >>
rect 274 131 275 132 
<< m1 >>
rect 276 131 277 132 
<< m2 >>
rect 276 131 277 132 
<< m2c >>
rect 276 131 277 132 
<< m1 >>
rect 276 131 277 132 
<< m2 >>
rect 276 131 277 132 
<< m1 >>
rect 278 131 279 132 
<< m2 >>
rect 278 131 279 132 
<< m2c >>
rect 278 131 279 132 
<< m1 >>
rect 278 131 279 132 
<< m2 >>
rect 278 131 279 132 
<< m1 >>
rect 283 131 284 132 
<< m2 >>
rect 283 131 284 132 
<< m2c >>
rect 283 131 284 132 
<< m1 >>
rect 283 131 284 132 
<< m2 >>
rect 283 131 284 132 
<< m1 >>
rect 286 131 287 132 
<< m1 >>
rect 289 131 290 132 
<< m1 >>
rect 296 131 297 132 
<< m1 >>
rect 298 131 299 132 
<< m1 >>
rect 307 131 308 132 
<< m2 >>
rect 308 131 309 132 
<< m1 >>
rect 325 131 326 132 
<< m1 >>
rect 327 131 328 132 
<< m1 >>
rect 329 131 330 132 
<< m1 >>
rect 338 131 339 132 
<< m1 >>
rect 345 131 346 132 
<< m1 >>
rect 10 132 11 133 
<< m1 >>
rect 19 132 20 133 
<< m2 >>
rect 19 132 20 133 
<< m1 >>
rect 21 132 22 133 
<< m1 >>
rect 23 132 24 133 
<< m2 >>
rect 27 132 28 133 
<< m1 >>
rect 28 132 29 133 
<< m1 >>
rect 37 132 38 133 
<< m1 >>
rect 42 132 43 133 
<< m1 >>
rect 46 132 47 133 
<< m1 >>
rect 58 132 59 133 
<< m2 >>
rect 59 132 60 133 
<< m2 >>
rect 61 132 62 133 
<< m1 >>
rect 62 132 63 133 
<< m1 >>
rect 64 132 65 133 
<< m1 >>
rect 73 132 74 133 
<< m1 >>
rect 78 132 79 133 
<< m1 >>
rect 82 132 83 133 
<< m1 >>
rect 85 132 86 133 
<< m1 >>
rect 91 132 92 133 
<< m2 >>
rect 92 132 93 133 
<< m1 >>
rect 106 132 107 133 
<< m1 >>
rect 109 132 110 133 
<< m1 >>
rect 130 132 131 133 
<< m1 >>
rect 132 132 133 133 
<< m1 >>
rect 136 132 137 133 
<< m2 >>
rect 136 132 137 133 
<< m1 >>
rect 145 132 146 133 
<< m2 >>
rect 145 132 146 133 
<< m1 >>
rect 147 132 148 133 
<< m1 >>
rect 154 132 155 133 
<< m1 >>
rect 163 132 164 133 
<< m2 >>
rect 164 132 165 133 
<< m1 >>
rect 168 132 169 133 
<< m1 >>
rect 170 132 171 133 
<< m1 >>
rect 172 132 173 133 
<< m2 >>
rect 176 132 177 133 
<< m2 >>
rect 178 132 179 133 
<< m2 >>
rect 179 132 180 133 
<< m2 >>
rect 180 132 181 133 
<< m2 >>
rect 181 132 182 133 
<< m2 >>
rect 182 132 183 133 
<< m2 >>
rect 183 132 184 133 
<< m2 >>
rect 184 132 185 133 
<< m2 >>
rect 185 132 186 133 
<< m2 >>
rect 186 132 187 133 
<< m2 >>
rect 187 132 188 133 
<< m2 >>
rect 188 132 189 133 
<< m2 >>
rect 189 132 190 133 
<< m1 >>
rect 190 132 191 133 
<< m2 >>
rect 190 132 191 133 
<< m2c >>
rect 190 132 191 133 
<< m1 >>
rect 190 132 191 133 
<< m2 >>
rect 190 132 191 133 
<< m1 >>
rect 191 132 192 133 
<< m1 >>
rect 192 132 193 133 
<< m2 >>
rect 192 132 193 133 
<< m1 >>
rect 193 132 194 133 
<< m1 >>
rect 194 132 195 133 
<< m1 >>
rect 195 132 196 133 
<< m1 >>
rect 196 132 197 133 
<< m1 >>
rect 197 132 198 133 
<< m1 >>
rect 199 132 200 133 
<< m1 >>
rect 201 132 202 133 
<< m1 >>
rect 205 132 206 133 
<< m1 >>
rect 226 132 227 133 
<< m2 >>
rect 226 132 227 133 
<< m1 >>
rect 235 132 236 133 
<< m2 >>
rect 235 132 236 133 
<< m2 >>
rect 241 132 242 133 
<< m2 >>
rect 242 132 243 133 
<< m2 >>
rect 243 132 244 133 
<< m2 >>
rect 244 132 245 133 
<< m2 >>
rect 245 132 246 133 
<< m2 >>
rect 246 132 247 133 
<< m2 >>
rect 247 132 248 133 
<< m2 >>
rect 248 132 249 133 
<< m2 >>
rect 249 132 250 133 
<< m2 >>
rect 250 132 251 133 
<< m2 >>
rect 251 132 252 133 
<< m2 >>
rect 253 132 254 133 
<< m2 >>
rect 255 132 256 133 
<< m2 >>
rect 258 132 259 133 
<< m2 >>
rect 262 132 263 133 
<< m2 >>
rect 268 132 269 133 
<< m2 >>
rect 272 132 273 133 
<< m2 >>
rect 274 132 275 133 
<< m2 >>
rect 276 132 277 133 
<< m2 >>
rect 278 132 279 133 
<< m2 >>
rect 279 132 280 133 
<< m2 >>
rect 280 132 281 133 
<< m2 >>
rect 282 132 283 133 
<< m2 >>
rect 283 132 284 133 
<< m1 >>
rect 286 132 287 133 
<< m1 >>
rect 289 132 290 133 
<< m1 >>
rect 296 132 297 133 
<< m1 >>
rect 298 132 299 133 
<< m1 >>
rect 307 132 308 133 
<< m2 >>
rect 308 132 309 133 
<< m1 >>
rect 325 132 326 133 
<< m1 >>
rect 327 132 328 133 
<< m1 >>
rect 329 132 330 133 
<< m1 >>
rect 338 132 339 133 
<< m1 >>
rect 345 132 346 133 
<< m1 >>
rect 10 133 11 134 
<< m1 >>
rect 19 133 20 134 
<< m2 >>
rect 19 133 20 134 
<< m1 >>
rect 21 133 22 134 
<< m1 >>
rect 23 133 24 134 
<< m2 >>
rect 27 133 28 134 
<< m1 >>
rect 28 133 29 134 
<< m1 >>
rect 37 133 38 134 
<< m2 >>
rect 38 133 39 134 
<< m1 >>
rect 39 133 40 134 
<< m2 >>
rect 39 133 40 134 
<< m1 >>
rect 40 133 41 134 
<< m2 >>
rect 40 133 41 134 
<< m2c >>
rect 40 133 41 134 
<< m1 >>
rect 40 133 41 134 
<< m2 >>
rect 40 133 41 134 
<< m2 >>
rect 41 133 42 134 
<< m1 >>
rect 42 133 43 134 
<< m2 >>
rect 42 133 43 134 
<< m2 >>
rect 43 133 44 134 
<< m1 >>
rect 44 133 45 134 
<< m2 >>
rect 44 133 45 134 
<< m2c >>
rect 44 133 45 134 
<< m1 >>
rect 44 133 45 134 
<< m2 >>
rect 44 133 45 134 
<< m2 >>
rect 45 133 46 134 
<< m1 >>
rect 46 133 47 134 
<< m2 >>
rect 46 133 47 134 
<< m2 >>
rect 47 133 48 134 
<< m1 >>
rect 48 133 49 134 
<< m2 >>
rect 48 133 49 134 
<< m2c >>
rect 48 133 49 134 
<< m1 >>
rect 48 133 49 134 
<< m2 >>
rect 48 133 49 134 
<< m1 >>
rect 49 133 50 134 
<< m1 >>
rect 50 133 51 134 
<< m1 >>
rect 51 133 52 134 
<< m1 >>
rect 52 133 53 134 
<< m1 >>
rect 58 133 59 134 
<< m2 >>
rect 59 133 60 134 
<< m2 >>
rect 61 133 62 134 
<< m1 >>
rect 62 133 63 134 
<< m1 >>
rect 64 133 65 134 
<< m1 >>
rect 73 133 74 134 
<< m1 >>
rect 78 133 79 134 
<< m1 >>
rect 82 133 83 134 
<< m1 >>
rect 85 133 86 134 
<< m1 >>
rect 91 133 92 134 
<< m2 >>
rect 92 133 93 134 
<< m1 >>
rect 106 133 107 134 
<< m1 >>
rect 109 133 110 134 
<< m1 >>
rect 130 133 131 134 
<< m1 >>
rect 132 133 133 134 
<< m1 >>
rect 136 133 137 134 
<< m2 >>
rect 136 133 137 134 
<< m1 >>
rect 145 133 146 134 
<< m2 >>
rect 145 133 146 134 
<< m1 >>
rect 147 133 148 134 
<< m1 >>
rect 154 133 155 134 
<< m1 >>
rect 156 133 157 134 
<< m1 >>
rect 157 133 158 134 
<< m1 >>
rect 158 133 159 134 
<< m1 >>
rect 159 133 160 134 
<< m1 >>
rect 160 133 161 134 
<< m1 >>
rect 163 133 164 134 
<< m2 >>
rect 164 133 165 134 
<< m1 >>
rect 168 133 169 134 
<< m2 >>
rect 168 133 169 134 
<< m2c >>
rect 168 133 169 134 
<< m1 >>
rect 168 133 169 134 
<< m2 >>
rect 168 133 169 134 
<< m2 >>
rect 169 133 170 134 
<< m1 >>
rect 170 133 171 134 
<< m2 >>
rect 170 133 171 134 
<< m2 >>
rect 171 133 172 134 
<< m1 >>
rect 172 133 173 134 
<< m2 >>
rect 172 133 173 134 
<< m2 >>
rect 173 133 174 134 
<< m1 >>
rect 174 133 175 134 
<< m2 >>
rect 174 133 175 134 
<< m2c >>
rect 174 133 175 134 
<< m1 >>
rect 174 133 175 134 
<< m2 >>
rect 174 133 175 134 
<< m1 >>
rect 175 133 176 134 
<< m1 >>
rect 176 133 177 134 
<< m2 >>
rect 176 133 177 134 
<< m1 >>
rect 177 133 178 134 
<< m1 >>
rect 178 133 179 134 
<< m2 >>
rect 178 133 179 134 
<< m1 >>
rect 179 133 180 134 
<< m1 >>
rect 180 133 181 134 
<< m1 >>
rect 181 133 182 134 
<< m1 >>
rect 182 133 183 134 
<< m1 >>
rect 183 133 184 134 
<< m1 >>
rect 184 133 185 134 
<< m1 >>
rect 185 133 186 134 
<< m1 >>
rect 186 133 187 134 
<< m1 >>
rect 187 133 188 134 
<< m1 >>
rect 188 133 189 134 
<< m2 >>
rect 192 133 193 134 
<< m1 >>
rect 199 133 200 134 
<< m1 >>
rect 201 133 202 134 
<< m1 >>
rect 205 133 206 134 
<< m1 >>
rect 226 133 227 134 
<< m2 >>
rect 226 133 227 134 
<< m1 >>
rect 235 133 236 134 
<< m2 >>
rect 235 133 236 134 
<< m1 >>
rect 237 133 238 134 
<< m1 >>
rect 238 133 239 134 
<< m1 >>
rect 239 133 240 134 
<< m1 >>
rect 240 133 241 134 
<< m1 >>
rect 241 133 242 134 
<< m2 >>
rect 241 133 242 134 
<< m1 >>
rect 242 133 243 134 
<< m1 >>
rect 243 133 244 134 
<< m1 >>
rect 244 133 245 134 
<< m1 >>
rect 245 133 246 134 
<< m1 >>
rect 246 133 247 134 
<< m1 >>
rect 247 133 248 134 
<< m1 >>
rect 248 133 249 134 
<< m1 >>
rect 249 133 250 134 
<< m1 >>
rect 250 133 251 134 
<< m1 >>
rect 251 133 252 134 
<< m1 >>
rect 252 133 253 134 
<< m1 >>
rect 253 133 254 134 
<< m2 >>
rect 253 133 254 134 
<< m1 >>
rect 254 133 255 134 
<< m1 >>
rect 255 133 256 134 
<< m2 >>
rect 255 133 256 134 
<< m1 >>
rect 256 133 257 134 
<< m1 >>
rect 257 133 258 134 
<< m1 >>
rect 258 133 259 134 
<< m2 >>
rect 258 133 259 134 
<< m1 >>
rect 259 133 260 134 
<< m1 >>
rect 260 133 261 134 
<< m1 >>
rect 261 133 262 134 
<< m1 >>
rect 262 133 263 134 
<< m2 >>
rect 262 133 263 134 
<< m1 >>
rect 263 133 264 134 
<< m1 >>
rect 264 133 265 134 
<< m1 >>
rect 265 133 266 134 
<< m1 >>
rect 266 133 267 134 
<< m1 >>
rect 267 133 268 134 
<< m1 >>
rect 268 133 269 134 
<< m2 >>
rect 268 133 269 134 
<< m1 >>
rect 269 133 270 134 
<< m1 >>
rect 270 133 271 134 
<< m1 >>
rect 271 133 272 134 
<< m1 >>
rect 272 133 273 134 
<< m2 >>
rect 272 133 273 134 
<< m1 >>
rect 273 133 274 134 
<< m1 >>
rect 274 133 275 134 
<< m2 >>
rect 274 133 275 134 
<< m1 >>
rect 275 133 276 134 
<< m1 >>
rect 276 133 277 134 
<< m2 >>
rect 276 133 277 134 
<< m1 >>
rect 277 133 278 134 
<< m1 >>
rect 278 133 279 134 
<< m1 >>
rect 279 133 280 134 
<< m1 >>
rect 280 133 281 134 
<< m2 >>
rect 280 133 281 134 
<< m1 >>
rect 281 133 282 134 
<< m1 >>
rect 282 133 283 134 
<< m2 >>
rect 282 133 283 134 
<< m1 >>
rect 283 133 284 134 
<< m1 >>
rect 284 133 285 134 
<< m1 >>
rect 285 133 286 134 
<< m1 >>
rect 286 133 287 134 
<< m1 >>
rect 289 133 290 134 
<< m1 >>
rect 296 133 297 134 
<< m1 >>
rect 298 133 299 134 
<< m1 >>
rect 307 133 308 134 
<< m2 >>
rect 308 133 309 134 
<< m1 >>
rect 325 133 326 134 
<< m1 >>
rect 327 133 328 134 
<< m1 >>
rect 329 133 330 134 
<< m1 >>
rect 338 133 339 134 
<< m2 >>
rect 338 133 339 134 
<< m2c >>
rect 338 133 339 134 
<< m1 >>
rect 338 133 339 134 
<< m2 >>
rect 338 133 339 134 
<< m1 >>
rect 345 133 346 134 
<< m1 >>
rect 10 134 11 135 
<< m1 >>
rect 19 134 20 135 
<< m2 >>
rect 19 134 20 135 
<< m1 >>
rect 21 134 22 135 
<< m1 >>
rect 23 134 24 135 
<< m2 >>
rect 27 134 28 135 
<< m1 >>
rect 28 134 29 135 
<< m1 >>
rect 37 134 38 135 
<< m2 >>
rect 38 134 39 135 
<< m1 >>
rect 42 134 43 135 
<< m1 >>
rect 46 134 47 135 
<< m1 >>
rect 52 134 53 135 
<< m1 >>
rect 58 134 59 135 
<< m2 >>
rect 59 134 60 135 
<< m2 >>
rect 61 134 62 135 
<< m1 >>
rect 62 134 63 135 
<< m1 >>
rect 64 134 65 135 
<< m1 >>
rect 73 134 74 135 
<< m1 >>
rect 78 134 79 135 
<< m1 >>
rect 82 134 83 135 
<< m1 >>
rect 85 134 86 135 
<< m1 >>
rect 91 134 92 135 
<< m2 >>
rect 92 134 93 135 
<< m1 >>
rect 106 134 107 135 
<< m1 >>
rect 109 134 110 135 
<< m1 >>
rect 130 134 131 135 
<< m1 >>
rect 132 134 133 135 
<< m1 >>
rect 136 134 137 135 
<< m2 >>
rect 136 134 137 135 
<< m1 >>
rect 145 134 146 135 
<< m2 >>
rect 145 134 146 135 
<< m1 >>
rect 147 134 148 135 
<< m1 >>
rect 154 134 155 135 
<< m1 >>
rect 156 134 157 135 
<< m1 >>
rect 160 134 161 135 
<< m1 >>
rect 163 134 164 135 
<< m2 >>
rect 164 134 165 135 
<< m1 >>
rect 170 134 171 135 
<< m1 >>
rect 172 134 173 135 
<< m2 >>
rect 176 134 177 135 
<< m2 >>
rect 178 134 179 135 
<< m1 >>
rect 188 134 189 135 
<< m2 >>
rect 189 134 190 135 
<< m1 >>
rect 190 134 191 135 
<< m2 >>
rect 190 134 191 135 
<< m2c >>
rect 190 134 191 135 
<< m1 >>
rect 190 134 191 135 
<< m2 >>
rect 190 134 191 135 
<< m1 >>
rect 191 134 192 135 
<< m1 >>
rect 192 134 193 135 
<< m2 >>
rect 192 134 193 135 
<< m2c >>
rect 192 134 193 135 
<< m1 >>
rect 192 134 193 135 
<< m2 >>
rect 192 134 193 135 
<< m1 >>
rect 199 134 200 135 
<< m1 >>
rect 201 134 202 135 
<< m1 >>
rect 205 134 206 135 
<< m1 >>
rect 226 134 227 135 
<< m2 >>
rect 226 134 227 135 
<< m1 >>
rect 235 134 236 135 
<< m2 >>
rect 235 134 236 135 
<< m1 >>
rect 237 134 238 135 
<< m2 >>
rect 241 134 242 135 
<< m2 >>
rect 253 134 254 135 
<< m2 >>
rect 255 134 256 135 
<< m2 >>
rect 258 134 259 135 
<< m2 >>
rect 259 134 260 135 
<< m2 >>
rect 260 134 261 135 
<< m2 >>
rect 262 134 263 135 
<< m2 >>
rect 268 134 269 135 
<< m2 >>
rect 272 134 273 135 
<< m2 >>
rect 274 134 275 135 
<< m2 >>
rect 276 134 277 135 
<< m2 >>
rect 280 134 281 135 
<< m2 >>
rect 282 134 283 135 
<< m1 >>
rect 289 134 290 135 
<< m1 >>
rect 296 134 297 135 
<< m1 >>
rect 298 134 299 135 
<< m1 >>
rect 307 134 308 135 
<< m2 >>
rect 308 134 309 135 
<< m1 >>
rect 325 134 326 135 
<< m1 >>
rect 327 134 328 135 
<< m1 >>
rect 329 134 330 135 
<< m2 >>
rect 338 134 339 135 
<< m2 >>
rect 339 134 340 135 
<< m2 >>
rect 340 134 341 135 
<< m2 >>
rect 341 134 342 135 
<< m2 >>
rect 342 134 343 135 
<< m2 >>
rect 343 134 344 135 
<< m1 >>
rect 345 134 346 135 
<< m1 >>
rect 10 135 11 136 
<< m1 >>
rect 13 135 14 136 
<< m1 >>
rect 14 135 15 136 
<< m1 >>
rect 15 135 16 136 
<< m1 >>
rect 16 135 17 136 
<< m1 >>
rect 17 135 18 136 
<< m2 >>
rect 17 135 18 136 
<< m2c >>
rect 17 135 18 136 
<< m1 >>
rect 17 135 18 136 
<< m2 >>
rect 17 135 18 136 
<< m2 >>
rect 18 135 19 136 
<< m1 >>
rect 19 135 20 136 
<< m2 >>
rect 19 135 20 136 
<< m1 >>
rect 21 135 22 136 
<< m1 >>
rect 23 135 24 136 
<< m2 >>
rect 27 135 28 136 
<< m1 >>
rect 28 135 29 136 
<< m1 >>
rect 37 135 38 136 
<< m2 >>
rect 38 135 39 136 
<< m1 >>
rect 42 135 43 136 
<< m1 >>
rect 46 135 47 136 
<< m1 >>
rect 52 135 53 136 
<< m1 >>
rect 58 135 59 136 
<< m2 >>
rect 59 135 60 136 
<< m2 >>
rect 61 135 62 136 
<< m1 >>
rect 62 135 63 136 
<< m1 >>
rect 64 135 65 136 
<< m1 >>
rect 67 135 68 136 
<< m1 >>
rect 68 135 69 136 
<< m1 >>
rect 69 135 70 136 
<< m1 >>
rect 70 135 71 136 
<< m1 >>
rect 71 135 72 136 
<< m1 >>
rect 72 135 73 136 
<< m1 >>
rect 73 135 74 136 
<< m1 >>
rect 78 135 79 136 
<< m1 >>
rect 82 135 83 136 
<< m1 >>
rect 85 135 86 136 
<< m1 >>
rect 91 135 92 136 
<< m2 >>
rect 92 135 93 136 
<< m1 >>
rect 106 135 107 136 
<< m1 >>
rect 109 135 110 136 
<< m1 >>
rect 130 135 131 136 
<< m1 >>
rect 132 135 133 136 
<< m1 >>
rect 136 135 137 136 
<< m2 >>
rect 136 135 137 136 
<< m1 >>
rect 145 135 146 136 
<< m2 >>
rect 145 135 146 136 
<< m1 >>
rect 147 135 148 136 
<< m1 >>
rect 154 135 155 136 
<< m1 >>
rect 156 135 157 136 
<< m1 >>
rect 160 135 161 136 
<< m1 >>
rect 163 135 164 136 
<< m2 >>
rect 164 135 165 136 
<< m1 >>
rect 170 135 171 136 
<< m1 >>
rect 172 135 173 136 
<< m1 >>
rect 176 135 177 136 
<< m2 >>
rect 176 135 177 136 
<< m2c >>
rect 176 135 177 136 
<< m1 >>
rect 176 135 177 136 
<< m2 >>
rect 176 135 177 136 
<< m1 >>
rect 177 135 178 136 
<< m1 >>
rect 178 135 179 136 
<< m2 >>
rect 178 135 179 136 
<< m1 >>
rect 179 135 180 136 
<< m1 >>
rect 180 135 181 136 
<< m1 >>
rect 181 135 182 136 
<< m1 >>
rect 184 135 185 136 
<< m1 >>
rect 185 135 186 136 
<< m1 >>
rect 186 135 187 136 
<< m2 >>
rect 186 135 187 136 
<< m2c >>
rect 186 135 187 136 
<< m1 >>
rect 186 135 187 136 
<< m2 >>
rect 186 135 187 136 
<< m2 >>
rect 187 135 188 136 
<< m1 >>
rect 188 135 189 136 
<< m2 >>
rect 188 135 189 136 
<< m2 >>
rect 189 135 190 136 
<< m1 >>
rect 199 135 200 136 
<< m1 >>
rect 201 135 202 136 
<< m1 >>
rect 205 135 206 136 
<< m1 >>
rect 226 135 227 136 
<< m2 >>
rect 226 135 227 136 
<< m1 >>
rect 235 135 236 136 
<< m2 >>
rect 235 135 236 136 
<< m2 >>
rect 236 135 237 136 
<< m1 >>
rect 237 135 238 136 
<< m2 >>
rect 237 135 238 136 
<< m2 >>
rect 238 135 239 136 
<< m1 >>
rect 239 135 240 136 
<< m2 >>
rect 239 135 240 136 
<< m2c >>
rect 239 135 240 136 
<< m1 >>
rect 239 135 240 136 
<< m2 >>
rect 239 135 240 136 
<< m1 >>
rect 240 135 241 136 
<< m2 >>
rect 241 135 242 136 
<< m1 >>
rect 253 135 254 136 
<< m2 >>
rect 253 135 254 136 
<< m2c >>
rect 253 135 254 136 
<< m1 >>
rect 253 135 254 136 
<< m2 >>
rect 253 135 254 136 
<< m1 >>
rect 255 135 256 136 
<< m2 >>
rect 255 135 256 136 
<< m2c >>
rect 255 135 256 136 
<< m1 >>
rect 255 135 256 136 
<< m2 >>
rect 255 135 256 136 
<< m1 >>
rect 260 135 261 136 
<< m2 >>
rect 260 135 261 136 
<< m2c >>
rect 260 135 261 136 
<< m1 >>
rect 260 135 261 136 
<< m2 >>
rect 260 135 261 136 
<< m1 >>
rect 262 135 263 136 
<< m2 >>
rect 262 135 263 136 
<< m2c >>
rect 262 135 263 136 
<< m1 >>
rect 262 135 263 136 
<< m2 >>
rect 262 135 263 136 
<< m1 >>
rect 268 135 269 136 
<< m2 >>
rect 268 135 269 136 
<< m2c >>
rect 268 135 269 136 
<< m1 >>
rect 268 135 269 136 
<< m2 >>
rect 268 135 269 136 
<< m1 >>
rect 272 135 273 136 
<< m2 >>
rect 272 135 273 136 
<< m2c >>
rect 272 135 273 136 
<< m1 >>
rect 272 135 273 136 
<< m2 >>
rect 272 135 273 136 
<< m1 >>
rect 274 135 275 136 
<< m2 >>
rect 274 135 275 136 
<< m2c >>
rect 274 135 275 136 
<< m1 >>
rect 274 135 275 136 
<< m2 >>
rect 274 135 275 136 
<< m1 >>
rect 276 135 277 136 
<< m2 >>
rect 276 135 277 136 
<< m2c >>
rect 276 135 277 136 
<< m1 >>
rect 276 135 277 136 
<< m2 >>
rect 276 135 277 136 
<< m1 >>
rect 280 135 281 136 
<< m2 >>
rect 280 135 281 136 
<< m1 >>
rect 281 135 282 136 
<< m1 >>
rect 282 135 283 136 
<< m2 >>
rect 282 135 283 136 
<< m2c >>
rect 282 135 283 136 
<< m1 >>
rect 282 135 283 136 
<< m2 >>
rect 282 135 283 136 
<< m1 >>
rect 289 135 290 136 
<< m1 >>
rect 296 135 297 136 
<< m1 >>
rect 298 135 299 136 
<< m1 >>
rect 307 135 308 136 
<< m2 >>
rect 308 135 309 136 
<< m1 >>
rect 325 135 326 136 
<< m1 >>
rect 327 135 328 136 
<< m1 >>
rect 329 135 330 136 
<< m1 >>
rect 337 135 338 136 
<< m1 >>
rect 338 135 339 136 
<< m1 >>
rect 339 135 340 136 
<< m1 >>
rect 340 135 341 136 
<< m1 >>
rect 341 135 342 136 
<< m1 >>
rect 342 135 343 136 
<< m1 >>
rect 343 135 344 136 
<< m2 >>
rect 343 135 344 136 
<< m1 >>
rect 345 135 346 136 
<< m1 >>
rect 10 136 11 137 
<< m1 >>
rect 13 136 14 137 
<< m1 >>
rect 19 136 20 137 
<< m1 >>
rect 21 136 22 137 
<< m1 >>
rect 23 136 24 137 
<< m2 >>
rect 27 136 28 137 
<< m1 >>
rect 28 136 29 137 
<< m1 >>
rect 37 136 38 137 
<< m2 >>
rect 38 136 39 137 
<< m1 >>
rect 42 136 43 137 
<< m1 >>
rect 46 136 47 137 
<< m1 >>
rect 52 136 53 137 
<< m1 >>
rect 58 136 59 137 
<< m2 >>
rect 59 136 60 137 
<< m2 >>
rect 61 136 62 137 
<< m1 >>
rect 62 136 63 137 
<< m1 >>
rect 64 136 65 137 
<< m1 >>
rect 67 136 68 137 
<< m1 >>
rect 78 136 79 137 
<< m1 >>
rect 82 136 83 137 
<< m1 >>
rect 85 136 86 137 
<< m1 >>
rect 91 136 92 137 
<< m2 >>
rect 92 136 93 137 
<< m1 >>
rect 106 136 107 137 
<< m1 >>
rect 109 136 110 137 
<< m1 >>
rect 130 136 131 137 
<< m1 >>
rect 132 136 133 137 
<< m1 >>
rect 136 136 137 137 
<< m2 >>
rect 136 136 137 137 
<< m1 >>
rect 142 136 143 137 
<< m1 >>
rect 143 136 144 137 
<< m2 >>
rect 143 136 144 137 
<< m2c >>
rect 143 136 144 137 
<< m1 >>
rect 143 136 144 137 
<< m2 >>
rect 143 136 144 137 
<< m2 >>
rect 144 136 145 137 
<< m1 >>
rect 145 136 146 137 
<< m2 >>
rect 145 136 146 137 
<< m1 >>
rect 147 136 148 137 
<< m2 >>
rect 153 136 154 137 
<< m1 >>
rect 154 136 155 137 
<< m2 >>
rect 154 136 155 137 
<< m2 >>
rect 155 136 156 137 
<< m1 >>
rect 156 136 157 137 
<< m2 >>
rect 156 136 157 137 
<< m2c >>
rect 156 136 157 137 
<< m1 >>
rect 156 136 157 137 
<< m2 >>
rect 156 136 157 137 
<< m1 >>
rect 160 136 161 137 
<< m1 >>
rect 163 136 164 137 
<< m2 >>
rect 164 136 165 137 
<< m1 >>
rect 170 136 171 137 
<< m1 >>
rect 172 136 173 137 
<< m2 >>
rect 178 136 179 137 
<< m1 >>
rect 181 136 182 137 
<< m1 >>
rect 184 136 185 137 
<< m1 >>
rect 188 136 189 137 
<< m1 >>
rect 199 136 200 137 
<< m1 >>
rect 201 136 202 137 
<< m1 >>
rect 205 136 206 137 
<< m1 >>
rect 226 136 227 137 
<< m2 >>
rect 226 136 227 137 
<< m1 >>
rect 235 136 236 137 
<< m1 >>
rect 237 136 238 137 
<< m1 >>
rect 240 136 241 137 
<< m2 >>
rect 241 136 242 137 
<< m1 >>
rect 253 136 254 137 
<< m1 >>
rect 255 136 256 137 
<< m1 >>
rect 260 136 261 137 
<< m1 >>
rect 262 136 263 137 
<< m1 >>
rect 268 136 269 137 
<< m1 >>
rect 272 136 273 137 
<< m1 >>
rect 274 136 275 137 
<< m1 >>
rect 276 136 277 137 
<< m1 >>
rect 280 136 281 137 
<< m2 >>
rect 280 136 281 137 
<< m1 >>
rect 289 136 290 137 
<< m1 >>
rect 296 136 297 137 
<< m1 >>
rect 298 136 299 137 
<< m1 >>
rect 307 136 308 137 
<< m2 >>
rect 308 136 309 137 
<< m1 >>
rect 325 136 326 137 
<< m1 >>
rect 327 136 328 137 
<< m1 >>
rect 329 136 330 137 
<< m1 >>
rect 337 136 338 137 
<< m1 >>
rect 343 136 344 137 
<< m2 >>
rect 343 136 344 137 
<< m1 >>
rect 345 136 346 137 
<< m1 >>
rect 10 137 11 138 
<< m1 >>
rect 13 137 14 138 
<< m1 >>
rect 19 137 20 138 
<< m1 >>
rect 21 137 22 138 
<< m1 >>
rect 23 137 24 138 
<< m2 >>
rect 27 137 28 138 
<< m1 >>
rect 28 137 29 138 
<< m1 >>
rect 37 137 38 138 
<< m2 >>
rect 38 137 39 138 
<< m1 >>
rect 42 137 43 138 
<< m1 >>
rect 46 137 47 138 
<< m1 >>
rect 52 137 53 138 
<< m1 >>
rect 58 137 59 138 
<< m2 >>
rect 59 137 60 138 
<< m2 >>
rect 61 137 62 138 
<< m1 >>
rect 62 137 63 138 
<< m1 >>
rect 64 137 65 138 
<< m1 >>
rect 67 137 68 138 
<< m1 >>
rect 78 137 79 138 
<< m1 >>
rect 82 137 83 138 
<< m1 >>
rect 85 137 86 138 
<< m1 >>
rect 91 137 92 138 
<< m2 >>
rect 92 137 93 138 
<< m1 >>
rect 106 137 107 138 
<< m1 >>
rect 109 137 110 138 
<< m1 >>
rect 130 137 131 138 
<< m1 >>
rect 132 137 133 138 
<< m1 >>
rect 136 137 137 138 
<< m2 >>
rect 136 137 137 138 
<< m1 >>
rect 142 137 143 138 
<< m1 >>
rect 145 137 146 138 
<< m1 >>
rect 147 137 148 138 
<< m2 >>
rect 153 137 154 138 
<< m1 >>
rect 154 137 155 138 
<< m1 >>
rect 160 137 161 138 
<< m1 >>
rect 163 137 164 138 
<< m2 >>
rect 164 137 165 138 
<< m1 >>
rect 170 137 171 138 
<< m1 >>
rect 172 137 173 138 
<< m1 >>
rect 178 137 179 138 
<< m2 >>
rect 178 137 179 138 
<< m2c >>
rect 178 137 179 138 
<< m1 >>
rect 178 137 179 138 
<< m2 >>
rect 178 137 179 138 
<< m1 >>
rect 181 137 182 138 
<< m1 >>
rect 184 137 185 138 
<< m1 >>
rect 188 137 189 138 
<< m1 >>
rect 199 137 200 138 
<< m1 >>
rect 201 137 202 138 
<< m1 >>
rect 205 137 206 138 
<< m1 >>
rect 226 137 227 138 
<< m2 >>
rect 226 137 227 138 
<< m1 >>
rect 235 137 236 138 
<< m1 >>
rect 237 137 238 138 
<< m2 >>
rect 238 137 239 138 
<< m2 >>
rect 239 137 240 138 
<< m1 >>
rect 240 137 241 138 
<< m2 >>
rect 240 137 241 138 
<< m2 >>
rect 241 137 242 138 
<< m1 >>
rect 253 137 254 138 
<< m1 >>
rect 255 137 256 138 
<< m1 >>
rect 260 137 261 138 
<< m1 >>
rect 262 137 263 138 
<< m1 >>
rect 268 137 269 138 
<< m1 >>
rect 272 137 273 138 
<< m1 >>
rect 274 137 275 138 
<< m1 >>
rect 276 137 277 138 
<< m2 >>
rect 277 137 278 138 
<< m1 >>
rect 278 137 279 138 
<< m2 >>
rect 278 137 279 138 
<< m2c >>
rect 278 137 279 138 
<< m1 >>
rect 278 137 279 138 
<< m2 >>
rect 278 137 279 138 
<< m1 >>
rect 279 137 280 138 
<< m1 >>
rect 280 137 281 138 
<< m2 >>
rect 280 137 281 138 
<< m1 >>
rect 289 137 290 138 
<< m1 >>
rect 296 137 297 138 
<< m1 >>
rect 298 137 299 138 
<< m1 >>
rect 307 137 308 138 
<< m2 >>
rect 308 137 309 138 
<< m1 >>
rect 325 137 326 138 
<< m1 >>
rect 327 137 328 138 
<< m1 >>
rect 329 137 330 138 
<< m1 >>
rect 337 137 338 138 
<< m1 >>
rect 343 137 344 138 
<< m2 >>
rect 343 137 344 138 
<< m1 >>
rect 345 137 346 138 
<< m1 >>
rect 10 138 11 139 
<< pdiffusion >>
rect 12 138 13 139 
<< m1 >>
rect 13 138 14 139 
<< pdiffusion >>
rect 13 138 14 139 
<< pdiffusion >>
rect 14 138 15 139 
<< pdiffusion >>
rect 15 138 16 139 
<< pdiffusion >>
rect 16 138 17 139 
<< pdiffusion >>
rect 17 138 18 139 
<< m1 >>
rect 19 138 20 139 
<< m1 >>
rect 21 138 22 139 
<< m1 >>
rect 23 138 24 139 
<< m2 >>
rect 27 138 28 139 
<< m1 >>
rect 28 138 29 139 
<< pdiffusion >>
rect 30 138 31 139 
<< pdiffusion >>
rect 31 138 32 139 
<< pdiffusion >>
rect 32 138 33 139 
<< pdiffusion >>
rect 33 138 34 139 
<< pdiffusion >>
rect 34 138 35 139 
<< pdiffusion >>
rect 35 138 36 139 
<< m1 >>
rect 37 138 38 139 
<< m2 >>
rect 38 138 39 139 
<< m1 >>
rect 42 138 43 139 
<< m1 >>
rect 46 138 47 139 
<< pdiffusion >>
rect 48 138 49 139 
<< pdiffusion >>
rect 49 138 50 139 
<< pdiffusion >>
rect 50 138 51 139 
<< pdiffusion >>
rect 51 138 52 139 
<< m1 >>
rect 52 138 53 139 
<< pdiffusion >>
rect 52 138 53 139 
<< pdiffusion >>
rect 53 138 54 139 
<< m1 >>
rect 58 138 59 139 
<< m2 >>
rect 59 138 60 139 
<< m2 >>
rect 61 138 62 139 
<< m1 >>
rect 62 138 63 139 
<< m1 >>
rect 64 138 65 139 
<< pdiffusion >>
rect 66 138 67 139 
<< m1 >>
rect 67 138 68 139 
<< pdiffusion >>
rect 67 138 68 139 
<< pdiffusion >>
rect 68 138 69 139 
<< pdiffusion >>
rect 69 138 70 139 
<< pdiffusion >>
rect 70 138 71 139 
<< pdiffusion >>
rect 71 138 72 139 
<< m1 >>
rect 78 138 79 139 
<< m1 >>
rect 82 138 83 139 
<< pdiffusion >>
rect 84 138 85 139 
<< m1 >>
rect 85 138 86 139 
<< pdiffusion >>
rect 85 138 86 139 
<< pdiffusion >>
rect 86 138 87 139 
<< pdiffusion >>
rect 87 138 88 139 
<< pdiffusion >>
rect 88 138 89 139 
<< pdiffusion >>
rect 89 138 90 139 
<< m1 >>
rect 91 138 92 139 
<< m2 >>
rect 92 138 93 139 
<< pdiffusion >>
rect 102 138 103 139 
<< pdiffusion >>
rect 103 138 104 139 
<< pdiffusion >>
rect 104 138 105 139 
<< pdiffusion >>
rect 105 138 106 139 
<< m1 >>
rect 106 138 107 139 
<< pdiffusion >>
rect 106 138 107 139 
<< pdiffusion >>
rect 107 138 108 139 
<< m1 >>
rect 109 138 110 139 
<< pdiffusion >>
rect 120 138 121 139 
<< pdiffusion >>
rect 121 138 122 139 
<< pdiffusion >>
rect 122 138 123 139 
<< pdiffusion >>
rect 123 138 124 139 
<< pdiffusion >>
rect 124 138 125 139 
<< pdiffusion >>
rect 125 138 126 139 
<< m1 >>
rect 130 138 131 139 
<< m1 >>
rect 132 138 133 139 
<< m1 >>
rect 136 138 137 139 
<< m2 >>
rect 136 138 137 139 
<< pdiffusion >>
rect 138 138 139 139 
<< pdiffusion >>
rect 139 138 140 139 
<< pdiffusion >>
rect 140 138 141 139 
<< pdiffusion >>
rect 141 138 142 139 
<< m1 >>
rect 142 138 143 139 
<< pdiffusion >>
rect 142 138 143 139 
<< pdiffusion >>
rect 143 138 144 139 
<< m1 >>
rect 145 138 146 139 
<< m1 >>
rect 147 138 148 139 
<< m2 >>
rect 153 138 154 139 
<< m1 >>
rect 154 138 155 139 
<< pdiffusion >>
rect 156 138 157 139 
<< pdiffusion >>
rect 157 138 158 139 
<< pdiffusion >>
rect 158 138 159 139 
<< pdiffusion >>
rect 159 138 160 139 
<< m1 >>
rect 160 138 161 139 
<< pdiffusion >>
rect 160 138 161 139 
<< pdiffusion >>
rect 161 138 162 139 
<< m1 >>
rect 163 138 164 139 
<< m2 >>
rect 164 138 165 139 
<< m1 >>
rect 170 138 171 139 
<< m1 >>
rect 172 138 173 139 
<< pdiffusion >>
rect 174 138 175 139 
<< pdiffusion >>
rect 175 138 176 139 
<< pdiffusion >>
rect 176 138 177 139 
<< pdiffusion >>
rect 177 138 178 139 
<< m1 >>
rect 178 138 179 139 
<< pdiffusion >>
rect 178 138 179 139 
<< pdiffusion >>
rect 179 138 180 139 
<< m1 >>
rect 181 138 182 139 
<< m1 >>
rect 184 138 185 139 
<< m1 >>
rect 188 138 189 139 
<< pdiffusion >>
rect 192 138 193 139 
<< pdiffusion >>
rect 193 138 194 139 
<< pdiffusion >>
rect 194 138 195 139 
<< pdiffusion >>
rect 195 138 196 139 
<< pdiffusion >>
rect 196 138 197 139 
<< pdiffusion >>
rect 197 138 198 139 
<< m1 >>
rect 199 138 200 139 
<< m1 >>
rect 201 138 202 139 
<< m1 >>
rect 205 138 206 139 
<< pdiffusion >>
rect 210 138 211 139 
<< pdiffusion >>
rect 211 138 212 139 
<< pdiffusion >>
rect 212 138 213 139 
<< pdiffusion >>
rect 213 138 214 139 
<< pdiffusion >>
rect 214 138 215 139 
<< pdiffusion >>
rect 215 138 216 139 
<< m1 >>
rect 226 138 227 139 
<< m2 >>
rect 226 138 227 139 
<< pdiffusion >>
rect 228 138 229 139 
<< pdiffusion >>
rect 229 138 230 139 
<< pdiffusion >>
rect 230 138 231 139 
<< pdiffusion >>
rect 231 138 232 139 
<< pdiffusion >>
rect 232 138 233 139 
<< pdiffusion >>
rect 233 138 234 139 
<< m1 >>
rect 235 138 236 139 
<< m1 >>
rect 237 138 238 139 
<< m2 >>
rect 238 138 239 139 
<< m1 >>
rect 240 138 241 139 
<< pdiffusion >>
rect 246 138 247 139 
<< pdiffusion >>
rect 247 138 248 139 
<< pdiffusion >>
rect 248 138 249 139 
<< pdiffusion >>
rect 249 138 250 139 
<< pdiffusion >>
rect 250 138 251 139 
<< pdiffusion >>
rect 251 138 252 139 
<< m1 >>
rect 253 138 254 139 
<< m1 >>
rect 255 138 256 139 
<< m1 >>
rect 260 138 261 139 
<< m1 >>
rect 262 138 263 139 
<< pdiffusion >>
rect 264 138 265 139 
<< pdiffusion >>
rect 265 138 266 139 
<< pdiffusion >>
rect 266 138 267 139 
<< pdiffusion >>
rect 267 138 268 139 
<< m1 >>
rect 268 138 269 139 
<< pdiffusion >>
rect 268 138 269 139 
<< pdiffusion >>
rect 269 138 270 139 
<< m1 >>
rect 272 138 273 139 
<< m1 >>
rect 274 138 275 139 
<< m1 >>
rect 276 138 277 139 
<< m2 >>
rect 277 138 278 139 
<< m2 >>
rect 280 138 281 139 
<< pdiffusion >>
rect 282 138 283 139 
<< pdiffusion >>
rect 283 138 284 139 
<< pdiffusion >>
rect 284 138 285 139 
<< pdiffusion >>
rect 285 138 286 139 
<< pdiffusion >>
rect 286 138 287 139 
<< pdiffusion >>
rect 287 138 288 139 
<< m1 >>
rect 289 138 290 139 
<< m1 >>
rect 296 138 297 139 
<< m1 >>
rect 298 138 299 139 
<< pdiffusion >>
rect 300 138 301 139 
<< pdiffusion >>
rect 301 138 302 139 
<< pdiffusion >>
rect 302 138 303 139 
<< pdiffusion >>
rect 303 138 304 139 
<< pdiffusion >>
rect 304 138 305 139 
<< pdiffusion >>
rect 305 138 306 139 
<< m1 >>
rect 307 138 308 139 
<< m2 >>
rect 308 138 309 139 
<< pdiffusion >>
rect 318 138 319 139 
<< pdiffusion >>
rect 319 138 320 139 
<< pdiffusion >>
rect 320 138 321 139 
<< pdiffusion >>
rect 321 138 322 139 
<< pdiffusion >>
rect 322 138 323 139 
<< pdiffusion >>
rect 323 138 324 139 
<< m1 >>
rect 325 138 326 139 
<< m1 >>
rect 327 138 328 139 
<< m1 >>
rect 329 138 330 139 
<< pdiffusion >>
rect 336 138 337 139 
<< m1 >>
rect 337 138 338 139 
<< pdiffusion >>
rect 337 138 338 139 
<< pdiffusion >>
rect 338 138 339 139 
<< pdiffusion >>
rect 339 138 340 139 
<< pdiffusion >>
rect 340 138 341 139 
<< pdiffusion >>
rect 341 138 342 139 
<< m1 >>
rect 343 138 344 139 
<< m2 >>
rect 343 138 344 139 
<< m1 >>
rect 345 138 346 139 
<< m1 >>
rect 10 139 11 140 
<< pdiffusion >>
rect 12 139 13 140 
<< pdiffusion >>
rect 13 139 14 140 
<< pdiffusion >>
rect 14 139 15 140 
<< pdiffusion >>
rect 15 139 16 140 
<< pdiffusion >>
rect 16 139 17 140 
<< pdiffusion >>
rect 17 139 18 140 
<< m1 >>
rect 19 139 20 140 
<< m1 >>
rect 21 139 22 140 
<< m1 >>
rect 23 139 24 140 
<< m2 >>
rect 27 139 28 140 
<< m1 >>
rect 28 139 29 140 
<< pdiffusion >>
rect 30 139 31 140 
<< pdiffusion >>
rect 31 139 32 140 
<< pdiffusion >>
rect 32 139 33 140 
<< pdiffusion >>
rect 33 139 34 140 
<< pdiffusion >>
rect 34 139 35 140 
<< pdiffusion >>
rect 35 139 36 140 
<< m1 >>
rect 37 139 38 140 
<< m2 >>
rect 38 139 39 140 
<< m1 >>
rect 42 139 43 140 
<< m1 >>
rect 46 139 47 140 
<< pdiffusion >>
rect 48 139 49 140 
<< pdiffusion >>
rect 49 139 50 140 
<< pdiffusion >>
rect 50 139 51 140 
<< pdiffusion >>
rect 51 139 52 140 
<< pdiffusion >>
rect 52 139 53 140 
<< pdiffusion >>
rect 53 139 54 140 
<< m1 >>
rect 58 139 59 140 
<< m2 >>
rect 59 139 60 140 
<< m2 >>
rect 61 139 62 140 
<< m1 >>
rect 62 139 63 140 
<< m1 >>
rect 64 139 65 140 
<< pdiffusion >>
rect 66 139 67 140 
<< pdiffusion >>
rect 67 139 68 140 
<< pdiffusion >>
rect 68 139 69 140 
<< pdiffusion >>
rect 69 139 70 140 
<< pdiffusion >>
rect 70 139 71 140 
<< pdiffusion >>
rect 71 139 72 140 
<< m1 >>
rect 78 139 79 140 
<< m1 >>
rect 82 139 83 140 
<< pdiffusion >>
rect 84 139 85 140 
<< pdiffusion >>
rect 85 139 86 140 
<< pdiffusion >>
rect 86 139 87 140 
<< pdiffusion >>
rect 87 139 88 140 
<< pdiffusion >>
rect 88 139 89 140 
<< pdiffusion >>
rect 89 139 90 140 
<< m1 >>
rect 91 139 92 140 
<< m2 >>
rect 92 139 93 140 
<< pdiffusion >>
rect 102 139 103 140 
<< pdiffusion >>
rect 103 139 104 140 
<< pdiffusion >>
rect 104 139 105 140 
<< pdiffusion >>
rect 105 139 106 140 
<< pdiffusion >>
rect 106 139 107 140 
<< pdiffusion >>
rect 107 139 108 140 
<< m1 >>
rect 109 139 110 140 
<< pdiffusion >>
rect 120 139 121 140 
<< pdiffusion >>
rect 121 139 122 140 
<< pdiffusion >>
rect 122 139 123 140 
<< pdiffusion >>
rect 123 139 124 140 
<< pdiffusion >>
rect 124 139 125 140 
<< pdiffusion >>
rect 125 139 126 140 
<< m1 >>
rect 130 139 131 140 
<< m1 >>
rect 132 139 133 140 
<< m1 >>
rect 136 139 137 140 
<< m2 >>
rect 136 139 137 140 
<< pdiffusion >>
rect 138 139 139 140 
<< pdiffusion >>
rect 139 139 140 140 
<< pdiffusion >>
rect 140 139 141 140 
<< pdiffusion >>
rect 141 139 142 140 
<< pdiffusion >>
rect 142 139 143 140 
<< pdiffusion >>
rect 143 139 144 140 
<< m1 >>
rect 145 139 146 140 
<< m1 >>
rect 147 139 148 140 
<< m2 >>
rect 153 139 154 140 
<< m1 >>
rect 154 139 155 140 
<< pdiffusion >>
rect 156 139 157 140 
<< pdiffusion >>
rect 157 139 158 140 
<< pdiffusion >>
rect 158 139 159 140 
<< pdiffusion >>
rect 159 139 160 140 
<< pdiffusion >>
rect 160 139 161 140 
<< pdiffusion >>
rect 161 139 162 140 
<< m1 >>
rect 163 139 164 140 
<< m2 >>
rect 164 139 165 140 
<< m1 >>
rect 170 139 171 140 
<< m1 >>
rect 172 139 173 140 
<< pdiffusion >>
rect 174 139 175 140 
<< pdiffusion >>
rect 175 139 176 140 
<< pdiffusion >>
rect 176 139 177 140 
<< pdiffusion >>
rect 177 139 178 140 
<< pdiffusion >>
rect 178 139 179 140 
<< pdiffusion >>
rect 179 139 180 140 
<< m1 >>
rect 181 139 182 140 
<< m1 >>
rect 184 139 185 140 
<< m1 >>
rect 188 139 189 140 
<< pdiffusion >>
rect 192 139 193 140 
<< pdiffusion >>
rect 193 139 194 140 
<< pdiffusion >>
rect 194 139 195 140 
<< pdiffusion >>
rect 195 139 196 140 
<< pdiffusion >>
rect 196 139 197 140 
<< pdiffusion >>
rect 197 139 198 140 
<< m1 >>
rect 199 139 200 140 
<< m1 >>
rect 201 139 202 140 
<< m1 >>
rect 205 139 206 140 
<< pdiffusion >>
rect 210 139 211 140 
<< pdiffusion >>
rect 211 139 212 140 
<< pdiffusion >>
rect 212 139 213 140 
<< pdiffusion >>
rect 213 139 214 140 
<< pdiffusion >>
rect 214 139 215 140 
<< pdiffusion >>
rect 215 139 216 140 
<< m1 >>
rect 226 139 227 140 
<< m2 >>
rect 226 139 227 140 
<< pdiffusion >>
rect 228 139 229 140 
<< pdiffusion >>
rect 229 139 230 140 
<< pdiffusion >>
rect 230 139 231 140 
<< pdiffusion >>
rect 231 139 232 140 
<< pdiffusion >>
rect 232 139 233 140 
<< pdiffusion >>
rect 233 139 234 140 
<< m1 >>
rect 235 139 236 140 
<< m1 >>
rect 237 139 238 140 
<< m2 >>
rect 238 139 239 140 
<< m1 >>
rect 240 139 241 140 
<< pdiffusion >>
rect 246 139 247 140 
<< pdiffusion >>
rect 247 139 248 140 
<< pdiffusion >>
rect 248 139 249 140 
<< pdiffusion >>
rect 249 139 250 140 
<< pdiffusion >>
rect 250 139 251 140 
<< pdiffusion >>
rect 251 139 252 140 
<< m1 >>
rect 253 139 254 140 
<< m1 >>
rect 255 139 256 140 
<< m1 >>
rect 260 139 261 140 
<< m1 >>
rect 262 139 263 140 
<< pdiffusion >>
rect 264 139 265 140 
<< pdiffusion >>
rect 265 139 266 140 
<< pdiffusion >>
rect 266 139 267 140 
<< pdiffusion >>
rect 267 139 268 140 
<< pdiffusion >>
rect 268 139 269 140 
<< pdiffusion >>
rect 269 139 270 140 
<< m1 >>
rect 272 139 273 140 
<< m1 >>
rect 274 139 275 140 
<< m1 >>
rect 276 139 277 140 
<< m2 >>
rect 277 139 278 140 
<< m1 >>
rect 280 139 281 140 
<< m2 >>
rect 280 139 281 140 
<< m2c >>
rect 280 139 281 140 
<< m1 >>
rect 280 139 281 140 
<< m2 >>
rect 280 139 281 140 
<< pdiffusion >>
rect 282 139 283 140 
<< pdiffusion >>
rect 283 139 284 140 
<< pdiffusion >>
rect 284 139 285 140 
<< pdiffusion >>
rect 285 139 286 140 
<< pdiffusion >>
rect 286 139 287 140 
<< pdiffusion >>
rect 287 139 288 140 
<< m1 >>
rect 289 139 290 140 
<< m1 >>
rect 296 139 297 140 
<< m1 >>
rect 298 139 299 140 
<< pdiffusion >>
rect 300 139 301 140 
<< pdiffusion >>
rect 301 139 302 140 
<< pdiffusion >>
rect 302 139 303 140 
<< pdiffusion >>
rect 303 139 304 140 
<< pdiffusion >>
rect 304 139 305 140 
<< pdiffusion >>
rect 305 139 306 140 
<< m1 >>
rect 307 139 308 140 
<< m2 >>
rect 308 139 309 140 
<< pdiffusion >>
rect 318 139 319 140 
<< pdiffusion >>
rect 319 139 320 140 
<< pdiffusion >>
rect 320 139 321 140 
<< pdiffusion >>
rect 321 139 322 140 
<< pdiffusion >>
rect 322 139 323 140 
<< pdiffusion >>
rect 323 139 324 140 
<< m1 >>
rect 325 139 326 140 
<< m1 >>
rect 327 139 328 140 
<< m1 >>
rect 329 139 330 140 
<< pdiffusion >>
rect 336 139 337 140 
<< pdiffusion >>
rect 337 139 338 140 
<< pdiffusion >>
rect 338 139 339 140 
<< pdiffusion >>
rect 339 139 340 140 
<< pdiffusion >>
rect 340 139 341 140 
<< pdiffusion >>
rect 341 139 342 140 
<< m1 >>
rect 343 139 344 140 
<< m2 >>
rect 343 139 344 140 
<< m1 >>
rect 345 139 346 140 
<< m1 >>
rect 10 140 11 141 
<< pdiffusion >>
rect 12 140 13 141 
<< pdiffusion >>
rect 13 140 14 141 
<< pdiffusion >>
rect 14 140 15 141 
<< pdiffusion >>
rect 15 140 16 141 
<< pdiffusion >>
rect 16 140 17 141 
<< pdiffusion >>
rect 17 140 18 141 
<< m1 >>
rect 19 140 20 141 
<< m1 >>
rect 21 140 22 141 
<< m1 >>
rect 23 140 24 141 
<< m2 >>
rect 27 140 28 141 
<< m1 >>
rect 28 140 29 141 
<< pdiffusion >>
rect 30 140 31 141 
<< pdiffusion >>
rect 31 140 32 141 
<< pdiffusion >>
rect 32 140 33 141 
<< pdiffusion >>
rect 33 140 34 141 
<< pdiffusion >>
rect 34 140 35 141 
<< pdiffusion >>
rect 35 140 36 141 
<< m1 >>
rect 37 140 38 141 
<< m2 >>
rect 38 140 39 141 
<< m1 >>
rect 42 140 43 141 
<< m1 >>
rect 46 140 47 141 
<< pdiffusion >>
rect 48 140 49 141 
<< pdiffusion >>
rect 49 140 50 141 
<< pdiffusion >>
rect 50 140 51 141 
<< pdiffusion >>
rect 51 140 52 141 
<< pdiffusion >>
rect 52 140 53 141 
<< pdiffusion >>
rect 53 140 54 141 
<< m1 >>
rect 58 140 59 141 
<< m2 >>
rect 59 140 60 141 
<< m2 >>
rect 61 140 62 141 
<< m1 >>
rect 62 140 63 141 
<< m1 >>
rect 64 140 65 141 
<< pdiffusion >>
rect 66 140 67 141 
<< pdiffusion >>
rect 67 140 68 141 
<< pdiffusion >>
rect 68 140 69 141 
<< pdiffusion >>
rect 69 140 70 141 
<< pdiffusion >>
rect 70 140 71 141 
<< pdiffusion >>
rect 71 140 72 141 
<< m1 >>
rect 78 140 79 141 
<< m1 >>
rect 82 140 83 141 
<< pdiffusion >>
rect 84 140 85 141 
<< pdiffusion >>
rect 85 140 86 141 
<< pdiffusion >>
rect 86 140 87 141 
<< pdiffusion >>
rect 87 140 88 141 
<< pdiffusion >>
rect 88 140 89 141 
<< pdiffusion >>
rect 89 140 90 141 
<< m1 >>
rect 91 140 92 141 
<< m2 >>
rect 92 140 93 141 
<< pdiffusion >>
rect 102 140 103 141 
<< pdiffusion >>
rect 103 140 104 141 
<< pdiffusion >>
rect 104 140 105 141 
<< pdiffusion >>
rect 105 140 106 141 
<< pdiffusion >>
rect 106 140 107 141 
<< pdiffusion >>
rect 107 140 108 141 
<< m1 >>
rect 109 140 110 141 
<< pdiffusion >>
rect 120 140 121 141 
<< pdiffusion >>
rect 121 140 122 141 
<< pdiffusion >>
rect 122 140 123 141 
<< pdiffusion >>
rect 123 140 124 141 
<< pdiffusion >>
rect 124 140 125 141 
<< pdiffusion >>
rect 125 140 126 141 
<< m1 >>
rect 130 140 131 141 
<< m1 >>
rect 132 140 133 141 
<< m1 >>
rect 136 140 137 141 
<< m2 >>
rect 136 140 137 141 
<< pdiffusion >>
rect 138 140 139 141 
<< pdiffusion >>
rect 139 140 140 141 
<< pdiffusion >>
rect 140 140 141 141 
<< pdiffusion >>
rect 141 140 142 141 
<< pdiffusion >>
rect 142 140 143 141 
<< pdiffusion >>
rect 143 140 144 141 
<< m1 >>
rect 145 140 146 141 
<< m1 >>
rect 147 140 148 141 
<< m2 >>
rect 153 140 154 141 
<< m1 >>
rect 154 140 155 141 
<< pdiffusion >>
rect 156 140 157 141 
<< pdiffusion >>
rect 157 140 158 141 
<< pdiffusion >>
rect 158 140 159 141 
<< pdiffusion >>
rect 159 140 160 141 
<< pdiffusion >>
rect 160 140 161 141 
<< pdiffusion >>
rect 161 140 162 141 
<< m1 >>
rect 163 140 164 141 
<< m2 >>
rect 164 140 165 141 
<< m1 >>
rect 170 140 171 141 
<< m1 >>
rect 172 140 173 141 
<< pdiffusion >>
rect 174 140 175 141 
<< pdiffusion >>
rect 175 140 176 141 
<< pdiffusion >>
rect 176 140 177 141 
<< pdiffusion >>
rect 177 140 178 141 
<< pdiffusion >>
rect 178 140 179 141 
<< pdiffusion >>
rect 179 140 180 141 
<< m1 >>
rect 181 140 182 141 
<< m1 >>
rect 184 140 185 141 
<< m1 >>
rect 188 140 189 141 
<< pdiffusion >>
rect 192 140 193 141 
<< pdiffusion >>
rect 193 140 194 141 
<< pdiffusion >>
rect 194 140 195 141 
<< pdiffusion >>
rect 195 140 196 141 
<< pdiffusion >>
rect 196 140 197 141 
<< pdiffusion >>
rect 197 140 198 141 
<< m1 >>
rect 199 140 200 141 
<< m1 >>
rect 201 140 202 141 
<< m1 >>
rect 205 140 206 141 
<< pdiffusion >>
rect 210 140 211 141 
<< pdiffusion >>
rect 211 140 212 141 
<< pdiffusion >>
rect 212 140 213 141 
<< pdiffusion >>
rect 213 140 214 141 
<< pdiffusion >>
rect 214 140 215 141 
<< pdiffusion >>
rect 215 140 216 141 
<< m1 >>
rect 226 140 227 141 
<< m2 >>
rect 226 140 227 141 
<< pdiffusion >>
rect 228 140 229 141 
<< pdiffusion >>
rect 229 140 230 141 
<< pdiffusion >>
rect 230 140 231 141 
<< pdiffusion >>
rect 231 140 232 141 
<< pdiffusion >>
rect 232 140 233 141 
<< pdiffusion >>
rect 233 140 234 141 
<< m1 >>
rect 235 140 236 141 
<< m1 >>
rect 237 140 238 141 
<< m2 >>
rect 238 140 239 141 
<< m1 >>
rect 240 140 241 141 
<< pdiffusion >>
rect 246 140 247 141 
<< pdiffusion >>
rect 247 140 248 141 
<< pdiffusion >>
rect 248 140 249 141 
<< pdiffusion >>
rect 249 140 250 141 
<< pdiffusion >>
rect 250 140 251 141 
<< pdiffusion >>
rect 251 140 252 141 
<< m1 >>
rect 253 140 254 141 
<< m1 >>
rect 255 140 256 141 
<< m1 >>
rect 260 140 261 141 
<< m1 >>
rect 262 140 263 141 
<< pdiffusion >>
rect 264 140 265 141 
<< pdiffusion >>
rect 265 140 266 141 
<< pdiffusion >>
rect 266 140 267 141 
<< pdiffusion >>
rect 267 140 268 141 
<< pdiffusion >>
rect 268 140 269 141 
<< pdiffusion >>
rect 269 140 270 141 
<< m1 >>
rect 272 140 273 141 
<< m1 >>
rect 274 140 275 141 
<< m1 >>
rect 276 140 277 141 
<< m2 >>
rect 277 140 278 141 
<< m1 >>
rect 280 140 281 141 
<< pdiffusion >>
rect 282 140 283 141 
<< pdiffusion >>
rect 283 140 284 141 
<< pdiffusion >>
rect 284 140 285 141 
<< pdiffusion >>
rect 285 140 286 141 
<< pdiffusion >>
rect 286 140 287 141 
<< pdiffusion >>
rect 287 140 288 141 
<< m1 >>
rect 289 140 290 141 
<< m1 >>
rect 296 140 297 141 
<< m1 >>
rect 298 140 299 141 
<< pdiffusion >>
rect 300 140 301 141 
<< pdiffusion >>
rect 301 140 302 141 
<< pdiffusion >>
rect 302 140 303 141 
<< pdiffusion >>
rect 303 140 304 141 
<< pdiffusion >>
rect 304 140 305 141 
<< pdiffusion >>
rect 305 140 306 141 
<< m1 >>
rect 307 140 308 141 
<< m2 >>
rect 308 140 309 141 
<< pdiffusion >>
rect 318 140 319 141 
<< pdiffusion >>
rect 319 140 320 141 
<< pdiffusion >>
rect 320 140 321 141 
<< pdiffusion >>
rect 321 140 322 141 
<< pdiffusion >>
rect 322 140 323 141 
<< pdiffusion >>
rect 323 140 324 141 
<< m1 >>
rect 325 140 326 141 
<< m1 >>
rect 327 140 328 141 
<< m1 >>
rect 329 140 330 141 
<< pdiffusion >>
rect 336 140 337 141 
<< pdiffusion >>
rect 337 140 338 141 
<< pdiffusion >>
rect 338 140 339 141 
<< pdiffusion >>
rect 339 140 340 141 
<< pdiffusion >>
rect 340 140 341 141 
<< pdiffusion >>
rect 341 140 342 141 
<< m1 >>
rect 343 140 344 141 
<< m2 >>
rect 343 140 344 141 
<< m1 >>
rect 345 140 346 141 
<< m1 >>
rect 10 141 11 142 
<< pdiffusion >>
rect 12 141 13 142 
<< pdiffusion >>
rect 13 141 14 142 
<< pdiffusion >>
rect 14 141 15 142 
<< pdiffusion >>
rect 15 141 16 142 
<< pdiffusion >>
rect 16 141 17 142 
<< pdiffusion >>
rect 17 141 18 142 
<< m1 >>
rect 19 141 20 142 
<< m1 >>
rect 21 141 22 142 
<< m1 >>
rect 23 141 24 142 
<< m2 >>
rect 27 141 28 142 
<< m1 >>
rect 28 141 29 142 
<< pdiffusion >>
rect 30 141 31 142 
<< pdiffusion >>
rect 31 141 32 142 
<< pdiffusion >>
rect 32 141 33 142 
<< pdiffusion >>
rect 33 141 34 142 
<< pdiffusion >>
rect 34 141 35 142 
<< pdiffusion >>
rect 35 141 36 142 
<< m1 >>
rect 37 141 38 142 
<< m2 >>
rect 38 141 39 142 
<< m1 >>
rect 42 141 43 142 
<< m1 >>
rect 46 141 47 142 
<< pdiffusion >>
rect 48 141 49 142 
<< pdiffusion >>
rect 49 141 50 142 
<< pdiffusion >>
rect 50 141 51 142 
<< pdiffusion >>
rect 51 141 52 142 
<< pdiffusion >>
rect 52 141 53 142 
<< pdiffusion >>
rect 53 141 54 142 
<< m1 >>
rect 58 141 59 142 
<< m2 >>
rect 59 141 60 142 
<< m2 >>
rect 61 141 62 142 
<< m1 >>
rect 62 141 63 142 
<< m1 >>
rect 64 141 65 142 
<< pdiffusion >>
rect 66 141 67 142 
<< pdiffusion >>
rect 67 141 68 142 
<< pdiffusion >>
rect 68 141 69 142 
<< pdiffusion >>
rect 69 141 70 142 
<< pdiffusion >>
rect 70 141 71 142 
<< pdiffusion >>
rect 71 141 72 142 
<< m1 >>
rect 78 141 79 142 
<< m1 >>
rect 82 141 83 142 
<< pdiffusion >>
rect 84 141 85 142 
<< pdiffusion >>
rect 85 141 86 142 
<< pdiffusion >>
rect 86 141 87 142 
<< pdiffusion >>
rect 87 141 88 142 
<< pdiffusion >>
rect 88 141 89 142 
<< pdiffusion >>
rect 89 141 90 142 
<< m1 >>
rect 91 141 92 142 
<< m2 >>
rect 92 141 93 142 
<< pdiffusion >>
rect 102 141 103 142 
<< pdiffusion >>
rect 103 141 104 142 
<< pdiffusion >>
rect 104 141 105 142 
<< pdiffusion >>
rect 105 141 106 142 
<< pdiffusion >>
rect 106 141 107 142 
<< pdiffusion >>
rect 107 141 108 142 
<< m1 >>
rect 109 141 110 142 
<< pdiffusion >>
rect 120 141 121 142 
<< pdiffusion >>
rect 121 141 122 142 
<< pdiffusion >>
rect 122 141 123 142 
<< pdiffusion >>
rect 123 141 124 142 
<< pdiffusion >>
rect 124 141 125 142 
<< pdiffusion >>
rect 125 141 126 142 
<< m1 >>
rect 130 141 131 142 
<< m1 >>
rect 132 141 133 142 
<< m1 >>
rect 136 141 137 142 
<< m2 >>
rect 136 141 137 142 
<< pdiffusion >>
rect 138 141 139 142 
<< pdiffusion >>
rect 139 141 140 142 
<< pdiffusion >>
rect 140 141 141 142 
<< pdiffusion >>
rect 141 141 142 142 
<< pdiffusion >>
rect 142 141 143 142 
<< pdiffusion >>
rect 143 141 144 142 
<< m1 >>
rect 145 141 146 142 
<< m1 >>
rect 147 141 148 142 
<< m2 >>
rect 153 141 154 142 
<< m1 >>
rect 154 141 155 142 
<< pdiffusion >>
rect 156 141 157 142 
<< pdiffusion >>
rect 157 141 158 142 
<< pdiffusion >>
rect 158 141 159 142 
<< pdiffusion >>
rect 159 141 160 142 
<< pdiffusion >>
rect 160 141 161 142 
<< pdiffusion >>
rect 161 141 162 142 
<< m1 >>
rect 163 141 164 142 
<< m2 >>
rect 164 141 165 142 
<< m1 >>
rect 170 141 171 142 
<< m1 >>
rect 172 141 173 142 
<< pdiffusion >>
rect 174 141 175 142 
<< pdiffusion >>
rect 175 141 176 142 
<< pdiffusion >>
rect 176 141 177 142 
<< pdiffusion >>
rect 177 141 178 142 
<< pdiffusion >>
rect 178 141 179 142 
<< pdiffusion >>
rect 179 141 180 142 
<< m1 >>
rect 181 141 182 142 
<< m1 >>
rect 184 141 185 142 
<< m1 >>
rect 188 141 189 142 
<< pdiffusion >>
rect 192 141 193 142 
<< pdiffusion >>
rect 193 141 194 142 
<< pdiffusion >>
rect 194 141 195 142 
<< pdiffusion >>
rect 195 141 196 142 
<< pdiffusion >>
rect 196 141 197 142 
<< pdiffusion >>
rect 197 141 198 142 
<< m1 >>
rect 199 141 200 142 
<< m1 >>
rect 201 141 202 142 
<< m1 >>
rect 205 141 206 142 
<< pdiffusion >>
rect 210 141 211 142 
<< pdiffusion >>
rect 211 141 212 142 
<< pdiffusion >>
rect 212 141 213 142 
<< pdiffusion >>
rect 213 141 214 142 
<< pdiffusion >>
rect 214 141 215 142 
<< pdiffusion >>
rect 215 141 216 142 
<< m1 >>
rect 226 141 227 142 
<< m2 >>
rect 226 141 227 142 
<< pdiffusion >>
rect 228 141 229 142 
<< pdiffusion >>
rect 229 141 230 142 
<< pdiffusion >>
rect 230 141 231 142 
<< pdiffusion >>
rect 231 141 232 142 
<< pdiffusion >>
rect 232 141 233 142 
<< pdiffusion >>
rect 233 141 234 142 
<< m1 >>
rect 235 141 236 142 
<< m1 >>
rect 237 141 238 142 
<< m2 >>
rect 238 141 239 142 
<< m1 >>
rect 240 141 241 142 
<< pdiffusion >>
rect 246 141 247 142 
<< pdiffusion >>
rect 247 141 248 142 
<< pdiffusion >>
rect 248 141 249 142 
<< pdiffusion >>
rect 249 141 250 142 
<< pdiffusion >>
rect 250 141 251 142 
<< pdiffusion >>
rect 251 141 252 142 
<< m1 >>
rect 253 141 254 142 
<< m1 >>
rect 255 141 256 142 
<< m1 >>
rect 260 141 261 142 
<< m1 >>
rect 262 141 263 142 
<< pdiffusion >>
rect 264 141 265 142 
<< pdiffusion >>
rect 265 141 266 142 
<< pdiffusion >>
rect 266 141 267 142 
<< pdiffusion >>
rect 267 141 268 142 
<< pdiffusion >>
rect 268 141 269 142 
<< pdiffusion >>
rect 269 141 270 142 
<< m1 >>
rect 272 141 273 142 
<< m1 >>
rect 274 141 275 142 
<< m1 >>
rect 276 141 277 142 
<< m2 >>
rect 277 141 278 142 
<< m1 >>
rect 280 141 281 142 
<< pdiffusion >>
rect 282 141 283 142 
<< pdiffusion >>
rect 283 141 284 142 
<< pdiffusion >>
rect 284 141 285 142 
<< pdiffusion >>
rect 285 141 286 142 
<< pdiffusion >>
rect 286 141 287 142 
<< pdiffusion >>
rect 287 141 288 142 
<< m1 >>
rect 289 141 290 142 
<< m1 >>
rect 296 141 297 142 
<< m1 >>
rect 298 141 299 142 
<< pdiffusion >>
rect 300 141 301 142 
<< pdiffusion >>
rect 301 141 302 142 
<< pdiffusion >>
rect 302 141 303 142 
<< pdiffusion >>
rect 303 141 304 142 
<< pdiffusion >>
rect 304 141 305 142 
<< pdiffusion >>
rect 305 141 306 142 
<< m1 >>
rect 307 141 308 142 
<< m2 >>
rect 308 141 309 142 
<< pdiffusion >>
rect 318 141 319 142 
<< pdiffusion >>
rect 319 141 320 142 
<< pdiffusion >>
rect 320 141 321 142 
<< pdiffusion >>
rect 321 141 322 142 
<< pdiffusion >>
rect 322 141 323 142 
<< pdiffusion >>
rect 323 141 324 142 
<< m1 >>
rect 325 141 326 142 
<< m1 >>
rect 327 141 328 142 
<< m1 >>
rect 329 141 330 142 
<< pdiffusion >>
rect 336 141 337 142 
<< pdiffusion >>
rect 337 141 338 142 
<< pdiffusion >>
rect 338 141 339 142 
<< pdiffusion >>
rect 339 141 340 142 
<< pdiffusion >>
rect 340 141 341 142 
<< pdiffusion >>
rect 341 141 342 142 
<< m1 >>
rect 343 141 344 142 
<< m2 >>
rect 343 141 344 142 
<< m1 >>
rect 345 141 346 142 
<< m1 >>
rect 10 142 11 143 
<< pdiffusion >>
rect 12 142 13 143 
<< pdiffusion >>
rect 13 142 14 143 
<< pdiffusion >>
rect 14 142 15 143 
<< pdiffusion >>
rect 15 142 16 143 
<< pdiffusion >>
rect 16 142 17 143 
<< pdiffusion >>
rect 17 142 18 143 
<< m1 >>
rect 19 142 20 143 
<< m1 >>
rect 21 142 22 143 
<< m1 >>
rect 23 142 24 143 
<< m2 >>
rect 27 142 28 143 
<< m1 >>
rect 28 142 29 143 
<< pdiffusion >>
rect 30 142 31 143 
<< pdiffusion >>
rect 31 142 32 143 
<< pdiffusion >>
rect 32 142 33 143 
<< pdiffusion >>
rect 33 142 34 143 
<< pdiffusion >>
rect 34 142 35 143 
<< pdiffusion >>
rect 35 142 36 143 
<< m1 >>
rect 37 142 38 143 
<< m2 >>
rect 38 142 39 143 
<< m1 >>
rect 42 142 43 143 
<< m1 >>
rect 46 142 47 143 
<< pdiffusion >>
rect 48 142 49 143 
<< pdiffusion >>
rect 49 142 50 143 
<< pdiffusion >>
rect 50 142 51 143 
<< pdiffusion >>
rect 51 142 52 143 
<< pdiffusion >>
rect 52 142 53 143 
<< pdiffusion >>
rect 53 142 54 143 
<< m1 >>
rect 58 142 59 143 
<< m2 >>
rect 59 142 60 143 
<< m2 >>
rect 61 142 62 143 
<< m1 >>
rect 62 142 63 143 
<< m1 >>
rect 64 142 65 143 
<< pdiffusion >>
rect 66 142 67 143 
<< pdiffusion >>
rect 67 142 68 143 
<< pdiffusion >>
rect 68 142 69 143 
<< pdiffusion >>
rect 69 142 70 143 
<< pdiffusion >>
rect 70 142 71 143 
<< pdiffusion >>
rect 71 142 72 143 
<< m1 >>
rect 78 142 79 143 
<< m1 >>
rect 82 142 83 143 
<< pdiffusion >>
rect 84 142 85 143 
<< pdiffusion >>
rect 85 142 86 143 
<< pdiffusion >>
rect 86 142 87 143 
<< pdiffusion >>
rect 87 142 88 143 
<< pdiffusion >>
rect 88 142 89 143 
<< pdiffusion >>
rect 89 142 90 143 
<< m1 >>
rect 91 142 92 143 
<< m2 >>
rect 92 142 93 143 
<< pdiffusion >>
rect 102 142 103 143 
<< pdiffusion >>
rect 103 142 104 143 
<< pdiffusion >>
rect 104 142 105 143 
<< pdiffusion >>
rect 105 142 106 143 
<< pdiffusion >>
rect 106 142 107 143 
<< pdiffusion >>
rect 107 142 108 143 
<< m1 >>
rect 109 142 110 143 
<< pdiffusion >>
rect 120 142 121 143 
<< pdiffusion >>
rect 121 142 122 143 
<< pdiffusion >>
rect 122 142 123 143 
<< pdiffusion >>
rect 123 142 124 143 
<< pdiffusion >>
rect 124 142 125 143 
<< pdiffusion >>
rect 125 142 126 143 
<< m1 >>
rect 130 142 131 143 
<< m1 >>
rect 132 142 133 143 
<< m1 >>
rect 136 142 137 143 
<< m2 >>
rect 136 142 137 143 
<< pdiffusion >>
rect 138 142 139 143 
<< pdiffusion >>
rect 139 142 140 143 
<< pdiffusion >>
rect 140 142 141 143 
<< pdiffusion >>
rect 141 142 142 143 
<< pdiffusion >>
rect 142 142 143 143 
<< pdiffusion >>
rect 143 142 144 143 
<< m1 >>
rect 145 142 146 143 
<< m1 >>
rect 147 142 148 143 
<< m2 >>
rect 153 142 154 143 
<< m1 >>
rect 154 142 155 143 
<< pdiffusion >>
rect 156 142 157 143 
<< pdiffusion >>
rect 157 142 158 143 
<< pdiffusion >>
rect 158 142 159 143 
<< pdiffusion >>
rect 159 142 160 143 
<< pdiffusion >>
rect 160 142 161 143 
<< pdiffusion >>
rect 161 142 162 143 
<< m1 >>
rect 163 142 164 143 
<< m2 >>
rect 164 142 165 143 
<< m1 >>
rect 170 142 171 143 
<< m1 >>
rect 172 142 173 143 
<< pdiffusion >>
rect 174 142 175 143 
<< pdiffusion >>
rect 175 142 176 143 
<< pdiffusion >>
rect 176 142 177 143 
<< pdiffusion >>
rect 177 142 178 143 
<< pdiffusion >>
rect 178 142 179 143 
<< pdiffusion >>
rect 179 142 180 143 
<< m1 >>
rect 181 142 182 143 
<< m1 >>
rect 184 142 185 143 
<< m1 >>
rect 188 142 189 143 
<< pdiffusion >>
rect 192 142 193 143 
<< pdiffusion >>
rect 193 142 194 143 
<< pdiffusion >>
rect 194 142 195 143 
<< pdiffusion >>
rect 195 142 196 143 
<< pdiffusion >>
rect 196 142 197 143 
<< pdiffusion >>
rect 197 142 198 143 
<< m1 >>
rect 199 142 200 143 
<< m1 >>
rect 201 142 202 143 
<< m1 >>
rect 205 142 206 143 
<< pdiffusion >>
rect 210 142 211 143 
<< pdiffusion >>
rect 211 142 212 143 
<< pdiffusion >>
rect 212 142 213 143 
<< pdiffusion >>
rect 213 142 214 143 
<< pdiffusion >>
rect 214 142 215 143 
<< pdiffusion >>
rect 215 142 216 143 
<< m1 >>
rect 226 142 227 143 
<< m2 >>
rect 226 142 227 143 
<< pdiffusion >>
rect 228 142 229 143 
<< pdiffusion >>
rect 229 142 230 143 
<< pdiffusion >>
rect 230 142 231 143 
<< pdiffusion >>
rect 231 142 232 143 
<< pdiffusion >>
rect 232 142 233 143 
<< pdiffusion >>
rect 233 142 234 143 
<< m1 >>
rect 235 142 236 143 
<< m1 >>
rect 237 142 238 143 
<< m2 >>
rect 238 142 239 143 
<< m1 >>
rect 240 142 241 143 
<< pdiffusion >>
rect 246 142 247 143 
<< pdiffusion >>
rect 247 142 248 143 
<< pdiffusion >>
rect 248 142 249 143 
<< pdiffusion >>
rect 249 142 250 143 
<< pdiffusion >>
rect 250 142 251 143 
<< pdiffusion >>
rect 251 142 252 143 
<< m1 >>
rect 253 142 254 143 
<< m1 >>
rect 255 142 256 143 
<< m1 >>
rect 260 142 261 143 
<< m1 >>
rect 262 142 263 143 
<< pdiffusion >>
rect 264 142 265 143 
<< pdiffusion >>
rect 265 142 266 143 
<< pdiffusion >>
rect 266 142 267 143 
<< pdiffusion >>
rect 267 142 268 143 
<< pdiffusion >>
rect 268 142 269 143 
<< pdiffusion >>
rect 269 142 270 143 
<< m1 >>
rect 272 142 273 143 
<< m1 >>
rect 274 142 275 143 
<< m1 >>
rect 276 142 277 143 
<< m2 >>
rect 277 142 278 143 
<< m1 >>
rect 280 142 281 143 
<< pdiffusion >>
rect 282 142 283 143 
<< pdiffusion >>
rect 283 142 284 143 
<< pdiffusion >>
rect 284 142 285 143 
<< pdiffusion >>
rect 285 142 286 143 
<< pdiffusion >>
rect 286 142 287 143 
<< pdiffusion >>
rect 287 142 288 143 
<< m1 >>
rect 289 142 290 143 
<< m1 >>
rect 296 142 297 143 
<< m1 >>
rect 298 142 299 143 
<< pdiffusion >>
rect 300 142 301 143 
<< pdiffusion >>
rect 301 142 302 143 
<< pdiffusion >>
rect 302 142 303 143 
<< pdiffusion >>
rect 303 142 304 143 
<< pdiffusion >>
rect 304 142 305 143 
<< pdiffusion >>
rect 305 142 306 143 
<< m1 >>
rect 307 142 308 143 
<< m2 >>
rect 308 142 309 143 
<< pdiffusion >>
rect 318 142 319 143 
<< pdiffusion >>
rect 319 142 320 143 
<< pdiffusion >>
rect 320 142 321 143 
<< pdiffusion >>
rect 321 142 322 143 
<< pdiffusion >>
rect 322 142 323 143 
<< pdiffusion >>
rect 323 142 324 143 
<< m1 >>
rect 325 142 326 143 
<< m1 >>
rect 327 142 328 143 
<< m1 >>
rect 329 142 330 143 
<< pdiffusion >>
rect 336 142 337 143 
<< pdiffusion >>
rect 337 142 338 143 
<< pdiffusion >>
rect 338 142 339 143 
<< pdiffusion >>
rect 339 142 340 143 
<< pdiffusion >>
rect 340 142 341 143 
<< pdiffusion >>
rect 341 142 342 143 
<< m1 >>
rect 343 142 344 143 
<< m2 >>
rect 343 142 344 143 
<< m1 >>
rect 345 142 346 143 
<< m1 >>
rect 10 143 11 144 
<< pdiffusion >>
rect 12 143 13 144 
<< pdiffusion >>
rect 13 143 14 144 
<< pdiffusion >>
rect 14 143 15 144 
<< pdiffusion >>
rect 15 143 16 144 
<< m1 >>
rect 16 143 17 144 
<< pdiffusion >>
rect 16 143 17 144 
<< pdiffusion >>
rect 17 143 18 144 
<< m1 >>
rect 19 143 20 144 
<< m1 >>
rect 21 143 22 144 
<< m1 >>
rect 23 143 24 144 
<< m2 >>
rect 27 143 28 144 
<< m1 >>
rect 28 143 29 144 
<< pdiffusion >>
rect 30 143 31 144 
<< pdiffusion >>
rect 31 143 32 144 
<< pdiffusion >>
rect 32 143 33 144 
<< pdiffusion >>
rect 33 143 34 144 
<< pdiffusion >>
rect 34 143 35 144 
<< pdiffusion >>
rect 35 143 36 144 
<< m1 >>
rect 37 143 38 144 
<< m2 >>
rect 38 143 39 144 
<< m1 >>
rect 42 143 43 144 
<< m1 >>
rect 46 143 47 144 
<< pdiffusion >>
rect 48 143 49 144 
<< pdiffusion >>
rect 49 143 50 144 
<< pdiffusion >>
rect 50 143 51 144 
<< pdiffusion >>
rect 51 143 52 144 
<< pdiffusion >>
rect 52 143 53 144 
<< pdiffusion >>
rect 53 143 54 144 
<< m1 >>
rect 58 143 59 144 
<< m2 >>
rect 59 143 60 144 
<< m2 >>
rect 61 143 62 144 
<< m1 >>
rect 62 143 63 144 
<< m1 >>
rect 64 143 65 144 
<< pdiffusion >>
rect 66 143 67 144 
<< pdiffusion >>
rect 67 143 68 144 
<< pdiffusion >>
rect 68 143 69 144 
<< pdiffusion >>
rect 69 143 70 144 
<< pdiffusion >>
rect 70 143 71 144 
<< pdiffusion >>
rect 71 143 72 144 
<< m1 >>
rect 78 143 79 144 
<< m1 >>
rect 82 143 83 144 
<< pdiffusion >>
rect 84 143 85 144 
<< pdiffusion >>
rect 85 143 86 144 
<< pdiffusion >>
rect 86 143 87 144 
<< pdiffusion >>
rect 87 143 88 144 
<< pdiffusion >>
rect 88 143 89 144 
<< pdiffusion >>
rect 89 143 90 144 
<< m1 >>
rect 91 143 92 144 
<< m2 >>
rect 92 143 93 144 
<< pdiffusion >>
rect 102 143 103 144 
<< pdiffusion >>
rect 103 143 104 144 
<< pdiffusion >>
rect 104 143 105 144 
<< pdiffusion >>
rect 105 143 106 144 
<< pdiffusion >>
rect 106 143 107 144 
<< pdiffusion >>
rect 107 143 108 144 
<< m1 >>
rect 109 143 110 144 
<< pdiffusion >>
rect 120 143 121 144 
<< pdiffusion >>
rect 121 143 122 144 
<< pdiffusion >>
rect 122 143 123 144 
<< pdiffusion >>
rect 123 143 124 144 
<< pdiffusion >>
rect 124 143 125 144 
<< pdiffusion >>
rect 125 143 126 144 
<< m1 >>
rect 130 143 131 144 
<< m1 >>
rect 132 143 133 144 
<< m1 >>
rect 136 143 137 144 
<< m2 >>
rect 136 143 137 144 
<< pdiffusion >>
rect 138 143 139 144 
<< pdiffusion >>
rect 139 143 140 144 
<< pdiffusion >>
rect 140 143 141 144 
<< pdiffusion >>
rect 141 143 142 144 
<< pdiffusion >>
rect 142 143 143 144 
<< pdiffusion >>
rect 143 143 144 144 
<< m1 >>
rect 145 143 146 144 
<< m1 >>
rect 147 143 148 144 
<< m2 >>
rect 153 143 154 144 
<< m1 >>
rect 154 143 155 144 
<< pdiffusion >>
rect 156 143 157 144 
<< pdiffusion >>
rect 157 143 158 144 
<< pdiffusion >>
rect 158 143 159 144 
<< pdiffusion >>
rect 159 143 160 144 
<< pdiffusion >>
rect 160 143 161 144 
<< pdiffusion >>
rect 161 143 162 144 
<< m1 >>
rect 163 143 164 144 
<< m2 >>
rect 164 143 165 144 
<< m1 >>
rect 170 143 171 144 
<< m1 >>
rect 172 143 173 144 
<< pdiffusion >>
rect 174 143 175 144 
<< pdiffusion >>
rect 175 143 176 144 
<< pdiffusion >>
rect 176 143 177 144 
<< pdiffusion >>
rect 177 143 178 144 
<< m1 >>
rect 178 143 179 144 
<< pdiffusion >>
rect 178 143 179 144 
<< pdiffusion >>
rect 179 143 180 144 
<< m1 >>
rect 181 143 182 144 
<< m1 >>
rect 184 143 185 144 
<< m2 >>
rect 184 143 185 144 
<< m2c >>
rect 184 143 185 144 
<< m1 >>
rect 184 143 185 144 
<< m2 >>
rect 184 143 185 144 
<< m1 >>
rect 188 143 189 144 
<< pdiffusion >>
rect 192 143 193 144 
<< pdiffusion >>
rect 193 143 194 144 
<< pdiffusion >>
rect 194 143 195 144 
<< pdiffusion >>
rect 195 143 196 144 
<< m1 >>
rect 196 143 197 144 
<< pdiffusion >>
rect 196 143 197 144 
<< pdiffusion >>
rect 197 143 198 144 
<< m1 >>
rect 199 143 200 144 
<< m1 >>
rect 201 143 202 144 
<< m1 >>
rect 205 143 206 144 
<< pdiffusion >>
rect 210 143 211 144 
<< m1 >>
rect 211 143 212 144 
<< pdiffusion >>
rect 211 143 212 144 
<< pdiffusion >>
rect 212 143 213 144 
<< pdiffusion >>
rect 213 143 214 144 
<< pdiffusion >>
rect 214 143 215 144 
<< pdiffusion >>
rect 215 143 216 144 
<< m1 >>
rect 226 143 227 144 
<< m2 >>
rect 226 143 227 144 
<< pdiffusion >>
rect 228 143 229 144 
<< pdiffusion >>
rect 229 143 230 144 
<< pdiffusion >>
rect 230 143 231 144 
<< pdiffusion >>
rect 231 143 232 144 
<< m1 >>
rect 232 143 233 144 
<< pdiffusion >>
rect 232 143 233 144 
<< pdiffusion >>
rect 233 143 234 144 
<< m1 >>
rect 235 143 236 144 
<< m1 >>
rect 237 143 238 144 
<< m2 >>
rect 238 143 239 144 
<< m1 >>
rect 240 143 241 144 
<< pdiffusion >>
rect 246 143 247 144 
<< pdiffusion >>
rect 247 143 248 144 
<< pdiffusion >>
rect 248 143 249 144 
<< pdiffusion >>
rect 249 143 250 144 
<< pdiffusion >>
rect 250 143 251 144 
<< pdiffusion >>
rect 251 143 252 144 
<< m1 >>
rect 253 143 254 144 
<< m1 >>
rect 255 143 256 144 
<< m1 >>
rect 260 143 261 144 
<< m1 >>
rect 262 143 263 144 
<< pdiffusion >>
rect 264 143 265 144 
<< m1 >>
rect 265 143 266 144 
<< pdiffusion >>
rect 265 143 266 144 
<< pdiffusion >>
rect 266 143 267 144 
<< pdiffusion >>
rect 267 143 268 144 
<< pdiffusion >>
rect 268 143 269 144 
<< pdiffusion >>
rect 269 143 270 144 
<< m1 >>
rect 272 143 273 144 
<< m1 >>
rect 274 143 275 144 
<< m1 >>
rect 276 143 277 144 
<< m2 >>
rect 277 143 278 144 
<< m1 >>
rect 280 143 281 144 
<< pdiffusion >>
rect 282 143 283 144 
<< pdiffusion >>
rect 283 143 284 144 
<< pdiffusion >>
rect 284 143 285 144 
<< pdiffusion >>
rect 285 143 286 144 
<< pdiffusion >>
rect 286 143 287 144 
<< pdiffusion >>
rect 287 143 288 144 
<< m1 >>
rect 289 143 290 144 
<< m1 >>
rect 296 143 297 144 
<< m1 >>
rect 298 143 299 144 
<< pdiffusion >>
rect 300 143 301 144 
<< pdiffusion >>
rect 301 143 302 144 
<< pdiffusion >>
rect 302 143 303 144 
<< pdiffusion >>
rect 303 143 304 144 
<< pdiffusion >>
rect 304 143 305 144 
<< pdiffusion >>
rect 305 143 306 144 
<< m1 >>
rect 307 143 308 144 
<< m2 >>
rect 308 143 309 144 
<< pdiffusion >>
rect 318 143 319 144 
<< pdiffusion >>
rect 319 143 320 144 
<< pdiffusion >>
rect 320 143 321 144 
<< pdiffusion >>
rect 321 143 322 144 
<< pdiffusion >>
rect 322 143 323 144 
<< pdiffusion >>
rect 323 143 324 144 
<< m1 >>
rect 325 143 326 144 
<< m1 >>
rect 327 143 328 144 
<< m1 >>
rect 329 143 330 144 
<< pdiffusion >>
rect 336 143 337 144 
<< pdiffusion >>
rect 337 143 338 144 
<< pdiffusion >>
rect 338 143 339 144 
<< pdiffusion >>
rect 339 143 340 144 
<< pdiffusion >>
rect 340 143 341 144 
<< pdiffusion >>
rect 341 143 342 144 
<< m1 >>
rect 343 143 344 144 
<< m2 >>
rect 343 143 344 144 
<< m1 >>
rect 345 143 346 144 
<< m1 >>
rect 10 144 11 145 
<< m1 >>
rect 16 144 17 145 
<< m1 >>
rect 19 144 20 145 
<< m1 >>
rect 21 144 22 145 
<< m1 >>
rect 23 144 24 145 
<< m2 >>
rect 27 144 28 145 
<< m1 >>
rect 28 144 29 145 
<< m1 >>
rect 37 144 38 145 
<< m2 >>
rect 38 144 39 145 
<< m1 >>
rect 42 144 43 145 
<< m1 >>
rect 46 144 47 145 
<< m1 >>
rect 58 144 59 145 
<< m2 >>
rect 59 144 60 145 
<< m2 >>
rect 61 144 62 145 
<< m1 >>
rect 62 144 63 145 
<< m1 >>
rect 64 144 65 145 
<< m1 >>
rect 78 144 79 145 
<< m1 >>
rect 82 144 83 145 
<< m1 >>
rect 91 144 92 145 
<< m2 >>
rect 92 144 93 145 
<< m1 >>
rect 109 144 110 145 
<< m1 >>
rect 130 144 131 145 
<< m1 >>
rect 132 144 133 145 
<< m1 >>
rect 136 144 137 145 
<< m2 >>
rect 136 144 137 145 
<< m1 >>
rect 145 144 146 145 
<< m1 >>
rect 147 144 148 145 
<< m1 >>
rect 149 144 150 145 
<< m1 >>
rect 150 144 151 145 
<< m1 >>
rect 151 144 152 145 
<< m1 >>
rect 152 144 153 145 
<< m2 >>
rect 152 144 153 145 
<< m2c >>
rect 152 144 153 145 
<< m1 >>
rect 152 144 153 145 
<< m2 >>
rect 152 144 153 145 
<< m2 >>
rect 153 144 154 145 
<< m1 >>
rect 154 144 155 145 
<< m1 >>
rect 163 144 164 145 
<< m2 >>
rect 164 144 165 145 
<< m1 >>
rect 170 144 171 145 
<< m1 >>
rect 172 144 173 145 
<< m1 >>
rect 178 144 179 145 
<< m1 >>
rect 181 144 182 145 
<< m2 >>
rect 184 144 185 145 
<< m1 >>
rect 188 144 189 145 
<< m1 >>
rect 196 144 197 145 
<< m1 >>
rect 199 144 200 145 
<< m1 >>
rect 201 144 202 145 
<< m1 >>
rect 205 144 206 145 
<< m1 >>
rect 211 144 212 145 
<< m1 >>
rect 226 144 227 145 
<< m2 >>
rect 226 144 227 145 
<< m1 >>
rect 232 144 233 145 
<< m1 >>
rect 235 144 236 145 
<< m1 >>
rect 237 144 238 145 
<< m2 >>
rect 238 144 239 145 
<< m1 >>
rect 240 144 241 145 
<< m1 >>
rect 253 144 254 145 
<< m1 >>
rect 255 144 256 145 
<< m1 >>
rect 260 144 261 145 
<< m1 >>
rect 262 144 263 145 
<< m1 >>
rect 265 144 266 145 
<< m1 >>
rect 272 144 273 145 
<< m1 >>
rect 274 144 275 145 
<< m1 >>
rect 276 144 277 145 
<< m2 >>
rect 277 144 278 145 
<< m1 >>
rect 280 144 281 145 
<< m1 >>
rect 289 144 290 145 
<< m1 >>
rect 296 144 297 145 
<< m1 >>
rect 298 144 299 145 
<< m1 >>
rect 307 144 308 145 
<< m2 >>
rect 308 144 309 145 
<< m1 >>
rect 325 144 326 145 
<< m1 >>
rect 327 144 328 145 
<< m1 >>
rect 329 144 330 145 
<< m1 >>
rect 343 144 344 145 
<< m2 >>
rect 343 144 344 145 
<< m1 >>
rect 345 144 346 145 
<< m1 >>
rect 10 145 11 146 
<< m1 >>
rect 16 145 17 146 
<< m1 >>
rect 17 145 18 146 
<< m1 >>
rect 18 145 19 146 
<< m1 >>
rect 19 145 20 146 
<< m1 >>
rect 21 145 22 146 
<< m1 >>
rect 23 145 24 146 
<< m2 >>
rect 27 145 28 146 
<< m1 >>
rect 28 145 29 146 
<< m1 >>
rect 35 145 36 146 
<< m2 >>
rect 35 145 36 146 
<< m2c >>
rect 35 145 36 146 
<< m1 >>
rect 35 145 36 146 
<< m2 >>
rect 35 145 36 146 
<< m2 >>
rect 36 145 37 146 
<< m1 >>
rect 37 145 38 146 
<< m2 >>
rect 37 145 38 146 
<< m2 >>
rect 38 145 39 146 
<< m1 >>
rect 42 145 43 146 
<< m1 >>
rect 46 145 47 146 
<< m1 >>
rect 58 145 59 146 
<< m2 >>
rect 59 145 60 146 
<< m2 >>
rect 61 145 62 146 
<< m1 >>
rect 62 145 63 146 
<< m1 >>
rect 64 145 65 146 
<< m1 >>
rect 78 145 79 146 
<< m1 >>
rect 82 145 83 146 
<< m1 >>
rect 91 145 92 146 
<< m2 >>
rect 92 145 93 146 
<< m1 >>
rect 109 145 110 146 
<< m1 >>
rect 130 145 131 146 
<< m1 >>
rect 132 145 133 146 
<< m1 >>
rect 136 145 137 146 
<< m2 >>
rect 136 145 137 146 
<< m1 >>
rect 145 145 146 146 
<< m1 >>
rect 147 145 148 146 
<< m1 >>
rect 149 145 150 146 
<< m1 >>
rect 154 145 155 146 
<< m1 >>
rect 163 145 164 146 
<< m2 >>
rect 164 145 165 146 
<< m1 >>
rect 170 145 171 146 
<< m1 >>
rect 172 145 173 146 
<< m1 >>
rect 178 145 179 146 
<< m1 >>
rect 179 145 180 146 
<< m2 >>
rect 179 145 180 146 
<< m2c >>
rect 179 145 180 146 
<< m1 >>
rect 179 145 180 146 
<< m2 >>
rect 179 145 180 146 
<< m2 >>
rect 180 145 181 146 
<< m1 >>
rect 181 145 182 146 
<< m2 >>
rect 181 145 182 146 
<< m2 >>
rect 182 145 183 146 
<< m1 >>
rect 183 145 184 146 
<< m2 >>
rect 183 145 184 146 
<< m1 >>
rect 184 145 185 146 
<< m2 >>
rect 184 145 185 146 
<< m1 >>
rect 185 145 186 146 
<< m1 >>
rect 186 145 187 146 
<< m2 >>
rect 186 145 187 146 
<< m2c >>
rect 186 145 187 146 
<< m1 >>
rect 186 145 187 146 
<< m2 >>
rect 186 145 187 146 
<< m2 >>
rect 187 145 188 146 
<< m1 >>
rect 188 145 189 146 
<< m2 >>
rect 188 145 189 146 
<< m2 >>
rect 189 145 190 146 
<< m1 >>
rect 190 145 191 146 
<< m2 >>
rect 190 145 191 146 
<< m2c >>
rect 190 145 191 146 
<< m1 >>
rect 190 145 191 146 
<< m2 >>
rect 190 145 191 146 
<< m1 >>
rect 191 145 192 146 
<< m1 >>
rect 192 145 193 146 
<< m1 >>
rect 196 145 197 146 
<< m1 >>
rect 199 145 200 146 
<< m1 >>
rect 201 145 202 146 
<< m1 >>
rect 205 145 206 146 
<< m1 >>
rect 206 145 207 146 
<< m1 >>
rect 207 145 208 146 
<< m1 >>
rect 208 145 209 146 
<< m1 >>
rect 209 145 210 146 
<< m1 >>
rect 210 145 211 146 
<< m1 >>
rect 211 145 212 146 
<< m1 >>
rect 226 145 227 146 
<< m2 >>
rect 226 145 227 146 
<< m1 >>
rect 232 145 233 146 
<< m1 >>
rect 235 145 236 146 
<< m1 >>
rect 237 145 238 146 
<< m2 >>
rect 238 145 239 146 
<< m1 >>
rect 240 145 241 146 
<< m1 >>
rect 253 145 254 146 
<< m1 >>
rect 255 145 256 146 
<< m1 >>
rect 260 145 261 146 
<< m1 >>
rect 262 145 263 146 
<< m1 >>
rect 265 145 266 146 
<< m1 >>
rect 270 145 271 146 
<< m2 >>
rect 270 145 271 146 
<< m2c >>
rect 270 145 271 146 
<< m1 >>
rect 270 145 271 146 
<< m2 >>
rect 270 145 271 146 
<< m2 >>
rect 271 145 272 146 
<< m1 >>
rect 272 145 273 146 
<< m2 >>
rect 272 145 273 146 
<< m2 >>
rect 273 145 274 146 
<< m1 >>
rect 274 145 275 146 
<< m2 >>
rect 274 145 275 146 
<< m2 >>
rect 275 145 276 146 
<< m1 >>
rect 276 145 277 146 
<< m2 >>
rect 276 145 277 146 
<< m2 >>
rect 277 145 278 146 
<< m1 >>
rect 280 145 281 146 
<< m1 >>
rect 289 145 290 146 
<< m1 >>
rect 296 145 297 146 
<< m1 >>
rect 298 145 299 146 
<< m1 >>
rect 307 145 308 146 
<< m2 >>
rect 308 145 309 146 
<< m1 >>
rect 325 145 326 146 
<< m1 >>
rect 327 145 328 146 
<< m1 >>
rect 329 145 330 146 
<< m1 >>
rect 343 145 344 146 
<< m2 >>
rect 343 145 344 146 
<< m1 >>
rect 345 145 346 146 
<< m1 >>
rect 10 146 11 147 
<< m1 >>
rect 21 146 22 147 
<< m1 >>
rect 23 146 24 147 
<< m2 >>
rect 27 146 28 147 
<< m1 >>
rect 28 146 29 147 
<< m1 >>
rect 35 146 36 147 
<< m1 >>
rect 37 146 38 147 
<< m1 >>
rect 42 146 43 147 
<< m1 >>
rect 46 146 47 147 
<< m1 >>
rect 58 146 59 147 
<< m2 >>
rect 59 146 60 147 
<< m2 >>
rect 61 146 62 147 
<< m1 >>
rect 62 146 63 147 
<< m1 >>
rect 64 146 65 147 
<< m1 >>
rect 78 146 79 147 
<< m1 >>
rect 82 146 83 147 
<< m1 >>
rect 91 146 92 147 
<< m2 >>
rect 92 146 93 147 
<< m1 >>
rect 109 146 110 147 
<< m1 >>
rect 130 146 131 147 
<< m1 >>
rect 132 146 133 147 
<< m1 >>
rect 136 146 137 147 
<< m2 >>
rect 136 146 137 147 
<< m1 >>
rect 145 146 146 147 
<< m2 >>
rect 145 146 146 147 
<< m2 >>
rect 146 146 147 147 
<< m1 >>
rect 147 146 148 147 
<< m2 >>
rect 147 146 148 147 
<< m2 >>
rect 148 146 149 147 
<< m1 >>
rect 149 146 150 147 
<< m2 >>
rect 149 146 150 147 
<< m2c >>
rect 149 146 150 147 
<< m1 >>
rect 149 146 150 147 
<< m2 >>
rect 149 146 150 147 
<< m1 >>
rect 154 146 155 147 
<< m2 >>
rect 154 146 155 147 
<< m2c >>
rect 154 146 155 147 
<< m1 >>
rect 154 146 155 147 
<< m2 >>
rect 154 146 155 147 
<< m1 >>
rect 163 146 164 147 
<< m2 >>
rect 164 146 165 147 
<< m1 >>
rect 170 146 171 147 
<< m1 >>
rect 172 146 173 147 
<< m1 >>
rect 181 146 182 147 
<< m1 >>
rect 183 146 184 147 
<< m1 >>
rect 188 146 189 147 
<< m1 >>
rect 192 146 193 147 
<< m1 >>
rect 196 146 197 147 
<< m1 >>
rect 199 146 200 147 
<< m1 >>
rect 201 146 202 147 
<< m1 >>
rect 226 146 227 147 
<< m2 >>
rect 226 146 227 147 
<< m1 >>
rect 232 146 233 147 
<< m1 >>
rect 235 146 236 147 
<< m1 >>
rect 237 146 238 147 
<< m2 >>
rect 238 146 239 147 
<< m1 >>
rect 240 146 241 147 
<< m1 >>
rect 253 146 254 147 
<< m1 >>
rect 255 146 256 147 
<< m1 >>
rect 260 146 261 147 
<< m1 >>
rect 262 146 263 147 
<< m1 >>
rect 265 146 266 147 
<< m2 >>
rect 266 146 267 147 
<< m1 >>
rect 267 146 268 147 
<< m2 >>
rect 267 146 268 147 
<< m2c >>
rect 267 146 268 147 
<< m1 >>
rect 267 146 268 147 
<< m2 >>
rect 267 146 268 147 
<< m1 >>
rect 268 146 269 147 
<< m1 >>
rect 269 146 270 147 
<< m1 >>
rect 270 146 271 147 
<< m1 >>
rect 272 146 273 147 
<< m1 >>
rect 274 146 275 147 
<< m1 >>
rect 276 146 277 147 
<< m1 >>
rect 280 146 281 147 
<< m1 >>
rect 289 146 290 147 
<< m1 >>
rect 296 146 297 147 
<< m1 >>
rect 298 146 299 147 
<< m1 >>
rect 307 146 308 147 
<< m2 >>
rect 308 146 309 147 
<< m1 >>
rect 325 146 326 147 
<< m1 >>
rect 327 146 328 147 
<< m2 >>
rect 327 146 328 147 
<< m2c >>
rect 327 146 328 147 
<< m1 >>
rect 327 146 328 147 
<< m2 >>
rect 327 146 328 147 
<< m1 >>
rect 329 146 330 147 
<< m2 >>
rect 329 146 330 147 
<< m2c >>
rect 329 146 330 147 
<< m1 >>
rect 329 146 330 147 
<< m2 >>
rect 329 146 330 147 
<< m1 >>
rect 343 146 344 147 
<< m2 >>
rect 343 146 344 147 
<< m1 >>
rect 345 146 346 147 
<< m1 >>
rect 10 147 11 148 
<< m1 >>
rect 21 147 22 148 
<< m1 >>
rect 23 147 24 148 
<< m1 >>
rect 25 147 26 148 
<< m1 >>
rect 26 147 27 148 
<< m2 >>
rect 26 147 27 148 
<< m2c >>
rect 26 147 27 148 
<< m1 >>
rect 26 147 27 148 
<< m2 >>
rect 26 147 27 148 
<< m2 >>
rect 27 147 28 148 
<< m1 >>
rect 28 147 29 148 
<< m1 >>
rect 35 147 36 148 
<< m1 >>
rect 37 147 38 148 
<< m1 >>
rect 42 147 43 148 
<< m1 >>
rect 44 147 45 148 
<< m2 >>
rect 44 147 45 148 
<< m2c >>
rect 44 147 45 148 
<< m1 >>
rect 44 147 45 148 
<< m2 >>
rect 44 147 45 148 
<< m2 >>
rect 45 147 46 148 
<< m1 >>
rect 46 147 47 148 
<< m2 >>
rect 46 147 47 148 
<< m2 >>
rect 47 147 48 148 
<< m1 >>
rect 48 147 49 148 
<< m2 >>
rect 48 147 49 148 
<< m2c >>
rect 48 147 49 148 
<< m1 >>
rect 48 147 49 148 
<< m2 >>
rect 48 147 49 148 
<< m1 >>
rect 56 147 57 148 
<< m2 >>
rect 56 147 57 148 
<< m2c >>
rect 56 147 57 148 
<< m1 >>
rect 56 147 57 148 
<< m2 >>
rect 56 147 57 148 
<< m2 >>
rect 57 147 58 148 
<< m1 >>
rect 58 147 59 148 
<< m2 >>
rect 58 147 59 148 
<< m2 >>
rect 59 147 60 148 
<< m2 >>
rect 61 147 62 148 
<< m1 >>
rect 62 147 63 148 
<< m1 >>
rect 64 147 65 148 
<< m1 >>
rect 78 147 79 148 
<< m1 >>
rect 82 147 83 148 
<< m1 >>
rect 91 147 92 148 
<< m2 >>
rect 92 147 93 148 
<< m1 >>
rect 109 147 110 148 
<< m1 >>
rect 130 147 131 148 
<< m1 >>
rect 132 147 133 148 
<< m1 >>
rect 136 147 137 148 
<< m2 >>
rect 136 147 137 148 
<< m1 >>
rect 145 147 146 148 
<< m2 >>
rect 145 147 146 148 
<< m1 >>
rect 147 147 148 148 
<< m2 >>
rect 154 147 155 148 
<< m1 >>
rect 163 147 164 148 
<< m2 >>
rect 164 147 165 148 
<< m1 >>
rect 165 147 166 148 
<< m2 >>
rect 165 147 166 148 
<< m2c >>
rect 165 147 166 148 
<< m1 >>
rect 165 147 166 148 
<< m2 >>
rect 165 147 166 148 
<< m1 >>
rect 166 147 167 148 
<< m1 >>
rect 167 147 168 148 
<< m1 >>
rect 168 147 169 148 
<< m2 >>
rect 168 147 169 148 
<< m2c >>
rect 168 147 169 148 
<< m1 >>
rect 168 147 169 148 
<< m2 >>
rect 168 147 169 148 
<< m2 >>
rect 169 147 170 148 
<< m1 >>
rect 170 147 171 148 
<< m2 >>
rect 170 147 171 148 
<< m2 >>
rect 171 147 172 148 
<< m1 >>
rect 172 147 173 148 
<< m2 >>
rect 172 147 173 148 
<< m2 >>
rect 173 147 174 148 
<< m1 >>
rect 174 147 175 148 
<< m2 >>
rect 174 147 175 148 
<< m2c >>
rect 174 147 175 148 
<< m1 >>
rect 174 147 175 148 
<< m2 >>
rect 174 147 175 148 
<< m1 >>
rect 181 147 182 148 
<< m2 >>
rect 181 147 182 148 
<< m2c >>
rect 181 147 182 148 
<< m1 >>
rect 181 147 182 148 
<< m2 >>
rect 181 147 182 148 
<< m1 >>
rect 183 147 184 148 
<< m2 >>
rect 183 147 184 148 
<< m2c >>
rect 183 147 184 148 
<< m1 >>
rect 183 147 184 148 
<< m2 >>
rect 183 147 184 148 
<< m1 >>
rect 188 147 189 148 
<< m2 >>
rect 188 147 189 148 
<< m2c >>
rect 188 147 189 148 
<< m1 >>
rect 188 147 189 148 
<< m2 >>
rect 188 147 189 148 
<< m1 >>
rect 192 147 193 148 
<< m1 >>
rect 196 147 197 148 
<< m1 >>
rect 199 147 200 148 
<< m1 >>
rect 201 147 202 148 
<< m1 >>
rect 226 147 227 148 
<< m2 >>
rect 226 147 227 148 
<< m2 >>
rect 227 147 228 148 
<< m1 >>
rect 228 147 229 148 
<< m2 >>
rect 228 147 229 148 
<< m2c >>
rect 228 147 229 148 
<< m1 >>
rect 228 147 229 148 
<< m2 >>
rect 228 147 229 148 
<< m1 >>
rect 232 147 233 148 
<< m1 >>
rect 235 147 236 148 
<< m1 >>
rect 237 147 238 148 
<< m2 >>
rect 238 147 239 148 
<< m1 >>
rect 240 147 241 148 
<< m1 >>
rect 253 147 254 148 
<< m1 >>
rect 255 147 256 148 
<< m1 >>
rect 260 147 261 148 
<< m1 >>
rect 262 147 263 148 
<< m1 >>
rect 265 147 266 148 
<< m2 >>
rect 266 147 267 148 
<< m1 >>
rect 272 147 273 148 
<< m1 >>
rect 274 147 275 148 
<< m1 >>
rect 276 147 277 148 
<< m1 >>
rect 280 147 281 148 
<< m1 >>
rect 289 147 290 148 
<< m1 >>
rect 296 147 297 148 
<< m1 >>
rect 298 147 299 148 
<< m1 >>
rect 307 147 308 148 
<< m2 >>
rect 308 147 309 148 
<< m1 >>
rect 325 147 326 148 
<< m2 >>
rect 327 147 328 148 
<< m2 >>
rect 329 147 330 148 
<< m1 >>
rect 343 147 344 148 
<< m2 >>
rect 343 147 344 148 
<< m1 >>
rect 345 147 346 148 
<< m1 >>
rect 10 148 11 149 
<< m1 >>
rect 21 148 22 149 
<< m1 >>
rect 23 148 24 149 
<< m1 >>
rect 25 148 26 149 
<< m1 >>
rect 28 148 29 149 
<< m1 >>
rect 35 148 36 149 
<< m1 >>
rect 37 148 38 149 
<< m1 >>
rect 42 148 43 149 
<< m1 >>
rect 44 148 45 149 
<< m1 >>
rect 46 148 47 149 
<< m1 >>
rect 48 148 49 149 
<< m1 >>
rect 56 148 57 149 
<< m1 >>
rect 58 148 59 149 
<< m2 >>
rect 61 148 62 149 
<< m1 >>
rect 62 148 63 149 
<< m1 >>
rect 64 148 65 149 
<< m2 >>
rect 65 148 66 149 
<< m1 >>
rect 66 148 67 149 
<< m2 >>
rect 66 148 67 149 
<< m2c >>
rect 66 148 67 149 
<< m1 >>
rect 66 148 67 149 
<< m2 >>
rect 66 148 67 149 
<< m1 >>
rect 67 148 68 149 
<< m1 >>
rect 68 148 69 149 
<< m1 >>
rect 69 148 70 149 
<< m1 >>
rect 70 148 71 149 
<< m1 >>
rect 71 148 72 149 
<< m1 >>
rect 72 148 73 149 
<< m1 >>
rect 73 148 74 149 
<< m1 >>
rect 74 148 75 149 
<< m1 >>
rect 75 148 76 149 
<< m1 >>
rect 76 148 77 149 
<< m1 >>
rect 77 148 78 149 
<< m1 >>
rect 78 148 79 149 
<< m1 >>
rect 82 148 83 149 
<< m1 >>
rect 91 148 92 149 
<< m2 >>
rect 92 148 93 149 
<< m1 >>
rect 109 148 110 149 
<< m1 >>
rect 130 148 131 149 
<< m1 >>
rect 132 148 133 149 
<< m1 >>
rect 136 148 137 149 
<< m2 >>
rect 136 148 137 149 
<< m1 >>
rect 145 148 146 149 
<< m2 >>
rect 145 148 146 149 
<< m1 >>
rect 147 148 148 149 
<< m1 >>
rect 148 148 149 149 
<< m1 >>
rect 149 148 150 149 
<< m1 >>
rect 150 148 151 149 
<< m1 >>
rect 151 148 152 149 
<< m1 >>
rect 152 148 153 149 
<< m1 >>
rect 153 148 154 149 
<< m1 >>
rect 154 148 155 149 
<< m2 >>
rect 154 148 155 149 
<< m1 >>
rect 155 148 156 149 
<< m1 >>
rect 156 148 157 149 
<< m1 >>
rect 157 148 158 149 
<< m1 >>
rect 158 148 159 149 
<< m1 >>
rect 159 148 160 149 
<< m1 >>
rect 160 148 161 149 
<< m1 >>
rect 161 148 162 149 
<< m2 >>
rect 161 148 162 149 
<< m2c >>
rect 161 148 162 149 
<< m1 >>
rect 161 148 162 149 
<< m2 >>
rect 161 148 162 149 
<< m2 >>
rect 162 148 163 149 
<< m1 >>
rect 163 148 164 149 
<< m1 >>
rect 170 148 171 149 
<< m1 >>
rect 172 148 173 149 
<< m1 >>
rect 174 148 175 149 
<< m2 >>
rect 181 148 182 149 
<< m2 >>
rect 183 148 184 149 
<< m2 >>
rect 188 148 189 149 
<< m1 >>
rect 192 148 193 149 
<< m1 >>
rect 193 148 194 149 
<< m1 >>
rect 194 148 195 149 
<< m1 >>
rect 195 148 196 149 
<< m1 >>
rect 196 148 197 149 
<< m1 >>
rect 199 148 200 149 
<< m1 >>
rect 201 148 202 149 
<< m1 >>
rect 226 148 227 149 
<< m1 >>
rect 228 148 229 149 
<< m1 >>
rect 232 148 233 149 
<< m1 >>
rect 235 148 236 149 
<< m1 >>
rect 237 148 238 149 
<< m2 >>
rect 238 148 239 149 
<< m1 >>
rect 240 148 241 149 
<< m1 >>
rect 250 148 251 149 
<< m1 >>
rect 251 148 252 149 
<< m2 >>
rect 251 148 252 149 
<< m2c >>
rect 251 148 252 149 
<< m1 >>
rect 251 148 252 149 
<< m2 >>
rect 251 148 252 149 
<< m2 >>
rect 252 148 253 149 
<< m1 >>
rect 253 148 254 149 
<< m2 >>
rect 253 148 254 149 
<< m2 >>
rect 254 148 255 149 
<< m1 >>
rect 255 148 256 149 
<< m2 >>
rect 255 148 256 149 
<< m2 >>
rect 256 148 257 149 
<< m1 >>
rect 257 148 258 149 
<< m2 >>
rect 257 148 258 149 
<< m1 >>
rect 258 148 259 149 
<< m2 >>
rect 258 148 259 149 
<< m2c >>
rect 258 148 259 149 
<< m1 >>
rect 258 148 259 149 
<< m2 >>
rect 258 148 259 149 
<< m2 >>
rect 259 148 260 149 
<< m1 >>
rect 260 148 261 149 
<< m2 >>
rect 260 148 261 149 
<< m2 >>
rect 261 148 262 149 
<< m1 >>
rect 262 148 263 149 
<< m2 >>
rect 262 148 263 149 
<< m2 >>
rect 263 148 264 149 
<< m2 >>
rect 264 148 265 149 
<< m1 >>
rect 265 148 266 149 
<< m2 >>
rect 265 148 266 149 
<< m2 >>
rect 266 148 267 149 
<< m1 >>
rect 272 148 273 149 
<< m1 >>
rect 274 148 275 149 
<< m1 >>
rect 276 148 277 149 
<< m1 >>
rect 280 148 281 149 
<< m1 >>
rect 289 148 290 149 
<< m1 >>
rect 296 148 297 149 
<< m1 >>
rect 298 148 299 149 
<< m1 >>
rect 307 148 308 149 
<< m2 >>
rect 308 148 309 149 
<< m1 >>
rect 325 148 326 149 
<< m1 >>
rect 326 148 327 149 
<< m1 >>
rect 327 148 328 149 
<< m2 >>
rect 327 148 328 149 
<< m1 >>
rect 328 148 329 149 
<< m1 >>
rect 329 148 330 149 
<< m2 >>
rect 329 148 330 149 
<< m1 >>
rect 330 148 331 149 
<< m1 >>
rect 331 148 332 149 
<< m1 >>
rect 332 148 333 149 
<< m1 >>
rect 333 148 334 149 
<< m1 >>
rect 334 148 335 149 
<< m1 >>
rect 335 148 336 149 
<< m1 >>
rect 336 148 337 149 
<< m1 >>
rect 337 148 338 149 
<< m1 >>
rect 338 148 339 149 
<< m1 >>
rect 339 148 340 149 
<< m1 >>
rect 340 148 341 149 
<< m1 >>
rect 343 148 344 149 
<< m2 >>
rect 343 148 344 149 
<< m1 >>
rect 345 148 346 149 
<< m1 >>
rect 10 149 11 150 
<< m1 >>
rect 19 149 20 150 
<< m2 >>
rect 19 149 20 150 
<< m2c >>
rect 19 149 20 150 
<< m1 >>
rect 19 149 20 150 
<< m2 >>
rect 19 149 20 150 
<< m1 >>
rect 20 149 21 150 
<< m1 >>
rect 21 149 22 150 
<< m2 >>
rect 21 149 22 150 
<< m2 >>
rect 22 149 23 150 
<< m1 >>
rect 23 149 24 150 
<< m2 >>
rect 23 149 24 150 
<< m2c >>
rect 23 149 24 150 
<< m1 >>
rect 23 149 24 150 
<< m2 >>
rect 23 149 24 150 
<< m1 >>
rect 25 149 26 150 
<< m2 >>
rect 25 149 26 150 
<< m2c >>
rect 25 149 26 150 
<< m1 >>
rect 25 149 26 150 
<< m2 >>
rect 25 149 26 150 
<< m1 >>
rect 28 149 29 150 
<< m2 >>
rect 28 149 29 150 
<< m2c >>
rect 28 149 29 150 
<< m1 >>
rect 28 149 29 150 
<< m2 >>
rect 28 149 29 150 
<< m1 >>
rect 35 149 36 150 
<< m2 >>
rect 35 149 36 150 
<< m2c >>
rect 35 149 36 150 
<< m1 >>
rect 35 149 36 150 
<< m2 >>
rect 35 149 36 150 
<< m1 >>
rect 37 149 38 150 
<< m2 >>
rect 37 149 38 150 
<< m2c >>
rect 37 149 38 150 
<< m1 >>
rect 37 149 38 150 
<< m2 >>
rect 37 149 38 150 
<< m1 >>
rect 42 149 43 150 
<< m2 >>
rect 42 149 43 150 
<< m2c >>
rect 42 149 43 150 
<< m1 >>
rect 42 149 43 150 
<< m2 >>
rect 42 149 43 150 
<< m1 >>
rect 44 149 45 150 
<< m2 >>
rect 44 149 45 150 
<< m2c >>
rect 44 149 45 150 
<< m1 >>
rect 44 149 45 150 
<< m2 >>
rect 44 149 45 150 
<< m1 >>
rect 46 149 47 150 
<< m2 >>
rect 46 149 47 150 
<< m2c >>
rect 46 149 47 150 
<< m1 >>
rect 46 149 47 150 
<< m2 >>
rect 46 149 47 150 
<< m1 >>
rect 48 149 49 150 
<< m2 >>
rect 48 149 49 150 
<< m2c >>
rect 48 149 49 150 
<< m1 >>
rect 48 149 49 150 
<< m2 >>
rect 48 149 49 150 
<< m1 >>
rect 56 149 57 150 
<< m2 >>
rect 56 149 57 150 
<< m2c >>
rect 56 149 57 150 
<< m1 >>
rect 56 149 57 150 
<< m2 >>
rect 56 149 57 150 
<< m1 >>
rect 58 149 59 150 
<< m2 >>
rect 58 149 59 150 
<< m2c >>
rect 58 149 59 150 
<< m1 >>
rect 58 149 59 150 
<< m2 >>
rect 58 149 59 150 
<< m2 >>
rect 61 149 62 150 
<< m1 >>
rect 62 149 63 150 
<< m1 >>
rect 64 149 65 150 
<< m2 >>
rect 65 149 66 150 
<< m1 >>
rect 82 149 83 150 
<< m1 >>
rect 91 149 92 150 
<< m2 >>
rect 92 149 93 150 
<< m1 >>
rect 109 149 110 150 
<< m1 >>
rect 130 149 131 150 
<< m1 >>
rect 132 149 133 150 
<< m1 >>
rect 136 149 137 150 
<< m2 >>
rect 136 149 137 150 
<< m1 >>
rect 145 149 146 150 
<< m2 >>
rect 145 149 146 150 
<< m2 >>
rect 154 149 155 150 
<< m2 >>
rect 162 149 163 150 
<< m1 >>
rect 163 149 164 150 
<< m1 >>
rect 170 149 171 150 
<< m2 >>
rect 170 149 171 150 
<< m2c >>
rect 170 149 171 150 
<< m1 >>
rect 170 149 171 150 
<< m2 >>
rect 170 149 171 150 
<< m1 >>
rect 172 149 173 150 
<< m2 >>
rect 172 149 173 150 
<< m2c >>
rect 172 149 173 150 
<< m1 >>
rect 172 149 173 150 
<< m2 >>
rect 172 149 173 150 
<< m1 >>
rect 174 149 175 150 
<< m1 >>
rect 175 149 176 150 
<< m1 >>
rect 176 149 177 150 
<< m1 >>
rect 177 149 178 150 
<< m1 >>
rect 178 149 179 150 
<< m1 >>
rect 179 149 180 150 
<< m1 >>
rect 180 149 181 150 
<< m1 >>
rect 181 149 182 150 
<< m2 >>
rect 181 149 182 150 
<< m1 >>
rect 182 149 183 150 
<< m1 >>
rect 183 149 184 150 
<< m2 >>
rect 183 149 184 150 
<< m1 >>
rect 184 149 185 150 
<< m1 >>
rect 185 149 186 150 
<< m1 >>
rect 186 149 187 150 
<< m1 >>
rect 187 149 188 150 
<< m1 >>
rect 188 149 189 150 
<< m2 >>
rect 188 149 189 150 
<< m1 >>
rect 189 149 190 150 
<< m1 >>
rect 190 149 191 150 
<< m2 >>
rect 190 149 191 150 
<< m2c >>
rect 190 149 191 150 
<< m1 >>
rect 190 149 191 150 
<< m2 >>
rect 190 149 191 150 
<< m1 >>
rect 199 149 200 150 
<< m2 >>
rect 199 149 200 150 
<< m2c >>
rect 199 149 200 150 
<< m1 >>
rect 199 149 200 150 
<< m2 >>
rect 199 149 200 150 
<< m1 >>
rect 201 149 202 150 
<< m2 >>
rect 201 149 202 150 
<< m2c >>
rect 201 149 202 150 
<< m1 >>
rect 201 149 202 150 
<< m2 >>
rect 201 149 202 150 
<< m1 >>
rect 226 149 227 150 
<< m2 >>
rect 226 149 227 150 
<< m2c >>
rect 226 149 227 150 
<< m1 >>
rect 226 149 227 150 
<< m2 >>
rect 226 149 227 150 
<< m1 >>
rect 228 149 229 150 
<< m1 >>
rect 229 149 230 150 
<< m2 >>
rect 229 149 230 150 
<< m2c >>
rect 229 149 230 150 
<< m1 >>
rect 229 149 230 150 
<< m2 >>
rect 229 149 230 150 
<< m1 >>
rect 232 149 233 150 
<< m1 >>
rect 235 149 236 150 
<< m1 >>
rect 237 149 238 150 
<< m2 >>
rect 238 149 239 150 
<< m1 >>
rect 240 149 241 150 
<< m1 >>
rect 250 149 251 150 
<< m1 >>
rect 253 149 254 150 
<< m1 >>
rect 255 149 256 150 
<< m1 >>
rect 260 149 261 150 
<< m1 >>
rect 262 149 263 150 
<< m1 >>
rect 265 149 266 150 
<< m1 >>
rect 272 149 273 150 
<< m1 >>
rect 274 149 275 150 
<< m1 >>
rect 276 149 277 150 
<< m1 >>
rect 280 149 281 150 
<< m1 >>
rect 289 149 290 150 
<< m2 >>
rect 289 149 290 150 
<< m2c >>
rect 289 149 290 150 
<< m1 >>
rect 289 149 290 150 
<< m2 >>
rect 289 149 290 150 
<< m1 >>
rect 296 149 297 150 
<< m2 >>
rect 296 149 297 150 
<< m2c >>
rect 296 149 297 150 
<< m1 >>
rect 296 149 297 150 
<< m2 >>
rect 296 149 297 150 
<< m1 >>
rect 298 149 299 150 
<< m2 >>
rect 298 149 299 150 
<< m2c >>
rect 298 149 299 150 
<< m1 >>
rect 298 149 299 150 
<< m2 >>
rect 298 149 299 150 
<< m1 >>
rect 307 149 308 150 
<< m2 >>
rect 308 149 309 150 
<< m2 >>
rect 327 149 328 150 
<< m2 >>
rect 329 149 330 150 
<< m1 >>
rect 340 149 341 150 
<< m1 >>
rect 343 149 344 150 
<< m2 >>
rect 343 149 344 150 
<< m1 >>
rect 345 149 346 150 
<< m1 >>
rect 10 150 11 151 
<< m2 >>
rect 19 150 20 151 
<< m2 >>
rect 21 150 22 151 
<< m2 >>
rect 25 150 26 151 
<< m2 >>
rect 27 150 28 151 
<< m2 >>
rect 28 150 29 151 
<< m2 >>
rect 30 150 31 151 
<< m2 >>
rect 31 150 32 151 
<< m2 >>
rect 32 150 33 151 
<< m2 >>
rect 33 150 34 151 
<< m2 >>
rect 34 150 35 151 
<< m2 >>
rect 35 150 36 151 
<< m2 >>
rect 37 150 38 151 
<< m2 >>
rect 42 150 43 151 
<< m2 >>
rect 44 150 45 151 
<< m2 >>
rect 46 150 47 151 
<< m2 >>
rect 48 150 49 151 
<< m2 >>
rect 49 150 50 151 
<< m2 >>
rect 50 150 51 151 
<< m2 >>
rect 56 150 57 151 
<< m2 >>
rect 58 150 59 151 
<< m2 >>
rect 61 150 62 151 
<< m1 >>
rect 62 150 63 151 
<< m1 >>
rect 64 150 65 151 
<< m2 >>
rect 65 150 66 151 
<< m1 >>
rect 82 150 83 151 
<< m1 >>
rect 91 150 92 151 
<< m2 >>
rect 92 150 93 151 
<< m1 >>
rect 109 150 110 151 
<< m1 >>
rect 130 150 131 151 
<< m1 >>
rect 132 150 133 151 
<< m1 >>
rect 136 150 137 151 
<< m2 >>
rect 136 150 137 151 
<< m1 >>
rect 145 150 146 151 
<< m2 >>
rect 145 150 146 151 
<< m1 >>
rect 154 150 155 151 
<< m2 >>
rect 154 150 155 151 
<< m2c >>
rect 154 150 155 151 
<< m1 >>
rect 154 150 155 151 
<< m2 >>
rect 154 150 155 151 
<< m2 >>
rect 162 150 163 151 
<< m1 >>
rect 163 150 164 151 
<< m2 >>
rect 170 150 171 151 
<< m2 >>
rect 172 150 173 151 
<< m2 >>
rect 181 150 182 151 
<< m2 >>
rect 183 150 184 151 
<< m2 >>
rect 188 150 189 151 
<< m2 >>
rect 190 150 191 151 
<< m2 >>
rect 199 150 200 151 
<< m2 >>
rect 201 150 202 151 
<< m2 >>
rect 202 150 203 151 
<< m2 >>
rect 203 150 204 151 
<< m2 >>
rect 204 150 205 151 
<< m2 >>
rect 205 150 206 151 
<< m2 >>
rect 206 150 207 151 
<< m2 >>
rect 207 150 208 151 
<< m2 >>
rect 208 150 209 151 
<< m2 >>
rect 209 150 210 151 
<< m2 >>
rect 210 150 211 151 
<< m2 >>
rect 211 150 212 151 
<< m2 >>
rect 212 150 213 151 
<< m2 >>
rect 226 150 227 151 
<< m2 >>
rect 229 150 230 151 
<< m1 >>
rect 232 150 233 151 
<< m1 >>
rect 235 150 236 151 
<< m1 >>
rect 237 150 238 151 
<< m2 >>
rect 238 150 239 151 
<< m1 >>
rect 240 150 241 151 
<< m1 >>
rect 250 150 251 151 
<< m1 >>
rect 253 150 254 151 
<< m1 >>
rect 255 150 256 151 
<< m1 >>
rect 260 150 261 151 
<< m1 >>
rect 262 150 263 151 
<< m1 >>
rect 265 150 266 151 
<< m1 >>
rect 272 150 273 151 
<< m1 >>
rect 274 150 275 151 
<< m1 >>
rect 276 150 277 151 
<< m1 >>
rect 280 150 281 151 
<< m2 >>
rect 289 150 290 151 
<< m2 >>
rect 296 150 297 151 
<< m2 >>
rect 298 150 299 151 
<< m1 >>
rect 307 150 308 151 
<< m2 >>
rect 308 150 309 151 
<< m1 >>
rect 327 150 328 151 
<< m2 >>
rect 327 150 328 151 
<< m2c >>
rect 327 150 328 151 
<< m1 >>
rect 327 150 328 151 
<< m2 >>
rect 327 150 328 151 
<< m1 >>
rect 329 150 330 151 
<< m2 >>
rect 329 150 330 151 
<< m2c >>
rect 329 150 330 151 
<< m1 >>
rect 329 150 330 151 
<< m2 >>
rect 329 150 330 151 
<< m1 >>
rect 340 150 341 151 
<< m1 >>
rect 343 150 344 151 
<< m2 >>
rect 343 150 344 151 
<< m1 >>
rect 345 150 346 151 
<< m1 >>
rect 10 151 11 152 
<< m1 >>
rect 19 151 20 152 
<< m2 >>
rect 19 151 20 152 
<< m1 >>
rect 20 151 21 152 
<< m1 >>
rect 21 151 22 152 
<< m2 >>
rect 21 151 22 152 
<< m1 >>
rect 22 151 23 152 
<< m1 >>
rect 23 151 24 152 
<< m1 >>
rect 24 151 25 152 
<< m1 >>
rect 25 151 26 152 
<< m2 >>
rect 25 151 26 152 
<< m1 >>
rect 26 151 27 152 
<< m1 >>
rect 27 151 28 152 
<< m2 >>
rect 27 151 28 152 
<< m1 >>
rect 28 151 29 152 
<< m1 >>
rect 29 151 30 152 
<< m1 >>
rect 30 151 31 152 
<< m2 >>
rect 30 151 31 152 
<< m1 >>
rect 31 151 32 152 
<< m1 >>
rect 32 151 33 152 
<< m1 >>
rect 33 151 34 152 
<< m1 >>
rect 34 151 35 152 
<< m1 >>
rect 35 151 36 152 
<< m1 >>
rect 36 151 37 152 
<< m1 >>
rect 37 151 38 152 
<< m2 >>
rect 37 151 38 152 
<< m1 >>
rect 38 151 39 152 
<< m1 >>
rect 39 151 40 152 
<< m1 >>
rect 40 151 41 152 
<< m1 >>
rect 41 151 42 152 
<< m1 >>
rect 42 151 43 152 
<< m2 >>
rect 42 151 43 152 
<< m1 >>
rect 43 151 44 152 
<< m1 >>
rect 44 151 45 152 
<< m2 >>
rect 44 151 45 152 
<< m1 >>
rect 45 151 46 152 
<< m1 >>
rect 46 151 47 152 
<< m2 >>
rect 46 151 47 152 
<< m1 >>
rect 47 151 48 152 
<< m1 >>
rect 48 151 49 152 
<< m1 >>
rect 49 151 50 152 
<< m1 >>
rect 50 151 51 152 
<< m2 >>
rect 50 151 51 152 
<< m1 >>
rect 51 151 52 152 
<< m1 >>
rect 52 151 53 152 
<< m1 >>
rect 53 151 54 152 
<< m1 >>
rect 54 151 55 152 
<< m1 >>
rect 55 151 56 152 
<< m1 >>
rect 56 151 57 152 
<< m2 >>
rect 56 151 57 152 
<< m1 >>
rect 57 151 58 152 
<< m1 >>
rect 58 151 59 152 
<< m2 >>
rect 58 151 59 152 
<< m1 >>
rect 59 151 60 152 
<< m1 >>
rect 60 151 61 152 
<< m2 >>
rect 60 151 61 152 
<< m2c >>
rect 60 151 61 152 
<< m1 >>
rect 60 151 61 152 
<< m2 >>
rect 60 151 61 152 
<< m2 >>
rect 61 151 62 152 
<< m1 >>
rect 62 151 63 152 
<< m1 >>
rect 64 151 65 152 
<< m2 >>
rect 65 151 66 152 
<< m1 >>
rect 82 151 83 152 
<< m1 >>
rect 91 151 92 152 
<< m2 >>
rect 92 151 93 152 
<< m1 >>
rect 109 151 110 152 
<< m1 >>
rect 130 151 131 152 
<< m1 >>
rect 132 151 133 152 
<< m1 >>
rect 136 151 137 152 
<< m2 >>
rect 136 151 137 152 
<< m1 >>
rect 145 151 146 152 
<< m2 >>
rect 145 151 146 152 
<< m1 >>
rect 154 151 155 152 
<< m2 >>
rect 162 151 163 152 
<< m1 >>
rect 163 151 164 152 
<< m1 >>
rect 165 151 166 152 
<< m1 >>
rect 166 151 167 152 
<< m1 >>
rect 167 151 168 152 
<< m1 >>
rect 168 151 169 152 
<< m1 >>
rect 169 151 170 152 
<< m1 >>
rect 170 151 171 152 
<< m2 >>
rect 170 151 171 152 
<< m1 >>
rect 171 151 172 152 
<< m1 >>
rect 172 151 173 152 
<< m2 >>
rect 172 151 173 152 
<< m1 >>
rect 173 151 174 152 
<< m1 >>
rect 174 151 175 152 
<< m1 >>
rect 175 151 176 152 
<< m1 >>
rect 176 151 177 152 
<< m1 >>
rect 177 151 178 152 
<< m1 >>
rect 178 151 179 152 
<< m1 >>
rect 179 151 180 152 
<< m1 >>
rect 180 151 181 152 
<< m1 >>
rect 181 151 182 152 
<< m2 >>
rect 181 151 182 152 
<< m1 >>
rect 182 151 183 152 
<< m1 >>
rect 183 151 184 152 
<< m2 >>
rect 183 151 184 152 
<< m1 >>
rect 184 151 185 152 
<< m1 >>
rect 185 151 186 152 
<< m1 >>
rect 186 151 187 152 
<< m1 >>
rect 187 151 188 152 
<< m1 >>
rect 188 151 189 152 
<< m2 >>
rect 188 151 189 152 
<< m1 >>
rect 189 151 190 152 
<< m1 >>
rect 190 151 191 152 
<< m2 >>
rect 190 151 191 152 
<< m1 >>
rect 191 151 192 152 
<< m1 >>
rect 192 151 193 152 
<< m1 >>
rect 193 151 194 152 
<< m1 >>
rect 194 151 195 152 
<< m1 >>
rect 195 151 196 152 
<< m1 >>
rect 196 151 197 152 
<< m1 >>
rect 197 151 198 152 
<< m1 >>
rect 198 151 199 152 
<< m1 >>
rect 199 151 200 152 
<< m2 >>
rect 199 151 200 152 
<< m1 >>
rect 200 151 201 152 
<< m1 >>
rect 201 151 202 152 
<< m1 >>
rect 202 151 203 152 
<< m1 >>
rect 203 151 204 152 
<< m1 >>
rect 204 151 205 152 
<< m1 >>
rect 205 151 206 152 
<< m1 >>
rect 206 151 207 152 
<< m1 >>
rect 207 151 208 152 
<< m1 >>
rect 208 151 209 152 
<< m1 >>
rect 209 151 210 152 
<< m1 >>
rect 210 151 211 152 
<< m1 >>
rect 211 151 212 152 
<< m1 >>
rect 212 151 213 152 
<< m2 >>
rect 212 151 213 152 
<< m1 >>
rect 213 151 214 152 
<< m1 >>
rect 214 151 215 152 
<< m1 >>
rect 215 151 216 152 
<< m1 >>
rect 216 151 217 152 
<< m1 >>
rect 217 151 218 152 
<< m1 >>
rect 218 151 219 152 
<< m1 >>
rect 219 151 220 152 
<< m1 >>
rect 220 151 221 152 
<< m1 >>
rect 221 151 222 152 
<< m1 >>
rect 222 151 223 152 
<< m1 >>
rect 223 151 224 152 
<< m1 >>
rect 224 151 225 152 
<< m1 >>
rect 225 151 226 152 
<< m1 >>
rect 226 151 227 152 
<< m2 >>
rect 226 151 227 152 
<< m1 >>
rect 227 151 228 152 
<< m1 >>
rect 228 151 229 152 
<< m1 >>
rect 229 151 230 152 
<< m2 >>
rect 229 151 230 152 
<< m1 >>
rect 230 151 231 152 
<< m1 >>
rect 231 151 232 152 
<< m1 >>
rect 232 151 233 152 
<< m1 >>
rect 235 151 236 152 
<< m1 >>
rect 237 151 238 152 
<< m2 >>
rect 238 151 239 152 
<< m1 >>
rect 240 151 241 152 
<< m1 >>
rect 250 151 251 152 
<< m1 >>
rect 253 151 254 152 
<< m1 >>
rect 255 151 256 152 
<< m1 >>
rect 260 151 261 152 
<< m1 >>
rect 262 151 263 152 
<< m2 >>
rect 262 151 263 152 
<< m2 >>
rect 263 151 264 152 
<< m2 >>
rect 264 151 265 152 
<< m1 >>
rect 265 151 266 152 
<< m2 >>
rect 265 151 266 152 
<< m1 >>
rect 266 151 267 152 
<< m2 >>
rect 266 151 267 152 
<< m1 >>
rect 267 151 268 152 
<< m2 >>
rect 267 151 268 152 
<< m1 >>
rect 268 151 269 152 
<< m2 >>
rect 268 151 269 152 
<< m1 >>
rect 269 151 270 152 
<< m2 >>
rect 269 151 270 152 
<< m1 >>
rect 270 151 271 152 
<< m2 >>
rect 270 151 271 152 
<< m2 >>
rect 271 151 272 152 
<< m1 >>
rect 272 151 273 152 
<< m2 >>
rect 272 151 273 152 
<< m2 >>
rect 273 151 274 152 
<< m1 >>
rect 274 151 275 152 
<< m2 >>
rect 274 151 275 152 
<< m2 >>
rect 275 151 276 152 
<< m1 >>
rect 276 151 277 152 
<< m2 >>
rect 276 151 277 152 
<< m2 >>
rect 277 151 278 152 
<< m1 >>
rect 278 151 279 152 
<< m2 >>
rect 278 151 279 152 
<< m2c >>
rect 278 151 279 152 
<< m1 >>
rect 278 151 279 152 
<< m2 >>
rect 278 151 279 152 
<< m2 >>
rect 279 151 280 152 
<< m1 >>
rect 280 151 281 152 
<< m2 >>
rect 280 151 281 152 
<< m2 >>
rect 281 151 282 152 
<< m1 >>
rect 282 151 283 152 
<< m2 >>
rect 282 151 283 152 
<< m2c >>
rect 282 151 283 152 
<< m1 >>
rect 282 151 283 152 
<< m2 >>
rect 282 151 283 152 
<< m1 >>
rect 283 151 284 152 
<< m1 >>
rect 284 151 285 152 
<< m1 >>
rect 285 151 286 152 
<< m1 >>
rect 286 151 287 152 
<< m1 >>
rect 287 151 288 152 
<< m1 >>
rect 288 151 289 152 
<< m1 >>
rect 289 151 290 152 
<< m2 >>
rect 289 151 290 152 
<< m1 >>
rect 290 151 291 152 
<< m1 >>
rect 291 151 292 152 
<< m1 >>
rect 292 151 293 152 
<< m1 >>
rect 293 151 294 152 
<< m1 >>
rect 294 151 295 152 
<< m1 >>
rect 295 151 296 152 
<< m1 >>
rect 296 151 297 152 
<< m2 >>
rect 296 151 297 152 
<< m1 >>
rect 297 151 298 152 
<< m1 >>
rect 298 151 299 152 
<< m2 >>
rect 298 151 299 152 
<< m1 >>
rect 299 151 300 152 
<< m1 >>
rect 300 151 301 152 
<< m1 >>
rect 301 151 302 152 
<< m1 >>
rect 302 151 303 152 
<< m1 >>
rect 303 151 304 152 
<< m1 >>
rect 304 151 305 152 
<< m1 >>
rect 307 151 308 152 
<< m2 >>
rect 308 151 309 152 
<< m1 >>
rect 327 151 328 152 
<< m1 >>
rect 329 151 330 152 
<< m1 >>
rect 340 151 341 152 
<< m1 >>
rect 343 151 344 152 
<< m2 >>
rect 343 151 344 152 
<< m1 >>
rect 345 151 346 152 
<< m1 >>
rect 10 152 11 153 
<< m1 >>
rect 19 152 20 153 
<< m2 >>
rect 19 152 20 153 
<< m2 >>
rect 21 152 22 153 
<< m2 >>
rect 23 152 24 153 
<< m2 >>
rect 24 152 25 153 
<< m2 >>
rect 25 152 26 153 
<< m2 >>
rect 27 152 28 153 
<< m2 >>
rect 30 152 31 153 
<< m2 >>
rect 37 152 38 153 
<< m2 >>
rect 42 152 43 153 
<< m2 >>
rect 44 152 45 153 
<< m2 >>
rect 46 152 47 153 
<< m2 >>
rect 50 152 51 153 
<< m2 >>
rect 56 152 57 153 
<< m2 >>
rect 58 152 59 153 
<< m1 >>
rect 62 152 63 153 
<< m1 >>
rect 64 152 65 153 
<< m2 >>
rect 65 152 66 153 
<< m1 >>
rect 82 152 83 153 
<< m1 >>
rect 91 152 92 153 
<< m2 >>
rect 92 152 93 153 
<< m1 >>
rect 109 152 110 153 
<< m1 >>
rect 130 152 131 153 
<< m1 >>
rect 132 152 133 153 
<< m1 >>
rect 136 152 137 153 
<< m2 >>
rect 136 152 137 153 
<< m1 >>
rect 145 152 146 153 
<< m2 >>
rect 145 152 146 153 
<< m1 >>
rect 154 152 155 153 
<< m2 >>
rect 162 152 163 153 
<< m1 >>
rect 163 152 164 153 
<< m1 >>
rect 165 152 166 153 
<< m2 >>
rect 170 152 171 153 
<< m2 >>
rect 172 152 173 153 
<< m2 >>
rect 181 152 182 153 
<< m2 >>
rect 183 152 184 153 
<< m2 >>
rect 188 152 189 153 
<< m2 >>
rect 190 152 191 153 
<< m2 >>
rect 199 152 200 153 
<< m2 >>
rect 212 152 213 153 
<< m2 >>
rect 226 152 227 153 
<< m2 >>
rect 229 152 230 153 
<< m1 >>
rect 235 152 236 153 
<< m1 >>
rect 237 152 238 153 
<< m2 >>
rect 238 152 239 153 
<< m1 >>
rect 240 152 241 153 
<< m1 >>
rect 250 152 251 153 
<< m1 >>
rect 253 152 254 153 
<< m1 >>
rect 255 152 256 153 
<< m1 >>
rect 260 152 261 153 
<< m1 >>
rect 262 152 263 153 
<< m2 >>
rect 262 152 263 153 
<< m1 >>
rect 270 152 271 153 
<< m1 >>
rect 272 152 273 153 
<< m1 >>
rect 274 152 275 153 
<< m1 >>
rect 276 152 277 153 
<< m1 >>
rect 280 152 281 153 
<< m2 >>
rect 289 152 290 153 
<< m2 >>
rect 296 152 297 153 
<< m2 >>
rect 298 152 299 153 
<< m1 >>
rect 304 152 305 153 
<< m1 >>
rect 307 152 308 153 
<< m2 >>
rect 308 152 309 153 
<< m1 >>
rect 327 152 328 153 
<< m1 >>
rect 329 152 330 153 
<< m1 >>
rect 340 152 341 153 
<< m1 >>
rect 343 152 344 153 
<< m2 >>
rect 343 152 344 153 
<< m1 >>
rect 345 152 346 153 
<< m1 >>
rect 10 153 11 154 
<< m1 >>
rect 19 153 20 154 
<< m2 >>
rect 19 153 20 154 
<< m1 >>
rect 21 153 22 154 
<< m2 >>
rect 21 153 22 154 
<< m2c >>
rect 21 153 22 154 
<< m1 >>
rect 21 153 22 154 
<< m2 >>
rect 21 153 22 154 
<< m1 >>
rect 23 153 24 154 
<< m2 >>
rect 23 153 24 154 
<< m2c >>
rect 23 153 24 154 
<< m1 >>
rect 23 153 24 154 
<< m2 >>
rect 23 153 24 154 
<< m2 >>
rect 27 153 28 154 
<< m1 >>
rect 28 153 29 154 
<< m1 >>
rect 29 153 30 154 
<< m1 >>
rect 30 153 31 154 
<< m2 >>
rect 30 153 31 154 
<< m2c >>
rect 30 153 31 154 
<< m1 >>
rect 30 153 31 154 
<< m2 >>
rect 30 153 31 154 
<< m1 >>
rect 37 153 38 154 
<< m2 >>
rect 37 153 38 154 
<< m2c >>
rect 37 153 38 154 
<< m1 >>
rect 37 153 38 154 
<< m2 >>
rect 37 153 38 154 
<< m1 >>
rect 42 153 43 154 
<< m2 >>
rect 42 153 43 154 
<< m2c >>
rect 42 153 43 154 
<< m1 >>
rect 42 153 43 154 
<< m2 >>
rect 42 153 43 154 
<< m1 >>
rect 44 153 45 154 
<< m2 >>
rect 44 153 45 154 
<< m2c >>
rect 44 153 45 154 
<< m1 >>
rect 44 153 45 154 
<< m2 >>
rect 44 153 45 154 
<< m1 >>
rect 46 153 47 154 
<< m2 >>
rect 46 153 47 154 
<< m2c >>
rect 46 153 47 154 
<< m1 >>
rect 46 153 47 154 
<< m2 >>
rect 46 153 47 154 
<< m1 >>
rect 50 153 51 154 
<< m2 >>
rect 50 153 51 154 
<< m2c >>
rect 50 153 51 154 
<< m1 >>
rect 50 153 51 154 
<< m2 >>
rect 50 153 51 154 
<< m1 >>
rect 51 153 52 154 
<< m1 >>
rect 52 153 53 154 
<< m1 >>
rect 56 153 57 154 
<< m2 >>
rect 56 153 57 154 
<< m2c >>
rect 56 153 57 154 
<< m1 >>
rect 56 153 57 154 
<< m2 >>
rect 56 153 57 154 
<< m1 >>
rect 58 153 59 154 
<< m2 >>
rect 58 153 59 154 
<< m2c >>
rect 58 153 59 154 
<< m1 >>
rect 58 153 59 154 
<< m2 >>
rect 58 153 59 154 
<< m1 >>
rect 60 153 61 154 
<< m2 >>
rect 60 153 61 154 
<< m2c >>
rect 60 153 61 154 
<< m1 >>
rect 60 153 61 154 
<< m2 >>
rect 60 153 61 154 
<< m2 >>
rect 61 153 62 154 
<< m1 >>
rect 62 153 63 154 
<< m2 >>
rect 62 153 63 154 
<< m2 >>
rect 63 153 64 154 
<< m1 >>
rect 64 153 65 154 
<< m2 >>
rect 64 153 65 154 
<< m2 >>
rect 65 153 66 154 
<< m1 >>
rect 82 153 83 154 
<< m1 >>
rect 91 153 92 154 
<< m2 >>
rect 92 153 93 154 
<< m1 >>
rect 103 153 104 154 
<< m1 >>
rect 104 153 105 154 
<< m1 >>
rect 105 153 106 154 
<< m1 >>
rect 106 153 107 154 
<< m1 >>
rect 107 153 108 154 
<< m1 >>
rect 108 153 109 154 
<< m1 >>
rect 109 153 110 154 
<< m1 >>
rect 130 153 131 154 
<< m1 >>
rect 132 153 133 154 
<< m1 >>
rect 136 153 137 154 
<< m2 >>
rect 136 153 137 154 
<< m1 >>
rect 145 153 146 154 
<< m2 >>
rect 145 153 146 154 
<< m1 >>
rect 154 153 155 154 
<< m2 >>
rect 162 153 163 154 
<< m1 >>
rect 163 153 164 154 
<< m2 >>
rect 163 153 164 154 
<< m2 >>
rect 164 153 165 154 
<< m1 >>
rect 165 153 166 154 
<< m2 >>
rect 165 153 166 154 
<< m2 >>
rect 166 153 167 154 
<< m1 >>
rect 167 153 168 154 
<< m2 >>
rect 167 153 168 154 
<< m2c >>
rect 167 153 168 154 
<< m1 >>
rect 167 153 168 154 
<< m2 >>
rect 167 153 168 154 
<< m1 >>
rect 170 153 171 154 
<< m2 >>
rect 170 153 171 154 
<< m2c >>
rect 170 153 171 154 
<< m1 >>
rect 170 153 171 154 
<< m2 >>
rect 170 153 171 154 
<< m1 >>
rect 172 153 173 154 
<< m2 >>
rect 172 153 173 154 
<< m2c >>
rect 172 153 173 154 
<< m1 >>
rect 172 153 173 154 
<< m2 >>
rect 172 153 173 154 
<< m1 >>
rect 181 153 182 154 
<< m2 >>
rect 181 153 182 154 
<< m2c >>
rect 181 153 182 154 
<< m1 >>
rect 181 153 182 154 
<< m2 >>
rect 181 153 182 154 
<< m1 >>
rect 183 153 184 154 
<< m2 >>
rect 183 153 184 154 
<< m2c >>
rect 183 153 184 154 
<< m1 >>
rect 183 153 184 154 
<< m2 >>
rect 183 153 184 154 
<< m1 >>
rect 188 153 189 154 
<< m2 >>
rect 188 153 189 154 
<< m2c >>
rect 188 153 189 154 
<< m1 >>
rect 188 153 189 154 
<< m2 >>
rect 188 153 189 154 
<< m1 >>
rect 190 153 191 154 
<< m2 >>
rect 190 153 191 154 
<< m2c >>
rect 190 153 191 154 
<< m1 >>
rect 190 153 191 154 
<< m2 >>
rect 190 153 191 154 
<< m1 >>
rect 199 153 200 154 
<< m2 >>
rect 199 153 200 154 
<< m2c >>
rect 199 153 200 154 
<< m1 >>
rect 199 153 200 154 
<< m2 >>
rect 199 153 200 154 
<< m1 >>
rect 212 153 213 154 
<< m2 >>
rect 212 153 213 154 
<< m2c >>
rect 212 153 213 154 
<< m1 >>
rect 212 153 213 154 
<< m2 >>
rect 212 153 213 154 
<< m1 >>
rect 213 153 214 154 
<< m1 >>
rect 214 153 215 154 
<< m1 >>
rect 215 153 216 154 
<< m1 >>
rect 216 153 217 154 
<< m1 >>
rect 217 153 218 154 
<< m1 >>
rect 226 153 227 154 
<< m2 >>
rect 226 153 227 154 
<< m2c >>
rect 226 153 227 154 
<< m1 >>
rect 226 153 227 154 
<< m2 >>
rect 226 153 227 154 
<< m1 >>
rect 229 153 230 154 
<< m2 >>
rect 229 153 230 154 
<< m2c >>
rect 229 153 230 154 
<< m1 >>
rect 229 153 230 154 
<< m2 >>
rect 229 153 230 154 
<< m1 >>
rect 235 153 236 154 
<< m1 >>
rect 237 153 238 154 
<< m2 >>
rect 238 153 239 154 
<< m1 >>
rect 240 153 241 154 
<< m1 >>
rect 250 153 251 154 
<< m1 >>
rect 253 153 254 154 
<< m1 >>
rect 255 153 256 154 
<< m1 >>
rect 260 153 261 154 
<< m1 >>
rect 262 153 263 154 
<< m2 >>
rect 262 153 263 154 
<< m1 >>
rect 270 153 271 154 
<< m1 >>
rect 272 153 273 154 
<< m1 >>
rect 274 153 275 154 
<< m1 >>
rect 276 153 277 154 
<< m1 >>
rect 280 153 281 154 
<< m1 >>
rect 286 153 287 154 
<< m1 >>
rect 287 153 288 154 
<< m1 >>
rect 288 153 289 154 
<< m1 >>
rect 289 153 290 154 
<< m2 >>
rect 289 153 290 154 
<< m2c >>
rect 289 153 290 154 
<< m1 >>
rect 289 153 290 154 
<< m2 >>
rect 289 153 290 154 
<< m1 >>
rect 296 153 297 154 
<< m2 >>
rect 296 153 297 154 
<< m2c >>
rect 296 153 297 154 
<< m1 >>
rect 296 153 297 154 
<< m2 >>
rect 296 153 297 154 
<< m1 >>
rect 298 153 299 154 
<< m2 >>
rect 298 153 299 154 
<< m2c >>
rect 298 153 299 154 
<< m1 >>
rect 298 153 299 154 
<< m2 >>
rect 298 153 299 154 
<< m1 >>
rect 304 153 305 154 
<< m1 >>
rect 307 153 308 154 
<< m2 >>
rect 308 153 309 154 
<< m1 >>
rect 327 153 328 154 
<< m1 >>
rect 329 153 330 154 
<< m1 >>
rect 340 153 341 154 
<< m1 >>
rect 343 153 344 154 
<< m2 >>
rect 343 153 344 154 
<< m1 >>
rect 345 153 346 154 
<< m1 >>
rect 10 154 11 155 
<< m1 >>
rect 19 154 20 155 
<< m2 >>
rect 19 154 20 155 
<< m1 >>
rect 21 154 22 155 
<< m1 >>
rect 23 154 24 155 
<< m2 >>
rect 27 154 28 155 
<< m1 >>
rect 28 154 29 155 
<< m1 >>
rect 37 154 38 155 
<< m1 >>
rect 42 154 43 155 
<< m1 >>
rect 44 154 45 155 
<< m1 >>
rect 46 154 47 155 
<< m1 >>
rect 52 154 53 155 
<< m1 >>
rect 56 154 57 155 
<< m1 >>
rect 58 154 59 155 
<< m1 >>
rect 60 154 61 155 
<< m1 >>
rect 62 154 63 155 
<< m1 >>
rect 64 154 65 155 
<< m1 >>
rect 82 154 83 155 
<< m1 >>
rect 91 154 92 155 
<< m2 >>
rect 92 154 93 155 
<< m1 >>
rect 103 154 104 155 
<< m1 >>
rect 130 154 131 155 
<< m1 >>
rect 132 154 133 155 
<< m1 >>
rect 136 154 137 155 
<< m2 >>
rect 136 154 137 155 
<< m1 >>
rect 145 154 146 155 
<< m2 >>
rect 145 154 146 155 
<< m1 >>
rect 154 154 155 155 
<< m1 >>
rect 163 154 164 155 
<< m1 >>
rect 165 154 166 155 
<< m1 >>
rect 167 154 168 155 
<< m1 >>
rect 170 154 171 155 
<< m1 >>
rect 172 154 173 155 
<< m1 >>
rect 181 154 182 155 
<< m1 >>
rect 183 154 184 155 
<< m1 >>
rect 188 154 189 155 
<< m1 >>
rect 190 154 191 155 
<< m1 >>
rect 199 154 200 155 
<< m1 >>
rect 217 154 218 155 
<< m1 >>
rect 226 154 227 155 
<< m1 >>
rect 229 154 230 155 
<< m1 >>
rect 235 154 236 155 
<< m1 >>
rect 237 154 238 155 
<< m2 >>
rect 238 154 239 155 
<< m1 >>
rect 240 154 241 155 
<< m1 >>
rect 250 154 251 155 
<< m1 >>
rect 253 154 254 155 
<< m1 >>
rect 255 154 256 155 
<< m1 >>
rect 260 154 261 155 
<< m1 >>
rect 262 154 263 155 
<< m2 >>
rect 262 154 263 155 
<< m1 >>
rect 270 154 271 155 
<< m2 >>
rect 270 154 271 155 
<< m2c >>
rect 270 154 271 155 
<< m1 >>
rect 270 154 271 155 
<< m2 >>
rect 270 154 271 155 
<< m2 >>
rect 271 154 272 155 
<< m1 >>
rect 272 154 273 155 
<< m2 >>
rect 272 154 273 155 
<< m2 >>
rect 273 154 274 155 
<< m1 >>
rect 274 154 275 155 
<< m2 >>
rect 274 154 275 155 
<< m2 >>
rect 275 154 276 155 
<< m1 >>
rect 276 154 277 155 
<< m1 >>
rect 280 154 281 155 
<< m1 >>
rect 286 154 287 155 
<< m1 >>
rect 296 154 297 155 
<< m1 >>
rect 298 154 299 155 
<< m1 >>
rect 304 154 305 155 
<< m1 >>
rect 307 154 308 155 
<< m2 >>
rect 308 154 309 155 
<< m1 >>
rect 327 154 328 155 
<< m1 >>
rect 329 154 330 155 
<< m1 >>
rect 340 154 341 155 
<< m1 >>
rect 343 154 344 155 
<< m2 >>
rect 343 154 344 155 
<< m1 >>
rect 345 154 346 155 
<< m1 >>
rect 10 155 11 156 
<< m1 >>
rect 19 155 20 156 
<< m2 >>
rect 19 155 20 156 
<< m1 >>
rect 21 155 22 156 
<< m1 >>
rect 23 155 24 156 
<< m2 >>
rect 27 155 28 156 
<< m1 >>
rect 28 155 29 156 
<< m1 >>
rect 37 155 38 156 
<< m2 >>
rect 38 155 39 156 
<< m1 >>
rect 39 155 40 156 
<< m2 >>
rect 39 155 40 156 
<< m2c >>
rect 39 155 40 156 
<< m1 >>
rect 39 155 40 156 
<< m2 >>
rect 39 155 40 156 
<< m1 >>
rect 40 155 41 156 
<< m1 >>
rect 41 155 42 156 
<< m1 >>
rect 42 155 43 156 
<< m1 >>
rect 44 155 45 156 
<< m1 >>
rect 46 155 47 156 
<< m1 >>
rect 52 155 53 156 
<< m1 >>
rect 56 155 57 156 
<< m1 >>
rect 58 155 59 156 
<< m1 >>
rect 60 155 61 156 
<< m1 >>
rect 62 155 63 156 
<< m1 >>
rect 64 155 65 156 
<< m1 >>
rect 82 155 83 156 
<< m1 >>
rect 91 155 92 156 
<< m2 >>
rect 92 155 93 156 
<< m1 >>
rect 103 155 104 156 
<< m1 >>
rect 130 155 131 156 
<< m1 >>
rect 132 155 133 156 
<< m1 >>
rect 136 155 137 156 
<< m2 >>
rect 136 155 137 156 
<< m1 >>
rect 145 155 146 156 
<< m2 >>
rect 145 155 146 156 
<< m1 >>
rect 154 155 155 156 
<< m1 >>
rect 163 155 164 156 
<< m1 >>
rect 165 155 166 156 
<< m1 >>
rect 167 155 168 156 
<< m1 >>
rect 168 155 169 156 
<< m2 >>
rect 168 155 169 156 
<< m2c >>
rect 168 155 169 156 
<< m1 >>
rect 168 155 169 156 
<< m2 >>
rect 168 155 169 156 
<< m2 >>
rect 169 155 170 156 
<< m1 >>
rect 170 155 171 156 
<< m1 >>
rect 172 155 173 156 
<< m1 >>
rect 181 155 182 156 
<< m2 >>
rect 181 155 182 156 
<< m2c >>
rect 181 155 182 156 
<< m1 >>
rect 181 155 182 156 
<< m2 >>
rect 181 155 182 156 
<< m2 >>
rect 182 155 183 156 
<< m1 >>
rect 183 155 184 156 
<< m2 >>
rect 183 155 184 156 
<< m2 >>
rect 184 155 185 156 
<< m1 >>
rect 185 155 186 156 
<< m2 >>
rect 185 155 186 156 
<< m2c >>
rect 185 155 186 156 
<< m1 >>
rect 185 155 186 156 
<< m2 >>
rect 185 155 186 156 
<< m1 >>
rect 186 155 187 156 
<< m2 >>
rect 186 155 187 156 
<< m2 >>
rect 187 155 188 156 
<< m1 >>
rect 188 155 189 156 
<< m1 >>
rect 190 155 191 156 
<< m1 >>
rect 199 155 200 156 
<< m1 >>
rect 217 155 218 156 
<< m1 >>
rect 218 155 219 156 
<< m1 >>
rect 219 155 220 156 
<< m1 >>
rect 220 155 221 156 
<< m1 >>
rect 221 155 222 156 
<< m1 >>
rect 222 155 223 156 
<< m1 >>
rect 223 155 224 156 
<< m1 >>
rect 224 155 225 156 
<< m2 >>
rect 224 155 225 156 
<< m2c >>
rect 224 155 225 156 
<< m1 >>
rect 224 155 225 156 
<< m2 >>
rect 224 155 225 156 
<< m2 >>
rect 225 155 226 156 
<< m1 >>
rect 226 155 227 156 
<< m1 >>
rect 229 155 230 156 
<< m1 >>
rect 235 155 236 156 
<< m1 >>
rect 237 155 238 156 
<< m2 >>
rect 238 155 239 156 
<< m1 >>
rect 240 155 241 156 
<< m1 >>
rect 250 155 251 156 
<< m1 >>
rect 253 155 254 156 
<< m1 >>
rect 255 155 256 156 
<< m1 >>
rect 260 155 261 156 
<< m1 >>
rect 262 155 263 156 
<< m2 >>
rect 262 155 263 156 
<< m1 >>
rect 272 155 273 156 
<< m1 >>
rect 274 155 275 156 
<< m2 >>
rect 275 155 276 156 
<< m1 >>
rect 276 155 277 156 
<< m1 >>
rect 280 155 281 156 
<< m1 >>
rect 286 155 287 156 
<< m1 >>
rect 296 155 297 156 
<< m1 >>
rect 298 155 299 156 
<< m1 >>
rect 304 155 305 156 
<< m1 >>
rect 307 155 308 156 
<< m2 >>
rect 308 155 309 156 
<< m1 >>
rect 327 155 328 156 
<< m1 >>
rect 329 155 330 156 
<< m1 >>
rect 340 155 341 156 
<< m1 >>
rect 343 155 344 156 
<< m2 >>
rect 343 155 344 156 
<< m1 >>
rect 345 155 346 156 
<< m1 >>
rect 10 156 11 157 
<< pdiffusion >>
rect 12 156 13 157 
<< pdiffusion >>
rect 13 156 14 157 
<< pdiffusion >>
rect 14 156 15 157 
<< pdiffusion >>
rect 15 156 16 157 
<< pdiffusion >>
rect 16 156 17 157 
<< pdiffusion >>
rect 17 156 18 157 
<< m1 >>
rect 19 156 20 157 
<< m2 >>
rect 19 156 20 157 
<< m1 >>
rect 21 156 22 157 
<< m1 >>
rect 23 156 24 157 
<< m2 >>
rect 27 156 28 157 
<< m1 >>
rect 28 156 29 157 
<< pdiffusion >>
rect 30 156 31 157 
<< pdiffusion >>
rect 31 156 32 157 
<< pdiffusion >>
rect 32 156 33 157 
<< pdiffusion >>
rect 33 156 34 157 
<< pdiffusion >>
rect 34 156 35 157 
<< pdiffusion >>
rect 35 156 36 157 
<< m1 >>
rect 37 156 38 157 
<< m2 >>
rect 38 156 39 157 
<< m1 >>
rect 44 156 45 157 
<< m1 >>
rect 46 156 47 157 
<< pdiffusion >>
rect 48 156 49 157 
<< pdiffusion >>
rect 49 156 50 157 
<< pdiffusion >>
rect 50 156 51 157 
<< pdiffusion >>
rect 51 156 52 157 
<< m1 >>
rect 52 156 53 157 
<< pdiffusion >>
rect 52 156 53 157 
<< pdiffusion >>
rect 53 156 54 157 
<< m1 >>
rect 56 156 57 157 
<< m1 >>
rect 58 156 59 157 
<< m1 >>
rect 60 156 61 157 
<< m1 >>
rect 62 156 63 157 
<< m1 >>
rect 64 156 65 157 
<< pdiffusion >>
rect 66 156 67 157 
<< pdiffusion >>
rect 67 156 68 157 
<< pdiffusion >>
rect 68 156 69 157 
<< pdiffusion >>
rect 69 156 70 157 
<< pdiffusion >>
rect 70 156 71 157 
<< pdiffusion >>
rect 71 156 72 157 
<< m1 >>
rect 82 156 83 157 
<< pdiffusion >>
rect 84 156 85 157 
<< pdiffusion >>
rect 85 156 86 157 
<< pdiffusion >>
rect 86 156 87 157 
<< pdiffusion >>
rect 87 156 88 157 
<< pdiffusion >>
rect 88 156 89 157 
<< pdiffusion >>
rect 89 156 90 157 
<< m1 >>
rect 91 156 92 157 
<< m2 >>
rect 92 156 93 157 
<< pdiffusion >>
rect 102 156 103 157 
<< m1 >>
rect 103 156 104 157 
<< pdiffusion >>
rect 103 156 104 157 
<< pdiffusion >>
rect 104 156 105 157 
<< pdiffusion >>
rect 105 156 106 157 
<< pdiffusion >>
rect 106 156 107 157 
<< pdiffusion >>
rect 107 156 108 157 
<< pdiffusion >>
rect 120 156 121 157 
<< pdiffusion >>
rect 121 156 122 157 
<< pdiffusion >>
rect 122 156 123 157 
<< pdiffusion >>
rect 123 156 124 157 
<< pdiffusion >>
rect 124 156 125 157 
<< pdiffusion >>
rect 125 156 126 157 
<< m1 >>
rect 130 156 131 157 
<< m1 >>
rect 132 156 133 157 
<< m1 >>
rect 136 156 137 157 
<< m2 >>
rect 136 156 137 157 
<< pdiffusion >>
rect 138 156 139 157 
<< pdiffusion >>
rect 139 156 140 157 
<< pdiffusion >>
rect 140 156 141 157 
<< pdiffusion >>
rect 141 156 142 157 
<< pdiffusion >>
rect 142 156 143 157 
<< pdiffusion >>
rect 143 156 144 157 
<< m1 >>
rect 145 156 146 157 
<< m2 >>
rect 145 156 146 157 
<< m1 >>
rect 154 156 155 157 
<< pdiffusion >>
rect 156 156 157 157 
<< pdiffusion >>
rect 157 156 158 157 
<< pdiffusion >>
rect 158 156 159 157 
<< pdiffusion >>
rect 159 156 160 157 
<< pdiffusion >>
rect 160 156 161 157 
<< pdiffusion >>
rect 161 156 162 157 
<< m1 >>
rect 163 156 164 157 
<< m1 >>
rect 165 156 166 157 
<< m2 >>
rect 169 156 170 157 
<< m1 >>
rect 170 156 171 157 
<< m1 >>
rect 172 156 173 157 
<< pdiffusion >>
rect 174 156 175 157 
<< pdiffusion >>
rect 175 156 176 157 
<< pdiffusion >>
rect 176 156 177 157 
<< pdiffusion >>
rect 177 156 178 157 
<< pdiffusion >>
rect 178 156 179 157 
<< pdiffusion >>
rect 179 156 180 157 
<< m1 >>
rect 183 156 184 157 
<< m2 >>
rect 187 156 188 157 
<< m1 >>
rect 188 156 189 157 
<< m1 >>
rect 190 156 191 157 
<< pdiffusion >>
rect 192 156 193 157 
<< pdiffusion >>
rect 193 156 194 157 
<< pdiffusion >>
rect 194 156 195 157 
<< pdiffusion >>
rect 195 156 196 157 
<< pdiffusion >>
rect 196 156 197 157 
<< pdiffusion >>
rect 197 156 198 157 
<< m1 >>
rect 199 156 200 157 
<< pdiffusion >>
rect 210 156 211 157 
<< pdiffusion >>
rect 211 156 212 157 
<< pdiffusion >>
rect 212 156 213 157 
<< pdiffusion >>
rect 213 156 214 157 
<< pdiffusion >>
rect 214 156 215 157 
<< pdiffusion >>
rect 215 156 216 157 
<< m2 >>
rect 225 156 226 157 
<< m1 >>
rect 226 156 227 157 
<< pdiffusion >>
rect 228 156 229 157 
<< m1 >>
rect 229 156 230 157 
<< pdiffusion >>
rect 229 156 230 157 
<< pdiffusion >>
rect 230 156 231 157 
<< pdiffusion >>
rect 231 156 232 157 
<< pdiffusion >>
rect 232 156 233 157 
<< pdiffusion >>
rect 233 156 234 157 
<< m1 >>
rect 235 156 236 157 
<< m1 >>
rect 237 156 238 157 
<< m2 >>
rect 238 156 239 157 
<< m1 >>
rect 240 156 241 157 
<< pdiffusion >>
rect 246 156 247 157 
<< pdiffusion >>
rect 247 156 248 157 
<< pdiffusion >>
rect 248 156 249 157 
<< pdiffusion >>
rect 249 156 250 157 
<< m1 >>
rect 250 156 251 157 
<< pdiffusion >>
rect 250 156 251 157 
<< pdiffusion >>
rect 251 156 252 157 
<< m1 >>
rect 253 156 254 157 
<< m1 >>
rect 255 156 256 157 
<< m1 >>
rect 260 156 261 157 
<< m1 >>
rect 262 156 263 157 
<< m2 >>
rect 262 156 263 157 
<< pdiffusion >>
rect 264 156 265 157 
<< pdiffusion >>
rect 265 156 266 157 
<< pdiffusion >>
rect 266 156 267 157 
<< pdiffusion >>
rect 267 156 268 157 
<< pdiffusion >>
rect 268 156 269 157 
<< pdiffusion >>
rect 269 156 270 157 
<< m1 >>
rect 272 156 273 157 
<< m1 >>
rect 274 156 275 157 
<< m2 >>
rect 275 156 276 157 
<< m1 >>
rect 276 156 277 157 
<< m1 >>
rect 280 156 281 157 
<< pdiffusion >>
rect 282 156 283 157 
<< pdiffusion >>
rect 283 156 284 157 
<< pdiffusion >>
rect 284 156 285 157 
<< pdiffusion >>
rect 285 156 286 157 
<< m1 >>
rect 286 156 287 157 
<< pdiffusion >>
rect 286 156 287 157 
<< pdiffusion >>
rect 287 156 288 157 
<< m1 >>
rect 296 156 297 157 
<< m1 >>
rect 298 156 299 157 
<< pdiffusion >>
rect 300 156 301 157 
<< pdiffusion >>
rect 301 156 302 157 
<< pdiffusion >>
rect 302 156 303 157 
<< pdiffusion >>
rect 303 156 304 157 
<< m1 >>
rect 304 156 305 157 
<< pdiffusion >>
rect 304 156 305 157 
<< pdiffusion >>
rect 305 156 306 157 
<< m1 >>
rect 307 156 308 157 
<< m2 >>
rect 308 156 309 157 
<< pdiffusion >>
rect 318 156 319 157 
<< pdiffusion >>
rect 319 156 320 157 
<< pdiffusion >>
rect 320 156 321 157 
<< pdiffusion >>
rect 321 156 322 157 
<< pdiffusion >>
rect 322 156 323 157 
<< pdiffusion >>
rect 323 156 324 157 
<< m1 >>
rect 327 156 328 157 
<< m1 >>
rect 329 156 330 157 
<< pdiffusion >>
rect 336 156 337 157 
<< pdiffusion >>
rect 337 156 338 157 
<< pdiffusion >>
rect 338 156 339 157 
<< pdiffusion >>
rect 339 156 340 157 
<< m1 >>
rect 340 156 341 157 
<< pdiffusion >>
rect 340 156 341 157 
<< pdiffusion >>
rect 341 156 342 157 
<< m1 >>
rect 343 156 344 157 
<< m2 >>
rect 343 156 344 157 
<< m1 >>
rect 345 156 346 157 
<< m1 >>
rect 10 157 11 158 
<< pdiffusion >>
rect 12 157 13 158 
<< pdiffusion >>
rect 13 157 14 158 
<< pdiffusion >>
rect 14 157 15 158 
<< pdiffusion >>
rect 15 157 16 158 
<< pdiffusion >>
rect 16 157 17 158 
<< pdiffusion >>
rect 17 157 18 158 
<< m1 >>
rect 19 157 20 158 
<< m2 >>
rect 19 157 20 158 
<< m1 >>
rect 21 157 22 158 
<< m1 >>
rect 23 157 24 158 
<< m2 >>
rect 27 157 28 158 
<< m1 >>
rect 28 157 29 158 
<< pdiffusion >>
rect 30 157 31 158 
<< pdiffusion >>
rect 31 157 32 158 
<< pdiffusion >>
rect 32 157 33 158 
<< pdiffusion >>
rect 33 157 34 158 
<< pdiffusion >>
rect 34 157 35 158 
<< pdiffusion >>
rect 35 157 36 158 
<< m1 >>
rect 37 157 38 158 
<< m2 >>
rect 38 157 39 158 
<< m1 >>
rect 44 157 45 158 
<< m1 >>
rect 46 157 47 158 
<< pdiffusion >>
rect 48 157 49 158 
<< pdiffusion >>
rect 49 157 50 158 
<< pdiffusion >>
rect 50 157 51 158 
<< pdiffusion >>
rect 51 157 52 158 
<< pdiffusion >>
rect 52 157 53 158 
<< pdiffusion >>
rect 53 157 54 158 
<< m1 >>
rect 56 157 57 158 
<< m1 >>
rect 58 157 59 158 
<< m1 >>
rect 60 157 61 158 
<< m1 >>
rect 62 157 63 158 
<< m1 >>
rect 64 157 65 158 
<< pdiffusion >>
rect 66 157 67 158 
<< pdiffusion >>
rect 67 157 68 158 
<< pdiffusion >>
rect 68 157 69 158 
<< pdiffusion >>
rect 69 157 70 158 
<< pdiffusion >>
rect 70 157 71 158 
<< pdiffusion >>
rect 71 157 72 158 
<< m1 >>
rect 82 157 83 158 
<< pdiffusion >>
rect 84 157 85 158 
<< pdiffusion >>
rect 85 157 86 158 
<< pdiffusion >>
rect 86 157 87 158 
<< pdiffusion >>
rect 87 157 88 158 
<< pdiffusion >>
rect 88 157 89 158 
<< pdiffusion >>
rect 89 157 90 158 
<< m1 >>
rect 91 157 92 158 
<< m2 >>
rect 92 157 93 158 
<< pdiffusion >>
rect 102 157 103 158 
<< pdiffusion >>
rect 103 157 104 158 
<< pdiffusion >>
rect 104 157 105 158 
<< pdiffusion >>
rect 105 157 106 158 
<< pdiffusion >>
rect 106 157 107 158 
<< pdiffusion >>
rect 107 157 108 158 
<< pdiffusion >>
rect 120 157 121 158 
<< pdiffusion >>
rect 121 157 122 158 
<< pdiffusion >>
rect 122 157 123 158 
<< pdiffusion >>
rect 123 157 124 158 
<< pdiffusion >>
rect 124 157 125 158 
<< pdiffusion >>
rect 125 157 126 158 
<< m1 >>
rect 130 157 131 158 
<< m1 >>
rect 132 157 133 158 
<< m1 >>
rect 136 157 137 158 
<< m2 >>
rect 136 157 137 158 
<< pdiffusion >>
rect 138 157 139 158 
<< pdiffusion >>
rect 139 157 140 158 
<< pdiffusion >>
rect 140 157 141 158 
<< pdiffusion >>
rect 141 157 142 158 
<< pdiffusion >>
rect 142 157 143 158 
<< pdiffusion >>
rect 143 157 144 158 
<< m1 >>
rect 145 157 146 158 
<< m2 >>
rect 145 157 146 158 
<< m1 >>
rect 154 157 155 158 
<< pdiffusion >>
rect 156 157 157 158 
<< pdiffusion >>
rect 157 157 158 158 
<< pdiffusion >>
rect 158 157 159 158 
<< pdiffusion >>
rect 159 157 160 158 
<< pdiffusion >>
rect 160 157 161 158 
<< pdiffusion >>
rect 161 157 162 158 
<< m1 >>
rect 163 157 164 158 
<< m1 >>
rect 165 157 166 158 
<< m2 >>
rect 169 157 170 158 
<< m1 >>
rect 170 157 171 158 
<< m1 >>
rect 172 157 173 158 
<< pdiffusion >>
rect 174 157 175 158 
<< pdiffusion >>
rect 175 157 176 158 
<< pdiffusion >>
rect 176 157 177 158 
<< pdiffusion >>
rect 177 157 178 158 
<< pdiffusion >>
rect 178 157 179 158 
<< pdiffusion >>
rect 179 157 180 158 
<< m1 >>
rect 183 157 184 158 
<< m2 >>
rect 187 157 188 158 
<< m1 >>
rect 188 157 189 158 
<< m1 >>
rect 190 157 191 158 
<< pdiffusion >>
rect 192 157 193 158 
<< pdiffusion >>
rect 193 157 194 158 
<< pdiffusion >>
rect 194 157 195 158 
<< pdiffusion >>
rect 195 157 196 158 
<< pdiffusion >>
rect 196 157 197 158 
<< pdiffusion >>
rect 197 157 198 158 
<< m1 >>
rect 199 157 200 158 
<< pdiffusion >>
rect 210 157 211 158 
<< pdiffusion >>
rect 211 157 212 158 
<< pdiffusion >>
rect 212 157 213 158 
<< pdiffusion >>
rect 213 157 214 158 
<< pdiffusion >>
rect 214 157 215 158 
<< pdiffusion >>
rect 215 157 216 158 
<< m2 >>
rect 225 157 226 158 
<< m1 >>
rect 226 157 227 158 
<< pdiffusion >>
rect 228 157 229 158 
<< pdiffusion >>
rect 229 157 230 158 
<< pdiffusion >>
rect 230 157 231 158 
<< pdiffusion >>
rect 231 157 232 158 
<< pdiffusion >>
rect 232 157 233 158 
<< pdiffusion >>
rect 233 157 234 158 
<< m1 >>
rect 235 157 236 158 
<< m1 >>
rect 237 157 238 158 
<< m2 >>
rect 238 157 239 158 
<< m1 >>
rect 240 157 241 158 
<< pdiffusion >>
rect 246 157 247 158 
<< pdiffusion >>
rect 247 157 248 158 
<< pdiffusion >>
rect 248 157 249 158 
<< pdiffusion >>
rect 249 157 250 158 
<< pdiffusion >>
rect 250 157 251 158 
<< pdiffusion >>
rect 251 157 252 158 
<< m1 >>
rect 253 157 254 158 
<< m1 >>
rect 255 157 256 158 
<< m1 >>
rect 260 157 261 158 
<< m1 >>
rect 262 157 263 158 
<< m2 >>
rect 262 157 263 158 
<< pdiffusion >>
rect 264 157 265 158 
<< pdiffusion >>
rect 265 157 266 158 
<< pdiffusion >>
rect 266 157 267 158 
<< pdiffusion >>
rect 267 157 268 158 
<< pdiffusion >>
rect 268 157 269 158 
<< pdiffusion >>
rect 269 157 270 158 
<< m1 >>
rect 272 157 273 158 
<< m1 >>
rect 274 157 275 158 
<< m2 >>
rect 275 157 276 158 
<< m1 >>
rect 276 157 277 158 
<< m1 >>
rect 280 157 281 158 
<< pdiffusion >>
rect 282 157 283 158 
<< pdiffusion >>
rect 283 157 284 158 
<< pdiffusion >>
rect 284 157 285 158 
<< pdiffusion >>
rect 285 157 286 158 
<< pdiffusion >>
rect 286 157 287 158 
<< pdiffusion >>
rect 287 157 288 158 
<< m1 >>
rect 296 157 297 158 
<< m1 >>
rect 298 157 299 158 
<< pdiffusion >>
rect 300 157 301 158 
<< pdiffusion >>
rect 301 157 302 158 
<< pdiffusion >>
rect 302 157 303 158 
<< pdiffusion >>
rect 303 157 304 158 
<< pdiffusion >>
rect 304 157 305 158 
<< pdiffusion >>
rect 305 157 306 158 
<< m1 >>
rect 307 157 308 158 
<< m2 >>
rect 308 157 309 158 
<< pdiffusion >>
rect 318 157 319 158 
<< pdiffusion >>
rect 319 157 320 158 
<< pdiffusion >>
rect 320 157 321 158 
<< pdiffusion >>
rect 321 157 322 158 
<< pdiffusion >>
rect 322 157 323 158 
<< pdiffusion >>
rect 323 157 324 158 
<< m1 >>
rect 327 157 328 158 
<< m1 >>
rect 329 157 330 158 
<< pdiffusion >>
rect 336 157 337 158 
<< pdiffusion >>
rect 337 157 338 158 
<< pdiffusion >>
rect 338 157 339 158 
<< pdiffusion >>
rect 339 157 340 158 
<< pdiffusion >>
rect 340 157 341 158 
<< pdiffusion >>
rect 341 157 342 158 
<< m1 >>
rect 343 157 344 158 
<< m2 >>
rect 343 157 344 158 
<< m1 >>
rect 345 157 346 158 
<< m1 >>
rect 10 158 11 159 
<< pdiffusion >>
rect 12 158 13 159 
<< pdiffusion >>
rect 13 158 14 159 
<< pdiffusion >>
rect 14 158 15 159 
<< pdiffusion >>
rect 15 158 16 159 
<< pdiffusion >>
rect 16 158 17 159 
<< pdiffusion >>
rect 17 158 18 159 
<< m1 >>
rect 19 158 20 159 
<< m2 >>
rect 19 158 20 159 
<< m1 >>
rect 21 158 22 159 
<< m1 >>
rect 23 158 24 159 
<< m2 >>
rect 27 158 28 159 
<< m1 >>
rect 28 158 29 159 
<< pdiffusion >>
rect 30 158 31 159 
<< pdiffusion >>
rect 31 158 32 159 
<< pdiffusion >>
rect 32 158 33 159 
<< pdiffusion >>
rect 33 158 34 159 
<< pdiffusion >>
rect 34 158 35 159 
<< pdiffusion >>
rect 35 158 36 159 
<< m1 >>
rect 37 158 38 159 
<< m2 >>
rect 38 158 39 159 
<< m1 >>
rect 44 158 45 159 
<< m1 >>
rect 46 158 47 159 
<< pdiffusion >>
rect 48 158 49 159 
<< pdiffusion >>
rect 49 158 50 159 
<< pdiffusion >>
rect 50 158 51 159 
<< pdiffusion >>
rect 51 158 52 159 
<< pdiffusion >>
rect 52 158 53 159 
<< pdiffusion >>
rect 53 158 54 159 
<< m1 >>
rect 56 158 57 159 
<< m1 >>
rect 58 158 59 159 
<< m1 >>
rect 60 158 61 159 
<< m1 >>
rect 62 158 63 159 
<< m1 >>
rect 64 158 65 159 
<< pdiffusion >>
rect 66 158 67 159 
<< pdiffusion >>
rect 67 158 68 159 
<< pdiffusion >>
rect 68 158 69 159 
<< pdiffusion >>
rect 69 158 70 159 
<< pdiffusion >>
rect 70 158 71 159 
<< pdiffusion >>
rect 71 158 72 159 
<< m1 >>
rect 82 158 83 159 
<< pdiffusion >>
rect 84 158 85 159 
<< pdiffusion >>
rect 85 158 86 159 
<< pdiffusion >>
rect 86 158 87 159 
<< pdiffusion >>
rect 87 158 88 159 
<< pdiffusion >>
rect 88 158 89 159 
<< pdiffusion >>
rect 89 158 90 159 
<< m1 >>
rect 91 158 92 159 
<< m2 >>
rect 92 158 93 159 
<< pdiffusion >>
rect 102 158 103 159 
<< pdiffusion >>
rect 103 158 104 159 
<< pdiffusion >>
rect 104 158 105 159 
<< pdiffusion >>
rect 105 158 106 159 
<< pdiffusion >>
rect 106 158 107 159 
<< pdiffusion >>
rect 107 158 108 159 
<< pdiffusion >>
rect 120 158 121 159 
<< pdiffusion >>
rect 121 158 122 159 
<< pdiffusion >>
rect 122 158 123 159 
<< pdiffusion >>
rect 123 158 124 159 
<< pdiffusion >>
rect 124 158 125 159 
<< pdiffusion >>
rect 125 158 126 159 
<< m1 >>
rect 130 158 131 159 
<< m1 >>
rect 132 158 133 159 
<< m1 >>
rect 136 158 137 159 
<< m2 >>
rect 136 158 137 159 
<< pdiffusion >>
rect 138 158 139 159 
<< pdiffusion >>
rect 139 158 140 159 
<< pdiffusion >>
rect 140 158 141 159 
<< pdiffusion >>
rect 141 158 142 159 
<< pdiffusion >>
rect 142 158 143 159 
<< pdiffusion >>
rect 143 158 144 159 
<< m1 >>
rect 145 158 146 159 
<< m2 >>
rect 145 158 146 159 
<< m1 >>
rect 154 158 155 159 
<< pdiffusion >>
rect 156 158 157 159 
<< pdiffusion >>
rect 157 158 158 159 
<< pdiffusion >>
rect 158 158 159 159 
<< pdiffusion >>
rect 159 158 160 159 
<< pdiffusion >>
rect 160 158 161 159 
<< pdiffusion >>
rect 161 158 162 159 
<< m1 >>
rect 163 158 164 159 
<< m1 >>
rect 165 158 166 159 
<< m2 >>
rect 169 158 170 159 
<< m1 >>
rect 170 158 171 159 
<< m1 >>
rect 172 158 173 159 
<< pdiffusion >>
rect 174 158 175 159 
<< pdiffusion >>
rect 175 158 176 159 
<< pdiffusion >>
rect 176 158 177 159 
<< pdiffusion >>
rect 177 158 178 159 
<< pdiffusion >>
rect 178 158 179 159 
<< pdiffusion >>
rect 179 158 180 159 
<< m1 >>
rect 183 158 184 159 
<< m2 >>
rect 187 158 188 159 
<< m1 >>
rect 188 158 189 159 
<< m1 >>
rect 190 158 191 159 
<< pdiffusion >>
rect 192 158 193 159 
<< pdiffusion >>
rect 193 158 194 159 
<< pdiffusion >>
rect 194 158 195 159 
<< pdiffusion >>
rect 195 158 196 159 
<< pdiffusion >>
rect 196 158 197 159 
<< pdiffusion >>
rect 197 158 198 159 
<< m1 >>
rect 199 158 200 159 
<< pdiffusion >>
rect 210 158 211 159 
<< pdiffusion >>
rect 211 158 212 159 
<< pdiffusion >>
rect 212 158 213 159 
<< pdiffusion >>
rect 213 158 214 159 
<< pdiffusion >>
rect 214 158 215 159 
<< pdiffusion >>
rect 215 158 216 159 
<< m2 >>
rect 225 158 226 159 
<< m1 >>
rect 226 158 227 159 
<< pdiffusion >>
rect 228 158 229 159 
<< pdiffusion >>
rect 229 158 230 159 
<< pdiffusion >>
rect 230 158 231 159 
<< pdiffusion >>
rect 231 158 232 159 
<< pdiffusion >>
rect 232 158 233 159 
<< pdiffusion >>
rect 233 158 234 159 
<< m1 >>
rect 235 158 236 159 
<< m1 >>
rect 237 158 238 159 
<< m2 >>
rect 238 158 239 159 
<< m1 >>
rect 240 158 241 159 
<< pdiffusion >>
rect 246 158 247 159 
<< pdiffusion >>
rect 247 158 248 159 
<< pdiffusion >>
rect 248 158 249 159 
<< pdiffusion >>
rect 249 158 250 159 
<< pdiffusion >>
rect 250 158 251 159 
<< pdiffusion >>
rect 251 158 252 159 
<< m1 >>
rect 253 158 254 159 
<< m1 >>
rect 255 158 256 159 
<< m1 >>
rect 260 158 261 159 
<< m1 >>
rect 262 158 263 159 
<< m2 >>
rect 262 158 263 159 
<< pdiffusion >>
rect 264 158 265 159 
<< pdiffusion >>
rect 265 158 266 159 
<< pdiffusion >>
rect 266 158 267 159 
<< pdiffusion >>
rect 267 158 268 159 
<< pdiffusion >>
rect 268 158 269 159 
<< pdiffusion >>
rect 269 158 270 159 
<< m1 >>
rect 272 158 273 159 
<< m1 >>
rect 274 158 275 159 
<< m2 >>
rect 275 158 276 159 
<< m1 >>
rect 276 158 277 159 
<< m1 >>
rect 280 158 281 159 
<< pdiffusion >>
rect 282 158 283 159 
<< pdiffusion >>
rect 283 158 284 159 
<< pdiffusion >>
rect 284 158 285 159 
<< pdiffusion >>
rect 285 158 286 159 
<< pdiffusion >>
rect 286 158 287 159 
<< pdiffusion >>
rect 287 158 288 159 
<< m1 >>
rect 296 158 297 159 
<< m1 >>
rect 298 158 299 159 
<< pdiffusion >>
rect 300 158 301 159 
<< pdiffusion >>
rect 301 158 302 159 
<< pdiffusion >>
rect 302 158 303 159 
<< pdiffusion >>
rect 303 158 304 159 
<< pdiffusion >>
rect 304 158 305 159 
<< pdiffusion >>
rect 305 158 306 159 
<< m1 >>
rect 307 158 308 159 
<< m2 >>
rect 308 158 309 159 
<< pdiffusion >>
rect 318 158 319 159 
<< pdiffusion >>
rect 319 158 320 159 
<< pdiffusion >>
rect 320 158 321 159 
<< pdiffusion >>
rect 321 158 322 159 
<< pdiffusion >>
rect 322 158 323 159 
<< pdiffusion >>
rect 323 158 324 159 
<< m1 >>
rect 327 158 328 159 
<< m1 >>
rect 329 158 330 159 
<< pdiffusion >>
rect 336 158 337 159 
<< pdiffusion >>
rect 337 158 338 159 
<< pdiffusion >>
rect 338 158 339 159 
<< pdiffusion >>
rect 339 158 340 159 
<< pdiffusion >>
rect 340 158 341 159 
<< pdiffusion >>
rect 341 158 342 159 
<< m1 >>
rect 343 158 344 159 
<< m2 >>
rect 343 158 344 159 
<< m1 >>
rect 345 158 346 159 
<< m1 >>
rect 10 159 11 160 
<< pdiffusion >>
rect 12 159 13 160 
<< pdiffusion >>
rect 13 159 14 160 
<< pdiffusion >>
rect 14 159 15 160 
<< pdiffusion >>
rect 15 159 16 160 
<< pdiffusion >>
rect 16 159 17 160 
<< pdiffusion >>
rect 17 159 18 160 
<< m1 >>
rect 19 159 20 160 
<< m2 >>
rect 19 159 20 160 
<< m1 >>
rect 21 159 22 160 
<< m1 >>
rect 23 159 24 160 
<< m2 >>
rect 27 159 28 160 
<< m1 >>
rect 28 159 29 160 
<< pdiffusion >>
rect 30 159 31 160 
<< pdiffusion >>
rect 31 159 32 160 
<< pdiffusion >>
rect 32 159 33 160 
<< pdiffusion >>
rect 33 159 34 160 
<< pdiffusion >>
rect 34 159 35 160 
<< pdiffusion >>
rect 35 159 36 160 
<< m1 >>
rect 37 159 38 160 
<< m2 >>
rect 38 159 39 160 
<< m1 >>
rect 44 159 45 160 
<< m1 >>
rect 46 159 47 160 
<< pdiffusion >>
rect 48 159 49 160 
<< pdiffusion >>
rect 49 159 50 160 
<< pdiffusion >>
rect 50 159 51 160 
<< pdiffusion >>
rect 51 159 52 160 
<< pdiffusion >>
rect 52 159 53 160 
<< pdiffusion >>
rect 53 159 54 160 
<< m1 >>
rect 56 159 57 160 
<< m1 >>
rect 58 159 59 160 
<< m1 >>
rect 60 159 61 160 
<< m1 >>
rect 62 159 63 160 
<< m1 >>
rect 64 159 65 160 
<< pdiffusion >>
rect 66 159 67 160 
<< pdiffusion >>
rect 67 159 68 160 
<< pdiffusion >>
rect 68 159 69 160 
<< pdiffusion >>
rect 69 159 70 160 
<< pdiffusion >>
rect 70 159 71 160 
<< pdiffusion >>
rect 71 159 72 160 
<< m1 >>
rect 82 159 83 160 
<< pdiffusion >>
rect 84 159 85 160 
<< pdiffusion >>
rect 85 159 86 160 
<< pdiffusion >>
rect 86 159 87 160 
<< pdiffusion >>
rect 87 159 88 160 
<< pdiffusion >>
rect 88 159 89 160 
<< pdiffusion >>
rect 89 159 90 160 
<< m1 >>
rect 91 159 92 160 
<< m2 >>
rect 92 159 93 160 
<< pdiffusion >>
rect 102 159 103 160 
<< pdiffusion >>
rect 103 159 104 160 
<< pdiffusion >>
rect 104 159 105 160 
<< pdiffusion >>
rect 105 159 106 160 
<< pdiffusion >>
rect 106 159 107 160 
<< pdiffusion >>
rect 107 159 108 160 
<< pdiffusion >>
rect 120 159 121 160 
<< pdiffusion >>
rect 121 159 122 160 
<< pdiffusion >>
rect 122 159 123 160 
<< pdiffusion >>
rect 123 159 124 160 
<< pdiffusion >>
rect 124 159 125 160 
<< pdiffusion >>
rect 125 159 126 160 
<< m1 >>
rect 130 159 131 160 
<< m1 >>
rect 132 159 133 160 
<< m1 >>
rect 136 159 137 160 
<< m2 >>
rect 136 159 137 160 
<< pdiffusion >>
rect 138 159 139 160 
<< pdiffusion >>
rect 139 159 140 160 
<< pdiffusion >>
rect 140 159 141 160 
<< pdiffusion >>
rect 141 159 142 160 
<< pdiffusion >>
rect 142 159 143 160 
<< pdiffusion >>
rect 143 159 144 160 
<< m1 >>
rect 145 159 146 160 
<< m2 >>
rect 145 159 146 160 
<< m1 >>
rect 154 159 155 160 
<< pdiffusion >>
rect 156 159 157 160 
<< pdiffusion >>
rect 157 159 158 160 
<< pdiffusion >>
rect 158 159 159 160 
<< pdiffusion >>
rect 159 159 160 160 
<< pdiffusion >>
rect 160 159 161 160 
<< pdiffusion >>
rect 161 159 162 160 
<< m1 >>
rect 163 159 164 160 
<< m1 >>
rect 165 159 166 160 
<< m2 >>
rect 169 159 170 160 
<< m1 >>
rect 170 159 171 160 
<< m1 >>
rect 172 159 173 160 
<< pdiffusion >>
rect 174 159 175 160 
<< pdiffusion >>
rect 175 159 176 160 
<< pdiffusion >>
rect 176 159 177 160 
<< pdiffusion >>
rect 177 159 178 160 
<< pdiffusion >>
rect 178 159 179 160 
<< pdiffusion >>
rect 179 159 180 160 
<< m1 >>
rect 183 159 184 160 
<< m2 >>
rect 187 159 188 160 
<< m1 >>
rect 188 159 189 160 
<< m1 >>
rect 190 159 191 160 
<< pdiffusion >>
rect 192 159 193 160 
<< pdiffusion >>
rect 193 159 194 160 
<< pdiffusion >>
rect 194 159 195 160 
<< pdiffusion >>
rect 195 159 196 160 
<< pdiffusion >>
rect 196 159 197 160 
<< pdiffusion >>
rect 197 159 198 160 
<< m1 >>
rect 199 159 200 160 
<< pdiffusion >>
rect 210 159 211 160 
<< pdiffusion >>
rect 211 159 212 160 
<< pdiffusion >>
rect 212 159 213 160 
<< pdiffusion >>
rect 213 159 214 160 
<< pdiffusion >>
rect 214 159 215 160 
<< pdiffusion >>
rect 215 159 216 160 
<< m2 >>
rect 225 159 226 160 
<< m1 >>
rect 226 159 227 160 
<< pdiffusion >>
rect 228 159 229 160 
<< pdiffusion >>
rect 229 159 230 160 
<< pdiffusion >>
rect 230 159 231 160 
<< pdiffusion >>
rect 231 159 232 160 
<< pdiffusion >>
rect 232 159 233 160 
<< pdiffusion >>
rect 233 159 234 160 
<< m1 >>
rect 235 159 236 160 
<< m1 >>
rect 237 159 238 160 
<< m2 >>
rect 238 159 239 160 
<< m1 >>
rect 240 159 241 160 
<< pdiffusion >>
rect 246 159 247 160 
<< pdiffusion >>
rect 247 159 248 160 
<< pdiffusion >>
rect 248 159 249 160 
<< pdiffusion >>
rect 249 159 250 160 
<< pdiffusion >>
rect 250 159 251 160 
<< pdiffusion >>
rect 251 159 252 160 
<< m1 >>
rect 253 159 254 160 
<< m1 >>
rect 255 159 256 160 
<< m1 >>
rect 260 159 261 160 
<< m1 >>
rect 262 159 263 160 
<< m2 >>
rect 262 159 263 160 
<< pdiffusion >>
rect 264 159 265 160 
<< pdiffusion >>
rect 265 159 266 160 
<< pdiffusion >>
rect 266 159 267 160 
<< pdiffusion >>
rect 267 159 268 160 
<< pdiffusion >>
rect 268 159 269 160 
<< pdiffusion >>
rect 269 159 270 160 
<< m1 >>
rect 272 159 273 160 
<< m1 >>
rect 274 159 275 160 
<< m2 >>
rect 275 159 276 160 
<< m1 >>
rect 276 159 277 160 
<< m1 >>
rect 280 159 281 160 
<< pdiffusion >>
rect 282 159 283 160 
<< pdiffusion >>
rect 283 159 284 160 
<< pdiffusion >>
rect 284 159 285 160 
<< pdiffusion >>
rect 285 159 286 160 
<< pdiffusion >>
rect 286 159 287 160 
<< pdiffusion >>
rect 287 159 288 160 
<< m1 >>
rect 296 159 297 160 
<< m1 >>
rect 298 159 299 160 
<< pdiffusion >>
rect 300 159 301 160 
<< pdiffusion >>
rect 301 159 302 160 
<< pdiffusion >>
rect 302 159 303 160 
<< pdiffusion >>
rect 303 159 304 160 
<< pdiffusion >>
rect 304 159 305 160 
<< pdiffusion >>
rect 305 159 306 160 
<< m1 >>
rect 307 159 308 160 
<< m2 >>
rect 308 159 309 160 
<< pdiffusion >>
rect 318 159 319 160 
<< pdiffusion >>
rect 319 159 320 160 
<< pdiffusion >>
rect 320 159 321 160 
<< pdiffusion >>
rect 321 159 322 160 
<< pdiffusion >>
rect 322 159 323 160 
<< pdiffusion >>
rect 323 159 324 160 
<< m1 >>
rect 327 159 328 160 
<< m1 >>
rect 329 159 330 160 
<< pdiffusion >>
rect 336 159 337 160 
<< pdiffusion >>
rect 337 159 338 160 
<< pdiffusion >>
rect 338 159 339 160 
<< pdiffusion >>
rect 339 159 340 160 
<< pdiffusion >>
rect 340 159 341 160 
<< pdiffusion >>
rect 341 159 342 160 
<< m1 >>
rect 343 159 344 160 
<< m2 >>
rect 343 159 344 160 
<< m1 >>
rect 345 159 346 160 
<< m1 >>
rect 10 160 11 161 
<< pdiffusion >>
rect 12 160 13 161 
<< pdiffusion >>
rect 13 160 14 161 
<< pdiffusion >>
rect 14 160 15 161 
<< pdiffusion >>
rect 15 160 16 161 
<< pdiffusion >>
rect 16 160 17 161 
<< pdiffusion >>
rect 17 160 18 161 
<< m1 >>
rect 19 160 20 161 
<< m2 >>
rect 19 160 20 161 
<< m1 >>
rect 21 160 22 161 
<< m1 >>
rect 23 160 24 161 
<< m2 >>
rect 27 160 28 161 
<< m1 >>
rect 28 160 29 161 
<< pdiffusion >>
rect 30 160 31 161 
<< pdiffusion >>
rect 31 160 32 161 
<< pdiffusion >>
rect 32 160 33 161 
<< pdiffusion >>
rect 33 160 34 161 
<< pdiffusion >>
rect 34 160 35 161 
<< pdiffusion >>
rect 35 160 36 161 
<< m1 >>
rect 37 160 38 161 
<< m2 >>
rect 38 160 39 161 
<< m1 >>
rect 44 160 45 161 
<< m1 >>
rect 46 160 47 161 
<< pdiffusion >>
rect 48 160 49 161 
<< pdiffusion >>
rect 49 160 50 161 
<< pdiffusion >>
rect 50 160 51 161 
<< pdiffusion >>
rect 51 160 52 161 
<< pdiffusion >>
rect 52 160 53 161 
<< pdiffusion >>
rect 53 160 54 161 
<< m1 >>
rect 56 160 57 161 
<< m1 >>
rect 58 160 59 161 
<< m1 >>
rect 60 160 61 161 
<< m1 >>
rect 62 160 63 161 
<< m1 >>
rect 64 160 65 161 
<< pdiffusion >>
rect 66 160 67 161 
<< pdiffusion >>
rect 67 160 68 161 
<< pdiffusion >>
rect 68 160 69 161 
<< pdiffusion >>
rect 69 160 70 161 
<< pdiffusion >>
rect 70 160 71 161 
<< pdiffusion >>
rect 71 160 72 161 
<< m1 >>
rect 82 160 83 161 
<< pdiffusion >>
rect 84 160 85 161 
<< pdiffusion >>
rect 85 160 86 161 
<< pdiffusion >>
rect 86 160 87 161 
<< pdiffusion >>
rect 87 160 88 161 
<< pdiffusion >>
rect 88 160 89 161 
<< pdiffusion >>
rect 89 160 90 161 
<< m1 >>
rect 91 160 92 161 
<< m2 >>
rect 92 160 93 161 
<< pdiffusion >>
rect 102 160 103 161 
<< pdiffusion >>
rect 103 160 104 161 
<< pdiffusion >>
rect 104 160 105 161 
<< pdiffusion >>
rect 105 160 106 161 
<< pdiffusion >>
rect 106 160 107 161 
<< pdiffusion >>
rect 107 160 108 161 
<< pdiffusion >>
rect 120 160 121 161 
<< pdiffusion >>
rect 121 160 122 161 
<< pdiffusion >>
rect 122 160 123 161 
<< pdiffusion >>
rect 123 160 124 161 
<< pdiffusion >>
rect 124 160 125 161 
<< pdiffusion >>
rect 125 160 126 161 
<< m1 >>
rect 130 160 131 161 
<< m1 >>
rect 132 160 133 161 
<< m1 >>
rect 136 160 137 161 
<< m2 >>
rect 136 160 137 161 
<< pdiffusion >>
rect 138 160 139 161 
<< pdiffusion >>
rect 139 160 140 161 
<< pdiffusion >>
rect 140 160 141 161 
<< pdiffusion >>
rect 141 160 142 161 
<< pdiffusion >>
rect 142 160 143 161 
<< pdiffusion >>
rect 143 160 144 161 
<< m1 >>
rect 145 160 146 161 
<< m2 >>
rect 145 160 146 161 
<< m1 >>
rect 154 160 155 161 
<< pdiffusion >>
rect 156 160 157 161 
<< pdiffusion >>
rect 157 160 158 161 
<< pdiffusion >>
rect 158 160 159 161 
<< pdiffusion >>
rect 159 160 160 161 
<< pdiffusion >>
rect 160 160 161 161 
<< pdiffusion >>
rect 161 160 162 161 
<< m1 >>
rect 163 160 164 161 
<< m1 >>
rect 165 160 166 161 
<< m2 >>
rect 169 160 170 161 
<< m1 >>
rect 170 160 171 161 
<< m1 >>
rect 172 160 173 161 
<< pdiffusion >>
rect 174 160 175 161 
<< pdiffusion >>
rect 175 160 176 161 
<< pdiffusion >>
rect 176 160 177 161 
<< pdiffusion >>
rect 177 160 178 161 
<< pdiffusion >>
rect 178 160 179 161 
<< pdiffusion >>
rect 179 160 180 161 
<< m1 >>
rect 183 160 184 161 
<< m2 >>
rect 187 160 188 161 
<< m1 >>
rect 188 160 189 161 
<< m1 >>
rect 190 160 191 161 
<< pdiffusion >>
rect 192 160 193 161 
<< pdiffusion >>
rect 193 160 194 161 
<< pdiffusion >>
rect 194 160 195 161 
<< pdiffusion >>
rect 195 160 196 161 
<< pdiffusion >>
rect 196 160 197 161 
<< pdiffusion >>
rect 197 160 198 161 
<< m1 >>
rect 199 160 200 161 
<< pdiffusion >>
rect 210 160 211 161 
<< pdiffusion >>
rect 211 160 212 161 
<< pdiffusion >>
rect 212 160 213 161 
<< pdiffusion >>
rect 213 160 214 161 
<< pdiffusion >>
rect 214 160 215 161 
<< pdiffusion >>
rect 215 160 216 161 
<< m2 >>
rect 225 160 226 161 
<< m1 >>
rect 226 160 227 161 
<< pdiffusion >>
rect 228 160 229 161 
<< pdiffusion >>
rect 229 160 230 161 
<< pdiffusion >>
rect 230 160 231 161 
<< pdiffusion >>
rect 231 160 232 161 
<< pdiffusion >>
rect 232 160 233 161 
<< pdiffusion >>
rect 233 160 234 161 
<< m1 >>
rect 235 160 236 161 
<< m1 >>
rect 237 160 238 161 
<< m2 >>
rect 238 160 239 161 
<< m1 >>
rect 240 160 241 161 
<< pdiffusion >>
rect 246 160 247 161 
<< pdiffusion >>
rect 247 160 248 161 
<< pdiffusion >>
rect 248 160 249 161 
<< pdiffusion >>
rect 249 160 250 161 
<< pdiffusion >>
rect 250 160 251 161 
<< pdiffusion >>
rect 251 160 252 161 
<< m1 >>
rect 253 160 254 161 
<< m1 >>
rect 255 160 256 161 
<< m1 >>
rect 260 160 261 161 
<< m1 >>
rect 262 160 263 161 
<< m2 >>
rect 262 160 263 161 
<< pdiffusion >>
rect 264 160 265 161 
<< pdiffusion >>
rect 265 160 266 161 
<< pdiffusion >>
rect 266 160 267 161 
<< pdiffusion >>
rect 267 160 268 161 
<< pdiffusion >>
rect 268 160 269 161 
<< pdiffusion >>
rect 269 160 270 161 
<< m1 >>
rect 272 160 273 161 
<< m1 >>
rect 274 160 275 161 
<< m2 >>
rect 275 160 276 161 
<< m1 >>
rect 276 160 277 161 
<< m1 >>
rect 280 160 281 161 
<< pdiffusion >>
rect 282 160 283 161 
<< pdiffusion >>
rect 283 160 284 161 
<< pdiffusion >>
rect 284 160 285 161 
<< pdiffusion >>
rect 285 160 286 161 
<< pdiffusion >>
rect 286 160 287 161 
<< pdiffusion >>
rect 287 160 288 161 
<< m1 >>
rect 296 160 297 161 
<< m1 >>
rect 298 160 299 161 
<< pdiffusion >>
rect 300 160 301 161 
<< pdiffusion >>
rect 301 160 302 161 
<< pdiffusion >>
rect 302 160 303 161 
<< pdiffusion >>
rect 303 160 304 161 
<< pdiffusion >>
rect 304 160 305 161 
<< pdiffusion >>
rect 305 160 306 161 
<< m1 >>
rect 307 160 308 161 
<< m2 >>
rect 308 160 309 161 
<< pdiffusion >>
rect 318 160 319 161 
<< pdiffusion >>
rect 319 160 320 161 
<< pdiffusion >>
rect 320 160 321 161 
<< pdiffusion >>
rect 321 160 322 161 
<< pdiffusion >>
rect 322 160 323 161 
<< pdiffusion >>
rect 323 160 324 161 
<< m1 >>
rect 327 160 328 161 
<< m1 >>
rect 329 160 330 161 
<< pdiffusion >>
rect 336 160 337 161 
<< pdiffusion >>
rect 337 160 338 161 
<< pdiffusion >>
rect 338 160 339 161 
<< pdiffusion >>
rect 339 160 340 161 
<< pdiffusion >>
rect 340 160 341 161 
<< pdiffusion >>
rect 341 160 342 161 
<< m1 >>
rect 343 160 344 161 
<< m2 >>
rect 343 160 344 161 
<< m1 >>
rect 345 160 346 161 
<< m1 >>
rect 10 161 11 162 
<< pdiffusion >>
rect 12 161 13 162 
<< pdiffusion >>
rect 13 161 14 162 
<< pdiffusion >>
rect 14 161 15 162 
<< pdiffusion >>
rect 15 161 16 162 
<< m1 >>
rect 16 161 17 162 
<< pdiffusion >>
rect 16 161 17 162 
<< pdiffusion >>
rect 17 161 18 162 
<< m1 >>
rect 19 161 20 162 
<< m2 >>
rect 19 161 20 162 
<< m1 >>
rect 21 161 22 162 
<< m1 >>
rect 23 161 24 162 
<< m2 >>
rect 27 161 28 162 
<< m1 >>
rect 28 161 29 162 
<< pdiffusion >>
rect 30 161 31 162 
<< pdiffusion >>
rect 31 161 32 162 
<< pdiffusion >>
rect 32 161 33 162 
<< pdiffusion >>
rect 33 161 34 162 
<< pdiffusion >>
rect 34 161 35 162 
<< pdiffusion >>
rect 35 161 36 162 
<< m1 >>
rect 37 161 38 162 
<< m2 >>
rect 38 161 39 162 
<< m1 >>
rect 44 161 45 162 
<< m1 >>
rect 46 161 47 162 
<< pdiffusion >>
rect 48 161 49 162 
<< m1 >>
rect 49 161 50 162 
<< pdiffusion >>
rect 49 161 50 162 
<< pdiffusion >>
rect 50 161 51 162 
<< pdiffusion >>
rect 51 161 52 162 
<< pdiffusion >>
rect 52 161 53 162 
<< pdiffusion >>
rect 53 161 54 162 
<< m1 >>
rect 56 161 57 162 
<< m1 >>
rect 58 161 59 162 
<< m1 >>
rect 60 161 61 162 
<< m1 >>
rect 62 161 63 162 
<< m1 >>
rect 64 161 65 162 
<< pdiffusion >>
rect 66 161 67 162 
<< pdiffusion >>
rect 67 161 68 162 
<< pdiffusion >>
rect 68 161 69 162 
<< pdiffusion >>
rect 69 161 70 162 
<< pdiffusion >>
rect 70 161 71 162 
<< pdiffusion >>
rect 71 161 72 162 
<< m1 >>
rect 82 161 83 162 
<< pdiffusion >>
rect 84 161 85 162 
<< pdiffusion >>
rect 85 161 86 162 
<< pdiffusion >>
rect 86 161 87 162 
<< pdiffusion >>
rect 87 161 88 162 
<< pdiffusion >>
rect 88 161 89 162 
<< pdiffusion >>
rect 89 161 90 162 
<< m1 >>
rect 91 161 92 162 
<< m2 >>
rect 92 161 93 162 
<< pdiffusion >>
rect 102 161 103 162 
<< m1 >>
rect 103 161 104 162 
<< pdiffusion >>
rect 103 161 104 162 
<< pdiffusion >>
rect 104 161 105 162 
<< pdiffusion >>
rect 105 161 106 162 
<< pdiffusion >>
rect 106 161 107 162 
<< pdiffusion >>
rect 107 161 108 162 
<< pdiffusion >>
rect 120 161 121 162 
<< pdiffusion >>
rect 121 161 122 162 
<< pdiffusion >>
rect 122 161 123 162 
<< pdiffusion >>
rect 123 161 124 162 
<< pdiffusion >>
rect 124 161 125 162 
<< pdiffusion >>
rect 125 161 126 162 
<< m1 >>
rect 130 161 131 162 
<< m1 >>
rect 132 161 133 162 
<< m1 >>
rect 136 161 137 162 
<< m2 >>
rect 136 161 137 162 
<< pdiffusion >>
rect 138 161 139 162 
<< pdiffusion >>
rect 139 161 140 162 
<< pdiffusion >>
rect 140 161 141 162 
<< pdiffusion >>
rect 141 161 142 162 
<< pdiffusion >>
rect 142 161 143 162 
<< pdiffusion >>
rect 143 161 144 162 
<< m1 >>
rect 145 161 146 162 
<< m2 >>
rect 145 161 146 162 
<< m1 >>
rect 154 161 155 162 
<< pdiffusion >>
rect 156 161 157 162 
<< pdiffusion >>
rect 157 161 158 162 
<< pdiffusion >>
rect 158 161 159 162 
<< pdiffusion >>
rect 159 161 160 162 
<< pdiffusion >>
rect 160 161 161 162 
<< pdiffusion >>
rect 161 161 162 162 
<< m1 >>
rect 163 161 164 162 
<< m1 >>
rect 165 161 166 162 
<< m2 >>
rect 169 161 170 162 
<< m1 >>
rect 170 161 171 162 
<< m1 >>
rect 172 161 173 162 
<< pdiffusion >>
rect 174 161 175 162 
<< pdiffusion >>
rect 175 161 176 162 
<< pdiffusion >>
rect 176 161 177 162 
<< pdiffusion >>
rect 177 161 178 162 
<< pdiffusion >>
rect 178 161 179 162 
<< pdiffusion >>
rect 179 161 180 162 
<< m1 >>
rect 183 161 184 162 
<< m2 >>
rect 187 161 188 162 
<< m1 >>
rect 188 161 189 162 
<< m1 >>
rect 190 161 191 162 
<< pdiffusion >>
rect 192 161 193 162 
<< pdiffusion >>
rect 193 161 194 162 
<< pdiffusion >>
rect 194 161 195 162 
<< pdiffusion >>
rect 195 161 196 162 
<< m1 >>
rect 196 161 197 162 
<< pdiffusion >>
rect 196 161 197 162 
<< pdiffusion >>
rect 197 161 198 162 
<< m1 >>
rect 199 161 200 162 
<< pdiffusion >>
rect 210 161 211 162 
<< m1 >>
rect 211 161 212 162 
<< pdiffusion >>
rect 211 161 212 162 
<< pdiffusion >>
rect 212 161 213 162 
<< pdiffusion >>
rect 213 161 214 162 
<< pdiffusion >>
rect 214 161 215 162 
<< pdiffusion >>
rect 215 161 216 162 
<< m2 >>
rect 225 161 226 162 
<< m1 >>
rect 226 161 227 162 
<< pdiffusion >>
rect 228 161 229 162 
<< pdiffusion >>
rect 229 161 230 162 
<< pdiffusion >>
rect 230 161 231 162 
<< pdiffusion >>
rect 231 161 232 162 
<< pdiffusion >>
rect 232 161 233 162 
<< pdiffusion >>
rect 233 161 234 162 
<< m1 >>
rect 235 161 236 162 
<< m1 >>
rect 237 161 238 162 
<< m2 >>
rect 238 161 239 162 
<< m1 >>
rect 240 161 241 162 
<< pdiffusion >>
rect 246 161 247 162 
<< pdiffusion >>
rect 247 161 248 162 
<< pdiffusion >>
rect 248 161 249 162 
<< pdiffusion >>
rect 249 161 250 162 
<< pdiffusion >>
rect 250 161 251 162 
<< pdiffusion >>
rect 251 161 252 162 
<< m1 >>
rect 253 161 254 162 
<< m1 >>
rect 255 161 256 162 
<< m1 >>
rect 260 161 261 162 
<< m1 >>
rect 262 161 263 162 
<< m2 >>
rect 262 161 263 162 
<< pdiffusion >>
rect 264 161 265 162 
<< pdiffusion >>
rect 265 161 266 162 
<< pdiffusion >>
rect 266 161 267 162 
<< pdiffusion >>
rect 267 161 268 162 
<< pdiffusion >>
rect 268 161 269 162 
<< pdiffusion >>
rect 269 161 270 162 
<< m1 >>
rect 272 161 273 162 
<< m1 >>
rect 274 161 275 162 
<< m2 >>
rect 275 161 276 162 
<< m1 >>
rect 276 161 277 162 
<< m1 >>
rect 280 161 281 162 
<< pdiffusion >>
rect 282 161 283 162 
<< pdiffusion >>
rect 283 161 284 162 
<< pdiffusion >>
rect 284 161 285 162 
<< pdiffusion >>
rect 285 161 286 162 
<< pdiffusion >>
rect 286 161 287 162 
<< pdiffusion >>
rect 287 161 288 162 
<< m1 >>
rect 296 161 297 162 
<< m1 >>
rect 298 161 299 162 
<< pdiffusion >>
rect 300 161 301 162 
<< pdiffusion >>
rect 301 161 302 162 
<< pdiffusion >>
rect 302 161 303 162 
<< pdiffusion >>
rect 303 161 304 162 
<< m1 >>
rect 304 161 305 162 
<< pdiffusion >>
rect 304 161 305 162 
<< pdiffusion >>
rect 305 161 306 162 
<< m1 >>
rect 307 161 308 162 
<< m2 >>
rect 308 161 309 162 
<< pdiffusion >>
rect 318 161 319 162 
<< pdiffusion >>
rect 319 161 320 162 
<< pdiffusion >>
rect 320 161 321 162 
<< pdiffusion >>
rect 321 161 322 162 
<< pdiffusion >>
rect 322 161 323 162 
<< pdiffusion >>
rect 323 161 324 162 
<< m1 >>
rect 327 161 328 162 
<< m1 >>
rect 329 161 330 162 
<< pdiffusion >>
rect 336 161 337 162 
<< pdiffusion >>
rect 337 161 338 162 
<< pdiffusion >>
rect 338 161 339 162 
<< pdiffusion >>
rect 339 161 340 162 
<< m1 >>
rect 340 161 341 162 
<< pdiffusion >>
rect 340 161 341 162 
<< pdiffusion >>
rect 341 161 342 162 
<< m1 >>
rect 343 161 344 162 
<< m2 >>
rect 343 161 344 162 
<< m1 >>
rect 345 161 346 162 
<< m1 >>
rect 10 162 11 163 
<< m1 >>
rect 16 162 17 163 
<< m1 >>
rect 19 162 20 163 
<< m2 >>
rect 19 162 20 163 
<< m1 >>
rect 21 162 22 163 
<< m1 >>
rect 23 162 24 163 
<< m2 >>
rect 27 162 28 163 
<< m1 >>
rect 28 162 29 163 
<< m1 >>
rect 37 162 38 163 
<< m2 >>
rect 38 162 39 163 
<< m1 >>
rect 44 162 45 163 
<< m1 >>
rect 46 162 47 163 
<< m1 >>
rect 49 162 50 163 
<< m1 >>
rect 56 162 57 163 
<< m2 >>
rect 56 162 57 163 
<< m2c >>
rect 56 162 57 163 
<< m1 >>
rect 56 162 57 163 
<< m2 >>
rect 56 162 57 163 
<< m1 >>
rect 58 162 59 163 
<< m2 >>
rect 58 162 59 163 
<< m2c >>
rect 58 162 59 163 
<< m1 >>
rect 58 162 59 163 
<< m2 >>
rect 58 162 59 163 
<< m1 >>
rect 60 162 61 163 
<< m2 >>
rect 60 162 61 163 
<< m2c >>
rect 60 162 61 163 
<< m1 >>
rect 60 162 61 163 
<< m2 >>
rect 60 162 61 163 
<< m1 >>
rect 62 162 63 163 
<< m2 >>
rect 62 162 63 163 
<< m2c >>
rect 62 162 63 163 
<< m1 >>
rect 62 162 63 163 
<< m2 >>
rect 62 162 63 163 
<< m1 >>
rect 64 162 65 163 
<< m2 >>
rect 64 162 65 163 
<< m2c >>
rect 64 162 65 163 
<< m1 >>
rect 64 162 65 163 
<< m2 >>
rect 64 162 65 163 
<< m1 >>
rect 82 162 83 163 
<< m1 >>
rect 91 162 92 163 
<< m2 >>
rect 92 162 93 163 
<< m1 >>
rect 103 162 104 163 
<< m1 >>
rect 130 162 131 163 
<< m1 >>
rect 132 162 133 163 
<< m1 >>
rect 136 162 137 163 
<< m2 >>
rect 136 162 137 163 
<< m1 >>
rect 145 162 146 163 
<< m2 >>
rect 145 162 146 163 
<< m1 >>
rect 154 162 155 163 
<< m1 >>
rect 163 162 164 163 
<< m1 >>
rect 165 162 166 163 
<< m2 >>
rect 169 162 170 163 
<< m1 >>
rect 170 162 171 163 
<< m1 >>
rect 172 162 173 163 
<< m1 >>
rect 183 162 184 163 
<< m2 >>
rect 187 162 188 163 
<< m1 >>
rect 188 162 189 163 
<< m1 >>
rect 190 162 191 163 
<< m1 >>
rect 196 162 197 163 
<< m1 >>
rect 199 162 200 163 
<< m1 >>
rect 211 162 212 163 
<< m2 >>
rect 225 162 226 163 
<< m1 >>
rect 226 162 227 163 
<< m1 >>
rect 235 162 236 163 
<< m1 >>
rect 237 162 238 163 
<< m2 >>
rect 238 162 239 163 
<< m1 >>
rect 240 162 241 163 
<< m1 >>
rect 253 162 254 163 
<< m1 >>
rect 255 162 256 163 
<< m1 >>
rect 260 162 261 163 
<< m1 >>
rect 262 162 263 163 
<< m2 >>
rect 262 162 263 163 
<< m1 >>
rect 272 162 273 163 
<< m1 >>
rect 274 162 275 163 
<< m2 >>
rect 275 162 276 163 
<< m1 >>
rect 276 162 277 163 
<< m1 >>
rect 280 162 281 163 
<< m1 >>
rect 296 162 297 163 
<< m1 >>
rect 298 162 299 163 
<< m1 >>
rect 304 162 305 163 
<< m1 >>
rect 307 162 308 163 
<< m2 >>
rect 308 162 309 163 
<< m1 >>
rect 327 162 328 163 
<< m1 >>
rect 329 162 330 163 
<< m1 >>
rect 340 162 341 163 
<< m1 >>
rect 343 162 344 163 
<< m2 >>
rect 343 162 344 163 
<< m1 >>
rect 345 162 346 163 
<< m1 >>
rect 10 163 11 164 
<< m1 >>
rect 16 163 17 164 
<< m1 >>
rect 17 163 18 164 
<< m1 >>
rect 18 163 19 164 
<< m1 >>
rect 19 163 20 164 
<< m2 >>
rect 19 163 20 164 
<< m1 >>
rect 21 163 22 164 
<< m1 >>
rect 23 163 24 164 
<< m2 >>
rect 27 163 28 164 
<< m1 >>
rect 28 163 29 164 
<< m1 >>
rect 37 163 38 164 
<< m2 >>
rect 38 163 39 164 
<< m1 >>
rect 44 163 45 164 
<< m1 >>
rect 46 163 47 164 
<< m1 >>
rect 49 163 50 164 
<< m2 >>
rect 56 163 57 164 
<< m2 >>
rect 58 163 59 164 
<< m2 >>
rect 60 163 61 164 
<< m2 >>
rect 62 163 63 164 
<< m2 >>
rect 64 163 65 164 
<< m1 >>
rect 82 163 83 164 
<< m1 >>
rect 89 163 90 164 
<< m2 >>
rect 89 163 90 164 
<< m2c >>
rect 89 163 90 164 
<< m1 >>
rect 89 163 90 164 
<< m2 >>
rect 89 163 90 164 
<< m2 >>
rect 90 163 91 164 
<< m1 >>
rect 91 163 92 164 
<< m2 >>
rect 91 163 92 164 
<< m2 >>
rect 92 163 93 164 
<< m1 >>
rect 103 163 104 164 
<< m1 >>
rect 130 163 131 164 
<< m1 >>
rect 132 163 133 164 
<< m1 >>
rect 136 163 137 164 
<< m2 >>
rect 136 163 137 164 
<< m1 >>
rect 145 163 146 164 
<< m2 >>
rect 145 163 146 164 
<< m1 >>
rect 154 163 155 164 
<< m1 >>
rect 163 163 164 164 
<< m1 >>
rect 165 163 166 164 
<< m2 >>
rect 169 163 170 164 
<< m1 >>
rect 170 163 171 164 
<< m2 >>
rect 170 163 171 164 
<< m2 >>
rect 171 163 172 164 
<< m1 >>
rect 172 163 173 164 
<< m2 >>
rect 172 163 173 164 
<< m2 >>
rect 173 163 174 164 
<< m1 >>
rect 174 163 175 164 
<< m2 >>
rect 174 163 175 164 
<< m2c >>
rect 174 163 175 164 
<< m1 >>
rect 174 163 175 164 
<< m2 >>
rect 174 163 175 164 
<< m1 >>
rect 183 163 184 164 
<< m2 >>
rect 187 163 188 164 
<< m1 >>
rect 188 163 189 164 
<< m2 >>
rect 188 163 189 164 
<< m2 >>
rect 189 163 190 164 
<< m1 >>
rect 190 163 191 164 
<< m2 >>
rect 190 163 191 164 
<< m2 >>
rect 191 163 192 164 
<< m1 >>
rect 192 163 193 164 
<< m2 >>
rect 192 163 193 164 
<< m2c >>
rect 192 163 193 164 
<< m1 >>
rect 192 163 193 164 
<< m2 >>
rect 192 163 193 164 
<< m1 >>
rect 196 163 197 164 
<< m1 >>
rect 199 163 200 164 
<< m1 >>
rect 211 163 212 164 
<< m2 >>
rect 225 163 226 164 
<< m1 >>
rect 226 163 227 164 
<< m1 >>
rect 235 163 236 164 
<< m1 >>
rect 237 163 238 164 
<< m2 >>
rect 238 163 239 164 
<< m1 >>
rect 240 163 241 164 
<< m1 >>
rect 253 163 254 164 
<< m1 >>
rect 255 163 256 164 
<< m1 >>
rect 260 163 261 164 
<< m1 >>
rect 262 163 263 164 
<< m2 >>
rect 262 163 263 164 
<< m2 >>
rect 263 163 264 164 
<< m1 >>
rect 264 163 265 164 
<< m2 >>
rect 264 163 265 164 
<< m2c >>
rect 264 163 265 164 
<< m1 >>
rect 264 163 265 164 
<< m2 >>
rect 264 163 265 164 
<< m1 >>
rect 272 163 273 164 
<< m1 >>
rect 274 163 275 164 
<< m2 >>
rect 275 163 276 164 
<< m1 >>
rect 276 163 277 164 
<< m1 >>
rect 280 163 281 164 
<< m1 >>
rect 296 163 297 164 
<< m1 >>
rect 298 163 299 164 
<< m1 >>
rect 304 163 305 164 
<< m1 >>
rect 307 163 308 164 
<< m2 >>
rect 308 163 309 164 
<< m1 >>
rect 327 163 328 164 
<< m1 >>
rect 329 163 330 164 
<< m1 >>
rect 340 163 341 164 
<< m1 >>
rect 343 163 344 164 
<< m2 >>
rect 343 163 344 164 
<< m1 >>
rect 345 163 346 164 
<< m1 >>
rect 10 164 11 165 
<< m2 >>
rect 19 164 20 165 
<< m1 >>
rect 21 164 22 165 
<< m1 >>
rect 23 164 24 165 
<< m2 >>
rect 27 164 28 165 
<< m1 >>
rect 28 164 29 165 
<< m1 >>
rect 37 164 38 165 
<< m2 >>
rect 38 164 39 165 
<< m1 >>
rect 44 164 45 165 
<< m1 >>
rect 46 164 47 165 
<< m1 >>
rect 49 164 50 165 
<< m1 >>
rect 50 164 51 165 
<< m1 >>
rect 51 164 52 165 
<< m1 >>
rect 52 164 53 165 
<< m1 >>
rect 53 164 54 165 
<< m1 >>
rect 54 164 55 165 
<< m1 >>
rect 55 164 56 165 
<< m1 >>
rect 56 164 57 165 
<< m2 >>
rect 56 164 57 165 
<< m1 >>
rect 57 164 58 165 
<< m1 >>
rect 58 164 59 165 
<< m2 >>
rect 58 164 59 165 
<< m1 >>
rect 59 164 60 165 
<< m1 >>
rect 60 164 61 165 
<< m2 >>
rect 60 164 61 165 
<< m1 >>
rect 61 164 62 165 
<< m1 >>
rect 62 164 63 165 
<< m2 >>
rect 62 164 63 165 
<< m1 >>
rect 63 164 64 165 
<< m1 >>
rect 64 164 65 165 
<< m2 >>
rect 64 164 65 165 
<< m1 >>
rect 65 164 66 165 
<< m1 >>
rect 66 164 67 165 
<< m2 >>
rect 66 164 67 165 
<< m2c >>
rect 66 164 67 165 
<< m1 >>
rect 66 164 67 165 
<< m2 >>
rect 66 164 67 165 
<< m1 >>
rect 82 164 83 165 
<< m1 >>
rect 83 164 84 165 
<< m1 >>
rect 84 164 85 165 
<< m2 >>
rect 84 164 85 165 
<< m2c >>
rect 84 164 85 165 
<< m1 >>
rect 84 164 85 165 
<< m2 >>
rect 84 164 85 165 
<< m1 >>
rect 89 164 90 165 
<< m1 >>
rect 91 164 92 165 
<< m1 >>
rect 103 164 104 165 
<< m1 >>
rect 130 164 131 165 
<< m1 >>
rect 132 164 133 165 
<< m1 >>
rect 136 164 137 165 
<< m2 >>
rect 136 164 137 165 
<< m1 >>
rect 145 164 146 165 
<< m2 >>
rect 145 164 146 165 
<< m1 >>
rect 154 164 155 165 
<< m1 >>
rect 163 164 164 165 
<< m1 >>
rect 165 164 166 165 
<< m1 >>
rect 170 164 171 165 
<< m1 >>
rect 172 164 173 165 
<< m1 >>
rect 174 164 175 165 
<< m1 >>
rect 183 164 184 165 
<< m1 >>
rect 188 164 189 165 
<< m1 >>
rect 190 164 191 165 
<< m1 >>
rect 192 164 193 165 
<< m1 >>
rect 196 164 197 165 
<< m1 >>
rect 199 164 200 165 
<< m1 >>
rect 211 164 212 165 
<< m2 >>
rect 225 164 226 165 
<< m1 >>
rect 226 164 227 165 
<< m1 >>
rect 235 164 236 165 
<< m1 >>
rect 237 164 238 165 
<< m2 >>
rect 238 164 239 165 
<< m1 >>
rect 240 164 241 165 
<< m1 >>
rect 253 164 254 165 
<< m1 >>
rect 255 164 256 165 
<< m1 >>
rect 260 164 261 165 
<< m1 >>
rect 262 164 263 165 
<< m1 >>
rect 264 164 265 165 
<< m1 >>
rect 272 164 273 165 
<< m1 >>
rect 274 164 275 165 
<< m2 >>
rect 275 164 276 165 
<< m1 >>
rect 276 164 277 165 
<< m1 >>
rect 280 164 281 165 
<< m2 >>
rect 280 164 281 165 
<< m2c >>
rect 280 164 281 165 
<< m1 >>
rect 280 164 281 165 
<< m2 >>
rect 280 164 281 165 
<< m1 >>
rect 296 164 297 165 
<< m2 >>
rect 296 164 297 165 
<< m2c >>
rect 296 164 297 165 
<< m1 >>
rect 296 164 297 165 
<< m2 >>
rect 296 164 297 165 
<< m1 >>
rect 298 164 299 165 
<< m2 >>
rect 298 164 299 165 
<< m2c >>
rect 298 164 299 165 
<< m1 >>
rect 298 164 299 165 
<< m2 >>
rect 298 164 299 165 
<< m1 >>
rect 304 164 305 165 
<< m1 >>
rect 307 164 308 165 
<< m2 >>
rect 308 164 309 165 
<< m1 >>
rect 327 164 328 165 
<< m1 >>
rect 329 164 330 165 
<< m1 >>
rect 338 164 339 165 
<< m2 >>
rect 338 164 339 165 
<< m2c >>
rect 338 164 339 165 
<< m1 >>
rect 338 164 339 165 
<< m2 >>
rect 338 164 339 165 
<< m1 >>
rect 339 164 340 165 
<< m1 >>
rect 340 164 341 165 
<< m1 >>
rect 343 164 344 165 
<< m2 >>
rect 343 164 344 165 
<< m1 >>
rect 345 164 346 165 
<< m1 >>
rect 10 165 11 166 
<< m1 >>
rect 19 165 20 166 
<< m2 >>
rect 19 165 20 166 
<< m2c >>
rect 19 165 20 166 
<< m1 >>
rect 19 165 20 166 
<< m2 >>
rect 19 165 20 166 
<< m1 >>
rect 21 165 22 166 
<< m1 >>
rect 23 165 24 166 
<< m2 >>
rect 27 165 28 166 
<< m1 >>
rect 28 165 29 166 
<< m1 >>
rect 37 165 38 166 
<< m2 >>
rect 38 165 39 166 
<< m1 >>
rect 44 165 45 166 
<< m1 >>
rect 46 165 47 166 
<< m2 >>
rect 56 165 57 166 
<< m2 >>
rect 58 165 59 166 
<< m2 >>
rect 60 165 61 166 
<< m2 >>
rect 62 165 63 166 
<< m2 >>
rect 64 165 65 166 
<< m2 >>
rect 66 165 67 166 
<< m2 >>
rect 84 165 85 166 
<< m1 >>
rect 89 165 90 166 
<< m1 >>
rect 91 165 92 166 
<< m1 >>
rect 103 165 104 166 
<< m1 >>
rect 130 165 131 166 
<< m1 >>
rect 132 165 133 166 
<< m1 >>
rect 136 165 137 166 
<< m2 >>
rect 136 165 137 166 
<< m1 >>
rect 145 165 146 166 
<< m2 >>
rect 145 165 146 166 
<< m1 >>
rect 154 165 155 166 
<< m1 >>
rect 163 165 164 166 
<< m1 >>
rect 165 165 166 166 
<< m1 >>
rect 170 165 171 166 
<< m1 >>
rect 172 165 173 166 
<< m1 >>
rect 174 165 175 166 
<< m1 >>
rect 183 165 184 166 
<< m1 >>
rect 188 165 189 166 
<< m1 >>
rect 190 165 191 166 
<< m1 >>
rect 192 165 193 166 
<< m1 >>
rect 196 165 197 166 
<< m1 >>
rect 199 165 200 166 
<< m1 >>
rect 211 165 212 166 
<< m2 >>
rect 225 165 226 166 
<< m1 >>
rect 226 165 227 166 
<< m1 >>
rect 235 165 236 166 
<< m1 >>
rect 237 165 238 166 
<< m2 >>
rect 238 165 239 166 
<< m1 >>
rect 240 165 241 166 
<< m1 >>
rect 253 165 254 166 
<< m1 >>
rect 255 165 256 166 
<< m1 >>
rect 260 165 261 166 
<< m1 >>
rect 262 165 263 166 
<< m1 >>
rect 264 165 265 166 
<< m1 >>
rect 272 165 273 166 
<< m1 >>
rect 274 165 275 166 
<< m2 >>
rect 275 165 276 166 
<< m1 >>
rect 276 165 277 166 
<< m2 >>
rect 280 165 281 166 
<< m2 >>
rect 296 165 297 166 
<< m2 >>
rect 298 165 299 166 
<< m1 >>
rect 304 165 305 166 
<< m1 >>
rect 307 165 308 166 
<< m2 >>
rect 308 165 309 166 
<< m1 >>
rect 327 165 328 166 
<< m1 >>
rect 329 165 330 166 
<< m2 >>
rect 338 165 339 166 
<< m1 >>
rect 343 165 344 166 
<< m2 >>
rect 343 165 344 166 
<< m1 >>
rect 345 165 346 166 
<< m1 >>
rect 10 166 11 167 
<< m1 >>
rect 19 166 20 167 
<< m1 >>
rect 21 166 22 167 
<< m1 >>
rect 23 166 24 167 
<< m2 >>
rect 27 166 28 167 
<< m1 >>
rect 28 166 29 167 
<< m1 >>
rect 37 166 38 167 
<< m2 >>
rect 38 166 39 167 
<< m1 >>
rect 44 166 45 167 
<< m1 >>
rect 46 166 47 167 
<< m1 >>
rect 49 166 50 167 
<< m1 >>
rect 50 166 51 167 
<< m1 >>
rect 51 166 52 167 
<< m1 >>
rect 52 166 53 167 
<< m1 >>
rect 53 166 54 167 
<< m1 >>
rect 54 166 55 167 
<< m1 >>
rect 55 166 56 167 
<< m1 >>
rect 56 166 57 167 
<< m2 >>
rect 56 166 57 167 
<< m1 >>
rect 57 166 58 167 
<< m1 >>
rect 58 166 59 167 
<< m2 >>
rect 58 166 59 167 
<< m1 >>
rect 59 166 60 167 
<< m1 >>
rect 60 166 61 167 
<< m2 >>
rect 60 166 61 167 
<< m1 >>
rect 61 166 62 167 
<< m1 >>
rect 62 166 63 167 
<< m2 >>
rect 62 166 63 167 
<< m1 >>
rect 63 166 64 167 
<< m1 >>
rect 64 166 65 167 
<< m2 >>
rect 64 166 65 167 
<< m1 >>
rect 65 166 66 167 
<< m1 >>
rect 66 166 67 167 
<< m2 >>
rect 66 166 67 167 
<< m1 >>
rect 67 166 68 167 
<< m1 >>
rect 68 166 69 167 
<< m1 >>
rect 69 166 70 167 
<< m1 >>
rect 70 166 71 167 
<< m1 >>
rect 71 166 72 167 
<< m1 >>
rect 72 166 73 167 
<< m1 >>
rect 73 166 74 167 
<< m1 >>
rect 74 166 75 167 
<< m1 >>
rect 75 166 76 167 
<< m1 >>
rect 76 166 77 167 
<< m1 >>
rect 77 166 78 167 
<< m1 >>
rect 78 166 79 167 
<< m1 >>
rect 79 166 80 167 
<< m1 >>
rect 80 166 81 167 
<< m1 >>
rect 81 166 82 167 
<< m1 >>
rect 82 166 83 167 
<< m1 >>
rect 83 166 84 167 
<< m1 >>
rect 84 166 85 167 
<< m2 >>
rect 84 166 85 167 
<< m1 >>
rect 85 166 86 167 
<< m1 >>
rect 86 166 87 167 
<< m1 >>
rect 87 166 88 167 
<< m1 >>
rect 88 166 89 167 
<< m1 >>
rect 89 166 90 167 
<< m1 >>
rect 91 166 92 167 
<< m1 >>
rect 103 166 104 167 
<< m1 >>
rect 104 166 105 167 
<< m1 >>
rect 105 166 106 167 
<< m1 >>
rect 106 166 107 167 
<< m1 >>
rect 107 166 108 167 
<< m1 >>
rect 108 166 109 167 
<< m1 >>
rect 109 166 110 167 
<< m1 >>
rect 110 166 111 167 
<< m1 >>
rect 111 166 112 167 
<< m1 >>
rect 112 166 113 167 
<< m1 >>
rect 113 166 114 167 
<< m1 >>
rect 114 166 115 167 
<< m1 >>
rect 115 166 116 167 
<< m1 >>
rect 116 166 117 167 
<< m1 >>
rect 117 166 118 167 
<< m1 >>
rect 118 166 119 167 
<< m1 >>
rect 119 166 120 167 
<< m1 >>
rect 120 166 121 167 
<< m1 >>
rect 121 166 122 167 
<< m1 >>
rect 122 166 123 167 
<< m1 >>
rect 123 166 124 167 
<< m1 >>
rect 124 166 125 167 
<< m1 >>
rect 125 166 126 167 
<< m1 >>
rect 126 166 127 167 
<< m1 >>
rect 127 166 128 167 
<< m1 >>
rect 130 166 131 167 
<< m1 >>
rect 132 166 133 167 
<< m1 >>
rect 136 166 137 167 
<< m2 >>
rect 136 166 137 167 
<< m1 >>
rect 145 166 146 167 
<< m2 >>
rect 145 166 146 167 
<< m1 >>
rect 154 166 155 167 
<< m1 >>
rect 155 166 156 167 
<< m1 >>
rect 156 166 157 167 
<< m1 >>
rect 157 166 158 167 
<< m1 >>
rect 158 166 159 167 
<< m1 >>
rect 159 166 160 167 
<< m1 >>
rect 160 166 161 167 
<< m1 >>
rect 163 166 164 167 
<< m1 >>
rect 165 166 166 167 
<< m1 >>
rect 170 166 171 167 
<< m1 >>
rect 172 166 173 167 
<< m1 >>
rect 174 166 175 167 
<< m1 >>
rect 183 166 184 167 
<< m1 >>
rect 188 166 189 167 
<< m1 >>
rect 190 166 191 167 
<< m1 >>
rect 192 166 193 167 
<< m1 >>
rect 193 166 194 167 
<< m1 >>
rect 194 166 195 167 
<< m2 >>
rect 194 166 195 167 
<< m2c >>
rect 194 166 195 167 
<< m1 >>
rect 194 166 195 167 
<< m2 >>
rect 194 166 195 167 
<< m2 >>
rect 195 166 196 167 
<< m1 >>
rect 196 166 197 167 
<< m2 >>
rect 196 166 197 167 
<< m2 >>
rect 197 166 198 167 
<< m2 >>
rect 198 166 199 167 
<< m1 >>
rect 199 166 200 167 
<< m2 >>
rect 199 166 200 167 
<< m2 >>
rect 200 166 201 167 
<< m1 >>
rect 201 166 202 167 
<< m2 >>
rect 201 166 202 167 
<< m2c >>
rect 201 166 202 167 
<< m1 >>
rect 201 166 202 167 
<< m2 >>
rect 201 166 202 167 
<< m1 >>
rect 202 166 203 167 
<< m1 >>
rect 203 166 204 167 
<< m1 >>
rect 204 166 205 167 
<< m1 >>
rect 205 166 206 167 
<< m1 >>
rect 206 166 207 167 
<< m1 >>
rect 207 166 208 167 
<< m1 >>
rect 208 166 209 167 
<< m1 >>
rect 209 166 210 167 
<< m1 >>
rect 210 166 211 167 
<< m1 >>
rect 211 166 212 167 
<< m2 >>
rect 225 166 226 167 
<< m1 >>
rect 226 166 227 167 
<< m1 >>
rect 235 166 236 167 
<< m1 >>
rect 237 166 238 167 
<< m2 >>
rect 238 166 239 167 
<< m1 >>
rect 240 166 241 167 
<< m1 >>
rect 253 166 254 167 
<< m1 >>
rect 255 166 256 167 
<< m1 >>
rect 260 166 261 167 
<< m1 >>
rect 262 166 263 167 
<< m1 >>
rect 264 166 265 167 
<< m1 >>
rect 265 166 266 167 
<< m1 >>
rect 266 166 267 167 
<< m1 >>
rect 267 166 268 167 
<< m1 >>
rect 268 166 269 167 
<< m1 >>
rect 269 166 270 167 
<< m1 >>
rect 270 166 271 167 
<< m2 >>
rect 270 166 271 167 
<< m2c >>
rect 270 166 271 167 
<< m1 >>
rect 270 166 271 167 
<< m2 >>
rect 270 166 271 167 
<< m2 >>
rect 271 166 272 167 
<< m1 >>
rect 272 166 273 167 
<< m1 >>
rect 274 166 275 167 
<< m2 >>
rect 275 166 276 167 
<< m1 >>
rect 276 166 277 167 
<< m1 >>
rect 277 166 278 167 
<< m1 >>
rect 278 166 279 167 
<< m1 >>
rect 279 166 280 167 
<< m1 >>
rect 280 166 281 167 
<< m2 >>
rect 280 166 281 167 
<< m1 >>
rect 281 166 282 167 
<< m1 >>
rect 282 166 283 167 
<< m1 >>
rect 283 166 284 167 
<< m1 >>
rect 284 166 285 167 
<< m1 >>
rect 285 166 286 167 
<< m1 >>
rect 286 166 287 167 
<< m1 >>
rect 287 166 288 167 
<< m1 >>
rect 288 166 289 167 
<< m1 >>
rect 289 166 290 167 
<< m1 >>
rect 290 166 291 167 
<< m1 >>
rect 291 166 292 167 
<< m1 >>
rect 292 166 293 167 
<< m1 >>
rect 293 166 294 167 
<< m1 >>
rect 294 166 295 167 
<< m1 >>
rect 295 166 296 167 
<< m1 >>
rect 296 166 297 167 
<< m2 >>
rect 296 166 297 167 
<< m1 >>
rect 297 166 298 167 
<< m1 >>
rect 298 166 299 167 
<< m2 >>
rect 298 166 299 167 
<< m1 >>
rect 299 166 300 167 
<< m1 >>
rect 300 166 301 167 
<< m1 >>
rect 301 166 302 167 
<< m1 >>
rect 302 166 303 167 
<< m1 >>
rect 303 166 304 167 
<< m1 >>
rect 304 166 305 167 
<< m1 >>
rect 307 166 308 167 
<< m2 >>
rect 308 166 309 167 
<< m1 >>
rect 327 166 328 167 
<< m1 >>
rect 329 166 330 167 
<< m1 >>
rect 330 166 331 167 
<< m1 >>
rect 331 166 332 167 
<< m1 >>
rect 332 166 333 167 
<< m1 >>
rect 333 166 334 167 
<< m1 >>
rect 334 166 335 167 
<< m1 >>
rect 335 166 336 167 
<< m1 >>
rect 336 166 337 167 
<< m1 >>
rect 337 166 338 167 
<< m1 >>
rect 338 166 339 167 
<< m2 >>
rect 338 166 339 167 
<< m1 >>
rect 339 166 340 167 
<< m1 >>
rect 340 166 341 167 
<< m1 >>
rect 343 166 344 167 
<< m2 >>
rect 343 166 344 167 
<< m1 >>
rect 345 166 346 167 
<< m1 >>
rect 10 167 11 168 
<< m1 >>
rect 19 167 20 168 
<< m1 >>
rect 21 167 22 168 
<< m1 >>
rect 23 167 24 168 
<< m2 >>
rect 27 167 28 168 
<< m1 >>
rect 28 167 29 168 
<< m1 >>
rect 37 167 38 168 
<< m2 >>
rect 38 167 39 168 
<< m1 >>
rect 44 167 45 168 
<< m1 >>
rect 46 167 47 168 
<< m1 >>
rect 49 167 50 168 
<< m2 >>
rect 56 167 57 168 
<< m2 >>
rect 58 167 59 168 
<< m2 >>
rect 60 167 61 168 
<< m2 >>
rect 62 167 63 168 
<< m2 >>
rect 64 167 65 168 
<< m2 >>
rect 66 167 67 168 
<< m2 >>
rect 67 167 68 168 
<< m2 >>
rect 68 167 69 168 
<< m2 >>
rect 69 167 70 168 
<< m2 >>
rect 70 167 71 168 
<< m2 >>
rect 71 167 72 168 
<< m2 >>
rect 72 167 73 168 
<< m2 >>
rect 73 167 74 168 
<< m2 >>
rect 74 167 75 168 
<< m2 >>
rect 75 167 76 168 
<< m2 >>
rect 76 167 77 168 
<< m2 >>
rect 77 167 78 168 
<< m2 >>
rect 78 167 79 168 
<< m2 >>
rect 79 167 80 168 
<< m2 >>
rect 80 167 81 168 
<< m2 >>
rect 81 167 82 168 
<< m2 >>
rect 82 167 83 168 
<< m2 >>
rect 84 167 85 168 
<< m1 >>
rect 91 167 92 168 
<< m1 >>
rect 127 167 128 168 
<< m1 >>
rect 130 167 131 168 
<< m1 >>
rect 132 167 133 168 
<< m1 >>
rect 136 167 137 168 
<< m2 >>
rect 136 167 137 168 
<< m1 >>
rect 145 167 146 168 
<< m2 >>
rect 145 167 146 168 
<< m1 >>
rect 160 167 161 168 
<< m1 >>
rect 163 167 164 168 
<< m1 >>
rect 165 167 166 168 
<< m1 >>
rect 170 167 171 168 
<< m2 >>
rect 170 167 171 168 
<< m2c >>
rect 170 167 171 168 
<< m1 >>
rect 170 167 171 168 
<< m2 >>
rect 170 167 171 168 
<< m1 >>
rect 172 167 173 168 
<< m2 >>
rect 172 167 173 168 
<< m2c >>
rect 172 167 173 168 
<< m1 >>
rect 172 167 173 168 
<< m2 >>
rect 172 167 173 168 
<< m1 >>
rect 174 167 175 168 
<< m2 >>
rect 174 167 175 168 
<< m2c >>
rect 174 167 175 168 
<< m1 >>
rect 174 167 175 168 
<< m2 >>
rect 174 167 175 168 
<< m1 >>
rect 183 167 184 168 
<< m2 >>
rect 183 167 184 168 
<< m2c >>
rect 183 167 184 168 
<< m1 >>
rect 183 167 184 168 
<< m2 >>
rect 183 167 184 168 
<< m1 >>
rect 188 167 189 168 
<< m2 >>
rect 188 167 189 168 
<< m2c >>
rect 188 167 189 168 
<< m1 >>
rect 188 167 189 168 
<< m2 >>
rect 188 167 189 168 
<< m1 >>
rect 190 167 191 168 
<< m2 >>
rect 190 167 191 168 
<< m2c >>
rect 190 167 191 168 
<< m1 >>
rect 190 167 191 168 
<< m2 >>
rect 190 167 191 168 
<< m1 >>
rect 196 167 197 168 
<< m1 >>
rect 199 167 200 168 
<< m2 >>
rect 225 167 226 168 
<< m1 >>
rect 226 167 227 168 
<< m1 >>
rect 235 167 236 168 
<< m1 >>
rect 237 167 238 168 
<< m2 >>
rect 238 167 239 168 
<< m1 >>
rect 240 167 241 168 
<< m1 >>
rect 253 167 254 168 
<< m1 >>
rect 255 167 256 168 
<< m1 >>
rect 260 167 261 168 
<< m1 >>
rect 262 167 263 168 
<< m2 >>
rect 271 167 272 168 
<< m1 >>
rect 272 167 273 168 
<< m1 >>
rect 274 167 275 168 
<< m2 >>
rect 275 167 276 168 
<< m2 >>
rect 280 167 281 168 
<< m2 >>
rect 296 167 297 168 
<< m2 >>
rect 298 167 299 168 
<< m1 >>
rect 307 167 308 168 
<< m2 >>
rect 308 167 309 168 
<< m2 >>
rect 326 167 327 168 
<< m1 >>
rect 327 167 328 168 
<< m2 >>
rect 327 167 328 168 
<< m2 >>
rect 328 167 329 168 
<< m2 >>
rect 329 167 330 168 
<< m2 >>
rect 330 167 331 168 
<< m2 >>
rect 331 167 332 168 
<< m2 >>
rect 332 167 333 168 
<< m2 >>
rect 333 167 334 168 
<< m2 >>
rect 334 167 335 168 
<< m2 >>
rect 335 167 336 168 
<< m2 >>
rect 336 167 337 168 
<< m2 >>
rect 337 167 338 168 
<< m2 >>
rect 338 167 339 168 
<< m1 >>
rect 340 167 341 168 
<< m1 >>
rect 343 167 344 168 
<< m2 >>
rect 343 167 344 168 
<< m1 >>
rect 345 167 346 168 
<< m1 >>
rect 10 168 11 169 
<< m1 >>
rect 19 168 20 169 
<< m1 >>
rect 21 168 22 169 
<< m1 >>
rect 23 168 24 169 
<< m2 >>
rect 27 168 28 169 
<< m1 >>
rect 28 168 29 169 
<< m1 >>
rect 37 168 38 169 
<< m2 >>
rect 38 168 39 169 
<< m1 >>
rect 44 168 45 169 
<< m1 >>
rect 46 168 47 169 
<< m1 >>
rect 49 168 50 169 
<< m1 >>
rect 56 168 57 169 
<< m2 >>
rect 56 168 57 169 
<< m2c >>
rect 56 168 57 169 
<< m1 >>
rect 56 168 57 169 
<< m2 >>
rect 56 168 57 169 
<< m1 >>
rect 58 168 59 169 
<< m2 >>
rect 58 168 59 169 
<< m2c >>
rect 58 168 59 169 
<< m1 >>
rect 58 168 59 169 
<< m2 >>
rect 58 168 59 169 
<< m1 >>
rect 60 168 61 169 
<< m2 >>
rect 60 168 61 169 
<< m2c >>
rect 60 168 61 169 
<< m1 >>
rect 60 168 61 169 
<< m2 >>
rect 60 168 61 169 
<< m1 >>
rect 62 168 63 169 
<< m2 >>
rect 62 168 63 169 
<< m2c >>
rect 62 168 63 169 
<< m1 >>
rect 62 168 63 169 
<< m2 >>
rect 62 168 63 169 
<< m1 >>
rect 64 168 65 169 
<< m2 >>
rect 64 168 65 169 
<< m2c >>
rect 64 168 65 169 
<< m1 >>
rect 64 168 65 169 
<< m2 >>
rect 64 168 65 169 
<< m1 >>
rect 82 168 83 169 
<< m2 >>
rect 82 168 83 169 
<< m2c >>
rect 82 168 83 169 
<< m1 >>
rect 82 168 83 169 
<< m2 >>
rect 82 168 83 169 
<< m2 >>
rect 84 168 85 169 
<< m1 >>
rect 91 168 92 169 
<< m1 >>
rect 127 168 128 169 
<< m1 >>
rect 130 168 131 169 
<< m1 >>
rect 132 168 133 169 
<< m1 >>
rect 136 168 137 169 
<< m2 >>
rect 136 168 137 169 
<< m1 >>
rect 145 168 146 169 
<< m2 >>
rect 145 168 146 169 
<< m1 >>
rect 160 168 161 169 
<< m1 >>
rect 163 168 164 169 
<< m1 >>
rect 165 168 166 169 
<< m2 >>
rect 170 168 171 169 
<< m2 >>
rect 172 168 173 169 
<< m2 >>
rect 174 168 175 169 
<< m2 >>
rect 175 168 176 169 
<< m2 >>
rect 176 168 177 169 
<< m2 >>
rect 183 168 184 169 
<< m2 >>
rect 188 168 189 169 
<< m2 >>
rect 190 168 191 169 
<< m1 >>
rect 196 168 197 169 
<< m1 >>
rect 199 168 200 169 
<< m2 >>
rect 225 168 226 169 
<< m1 >>
rect 226 168 227 169 
<< m1 >>
rect 235 168 236 169 
<< m1 >>
rect 237 168 238 169 
<< m2 >>
rect 238 168 239 169 
<< m1 >>
rect 240 168 241 169 
<< m1 >>
rect 253 168 254 169 
<< m1 >>
rect 255 168 256 169 
<< m1 >>
rect 260 168 261 169 
<< m1 >>
rect 262 168 263 169 
<< m2 >>
rect 271 168 272 169 
<< m1 >>
rect 272 168 273 169 
<< m1 >>
rect 274 168 275 169 
<< m2 >>
rect 275 168 276 169 
<< m1 >>
rect 280 168 281 169 
<< m2 >>
rect 280 168 281 169 
<< m2c >>
rect 280 168 281 169 
<< m1 >>
rect 280 168 281 169 
<< m2 >>
rect 280 168 281 169 
<< m1 >>
rect 281 168 282 169 
<< m1 >>
rect 282 168 283 169 
<< m1 >>
rect 283 168 284 169 
<< m1 >>
rect 284 168 285 169 
<< m1 >>
rect 285 168 286 169 
<< m1 >>
rect 286 168 287 169 
<< m1 >>
rect 287 168 288 169 
<< m1 >>
rect 288 168 289 169 
<< m1 >>
rect 289 168 290 169 
<< m1 >>
rect 296 168 297 169 
<< m2 >>
rect 296 168 297 169 
<< m2c >>
rect 296 168 297 169 
<< m1 >>
rect 296 168 297 169 
<< m2 >>
rect 296 168 297 169 
<< m1 >>
rect 298 168 299 169 
<< m2 >>
rect 298 168 299 169 
<< m2c >>
rect 298 168 299 169 
<< m1 >>
rect 298 168 299 169 
<< m2 >>
rect 298 168 299 169 
<< m1 >>
rect 307 168 308 169 
<< m2 >>
rect 308 168 309 169 
<< m2 >>
rect 326 168 327 169 
<< m1 >>
rect 327 168 328 169 
<< m1 >>
rect 340 168 341 169 
<< m1 >>
rect 343 168 344 169 
<< m2 >>
rect 343 168 344 169 
<< m1 >>
rect 345 168 346 169 
<< m1 >>
rect 10 169 11 170 
<< m1 >>
rect 19 169 20 170 
<< m1 >>
rect 21 169 22 170 
<< m1 >>
rect 23 169 24 170 
<< m2 >>
rect 27 169 28 170 
<< m1 >>
rect 28 169 29 170 
<< m1 >>
rect 37 169 38 170 
<< m2 >>
rect 38 169 39 170 
<< m1 >>
rect 44 169 45 170 
<< m1 >>
rect 46 169 47 170 
<< m1 >>
rect 49 169 50 170 
<< m1 >>
rect 56 169 57 170 
<< m1 >>
rect 58 169 59 170 
<< m1 >>
rect 60 169 61 170 
<< m1 >>
rect 62 169 63 170 
<< m1 >>
rect 64 169 65 170 
<< m1 >>
rect 82 169 83 170 
<< m1 >>
rect 84 169 85 170 
<< m2 >>
rect 84 169 85 170 
<< m1 >>
rect 85 169 86 170 
<< m1 >>
rect 86 169 87 170 
<< m1 >>
rect 87 169 88 170 
<< m1 >>
rect 88 169 89 170 
<< m1 >>
rect 91 169 92 170 
<< m1 >>
rect 127 169 128 170 
<< m1 >>
rect 130 169 131 170 
<< m1 >>
rect 132 169 133 170 
<< m1 >>
rect 136 169 137 170 
<< m2 >>
rect 136 169 137 170 
<< m1 >>
rect 145 169 146 170 
<< m2 >>
rect 145 169 146 170 
<< m1 >>
rect 160 169 161 170 
<< m1 >>
rect 163 169 164 170 
<< m1 >>
rect 165 169 166 170 
<< m1 >>
rect 167 169 168 170 
<< m1 >>
rect 168 169 169 170 
<< m1 >>
rect 169 169 170 170 
<< m1 >>
rect 170 169 171 170 
<< m2 >>
rect 170 169 171 170 
<< m1 >>
rect 171 169 172 170 
<< m1 >>
rect 172 169 173 170 
<< m2 >>
rect 172 169 173 170 
<< m1 >>
rect 173 169 174 170 
<< m1 >>
rect 174 169 175 170 
<< m1 >>
rect 175 169 176 170 
<< m1 >>
rect 176 169 177 170 
<< m2 >>
rect 176 169 177 170 
<< m1 >>
rect 177 169 178 170 
<< m1 >>
rect 178 169 179 170 
<< m1 >>
rect 179 169 180 170 
<< m1 >>
rect 180 169 181 170 
<< m1 >>
rect 181 169 182 170 
<< m1 >>
rect 182 169 183 170 
<< m1 >>
rect 183 169 184 170 
<< m2 >>
rect 183 169 184 170 
<< m1 >>
rect 184 169 185 170 
<< m1 >>
rect 185 169 186 170 
<< m1 >>
rect 186 169 187 170 
<< m1 >>
rect 187 169 188 170 
<< m1 >>
rect 188 169 189 170 
<< m2 >>
rect 188 169 189 170 
<< m1 >>
rect 189 169 190 170 
<< m1 >>
rect 190 169 191 170 
<< m2 >>
rect 190 169 191 170 
<< m1 >>
rect 191 169 192 170 
<< m1 >>
rect 192 169 193 170 
<< m1 >>
rect 193 169 194 170 
<< m1 >>
rect 194 169 195 170 
<< m1 >>
rect 195 169 196 170 
<< m1 >>
rect 196 169 197 170 
<< m1 >>
rect 199 169 200 170 
<< m2 >>
rect 225 169 226 170 
<< m1 >>
rect 226 169 227 170 
<< m1 >>
rect 235 169 236 170 
<< m1 >>
rect 237 169 238 170 
<< m2 >>
rect 238 169 239 170 
<< m1 >>
rect 240 169 241 170 
<< m1 >>
rect 253 169 254 170 
<< m1 >>
rect 255 169 256 170 
<< m1 >>
rect 260 169 261 170 
<< m1 >>
rect 262 169 263 170 
<< m2 >>
rect 271 169 272 170 
<< m1 >>
rect 272 169 273 170 
<< m1 >>
rect 274 169 275 170 
<< m2 >>
rect 275 169 276 170 
<< m1 >>
rect 289 169 290 170 
<< m1 >>
rect 296 169 297 170 
<< m1 >>
rect 298 169 299 170 
<< m1 >>
rect 300 169 301 170 
<< m1 >>
rect 301 169 302 170 
<< m1 >>
rect 302 169 303 170 
<< m1 >>
rect 303 169 304 170 
<< m1 >>
rect 304 169 305 170 
<< m1 >>
rect 307 169 308 170 
<< m2 >>
rect 308 169 309 170 
<< m2 >>
rect 326 169 327 170 
<< m1 >>
rect 327 169 328 170 
<< m1 >>
rect 340 169 341 170 
<< m1 >>
rect 343 169 344 170 
<< m2 >>
rect 343 169 344 170 
<< m1 >>
rect 345 169 346 170 
<< m1 >>
rect 10 170 11 171 
<< m1 >>
rect 19 170 20 171 
<< m1 >>
rect 21 170 22 171 
<< m1 >>
rect 23 170 24 171 
<< m2 >>
rect 27 170 28 171 
<< m1 >>
rect 28 170 29 171 
<< m1 >>
rect 37 170 38 171 
<< m2 >>
rect 38 170 39 171 
<< m1 >>
rect 44 170 45 171 
<< m1 >>
rect 46 170 47 171 
<< m1 >>
rect 49 170 50 171 
<< m1 >>
rect 56 170 57 171 
<< m1 >>
rect 58 170 59 171 
<< m1 >>
rect 60 170 61 171 
<< m2 >>
rect 60 170 61 171 
<< m2c >>
rect 60 170 61 171 
<< m1 >>
rect 60 170 61 171 
<< m2 >>
rect 60 170 61 171 
<< m2 >>
rect 61 170 62 171 
<< m1 >>
rect 62 170 63 171 
<< m1 >>
rect 64 170 65 171 
<< m1 >>
rect 80 170 81 171 
<< m2 >>
rect 80 170 81 171 
<< m2c >>
rect 80 170 81 171 
<< m1 >>
rect 80 170 81 171 
<< m2 >>
rect 80 170 81 171 
<< m2 >>
rect 81 170 82 171 
<< m1 >>
rect 82 170 83 171 
<< m2 >>
rect 82 170 83 171 
<< m2 >>
rect 83 170 84 171 
<< m1 >>
rect 84 170 85 171 
<< m2 >>
rect 84 170 85 171 
<< m1 >>
rect 88 170 89 171 
<< m1 >>
rect 91 170 92 171 
<< m1 >>
rect 127 170 128 171 
<< m1 >>
rect 130 170 131 171 
<< m1 >>
rect 132 170 133 171 
<< m1 >>
rect 136 170 137 171 
<< m2 >>
rect 136 170 137 171 
<< m1 >>
rect 145 170 146 171 
<< m2 >>
rect 145 170 146 171 
<< m1 >>
rect 160 170 161 171 
<< m1 >>
rect 163 170 164 171 
<< m1 >>
rect 165 170 166 171 
<< m1 >>
rect 167 170 168 171 
<< m2 >>
rect 170 170 171 171 
<< m2 >>
rect 172 170 173 171 
<< m2 >>
rect 176 170 177 171 
<< m2 >>
rect 183 170 184 171 
<< m2 >>
rect 188 170 189 171 
<< m2 >>
rect 190 170 191 171 
<< m1 >>
rect 199 170 200 171 
<< m2 >>
rect 225 170 226 171 
<< m1 >>
rect 226 170 227 171 
<< m1 >>
rect 235 170 236 171 
<< m1 >>
rect 237 170 238 171 
<< m2 >>
rect 238 170 239 171 
<< m1 >>
rect 240 170 241 171 
<< m2 >>
rect 240 170 241 171 
<< m2c >>
rect 240 170 241 171 
<< m1 >>
rect 240 170 241 171 
<< m2 >>
rect 240 170 241 171 
<< m1 >>
rect 253 170 254 171 
<< m1 >>
rect 255 170 256 171 
<< m1 >>
rect 260 170 261 171 
<< m1 >>
rect 262 170 263 171 
<< m2 >>
rect 271 170 272 171 
<< m1 >>
rect 272 170 273 171 
<< m1 >>
rect 274 170 275 171 
<< m2 >>
rect 275 170 276 171 
<< m1 >>
rect 289 170 290 171 
<< m1 >>
rect 296 170 297 171 
<< m2 >>
rect 296 170 297 171 
<< m2c >>
rect 296 170 297 171 
<< m1 >>
rect 296 170 297 171 
<< m2 >>
rect 296 170 297 171 
<< m2 >>
rect 297 170 298 171 
<< m1 >>
rect 298 170 299 171 
<< m2 >>
rect 298 170 299 171 
<< m2 >>
rect 299 170 300 171 
<< m1 >>
rect 300 170 301 171 
<< m2 >>
rect 300 170 301 171 
<< m2c >>
rect 300 170 301 171 
<< m1 >>
rect 300 170 301 171 
<< m2 >>
rect 300 170 301 171 
<< m1 >>
rect 304 170 305 171 
<< m1 >>
rect 307 170 308 171 
<< m2 >>
rect 308 170 309 171 
<< m2 >>
rect 326 170 327 171 
<< m1 >>
rect 327 170 328 171 
<< m1 >>
rect 340 170 341 171 
<< m1 >>
rect 343 170 344 171 
<< m2 >>
rect 343 170 344 171 
<< m1 >>
rect 345 170 346 171 
<< m1 >>
rect 10 171 11 172 
<< m1 >>
rect 19 171 20 172 
<< m1 >>
rect 21 171 22 172 
<< m1 >>
rect 23 171 24 172 
<< m2 >>
rect 27 171 28 172 
<< m1 >>
rect 28 171 29 172 
<< m1 >>
rect 37 171 38 172 
<< m2 >>
rect 38 171 39 172 
<< m1 >>
rect 44 171 45 172 
<< m1 >>
rect 46 171 47 172 
<< m1 >>
rect 49 171 50 172 
<< m1 >>
rect 56 171 57 172 
<< m1 >>
rect 58 171 59 172 
<< m2 >>
rect 61 171 62 172 
<< m1 >>
rect 62 171 63 172 
<< m1 >>
rect 64 171 65 172 
<< m1 >>
rect 80 171 81 172 
<< m1 >>
rect 82 171 83 172 
<< m1 >>
rect 84 171 85 172 
<< m1 >>
rect 88 171 89 172 
<< m1 >>
rect 91 171 92 172 
<< m1 >>
rect 127 171 128 172 
<< m1 >>
rect 130 171 131 172 
<< m1 >>
rect 132 171 133 172 
<< m1 >>
rect 136 171 137 172 
<< m2 >>
rect 136 171 137 172 
<< m1 >>
rect 145 171 146 172 
<< m2 >>
rect 145 171 146 172 
<< m1 >>
rect 160 171 161 172 
<< m1 >>
rect 163 171 164 172 
<< m1 >>
rect 165 171 166 172 
<< m1 >>
rect 167 171 168 172 
<< m1 >>
rect 170 171 171 172 
<< m2 >>
rect 170 171 171 172 
<< m2c >>
rect 170 171 171 172 
<< m1 >>
rect 170 171 171 172 
<< m2 >>
rect 170 171 171 172 
<< m1 >>
rect 172 171 173 172 
<< m2 >>
rect 172 171 173 172 
<< m2c >>
rect 172 171 173 172 
<< m1 >>
rect 172 171 173 172 
<< m2 >>
rect 172 171 173 172 
<< m1 >>
rect 176 171 177 172 
<< m2 >>
rect 176 171 177 172 
<< m2c >>
rect 176 171 177 172 
<< m1 >>
rect 176 171 177 172 
<< m2 >>
rect 176 171 177 172 
<< m1 >>
rect 177 171 178 172 
<< m1 >>
rect 178 171 179 172 
<< m1 >>
rect 179 171 180 172 
<< m1 >>
rect 180 171 181 172 
<< m1 >>
rect 181 171 182 172 
<< m1 >>
rect 183 171 184 172 
<< m2 >>
rect 183 171 184 172 
<< m2c >>
rect 183 171 184 172 
<< m1 >>
rect 183 171 184 172 
<< m2 >>
rect 183 171 184 172 
<< m1 >>
rect 188 171 189 172 
<< m2 >>
rect 188 171 189 172 
<< m2c >>
rect 188 171 189 172 
<< m1 >>
rect 188 171 189 172 
<< m2 >>
rect 188 171 189 172 
<< m2 >>
rect 190 171 191 172 
<< m1 >>
rect 199 171 200 172 
<< m2 >>
rect 225 171 226 172 
<< m1 >>
rect 226 171 227 172 
<< m1 >>
rect 235 171 236 172 
<< m1 >>
rect 237 171 238 172 
<< m2 >>
rect 238 171 239 172 
<< m2 >>
rect 240 171 241 172 
<< m1 >>
rect 253 171 254 172 
<< m1 >>
rect 255 171 256 172 
<< m1 >>
rect 260 171 261 172 
<< m1 >>
rect 262 171 263 172 
<< m2 >>
rect 271 171 272 172 
<< m1 >>
rect 272 171 273 172 
<< m1 >>
rect 274 171 275 172 
<< m2 >>
rect 275 171 276 172 
<< m1 >>
rect 289 171 290 172 
<< m1 >>
rect 298 171 299 172 
<< m1 >>
rect 304 171 305 172 
<< m1 >>
rect 307 171 308 172 
<< m2 >>
rect 308 171 309 172 
<< m2 >>
rect 326 171 327 172 
<< m1 >>
rect 327 171 328 172 
<< m1 >>
rect 340 171 341 172 
<< m1 >>
rect 343 171 344 172 
<< m2 >>
rect 343 171 344 172 
<< m1 >>
rect 345 171 346 172 
<< m1 >>
rect 10 172 11 173 
<< m1 >>
rect 19 172 20 173 
<< m1 >>
rect 21 172 22 173 
<< m1 >>
rect 23 172 24 173 
<< m2 >>
rect 27 172 28 173 
<< m1 >>
rect 28 172 29 173 
<< m1 >>
rect 37 172 38 173 
<< m2 >>
rect 38 172 39 173 
<< m1 >>
rect 44 172 45 173 
<< m1 >>
rect 46 172 47 173 
<< m1 >>
rect 49 172 50 173 
<< m1 >>
rect 56 172 57 173 
<< m1 >>
rect 58 172 59 173 
<< m2 >>
rect 61 172 62 173 
<< m1 >>
rect 62 172 63 173 
<< m1 >>
rect 64 172 65 173 
<< m1 >>
rect 80 172 81 173 
<< m1 >>
rect 82 172 83 173 
<< m2 >>
rect 82 172 83 173 
<< m2 >>
rect 83 172 84 173 
<< m1 >>
rect 84 172 85 173 
<< m2 >>
rect 84 172 85 173 
<< m2c >>
rect 84 172 85 173 
<< m1 >>
rect 84 172 85 173 
<< m2 >>
rect 84 172 85 173 
<< m1 >>
rect 88 172 89 173 
<< m1 >>
rect 91 172 92 173 
<< m1 >>
rect 127 172 128 173 
<< m1 >>
rect 130 172 131 173 
<< m1 >>
rect 132 172 133 173 
<< m1 >>
rect 136 172 137 173 
<< m2 >>
rect 136 172 137 173 
<< m1 >>
rect 145 172 146 173 
<< m2 >>
rect 145 172 146 173 
<< m1 >>
rect 160 172 161 173 
<< m1 >>
rect 163 172 164 173 
<< m1 >>
rect 165 172 166 173 
<< m1 >>
rect 167 172 168 173 
<< m1 >>
rect 170 172 171 173 
<< m1 >>
rect 172 172 173 173 
<< m1 >>
rect 181 172 182 173 
<< m1 >>
rect 183 172 184 173 
<< m1 >>
rect 188 172 189 173 
<< m1 >>
rect 190 172 191 173 
<< m2 >>
rect 190 172 191 173 
<< m1 >>
rect 191 172 192 173 
<< m1 >>
rect 192 172 193 173 
<< m1 >>
rect 193 172 194 173 
<< m1 >>
rect 196 172 197 173 
<< m1 >>
rect 197 172 198 173 
<< m2 >>
rect 197 172 198 173 
<< m2c >>
rect 197 172 198 173 
<< m1 >>
rect 197 172 198 173 
<< m2 >>
rect 197 172 198 173 
<< m2 >>
rect 198 172 199 173 
<< m1 >>
rect 199 172 200 173 
<< m2 >>
rect 199 172 200 173 
<< m2 >>
rect 200 172 201 173 
<< m1 >>
rect 201 172 202 173 
<< m2 >>
rect 201 172 202 173 
<< m2c >>
rect 201 172 202 173 
<< m1 >>
rect 201 172 202 173 
<< m2 >>
rect 201 172 202 173 
<< m2 >>
rect 225 172 226 173 
<< m1 >>
rect 226 172 227 173 
<< m1 >>
rect 235 172 236 173 
<< m1 >>
rect 237 172 238 173 
<< m2 >>
rect 238 172 239 173 
<< m2 >>
rect 240 172 241 173 
<< m1 >>
rect 241 172 242 173 
<< m1 >>
rect 242 172 243 173 
<< m1 >>
rect 243 172 244 173 
<< m1 >>
rect 244 172 245 173 
<< m1 >>
rect 245 172 246 173 
<< m1 >>
rect 246 172 247 173 
<< m1 >>
rect 247 172 248 173 
<< m1 >>
rect 253 172 254 173 
<< m1 >>
rect 255 172 256 173 
<< m1 >>
rect 260 172 261 173 
<< m1 >>
rect 262 172 263 173 
<< m2 >>
rect 271 172 272 173 
<< m1 >>
rect 272 172 273 173 
<< m1 >>
rect 274 172 275 173 
<< m2 >>
rect 275 172 276 173 
<< m1 >>
rect 289 172 290 173 
<< m1 >>
rect 298 172 299 173 
<< m1 >>
rect 304 172 305 173 
<< m1 >>
rect 307 172 308 173 
<< m2 >>
rect 308 172 309 173 
<< m2 >>
rect 326 172 327 173 
<< m1 >>
rect 327 172 328 173 
<< m1 >>
rect 340 172 341 173 
<< m1 >>
rect 343 172 344 173 
<< m2 >>
rect 343 172 344 173 
<< m1 >>
rect 345 172 346 173 
<< m1 >>
rect 10 173 11 174 
<< m1 >>
rect 19 173 20 174 
<< m1 >>
rect 21 173 22 174 
<< m1 >>
rect 23 173 24 174 
<< m2 >>
rect 27 173 28 174 
<< m1 >>
rect 28 173 29 174 
<< m1 >>
rect 37 173 38 174 
<< m2 >>
rect 38 173 39 174 
<< m1 >>
rect 44 173 45 174 
<< m1 >>
rect 46 173 47 174 
<< m1 >>
rect 49 173 50 174 
<< m1 >>
rect 56 173 57 174 
<< m1 >>
rect 58 173 59 174 
<< m2 >>
rect 61 173 62 174 
<< m1 >>
rect 62 173 63 174 
<< m1 >>
rect 64 173 65 174 
<< m1 >>
rect 80 173 81 174 
<< m1 >>
rect 82 173 83 174 
<< m2 >>
rect 82 173 83 174 
<< m1 >>
rect 88 173 89 174 
<< m1 >>
rect 91 173 92 174 
<< m1 >>
rect 127 173 128 174 
<< m1 >>
rect 130 173 131 174 
<< m1 >>
rect 132 173 133 174 
<< m1 >>
rect 136 173 137 174 
<< m2 >>
rect 136 173 137 174 
<< m1 >>
rect 145 173 146 174 
<< m2 >>
rect 145 173 146 174 
<< m1 >>
rect 160 173 161 174 
<< m1 >>
rect 163 173 164 174 
<< m1 >>
rect 165 173 166 174 
<< m1 >>
rect 167 173 168 174 
<< m1 >>
rect 170 173 171 174 
<< m1 >>
rect 172 173 173 174 
<< m1 >>
rect 181 173 182 174 
<< m1 >>
rect 183 173 184 174 
<< m1 >>
rect 188 173 189 174 
<< m1 >>
rect 190 173 191 174 
<< m2 >>
rect 190 173 191 174 
<< m1 >>
rect 193 173 194 174 
<< m1 >>
rect 196 173 197 174 
<< m1 >>
rect 199 173 200 174 
<< m1 >>
rect 201 173 202 174 
<< m2 >>
rect 225 173 226 174 
<< m1 >>
rect 226 173 227 174 
<< m1 >>
rect 235 173 236 174 
<< m1 >>
rect 237 173 238 174 
<< m2 >>
rect 238 173 239 174 
<< m2 >>
rect 240 173 241 174 
<< m1 >>
rect 241 173 242 174 
<< m1 >>
rect 247 173 248 174 
<< m1 >>
rect 253 173 254 174 
<< m1 >>
rect 255 173 256 174 
<< m1 >>
rect 260 173 261 174 
<< m1 >>
rect 262 173 263 174 
<< m2 >>
rect 271 173 272 174 
<< m1 >>
rect 272 173 273 174 
<< m1 >>
rect 274 173 275 174 
<< m2 >>
rect 275 173 276 174 
<< m1 >>
rect 289 173 290 174 
<< m1 >>
rect 298 173 299 174 
<< m1 >>
rect 304 173 305 174 
<< m1 >>
rect 307 173 308 174 
<< m2 >>
rect 308 173 309 174 
<< m2 >>
rect 326 173 327 174 
<< m1 >>
rect 327 173 328 174 
<< m1 >>
rect 340 173 341 174 
<< m1 >>
rect 343 173 344 174 
<< m2 >>
rect 343 173 344 174 
<< m1 >>
rect 345 173 346 174 
<< m1 >>
rect 10 174 11 175 
<< pdiffusion >>
rect 12 174 13 175 
<< pdiffusion >>
rect 13 174 14 175 
<< pdiffusion >>
rect 14 174 15 175 
<< pdiffusion >>
rect 15 174 16 175 
<< pdiffusion >>
rect 16 174 17 175 
<< pdiffusion >>
rect 17 174 18 175 
<< m1 >>
rect 19 174 20 175 
<< m1 >>
rect 21 174 22 175 
<< m1 >>
rect 23 174 24 175 
<< m2 >>
rect 27 174 28 175 
<< m1 >>
rect 28 174 29 175 
<< pdiffusion >>
rect 30 174 31 175 
<< pdiffusion >>
rect 31 174 32 175 
<< pdiffusion >>
rect 32 174 33 175 
<< pdiffusion >>
rect 33 174 34 175 
<< pdiffusion >>
rect 34 174 35 175 
<< pdiffusion >>
rect 35 174 36 175 
<< m1 >>
rect 37 174 38 175 
<< m2 >>
rect 38 174 39 175 
<< m1 >>
rect 44 174 45 175 
<< m1 >>
rect 46 174 47 175 
<< pdiffusion >>
rect 48 174 49 175 
<< m1 >>
rect 49 174 50 175 
<< pdiffusion >>
rect 49 174 50 175 
<< pdiffusion >>
rect 50 174 51 175 
<< pdiffusion >>
rect 51 174 52 175 
<< pdiffusion >>
rect 52 174 53 175 
<< pdiffusion >>
rect 53 174 54 175 
<< m1 >>
rect 56 174 57 175 
<< m1 >>
rect 58 174 59 175 
<< m2 >>
rect 61 174 62 175 
<< m1 >>
rect 62 174 63 175 
<< m1 >>
rect 64 174 65 175 
<< pdiffusion >>
rect 66 174 67 175 
<< pdiffusion >>
rect 67 174 68 175 
<< pdiffusion >>
rect 68 174 69 175 
<< pdiffusion >>
rect 69 174 70 175 
<< pdiffusion >>
rect 70 174 71 175 
<< pdiffusion >>
rect 71 174 72 175 
<< m1 >>
rect 80 174 81 175 
<< m1 >>
rect 82 174 83 175 
<< m2 >>
rect 82 174 83 175 
<< pdiffusion >>
rect 84 174 85 175 
<< pdiffusion >>
rect 85 174 86 175 
<< pdiffusion >>
rect 86 174 87 175 
<< pdiffusion >>
rect 87 174 88 175 
<< m1 >>
rect 88 174 89 175 
<< pdiffusion >>
rect 88 174 89 175 
<< pdiffusion >>
rect 89 174 90 175 
<< m1 >>
rect 91 174 92 175 
<< pdiffusion >>
rect 102 174 103 175 
<< pdiffusion >>
rect 103 174 104 175 
<< pdiffusion >>
rect 104 174 105 175 
<< pdiffusion >>
rect 105 174 106 175 
<< pdiffusion >>
rect 106 174 107 175 
<< pdiffusion >>
rect 107 174 108 175 
<< pdiffusion >>
rect 120 174 121 175 
<< pdiffusion >>
rect 121 174 122 175 
<< pdiffusion >>
rect 122 174 123 175 
<< pdiffusion >>
rect 123 174 124 175 
<< pdiffusion >>
rect 124 174 125 175 
<< pdiffusion >>
rect 125 174 126 175 
<< m1 >>
rect 127 174 128 175 
<< m1 >>
rect 130 174 131 175 
<< m1 >>
rect 132 174 133 175 
<< m1 >>
rect 136 174 137 175 
<< m2 >>
rect 136 174 137 175 
<< pdiffusion >>
rect 138 174 139 175 
<< pdiffusion >>
rect 139 174 140 175 
<< pdiffusion >>
rect 140 174 141 175 
<< pdiffusion >>
rect 141 174 142 175 
<< pdiffusion >>
rect 142 174 143 175 
<< pdiffusion >>
rect 143 174 144 175 
<< m1 >>
rect 145 174 146 175 
<< m2 >>
rect 145 174 146 175 
<< pdiffusion >>
rect 156 174 157 175 
<< pdiffusion >>
rect 157 174 158 175 
<< pdiffusion >>
rect 158 174 159 175 
<< pdiffusion >>
rect 159 174 160 175 
<< m1 >>
rect 160 174 161 175 
<< pdiffusion >>
rect 160 174 161 175 
<< pdiffusion >>
rect 161 174 162 175 
<< m1 >>
rect 163 174 164 175 
<< m1 >>
rect 165 174 166 175 
<< m1 >>
rect 167 174 168 175 
<< m1 >>
rect 170 174 171 175 
<< m1 >>
rect 172 174 173 175 
<< pdiffusion >>
rect 174 174 175 175 
<< pdiffusion >>
rect 175 174 176 175 
<< pdiffusion >>
rect 176 174 177 175 
<< pdiffusion >>
rect 177 174 178 175 
<< pdiffusion >>
rect 178 174 179 175 
<< pdiffusion >>
rect 179 174 180 175 
<< m1 >>
rect 181 174 182 175 
<< m1 >>
rect 183 174 184 175 
<< m1 >>
rect 188 174 189 175 
<< m1 >>
rect 190 174 191 175 
<< m2 >>
rect 190 174 191 175 
<< pdiffusion >>
rect 192 174 193 175 
<< m1 >>
rect 193 174 194 175 
<< pdiffusion >>
rect 193 174 194 175 
<< pdiffusion >>
rect 194 174 195 175 
<< pdiffusion >>
rect 195 174 196 175 
<< m1 >>
rect 196 174 197 175 
<< pdiffusion >>
rect 196 174 197 175 
<< pdiffusion >>
rect 197 174 198 175 
<< m1 >>
rect 199 174 200 175 
<< m1 >>
rect 201 174 202 175 
<< pdiffusion >>
rect 210 174 211 175 
<< pdiffusion >>
rect 211 174 212 175 
<< pdiffusion >>
rect 212 174 213 175 
<< pdiffusion >>
rect 213 174 214 175 
<< pdiffusion >>
rect 214 174 215 175 
<< pdiffusion >>
rect 215 174 216 175 
<< m2 >>
rect 225 174 226 175 
<< m1 >>
rect 226 174 227 175 
<< pdiffusion >>
rect 228 174 229 175 
<< pdiffusion >>
rect 229 174 230 175 
<< pdiffusion >>
rect 230 174 231 175 
<< pdiffusion >>
rect 231 174 232 175 
<< pdiffusion >>
rect 232 174 233 175 
<< pdiffusion >>
rect 233 174 234 175 
<< m1 >>
rect 235 174 236 175 
<< m1 >>
rect 237 174 238 175 
<< m2 >>
rect 238 174 239 175 
<< m2 >>
rect 240 174 241 175 
<< m1 >>
rect 241 174 242 175 
<< m2 >>
rect 241 174 242 175 
<< m2 >>
rect 242 174 243 175 
<< m1 >>
rect 243 174 244 175 
<< m2 >>
rect 243 174 244 175 
<< m2c >>
rect 243 174 244 175 
<< m1 >>
rect 243 174 244 175 
<< m2 >>
rect 243 174 244 175 
<< pdiffusion >>
rect 246 174 247 175 
<< m1 >>
rect 247 174 248 175 
<< pdiffusion >>
rect 247 174 248 175 
<< pdiffusion >>
rect 248 174 249 175 
<< pdiffusion >>
rect 249 174 250 175 
<< pdiffusion >>
rect 250 174 251 175 
<< pdiffusion >>
rect 251 174 252 175 
<< m1 >>
rect 253 174 254 175 
<< m1 >>
rect 255 174 256 175 
<< m1 >>
rect 260 174 261 175 
<< m1 >>
rect 262 174 263 175 
<< pdiffusion >>
rect 264 174 265 175 
<< pdiffusion >>
rect 265 174 266 175 
<< pdiffusion >>
rect 266 174 267 175 
<< pdiffusion >>
rect 267 174 268 175 
<< pdiffusion >>
rect 268 174 269 175 
<< pdiffusion >>
rect 269 174 270 175 
<< m2 >>
rect 271 174 272 175 
<< m1 >>
rect 272 174 273 175 
<< m1 >>
rect 274 174 275 175 
<< m2 >>
rect 275 174 276 175 
<< pdiffusion >>
rect 282 174 283 175 
<< pdiffusion >>
rect 283 174 284 175 
<< pdiffusion >>
rect 284 174 285 175 
<< pdiffusion >>
rect 285 174 286 175 
<< pdiffusion >>
rect 286 174 287 175 
<< pdiffusion >>
rect 287 174 288 175 
<< m1 >>
rect 289 174 290 175 
<< m1 >>
rect 298 174 299 175 
<< pdiffusion >>
rect 300 174 301 175 
<< pdiffusion >>
rect 301 174 302 175 
<< pdiffusion >>
rect 302 174 303 175 
<< pdiffusion >>
rect 303 174 304 175 
<< m1 >>
rect 304 174 305 175 
<< pdiffusion >>
rect 304 174 305 175 
<< pdiffusion >>
rect 305 174 306 175 
<< m1 >>
rect 307 174 308 175 
<< m2 >>
rect 308 174 309 175 
<< pdiffusion >>
rect 318 174 319 175 
<< pdiffusion >>
rect 319 174 320 175 
<< pdiffusion >>
rect 320 174 321 175 
<< pdiffusion >>
rect 321 174 322 175 
<< pdiffusion >>
rect 322 174 323 175 
<< pdiffusion >>
rect 323 174 324 175 
<< m2 >>
rect 326 174 327 175 
<< m1 >>
rect 327 174 328 175 
<< pdiffusion >>
rect 336 174 337 175 
<< pdiffusion >>
rect 337 174 338 175 
<< pdiffusion >>
rect 338 174 339 175 
<< pdiffusion >>
rect 339 174 340 175 
<< m1 >>
rect 340 174 341 175 
<< pdiffusion >>
rect 340 174 341 175 
<< pdiffusion >>
rect 341 174 342 175 
<< m1 >>
rect 343 174 344 175 
<< m2 >>
rect 343 174 344 175 
<< m1 >>
rect 345 174 346 175 
<< m1 >>
rect 10 175 11 176 
<< pdiffusion >>
rect 12 175 13 176 
<< pdiffusion >>
rect 13 175 14 176 
<< pdiffusion >>
rect 14 175 15 176 
<< pdiffusion >>
rect 15 175 16 176 
<< pdiffusion >>
rect 16 175 17 176 
<< pdiffusion >>
rect 17 175 18 176 
<< m1 >>
rect 19 175 20 176 
<< m1 >>
rect 21 175 22 176 
<< m1 >>
rect 23 175 24 176 
<< m2 >>
rect 27 175 28 176 
<< m1 >>
rect 28 175 29 176 
<< pdiffusion >>
rect 30 175 31 176 
<< pdiffusion >>
rect 31 175 32 176 
<< pdiffusion >>
rect 32 175 33 176 
<< pdiffusion >>
rect 33 175 34 176 
<< pdiffusion >>
rect 34 175 35 176 
<< pdiffusion >>
rect 35 175 36 176 
<< m1 >>
rect 37 175 38 176 
<< m2 >>
rect 38 175 39 176 
<< m1 >>
rect 44 175 45 176 
<< m1 >>
rect 46 175 47 176 
<< pdiffusion >>
rect 48 175 49 176 
<< pdiffusion >>
rect 49 175 50 176 
<< pdiffusion >>
rect 50 175 51 176 
<< pdiffusion >>
rect 51 175 52 176 
<< pdiffusion >>
rect 52 175 53 176 
<< pdiffusion >>
rect 53 175 54 176 
<< m1 >>
rect 56 175 57 176 
<< m1 >>
rect 58 175 59 176 
<< m2 >>
rect 61 175 62 176 
<< m1 >>
rect 62 175 63 176 
<< m1 >>
rect 64 175 65 176 
<< pdiffusion >>
rect 66 175 67 176 
<< pdiffusion >>
rect 67 175 68 176 
<< pdiffusion >>
rect 68 175 69 176 
<< pdiffusion >>
rect 69 175 70 176 
<< pdiffusion >>
rect 70 175 71 176 
<< pdiffusion >>
rect 71 175 72 176 
<< m1 >>
rect 80 175 81 176 
<< m1 >>
rect 82 175 83 176 
<< m2 >>
rect 82 175 83 176 
<< pdiffusion >>
rect 84 175 85 176 
<< pdiffusion >>
rect 85 175 86 176 
<< pdiffusion >>
rect 86 175 87 176 
<< pdiffusion >>
rect 87 175 88 176 
<< pdiffusion >>
rect 88 175 89 176 
<< pdiffusion >>
rect 89 175 90 176 
<< m1 >>
rect 91 175 92 176 
<< pdiffusion >>
rect 102 175 103 176 
<< pdiffusion >>
rect 103 175 104 176 
<< pdiffusion >>
rect 104 175 105 176 
<< pdiffusion >>
rect 105 175 106 176 
<< pdiffusion >>
rect 106 175 107 176 
<< pdiffusion >>
rect 107 175 108 176 
<< pdiffusion >>
rect 120 175 121 176 
<< pdiffusion >>
rect 121 175 122 176 
<< pdiffusion >>
rect 122 175 123 176 
<< pdiffusion >>
rect 123 175 124 176 
<< pdiffusion >>
rect 124 175 125 176 
<< pdiffusion >>
rect 125 175 126 176 
<< m1 >>
rect 127 175 128 176 
<< m1 >>
rect 130 175 131 176 
<< m1 >>
rect 132 175 133 176 
<< m1 >>
rect 136 175 137 176 
<< m2 >>
rect 136 175 137 176 
<< pdiffusion >>
rect 138 175 139 176 
<< pdiffusion >>
rect 139 175 140 176 
<< pdiffusion >>
rect 140 175 141 176 
<< pdiffusion >>
rect 141 175 142 176 
<< pdiffusion >>
rect 142 175 143 176 
<< pdiffusion >>
rect 143 175 144 176 
<< m1 >>
rect 145 175 146 176 
<< m2 >>
rect 145 175 146 176 
<< pdiffusion >>
rect 156 175 157 176 
<< pdiffusion >>
rect 157 175 158 176 
<< pdiffusion >>
rect 158 175 159 176 
<< pdiffusion >>
rect 159 175 160 176 
<< pdiffusion >>
rect 160 175 161 176 
<< pdiffusion >>
rect 161 175 162 176 
<< m1 >>
rect 163 175 164 176 
<< m1 >>
rect 165 175 166 176 
<< m1 >>
rect 167 175 168 176 
<< m1 >>
rect 170 175 171 176 
<< m1 >>
rect 172 175 173 176 
<< pdiffusion >>
rect 174 175 175 176 
<< pdiffusion >>
rect 175 175 176 176 
<< pdiffusion >>
rect 176 175 177 176 
<< pdiffusion >>
rect 177 175 178 176 
<< pdiffusion >>
rect 178 175 179 176 
<< pdiffusion >>
rect 179 175 180 176 
<< m1 >>
rect 181 175 182 176 
<< m1 >>
rect 183 175 184 176 
<< m1 >>
rect 188 175 189 176 
<< m1 >>
rect 190 175 191 176 
<< m2 >>
rect 190 175 191 176 
<< pdiffusion >>
rect 192 175 193 176 
<< pdiffusion >>
rect 193 175 194 176 
<< pdiffusion >>
rect 194 175 195 176 
<< pdiffusion >>
rect 195 175 196 176 
<< pdiffusion >>
rect 196 175 197 176 
<< pdiffusion >>
rect 197 175 198 176 
<< m1 >>
rect 199 175 200 176 
<< m1 >>
rect 201 175 202 176 
<< pdiffusion >>
rect 210 175 211 176 
<< pdiffusion >>
rect 211 175 212 176 
<< pdiffusion >>
rect 212 175 213 176 
<< pdiffusion >>
rect 213 175 214 176 
<< pdiffusion >>
rect 214 175 215 176 
<< pdiffusion >>
rect 215 175 216 176 
<< m2 >>
rect 225 175 226 176 
<< m1 >>
rect 226 175 227 176 
<< pdiffusion >>
rect 228 175 229 176 
<< pdiffusion >>
rect 229 175 230 176 
<< pdiffusion >>
rect 230 175 231 176 
<< pdiffusion >>
rect 231 175 232 176 
<< pdiffusion >>
rect 232 175 233 176 
<< pdiffusion >>
rect 233 175 234 176 
<< m1 >>
rect 235 175 236 176 
<< m1 >>
rect 237 175 238 176 
<< m2 >>
rect 238 175 239 176 
<< m1 >>
rect 241 175 242 176 
<< m1 >>
rect 243 175 244 176 
<< pdiffusion >>
rect 246 175 247 176 
<< pdiffusion >>
rect 247 175 248 176 
<< pdiffusion >>
rect 248 175 249 176 
<< pdiffusion >>
rect 249 175 250 176 
<< pdiffusion >>
rect 250 175 251 176 
<< pdiffusion >>
rect 251 175 252 176 
<< m1 >>
rect 253 175 254 176 
<< m1 >>
rect 255 175 256 176 
<< m1 >>
rect 260 175 261 176 
<< m1 >>
rect 262 175 263 176 
<< pdiffusion >>
rect 264 175 265 176 
<< pdiffusion >>
rect 265 175 266 176 
<< pdiffusion >>
rect 266 175 267 176 
<< pdiffusion >>
rect 267 175 268 176 
<< pdiffusion >>
rect 268 175 269 176 
<< pdiffusion >>
rect 269 175 270 176 
<< m2 >>
rect 271 175 272 176 
<< m1 >>
rect 272 175 273 176 
<< m1 >>
rect 274 175 275 176 
<< m2 >>
rect 275 175 276 176 
<< pdiffusion >>
rect 282 175 283 176 
<< pdiffusion >>
rect 283 175 284 176 
<< pdiffusion >>
rect 284 175 285 176 
<< pdiffusion >>
rect 285 175 286 176 
<< pdiffusion >>
rect 286 175 287 176 
<< pdiffusion >>
rect 287 175 288 176 
<< m1 >>
rect 289 175 290 176 
<< m1 >>
rect 298 175 299 176 
<< pdiffusion >>
rect 300 175 301 176 
<< pdiffusion >>
rect 301 175 302 176 
<< pdiffusion >>
rect 302 175 303 176 
<< pdiffusion >>
rect 303 175 304 176 
<< pdiffusion >>
rect 304 175 305 176 
<< pdiffusion >>
rect 305 175 306 176 
<< m1 >>
rect 307 175 308 176 
<< m2 >>
rect 308 175 309 176 
<< pdiffusion >>
rect 318 175 319 176 
<< pdiffusion >>
rect 319 175 320 176 
<< pdiffusion >>
rect 320 175 321 176 
<< pdiffusion >>
rect 321 175 322 176 
<< pdiffusion >>
rect 322 175 323 176 
<< pdiffusion >>
rect 323 175 324 176 
<< m2 >>
rect 326 175 327 176 
<< m1 >>
rect 327 175 328 176 
<< pdiffusion >>
rect 336 175 337 176 
<< pdiffusion >>
rect 337 175 338 176 
<< pdiffusion >>
rect 338 175 339 176 
<< pdiffusion >>
rect 339 175 340 176 
<< pdiffusion >>
rect 340 175 341 176 
<< pdiffusion >>
rect 341 175 342 176 
<< m1 >>
rect 343 175 344 176 
<< m2 >>
rect 343 175 344 176 
<< m1 >>
rect 345 175 346 176 
<< m1 >>
rect 10 176 11 177 
<< pdiffusion >>
rect 12 176 13 177 
<< pdiffusion >>
rect 13 176 14 177 
<< pdiffusion >>
rect 14 176 15 177 
<< pdiffusion >>
rect 15 176 16 177 
<< pdiffusion >>
rect 16 176 17 177 
<< pdiffusion >>
rect 17 176 18 177 
<< m1 >>
rect 19 176 20 177 
<< m1 >>
rect 21 176 22 177 
<< m1 >>
rect 23 176 24 177 
<< m2 >>
rect 27 176 28 177 
<< m1 >>
rect 28 176 29 177 
<< pdiffusion >>
rect 30 176 31 177 
<< pdiffusion >>
rect 31 176 32 177 
<< pdiffusion >>
rect 32 176 33 177 
<< pdiffusion >>
rect 33 176 34 177 
<< pdiffusion >>
rect 34 176 35 177 
<< pdiffusion >>
rect 35 176 36 177 
<< m1 >>
rect 37 176 38 177 
<< m2 >>
rect 38 176 39 177 
<< m1 >>
rect 44 176 45 177 
<< m1 >>
rect 46 176 47 177 
<< pdiffusion >>
rect 48 176 49 177 
<< pdiffusion >>
rect 49 176 50 177 
<< pdiffusion >>
rect 50 176 51 177 
<< pdiffusion >>
rect 51 176 52 177 
<< pdiffusion >>
rect 52 176 53 177 
<< pdiffusion >>
rect 53 176 54 177 
<< m1 >>
rect 56 176 57 177 
<< m1 >>
rect 58 176 59 177 
<< m2 >>
rect 61 176 62 177 
<< m1 >>
rect 62 176 63 177 
<< m1 >>
rect 64 176 65 177 
<< pdiffusion >>
rect 66 176 67 177 
<< pdiffusion >>
rect 67 176 68 177 
<< pdiffusion >>
rect 68 176 69 177 
<< pdiffusion >>
rect 69 176 70 177 
<< pdiffusion >>
rect 70 176 71 177 
<< pdiffusion >>
rect 71 176 72 177 
<< m1 >>
rect 80 176 81 177 
<< m1 >>
rect 82 176 83 177 
<< m2 >>
rect 82 176 83 177 
<< pdiffusion >>
rect 84 176 85 177 
<< pdiffusion >>
rect 85 176 86 177 
<< pdiffusion >>
rect 86 176 87 177 
<< pdiffusion >>
rect 87 176 88 177 
<< pdiffusion >>
rect 88 176 89 177 
<< pdiffusion >>
rect 89 176 90 177 
<< m1 >>
rect 91 176 92 177 
<< pdiffusion >>
rect 102 176 103 177 
<< pdiffusion >>
rect 103 176 104 177 
<< pdiffusion >>
rect 104 176 105 177 
<< pdiffusion >>
rect 105 176 106 177 
<< pdiffusion >>
rect 106 176 107 177 
<< pdiffusion >>
rect 107 176 108 177 
<< pdiffusion >>
rect 120 176 121 177 
<< pdiffusion >>
rect 121 176 122 177 
<< pdiffusion >>
rect 122 176 123 177 
<< pdiffusion >>
rect 123 176 124 177 
<< pdiffusion >>
rect 124 176 125 177 
<< pdiffusion >>
rect 125 176 126 177 
<< m1 >>
rect 127 176 128 177 
<< m1 >>
rect 130 176 131 177 
<< m1 >>
rect 132 176 133 177 
<< m1 >>
rect 136 176 137 177 
<< m2 >>
rect 136 176 137 177 
<< pdiffusion >>
rect 138 176 139 177 
<< pdiffusion >>
rect 139 176 140 177 
<< pdiffusion >>
rect 140 176 141 177 
<< pdiffusion >>
rect 141 176 142 177 
<< pdiffusion >>
rect 142 176 143 177 
<< pdiffusion >>
rect 143 176 144 177 
<< m1 >>
rect 145 176 146 177 
<< m2 >>
rect 145 176 146 177 
<< pdiffusion >>
rect 156 176 157 177 
<< pdiffusion >>
rect 157 176 158 177 
<< pdiffusion >>
rect 158 176 159 177 
<< pdiffusion >>
rect 159 176 160 177 
<< pdiffusion >>
rect 160 176 161 177 
<< pdiffusion >>
rect 161 176 162 177 
<< m1 >>
rect 163 176 164 177 
<< m1 >>
rect 165 176 166 177 
<< m1 >>
rect 167 176 168 177 
<< m1 >>
rect 170 176 171 177 
<< m1 >>
rect 172 176 173 177 
<< pdiffusion >>
rect 174 176 175 177 
<< pdiffusion >>
rect 175 176 176 177 
<< pdiffusion >>
rect 176 176 177 177 
<< pdiffusion >>
rect 177 176 178 177 
<< pdiffusion >>
rect 178 176 179 177 
<< pdiffusion >>
rect 179 176 180 177 
<< m1 >>
rect 181 176 182 177 
<< m1 >>
rect 183 176 184 177 
<< m1 >>
rect 188 176 189 177 
<< m1 >>
rect 190 176 191 177 
<< m2 >>
rect 190 176 191 177 
<< pdiffusion >>
rect 192 176 193 177 
<< pdiffusion >>
rect 193 176 194 177 
<< pdiffusion >>
rect 194 176 195 177 
<< pdiffusion >>
rect 195 176 196 177 
<< pdiffusion >>
rect 196 176 197 177 
<< pdiffusion >>
rect 197 176 198 177 
<< m1 >>
rect 199 176 200 177 
<< m1 >>
rect 201 176 202 177 
<< pdiffusion >>
rect 210 176 211 177 
<< pdiffusion >>
rect 211 176 212 177 
<< pdiffusion >>
rect 212 176 213 177 
<< pdiffusion >>
rect 213 176 214 177 
<< pdiffusion >>
rect 214 176 215 177 
<< pdiffusion >>
rect 215 176 216 177 
<< m2 >>
rect 225 176 226 177 
<< m1 >>
rect 226 176 227 177 
<< pdiffusion >>
rect 228 176 229 177 
<< pdiffusion >>
rect 229 176 230 177 
<< pdiffusion >>
rect 230 176 231 177 
<< pdiffusion >>
rect 231 176 232 177 
<< pdiffusion >>
rect 232 176 233 177 
<< pdiffusion >>
rect 233 176 234 177 
<< m1 >>
rect 235 176 236 177 
<< m1 >>
rect 237 176 238 177 
<< m2 >>
rect 238 176 239 177 
<< m1 >>
rect 241 176 242 177 
<< m1 >>
rect 243 176 244 177 
<< pdiffusion >>
rect 246 176 247 177 
<< pdiffusion >>
rect 247 176 248 177 
<< pdiffusion >>
rect 248 176 249 177 
<< pdiffusion >>
rect 249 176 250 177 
<< pdiffusion >>
rect 250 176 251 177 
<< pdiffusion >>
rect 251 176 252 177 
<< m1 >>
rect 253 176 254 177 
<< m1 >>
rect 255 176 256 177 
<< m1 >>
rect 260 176 261 177 
<< m1 >>
rect 262 176 263 177 
<< pdiffusion >>
rect 264 176 265 177 
<< pdiffusion >>
rect 265 176 266 177 
<< pdiffusion >>
rect 266 176 267 177 
<< pdiffusion >>
rect 267 176 268 177 
<< pdiffusion >>
rect 268 176 269 177 
<< pdiffusion >>
rect 269 176 270 177 
<< m2 >>
rect 271 176 272 177 
<< m1 >>
rect 272 176 273 177 
<< m1 >>
rect 274 176 275 177 
<< m2 >>
rect 275 176 276 177 
<< pdiffusion >>
rect 282 176 283 177 
<< pdiffusion >>
rect 283 176 284 177 
<< pdiffusion >>
rect 284 176 285 177 
<< pdiffusion >>
rect 285 176 286 177 
<< pdiffusion >>
rect 286 176 287 177 
<< pdiffusion >>
rect 287 176 288 177 
<< m1 >>
rect 289 176 290 177 
<< m1 >>
rect 298 176 299 177 
<< pdiffusion >>
rect 300 176 301 177 
<< pdiffusion >>
rect 301 176 302 177 
<< pdiffusion >>
rect 302 176 303 177 
<< pdiffusion >>
rect 303 176 304 177 
<< pdiffusion >>
rect 304 176 305 177 
<< pdiffusion >>
rect 305 176 306 177 
<< m1 >>
rect 307 176 308 177 
<< m2 >>
rect 308 176 309 177 
<< pdiffusion >>
rect 318 176 319 177 
<< pdiffusion >>
rect 319 176 320 177 
<< pdiffusion >>
rect 320 176 321 177 
<< pdiffusion >>
rect 321 176 322 177 
<< pdiffusion >>
rect 322 176 323 177 
<< pdiffusion >>
rect 323 176 324 177 
<< m2 >>
rect 326 176 327 177 
<< m1 >>
rect 327 176 328 177 
<< pdiffusion >>
rect 336 176 337 177 
<< pdiffusion >>
rect 337 176 338 177 
<< pdiffusion >>
rect 338 176 339 177 
<< pdiffusion >>
rect 339 176 340 177 
<< pdiffusion >>
rect 340 176 341 177 
<< pdiffusion >>
rect 341 176 342 177 
<< m1 >>
rect 343 176 344 177 
<< m2 >>
rect 343 176 344 177 
<< m1 >>
rect 345 176 346 177 
<< m1 >>
rect 10 177 11 178 
<< pdiffusion >>
rect 12 177 13 178 
<< pdiffusion >>
rect 13 177 14 178 
<< pdiffusion >>
rect 14 177 15 178 
<< pdiffusion >>
rect 15 177 16 178 
<< pdiffusion >>
rect 16 177 17 178 
<< pdiffusion >>
rect 17 177 18 178 
<< m1 >>
rect 19 177 20 178 
<< m1 >>
rect 21 177 22 178 
<< m1 >>
rect 23 177 24 178 
<< m2 >>
rect 27 177 28 178 
<< m1 >>
rect 28 177 29 178 
<< pdiffusion >>
rect 30 177 31 178 
<< pdiffusion >>
rect 31 177 32 178 
<< pdiffusion >>
rect 32 177 33 178 
<< pdiffusion >>
rect 33 177 34 178 
<< pdiffusion >>
rect 34 177 35 178 
<< pdiffusion >>
rect 35 177 36 178 
<< m1 >>
rect 37 177 38 178 
<< m2 >>
rect 38 177 39 178 
<< m1 >>
rect 44 177 45 178 
<< m1 >>
rect 46 177 47 178 
<< pdiffusion >>
rect 48 177 49 178 
<< pdiffusion >>
rect 49 177 50 178 
<< pdiffusion >>
rect 50 177 51 178 
<< pdiffusion >>
rect 51 177 52 178 
<< pdiffusion >>
rect 52 177 53 178 
<< pdiffusion >>
rect 53 177 54 178 
<< m1 >>
rect 56 177 57 178 
<< m1 >>
rect 58 177 59 178 
<< m2 >>
rect 61 177 62 178 
<< m1 >>
rect 62 177 63 178 
<< m1 >>
rect 64 177 65 178 
<< pdiffusion >>
rect 66 177 67 178 
<< pdiffusion >>
rect 67 177 68 178 
<< pdiffusion >>
rect 68 177 69 178 
<< pdiffusion >>
rect 69 177 70 178 
<< pdiffusion >>
rect 70 177 71 178 
<< pdiffusion >>
rect 71 177 72 178 
<< m1 >>
rect 80 177 81 178 
<< m1 >>
rect 82 177 83 178 
<< m2 >>
rect 82 177 83 178 
<< pdiffusion >>
rect 84 177 85 178 
<< pdiffusion >>
rect 85 177 86 178 
<< pdiffusion >>
rect 86 177 87 178 
<< pdiffusion >>
rect 87 177 88 178 
<< pdiffusion >>
rect 88 177 89 178 
<< pdiffusion >>
rect 89 177 90 178 
<< m1 >>
rect 91 177 92 178 
<< pdiffusion >>
rect 102 177 103 178 
<< pdiffusion >>
rect 103 177 104 178 
<< pdiffusion >>
rect 104 177 105 178 
<< pdiffusion >>
rect 105 177 106 178 
<< pdiffusion >>
rect 106 177 107 178 
<< pdiffusion >>
rect 107 177 108 178 
<< pdiffusion >>
rect 120 177 121 178 
<< pdiffusion >>
rect 121 177 122 178 
<< pdiffusion >>
rect 122 177 123 178 
<< pdiffusion >>
rect 123 177 124 178 
<< pdiffusion >>
rect 124 177 125 178 
<< pdiffusion >>
rect 125 177 126 178 
<< m1 >>
rect 127 177 128 178 
<< m1 >>
rect 130 177 131 178 
<< m1 >>
rect 132 177 133 178 
<< m1 >>
rect 136 177 137 178 
<< m2 >>
rect 136 177 137 178 
<< pdiffusion >>
rect 138 177 139 178 
<< pdiffusion >>
rect 139 177 140 178 
<< pdiffusion >>
rect 140 177 141 178 
<< pdiffusion >>
rect 141 177 142 178 
<< pdiffusion >>
rect 142 177 143 178 
<< pdiffusion >>
rect 143 177 144 178 
<< m1 >>
rect 145 177 146 178 
<< m2 >>
rect 145 177 146 178 
<< pdiffusion >>
rect 156 177 157 178 
<< pdiffusion >>
rect 157 177 158 178 
<< pdiffusion >>
rect 158 177 159 178 
<< pdiffusion >>
rect 159 177 160 178 
<< pdiffusion >>
rect 160 177 161 178 
<< pdiffusion >>
rect 161 177 162 178 
<< m1 >>
rect 163 177 164 178 
<< m1 >>
rect 165 177 166 178 
<< m1 >>
rect 167 177 168 178 
<< m1 >>
rect 170 177 171 178 
<< m1 >>
rect 172 177 173 178 
<< pdiffusion >>
rect 174 177 175 178 
<< pdiffusion >>
rect 175 177 176 178 
<< pdiffusion >>
rect 176 177 177 178 
<< pdiffusion >>
rect 177 177 178 178 
<< pdiffusion >>
rect 178 177 179 178 
<< pdiffusion >>
rect 179 177 180 178 
<< m1 >>
rect 181 177 182 178 
<< m1 >>
rect 183 177 184 178 
<< m1 >>
rect 188 177 189 178 
<< m1 >>
rect 190 177 191 178 
<< m2 >>
rect 190 177 191 178 
<< pdiffusion >>
rect 192 177 193 178 
<< pdiffusion >>
rect 193 177 194 178 
<< pdiffusion >>
rect 194 177 195 178 
<< pdiffusion >>
rect 195 177 196 178 
<< pdiffusion >>
rect 196 177 197 178 
<< pdiffusion >>
rect 197 177 198 178 
<< m1 >>
rect 199 177 200 178 
<< m1 >>
rect 201 177 202 178 
<< pdiffusion >>
rect 210 177 211 178 
<< pdiffusion >>
rect 211 177 212 178 
<< pdiffusion >>
rect 212 177 213 178 
<< pdiffusion >>
rect 213 177 214 178 
<< pdiffusion >>
rect 214 177 215 178 
<< pdiffusion >>
rect 215 177 216 178 
<< m2 >>
rect 225 177 226 178 
<< m1 >>
rect 226 177 227 178 
<< pdiffusion >>
rect 228 177 229 178 
<< pdiffusion >>
rect 229 177 230 178 
<< pdiffusion >>
rect 230 177 231 178 
<< pdiffusion >>
rect 231 177 232 178 
<< pdiffusion >>
rect 232 177 233 178 
<< pdiffusion >>
rect 233 177 234 178 
<< m1 >>
rect 235 177 236 178 
<< m1 >>
rect 237 177 238 178 
<< m2 >>
rect 238 177 239 178 
<< m1 >>
rect 241 177 242 178 
<< m1 >>
rect 243 177 244 178 
<< pdiffusion >>
rect 246 177 247 178 
<< pdiffusion >>
rect 247 177 248 178 
<< pdiffusion >>
rect 248 177 249 178 
<< pdiffusion >>
rect 249 177 250 178 
<< pdiffusion >>
rect 250 177 251 178 
<< pdiffusion >>
rect 251 177 252 178 
<< m1 >>
rect 253 177 254 178 
<< m1 >>
rect 255 177 256 178 
<< m1 >>
rect 260 177 261 178 
<< m1 >>
rect 262 177 263 178 
<< pdiffusion >>
rect 264 177 265 178 
<< pdiffusion >>
rect 265 177 266 178 
<< pdiffusion >>
rect 266 177 267 178 
<< pdiffusion >>
rect 267 177 268 178 
<< pdiffusion >>
rect 268 177 269 178 
<< pdiffusion >>
rect 269 177 270 178 
<< m2 >>
rect 271 177 272 178 
<< m1 >>
rect 272 177 273 178 
<< m1 >>
rect 274 177 275 178 
<< m2 >>
rect 275 177 276 178 
<< pdiffusion >>
rect 282 177 283 178 
<< pdiffusion >>
rect 283 177 284 178 
<< pdiffusion >>
rect 284 177 285 178 
<< pdiffusion >>
rect 285 177 286 178 
<< pdiffusion >>
rect 286 177 287 178 
<< pdiffusion >>
rect 287 177 288 178 
<< m1 >>
rect 289 177 290 178 
<< m1 >>
rect 298 177 299 178 
<< pdiffusion >>
rect 300 177 301 178 
<< pdiffusion >>
rect 301 177 302 178 
<< pdiffusion >>
rect 302 177 303 178 
<< pdiffusion >>
rect 303 177 304 178 
<< pdiffusion >>
rect 304 177 305 178 
<< pdiffusion >>
rect 305 177 306 178 
<< m1 >>
rect 307 177 308 178 
<< m2 >>
rect 308 177 309 178 
<< pdiffusion >>
rect 318 177 319 178 
<< pdiffusion >>
rect 319 177 320 178 
<< pdiffusion >>
rect 320 177 321 178 
<< pdiffusion >>
rect 321 177 322 178 
<< pdiffusion >>
rect 322 177 323 178 
<< pdiffusion >>
rect 323 177 324 178 
<< m2 >>
rect 326 177 327 178 
<< m1 >>
rect 327 177 328 178 
<< pdiffusion >>
rect 336 177 337 178 
<< pdiffusion >>
rect 337 177 338 178 
<< pdiffusion >>
rect 338 177 339 178 
<< pdiffusion >>
rect 339 177 340 178 
<< pdiffusion >>
rect 340 177 341 178 
<< pdiffusion >>
rect 341 177 342 178 
<< m1 >>
rect 343 177 344 178 
<< m2 >>
rect 343 177 344 178 
<< m1 >>
rect 345 177 346 178 
<< m1 >>
rect 10 178 11 179 
<< pdiffusion >>
rect 12 178 13 179 
<< pdiffusion >>
rect 13 178 14 179 
<< pdiffusion >>
rect 14 178 15 179 
<< pdiffusion >>
rect 15 178 16 179 
<< pdiffusion >>
rect 16 178 17 179 
<< pdiffusion >>
rect 17 178 18 179 
<< m1 >>
rect 19 178 20 179 
<< m1 >>
rect 21 178 22 179 
<< m1 >>
rect 23 178 24 179 
<< m2 >>
rect 27 178 28 179 
<< m1 >>
rect 28 178 29 179 
<< pdiffusion >>
rect 30 178 31 179 
<< pdiffusion >>
rect 31 178 32 179 
<< pdiffusion >>
rect 32 178 33 179 
<< pdiffusion >>
rect 33 178 34 179 
<< pdiffusion >>
rect 34 178 35 179 
<< pdiffusion >>
rect 35 178 36 179 
<< m1 >>
rect 37 178 38 179 
<< m2 >>
rect 38 178 39 179 
<< m1 >>
rect 44 178 45 179 
<< m1 >>
rect 46 178 47 179 
<< pdiffusion >>
rect 48 178 49 179 
<< pdiffusion >>
rect 49 178 50 179 
<< pdiffusion >>
rect 50 178 51 179 
<< pdiffusion >>
rect 51 178 52 179 
<< pdiffusion >>
rect 52 178 53 179 
<< pdiffusion >>
rect 53 178 54 179 
<< m1 >>
rect 56 178 57 179 
<< m1 >>
rect 58 178 59 179 
<< m2 >>
rect 61 178 62 179 
<< m1 >>
rect 62 178 63 179 
<< m1 >>
rect 64 178 65 179 
<< pdiffusion >>
rect 66 178 67 179 
<< pdiffusion >>
rect 67 178 68 179 
<< pdiffusion >>
rect 68 178 69 179 
<< pdiffusion >>
rect 69 178 70 179 
<< pdiffusion >>
rect 70 178 71 179 
<< pdiffusion >>
rect 71 178 72 179 
<< m1 >>
rect 80 178 81 179 
<< m1 >>
rect 82 178 83 179 
<< m2 >>
rect 82 178 83 179 
<< pdiffusion >>
rect 84 178 85 179 
<< pdiffusion >>
rect 85 178 86 179 
<< pdiffusion >>
rect 86 178 87 179 
<< pdiffusion >>
rect 87 178 88 179 
<< pdiffusion >>
rect 88 178 89 179 
<< pdiffusion >>
rect 89 178 90 179 
<< m1 >>
rect 91 178 92 179 
<< pdiffusion >>
rect 102 178 103 179 
<< pdiffusion >>
rect 103 178 104 179 
<< pdiffusion >>
rect 104 178 105 179 
<< pdiffusion >>
rect 105 178 106 179 
<< pdiffusion >>
rect 106 178 107 179 
<< pdiffusion >>
rect 107 178 108 179 
<< pdiffusion >>
rect 120 178 121 179 
<< pdiffusion >>
rect 121 178 122 179 
<< pdiffusion >>
rect 122 178 123 179 
<< pdiffusion >>
rect 123 178 124 179 
<< pdiffusion >>
rect 124 178 125 179 
<< pdiffusion >>
rect 125 178 126 179 
<< m1 >>
rect 127 178 128 179 
<< m1 >>
rect 130 178 131 179 
<< m1 >>
rect 132 178 133 179 
<< m1 >>
rect 136 178 137 179 
<< m2 >>
rect 136 178 137 179 
<< pdiffusion >>
rect 138 178 139 179 
<< pdiffusion >>
rect 139 178 140 179 
<< pdiffusion >>
rect 140 178 141 179 
<< pdiffusion >>
rect 141 178 142 179 
<< pdiffusion >>
rect 142 178 143 179 
<< pdiffusion >>
rect 143 178 144 179 
<< m1 >>
rect 145 178 146 179 
<< m2 >>
rect 145 178 146 179 
<< pdiffusion >>
rect 156 178 157 179 
<< pdiffusion >>
rect 157 178 158 179 
<< pdiffusion >>
rect 158 178 159 179 
<< pdiffusion >>
rect 159 178 160 179 
<< pdiffusion >>
rect 160 178 161 179 
<< pdiffusion >>
rect 161 178 162 179 
<< m1 >>
rect 163 178 164 179 
<< m1 >>
rect 165 178 166 179 
<< m1 >>
rect 167 178 168 179 
<< m1 >>
rect 170 178 171 179 
<< m1 >>
rect 172 178 173 179 
<< pdiffusion >>
rect 174 178 175 179 
<< pdiffusion >>
rect 175 178 176 179 
<< pdiffusion >>
rect 176 178 177 179 
<< pdiffusion >>
rect 177 178 178 179 
<< pdiffusion >>
rect 178 178 179 179 
<< pdiffusion >>
rect 179 178 180 179 
<< m1 >>
rect 181 178 182 179 
<< m1 >>
rect 183 178 184 179 
<< m1 >>
rect 188 178 189 179 
<< m1 >>
rect 190 178 191 179 
<< m2 >>
rect 190 178 191 179 
<< pdiffusion >>
rect 192 178 193 179 
<< pdiffusion >>
rect 193 178 194 179 
<< pdiffusion >>
rect 194 178 195 179 
<< pdiffusion >>
rect 195 178 196 179 
<< pdiffusion >>
rect 196 178 197 179 
<< pdiffusion >>
rect 197 178 198 179 
<< m1 >>
rect 199 178 200 179 
<< m1 >>
rect 201 178 202 179 
<< pdiffusion >>
rect 210 178 211 179 
<< pdiffusion >>
rect 211 178 212 179 
<< pdiffusion >>
rect 212 178 213 179 
<< pdiffusion >>
rect 213 178 214 179 
<< pdiffusion >>
rect 214 178 215 179 
<< pdiffusion >>
rect 215 178 216 179 
<< m2 >>
rect 225 178 226 179 
<< m1 >>
rect 226 178 227 179 
<< pdiffusion >>
rect 228 178 229 179 
<< pdiffusion >>
rect 229 178 230 179 
<< pdiffusion >>
rect 230 178 231 179 
<< pdiffusion >>
rect 231 178 232 179 
<< pdiffusion >>
rect 232 178 233 179 
<< pdiffusion >>
rect 233 178 234 179 
<< m1 >>
rect 235 178 236 179 
<< m1 >>
rect 237 178 238 179 
<< m2 >>
rect 238 178 239 179 
<< m1 >>
rect 241 178 242 179 
<< m1 >>
rect 243 178 244 179 
<< pdiffusion >>
rect 246 178 247 179 
<< pdiffusion >>
rect 247 178 248 179 
<< pdiffusion >>
rect 248 178 249 179 
<< pdiffusion >>
rect 249 178 250 179 
<< pdiffusion >>
rect 250 178 251 179 
<< pdiffusion >>
rect 251 178 252 179 
<< m1 >>
rect 253 178 254 179 
<< m1 >>
rect 255 178 256 179 
<< m1 >>
rect 260 178 261 179 
<< m1 >>
rect 262 178 263 179 
<< pdiffusion >>
rect 264 178 265 179 
<< pdiffusion >>
rect 265 178 266 179 
<< pdiffusion >>
rect 266 178 267 179 
<< pdiffusion >>
rect 267 178 268 179 
<< pdiffusion >>
rect 268 178 269 179 
<< pdiffusion >>
rect 269 178 270 179 
<< m2 >>
rect 271 178 272 179 
<< m1 >>
rect 272 178 273 179 
<< m1 >>
rect 274 178 275 179 
<< m2 >>
rect 275 178 276 179 
<< pdiffusion >>
rect 282 178 283 179 
<< pdiffusion >>
rect 283 178 284 179 
<< pdiffusion >>
rect 284 178 285 179 
<< pdiffusion >>
rect 285 178 286 179 
<< pdiffusion >>
rect 286 178 287 179 
<< pdiffusion >>
rect 287 178 288 179 
<< m1 >>
rect 289 178 290 179 
<< m1 >>
rect 298 178 299 179 
<< pdiffusion >>
rect 300 178 301 179 
<< pdiffusion >>
rect 301 178 302 179 
<< pdiffusion >>
rect 302 178 303 179 
<< pdiffusion >>
rect 303 178 304 179 
<< pdiffusion >>
rect 304 178 305 179 
<< pdiffusion >>
rect 305 178 306 179 
<< m1 >>
rect 307 178 308 179 
<< m2 >>
rect 308 178 309 179 
<< pdiffusion >>
rect 318 178 319 179 
<< pdiffusion >>
rect 319 178 320 179 
<< pdiffusion >>
rect 320 178 321 179 
<< pdiffusion >>
rect 321 178 322 179 
<< pdiffusion >>
rect 322 178 323 179 
<< pdiffusion >>
rect 323 178 324 179 
<< m2 >>
rect 326 178 327 179 
<< m1 >>
rect 327 178 328 179 
<< pdiffusion >>
rect 336 178 337 179 
<< pdiffusion >>
rect 337 178 338 179 
<< pdiffusion >>
rect 338 178 339 179 
<< pdiffusion >>
rect 339 178 340 179 
<< pdiffusion >>
rect 340 178 341 179 
<< pdiffusion >>
rect 341 178 342 179 
<< m1 >>
rect 343 178 344 179 
<< m2 >>
rect 343 178 344 179 
<< m1 >>
rect 345 178 346 179 
<< m1 >>
rect 10 179 11 180 
<< pdiffusion >>
rect 12 179 13 180 
<< pdiffusion >>
rect 13 179 14 180 
<< pdiffusion >>
rect 14 179 15 180 
<< pdiffusion >>
rect 15 179 16 180 
<< pdiffusion >>
rect 16 179 17 180 
<< pdiffusion >>
rect 17 179 18 180 
<< m1 >>
rect 19 179 20 180 
<< m1 >>
rect 21 179 22 180 
<< m1 >>
rect 23 179 24 180 
<< m2 >>
rect 27 179 28 180 
<< m1 >>
rect 28 179 29 180 
<< pdiffusion >>
rect 30 179 31 180 
<< pdiffusion >>
rect 31 179 32 180 
<< pdiffusion >>
rect 32 179 33 180 
<< pdiffusion >>
rect 33 179 34 180 
<< pdiffusion >>
rect 34 179 35 180 
<< pdiffusion >>
rect 35 179 36 180 
<< m1 >>
rect 37 179 38 180 
<< m2 >>
rect 38 179 39 180 
<< m1 >>
rect 44 179 45 180 
<< m1 >>
rect 46 179 47 180 
<< pdiffusion >>
rect 48 179 49 180 
<< pdiffusion >>
rect 49 179 50 180 
<< pdiffusion >>
rect 50 179 51 180 
<< pdiffusion >>
rect 51 179 52 180 
<< pdiffusion >>
rect 52 179 53 180 
<< pdiffusion >>
rect 53 179 54 180 
<< m1 >>
rect 56 179 57 180 
<< m1 >>
rect 58 179 59 180 
<< m2 >>
rect 61 179 62 180 
<< m1 >>
rect 62 179 63 180 
<< m1 >>
rect 64 179 65 180 
<< pdiffusion >>
rect 66 179 67 180 
<< pdiffusion >>
rect 67 179 68 180 
<< pdiffusion >>
rect 68 179 69 180 
<< pdiffusion >>
rect 69 179 70 180 
<< pdiffusion >>
rect 70 179 71 180 
<< pdiffusion >>
rect 71 179 72 180 
<< m1 >>
rect 80 179 81 180 
<< m1 >>
rect 82 179 83 180 
<< m2 >>
rect 82 179 83 180 
<< pdiffusion >>
rect 84 179 85 180 
<< pdiffusion >>
rect 85 179 86 180 
<< pdiffusion >>
rect 86 179 87 180 
<< pdiffusion >>
rect 87 179 88 180 
<< pdiffusion >>
rect 88 179 89 180 
<< pdiffusion >>
rect 89 179 90 180 
<< m1 >>
rect 91 179 92 180 
<< pdiffusion >>
rect 102 179 103 180 
<< pdiffusion >>
rect 103 179 104 180 
<< pdiffusion >>
rect 104 179 105 180 
<< pdiffusion >>
rect 105 179 106 180 
<< pdiffusion >>
rect 106 179 107 180 
<< pdiffusion >>
rect 107 179 108 180 
<< pdiffusion >>
rect 120 179 121 180 
<< m1 >>
rect 121 179 122 180 
<< pdiffusion >>
rect 121 179 122 180 
<< pdiffusion >>
rect 122 179 123 180 
<< pdiffusion >>
rect 123 179 124 180 
<< pdiffusion >>
rect 124 179 125 180 
<< pdiffusion >>
rect 125 179 126 180 
<< m1 >>
rect 127 179 128 180 
<< m1 >>
rect 130 179 131 180 
<< m1 >>
rect 132 179 133 180 
<< m1 >>
rect 136 179 137 180 
<< m2 >>
rect 136 179 137 180 
<< pdiffusion >>
rect 138 179 139 180 
<< pdiffusion >>
rect 139 179 140 180 
<< pdiffusion >>
rect 140 179 141 180 
<< pdiffusion >>
rect 141 179 142 180 
<< pdiffusion >>
rect 142 179 143 180 
<< pdiffusion >>
rect 143 179 144 180 
<< m1 >>
rect 145 179 146 180 
<< m2 >>
rect 145 179 146 180 
<< pdiffusion >>
rect 156 179 157 180 
<< pdiffusion >>
rect 157 179 158 180 
<< pdiffusion >>
rect 158 179 159 180 
<< pdiffusion >>
rect 159 179 160 180 
<< pdiffusion >>
rect 160 179 161 180 
<< pdiffusion >>
rect 161 179 162 180 
<< m1 >>
rect 163 179 164 180 
<< m1 >>
rect 165 179 166 180 
<< m1 >>
rect 167 179 168 180 
<< m1 >>
rect 170 179 171 180 
<< m1 >>
rect 172 179 173 180 
<< pdiffusion >>
rect 174 179 175 180 
<< pdiffusion >>
rect 175 179 176 180 
<< pdiffusion >>
rect 176 179 177 180 
<< pdiffusion >>
rect 177 179 178 180 
<< pdiffusion >>
rect 178 179 179 180 
<< pdiffusion >>
rect 179 179 180 180 
<< m1 >>
rect 181 179 182 180 
<< m1 >>
rect 183 179 184 180 
<< m1 >>
rect 188 179 189 180 
<< m1 >>
rect 190 179 191 180 
<< m2 >>
rect 190 179 191 180 
<< pdiffusion >>
rect 192 179 193 180 
<< pdiffusion >>
rect 193 179 194 180 
<< pdiffusion >>
rect 194 179 195 180 
<< pdiffusion >>
rect 195 179 196 180 
<< pdiffusion >>
rect 196 179 197 180 
<< pdiffusion >>
rect 197 179 198 180 
<< m1 >>
rect 199 179 200 180 
<< m1 >>
rect 201 179 202 180 
<< pdiffusion >>
rect 210 179 211 180 
<< pdiffusion >>
rect 211 179 212 180 
<< pdiffusion >>
rect 212 179 213 180 
<< pdiffusion >>
rect 213 179 214 180 
<< pdiffusion >>
rect 214 179 215 180 
<< pdiffusion >>
rect 215 179 216 180 
<< m2 >>
rect 225 179 226 180 
<< m1 >>
rect 226 179 227 180 
<< pdiffusion >>
rect 228 179 229 180 
<< pdiffusion >>
rect 229 179 230 180 
<< pdiffusion >>
rect 230 179 231 180 
<< pdiffusion >>
rect 231 179 232 180 
<< pdiffusion >>
rect 232 179 233 180 
<< pdiffusion >>
rect 233 179 234 180 
<< m1 >>
rect 235 179 236 180 
<< m1 >>
rect 237 179 238 180 
<< m2 >>
rect 238 179 239 180 
<< m1 >>
rect 241 179 242 180 
<< m1 >>
rect 243 179 244 180 
<< pdiffusion >>
rect 246 179 247 180 
<< pdiffusion >>
rect 247 179 248 180 
<< pdiffusion >>
rect 248 179 249 180 
<< pdiffusion >>
rect 249 179 250 180 
<< pdiffusion >>
rect 250 179 251 180 
<< pdiffusion >>
rect 251 179 252 180 
<< m1 >>
rect 253 179 254 180 
<< m1 >>
rect 255 179 256 180 
<< m1 >>
rect 260 179 261 180 
<< m1 >>
rect 262 179 263 180 
<< pdiffusion >>
rect 264 179 265 180 
<< pdiffusion >>
rect 265 179 266 180 
<< pdiffusion >>
rect 266 179 267 180 
<< pdiffusion >>
rect 267 179 268 180 
<< m1 >>
rect 268 179 269 180 
<< pdiffusion >>
rect 268 179 269 180 
<< pdiffusion >>
rect 269 179 270 180 
<< m2 >>
rect 271 179 272 180 
<< m1 >>
rect 272 179 273 180 
<< m1 >>
rect 274 179 275 180 
<< m2 >>
rect 275 179 276 180 
<< pdiffusion >>
rect 282 179 283 180 
<< pdiffusion >>
rect 283 179 284 180 
<< pdiffusion >>
rect 284 179 285 180 
<< pdiffusion >>
rect 285 179 286 180 
<< pdiffusion >>
rect 286 179 287 180 
<< pdiffusion >>
rect 287 179 288 180 
<< m1 >>
rect 289 179 290 180 
<< m1 >>
rect 298 179 299 180 
<< pdiffusion >>
rect 300 179 301 180 
<< m1 >>
rect 301 179 302 180 
<< pdiffusion >>
rect 301 179 302 180 
<< pdiffusion >>
rect 302 179 303 180 
<< pdiffusion >>
rect 303 179 304 180 
<< pdiffusion >>
rect 304 179 305 180 
<< pdiffusion >>
rect 305 179 306 180 
<< m1 >>
rect 307 179 308 180 
<< m2 >>
rect 308 179 309 180 
<< pdiffusion >>
rect 318 179 319 180 
<< pdiffusion >>
rect 319 179 320 180 
<< pdiffusion >>
rect 320 179 321 180 
<< pdiffusion >>
rect 321 179 322 180 
<< pdiffusion >>
rect 322 179 323 180 
<< pdiffusion >>
rect 323 179 324 180 
<< m2 >>
rect 326 179 327 180 
<< m1 >>
rect 327 179 328 180 
<< pdiffusion >>
rect 336 179 337 180 
<< pdiffusion >>
rect 337 179 338 180 
<< pdiffusion >>
rect 338 179 339 180 
<< pdiffusion >>
rect 339 179 340 180 
<< pdiffusion >>
rect 340 179 341 180 
<< pdiffusion >>
rect 341 179 342 180 
<< m1 >>
rect 343 179 344 180 
<< m2 >>
rect 343 179 344 180 
<< m1 >>
rect 345 179 346 180 
<< m1 >>
rect 10 180 11 181 
<< m1 >>
rect 19 180 20 181 
<< m1 >>
rect 21 180 22 181 
<< m1 >>
rect 23 180 24 181 
<< m2 >>
rect 27 180 28 181 
<< m1 >>
rect 28 180 29 181 
<< m1 >>
rect 37 180 38 181 
<< m2 >>
rect 38 180 39 181 
<< m1 >>
rect 44 180 45 181 
<< m1 >>
rect 46 180 47 181 
<< m1 >>
rect 56 180 57 181 
<< m1 >>
rect 58 180 59 181 
<< m2 >>
rect 61 180 62 181 
<< m1 >>
rect 62 180 63 181 
<< m1 >>
rect 64 180 65 181 
<< m1 >>
rect 80 180 81 181 
<< m1 >>
rect 82 180 83 181 
<< m2 >>
rect 82 180 83 181 
<< m1 >>
rect 91 180 92 181 
<< m1 >>
rect 121 180 122 181 
<< m1 >>
rect 127 180 128 181 
<< m2 >>
rect 127 180 128 181 
<< m2c >>
rect 127 180 128 181 
<< m1 >>
rect 127 180 128 181 
<< m2 >>
rect 127 180 128 181 
<< m1 >>
rect 130 180 131 181 
<< m2 >>
rect 130 180 131 181 
<< m2c >>
rect 130 180 131 181 
<< m1 >>
rect 130 180 131 181 
<< m2 >>
rect 130 180 131 181 
<< m1 >>
rect 132 180 133 181 
<< m2 >>
rect 132 180 133 181 
<< m2c >>
rect 132 180 133 181 
<< m1 >>
rect 132 180 133 181 
<< m2 >>
rect 132 180 133 181 
<< m1 >>
rect 136 180 137 181 
<< m2 >>
rect 136 180 137 181 
<< m1 >>
rect 145 180 146 181 
<< m2 >>
rect 145 180 146 181 
<< m1 >>
rect 163 180 164 181 
<< m1 >>
rect 165 180 166 181 
<< m1 >>
rect 167 180 168 181 
<< m1 >>
rect 170 180 171 181 
<< m1 >>
rect 172 180 173 181 
<< m1 >>
rect 181 180 182 181 
<< m1 >>
rect 183 180 184 181 
<< m1 >>
rect 188 180 189 181 
<< m1 >>
rect 190 180 191 181 
<< m2 >>
rect 190 180 191 181 
<< m1 >>
rect 199 180 200 181 
<< m1 >>
rect 201 180 202 181 
<< m2 >>
rect 225 180 226 181 
<< m1 >>
rect 226 180 227 181 
<< m1 >>
rect 235 180 236 181 
<< m1 >>
rect 237 180 238 181 
<< m2 >>
rect 238 180 239 181 
<< m1 >>
rect 241 180 242 181 
<< m1 >>
rect 243 180 244 181 
<< m1 >>
rect 253 180 254 181 
<< m1 >>
rect 255 180 256 181 
<< m1 >>
rect 260 180 261 181 
<< m1 >>
rect 262 180 263 181 
<< m1 >>
rect 268 180 269 181 
<< m2 >>
rect 271 180 272 181 
<< m1 >>
rect 272 180 273 181 
<< m1 >>
rect 274 180 275 181 
<< m2 >>
rect 275 180 276 181 
<< m1 >>
rect 289 180 290 181 
<< m1 >>
rect 298 180 299 181 
<< m1 >>
rect 301 180 302 181 
<< m1 >>
rect 307 180 308 181 
<< m2 >>
rect 308 180 309 181 
<< m2 >>
rect 326 180 327 181 
<< m1 >>
rect 327 180 328 181 
<< m1 >>
rect 343 180 344 181 
<< m2 >>
rect 343 180 344 181 
<< m1 >>
rect 345 180 346 181 
<< m1 >>
rect 10 181 11 182 
<< m1 >>
rect 19 181 20 182 
<< m1 >>
rect 21 181 22 182 
<< m1 >>
rect 23 181 24 182 
<< m2 >>
rect 27 181 28 182 
<< m1 >>
rect 28 181 29 182 
<< m1 >>
rect 37 181 38 182 
<< m2 >>
rect 38 181 39 182 
<< m1 >>
rect 44 181 45 182 
<< m1 >>
rect 46 181 47 182 
<< m1 >>
rect 56 181 57 182 
<< m1 >>
rect 58 181 59 182 
<< m2 >>
rect 61 181 62 182 
<< m1 >>
rect 62 181 63 182 
<< m2 >>
rect 62 181 63 182 
<< m2 >>
rect 63 181 64 182 
<< m1 >>
rect 64 181 65 182 
<< m2 >>
rect 64 181 65 182 
<< m2 >>
rect 65 181 66 182 
<< m1 >>
rect 66 181 67 182 
<< m2 >>
rect 66 181 67 182 
<< m2c >>
rect 66 181 67 182 
<< m1 >>
rect 66 181 67 182 
<< m2 >>
rect 66 181 67 182 
<< m1 >>
rect 80 181 81 182 
<< m1 >>
rect 82 181 83 182 
<< m2 >>
rect 82 181 83 182 
<< m1 >>
rect 91 181 92 182 
<< m1 >>
rect 121 181 122 182 
<< m2 >>
rect 127 181 128 182 
<< m2 >>
rect 130 181 131 182 
<< m2 >>
rect 132 181 133 182 
<< m1 >>
rect 136 181 137 182 
<< m2 >>
rect 136 181 137 182 
<< m1 >>
rect 145 181 146 182 
<< m2 >>
rect 145 181 146 182 
<< m1 >>
rect 163 181 164 182 
<< m1 >>
rect 165 181 166 182 
<< m1 >>
rect 167 181 168 182 
<< m1 >>
rect 170 181 171 182 
<< m1 >>
rect 172 181 173 182 
<< m1 >>
rect 181 181 182 182 
<< m1 >>
rect 183 181 184 182 
<< m1 >>
rect 188 181 189 182 
<< m1 >>
rect 190 181 191 182 
<< m2 >>
rect 190 181 191 182 
<< m1 >>
rect 199 181 200 182 
<< m1 >>
rect 201 181 202 182 
<< m2 >>
rect 225 181 226 182 
<< m1 >>
rect 226 181 227 182 
<< m1 >>
rect 233 181 234 182 
<< m2 >>
rect 233 181 234 182 
<< m2c >>
rect 233 181 234 182 
<< m1 >>
rect 233 181 234 182 
<< m2 >>
rect 233 181 234 182 
<< m2 >>
rect 234 181 235 182 
<< m1 >>
rect 235 181 236 182 
<< m2 >>
rect 235 181 236 182 
<< m2 >>
rect 236 181 237 182 
<< m1 >>
rect 237 181 238 182 
<< m2 >>
rect 237 181 238 182 
<< m2 >>
rect 238 181 239 182 
<< m1 >>
rect 241 181 242 182 
<< m1 >>
rect 243 181 244 182 
<< m1 >>
rect 253 181 254 182 
<< m1 >>
rect 255 181 256 182 
<< m1 >>
rect 260 181 261 182 
<< m1 >>
rect 262 181 263 182 
<< m1 >>
rect 268 181 269 182 
<< m2 >>
rect 271 181 272 182 
<< m1 >>
rect 272 181 273 182 
<< m1 >>
rect 274 181 275 182 
<< m2 >>
rect 275 181 276 182 
<< m1 >>
rect 289 181 290 182 
<< m1 >>
rect 298 181 299 182 
<< m1 >>
rect 299 181 300 182 
<< m1 >>
rect 300 181 301 182 
<< m1 >>
rect 301 181 302 182 
<< m1 >>
rect 307 181 308 182 
<< m2 >>
rect 308 181 309 182 
<< m2 >>
rect 326 181 327 182 
<< m1 >>
rect 327 181 328 182 
<< m1 >>
rect 343 181 344 182 
<< m2 >>
rect 343 181 344 182 
<< m1 >>
rect 345 181 346 182 
<< m1 >>
rect 10 182 11 183 
<< m1 >>
rect 19 182 20 183 
<< m1 >>
rect 21 182 22 183 
<< m1 >>
rect 23 182 24 183 
<< m2 >>
rect 27 182 28 183 
<< m1 >>
rect 28 182 29 183 
<< m1 >>
rect 37 182 38 183 
<< m2 >>
rect 38 182 39 183 
<< m1 >>
rect 44 182 45 183 
<< m1 >>
rect 46 182 47 183 
<< m1 >>
rect 56 182 57 183 
<< m1 >>
rect 58 182 59 183 
<< m1 >>
rect 62 182 63 183 
<< m1 >>
rect 64 182 65 183 
<< m1 >>
rect 66 182 67 183 
<< m1 >>
rect 80 182 81 183 
<< m2 >>
rect 80 182 81 183 
<< m2c >>
rect 80 182 81 183 
<< m1 >>
rect 80 182 81 183 
<< m2 >>
rect 80 182 81 183 
<< m1 >>
rect 82 182 83 183 
<< m2 >>
rect 82 182 83 183 
<< m1 >>
rect 83 182 84 183 
<< m1 >>
rect 84 182 85 183 
<< m2 >>
rect 84 182 85 183 
<< m2c >>
rect 84 182 85 183 
<< m1 >>
rect 84 182 85 183 
<< m2 >>
rect 84 182 85 183 
<< m1 >>
rect 91 182 92 183 
<< m2 >>
rect 91 182 92 183 
<< m2c >>
rect 91 182 92 183 
<< m1 >>
rect 91 182 92 183 
<< m2 >>
rect 91 182 92 183 
<< m1 >>
rect 121 182 122 183 
<< m1 >>
rect 122 182 123 183 
<< m1 >>
rect 123 182 124 183 
<< m1 >>
rect 124 182 125 183 
<< m1 >>
rect 125 182 126 183 
<< m1 >>
rect 126 182 127 183 
<< m1 >>
rect 127 182 128 183 
<< m2 >>
rect 127 182 128 183 
<< m1 >>
rect 128 182 129 183 
<< m1 >>
rect 129 182 130 183 
<< m1 >>
rect 130 182 131 183 
<< m2 >>
rect 130 182 131 183 
<< m1 >>
rect 131 182 132 183 
<< m1 >>
rect 132 182 133 183 
<< m2 >>
rect 132 182 133 183 
<< m1 >>
rect 133 182 134 183 
<< m1 >>
rect 134 182 135 183 
<< m1 >>
rect 135 182 136 183 
<< m1 >>
rect 136 182 137 183 
<< m2 >>
rect 136 182 137 183 
<< m1 >>
rect 141 182 142 183 
<< m2 >>
rect 141 182 142 183 
<< m2c >>
rect 141 182 142 183 
<< m1 >>
rect 141 182 142 183 
<< m2 >>
rect 141 182 142 183 
<< m1 >>
rect 142 182 143 183 
<< m1 >>
rect 143 182 144 183 
<< m2 >>
rect 143 182 144 183 
<< m2c >>
rect 143 182 144 183 
<< m1 >>
rect 143 182 144 183 
<< m2 >>
rect 143 182 144 183 
<< m2 >>
rect 144 182 145 183 
<< m1 >>
rect 145 182 146 183 
<< m2 >>
rect 145 182 146 183 
<< m1 >>
rect 158 182 159 183 
<< m2 >>
rect 158 182 159 183 
<< m2c >>
rect 158 182 159 183 
<< m1 >>
rect 158 182 159 183 
<< m2 >>
rect 158 182 159 183 
<< m1 >>
rect 159 182 160 183 
<< m1 >>
rect 160 182 161 183 
<< m1 >>
rect 161 182 162 183 
<< m2 >>
rect 161 182 162 183 
<< m2c >>
rect 161 182 162 183 
<< m1 >>
rect 161 182 162 183 
<< m2 >>
rect 161 182 162 183 
<< m2 >>
rect 162 182 163 183 
<< m1 >>
rect 163 182 164 183 
<< m2 >>
rect 163 182 164 183 
<< m2 >>
rect 164 182 165 183 
<< m1 >>
rect 165 182 166 183 
<< m2 >>
rect 165 182 166 183 
<< m2 >>
rect 166 182 167 183 
<< m1 >>
rect 167 182 168 183 
<< m2 >>
rect 167 182 168 183 
<< m2c >>
rect 167 182 168 183 
<< m1 >>
rect 167 182 168 183 
<< m2 >>
rect 167 182 168 183 
<< m1 >>
rect 170 182 171 183 
<< m2 >>
rect 170 182 171 183 
<< m2c >>
rect 170 182 171 183 
<< m1 >>
rect 170 182 171 183 
<< m2 >>
rect 170 182 171 183 
<< m1 >>
rect 172 182 173 183 
<< m2 >>
rect 172 182 173 183 
<< m2c >>
rect 172 182 173 183 
<< m1 >>
rect 172 182 173 183 
<< m2 >>
rect 172 182 173 183 
<< m1 >>
rect 181 182 182 183 
<< m2 >>
rect 181 182 182 183 
<< m2c >>
rect 181 182 182 183 
<< m1 >>
rect 181 182 182 183 
<< m2 >>
rect 181 182 182 183 
<< m1 >>
rect 183 182 184 183 
<< m2 >>
rect 183 182 184 183 
<< m2c >>
rect 183 182 184 183 
<< m1 >>
rect 183 182 184 183 
<< m2 >>
rect 183 182 184 183 
<< m1 >>
rect 188 182 189 183 
<< m2 >>
rect 188 182 189 183 
<< m2c >>
rect 188 182 189 183 
<< m1 >>
rect 188 182 189 183 
<< m2 >>
rect 188 182 189 183 
<< m1 >>
rect 190 182 191 183 
<< m2 >>
rect 190 182 191 183 
<< m1 >>
rect 199 182 200 183 
<< m1 >>
rect 201 182 202 183 
<< m2 >>
rect 225 182 226 183 
<< m1 >>
rect 226 182 227 183 
<< m1 >>
rect 232 182 233 183 
<< m1 >>
rect 233 182 234 183 
<< m1 >>
rect 235 182 236 183 
<< m1 >>
rect 237 182 238 183 
<< m1 >>
rect 241 182 242 183 
<< m1 >>
rect 243 182 244 183 
<< m1 >>
rect 253 182 254 183 
<< m1 >>
rect 255 182 256 183 
<< m1 >>
rect 260 182 261 183 
<< m1 >>
rect 262 182 263 183 
<< m1 >>
rect 268 182 269 183 
<< m2 >>
rect 271 182 272 183 
<< m1 >>
rect 272 182 273 183 
<< m1 >>
rect 274 182 275 183 
<< m2 >>
rect 275 182 276 183 
<< m1 >>
rect 289 182 290 183 
<< m1 >>
rect 307 182 308 183 
<< m2 >>
rect 308 182 309 183 
<< m2 >>
rect 326 182 327 183 
<< m1 >>
rect 327 182 328 183 
<< m1 >>
rect 343 182 344 183 
<< m2 >>
rect 343 182 344 183 
<< m1 >>
rect 345 182 346 183 
<< m1 >>
rect 10 183 11 184 
<< m1 >>
rect 19 183 20 184 
<< m1 >>
rect 21 183 22 184 
<< m1 >>
rect 23 183 24 184 
<< m2 >>
rect 27 183 28 184 
<< m1 >>
rect 28 183 29 184 
<< m1 >>
rect 37 183 38 184 
<< m2 >>
rect 38 183 39 184 
<< m1 >>
rect 44 183 45 184 
<< m1 >>
rect 46 183 47 184 
<< m1 >>
rect 56 183 57 184 
<< m1 >>
rect 58 183 59 184 
<< m1 >>
rect 62 183 63 184 
<< m1 >>
rect 64 183 65 184 
<< m1 >>
rect 66 183 67 184 
<< m2 >>
rect 80 183 81 184 
<< m2 >>
rect 82 183 83 184 
<< m2 >>
rect 84 183 85 184 
<< m2 >>
rect 91 183 92 184 
<< m2 >>
rect 127 183 128 184 
<< m2 >>
rect 130 183 131 184 
<< m2 >>
rect 132 183 133 184 
<< m2 >>
rect 136 183 137 184 
<< m2 >>
rect 141 183 142 184 
<< m1 >>
rect 145 183 146 184 
<< m2 >>
rect 158 183 159 184 
<< m1 >>
rect 163 183 164 184 
<< m1 >>
rect 165 183 166 184 
<< m2 >>
rect 170 183 171 184 
<< m2 >>
rect 172 183 173 184 
<< m2 >>
rect 181 183 182 184 
<< m2 >>
rect 183 183 184 184 
<< m2 >>
rect 188 183 189 184 
<< m1 >>
rect 190 183 191 184 
<< m2 >>
rect 190 183 191 184 
<< m1 >>
rect 199 183 200 184 
<< m1 >>
rect 201 183 202 184 
<< m2 >>
rect 225 183 226 184 
<< m1 >>
rect 226 183 227 184 
<< m1 >>
rect 232 183 233 184 
<< m1 >>
rect 235 183 236 184 
<< m1 >>
rect 237 183 238 184 
<< m1 >>
rect 241 183 242 184 
<< m1 >>
rect 243 183 244 184 
<< m1 >>
rect 253 183 254 184 
<< m1 >>
rect 255 183 256 184 
<< m1 >>
rect 260 183 261 184 
<< m1 >>
rect 262 183 263 184 
<< m1 >>
rect 268 183 269 184 
<< m2 >>
rect 271 183 272 184 
<< m1 >>
rect 272 183 273 184 
<< m1 >>
rect 274 183 275 184 
<< m2 >>
rect 275 183 276 184 
<< m1 >>
rect 289 183 290 184 
<< m1 >>
rect 307 183 308 184 
<< m2 >>
rect 308 183 309 184 
<< m2 >>
rect 326 183 327 184 
<< m1 >>
rect 327 183 328 184 
<< m1 >>
rect 343 183 344 184 
<< m2 >>
rect 343 183 344 184 
<< m1 >>
rect 345 183 346 184 
<< m1 >>
rect 10 184 11 185 
<< m1 >>
rect 19 184 20 185 
<< m1 >>
rect 21 184 22 185 
<< m1 >>
rect 23 184 24 185 
<< m2 >>
rect 27 184 28 185 
<< m1 >>
rect 28 184 29 185 
<< m1 >>
rect 37 184 38 185 
<< m2 >>
rect 38 184 39 185 
<< m1 >>
rect 44 184 45 185 
<< m1 >>
rect 46 184 47 185 
<< m1 >>
rect 56 184 57 185 
<< m1 >>
rect 58 184 59 185 
<< m1 >>
rect 62 184 63 185 
<< m1 >>
rect 64 184 65 185 
<< m1 >>
rect 66 184 67 185 
<< m1 >>
rect 67 184 68 185 
<< m1 >>
rect 68 184 69 185 
<< m2 >>
rect 68 184 69 185 
<< m2c >>
rect 68 184 69 185 
<< m1 >>
rect 68 184 69 185 
<< m2 >>
rect 68 184 69 185 
<< m2 >>
rect 69 184 70 185 
<< m1 >>
rect 70 184 71 185 
<< m2 >>
rect 70 184 71 185 
<< m1 >>
rect 71 184 72 185 
<< m2 >>
rect 71 184 72 185 
<< m1 >>
rect 72 184 73 185 
<< m2 >>
rect 72 184 73 185 
<< m1 >>
rect 73 184 74 185 
<< m2 >>
rect 73 184 74 185 
<< m1 >>
rect 74 184 75 185 
<< m2 >>
rect 74 184 75 185 
<< m1 >>
rect 75 184 76 185 
<< m1 >>
rect 76 184 77 185 
<< m1 >>
rect 77 184 78 185 
<< m1 >>
rect 78 184 79 185 
<< m1 >>
rect 79 184 80 185 
<< m1 >>
rect 80 184 81 185 
<< m2 >>
rect 80 184 81 185 
<< m1 >>
rect 81 184 82 185 
<< m1 >>
rect 82 184 83 185 
<< m2 >>
rect 82 184 83 185 
<< m1 >>
rect 83 184 84 185 
<< m1 >>
rect 84 184 85 185 
<< m2 >>
rect 84 184 85 185 
<< m1 >>
rect 85 184 86 185 
<< m1 >>
rect 86 184 87 185 
<< m1 >>
rect 87 184 88 185 
<< m1 >>
rect 88 184 89 185 
<< m1 >>
rect 89 184 90 185 
<< m1 >>
rect 90 184 91 185 
<< m1 >>
rect 91 184 92 185 
<< m2 >>
rect 91 184 92 185 
<< m1 >>
rect 92 184 93 185 
<< m2 >>
rect 92 184 93 185 
<< m1 >>
rect 93 184 94 185 
<< m2 >>
rect 93 184 94 185 
<< m1 >>
rect 94 184 95 185 
<< m2 >>
rect 94 184 95 185 
<< m1 >>
rect 95 184 96 185 
<< m2 >>
rect 95 184 96 185 
<< m1 >>
rect 96 184 97 185 
<< m2 >>
rect 96 184 97 185 
<< m1 >>
rect 97 184 98 185 
<< m2 >>
rect 97 184 98 185 
<< m1 >>
rect 98 184 99 185 
<< m2 >>
rect 98 184 99 185 
<< m1 >>
rect 99 184 100 185 
<< m2 >>
rect 99 184 100 185 
<< m1 >>
rect 100 184 101 185 
<< m2 >>
rect 100 184 101 185 
<< m1 >>
rect 101 184 102 185 
<< m2 >>
rect 101 184 102 185 
<< m1 >>
rect 102 184 103 185 
<< m2 >>
rect 102 184 103 185 
<< m1 >>
rect 103 184 104 185 
<< m2 >>
rect 103 184 104 185 
<< m1 >>
rect 104 184 105 185 
<< m2 >>
rect 104 184 105 185 
<< m1 >>
rect 105 184 106 185 
<< m2 >>
rect 105 184 106 185 
<< m1 >>
rect 106 184 107 185 
<< m2 >>
rect 106 184 107 185 
<< m1 >>
rect 107 184 108 185 
<< m2 >>
rect 107 184 108 185 
<< m1 >>
rect 108 184 109 185 
<< m2 >>
rect 108 184 109 185 
<< m1 >>
rect 109 184 110 185 
<< m2 >>
rect 109 184 110 185 
<< m1 >>
rect 110 184 111 185 
<< m2 >>
rect 110 184 111 185 
<< m1 >>
rect 111 184 112 185 
<< m2 >>
rect 111 184 112 185 
<< m1 >>
rect 112 184 113 185 
<< m2 >>
rect 112 184 113 185 
<< m1 >>
rect 113 184 114 185 
<< m2 >>
rect 113 184 114 185 
<< m1 >>
rect 114 184 115 185 
<< m2 >>
rect 114 184 115 185 
<< m1 >>
rect 115 184 116 185 
<< m2 >>
rect 115 184 116 185 
<< m1 >>
rect 116 184 117 185 
<< m2 >>
rect 116 184 117 185 
<< m1 >>
rect 117 184 118 185 
<< m2 >>
rect 117 184 118 185 
<< m1 >>
rect 118 184 119 185 
<< m2 >>
rect 118 184 119 185 
<< m1 >>
rect 119 184 120 185 
<< m2 >>
rect 119 184 120 185 
<< m1 >>
rect 120 184 121 185 
<< m2 >>
rect 120 184 121 185 
<< m1 >>
rect 121 184 122 185 
<< m2 >>
rect 121 184 122 185 
<< m1 >>
rect 122 184 123 185 
<< m2 >>
rect 122 184 123 185 
<< m1 >>
rect 123 184 124 185 
<< m1 >>
rect 124 184 125 185 
<< m1 >>
rect 125 184 126 185 
<< m1 >>
rect 126 184 127 185 
<< m1 >>
rect 127 184 128 185 
<< m2 >>
rect 127 184 128 185 
<< m1 >>
rect 128 184 129 185 
<< m1 >>
rect 129 184 130 185 
<< m1 >>
rect 130 184 131 185 
<< m2 >>
rect 130 184 131 185 
<< m1 >>
rect 131 184 132 185 
<< m1 >>
rect 132 184 133 185 
<< m2 >>
rect 132 184 133 185 
<< m1 >>
rect 133 184 134 185 
<< m1 >>
rect 134 184 135 185 
<< m1 >>
rect 135 184 136 185 
<< m1 >>
rect 136 184 137 185 
<< m2 >>
rect 136 184 137 185 
<< m1 >>
rect 137 184 138 185 
<< m1 >>
rect 138 184 139 185 
<< m1 >>
rect 139 184 140 185 
<< m1 >>
rect 140 184 141 185 
<< m1 >>
rect 141 184 142 185 
<< m2 >>
rect 141 184 142 185 
<< m1 >>
rect 142 184 143 185 
<< m1 >>
rect 143 184 144 185 
<< m2 >>
rect 143 184 144 185 
<< m2c >>
rect 143 184 144 185 
<< m1 >>
rect 143 184 144 185 
<< m2 >>
rect 143 184 144 185 
<< m2 >>
rect 144 184 145 185 
<< m1 >>
rect 145 184 146 185 
<< m2 >>
rect 145 184 146 185 
<< m2 >>
rect 146 184 147 185 
<< m1 >>
rect 147 184 148 185 
<< m2 >>
rect 147 184 148 185 
<< m2c >>
rect 147 184 148 185 
<< m1 >>
rect 147 184 148 185 
<< m2 >>
rect 147 184 148 185 
<< m1 >>
rect 148 184 149 185 
<< m1 >>
rect 149 184 150 185 
<< m1 >>
rect 150 184 151 185 
<< m1 >>
rect 151 184 152 185 
<< m1 >>
rect 152 184 153 185 
<< m1 >>
rect 153 184 154 185 
<< m1 >>
rect 154 184 155 185 
<< m1 >>
rect 155 184 156 185 
<< m1 >>
rect 156 184 157 185 
<< m1 >>
rect 157 184 158 185 
<< m1 >>
rect 158 184 159 185 
<< m2 >>
rect 158 184 159 185 
<< m1 >>
rect 159 184 160 185 
<< m1 >>
rect 160 184 161 185 
<< m1 >>
rect 161 184 162 185 
<< m2 >>
rect 161 184 162 185 
<< m2c >>
rect 161 184 162 185 
<< m1 >>
rect 161 184 162 185 
<< m2 >>
rect 161 184 162 185 
<< m2 >>
rect 162 184 163 185 
<< m1 >>
rect 163 184 164 185 
<< m2 >>
rect 163 184 164 185 
<< m2 >>
rect 164 184 165 185 
<< m1 >>
rect 165 184 166 185 
<< m2 >>
rect 165 184 166 185 
<< m2 >>
rect 166 184 167 185 
<< m1 >>
rect 167 184 168 185 
<< m2 >>
rect 167 184 168 185 
<< m2c >>
rect 167 184 168 185 
<< m1 >>
rect 167 184 168 185 
<< m2 >>
rect 167 184 168 185 
<< m1 >>
rect 168 184 169 185 
<< m1 >>
rect 169 184 170 185 
<< m1 >>
rect 170 184 171 185 
<< m2 >>
rect 170 184 171 185 
<< m1 >>
rect 171 184 172 185 
<< m1 >>
rect 172 184 173 185 
<< m2 >>
rect 172 184 173 185 
<< m1 >>
rect 173 184 174 185 
<< m1 >>
rect 174 184 175 185 
<< m1 >>
rect 175 184 176 185 
<< m1 >>
rect 176 184 177 185 
<< m1 >>
rect 177 184 178 185 
<< m1 >>
rect 178 184 179 185 
<< m1 >>
rect 179 184 180 185 
<< m1 >>
rect 180 184 181 185 
<< m1 >>
rect 181 184 182 185 
<< m2 >>
rect 181 184 182 185 
<< m1 >>
rect 182 184 183 185 
<< m1 >>
rect 183 184 184 185 
<< m2 >>
rect 183 184 184 185 
<< m1 >>
rect 184 184 185 185 
<< m1 >>
rect 185 184 186 185 
<< m1 >>
rect 186 184 187 185 
<< m1 >>
rect 187 184 188 185 
<< m1 >>
rect 188 184 189 185 
<< m2 >>
rect 188 184 189 185 
<< m1 >>
rect 189 184 190 185 
<< m1 >>
rect 190 184 191 185 
<< m2 >>
rect 190 184 191 185 
<< m1 >>
rect 199 184 200 185 
<< m1 >>
rect 201 184 202 185 
<< m2 >>
rect 225 184 226 185 
<< m1 >>
rect 226 184 227 185 
<< m1 >>
rect 232 184 233 185 
<< m1 >>
rect 235 184 236 185 
<< m1 >>
rect 237 184 238 185 
<< m1 >>
rect 241 184 242 185 
<< m1 >>
rect 243 184 244 185 
<< m1 >>
rect 253 184 254 185 
<< m1 >>
rect 255 184 256 185 
<< m1 >>
rect 260 184 261 185 
<< m1 >>
rect 262 184 263 185 
<< m2 >>
rect 262 184 263 185 
<< m2 >>
rect 263 184 264 185 
<< m1 >>
rect 264 184 265 185 
<< m2 >>
rect 264 184 265 185 
<< m2c >>
rect 264 184 265 185 
<< m1 >>
rect 264 184 265 185 
<< m2 >>
rect 264 184 265 185 
<< m1 >>
rect 265 184 266 185 
<< m1 >>
rect 266 184 267 185 
<< m1 >>
rect 267 184 268 185 
<< m1 >>
rect 268 184 269 185 
<< m2 >>
rect 271 184 272 185 
<< m1 >>
rect 272 184 273 185 
<< m1 >>
rect 274 184 275 185 
<< m2 >>
rect 275 184 276 185 
<< m1 >>
rect 289 184 290 185 
<< m1 >>
rect 307 184 308 185 
<< m2 >>
rect 308 184 309 185 
<< m2 >>
rect 326 184 327 185 
<< m1 >>
rect 327 184 328 185 
<< m1 >>
rect 343 184 344 185 
<< m2 >>
rect 343 184 344 185 
<< m1 >>
rect 345 184 346 185 
<< m1 >>
rect 10 185 11 186 
<< m1 >>
rect 19 185 20 186 
<< m1 >>
rect 21 185 22 186 
<< m1 >>
rect 23 185 24 186 
<< m2 >>
rect 27 185 28 186 
<< m1 >>
rect 28 185 29 186 
<< m1 >>
rect 37 185 38 186 
<< m2 >>
rect 38 185 39 186 
<< m1 >>
rect 44 185 45 186 
<< m1 >>
rect 46 185 47 186 
<< m1 >>
rect 56 185 57 186 
<< m1 >>
rect 58 185 59 186 
<< m1 >>
rect 62 185 63 186 
<< m1 >>
rect 64 185 65 186 
<< m1 >>
rect 70 185 71 186 
<< m2 >>
rect 74 185 75 186 
<< m2 >>
rect 80 185 81 186 
<< m2 >>
rect 82 185 83 186 
<< m2 >>
rect 84 185 85 186 
<< m2 >>
rect 122 185 123 186 
<< m2 >>
rect 127 185 128 186 
<< m2 >>
rect 130 185 131 186 
<< m2 >>
rect 132 185 133 186 
<< m2 >>
rect 136 185 137 186 
<< m2 >>
rect 141 185 142 186 
<< m1 >>
rect 145 185 146 186 
<< m2 >>
rect 149 185 150 186 
<< m2 >>
rect 150 185 151 186 
<< m2 >>
rect 151 185 152 186 
<< m2 >>
rect 152 185 153 186 
<< m2 >>
rect 153 185 154 186 
<< m2 >>
rect 154 185 155 186 
<< m2 >>
rect 155 185 156 186 
<< m2 >>
rect 156 185 157 186 
<< m2 >>
rect 157 185 158 186 
<< m2 >>
rect 158 185 159 186 
<< m1 >>
rect 163 185 164 186 
<< m1 >>
rect 165 185 166 186 
<< m2 >>
rect 170 185 171 186 
<< m2 >>
rect 172 185 173 186 
<< m2 >>
rect 181 185 182 186 
<< m2 >>
rect 183 185 184 186 
<< m2 >>
rect 188 185 189 186 
<< m2 >>
rect 190 185 191 186 
<< m1 >>
rect 199 185 200 186 
<< m1 >>
rect 201 185 202 186 
<< m2 >>
rect 225 185 226 186 
<< m1 >>
rect 226 185 227 186 
<< m1 >>
rect 232 185 233 186 
<< m1 >>
rect 235 185 236 186 
<< m1 >>
rect 237 185 238 186 
<< m1 >>
rect 241 185 242 186 
<< m1 >>
rect 243 185 244 186 
<< m1 >>
rect 253 185 254 186 
<< m1 >>
rect 255 185 256 186 
<< m1 >>
rect 260 185 261 186 
<< m1 >>
rect 262 185 263 186 
<< m2 >>
rect 262 185 263 186 
<< m2 >>
rect 271 185 272 186 
<< m1 >>
rect 272 185 273 186 
<< m1 >>
rect 274 185 275 186 
<< m2 >>
rect 275 185 276 186 
<< m1 >>
rect 289 185 290 186 
<< m1 >>
rect 307 185 308 186 
<< m2 >>
rect 308 185 309 186 
<< m2 >>
rect 326 185 327 186 
<< m1 >>
rect 327 185 328 186 
<< m1 >>
rect 343 185 344 186 
<< m2 >>
rect 343 185 344 186 
<< m1 >>
rect 345 185 346 186 
<< m1 >>
rect 10 186 11 187 
<< m1 >>
rect 19 186 20 187 
<< m1 >>
rect 21 186 22 187 
<< m1 >>
rect 23 186 24 187 
<< m2 >>
rect 27 186 28 187 
<< m1 >>
rect 28 186 29 187 
<< m1 >>
rect 37 186 38 187 
<< m2 >>
rect 38 186 39 187 
<< m1 >>
rect 44 186 45 187 
<< m1 >>
rect 46 186 47 187 
<< m1 >>
rect 56 186 57 187 
<< m1 >>
rect 58 186 59 187 
<< m1 >>
rect 62 186 63 187 
<< m1 >>
rect 64 186 65 187 
<< m1 >>
rect 70 186 71 187 
<< m2 >>
rect 74 186 75 187 
<< m2 >>
rect 80 186 81 187 
<< m2 >>
rect 82 186 83 187 
<< m2 >>
rect 84 186 85 187 
<< m2 >>
rect 122 186 123 187 
<< m2 >>
rect 127 186 128 187 
<< m2 >>
rect 130 186 131 187 
<< m2 >>
rect 132 186 133 187 
<< m2 >>
rect 136 186 137 187 
<< m2 >>
rect 141 186 142 187 
<< m1 >>
rect 145 186 146 187 
<< m1 >>
rect 149 186 150 187 
<< m2 >>
rect 149 186 150 187 
<< m2c >>
rect 149 186 150 187 
<< m1 >>
rect 149 186 150 187 
<< m2 >>
rect 149 186 150 187 
<< m1 >>
rect 163 186 164 187 
<< m1 >>
rect 165 186 166 187 
<< m1 >>
rect 170 186 171 187 
<< m2 >>
rect 170 186 171 187 
<< m2c >>
rect 170 186 171 187 
<< m1 >>
rect 170 186 171 187 
<< m2 >>
rect 170 186 171 187 
<< m1 >>
rect 172 186 173 187 
<< m2 >>
rect 172 186 173 187 
<< m2c >>
rect 172 186 173 187 
<< m1 >>
rect 172 186 173 187 
<< m2 >>
rect 172 186 173 187 
<< m1 >>
rect 181 186 182 187 
<< m2 >>
rect 181 186 182 187 
<< m2c >>
rect 181 186 182 187 
<< m1 >>
rect 181 186 182 187 
<< m2 >>
rect 181 186 182 187 
<< m1 >>
rect 183 186 184 187 
<< m2 >>
rect 183 186 184 187 
<< m2c >>
rect 183 186 184 187 
<< m1 >>
rect 183 186 184 187 
<< m2 >>
rect 183 186 184 187 
<< m1 >>
rect 188 186 189 187 
<< m2 >>
rect 188 186 189 187 
<< m2c >>
rect 188 186 189 187 
<< m1 >>
rect 188 186 189 187 
<< m2 >>
rect 188 186 189 187 
<< m1 >>
rect 190 186 191 187 
<< m2 >>
rect 190 186 191 187 
<< m2c >>
rect 190 186 191 187 
<< m1 >>
rect 190 186 191 187 
<< m2 >>
rect 190 186 191 187 
<< m1 >>
rect 199 186 200 187 
<< m1 >>
rect 201 186 202 187 
<< m2 >>
rect 225 186 226 187 
<< m1 >>
rect 226 186 227 187 
<< m1 >>
rect 232 186 233 187 
<< m1 >>
rect 235 186 236 187 
<< m1 >>
rect 237 186 238 187 
<< m1 >>
rect 241 186 242 187 
<< m1 >>
rect 243 186 244 187 
<< m1 >>
rect 253 186 254 187 
<< m1 >>
rect 255 186 256 187 
<< m1 >>
rect 260 186 261 187 
<< m1 >>
rect 262 186 263 187 
<< m2 >>
rect 262 186 263 187 
<< m2 >>
rect 271 186 272 187 
<< m1 >>
rect 272 186 273 187 
<< m1 >>
rect 274 186 275 187 
<< m2 >>
rect 275 186 276 187 
<< m1 >>
rect 289 186 290 187 
<< m1 >>
rect 307 186 308 187 
<< m2 >>
rect 308 186 309 187 
<< m2 >>
rect 326 186 327 187 
<< m1 >>
rect 327 186 328 187 
<< m1 >>
rect 343 186 344 187 
<< m2 >>
rect 343 186 344 187 
<< m1 >>
rect 345 186 346 187 
<< m1 >>
rect 10 187 11 188 
<< m1 >>
rect 19 187 20 188 
<< m1 >>
rect 21 187 22 188 
<< m1 >>
rect 23 187 24 188 
<< m2 >>
rect 27 187 28 188 
<< m1 >>
rect 28 187 29 188 
<< m1 >>
rect 37 187 38 188 
<< m2 >>
rect 38 187 39 188 
<< m1 >>
rect 44 187 45 188 
<< m1 >>
rect 46 187 47 188 
<< m1 >>
rect 56 187 57 188 
<< m1 >>
rect 58 187 59 188 
<< m1 >>
rect 62 187 63 188 
<< m1 >>
rect 64 187 65 188 
<< m1 >>
rect 70 187 71 188 
<< m1 >>
rect 72 187 73 188 
<< m1 >>
rect 73 187 74 188 
<< m1 >>
rect 74 187 75 188 
<< m2 >>
rect 74 187 75 188 
<< m1 >>
rect 75 187 76 188 
<< m1 >>
rect 76 187 77 188 
<< m1 >>
rect 77 187 78 188 
<< m1 >>
rect 78 187 79 188 
<< m1 >>
rect 79 187 80 188 
<< m1 >>
rect 80 187 81 188 
<< m2 >>
rect 80 187 81 188 
<< m1 >>
rect 81 187 82 188 
<< m1 >>
rect 82 187 83 188 
<< m2 >>
rect 82 187 83 188 
<< m1 >>
rect 83 187 84 188 
<< m1 >>
rect 84 187 85 188 
<< m2 >>
rect 84 187 85 188 
<< m1 >>
rect 85 187 86 188 
<< m2 >>
rect 85 187 86 188 
<< m1 >>
rect 86 187 87 188 
<< m2 >>
rect 86 187 87 188 
<< m1 >>
rect 87 187 88 188 
<< m2 >>
rect 87 187 88 188 
<< m1 >>
rect 88 187 89 188 
<< m2 >>
rect 88 187 89 188 
<< m1 >>
rect 89 187 90 188 
<< m2 >>
rect 89 187 90 188 
<< m1 >>
rect 90 187 91 188 
<< m2 >>
rect 90 187 91 188 
<< m1 >>
rect 91 187 92 188 
<< m2 >>
rect 91 187 92 188 
<< m1 >>
rect 92 187 93 188 
<< m2 >>
rect 92 187 93 188 
<< m1 >>
rect 93 187 94 188 
<< m2 >>
rect 93 187 94 188 
<< m1 >>
rect 94 187 95 188 
<< m2 >>
rect 94 187 95 188 
<< m1 >>
rect 95 187 96 188 
<< m2 >>
rect 95 187 96 188 
<< m1 >>
rect 96 187 97 188 
<< m2 >>
rect 96 187 97 188 
<< m1 >>
rect 97 187 98 188 
<< m2 >>
rect 97 187 98 188 
<< m1 >>
rect 98 187 99 188 
<< m2 >>
rect 98 187 99 188 
<< m1 >>
rect 99 187 100 188 
<< m2 >>
rect 99 187 100 188 
<< m1 >>
rect 100 187 101 188 
<< m2 >>
rect 100 187 101 188 
<< m1 >>
rect 101 187 102 188 
<< m2 >>
rect 101 187 102 188 
<< m1 >>
rect 102 187 103 188 
<< m2 >>
rect 102 187 103 188 
<< m1 >>
rect 103 187 104 188 
<< m2 >>
rect 103 187 104 188 
<< m1 >>
rect 104 187 105 188 
<< m2 >>
rect 104 187 105 188 
<< m1 >>
rect 105 187 106 188 
<< m2 >>
rect 105 187 106 188 
<< m1 >>
rect 106 187 107 188 
<< m2 >>
rect 106 187 107 188 
<< m1 >>
rect 107 187 108 188 
<< m2 >>
rect 107 187 108 188 
<< m1 >>
rect 108 187 109 188 
<< m2 >>
rect 108 187 109 188 
<< m1 >>
rect 109 187 110 188 
<< m2 >>
rect 109 187 110 188 
<< m1 >>
rect 110 187 111 188 
<< m2 >>
rect 110 187 111 188 
<< m1 >>
rect 111 187 112 188 
<< m2 >>
rect 111 187 112 188 
<< m1 >>
rect 112 187 113 188 
<< m2 >>
rect 112 187 113 188 
<< m1 >>
rect 113 187 114 188 
<< m2 >>
rect 113 187 114 188 
<< m1 >>
rect 114 187 115 188 
<< m2 >>
rect 114 187 115 188 
<< m1 >>
rect 115 187 116 188 
<< m2 >>
rect 115 187 116 188 
<< m1 >>
rect 116 187 117 188 
<< m2 >>
rect 116 187 117 188 
<< m1 >>
rect 117 187 118 188 
<< m2 >>
rect 117 187 118 188 
<< m1 >>
rect 118 187 119 188 
<< m2 >>
rect 118 187 119 188 
<< m1 >>
rect 119 187 120 188 
<< m1 >>
rect 120 187 121 188 
<< m1 >>
rect 121 187 122 188 
<< m1 >>
rect 122 187 123 188 
<< m2 >>
rect 122 187 123 188 
<< m1 >>
rect 123 187 124 188 
<< m1 >>
rect 124 187 125 188 
<< m1 >>
rect 125 187 126 188 
<< m1 >>
rect 126 187 127 188 
<< m1 >>
rect 127 187 128 188 
<< m2 >>
rect 127 187 128 188 
<< m1 >>
rect 128 187 129 188 
<< m1 >>
rect 129 187 130 188 
<< m1 >>
rect 130 187 131 188 
<< m2 >>
rect 130 187 131 188 
<< m1 >>
rect 131 187 132 188 
<< m1 >>
rect 132 187 133 188 
<< m2 >>
rect 132 187 133 188 
<< m1 >>
rect 133 187 134 188 
<< m1 >>
rect 134 187 135 188 
<< m1 >>
rect 135 187 136 188 
<< m1 >>
rect 136 187 137 188 
<< m2 >>
rect 136 187 137 188 
<< m1 >>
rect 137 187 138 188 
<< m1 >>
rect 138 187 139 188 
<< m1 >>
rect 139 187 140 188 
<< m1 >>
rect 140 187 141 188 
<< m1 >>
rect 141 187 142 188 
<< m2 >>
rect 141 187 142 188 
<< m1 >>
rect 142 187 143 188 
<< m1 >>
rect 143 187 144 188 
<< m2 >>
rect 143 187 144 188 
<< m2c >>
rect 143 187 144 188 
<< m1 >>
rect 143 187 144 188 
<< m2 >>
rect 143 187 144 188 
<< m2 >>
rect 144 187 145 188 
<< m1 >>
rect 145 187 146 188 
<< m2 >>
rect 145 187 146 188 
<< m2 >>
rect 146 187 147 188 
<< m1 >>
rect 147 187 148 188 
<< m2 >>
rect 147 187 148 188 
<< m2c >>
rect 147 187 148 188 
<< m1 >>
rect 147 187 148 188 
<< m2 >>
rect 147 187 148 188 
<< m1 >>
rect 148 187 149 188 
<< m1 >>
rect 149 187 150 188 
<< m1 >>
rect 163 187 164 188 
<< m1 >>
rect 165 187 166 188 
<< m1 >>
rect 170 187 171 188 
<< m1 >>
rect 172 187 173 188 
<< m1 >>
rect 181 187 182 188 
<< m1 >>
rect 183 187 184 188 
<< m1 >>
rect 188 187 189 188 
<< m1 >>
rect 190 187 191 188 
<< m1 >>
rect 199 187 200 188 
<< m1 >>
rect 201 187 202 188 
<< m2 >>
rect 225 187 226 188 
<< m1 >>
rect 226 187 227 188 
<< m1 >>
rect 232 187 233 188 
<< m1 >>
rect 235 187 236 188 
<< m1 >>
rect 237 187 238 188 
<< m1 >>
rect 241 187 242 188 
<< m1 >>
rect 243 187 244 188 
<< m1 >>
rect 253 187 254 188 
<< m1 >>
rect 255 187 256 188 
<< m1 >>
rect 260 187 261 188 
<< m1 >>
rect 262 187 263 188 
<< m2 >>
rect 262 187 263 188 
<< m2 >>
rect 271 187 272 188 
<< m1 >>
rect 272 187 273 188 
<< m1 >>
rect 274 187 275 188 
<< m2 >>
rect 275 187 276 188 
<< m1 >>
rect 289 187 290 188 
<< m1 >>
rect 291 187 292 188 
<< m1 >>
rect 292 187 293 188 
<< m1 >>
rect 293 187 294 188 
<< m1 >>
rect 294 187 295 188 
<< m1 >>
rect 295 187 296 188 
<< m1 >>
rect 296 187 297 188 
<< m1 >>
rect 297 187 298 188 
<< m1 >>
rect 298 187 299 188 
<< m1 >>
rect 299 187 300 188 
<< m1 >>
rect 300 187 301 188 
<< m1 >>
rect 301 187 302 188 
<< m1 >>
rect 302 187 303 188 
<< m1 >>
rect 303 187 304 188 
<< m1 >>
rect 304 187 305 188 
<< m1 >>
rect 305 187 306 188 
<< m2 >>
rect 305 187 306 188 
<< m2c >>
rect 305 187 306 188 
<< m1 >>
rect 305 187 306 188 
<< m2 >>
rect 305 187 306 188 
<< m2 >>
rect 306 187 307 188 
<< m1 >>
rect 307 187 308 188 
<< m2 >>
rect 308 187 309 188 
<< m1 >>
rect 309 187 310 188 
<< m2 >>
rect 309 187 310 188 
<< m2c >>
rect 309 187 310 188 
<< m1 >>
rect 309 187 310 188 
<< m2 >>
rect 309 187 310 188 
<< m1 >>
rect 310 187 311 188 
<< m1 >>
rect 311 187 312 188 
<< m2 >>
rect 311 187 312 188 
<< m1 >>
rect 312 187 313 188 
<< m2 >>
rect 312 187 313 188 
<< m1 >>
rect 313 187 314 188 
<< m2 >>
rect 313 187 314 188 
<< m1 >>
rect 314 187 315 188 
<< m2 >>
rect 314 187 315 188 
<< m1 >>
rect 315 187 316 188 
<< m2 >>
rect 315 187 316 188 
<< m1 >>
rect 316 187 317 188 
<< m2 >>
rect 316 187 317 188 
<< m1 >>
rect 317 187 318 188 
<< m2 >>
rect 317 187 318 188 
<< m1 >>
rect 318 187 319 188 
<< m2 >>
rect 318 187 319 188 
<< m1 >>
rect 319 187 320 188 
<< m2 >>
rect 319 187 320 188 
<< m1 >>
rect 320 187 321 188 
<< m2 >>
rect 320 187 321 188 
<< m1 >>
rect 321 187 322 188 
<< m2 >>
rect 321 187 322 188 
<< m1 >>
rect 322 187 323 188 
<< m2 >>
rect 322 187 323 188 
<< m1 >>
rect 323 187 324 188 
<< m2 >>
rect 323 187 324 188 
<< m1 >>
rect 324 187 325 188 
<< m2 >>
rect 324 187 325 188 
<< m1 >>
rect 325 187 326 188 
<< m2 >>
rect 325 187 326 188 
<< m2 >>
rect 326 187 327 188 
<< m1 >>
rect 327 187 328 188 
<< m1 >>
rect 343 187 344 188 
<< m2 >>
rect 343 187 344 188 
<< m1 >>
rect 345 187 346 188 
<< m1 >>
rect 10 188 11 189 
<< m1 >>
rect 19 188 20 189 
<< m1 >>
rect 21 188 22 189 
<< m1 >>
rect 23 188 24 189 
<< m2 >>
rect 27 188 28 189 
<< m1 >>
rect 28 188 29 189 
<< m1 >>
rect 37 188 38 189 
<< m2 >>
rect 38 188 39 189 
<< m1 >>
rect 44 188 45 189 
<< m1 >>
rect 46 188 47 189 
<< m1 >>
rect 56 188 57 189 
<< m1 >>
rect 58 188 59 189 
<< m1 >>
rect 62 188 63 189 
<< m1 >>
rect 64 188 65 189 
<< m1 >>
rect 70 188 71 189 
<< m1 >>
rect 72 188 73 189 
<< m2 >>
rect 74 188 75 189 
<< m2 >>
rect 80 188 81 189 
<< m2 >>
rect 82 188 83 189 
<< m2 >>
rect 118 188 119 189 
<< m2 >>
rect 122 188 123 189 
<< m2 >>
rect 127 188 128 189 
<< m2 >>
rect 130 188 131 189 
<< m2 >>
rect 132 188 133 189 
<< m2 >>
rect 136 188 137 189 
<< m2 >>
rect 141 188 142 189 
<< m1 >>
rect 145 188 146 189 
<< m1 >>
rect 163 188 164 189 
<< m1 >>
rect 165 188 166 189 
<< m1 >>
rect 170 188 171 189 
<< m1 >>
rect 172 188 173 189 
<< m1 >>
rect 181 188 182 189 
<< m2 >>
rect 181 188 182 189 
<< m2c >>
rect 181 188 182 189 
<< m1 >>
rect 181 188 182 189 
<< m2 >>
rect 181 188 182 189 
<< m1 >>
rect 183 188 184 189 
<< m2 >>
rect 183 188 184 189 
<< m2c >>
rect 183 188 184 189 
<< m1 >>
rect 183 188 184 189 
<< m2 >>
rect 183 188 184 189 
<< m1 >>
rect 188 188 189 189 
<< m2 >>
rect 188 188 189 189 
<< m2c >>
rect 188 188 189 189 
<< m1 >>
rect 188 188 189 189 
<< m2 >>
rect 188 188 189 189 
<< m1 >>
rect 190 188 191 189 
<< m2 >>
rect 190 188 191 189 
<< m2c >>
rect 190 188 191 189 
<< m1 >>
rect 190 188 191 189 
<< m2 >>
rect 190 188 191 189 
<< m1 >>
rect 199 188 200 189 
<< m1 >>
rect 201 188 202 189 
<< m2 >>
rect 225 188 226 189 
<< m1 >>
rect 226 188 227 189 
<< m1 >>
rect 232 188 233 189 
<< m1 >>
rect 235 188 236 189 
<< m1 >>
rect 237 188 238 189 
<< m1 >>
rect 241 188 242 189 
<< m1 >>
rect 243 188 244 189 
<< m1 >>
rect 253 188 254 189 
<< m1 >>
rect 255 188 256 189 
<< m1 >>
rect 260 188 261 189 
<< m1 >>
rect 262 188 263 189 
<< m2 >>
rect 262 188 263 189 
<< m2 >>
rect 271 188 272 189 
<< m1 >>
rect 272 188 273 189 
<< m1 >>
rect 274 188 275 189 
<< m2 >>
rect 275 188 276 189 
<< m1 >>
rect 289 188 290 189 
<< m1 >>
rect 291 188 292 189 
<< m2 >>
rect 306 188 307 189 
<< m1 >>
rect 307 188 308 189 
<< m2 >>
rect 311 188 312 189 
<< m1 >>
rect 325 188 326 189 
<< m1 >>
rect 327 188 328 189 
<< m1 >>
rect 343 188 344 189 
<< m2 >>
rect 343 188 344 189 
<< m1 >>
rect 345 188 346 189 
<< m1 >>
rect 10 189 11 190 
<< m1 >>
rect 19 189 20 190 
<< m1 >>
rect 21 189 22 190 
<< m1 >>
rect 23 189 24 190 
<< m2 >>
rect 27 189 28 190 
<< m1 >>
rect 28 189 29 190 
<< m1 >>
rect 37 189 38 190 
<< m2 >>
rect 38 189 39 190 
<< m1 >>
rect 44 189 45 190 
<< m1 >>
rect 46 189 47 190 
<< m1 >>
rect 56 189 57 190 
<< m1 >>
rect 58 189 59 190 
<< m1 >>
rect 62 189 63 190 
<< m1 >>
rect 64 189 65 190 
<< m2 >>
rect 69 189 70 190 
<< m1 >>
rect 70 189 71 190 
<< m2 >>
rect 70 189 71 190 
<< m2 >>
rect 71 189 72 190 
<< m1 >>
rect 72 189 73 190 
<< m2 >>
rect 72 189 73 190 
<< m2c >>
rect 72 189 73 190 
<< m1 >>
rect 72 189 73 190 
<< m2 >>
rect 72 189 73 190 
<< m1 >>
rect 74 189 75 190 
<< m2 >>
rect 74 189 75 190 
<< m2c >>
rect 74 189 75 190 
<< m1 >>
rect 74 189 75 190 
<< m2 >>
rect 74 189 75 190 
<< m1 >>
rect 80 189 81 190 
<< m2 >>
rect 80 189 81 190 
<< m2c >>
rect 80 189 81 190 
<< m1 >>
rect 80 189 81 190 
<< m2 >>
rect 80 189 81 190 
<< m1 >>
rect 82 189 83 190 
<< m2 >>
rect 82 189 83 190 
<< m2c >>
rect 82 189 83 190 
<< m1 >>
rect 82 189 83 190 
<< m2 >>
rect 82 189 83 190 
<< m1 >>
rect 118 189 119 190 
<< m2 >>
rect 118 189 119 190 
<< m2c >>
rect 118 189 119 190 
<< m1 >>
rect 118 189 119 190 
<< m2 >>
rect 118 189 119 190 
<< m1 >>
rect 122 189 123 190 
<< m2 >>
rect 122 189 123 190 
<< m2c >>
rect 122 189 123 190 
<< m1 >>
rect 122 189 123 190 
<< m2 >>
rect 122 189 123 190 
<< m1 >>
rect 123 189 124 190 
<< m1 >>
rect 124 189 125 190 
<< m1 >>
rect 125 189 126 190 
<< m1 >>
rect 126 189 127 190 
<< m1 >>
rect 127 189 128 190 
<< m2 >>
rect 127 189 128 190 
<< m1 >>
rect 130 189 131 190 
<< m2 >>
rect 130 189 131 190 
<< m2c >>
rect 130 189 131 190 
<< m1 >>
rect 130 189 131 190 
<< m2 >>
rect 130 189 131 190 
<< m1 >>
rect 132 189 133 190 
<< m2 >>
rect 132 189 133 190 
<< m2c >>
rect 132 189 133 190 
<< m1 >>
rect 132 189 133 190 
<< m2 >>
rect 132 189 133 190 
<< m1 >>
rect 136 189 137 190 
<< m2 >>
rect 136 189 137 190 
<< m2c >>
rect 136 189 137 190 
<< m1 >>
rect 136 189 137 190 
<< m2 >>
rect 136 189 137 190 
<< m1 >>
rect 141 189 142 190 
<< m2 >>
rect 141 189 142 190 
<< m2c >>
rect 141 189 142 190 
<< m1 >>
rect 141 189 142 190 
<< m2 >>
rect 141 189 142 190 
<< m1 >>
rect 142 189 143 190 
<< m1 >>
rect 143 189 144 190 
<< m1 >>
rect 145 189 146 190 
<< m1 >>
rect 163 189 164 190 
<< m1 >>
rect 165 189 166 190 
<< m1 >>
rect 170 189 171 190 
<< m1 >>
rect 172 189 173 190 
<< m2 >>
rect 181 189 182 190 
<< m2 >>
rect 183 189 184 190 
<< m2 >>
rect 188 189 189 190 
<< m2 >>
rect 190 189 191 190 
<< m1 >>
rect 199 189 200 190 
<< m1 >>
rect 201 189 202 190 
<< m1 >>
rect 211 189 212 190 
<< m1 >>
rect 212 189 213 190 
<< m1 >>
rect 213 189 214 190 
<< m1 >>
rect 214 189 215 190 
<< m1 >>
rect 215 189 216 190 
<< m1 >>
rect 216 189 217 190 
<< m1 >>
rect 217 189 218 190 
<< m1 >>
rect 218 189 219 190 
<< m2 >>
rect 225 189 226 190 
<< m1 >>
rect 226 189 227 190 
<< m1 >>
rect 232 189 233 190 
<< m1 >>
rect 235 189 236 190 
<< m1 >>
rect 237 189 238 190 
<< m1 >>
rect 241 189 242 190 
<< m1 >>
rect 243 189 244 190 
<< m1 >>
rect 253 189 254 190 
<< m1 >>
rect 255 189 256 190 
<< m1 >>
rect 260 189 261 190 
<< m1 >>
rect 262 189 263 190 
<< m2 >>
rect 262 189 263 190 
<< m2 >>
rect 271 189 272 190 
<< m1 >>
rect 272 189 273 190 
<< m1 >>
rect 274 189 275 190 
<< m2 >>
rect 275 189 276 190 
<< m1 >>
rect 283 189 284 190 
<< m1 >>
rect 284 189 285 190 
<< m1 >>
rect 285 189 286 190 
<< m1 >>
rect 286 189 287 190 
<< m1 >>
rect 287 189 288 190 
<< m2 >>
rect 287 189 288 190 
<< m2c >>
rect 287 189 288 190 
<< m1 >>
rect 287 189 288 190 
<< m2 >>
rect 287 189 288 190 
<< m2 >>
rect 288 189 289 190 
<< m1 >>
rect 289 189 290 190 
<< m2 >>
rect 289 189 290 190 
<< m2 >>
rect 290 189 291 190 
<< m1 >>
rect 291 189 292 190 
<< m2 >>
rect 291 189 292 190 
<< m2c >>
rect 291 189 292 190 
<< m1 >>
rect 291 189 292 190 
<< m2 >>
rect 291 189 292 190 
<< m2 >>
rect 306 189 307 190 
<< m1 >>
rect 307 189 308 190 
<< m2 >>
rect 307 189 308 190 
<< m2 >>
rect 308 189 309 190 
<< m1 >>
rect 309 189 310 190 
<< m2 >>
rect 309 189 310 190 
<< m2c >>
rect 309 189 310 190 
<< m1 >>
rect 309 189 310 190 
<< m2 >>
rect 309 189 310 190 
<< m1 >>
rect 310 189 311 190 
<< m1 >>
rect 311 189 312 190 
<< m2 >>
rect 311 189 312 190 
<< m2c >>
rect 311 189 312 190 
<< m1 >>
rect 311 189 312 190 
<< m2 >>
rect 311 189 312 190 
<< m1 >>
rect 325 189 326 190 
<< m1 >>
rect 327 189 328 190 
<< m1 >>
rect 343 189 344 190 
<< m2 >>
rect 343 189 344 190 
<< m1 >>
rect 345 189 346 190 
<< m1 >>
rect 10 190 11 191 
<< m1 >>
rect 16 190 17 191 
<< m1 >>
rect 17 190 18 191 
<< m2 >>
rect 17 190 18 191 
<< m2c >>
rect 17 190 18 191 
<< m1 >>
rect 17 190 18 191 
<< m2 >>
rect 17 190 18 191 
<< m2 >>
rect 18 190 19 191 
<< m1 >>
rect 19 190 20 191 
<< m2 >>
rect 19 190 20 191 
<< m2 >>
rect 20 190 21 191 
<< m1 >>
rect 21 190 22 191 
<< m2 >>
rect 21 190 22 191 
<< m2 >>
rect 22 190 23 191 
<< m1 >>
rect 23 190 24 191 
<< m2 >>
rect 23 190 24 191 
<< m2c >>
rect 23 190 24 191 
<< m1 >>
rect 23 190 24 191 
<< m2 >>
rect 23 190 24 191 
<< m2 >>
rect 27 190 28 191 
<< m1 >>
rect 28 190 29 191 
<< m1 >>
rect 37 190 38 191 
<< m2 >>
rect 38 190 39 191 
<< m1 >>
rect 44 190 45 191 
<< m1 >>
rect 46 190 47 191 
<< m1 >>
rect 56 190 57 191 
<< m1 >>
rect 58 190 59 191 
<< m1 >>
rect 62 190 63 191 
<< m1 >>
rect 64 190 65 191 
<< m1 >>
rect 67 190 68 191 
<< m1 >>
rect 68 190 69 191 
<< m2 >>
rect 68 190 69 191 
<< m2c >>
rect 68 190 69 191 
<< m1 >>
rect 68 190 69 191 
<< m2 >>
rect 68 190 69 191 
<< m2 >>
rect 69 190 70 191 
<< m1 >>
rect 70 190 71 191 
<< m1 >>
rect 74 190 75 191 
<< m1 >>
rect 80 190 81 191 
<< m1 >>
rect 82 190 83 191 
<< m1 >>
rect 118 190 119 191 
<< m1 >>
rect 127 190 128 191 
<< m2 >>
rect 127 190 128 191 
<< m2 >>
rect 130 190 131 191 
<< m2 >>
rect 132 190 133 191 
<< m1 >>
rect 136 190 137 191 
<< m1 >>
rect 143 190 144 191 
<< m2 >>
rect 143 190 144 191 
<< m2c >>
rect 143 190 144 191 
<< m1 >>
rect 143 190 144 191 
<< m2 >>
rect 143 190 144 191 
<< m2 >>
rect 144 190 145 191 
<< m1 >>
rect 145 190 146 191 
<< m2 >>
rect 145 190 146 191 
<< m2 >>
rect 146 190 147 191 
<< m1 >>
rect 163 190 164 191 
<< m1 >>
rect 165 190 166 191 
<< m1 >>
rect 170 190 171 191 
<< m1 >>
rect 172 190 173 191 
<< m1 >>
rect 181 190 182 191 
<< m2 >>
rect 181 190 182 191 
<< m1 >>
rect 182 190 183 191 
<< m1 >>
rect 183 190 184 191 
<< m2 >>
rect 183 190 184 191 
<< m1 >>
rect 184 190 185 191 
<< m1 >>
rect 185 190 186 191 
<< m1 >>
rect 186 190 187 191 
<< m1 >>
rect 187 190 188 191 
<< m1 >>
rect 188 190 189 191 
<< m2 >>
rect 188 190 189 191 
<< m1 >>
rect 189 190 190 191 
<< m1 >>
rect 190 190 191 191 
<< m2 >>
rect 190 190 191 191 
<< m1 >>
rect 191 190 192 191 
<< m1 >>
rect 192 190 193 191 
<< m1 >>
rect 193 190 194 191 
<< m1 >>
rect 196 190 197 191 
<< m1 >>
rect 197 190 198 191 
<< m2 >>
rect 197 190 198 191 
<< m2c >>
rect 197 190 198 191 
<< m1 >>
rect 197 190 198 191 
<< m2 >>
rect 197 190 198 191 
<< m2 >>
rect 198 190 199 191 
<< m1 >>
rect 199 190 200 191 
<< m2 >>
rect 199 190 200 191 
<< m1 >>
rect 201 190 202 191 
<< m1 >>
rect 211 190 212 191 
<< m1 >>
rect 218 190 219 191 
<< m2 >>
rect 225 190 226 191 
<< m1 >>
rect 226 190 227 191 
<< m1 >>
rect 232 190 233 191 
<< m1 >>
rect 235 190 236 191 
<< m1 >>
rect 237 190 238 191 
<< m1 >>
rect 241 190 242 191 
<< m1 >>
rect 243 190 244 191 
<< m1 >>
rect 253 190 254 191 
<< m1 >>
rect 255 190 256 191 
<< m1 >>
rect 260 190 261 191 
<< m1 >>
rect 262 190 263 191 
<< m2 >>
rect 262 190 263 191 
<< m2 >>
rect 271 190 272 191 
<< m1 >>
rect 272 190 273 191 
<< m1 >>
rect 274 190 275 191 
<< m2 >>
rect 275 190 276 191 
<< m1 >>
rect 283 190 284 191 
<< m1 >>
rect 289 190 290 191 
<< m1 >>
rect 307 190 308 191 
<< m1 >>
rect 325 190 326 191 
<< m1 >>
rect 327 190 328 191 
<< m1 >>
rect 343 190 344 191 
<< m2 >>
rect 343 190 344 191 
<< m1 >>
rect 345 190 346 191 
<< m1 >>
rect 10 191 11 192 
<< m1 >>
rect 16 191 17 192 
<< m1 >>
rect 19 191 20 192 
<< m1 >>
rect 21 191 22 192 
<< m2 >>
rect 27 191 28 192 
<< m1 >>
rect 28 191 29 192 
<< m1 >>
rect 37 191 38 192 
<< m2 >>
rect 38 191 39 192 
<< m1 >>
rect 44 191 45 192 
<< m1 >>
rect 46 191 47 192 
<< m1 >>
rect 56 191 57 192 
<< m1 >>
rect 58 191 59 192 
<< m1 >>
rect 62 191 63 192 
<< m1 >>
rect 64 191 65 192 
<< m1 >>
rect 67 191 68 192 
<< m1 >>
rect 70 191 71 192 
<< m1 >>
rect 74 191 75 192 
<< m1 >>
rect 75 191 76 192 
<< m1 >>
rect 76 191 77 192 
<< m1 >>
rect 77 191 78 192 
<< m1 >>
rect 78 191 79 192 
<< m2 >>
rect 78 191 79 192 
<< m2c >>
rect 78 191 79 192 
<< m1 >>
rect 78 191 79 192 
<< m2 >>
rect 78 191 79 192 
<< m2 >>
rect 79 191 80 192 
<< m1 >>
rect 80 191 81 192 
<< m1 >>
rect 82 191 83 192 
<< m1 >>
rect 118 191 119 192 
<< m1 >>
rect 127 191 128 192 
<< m2 >>
rect 127 191 128 192 
<< m1 >>
rect 128 191 129 192 
<< m1 >>
rect 129 191 130 192 
<< m1 >>
rect 130 191 131 192 
<< m2 >>
rect 130 191 131 192 
<< m1 >>
rect 131 191 132 192 
<< m1 >>
rect 132 191 133 192 
<< m2 >>
rect 132 191 133 192 
<< m1 >>
rect 133 191 134 192 
<< m1 >>
rect 134 191 135 192 
<< m2 >>
rect 134 191 135 192 
<< m2c >>
rect 134 191 135 192 
<< m1 >>
rect 134 191 135 192 
<< m2 >>
rect 134 191 135 192 
<< m2 >>
rect 135 191 136 192 
<< m1 >>
rect 136 191 137 192 
<< m1 >>
rect 145 191 146 192 
<< m2 >>
rect 146 191 147 192 
<< m1 >>
rect 163 191 164 192 
<< m1 >>
rect 165 191 166 192 
<< m1 >>
rect 170 191 171 192 
<< m1 >>
rect 172 191 173 192 
<< m1 >>
rect 181 191 182 192 
<< m2 >>
rect 181 191 182 192 
<< m2 >>
rect 183 191 184 192 
<< m2 >>
rect 188 191 189 192 
<< m2 >>
rect 190 191 191 192 
<< m1 >>
rect 193 191 194 192 
<< m1 >>
rect 196 191 197 192 
<< m1 >>
rect 199 191 200 192 
<< m2 >>
rect 199 191 200 192 
<< m1 >>
rect 201 191 202 192 
<< m1 >>
rect 211 191 212 192 
<< m1 >>
rect 218 191 219 192 
<< m2 >>
rect 225 191 226 192 
<< m1 >>
rect 226 191 227 192 
<< m1 >>
rect 232 191 233 192 
<< m1 >>
rect 235 191 236 192 
<< m1 >>
rect 237 191 238 192 
<< m1 >>
rect 241 191 242 192 
<< m1 >>
rect 243 191 244 192 
<< m1 >>
rect 253 191 254 192 
<< m1 >>
rect 255 191 256 192 
<< m1 >>
rect 260 191 261 192 
<< m1 >>
rect 262 191 263 192 
<< m2 >>
rect 262 191 263 192 
<< m2 >>
rect 271 191 272 192 
<< m1 >>
rect 272 191 273 192 
<< m1 >>
rect 274 191 275 192 
<< m2 >>
rect 275 191 276 192 
<< m1 >>
rect 283 191 284 192 
<< m1 >>
rect 289 191 290 192 
<< m1 >>
rect 307 191 308 192 
<< m1 >>
rect 325 191 326 192 
<< m1 >>
rect 327 191 328 192 
<< m1 >>
rect 343 191 344 192 
<< m2 >>
rect 343 191 344 192 
<< m1 >>
rect 345 191 346 192 
<< m1 >>
rect 10 192 11 193 
<< pdiffusion >>
rect 12 192 13 193 
<< pdiffusion >>
rect 13 192 14 193 
<< pdiffusion >>
rect 14 192 15 193 
<< pdiffusion >>
rect 15 192 16 193 
<< m1 >>
rect 16 192 17 193 
<< pdiffusion >>
rect 16 192 17 193 
<< pdiffusion >>
rect 17 192 18 193 
<< m1 >>
rect 19 192 20 193 
<< m1 >>
rect 21 192 22 193 
<< m2 >>
rect 27 192 28 193 
<< m1 >>
rect 28 192 29 193 
<< pdiffusion >>
rect 30 192 31 193 
<< pdiffusion >>
rect 31 192 32 193 
<< pdiffusion >>
rect 32 192 33 193 
<< pdiffusion >>
rect 33 192 34 193 
<< pdiffusion >>
rect 34 192 35 193 
<< pdiffusion >>
rect 35 192 36 193 
<< m1 >>
rect 37 192 38 193 
<< m2 >>
rect 38 192 39 193 
<< m1 >>
rect 44 192 45 193 
<< m1 >>
rect 46 192 47 193 
<< pdiffusion >>
rect 48 192 49 193 
<< pdiffusion >>
rect 49 192 50 193 
<< pdiffusion >>
rect 50 192 51 193 
<< pdiffusion >>
rect 51 192 52 193 
<< pdiffusion >>
rect 52 192 53 193 
<< pdiffusion >>
rect 53 192 54 193 
<< m1 >>
rect 56 192 57 193 
<< m1 >>
rect 58 192 59 193 
<< m1 >>
rect 62 192 63 193 
<< m1 >>
rect 64 192 65 193 
<< pdiffusion >>
rect 66 192 67 193 
<< m1 >>
rect 67 192 68 193 
<< pdiffusion >>
rect 67 192 68 193 
<< pdiffusion >>
rect 68 192 69 193 
<< pdiffusion >>
rect 69 192 70 193 
<< m1 >>
rect 70 192 71 193 
<< pdiffusion >>
rect 70 192 71 193 
<< pdiffusion >>
rect 71 192 72 193 
<< m2 >>
rect 79 192 80 193 
<< m1 >>
rect 80 192 81 193 
<< m1 >>
rect 82 192 83 193 
<< pdiffusion >>
rect 84 192 85 193 
<< pdiffusion >>
rect 85 192 86 193 
<< pdiffusion >>
rect 86 192 87 193 
<< pdiffusion >>
rect 87 192 88 193 
<< pdiffusion >>
rect 88 192 89 193 
<< pdiffusion >>
rect 89 192 90 193 
<< pdiffusion >>
rect 102 192 103 193 
<< pdiffusion >>
rect 103 192 104 193 
<< pdiffusion >>
rect 104 192 105 193 
<< pdiffusion >>
rect 105 192 106 193 
<< pdiffusion >>
rect 106 192 107 193 
<< pdiffusion >>
rect 107 192 108 193 
<< m1 >>
rect 118 192 119 193 
<< pdiffusion >>
rect 120 192 121 193 
<< pdiffusion >>
rect 121 192 122 193 
<< pdiffusion >>
rect 122 192 123 193 
<< pdiffusion >>
rect 123 192 124 193 
<< pdiffusion >>
rect 124 192 125 193 
<< pdiffusion >>
rect 125 192 126 193 
<< m2 >>
rect 127 192 128 193 
<< m2 >>
rect 130 192 131 193 
<< m2 >>
rect 132 192 133 193 
<< m2 >>
rect 135 192 136 193 
<< m1 >>
rect 136 192 137 193 
<< pdiffusion >>
rect 138 192 139 193 
<< pdiffusion >>
rect 139 192 140 193 
<< pdiffusion >>
rect 140 192 141 193 
<< pdiffusion >>
rect 141 192 142 193 
<< pdiffusion >>
rect 142 192 143 193 
<< pdiffusion >>
rect 143 192 144 193 
<< m1 >>
rect 145 192 146 193 
<< m2 >>
rect 146 192 147 193 
<< pdiffusion >>
rect 156 192 157 193 
<< pdiffusion >>
rect 157 192 158 193 
<< pdiffusion >>
rect 158 192 159 193 
<< pdiffusion >>
rect 159 192 160 193 
<< pdiffusion >>
rect 160 192 161 193 
<< pdiffusion >>
rect 161 192 162 193 
<< m1 >>
rect 163 192 164 193 
<< m1 >>
rect 165 192 166 193 
<< m1 >>
rect 170 192 171 193 
<< m1 >>
rect 172 192 173 193 
<< pdiffusion >>
rect 174 192 175 193 
<< pdiffusion >>
rect 175 192 176 193 
<< pdiffusion >>
rect 176 192 177 193 
<< pdiffusion >>
rect 177 192 178 193 
<< pdiffusion >>
rect 178 192 179 193 
<< pdiffusion >>
rect 179 192 180 193 
<< m1 >>
rect 181 192 182 193 
<< m2 >>
rect 181 192 182 193 
<< m1 >>
rect 183 192 184 193 
<< m2 >>
rect 183 192 184 193 
<< m2c >>
rect 183 192 184 193 
<< m1 >>
rect 183 192 184 193 
<< m2 >>
rect 183 192 184 193 
<< m1 >>
rect 188 192 189 193 
<< m2 >>
rect 188 192 189 193 
<< m2c >>
rect 188 192 189 193 
<< m1 >>
rect 188 192 189 193 
<< m2 >>
rect 188 192 189 193 
<< m1 >>
rect 190 192 191 193 
<< m2 >>
rect 190 192 191 193 
<< m2c >>
rect 190 192 191 193 
<< m1 >>
rect 190 192 191 193 
<< m2 >>
rect 190 192 191 193 
<< pdiffusion >>
rect 192 192 193 193 
<< m1 >>
rect 193 192 194 193 
<< pdiffusion >>
rect 193 192 194 193 
<< pdiffusion >>
rect 194 192 195 193 
<< pdiffusion >>
rect 195 192 196 193 
<< m1 >>
rect 196 192 197 193 
<< pdiffusion >>
rect 196 192 197 193 
<< pdiffusion >>
rect 197 192 198 193 
<< m1 >>
rect 199 192 200 193 
<< m2 >>
rect 199 192 200 193 
<< m1 >>
rect 201 192 202 193 
<< pdiffusion >>
rect 210 192 211 193 
<< m1 >>
rect 211 192 212 193 
<< pdiffusion >>
rect 211 192 212 193 
<< pdiffusion >>
rect 212 192 213 193 
<< pdiffusion >>
rect 213 192 214 193 
<< pdiffusion >>
rect 214 192 215 193 
<< pdiffusion >>
rect 215 192 216 193 
<< m1 >>
rect 218 192 219 193 
<< m2 >>
rect 225 192 226 193 
<< m1 >>
rect 226 192 227 193 
<< pdiffusion >>
rect 228 192 229 193 
<< pdiffusion >>
rect 229 192 230 193 
<< pdiffusion >>
rect 230 192 231 193 
<< pdiffusion >>
rect 231 192 232 193 
<< m1 >>
rect 232 192 233 193 
<< pdiffusion >>
rect 232 192 233 193 
<< pdiffusion >>
rect 233 192 234 193 
<< m1 >>
rect 235 192 236 193 
<< m1 >>
rect 237 192 238 193 
<< m1 >>
rect 241 192 242 193 
<< m1 >>
rect 243 192 244 193 
<< pdiffusion >>
rect 246 192 247 193 
<< pdiffusion >>
rect 247 192 248 193 
<< pdiffusion >>
rect 248 192 249 193 
<< pdiffusion >>
rect 249 192 250 193 
<< pdiffusion >>
rect 250 192 251 193 
<< pdiffusion >>
rect 251 192 252 193 
<< m1 >>
rect 253 192 254 193 
<< m1 >>
rect 255 192 256 193 
<< m1 >>
rect 260 192 261 193 
<< m1 >>
rect 262 192 263 193 
<< m2 >>
rect 262 192 263 193 
<< pdiffusion >>
rect 264 192 265 193 
<< pdiffusion >>
rect 265 192 266 193 
<< pdiffusion >>
rect 266 192 267 193 
<< pdiffusion >>
rect 267 192 268 193 
<< pdiffusion >>
rect 268 192 269 193 
<< pdiffusion >>
rect 269 192 270 193 
<< m2 >>
rect 271 192 272 193 
<< m1 >>
rect 272 192 273 193 
<< m1 >>
rect 274 192 275 193 
<< m2 >>
rect 275 192 276 193 
<< pdiffusion >>
rect 282 192 283 193 
<< m1 >>
rect 283 192 284 193 
<< pdiffusion >>
rect 283 192 284 193 
<< pdiffusion >>
rect 284 192 285 193 
<< pdiffusion >>
rect 285 192 286 193 
<< pdiffusion >>
rect 286 192 287 193 
<< pdiffusion >>
rect 287 192 288 193 
<< m1 >>
rect 289 192 290 193 
<< pdiffusion >>
rect 300 192 301 193 
<< pdiffusion >>
rect 301 192 302 193 
<< pdiffusion >>
rect 302 192 303 193 
<< pdiffusion >>
rect 303 192 304 193 
<< pdiffusion >>
rect 304 192 305 193 
<< pdiffusion >>
rect 305 192 306 193 
<< m1 >>
rect 307 192 308 193 
<< pdiffusion >>
rect 318 192 319 193 
<< pdiffusion >>
rect 319 192 320 193 
<< pdiffusion >>
rect 320 192 321 193 
<< pdiffusion >>
rect 321 192 322 193 
<< pdiffusion >>
rect 322 192 323 193 
<< pdiffusion >>
rect 323 192 324 193 
<< m1 >>
rect 325 192 326 193 
<< m1 >>
rect 327 192 328 193 
<< pdiffusion >>
rect 336 192 337 193 
<< pdiffusion >>
rect 337 192 338 193 
<< pdiffusion >>
rect 338 192 339 193 
<< pdiffusion >>
rect 339 192 340 193 
<< pdiffusion >>
rect 340 192 341 193 
<< pdiffusion >>
rect 341 192 342 193 
<< m1 >>
rect 343 192 344 193 
<< m2 >>
rect 343 192 344 193 
<< m1 >>
rect 345 192 346 193 
<< m1 >>
rect 10 193 11 194 
<< pdiffusion >>
rect 12 193 13 194 
<< pdiffusion >>
rect 13 193 14 194 
<< pdiffusion >>
rect 14 193 15 194 
<< pdiffusion >>
rect 15 193 16 194 
<< pdiffusion >>
rect 16 193 17 194 
<< pdiffusion >>
rect 17 193 18 194 
<< m1 >>
rect 19 193 20 194 
<< m1 >>
rect 21 193 22 194 
<< m2 >>
rect 27 193 28 194 
<< m1 >>
rect 28 193 29 194 
<< pdiffusion >>
rect 30 193 31 194 
<< pdiffusion >>
rect 31 193 32 194 
<< pdiffusion >>
rect 32 193 33 194 
<< pdiffusion >>
rect 33 193 34 194 
<< pdiffusion >>
rect 34 193 35 194 
<< pdiffusion >>
rect 35 193 36 194 
<< m1 >>
rect 37 193 38 194 
<< m2 >>
rect 38 193 39 194 
<< m1 >>
rect 44 193 45 194 
<< m1 >>
rect 46 193 47 194 
<< pdiffusion >>
rect 48 193 49 194 
<< pdiffusion >>
rect 49 193 50 194 
<< pdiffusion >>
rect 50 193 51 194 
<< pdiffusion >>
rect 51 193 52 194 
<< pdiffusion >>
rect 52 193 53 194 
<< pdiffusion >>
rect 53 193 54 194 
<< m1 >>
rect 56 193 57 194 
<< m1 >>
rect 58 193 59 194 
<< m1 >>
rect 62 193 63 194 
<< m1 >>
rect 64 193 65 194 
<< pdiffusion >>
rect 66 193 67 194 
<< pdiffusion >>
rect 67 193 68 194 
<< pdiffusion >>
rect 68 193 69 194 
<< pdiffusion >>
rect 69 193 70 194 
<< pdiffusion >>
rect 70 193 71 194 
<< pdiffusion >>
rect 71 193 72 194 
<< m2 >>
rect 79 193 80 194 
<< m1 >>
rect 80 193 81 194 
<< m1 >>
rect 82 193 83 194 
<< pdiffusion >>
rect 84 193 85 194 
<< pdiffusion >>
rect 85 193 86 194 
<< pdiffusion >>
rect 86 193 87 194 
<< pdiffusion >>
rect 87 193 88 194 
<< pdiffusion >>
rect 88 193 89 194 
<< pdiffusion >>
rect 89 193 90 194 
<< pdiffusion >>
rect 102 193 103 194 
<< pdiffusion >>
rect 103 193 104 194 
<< pdiffusion >>
rect 104 193 105 194 
<< pdiffusion >>
rect 105 193 106 194 
<< pdiffusion >>
rect 106 193 107 194 
<< pdiffusion >>
rect 107 193 108 194 
<< m1 >>
rect 118 193 119 194 
<< pdiffusion >>
rect 120 193 121 194 
<< pdiffusion >>
rect 121 193 122 194 
<< pdiffusion >>
rect 122 193 123 194 
<< pdiffusion >>
rect 123 193 124 194 
<< pdiffusion >>
rect 124 193 125 194 
<< pdiffusion >>
rect 125 193 126 194 
<< m1 >>
rect 127 193 128 194 
<< m2 >>
rect 127 193 128 194 
<< m2c >>
rect 127 193 128 194 
<< m1 >>
rect 127 193 128 194 
<< m2 >>
rect 127 193 128 194 
<< m1 >>
rect 130 193 131 194 
<< m2 >>
rect 130 193 131 194 
<< m2c >>
rect 130 193 131 194 
<< m1 >>
rect 130 193 131 194 
<< m2 >>
rect 130 193 131 194 
<< m1 >>
rect 132 193 133 194 
<< m2 >>
rect 132 193 133 194 
<< m2c >>
rect 132 193 133 194 
<< m1 >>
rect 132 193 133 194 
<< m2 >>
rect 132 193 133 194 
<< m2 >>
rect 135 193 136 194 
<< m1 >>
rect 136 193 137 194 
<< pdiffusion >>
rect 138 193 139 194 
<< pdiffusion >>
rect 139 193 140 194 
<< pdiffusion >>
rect 140 193 141 194 
<< pdiffusion >>
rect 141 193 142 194 
<< pdiffusion >>
rect 142 193 143 194 
<< pdiffusion >>
rect 143 193 144 194 
<< m1 >>
rect 145 193 146 194 
<< m2 >>
rect 146 193 147 194 
<< pdiffusion >>
rect 156 193 157 194 
<< pdiffusion >>
rect 157 193 158 194 
<< pdiffusion >>
rect 158 193 159 194 
<< pdiffusion >>
rect 159 193 160 194 
<< pdiffusion >>
rect 160 193 161 194 
<< pdiffusion >>
rect 161 193 162 194 
<< m1 >>
rect 163 193 164 194 
<< m1 >>
rect 165 193 166 194 
<< m1 >>
rect 170 193 171 194 
<< m1 >>
rect 172 193 173 194 
<< pdiffusion >>
rect 174 193 175 194 
<< pdiffusion >>
rect 175 193 176 194 
<< pdiffusion >>
rect 176 193 177 194 
<< pdiffusion >>
rect 177 193 178 194 
<< pdiffusion >>
rect 178 193 179 194 
<< pdiffusion >>
rect 179 193 180 194 
<< m1 >>
rect 181 193 182 194 
<< m2 >>
rect 181 193 182 194 
<< m1 >>
rect 183 193 184 194 
<< m1 >>
rect 188 193 189 194 
<< m1 >>
rect 190 193 191 194 
<< pdiffusion >>
rect 192 193 193 194 
<< pdiffusion >>
rect 193 193 194 194 
<< pdiffusion >>
rect 194 193 195 194 
<< pdiffusion >>
rect 195 193 196 194 
<< pdiffusion >>
rect 196 193 197 194 
<< pdiffusion >>
rect 197 193 198 194 
<< m1 >>
rect 199 193 200 194 
<< m2 >>
rect 199 193 200 194 
<< m1 >>
rect 201 193 202 194 
<< pdiffusion >>
rect 210 193 211 194 
<< pdiffusion >>
rect 211 193 212 194 
<< pdiffusion >>
rect 212 193 213 194 
<< pdiffusion >>
rect 213 193 214 194 
<< pdiffusion >>
rect 214 193 215 194 
<< pdiffusion >>
rect 215 193 216 194 
<< m1 >>
rect 218 193 219 194 
<< m2 >>
rect 225 193 226 194 
<< m1 >>
rect 226 193 227 194 
<< pdiffusion >>
rect 228 193 229 194 
<< pdiffusion >>
rect 229 193 230 194 
<< pdiffusion >>
rect 230 193 231 194 
<< pdiffusion >>
rect 231 193 232 194 
<< pdiffusion >>
rect 232 193 233 194 
<< pdiffusion >>
rect 233 193 234 194 
<< m1 >>
rect 235 193 236 194 
<< m1 >>
rect 237 193 238 194 
<< m1 >>
rect 241 193 242 194 
<< m1 >>
rect 243 193 244 194 
<< pdiffusion >>
rect 246 193 247 194 
<< pdiffusion >>
rect 247 193 248 194 
<< pdiffusion >>
rect 248 193 249 194 
<< pdiffusion >>
rect 249 193 250 194 
<< pdiffusion >>
rect 250 193 251 194 
<< pdiffusion >>
rect 251 193 252 194 
<< m1 >>
rect 253 193 254 194 
<< m1 >>
rect 255 193 256 194 
<< m1 >>
rect 260 193 261 194 
<< m1 >>
rect 262 193 263 194 
<< m2 >>
rect 262 193 263 194 
<< pdiffusion >>
rect 264 193 265 194 
<< pdiffusion >>
rect 265 193 266 194 
<< pdiffusion >>
rect 266 193 267 194 
<< pdiffusion >>
rect 267 193 268 194 
<< pdiffusion >>
rect 268 193 269 194 
<< pdiffusion >>
rect 269 193 270 194 
<< m2 >>
rect 271 193 272 194 
<< m1 >>
rect 272 193 273 194 
<< m1 >>
rect 274 193 275 194 
<< m2 >>
rect 275 193 276 194 
<< pdiffusion >>
rect 282 193 283 194 
<< pdiffusion >>
rect 283 193 284 194 
<< pdiffusion >>
rect 284 193 285 194 
<< pdiffusion >>
rect 285 193 286 194 
<< pdiffusion >>
rect 286 193 287 194 
<< pdiffusion >>
rect 287 193 288 194 
<< m1 >>
rect 289 193 290 194 
<< pdiffusion >>
rect 300 193 301 194 
<< pdiffusion >>
rect 301 193 302 194 
<< pdiffusion >>
rect 302 193 303 194 
<< pdiffusion >>
rect 303 193 304 194 
<< pdiffusion >>
rect 304 193 305 194 
<< pdiffusion >>
rect 305 193 306 194 
<< m1 >>
rect 307 193 308 194 
<< pdiffusion >>
rect 318 193 319 194 
<< pdiffusion >>
rect 319 193 320 194 
<< pdiffusion >>
rect 320 193 321 194 
<< pdiffusion >>
rect 321 193 322 194 
<< pdiffusion >>
rect 322 193 323 194 
<< pdiffusion >>
rect 323 193 324 194 
<< m1 >>
rect 325 193 326 194 
<< m1 >>
rect 327 193 328 194 
<< pdiffusion >>
rect 336 193 337 194 
<< pdiffusion >>
rect 337 193 338 194 
<< pdiffusion >>
rect 338 193 339 194 
<< pdiffusion >>
rect 339 193 340 194 
<< pdiffusion >>
rect 340 193 341 194 
<< pdiffusion >>
rect 341 193 342 194 
<< m1 >>
rect 343 193 344 194 
<< m2 >>
rect 343 193 344 194 
<< m1 >>
rect 345 193 346 194 
<< m1 >>
rect 10 194 11 195 
<< pdiffusion >>
rect 12 194 13 195 
<< pdiffusion >>
rect 13 194 14 195 
<< pdiffusion >>
rect 14 194 15 195 
<< pdiffusion >>
rect 15 194 16 195 
<< pdiffusion >>
rect 16 194 17 195 
<< pdiffusion >>
rect 17 194 18 195 
<< m1 >>
rect 19 194 20 195 
<< m1 >>
rect 21 194 22 195 
<< m2 >>
rect 27 194 28 195 
<< m1 >>
rect 28 194 29 195 
<< pdiffusion >>
rect 30 194 31 195 
<< pdiffusion >>
rect 31 194 32 195 
<< pdiffusion >>
rect 32 194 33 195 
<< pdiffusion >>
rect 33 194 34 195 
<< pdiffusion >>
rect 34 194 35 195 
<< pdiffusion >>
rect 35 194 36 195 
<< m1 >>
rect 37 194 38 195 
<< m2 >>
rect 38 194 39 195 
<< m1 >>
rect 44 194 45 195 
<< m1 >>
rect 46 194 47 195 
<< pdiffusion >>
rect 48 194 49 195 
<< pdiffusion >>
rect 49 194 50 195 
<< pdiffusion >>
rect 50 194 51 195 
<< pdiffusion >>
rect 51 194 52 195 
<< pdiffusion >>
rect 52 194 53 195 
<< pdiffusion >>
rect 53 194 54 195 
<< m1 >>
rect 56 194 57 195 
<< m1 >>
rect 58 194 59 195 
<< m1 >>
rect 62 194 63 195 
<< m1 >>
rect 64 194 65 195 
<< pdiffusion >>
rect 66 194 67 195 
<< pdiffusion >>
rect 67 194 68 195 
<< pdiffusion >>
rect 68 194 69 195 
<< pdiffusion >>
rect 69 194 70 195 
<< pdiffusion >>
rect 70 194 71 195 
<< pdiffusion >>
rect 71 194 72 195 
<< m2 >>
rect 79 194 80 195 
<< m1 >>
rect 80 194 81 195 
<< m1 >>
rect 82 194 83 195 
<< pdiffusion >>
rect 84 194 85 195 
<< pdiffusion >>
rect 85 194 86 195 
<< pdiffusion >>
rect 86 194 87 195 
<< pdiffusion >>
rect 87 194 88 195 
<< pdiffusion >>
rect 88 194 89 195 
<< pdiffusion >>
rect 89 194 90 195 
<< pdiffusion >>
rect 102 194 103 195 
<< pdiffusion >>
rect 103 194 104 195 
<< pdiffusion >>
rect 104 194 105 195 
<< pdiffusion >>
rect 105 194 106 195 
<< pdiffusion >>
rect 106 194 107 195 
<< pdiffusion >>
rect 107 194 108 195 
<< m1 >>
rect 118 194 119 195 
<< pdiffusion >>
rect 120 194 121 195 
<< pdiffusion >>
rect 121 194 122 195 
<< pdiffusion >>
rect 122 194 123 195 
<< pdiffusion >>
rect 123 194 124 195 
<< pdiffusion >>
rect 124 194 125 195 
<< pdiffusion >>
rect 125 194 126 195 
<< m1 >>
rect 127 194 128 195 
<< m1 >>
rect 130 194 131 195 
<< m1 >>
rect 132 194 133 195 
<< m2 >>
rect 135 194 136 195 
<< m1 >>
rect 136 194 137 195 
<< pdiffusion >>
rect 138 194 139 195 
<< pdiffusion >>
rect 139 194 140 195 
<< pdiffusion >>
rect 140 194 141 195 
<< pdiffusion >>
rect 141 194 142 195 
<< pdiffusion >>
rect 142 194 143 195 
<< pdiffusion >>
rect 143 194 144 195 
<< m1 >>
rect 145 194 146 195 
<< m2 >>
rect 146 194 147 195 
<< pdiffusion >>
rect 156 194 157 195 
<< pdiffusion >>
rect 157 194 158 195 
<< pdiffusion >>
rect 158 194 159 195 
<< pdiffusion >>
rect 159 194 160 195 
<< pdiffusion >>
rect 160 194 161 195 
<< pdiffusion >>
rect 161 194 162 195 
<< m1 >>
rect 163 194 164 195 
<< m1 >>
rect 165 194 166 195 
<< m1 >>
rect 170 194 171 195 
<< m1 >>
rect 172 194 173 195 
<< pdiffusion >>
rect 174 194 175 195 
<< pdiffusion >>
rect 175 194 176 195 
<< pdiffusion >>
rect 176 194 177 195 
<< pdiffusion >>
rect 177 194 178 195 
<< pdiffusion >>
rect 178 194 179 195 
<< pdiffusion >>
rect 179 194 180 195 
<< m1 >>
rect 181 194 182 195 
<< m2 >>
rect 181 194 182 195 
<< m1 >>
rect 183 194 184 195 
<< m1 >>
rect 188 194 189 195 
<< m1 >>
rect 190 194 191 195 
<< pdiffusion >>
rect 192 194 193 195 
<< pdiffusion >>
rect 193 194 194 195 
<< pdiffusion >>
rect 194 194 195 195 
<< pdiffusion >>
rect 195 194 196 195 
<< pdiffusion >>
rect 196 194 197 195 
<< pdiffusion >>
rect 197 194 198 195 
<< m1 >>
rect 199 194 200 195 
<< m2 >>
rect 199 194 200 195 
<< m1 >>
rect 201 194 202 195 
<< pdiffusion >>
rect 210 194 211 195 
<< pdiffusion >>
rect 211 194 212 195 
<< pdiffusion >>
rect 212 194 213 195 
<< pdiffusion >>
rect 213 194 214 195 
<< pdiffusion >>
rect 214 194 215 195 
<< pdiffusion >>
rect 215 194 216 195 
<< m1 >>
rect 218 194 219 195 
<< m2 >>
rect 225 194 226 195 
<< m1 >>
rect 226 194 227 195 
<< pdiffusion >>
rect 228 194 229 195 
<< pdiffusion >>
rect 229 194 230 195 
<< pdiffusion >>
rect 230 194 231 195 
<< pdiffusion >>
rect 231 194 232 195 
<< pdiffusion >>
rect 232 194 233 195 
<< pdiffusion >>
rect 233 194 234 195 
<< m1 >>
rect 235 194 236 195 
<< m1 >>
rect 237 194 238 195 
<< m1 >>
rect 241 194 242 195 
<< m1 >>
rect 243 194 244 195 
<< pdiffusion >>
rect 246 194 247 195 
<< pdiffusion >>
rect 247 194 248 195 
<< pdiffusion >>
rect 248 194 249 195 
<< pdiffusion >>
rect 249 194 250 195 
<< pdiffusion >>
rect 250 194 251 195 
<< pdiffusion >>
rect 251 194 252 195 
<< m1 >>
rect 253 194 254 195 
<< m1 >>
rect 255 194 256 195 
<< m1 >>
rect 260 194 261 195 
<< m1 >>
rect 262 194 263 195 
<< m2 >>
rect 262 194 263 195 
<< pdiffusion >>
rect 264 194 265 195 
<< pdiffusion >>
rect 265 194 266 195 
<< pdiffusion >>
rect 266 194 267 195 
<< pdiffusion >>
rect 267 194 268 195 
<< pdiffusion >>
rect 268 194 269 195 
<< pdiffusion >>
rect 269 194 270 195 
<< m2 >>
rect 271 194 272 195 
<< m1 >>
rect 272 194 273 195 
<< m1 >>
rect 274 194 275 195 
<< m2 >>
rect 275 194 276 195 
<< pdiffusion >>
rect 282 194 283 195 
<< pdiffusion >>
rect 283 194 284 195 
<< pdiffusion >>
rect 284 194 285 195 
<< pdiffusion >>
rect 285 194 286 195 
<< pdiffusion >>
rect 286 194 287 195 
<< pdiffusion >>
rect 287 194 288 195 
<< m1 >>
rect 289 194 290 195 
<< pdiffusion >>
rect 300 194 301 195 
<< pdiffusion >>
rect 301 194 302 195 
<< pdiffusion >>
rect 302 194 303 195 
<< pdiffusion >>
rect 303 194 304 195 
<< pdiffusion >>
rect 304 194 305 195 
<< pdiffusion >>
rect 305 194 306 195 
<< m1 >>
rect 307 194 308 195 
<< pdiffusion >>
rect 318 194 319 195 
<< pdiffusion >>
rect 319 194 320 195 
<< pdiffusion >>
rect 320 194 321 195 
<< pdiffusion >>
rect 321 194 322 195 
<< pdiffusion >>
rect 322 194 323 195 
<< pdiffusion >>
rect 323 194 324 195 
<< m1 >>
rect 325 194 326 195 
<< m1 >>
rect 327 194 328 195 
<< pdiffusion >>
rect 336 194 337 195 
<< pdiffusion >>
rect 337 194 338 195 
<< pdiffusion >>
rect 338 194 339 195 
<< pdiffusion >>
rect 339 194 340 195 
<< pdiffusion >>
rect 340 194 341 195 
<< pdiffusion >>
rect 341 194 342 195 
<< m1 >>
rect 343 194 344 195 
<< m2 >>
rect 343 194 344 195 
<< m1 >>
rect 345 194 346 195 
<< m1 >>
rect 10 195 11 196 
<< pdiffusion >>
rect 12 195 13 196 
<< pdiffusion >>
rect 13 195 14 196 
<< pdiffusion >>
rect 14 195 15 196 
<< pdiffusion >>
rect 15 195 16 196 
<< pdiffusion >>
rect 16 195 17 196 
<< pdiffusion >>
rect 17 195 18 196 
<< m1 >>
rect 19 195 20 196 
<< m1 >>
rect 21 195 22 196 
<< m2 >>
rect 27 195 28 196 
<< m1 >>
rect 28 195 29 196 
<< pdiffusion >>
rect 30 195 31 196 
<< pdiffusion >>
rect 31 195 32 196 
<< pdiffusion >>
rect 32 195 33 196 
<< pdiffusion >>
rect 33 195 34 196 
<< pdiffusion >>
rect 34 195 35 196 
<< pdiffusion >>
rect 35 195 36 196 
<< m1 >>
rect 37 195 38 196 
<< m2 >>
rect 38 195 39 196 
<< m1 >>
rect 44 195 45 196 
<< m1 >>
rect 46 195 47 196 
<< pdiffusion >>
rect 48 195 49 196 
<< pdiffusion >>
rect 49 195 50 196 
<< pdiffusion >>
rect 50 195 51 196 
<< pdiffusion >>
rect 51 195 52 196 
<< pdiffusion >>
rect 52 195 53 196 
<< pdiffusion >>
rect 53 195 54 196 
<< m1 >>
rect 56 195 57 196 
<< m1 >>
rect 58 195 59 196 
<< m1 >>
rect 62 195 63 196 
<< m1 >>
rect 64 195 65 196 
<< pdiffusion >>
rect 66 195 67 196 
<< pdiffusion >>
rect 67 195 68 196 
<< pdiffusion >>
rect 68 195 69 196 
<< pdiffusion >>
rect 69 195 70 196 
<< pdiffusion >>
rect 70 195 71 196 
<< pdiffusion >>
rect 71 195 72 196 
<< m2 >>
rect 79 195 80 196 
<< m1 >>
rect 80 195 81 196 
<< m1 >>
rect 82 195 83 196 
<< pdiffusion >>
rect 84 195 85 196 
<< pdiffusion >>
rect 85 195 86 196 
<< pdiffusion >>
rect 86 195 87 196 
<< pdiffusion >>
rect 87 195 88 196 
<< pdiffusion >>
rect 88 195 89 196 
<< pdiffusion >>
rect 89 195 90 196 
<< pdiffusion >>
rect 102 195 103 196 
<< pdiffusion >>
rect 103 195 104 196 
<< pdiffusion >>
rect 104 195 105 196 
<< pdiffusion >>
rect 105 195 106 196 
<< pdiffusion >>
rect 106 195 107 196 
<< pdiffusion >>
rect 107 195 108 196 
<< m1 >>
rect 118 195 119 196 
<< pdiffusion >>
rect 120 195 121 196 
<< pdiffusion >>
rect 121 195 122 196 
<< pdiffusion >>
rect 122 195 123 196 
<< pdiffusion >>
rect 123 195 124 196 
<< pdiffusion >>
rect 124 195 125 196 
<< pdiffusion >>
rect 125 195 126 196 
<< m1 >>
rect 127 195 128 196 
<< m1 >>
rect 128 195 129 196 
<< m2 >>
rect 128 195 129 196 
<< m2c >>
rect 128 195 129 196 
<< m1 >>
rect 128 195 129 196 
<< m2 >>
rect 128 195 129 196 
<< m2 >>
rect 129 195 130 196 
<< m1 >>
rect 130 195 131 196 
<< m2 >>
rect 130 195 131 196 
<< m2 >>
rect 131 195 132 196 
<< m1 >>
rect 132 195 133 196 
<< m2 >>
rect 132 195 133 196 
<< m2 >>
rect 133 195 134 196 
<< m1 >>
rect 134 195 135 196 
<< m2 >>
rect 134 195 135 196 
<< m2c >>
rect 134 195 135 196 
<< m1 >>
rect 134 195 135 196 
<< m2 >>
rect 134 195 135 196 
<< m2 >>
rect 135 195 136 196 
<< m1 >>
rect 136 195 137 196 
<< pdiffusion >>
rect 138 195 139 196 
<< pdiffusion >>
rect 139 195 140 196 
<< pdiffusion >>
rect 140 195 141 196 
<< pdiffusion >>
rect 141 195 142 196 
<< pdiffusion >>
rect 142 195 143 196 
<< pdiffusion >>
rect 143 195 144 196 
<< m1 >>
rect 145 195 146 196 
<< m2 >>
rect 146 195 147 196 
<< pdiffusion >>
rect 156 195 157 196 
<< pdiffusion >>
rect 157 195 158 196 
<< pdiffusion >>
rect 158 195 159 196 
<< pdiffusion >>
rect 159 195 160 196 
<< pdiffusion >>
rect 160 195 161 196 
<< pdiffusion >>
rect 161 195 162 196 
<< m1 >>
rect 163 195 164 196 
<< m1 >>
rect 165 195 166 196 
<< m1 >>
rect 170 195 171 196 
<< m1 >>
rect 172 195 173 196 
<< pdiffusion >>
rect 174 195 175 196 
<< pdiffusion >>
rect 175 195 176 196 
<< pdiffusion >>
rect 176 195 177 196 
<< pdiffusion >>
rect 177 195 178 196 
<< pdiffusion >>
rect 178 195 179 196 
<< pdiffusion >>
rect 179 195 180 196 
<< m1 >>
rect 181 195 182 196 
<< m2 >>
rect 181 195 182 196 
<< m1 >>
rect 183 195 184 196 
<< m1 >>
rect 188 195 189 196 
<< m1 >>
rect 190 195 191 196 
<< pdiffusion >>
rect 192 195 193 196 
<< pdiffusion >>
rect 193 195 194 196 
<< pdiffusion >>
rect 194 195 195 196 
<< pdiffusion >>
rect 195 195 196 196 
<< pdiffusion >>
rect 196 195 197 196 
<< pdiffusion >>
rect 197 195 198 196 
<< m1 >>
rect 199 195 200 196 
<< m2 >>
rect 199 195 200 196 
<< m1 >>
rect 201 195 202 196 
<< pdiffusion >>
rect 210 195 211 196 
<< pdiffusion >>
rect 211 195 212 196 
<< pdiffusion >>
rect 212 195 213 196 
<< pdiffusion >>
rect 213 195 214 196 
<< pdiffusion >>
rect 214 195 215 196 
<< pdiffusion >>
rect 215 195 216 196 
<< m1 >>
rect 218 195 219 196 
<< m2 >>
rect 225 195 226 196 
<< m1 >>
rect 226 195 227 196 
<< pdiffusion >>
rect 228 195 229 196 
<< pdiffusion >>
rect 229 195 230 196 
<< pdiffusion >>
rect 230 195 231 196 
<< pdiffusion >>
rect 231 195 232 196 
<< pdiffusion >>
rect 232 195 233 196 
<< pdiffusion >>
rect 233 195 234 196 
<< m1 >>
rect 235 195 236 196 
<< m1 >>
rect 237 195 238 196 
<< m1 >>
rect 241 195 242 196 
<< m1 >>
rect 243 195 244 196 
<< pdiffusion >>
rect 246 195 247 196 
<< pdiffusion >>
rect 247 195 248 196 
<< pdiffusion >>
rect 248 195 249 196 
<< pdiffusion >>
rect 249 195 250 196 
<< pdiffusion >>
rect 250 195 251 196 
<< pdiffusion >>
rect 251 195 252 196 
<< m1 >>
rect 253 195 254 196 
<< m1 >>
rect 255 195 256 196 
<< m1 >>
rect 260 195 261 196 
<< m1 >>
rect 262 195 263 196 
<< m2 >>
rect 262 195 263 196 
<< pdiffusion >>
rect 264 195 265 196 
<< pdiffusion >>
rect 265 195 266 196 
<< pdiffusion >>
rect 266 195 267 196 
<< pdiffusion >>
rect 267 195 268 196 
<< pdiffusion >>
rect 268 195 269 196 
<< pdiffusion >>
rect 269 195 270 196 
<< m2 >>
rect 271 195 272 196 
<< m1 >>
rect 272 195 273 196 
<< m1 >>
rect 274 195 275 196 
<< m2 >>
rect 275 195 276 196 
<< pdiffusion >>
rect 282 195 283 196 
<< pdiffusion >>
rect 283 195 284 196 
<< pdiffusion >>
rect 284 195 285 196 
<< pdiffusion >>
rect 285 195 286 196 
<< pdiffusion >>
rect 286 195 287 196 
<< pdiffusion >>
rect 287 195 288 196 
<< m1 >>
rect 289 195 290 196 
<< pdiffusion >>
rect 300 195 301 196 
<< pdiffusion >>
rect 301 195 302 196 
<< pdiffusion >>
rect 302 195 303 196 
<< pdiffusion >>
rect 303 195 304 196 
<< pdiffusion >>
rect 304 195 305 196 
<< pdiffusion >>
rect 305 195 306 196 
<< m1 >>
rect 307 195 308 196 
<< pdiffusion >>
rect 318 195 319 196 
<< pdiffusion >>
rect 319 195 320 196 
<< pdiffusion >>
rect 320 195 321 196 
<< pdiffusion >>
rect 321 195 322 196 
<< pdiffusion >>
rect 322 195 323 196 
<< pdiffusion >>
rect 323 195 324 196 
<< m1 >>
rect 325 195 326 196 
<< m1 >>
rect 327 195 328 196 
<< pdiffusion >>
rect 336 195 337 196 
<< pdiffusion >>
rect 337 195 338 196 
<< pdiffusion >>
rect 338 195 339 196 
<< pdiffusion >>
rect 339 195 340 196 
<< pdiffusion >>
rect 340 195 341 196 
<< pdiffusion >>
rect 341 195 342 196 
<< m1 >>
rect 343 195 344 196 
<< m2 >>
rect 343 195 344 196 
<< m1 >>
rect 345 195 346 196 
<< m1 >>
rect 10 196 11 197 
<< pdiffusion >>
rect 12 196 13 197 
<< pdiffusion >>
rect 13 196 14 197 
<< pdiffusion >>
rect 14 196 15 197 
<< pdiffusion >>
rect 15 196 16 197 
<< pdiffusion >>
rect 16 196 17 197 
<< pdiffusion >>
rect 17 196 18 197 
<< m1 >>
rect 19 196 20 197 
<< m1 >>
rect 21 196 22 197 
<< m2 >>
rect 27 196 28 197 
<< m1 >>
rect 28 196 29 197 
<< pdiffusion >>
rect 30 196 31 197 
<< pdiffusion >>
rect 31 196 32 197 
<< pdiffusion >>
rect 32 196 33 197 
<< pdiffusion >>
rect 33 196 34 197 
<< pdiffusion >>
rect 34 196 35 197 
<< pdiffusion >>
rect 35 196 36 197 
<< m1 >>
rect 37 196 38 197 
<< m2 >>
rect 38 196 39 197 
<< m1 >>
rect 44 196 45 197 
<< m1 >>
rect 46 196 47 197 
<< pdiffusion >>
rect 48 196 49 197 
<< pdiffusion >>
rect 49 196 50 197 
<< pdiffusion >>
rect 50 196 51 197 
<< pdiffusion >>
rect 51 196 52 197 
<< pdiffusion >>
rect 52 196 53 197 
<< pdiffusion >>
rect 53 196 54 197 
<< m1 >>
rect 56 196 57 197 
<< m1 >>
rect 58 196 59 197 
<< m1 >>
rect 62 196 63 197 
<< m1 >>
rect 64 196 65 197 
<< pdiffusion >>
rect 66 196 67 197 
<< pdiffusion >>
rect 67 196 68 197 
<< pdiffusion >>
rect 68 196 69 197 
<< pdiffusion >>
rect 69 196 70 197 
<< pdiffusion >>
rect 70 196 71 197 
<< pdiffusion >>
rect 71 196 72 197 
<< m2 >>
rect 79 196 80 197 
<< m1 >>
rect 80 196 81 197 
<< m1 >>
rect 82 196 83 197 
<< pdiffusion >>
rect 84 196 85 197 
<< pdiffusion >>
rect 85 196 86 197 
<< pdiffusion >>
rect 86 196 87 197 
<< pdiffusion >>
rect 87 196 88 197 
<< pdiffusion >>
rect 88 196 89 197 
<< pdiffusion >>
rect 89 196 90 197 
<< pdiffusion >>
rect 102 196 103 197 
<< pdiffusion >>
rect 103 196 104 197 
<< pdiffusion >>
rect 104 196 105 197 
<< pdiffusion >>
rect 105 196 106 197 
<< pdiffusion >>
rect 106 196 107 197 
<< pdiffusion >>
rect 107 196 108 197 
<< m1 >>
rect 118 196 119 197 
<< pdiffusion >>
rect 120 196 121 197 
<< pdiffusion >>
rect 121 196 122 197 
<< pdiffusion >>
rect 122 196 123 197 
<< pdiffusion >>
rect 123 196 124 197 
<< pdiffusion >>
rect 124 196 125 197 
<< pdiffusion >>
rect 125 196 126 197 
<< m1 >>
rect 130 196 131 197 
<< m1 >>
rect 132 196 133 197 
<< m1 >>
rect 134 196 135 197 
<< m2 >>
rect 135 196 136 197 
<< m1 >>
rect 136 196 137 197 
<< pdiffusion >>
rect 138 196 139 197 
<< pdiffusion >>
rect 139 196 140 197 
<< pdiffusion >>
rect 140 196 141 197 
<< pdiffusion >>
rect 141 196 142 197 
<< pdiffusion >>
rect 142 196 143 197 
<< pdiffusion >>
rect 143 196 144 197 
<< m1 >>
rect 145 196 146 197 
<< m2 >>
rect 146 196 147 197 
<< pdiffusion >>
rect 156 196 157 197 
<< pdiffusion >>
rect 157 196 158 197 
<< pdiffusion >>
rect 158 196 159 197 
<< pdiffusion >>
rect 159 196 160 197 
<< pdiffusion >>
rect 160 196 161 197 
<< pdiffusion >>
rect 161 196 162 197 
<< m1 >>
rect 163 196 164 197 
<< m1 >>
rect 165 196 166 197 
<< m1 >>
rect 170 196 171 197 
<< m1 >>
rect 172 196 173 197 
<< pdiffusion >>
rect 174 196 175 197 
<< pdiffusion >>
rect 175 196 176 197 
<< pdiffusion >>
rect 176 196 177 197 
<< pdiffusion >>
rect 177 196 178 197 
<< pdiffusion >>
rect 178 196 179 197 
<< pdiffusion >>
rect 179 196 180 197 
<< m1 >>
rect 181 196 182 197 
<< m2 >>
rect 181 196 182 197 
<< m1 >>
rect 183 196 184 197 
<< m1 >>
rect 188 196 189 197 
<< m1 >>
rect 190 196 191 197 
<< pdiffusion >>
rect 192 196 193 197 
<< pdiffusion >>
rect 193 196 194 197 
<< pdiffusion >>
rect 194 196 195 197 
<< pdiffusion >>
rect 195 196 196 197 
<< pdiffusion >>
rect 196 196 197 197 
<< pdiffusion >>
rect 197 196 198 197 
<< m1 >>
rect 199 196 200 197 
<< m2 >>
rect 199 196 200 197 
<< m1 >>
rect 201 196 202 197 
<< pdiffusion >>
rect 210 196 211 197 
<< pdiffusion >>
rect 211 196 212 197 
<< pdiffusion >>
rect 212 196 213 197 
<< pdiffusion >>
rect 213 196 214 197 
<< pdiffusion >>
rect 214 196 215 197 
<< pdiffusion >>
rect 215 196 216 197 
<< m1 >>
rect 218 196 219 197 
<< m2 >>
rect 225 196 226 197 
<< m1 >>
rect 226 196 227 197 
<< pdiffusion >>
rect 228 196 229 197 
<< pdiffusion >>
rect 229 196 230 197 
<< pdiffusion >>
rect 230 196 231 197 
<< pdiffusion >>
rect 231 196 232 197 
<< pdiffusion >>
rect 232 196 233 197 
<< pdiffusion >>
rect 233 196 234 197 
<< m1 >>
rect 235 196 236 197 
<< m1 >>
rect 237 196 238 197 
<< m1 >>
rect 241 196 242 197 
<< m1 >>
rect 243 196 244 197 
<< pdiffusion >>
rect 246 196 247 197 
<< pdiffusion >>
rect 247 196 248 197 
<< pdiffusion >>
rect 248 196 249 197 
<< pdiffusion >>
rect 249 196 250 197 
<< pdiffusion >>
rect 250 196 251 197 
<< pdiffusion >>
rect 251 196 252 197 
<< m1 >>
rect 253 196 254 197 
<< m1 >>
rect 255 196 256 197 
<< m1 >>
rect 260 196 261 197 
<< m1 >>
rect 262 196 263 197 
<< m2 >>
rect 262 196 263 197 
<< pdiffusion >>
rect 264 196 265 197 
<< pdiffusion >>
rect 265 196 266 197 
<< pdiffusion >>
rect 266 196 267 197 
<< pdiffusion >>
rect 267 196 268 197 
<< pdiffusion >>
rect 268 196 269 197 
<< pdiffusion >>
rect 269 196 270 197 
<< m2 >>
rect 271 196 272 197 
<< m1 >>
rect 272 196 273 197 
<< m1 >>
rect 274 196 275 197 
<< m2 >>
rect 275 196 276 197 
<< pdiffusion >>
rect 282 196 283 197 
<< pdiffusion >>
rect 283 196 284 197 
<< pdiffusion >>
rect 284 196 285 197 
<< pdiffusion >>
rect 285 196 286 197 
<< pdiffusion >>
rect 286 196 287 197 
<< pdiffusion >>
rect 287 196 288 197 
<< m1 >>
rect 289 196 290 197 
<< pdiffusion >>
rect 300 196 301 197 
<< pdiffusion >>
rect 301 196 302 197 
<< pdiffusion >>
rect 302 196 303 197 
<< pdiffusion >>
rect 303 196 304 197 
<< pdiffusion >>
rect 304 196 305 197 
<< pdiffusion >>
rect 305 196 306 197 
<< m1 >>
rect 307 196 308 197 
<< pdiffusion >>
rect 318 196 319 197 
<< pdiffusion >>
rect 319 196 320 197 
<< pdiffusion >>
rect 320 196 321 197 
<< pdiffusion >>
rect 321 196 322 197 
<< pdiffusion >>
rect 322 196 323 197 
<< pdiffusion >>
rect 323 196 324 197 
<< m1 >>
rect 325 196 326 197 
<< m1 >>
rect 327 196 328 197 
<< pdiffusion >>
rect 336 196 337 197 
<< pdiffusion >>
rect 337 196 338 197 
<< pdiffusion >>
rect 338 196 339 197 
<< pdiffusion >>
rect 339 196 340 197 
<< pdiffusion >>
rect 340 196 341 197 
<< pdiffusion >>
rect 341 196 342 197 
<< m1 >>
rect 343 196 344 197 
<< m2 >>
rect 343 196 344 197 
<< m1 >>
rect 345 196 346 197 
<< m1 >>
rect 10 197 11 198 
<< pdiffusion >>
rect 12 197 13 198 
<< pdiffusion >>
rect 13 197 14 198 
<< pdiffusion >>
rect 14 197 15 198 
<< pdiffusion >>
rect 15 197 16 198 
<< pdiffusion >>
rect 16 197 17 198 
<< pdiffusion >>
rect 17 197 18 198 
<< m1 >>
rect 19 197 20 198 
<< m1 >>
rect 21 197 22 198 
<< m2 >>
rect 27 197 28 198 
<< m1 >>
rect 28 197 29 198 
<< pdiffusion >>
rect 30 197 31 198 
<< pdiffusion >>
rect 31 197 32 198 
<< pdiffusion >>
rect 32 197 33 198 
<< pdiffusion >>
rect 33 197 34 198 
<< pdiffusion >>
rect 34 197 35 198 
<< pdiffusion >>
rect 35 197 36 198 
<< m1 >>
rect 37 197 38 198 
<< m2 >>
rect 38 197 39 198 
<< m1 >>
rect 44 197 45 198 
<< m1 >>
rect 46 197 47 198 
<< pdiffusion >>
rect 48 197 49 198 
<< pdiffusion >>
rect 49 197 50 198 
<< pdiffusion >>
rect 50 197 51 198 
<< pdiffusion >>
rect 51 197 52 198 
<< pdiffusion >>
rect 52 197 53 198 
<< pdiffusion >>
rect 53 197 54 198 
<< m1 >>
rect 56 197 57 198 
<< m1 >>
rect 58 197 59 198 
<< m1 >>
rect 62 197 63 198 
<< m1 >>
rect 64 197 65 198 
<< pdiffusion >>
rect 66 197 67 198 
<< pdiffusion >>
rect 67 197 68 198 
<< pdiffusion >>
rect 68 197 69 198 
<< pdiffusion >>
rect 69 197 70 198 
<< pdiffusion >>
rect 70 197 71 198 
<< pdiffusion >>
rect 71 197 72 198 
<< m2 >>
rect 79 197 80 198 
<< m1 >>
rect 80 197 81 198 
<< m1 >>
rect 82 197 83 198 
<< pdiffusion >>
rect 84 197 85 198 
<< pdiffusion >>
rect 85 197 86 198 
<< pdiffusion >>
rect 86 197 87 198 
<< pdiffusion >>
rect 87 197 88 198 
<< pdiffusion >>
rect 88 197 89 198 
<< pdiffusion >>
rect 89 197 90 198 
<< pdiffusion >>
rect 102 197 103 198 
<< pdiffusion >>
rect 103 197 104 198 
<< pdiffusion >>
rect 104 197 105 198 
<< pdiffusion >>
rect 105 197 106 198 
<< m1 >>
rect 106 197 107 198 
<< pdiffusion >>
rect 106 197 107 198 
<< pdiffusion >>
rect 107 197 108 198 
<< m1 >>
rect 118 197 119 198 
<< pdiffusion >>
rect 120 197 121 198 
<< pdiffusion >>
rect 121 197 122 198 
<< pdiffusion >>
rect 122 197 123 198 
<< pdiffusion >>
rect 123 197 124 198 
<< pdiffusion >>
rect 124 197 125 198 
<< pdiffusion >>
rect 125 197 126 198 
<< m1 >>
rect 130 197 131 198 
<< m1 >>
rect 132 197 133 198 
<< m1 >>
rect 134 197 135 198 
<< m2 >>
rect 135 197 136 198 
<< m1 >>
rect 136 197 137 198 
<< pdiffusion >>
rect 138 197 139 198 
<< pdiffusion >>
rect 139 197 140 198 
<< pdiffusion >>
rect 140 197 141 198 
<< pdiffusion >>
rect 141 197 142 198 
<< pdiffusion >>
rect 142 197 143 198 
<< pdiffusion >>
rect 143 197 144 198 
<< m1 >>
rect 145 197 146 198 
<< m2 >>
rect 146 197 147 198 
<< pdiffusion >>
rect 156 197 157 198 
<< pdiffusion >>
rect 157 197 158 198 
<< pdiffusion >>
rect 158 197 159 198 
<< pdiffusion >>
rect 159 197 160 198 
<< m1 >>
rect 160 197 161 198 
<< pdiffusion >>
rect 160 197 161 198 
<< pdiffusion >>
rect 161 197 162 198 
<< m1 >>
rect 163 197 164 198 
<< m1 >>
rect 165 197 166 198 
<< m1 >>
rect 170 197 171 198 
<< m1 >>
rect 172 197 173 198 
<< pdiffusion >>
rect 174 197 175 198 
<< pdiffusion >>
rect 175 197 176 198 
<< pdiffusion >>
rect 176 197 177 198 
<< pdiffusion >>
rect 177 197 178 198 
<< pdiffusion >>
rect 178 197 179 198 
<< pdiffusion >>
rect 179 197 180 198 
<< m1 >>
rect 181 197 182 198 
<< m2 >>
rect 181 197 182 198 
<< m1 >>
rect 183 197 184 198 
<< m1 >>
rect 188 197 189 198 
<< m1 >>
rect 190 197 191 198 
<< pdiffusion >>
rect 192 197 193 198 
<< m1 >>
rect 193 197 194 198 
<< pdiffusion >>
rect 193 197 194 198 
<< pdiffusion >>
rect 194 197 195 198 
<< pdiffusion >>
rect 195 197 196 198 
<< pdiffusion >>
rect 196 197 197 198 
<< pdiffusion >>
rect 197 197 198 198 
<< m1 >>
rect 199 197 200 198 
<< m2 >>
rect 199 197 200 198 
<< m1 >>
rect 201 197 202 198 
<< pdiffusion >>
rect 210 197 211 198 
<< pdiffusion >>
rect 211 197 212 198 
<< pdiffusion >>
rect 212 197 213 198 
<< pdiffusion >>
rect 213 197 214 198 
<< pdiffusion >>
rect 214 197 215 198 
<< pdiffusion >>
rect 215 197 216 198 
<< m1 >>
rect 218 197 219 198 
<< m2 >>
rect 225 197 226 198 
<< m1 >>
rect 226 197 227 198 
<< pdiffusion >>
rect 228 197 229 198 
<< pdiffusion >>
rect 229 197 230 198 
<< pdiffusion >>
rect 230 197 231 198 
<< pdiffusion >>
rect 231 197 232 198 
<< m1 >>
rect 232 197 233 198 
<< pdiffusion >>
rect 232 197 233 198 
<< pdiffusion >>
rect 233 197 234 198 
<< m1 >>
rect 235 197 236 198 
<< m1 >>
rect 237 197 238 198 
<< m1 >>
rect 241 197 242 198 
<< m1 >>
rect 243 197 244 198 
<< pdiffusion >>
rect 246 197 247 198 
<< pdiffusion >>
rect 247 197 248 198 
<< pdiffusion >>
rect 248 197 249 198 
<< pdiffusion >>
rect 249 197 250 198 
<< m1 >>
rect 250 197 251 198 
<< pdiffusion >>
rect 250 197 251 198 
<< pdiffusion >>
rect 251 197 252 198 
<< m1 >>
rect 253 197 254 198 
<< m1 >>
rect 255 197 256 198 
<< m1 >>
rect 260 197 261 198 
<< m1 >>
rect 262 197 263 198 
<< m2 >>
rect 262 197 263 198 
<< pdiffusion >>
rect 264 197 265 198 
<< m1 >>
rect 265 197 266 198 
<< pdiffusion >>
rect 265 197 266 198 
<< pdiffusion >>
rect 266 197 267 198 
<< pdiffusion >>
rect 267 197 268 198 
<< m1 >>
rect 268 197 269 198 
<< pdiffusion >>
rect 268 197 269 198 
<< pdiffusion >>
rect 269 197 270 198 
<< m2 >>
rect 271 197 272 198 
<< m1 >>
rect 272 197 273 198 
<< m1 >>
rect 274 197 275 198 
<< m2 >>
rect 275 197 276 198 
<< pdiffusion >>
rect 282 197 283 198 
<< pdiffusion >>
rect 283 197 284 198 
<< pdiffusion >>
rect 284 197 285 198 
<< pdiffusion >>
rect 285 197 286 198 
<< pdiffusion >>
rect 286 197 287 198 
<< pdiffusion >>
rect 287 197 288 198 
<< m1 >>
rect 289 197 290 198 
<< pdiffusion >>
rect 300 197 301 198 
<< pdiffusion >>
rect 301 197 302 198 
<< pdiffusion >>
rect 302 197 303 198 
<< pdiffusion >>
rect 303 197 304 198 
<< pdiffusion >>
rect 304 197 305 198 
<< pdiffusion >>
rect 305 197 306 198 
<< m1 >>
rect 307 197 308 198 
<< pdiffusion >>
rect 318 197 319 198 
<< pdiffusion >>
rect 319 197 320 198 
<< pdiffusion >>
rect 320 197 321 198 
<< pdiffusion >>
rect 321 197 322 198 
<< pdiffusion >>
rect 322 197 323 198 
<< pdiffusion >>
rect 323 197 324 198 
<< m1 >>
rect 325 197 326 198 
<< m1 >>
rect 327 197 328 198 
<< pdiffusion >>
rect 336 197 337 198 
<< pdiffusion >>
rect 337 197 338 198 
<< pdiffusion >>
rect 338 197 339 198 
<< pdiffusion >>
rect 339 197 340 198 
<< m1 >>
rect 340 197 341 198 
<< pdiffusion >>
rect 340 197 341 198 
<< pdiffusion >>
rect 341 197 342 198 
<< m1 >>
rect 343 197 344 198 
<< m2 >>
rect 343 197 344 198 
<< m1 >>
rect 345 197 346 198 
<< m1 >>
rect 10 198 11 199 
<< m1 >>
rect 19 198 20 199 
<< m1 >>
rect 21 198 22 199 
<< m2 >>
rect 27 198 28 199 
<< m1 >>
rect 28 198 29 199 
<< m1 >>
rect 37 198 38 199 
<< m2 >>
rect 38 198 39 199 
<< m1 >>
rect 44 198 45 199 
<< m1 >>
rect 46 198 47 199 
<< m1 >>
rect 56 198 57 199 
<< m1 >>
rect 58 198 59 199 
<< m1 >>
rect 62 198 63 199 
<< m1 >>
rect 64 198 65 199 
<< m2 >>
rect 79 198 80 199 
<< m1 >>
rect 80 198 81 199 
<< m1 >>
rect 82 198 83 199 
<< m1 >>
rect 106 198 107 199 
<< m1 >>
rect 118 198 119 199 
<< m1 >>
rect 130 198 131 199 
<< m1 >>
rect 132 198 133 199 
<< m1 >>
rect 134 198 135 199 
<< m2 >>
rect 135 198 136 199 
<< m1 >>
rect 136 198 137 199 
<< m1 >>
rect 145 198 146 199 
<< m2 >>
rect 146 198 147 199 
<< m1 >>
rect 160 198 161 199 
<< m1 >>
rect 163 198 164 199 
<< m1 >>
rect 165 198 166 199 
<< m1 >>
rect 170 198 171 199 
<< m1 >>
rect 172 198 173 199 
<< m1 >>
rect 181 198 182 199 
<< m2 >>
rect 181 198 182 199 
<< m1 >>
rect 183 198 184 199 
<< m1 >>
rect 188 198 189 199 
<< m1 >>
rect 190 198 191 199 
<< m1 >>
rect 193 198 194 199 
<< m1 >>
rect 199 198 200 199 
<< m2 >>
rect 199 198 200 199 
<< m1 >>
rect 201 198 202 199 
<< m1 >>
rect 218 198 219 199 
<< m2 >>
rect 225 198 226 199 
<< m1 >>
rect 226 198 227 199 
<< m1 >>
rect 232 198 233 199 
<< m1 >>
rect 235 198 236 199 
<< m1 >>
rect 237 198 238 199 
<< m1 >>
rect 241 198 242 199 
<< m1 >>
rect 243 198 244 199 
<< m1 >>
rect 250 198 251 199 
<< m1 >>
rect 253 198 254 199 
<< m1 >>
rect 255 198 256 199 
<< m1 >>
rect 260 198 261 199 
<< m1 >>
rect 262 198 263 199 
<< m2 >>
rect 262 198 263 199 
<< m1 >>
rect 265 198 266 199 
<< m1 >>
rect 268 198 269 199 
<< m2 >>
rect 271 198 272 199 
<< m1 >>
rect 272 198 273 199 
<< m1 >>
rect 274 198 275 199 
<< m2 >>
rect 275 198 276 199 
<< m1 >>
rect 289 198 290 199 
<< m1 >>
rect 307 198 308 199 
<< m1 >>
rect 325 198 326 199 
<< m1 >>
rect 327 198 328 199 
<< m1 >>
rect 340 198 341 199 
<< m1 >>
rect 343 198 344 199 
<< m2 >>
rect 343 198 344 199 
<< m1 >>
rect 345 198 346 199 
<< m1 >>
rect 10 199 11 200 
<< m1 >>
rect 19 199 20 200 
<< m1 >>
rect 21 199 22 200 
<< m2 >>
rect 27 199 28 200 
<< m1 >>
rect 28 199 29 200 
<< m1 >>
rect 37 199 38 200 
<< m2 >>
rect 38 199 39 200 
<< m1 >>
rect 44 199 45 200 
<< m1 >>
rect 46 199 47 200 
<< m1 >>
rect 56 199 57 200 
<< m1 >>
rect 58 199 59 200 
<< m1 >>
rect 62 199 63 200 
<< m1 >>
rect 64 199 65 200 
<< m2 >>
rect 79 199 80 200 
<< m1 >>
rect 80 199 81 200 
<< m1 >>
rect 82 199 83 200 
<< m1 >>
rect 106 199 107 200 
<< m1 >>
rect 118 199 119 200 
<< m1 >>
rect 130 199 131 200 
<< m1 >>
rect 132 199 133 200 
<< m1 >>
rect 134 199 135 200 
<< m2 >>
rect 135 199 136 200 
<< m1 >>
rect 136 199 137 200 
<< m2 >>
rect 136 199 137 200 
<< m2 >>
rect 137 199 138 200 
<< m1 >>
rect 138 199 139 200 
<< m2 >>
rect 138 199 139 200 
<< m2c >>
rect 138 199 139 200 
<< m1 >>
rect 138 199 139 200 
<< m2 >>
rect 138 199 139 200 
<< m1 >>
rect 145 199 146 200 
<< m2 >>
rect 146 199 147 200 
<< m1 >>
rect 160 199 161 200 
<< m1 >>
rect 163 199 164 200 
<< m1 >>
rect 165 199 166 200 
<< m1 >>
rect 170 199 171 200 
<< m1 >>
rect 172 199 173 200 
<< m1 >>
rect 179 199 180 200 
<< m2 >>
rect 179 199 180 200 
<< m2c >>
rect 179 199 180 200 
<< m1 >>
rect 179 199 180 200 
<< m2 >>
rect 179 199 180 200 
<< m2 >>
rect 180 199 181 200 
<< m1 >>
rect 181 199 182 200 
<< m2 >>
rect 181 199 182 200 
<< m1 >>
rect 183 199 184 200 
<< m1 >>
rect 188 199 189 200 
<< m1 >>
rect 190 199 191 200 
<< m1 >>
rect 193 199 194 200 
<< m1 >>
rect 197 199 198 200 
<< m2 >>
rect 197 199 198 200 
<< m2c >>
rect 197 199 198 200 
<< m1 >>
rect 197 199 198 200 
<< m2 >>
rect 197 199 198 200 
<< m2 >>
rect 198 199 199 200 
<< m1 >>
rect 199 199 200 200 
<< m2 >>
rect 199 199 200 200 
<< m1 >>
rect 201 199 202 200 
<< m1 >>
rect 218 199 219 200 
<< m2 >>
rect 225 199 226 200 
<< m1 >>
rect 226 199 227 200 
<< m1 >>
rect 232 199 233 200 
<< m1 >>
rect 235 199 236 200 
<< m1 >>
rect 237 199 238 200 
<< m1 >>
rect 241 199 242 200 
<< m1 >>
rect 243 199 244 200 
<< m1 >>
rect 250 199 251 200 
<< m1 >>
rect 251 199 252 200 
<< m1 >>
rect 252 199 253 200 
<< m1 >>
rect 253 199 254 200 
<< m1 >>
rect 255 199 256 200 
<< m1 >>
rect 260 199 261 200 
<< m1 >>
rect 262 199 263 200 
<< m2 >>
rect 262 199 263 200 
<< m1 >>
rect 265 199 266 200 
<< m1 >>
rect 268 199 269 200 
<< m2 >>
rect 269 199 270 200 
<< m1 >>
rect 270 199 271 200 
<< m2 >>
rect 270 199 271 200 
<< m2c >>
rect 270 199 271 200 
<< m1 >>
rect 270 199 271 200 
<< m2 >>
rect 270 199 271 200 
<< m2 >>
rect 271 199 272 200 
<< m1 >>
rect 272 199 273 200 
<< m1 >>
rect 274 199 275 200 
<< m2 >>
rect 275 199 276 200 
<< m1 >>
rect 289 199 290 200 
<< m1 >>
rect 307 199 308 200 
<< m1 >>
rect 325 199 326 200 
<< m1 >>
rect 327 199 328 200 
<< m1 >>
rect 340 199 341 200 
<< m1 >>
rect 343 199 344 200 
<< m2 >>
rect 343 199 344 200 
<< m1 >>
rect 345 199 346 200 
<< m1 >>
rect 10 200 11 201 
<< m1 >>
rect 19 200 20 201 
<< m1 >>
rect 21 200 22 201 
<< m2 >>
rect 27 200 28 201 
<< m1 >>
rect 28 200 29 201 
<< m1 >>
rect 37 200 38 201 
<< m2 >>
rect 38 200 39 201 
<< m1 >>
rect 44 200 45 201 
<< m1 >>
rect 46 200 47 201 
<< m1 >>
rect 56 200 57 201 
<< m1 >>
rect 58 200 59 201 
<< m1 >>
rect 62 200 63 201 
<< m1 >>
rect 64 200 65 201 
<< m2 >>
rect 79 200 80 201 
<< m1 >>
rect 80 200 81 201 
<< m1 >>
rect 82 200 83 201 
<< m1 >>
rect 106 200 107 201 
<< m1 >>
rect 118 200 119 201 
<< m1 >>
rect 130 200 131 201 
<< m1 >>
rect 132 200 133 201 
<< m1 >>
rect 134 200 135 201 
<< m1 >>
rect 136 200 137 201 
<< m1 >>
rect 138 200 139 201 
<< m1 >>
rect 145 200 146 201 
<< m2 >>
rect 146 200 147 201 
<< m1 >>
rect 147 200 148 201 
<< m2 >>
rect 147 200 148 201 
<< m2c >>
rect 147 200 148 201 
<< m1 >>
rect 147 200 148 201 
<< m2 >>
rect 147 200 148 201 
<< m1 >>
rect 148 200 149 201 
<< m1 >>
rect 149 200 150 201 
<< m2 >>
rect 149 200 150 201 
<< m2c >>
rect 149 200 150 201 
<< m1 >>
rect 149 200 150 201 
<< m2 >>
rect 149 200 150 201 
<< m1 >>
rect 158 200 159 201 
<< m2 >>
rect 158 200 159 201 
<< m2c >>
rect 158 200 159 201 
<< m1 >>
rect 158 200 159 201 
<< m2 >>
rect 158 200 159 201 
<< m1 >>
rect 159 200 160 201 
<< m1 >>
rect 160 200 161 201 
<< m1 >>
rect 163 200 164 201 
<< m1 >>
rect 165 200 166 201 
<< m1 >>
rect 170 200 171 201 
<< m2 >>
rect 170 200 171 201 
<< m2c >>
rect 170 200 171 201 
<< m1 >>
rect 170 200 171 201 
<< m2 >>
rect 170 200 171 201 
<< m2 >>
rect 171 200 172 201 
<< m1 >>
rect 172 200 173 201 
<< m2 >>
rect 172 200 173 201 
<< m2 >>
rect 173 200 174 201 
<< m1 >>
rect 174 200 175 201 
<< m2 >>
rect 174 200 175 201 
<< m2c >>
rect 174 200 175 201 
<< m1 >>
rect 174 200 175 201 
<< m2 >>
rect 174 200 175 201 
<< m1 >>
rect 177 200 178 201 
<< m2 >>
rect 177 200 178 201 
<< m2c >>
rect 177 200 178 201 
<< m1 >>
rect 177 200 178 201 
<< m2 >>
rect 177 200 178 201 
<< m1 >>
rect 178 200 179 201 
<< m1 >>
rect 179 200 180 201 
<< m1 >>
rect 181 200 182 201 
<< m1 >>
rect 183 200 184 201 
<< m1 >>
rect 188 200 189 201 
<< m1 >>
rect 190 200 191 201 
<< m1 >>
rect 193 200 194 201 
<< m1 >>
rect 194 200 195 201 
<< m2 >>
rect 194 200 195 201 
<< m2c >>
rect 194 200 195 201 
<< m1 >>
rect 194 200 195 201 
<< m2 >>
rect 194 200 195 201 
<< m1 >>
rect 197 200 198 201 
<< m1 >>
rect 199 200 200 201 
<< m1 >>
rect 201 200 202 201 
<< m1 >>
rect 218 200 219 201 
<< m2 >>
rect 225 200 226 201 
<< m1 >>
rect 226 200 227 201 
<< m1 >>
rect 232 200 233 201 
<< m1 >>
rect 235 200 236 201 
<< m1 >>
rect 237 200 238 201 
<< m1 >>
rect 241 200 242 201 
<< m1 >>
rect 243 200 244 201 
<< m1 >>
rect 255 200 256 201 
<< m1 >>
rect 260 200 261 201 
<< m1 >>
rect 262 200 263 201 
<< m2 >>
rect 262 200 263 201 
<< m1 >>
rect 265 200 266 201 
<< m1 >>
rect 266 200 267 201 
<< m2 >>
rect 266 200 267 201 
<< m2c >>
rect 266 200 267 201 
<< m1 >>
rect 266 200 267 201 
<< m2 >>
rect 266 200 267 201 
<< m2 >>
rect 267 200 268 201 
<< m1 >>
rect 268 200 269 201 
<< m2 >>
rect 268 200 269 201 
<< m2 >>
rect 269 200 270 201 
<< m1 >>
rect 272 200 273 201 
<< m1 >>
rect 274 200 275 201 
<< m2 >>
rect 275 200 276 201 
<< m1 >>
rect 289 200 290 201 
<< m2 >>
rect 289 200 290 201 
<< m2c >>
rect 289 200 290 201 
<< m1 >>
rect 289 200 290 201 
<< m2 >>
rect 289 200 290 201 
<< m1 >>
rect 307 200 308 201 
<< m2 >>
rect 307 200 308 201 
<< m2c >>
rect 307 200 308 201 
<< m1 >>
rect 307 200 308 201 
<< m2 >>
rect 307 200 308 201 
<< m1 >>
rect 323 200 324 201 
<< m2 >>
rect 323 200 324 201 
<< m2c >>
rect 323 200 324 201 
<< m1 >>
rect 323 200 324 201 
<< m2 >>
rect 323 200 324 201 
<< m1 >>
rect 324 200 325 201 
<< m1 >>
rect 325 200 326 201 
<< m1 >>
rect 327 200 328 201 
<< m2 >>
rect 327 200 328 201 
<< m2c >>
rect 327 200 328 201 
<< m1 >>
rect 327 200 328 201 
<< m2 >>
rect 327 200 328 201 
<< m1 >>
rect 340 200 341 201 
<< m1 >>
rect 343 200 344 201 
<< m2 >>
rect 343 200 344 201 
<< m1 >>
rect 345 200 346 201 
<< m1 >>
rect 10 201 11 202 
<< m1 >>
rect 19 201 20 202 
<< m1 >>
rect 21 201 22 202 
<< m2 >>
rect 27 201 28 202 
<< m1 >>
rect 28 201 29 202 
<< m1 >>
rect 37 201 38 202 
<< m2 >>
rect 38 201 39 202 
<< m1 >>
rect 44 201 45 202 
<< m1 >>
rect 46 201 47 202 
<< m1 >>
rect 56 201 57 202 
<< m1 >>
rect 58 201 59 202 
<< m1 >>
rect 62 201 63 202 
<< m1 >>
rect 64 201 65 202 
<< m2 >>
rect 79 201 80 202 
<< m1 >>
rect 80 201 81 202 
<< m1 >>
rect 82 201 83 202 
<< m1 >>
rect 106 201 107 202 
<< m1 >>
rect 118 201 119 202 
<< m1 >>
rect 130 201 131 202 
<< m1 >>
rect 132 201 133 202 
<< m1 >>
rect 134 201 135 202 
<< m2 >>
rect 134 201 135 202 
<< m2c >>
rect 134 201 135 202 
<< m1 >>
rect 134 201 135 202 
<< m2 >>
rect 134 201 135 202 
<< m2 >>
rect 135 201 136 202 
<< m1 >>
rect 136 201 137 202 
<< m1 >>
rect 138 201 139 202 
<< m1 >>
rect 145 201 146 202 
<< m2 >>
rect 149 201 150 202 
<< m2 >>
rect 158 201 159 202 
<< m1 >>
rect 163 201 164 202 
<< m1 >>
rect 165 201 166 202 
<< m1 >>
rect 172 201 173 202 
<< m1 >>
rect 174 201 175 202 
<< m2 >>
rect 177 201 178 202 
<< m1 >>
rect 181 201 182 202 
<< m1 >>
rect 183 201 184 202 
<< m1 >>
rect 188 201 189 202 
<< m1 >>
rect 190 201 191 202 
<< m2 >>
rect 194 201 195 202 
<< m1 >>
rect 197 201 198 202 
<< m1 >>
rect 199 201 200 202 
<< m1 >>
rect 201 201 202 202 
<< m1 >>
rect 218 201 219 202 
<< m2 >>
rect 225 201 226 202 
<< m1 >>
rect 226 201 227 202 
<< m1 >>
rect 232 201 233 202 
<< m1 >>
rect 235 201 236 202 
<< m1 >>
rect 237 201 238 202 
<< m1 >>
rect 241 201 242 202 
<< m1 >>
rect 243 201 244 202 
<< m1 >>
rect 255 201 256 202 
<< m1 >>
rect 260 201 261 202 
<< m1 >>
rect 262 201 263 202 
<< m2 >>
rect 262 201 263 202 
<< m1 >>
rect 268 201 269 202 
<< m1 >>
rect 272 201 273 202 
<< m1 >>
rect 274 201 275 202 
<< m2 >>
rect 275 201 276 202 
<< m2 >>
rect 289 201 290 202 
<< m2 >>
rect 290 201 291 202 
<< m2 >>
rect 291 201 292 202 
<< m2 >>
rect 292 201 293 202 
<< m2 >>
rect 293 201 294 202 
<< m2 >>
rect 294 201 295 202 
<< m2 >>
rect 295 201 296 202 
<< m2 >>
rect 296 201 297 202 
<< m2 >>
rect 297 201 298 202 
<< m2 >>
rect 298 201 299 202 
<< m2 >>
rect 307 201 308 202 
<< m2 >>
rect 323 201 324 202 
<< m2 >>
rect 327 201 328 202 
<< m1 >>
rect 340 201 341 202 
<< m1 >>
rect 343 201 344 202 
<< m2 >>
rect 343 201 344 202 
<< m1 >>
rect 345 201 346 202 
<< m1 >>
rect 10 202 11 203 
<< m1 >>
rect 19 202 20 203 
<< m1 >>
rect 21 202 22 203 
<< m2 >>
rect 27 202 28 203 
<< m1 >>
rect 28 202 29 203 
<< m1 >>
rect 37 202 38 203 
<< m2 >>
rect 38 202 39 203 
<< m1 >>
rect 44 202 45 203 
<< m1 >>
rect 46 202 47 203 
<< m1 >>
rect 56 202 57 203 
<< m1 >>
rect 58 202 59 203 
<< m1 >>
rect 62 202 63 203 
<< m1 >>
rect 64 202 65 203 
<< m2 >>
rect 79 202 80 203 
<< m1 >>
rect 80 202 81 203 
<< m1 >>
rect 82 202 83 203 
<< m1 >>
rect 100 202 101 203 
<< m1 >>
rect 101 202 102 203 
<< m1 >>
rect 102 202 103 203 
<< m1 >>
rect 103 202 104 203 
<< m1 >>
rect 104 202 105 203 
<< m1 >>
rect 105 202 106 203 
<< m1 >>
rect 106 202 107 203 
<< m1 >>
rect 118 202 119 203 
<< m1 >>
rect 130 202 131 203 
<< m1 >>
rect 132 202 133 203 
<< m2 >>
rect 135 202 136 203 
<< m1 >>
rect 136 202 137 203 
<< m1 >>
rect 138 202 139 203 
<< m1 >>
rect 139 202 140 203 
<< m1 >>
rect 140 202 141 203 
<< m1 >>
rect 141 202 142 203 
<< m1 >>
rect 142 202 143 203 
<< m1 >>
rect 143 202 144 203 
<< m2 >>
rect 143 202 144 203 
<< m2c >>
rect 143 202 144 203 
<< m1 >>
rect 143 202 144 203 
<< m2 >>
rect 143 202 144 203 
<< m2 >>
rect 144 202 145 203 
<< m1 >>
rect 145 202 146 203 
<< m2 >>
rect 145 202 146 203 
<< m2 >>
rect 146 202 147 203 
<< m1 >>
rect 147 202 148 203 
<< m2 >>
rect 147 202 148 203 
<< m2c >>
rect 147 202 148 203 
<< m1 >>
rect 147 202 148 203 
<< m2 >>
rect 147 202 148 203 
<< m1 >>
rect 148 202 149 203 
<< m1 >>
rect 149 202 150 203 
<< m2 >>
rect 149 202 150 203 
<< m1 >>
rect 150 202 151 203 
<< m1 >>
rect 151 202 152 203 
<< m1 >>
rect 152 202 153 203 
<< m1 >>
rect 153 202 154 203 
<< m1 >>
rect 154 202 155 203 
<< m1 >>
rect 155 202 156 203 
<< m1 >>
rect 156 202 157 203 
<< m1 >>
rect 157 202 158 203 
<< m1 >>
rect 158 202 159 203 
<< m2 >>
rect 158 202 159 203 
<< m1 >>
rect 159 202 160 203 
<< m1 >>
rect 160 202 161 203 
<< m1 >>
rect 161 202 162 203 
<< m2 >>
rect 161 202 162 203 
<< m2c >>
rect 161 202 162 203 
<< m1 >>
rect 161 202 162 203 
<< m2 >>
rect 161 202 162 203 
<< m2 >>
rect 162 202 163 203 
<< m1 >>
rect 163 202 164 203 
<< m2 >>
rect 163 202 164 203 
<< m2 >>
rect 164 202 165 203 
<< m1 >>
rect 165 202 166 203 
<< m2 >>
rect 165 202 166 203 
<< m2 >>
rect 166 202 167 203 
<< m1 >>
rect 167 202 168 203 
<< m2 >>
rect 167 202 168 203 
<< m2c >>
rect 167 202 168 203 
<< m1 >>
rect 167 202 168 203 
<< m2 >>
rect 167 202 168 203 
<< m1 >>
rect 172 202 173 203 
<< m2 >>
rect 172 202 173 203 
<< m2c >>
rect 172 202 173 203 
<< m1 >>
rect 172 202 173 203 
<< m2 >>
rect 172 202 173 203 
<< m1 >>
rect 174 202 175 203 
<< m1 >>
rect 175 202 176 203 
<< m1 >>
rect 176 202 177 203 
<< m1 >>
rect 177 202 178 203 
<< m2 >>
rect 177 202 178 203 
<< m1 >>
rect 178 202 179 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m2c >>
rect 179 202 180 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m2 >>
rect 180 202 181 203 
<< m1 >>
rect 181 202 182 203 
<< m2 >>
rect 181 202 182 203 
<< m1 >>
rect 183 202 184 203 
<< m1 >>
rect 186 202 187 203 
<< m2 >>
rect 186 202 187 203 
<< m2c >>
rect 186 202 187 203 
<< m1 >>
rect 186 202 187 203 
<< m2 >>
rect 186 202 187 203 
<< m2 >>
rect 187 202 188 203 
<< m1 >>
rect 188 202 189 203 
<< m2 >>
rect 188 202 189 203 
<< m2 >>
rect 189 202 190 203 
<< m1 >>
rect 190 202 191 203 
<< m2 >>
rect 190 202 191 203 
<< m2 >>
rect 191 202 192 203 
<< m1 >>
rect 192 202 193 203 
<< m2 >>
rect 192 202 193 203 
<< m2c >>
rect 192 202 193 203 
<< m1 >>
rect 192 202 193 203 
<< m2 >>
rect 192 202 193 203 
<< m1 >>
rect 193 202 194 203 
<< m1 >>
rect 194 202 195 203 
<< m2 >>
rect 194 202 195 203 
<< m1 >>
rect 195 202 196 203 
<< m1 >>
rect 196 202 197 203 
<< m1 >>
rect 197 202 198 203 
<< m1 >>
rect 199 202 200 203 
<< m1 >>
rect 201 202 202 203 
<< m1 >>
rect 218 202 219 203 
<< m2 >>
rect 225 202 226 203 
<< m1 >>
rect 226 202 227 203 
<< m1 >>
rect 232 202 233 203 
<< m1 >>
rect 235 202 236 203 
<< m1 >>
rect 237 202 238 203 
<< m1 >>
rect 241 202 242 203 
<< m1 >>
rect 243 202 244 203 
<< m1 >>
rect 255 202 256 203 
<< m1 >>
rect 260 202 261 203 
<< m1 >>
rect 262 202 263 203 
<< m2 >>
rect 262 202 263 203 
<< m1 >>
rect 268 202 269 203 
<< m1 >>
rect 272 202 273 203 
<< m1 >>
rect 274 202 275 203 
<< m1 >>
rect 275 202 276 203 
<< m2 >>
rect 275 202 276 203 
<< m1 >>
rect 276 202 277 203 
<< m1 >>
rect 277 202 278 203 
<< m1 >>
rect 278 202 279 203 
<< m1 >>
rect 279 202 280 203 
<< m1 >>
rect 280 202 281 203 
<< m1 >>
rect 281 202 282 203 
<< m1 >>
rect 282 202 283 203 
<< m1 >>
rect 283 202 284 203 
<< m1 >>
rect 284 202 285 203 
<< m1 >>
rect 285 202 286 203 
<< m1 >>
rect 286 202 287 203 
<< m1 >>
rect 287 202 288 203 
<< m1 >>
rect 288 202 289 203 
<< m1 >>
rect 289 202 290 203 
<< m1 >>
rect 290 202 291 203 
<< m1 >>
rect 291 202 292 203 
<< m1 >>
rect 292 202 293 203 
<< m1 >>
rect 293 202 294 203 
<< m1 >>
rect 294 202 295 203 
<< m1 >>
rect 295 202 296 203 
<< m1 >>
rect 296 202 297 203 
<< m1 >>
rect 297 202 298 203 
<< m1 >>
rect 298 202 299 203 
<< m2 >>
rect 298 202 299 203 
<< m1 >>
rect 299 202 300 203 
<< m2 >>
rect 299 202 300 203 
<< m1 >>
rect 300 202 301 203 
<< m2 >>
rect 300 202 301 203 
<< m1 >>
rect 301 202 302 203 
<< m2 >>
rect 301 202 302 203 
<< m1 >>
rect 302 202 303 203 
<< m2 >>
rect 302 202 303 203 
<< m1 >>
rect 303 202 304 203 
<< m1 >>
rect 304 202 305 203 
<< m1 >>
rect 305 202 306 203 
<< m1 >>
rect 306 202 307 203 
<< m1 >>
rect 307 202 308 203 
<< m2 >>
rect 307 202 308 203 
<< m1 >>
rect 308 202 309 203 
<< m2 >>
rect 308 202 309 203 
<< m1 >>
rect 309 202 310 203 
<< m2 >>
rect 309 202 310 203 
<< m1 >>
rect 310 202 311 203 
<< m2 >>
rect 310 202 311 203 
<< m1 >>
rect 311 202 312 203 
<< m2 >>
rect 311 202 312 203 
<< m1 >>
rect 312 202 313 203 
<< m2 >>
rect 312 202 313 203 
<< m1 >>
rect 313 202 314 203 
<< m2 >>
rect 313 202 314 203 
<< m1 >>
rect 314 202 315 203 
<< m2 >>
rect 314 202 315 203 
<< m1 >>
rect 315 202 316 203 
<< m2 >>
rect 315 202 316 203 
<< m1 >>
rect 316 202 317 203 
<< m2 >>
rect 316 202 317 203 
<< m1 >>
rect 317 202 318 203 
<< m2 >>
rect 317 202 318 203 
<< m1 >>
rect 318 202 319 203 
<< m2 >>
rect 318 202 319 203 
<< m1 >>
rect 319 202 320 203 
<< m2 >>
rect 319 202 320 203 
<< m1 >>
rect 320 202 321 203 
<< m2 >>
rect 320 202 321 203 
<< m1 >>
rect 321 202 322 203 
<< m1 >>
rect 322 202 323 203 
<< m1 >>
rect 323 202 324 203 
<< m2 >>
rect 323 202 324 203 
<< m1 >>
rect 324 202 325 203 
<< m1 >>
rect 325 202 326 203 
<< m1 >>
rect 326 202 327 203 
<< m1 >>
rect 327 202 328 203 
<< m2 >>
rect 327 202 328 203 
<< m1 >>
rect 328 202 329 203 
<< m1 >>
rect 329 202 330 203 
<< m1 >>
rect 330 202 331 203 
<< m1 >>
rect 331 202 332 203 
<< m1 >>
rect 332 202 333 203 
<< m1 >>
rect 333 202 334 203 
<< m1 >>
rect 334 202 335 203 
<< m1 >>
rect 335 202 336 203 
<< m1 >>
rect 336 202 337 203 
<< m1 >>
rect 337 202 338 203 
<< m1 >>
rect 338 202 339 203 
<< m1 >>
rect 339 202 340 203 
<< m1 >>
rect 340 202 341 203 
<< m1 >>
rect 343 202 344 203 
<< m2 >>
rect 343 202 344 203 
<< m1 >>
rect 345 202 346 203 
<< m1 >>
rect 10 203 11 204 
<< m1 >>
rect 19 203 20 204 
<< m1 >>
rect 21 203 22 204 
<< m2 >>
rect 27 203 28 204 
<< m1 >>
rect 28 203 29 204 
<< m1 >>
rect 37 203 38 204 
<< m2 >>
rect 38 203 39 204 
<< m1 >>
rect 44 203 45 204 
<< m1 >>
rect 46 203 47 204 
<< m1 >>
rect 56 203 57 204 
<< m1 >>
rect 58 203 59 204 
<< m1 >>
rect 62 203 63 204 
<< m1 >>
rect 64 203 65 204 
<< m2 >>
rect 79 203 80 204 
<< m1 >>
rect 80 203 81 204 
<< m1 >>
rect 82 203 83 204 
<< m1 >>
rect 100 203 101 204 
<< m1 >>
rect 118 203 119 204 
<< m1 >>
rect 130 203 131 204 
<< m1 >>
rect 132 203 133 204 
<< m2 >>
rect 135 203 136 204 
<< m1 >>
rect 136 203 137 204 
<< m1 >>
rect 145 203 146 204 
<< m2 >>
rect 149 203 150 204 
<< m2 >>
rect 158 203 159 204 
<< m1 >>
rect 163 203 164 204 
<< m1 >>
rect 165 203 166 204 
<< m1 >>
rect 167 203 168 204 
<< m2 >>
rect 172 203 173 204 
<< m2 >>
rect 177 203 178 204 
<< m1 >>
rect 181 203 182 204 
<< m2 >>
rect 181 203 182 204 
<< m1 >>
rect 183 203 184 204 
<< m1 >>
rect 186 203 187 204 
<< m1 >>
rect 188 203 189 204 
<< m1 >>
rect 190 203 191 204 
<< m2 >>
rect 194 203 195 204 
<< m1 >>
rect 199 203 200 204 
<< m1 >>
rect 201 203 202 204 
<< m1 >>
rect 218 203 219 204 
<< m2 >>
rect 225 203 226 204 
<< m1 >>
rect 226 203 227 204 
<< m1 >>
rect 232 203 233 204 
<< m1 >>
rect 235 203 236 204 
<< m1 >>
rect 237 203 238 204 
<< m1 >>
rect 241 203 242 204 
<< m1 >>
rect 243 203 244 204 
<< m1 >>
rect 253 203 254 204 
<< m2 >>
rect 253 203 254 204 
<< m2c >>
rect 253 203 254 204 
<< m1 >>
rect 253 203 254 204 
<< m2 >>
rect 253 203 254 204 
<< m1 >>
rect 254 203 255 204 
<< m1 >>
rect 255 203 256 204 
<< m1 >>
rect 260 203 261 204 
<< m1 >>
rect 262 203 263 204 
<< m2 >>
rect 262 203 263 204 
<< m1 >>
rect 268 203 269 204 
<< m1 >>
rect 272 203 273 204 
<< m2 >>
rect 275 203 276 204 
<< m2 >>
rect 276 203 277 204 
<< m2 >>
rect 277 203 278 204 
<< m2 >>
rect 278 203 279 204 
<< m2 >>
rect 279 203 280 204 
<< m2 >>
rect 280 203 281 204 
<< m2 >>
rect 281 203 282 204 
<< m2 >>
rect 282 203 283 204 
<< m2 >>
rect 283 203 284 204 
<< m2 >>
rect 284 203 285 204 
<< m2 >>
rect 285 203 286 204 
<< m2 >>
rect 286 203 287 204 
<< m2 >>
rect 287 203 288 204 
<< m2 >>
rect 288 203 289 204 
<< m2 >>
rect 289 203 290 204 
<< m2 >>
rect 290 203 291 204 
<< m2 >>
rect 291 203 292 204 
<< m2 >>
rect 292 203 293 204 
<< m2 >>
rect 293 203 294 204 
<< m2 >>
rect 294 203 295 204 
<< m2 >>
rect 295 203 296 204 
<< m2 >>
rect 296 203 297 204 
<< m2 >>
rect 297 203 298 204 
<< m2 >>
rect 298 203 299 204 
<< m2 >>
rect 302 203 303 204 
<< m2 >>
rect 320 203 321 204 
<< m2 >>
rect 323 203 324 204 
<< m2 >>
rect 327 203 328 204 
<< m1 >>
rect 343 203 344 204 
<< m2 >>
rect 343 203 344 204 
<< m1 >>
rect 345 203 346 204 
<< m1 >>
rect 10 204 11 205 
<< m1 >>
rect 19 204 20 205 
<< m1 >>
rect 21 204 22 205 
<< m2 >>
rect 27 204 28 205 
<< m1 >>
rect 28 204 29 205 
<< m1 >>
rect 37 204 38 205 
<< m2 >>
rect 38 204 39 205 
<< m1 >>
rect 44 204 45 205 
<< m1 >>
rect 46 204 47 205 
<< m1 >>
rect 56 204 57 205 
<< m1 >>
rect 58 204 59 205 
<< m1 >>
rect 62 204 63 205 
<< m1 >>
rect 64 204 65 205 
<< m2 >>
rect 79 204 80 205 
<< m1 >>
rect 80 204 81 205 
<< m1 >>
rect 82 204 83 205 
<< m1 >>
rect 100 204 101 205 
<< m1 >>
rect 118 204 119 205 
<< m1 >>
rect 130 204 131 205 
<< m1 >>
rect 132 204 133 205 
<< m2 >>
rect 135 204 136 205 
<< m1 >>
rect 136 204 137 205 
<< m2 >>
rect 136 204 137 205 
<< m2 >>
rect 137 204 138 205 
<< m1 >>
rect 138 204 139 205 
<< m2 >>
rect 138 204 139 205 
<< m2c >>
rect 138 204 139 205 
<< m1 >>
rect 138 204 139 205 
<< m2 >>
rect 138 204 139 205 
<< m1 >>
rect 139 204 140 205 
<< m1 >>
rect 140 204 141 205 
<< m1 >>
rect 141 204 142 205 
<< m1 >>
rect 142 204 143 205 
<< m1 >>
rect 143 204 144 205 
<< m2 >>
rect 143 204 144 205 
<< m2c >>
rect 143 204 144 205 
<< m1 >>
rect 143 204 144 205 
<< m2 >>
rect 143 204 144 205 
<< m2 >>
rect 144 204 145 205 
<< m1 >>
rect 145 204 146 205 
<< m2 >>
rect 145 204 146 205 
<< m2 >>
rect 146 204 147 205 
<< m1 >>
rect 147 204 148 205 
<< m2 >>
rect 147 204 148 205 
<< m2c >>
rect 147 204 148 205 
<< m1 >>
rect 147 204 148 205 
<< m2 >>
rect 147 204 148 205 
<< m1 >>
rect 148 204 149 205 
<< m1 >>
rect 149 204 150 205 
<< m2 >>
rect 149 204 150 205 
<< m1 >>
rect 150 204 151 205 
<< m1 >>
rect 151 204 152 205 
<< m1 >>
rect 152 204 153 205 
<< m1 >>
rect 153 204 154 205 
<< m1 >>
rect 154 204 155 205 
<< m1 >>
rect 155 204 156 205 
<< m1 >>
rect 156 204 157 205 
<< m1 >>
rect 157 204 158 205 
<< m1 >>
rect 158 204 159 205 
<< m2 >>
rect 158 204 159 205 
<< m1 >>
rect 159 204 160 205 
<< m1 >>
rect 160 204 161 205 
<< m1 >>
rect 161 204 162 205 
<< m2 >>
rect 161 204 162 205 
<< m2c >>
rect 161 204 162 205 
<< m1 >>
rect 161 204 162 205 
<< m2 >>
rect 161 204 162 205 
<< m2 >>
rect 162 204 163 205 
<< m1 >>
rect 163 204 164 205 
<< m2 >>
rect 163 204 164 205 
<< m2 >>
rect 164 204 165 205 
<< m1 >>
rect 165 204 166 205 
<< m2 >>
rect 165 204 166 205 
<< m2 >>
rect 166 204 167 205 
<< m1 >>
rect 167 204 168 205 
<< m2 >>
rect 167 204 168 205 
<< m2 >>
rect 168 204 169 205 
<< m1 >>
rect 169 204 170 205 
<< m2 >>
rect 169 204 170 205 
<< m2c >>
rect 169 204 170 205 
<< m1 >>
rect 169 204 170 205 
<< m2 >>
rect 169 204 170 205 
<< m1 >>
rect 170 204 171 205 
<< m1 >>
rect 171 204 172 205 
<< m1 >>
rect 172 204 173 205 
<< m2 >>
rect 172 204 173 205 
<< m1 >>
rect 173 204 174 205 
<< m1 >>
rect 174 204 175 205 
<< m1 >>
rect 175 204 176 205 
<< m1 >>
rect 176 204 177 205 
<< m1 >>
rect 177 204 178 205 
<< m2 >>
rect 177 204 178 205 
<< m1 >>
rect 178 204 179 205 
<< m1 >>
rect 179 204 180 205 
<< m1 >>
rect 180 204 181 205 
<< m1 >>
rect 181 204 182 205 
<< m2 >>
rect 181 204 182 205 
<< m1 >>
rect 183 204 184 205 
<< m1 >>
rect 186 204 187 205 
<< m1 >>
rect 188 204 189 205 
<< m1 >>
rect 190 204 191 205 
<< m1 >>
rect 194 204 195 205 
<< m2 >>
rect 194 204 195 205 
<< m2c >>
rect 194 204 195 205 
<< m1 >>
rect 194 204 195 205 
<< m2 >>
rect 194 204 195 205 
<< m1 >>
rect 199 204 200 205 
<< m1 >>
rect 201 204 202 205 
<< m1 >>
rect 218 204 219 205 
<< m2 >>
rect 225 204 226 205 
<< m1 >>
rect 226 204 227 205 
<< m1 >>
rect 232 204 233 205 
<< m1 >>
rect 235 204 236 205 
<< m1 >>
rect 237 204 238 205 
<< m1 >>
rect 241 204 242 205 
<< m1 >>
rect 243 204 244 205 
<< m2 >>
rect 253 204 254 205 
<< m1 >>
rect 260 204 261 205 
<< m1 >>
rect 262 204 263 205 
<< m2 >>
rect 262 204 263 205 
<< m1 >>
rect 268 204 269 205 
<< m1 >>
rect 272 204 273 205 
<< m1 >>
rect 298 204 299 205 
<< m2 >>
rect 298 204 299 205 
<< m2c >>
rect 298 204 299 205 
<< m1 >>
rect 298 204 299 205 
<< m2 >>
rect 298 204 299 205 
<< m2 >>
rect 302 204 303 205 
<< m2 >>
rect 320 204 321 205 
<< m1 >>
rect 323 204 324 205 
<< m2 >>
rect 323 204 324 205 
<< m2c >>
rect 323 204 324 205 
<< m1 >>
rect 323 204 324 205 
<< m2 >>
rect 323 204 324 205 
<< m1 >>
rect 327 204 328 205 
<< m2 >>
rect 327 204 328 205 
<< m2c >>
rect 327 204 328 205 
<< m1 >>
rect 327 204 328 205 
<< m2 >>
rect 327 204 328 205 
<< m1 >>
rect 343 204 344 205 
<< m2 >>
rect 343 204 344 205 
<< m1 >>
rect 345 204 346 205 
<< m1 >>
rect 10 205 11 206 
<< m1 >>
rect 19 205 20 206 
<< m1 >>
rect 21 205 22 206 
<< m2 >>
rect 27 205 28 206 
<< m1 >>
rect 28 205 29 206 
<< m1 >>
rect 37 205 38 206 
<< m2 >>
rect 38 205 39 206 
<< m1 >>
rect 44 205 45 206 
<< m1 >>
rect 46 205 47 206 
<< m1 >>
rect 56 205 57 206 
<< m1 >>
rect 58 205 59 206 
<< m1 >>
rect 62 205 63 206 
<< m1 >>
rect 64 205 65 206 
<< m2 >>
rect 79 205 80 206 
<< m1 >>
rect 80 205 81 206 
<< m1 >>
rect 82 205 83 206 
<< m1 >>
rect 100 205 101 206 
<< m1 >>
rect 118 205 119 206 
<< m1 >>
rect 130 205 131 206 
<< m1 >>
rect 132 205 133 206 
<< m1 >>
rect 136 205 137 206 
<< m1 >>
rect 145 205 146 206 
<< m2 >>
rect 149 205 150 206 
<< m2 >>
rect 154 205 155 206 
<< m2 >>
rect 155 205 156 206 
<< m2 >>
rect 156 205 157 206 
<< m2 >>
rect 157 205 158 206 
<< m2 >>
rect 158 205 159 206 
<< m1 >>
rect 163 205 164 206 
<< m1 >>
rect 165 205 166 206 
<< m1 >>
rect 167 205 168 206 
<< m2 >>
rect 172 205 173 206 
<< m2 >>
rect 177 205 178 206 
<< m2 >>
rect 181 205 182 206 
<< m1 >>
rect 183 205 184 206 
<< m1 >>
rect 186 205 187 206 
<< m1 >>
rect 188 205 189 206 
<< m1 >>
rect 190 205 191 206 
<< m1 >>
rect 194 205 195 206 
<< m1 >>
rect 199 205 200 206 
<< m1 >>
rect 201 205 202 206 
<< m1 >>
rect 218 205 219 206 
<< m2 >>
rect 225 205 226 206 
<< m1 >>
rect 226 205 227 206 
<< m1 >>
rect 232 205 233 206 
<< m1 >>
rect 233 205 234 206 
<< m2 >>
rect 233 205 234 206 
<< m2c >>
rect 233 205 234 206 
<< m1 >>
rect 233 205 234 206 
<< m2 >>
rect 233 205 234 206 
<< m2 >>
rect 234 205 235 206 
<< m1 >>
rect 235 205 236 206 
<< m2 >>
rect 235 205 236 206 
<< m2 >>
rect 236 205 237 206 
<< m1 >>
rect 237 205 238 206 
<< m2 >>
rect 237 205 238 206 
<< m2 >>
rect 238 205 239 206 
<< m1 >>
rect 239 205 240 206 
<< m2 >>
rect 239 205 240 206 
<< m2c >>
rect 239 205 240 206 
<< m1 >>
rect 239 205 240 206 
<< m2 >>
rect 239 205 240 206 
<< m2 >>
rect 240 205 241 206 
<< m1 >>
rect 241 205 242 206 
<< m2 >>
rect 241 205 242 206 
<< m2 >>
rect 242 205 243 206 
<< m1 >>
rect 243 205 244 206 
<< m2 >>
rect 243 205 244 206 
<< m2 >>
rect 244 205 245 206 
<< m1 >>
rect 245 205 246 206 
<< m2 >>
rect 245 205 246 206 
<< m2c >>
rect 245 205 246 206 
<< m1 >>
rect 245 205 246 206 
<< m2 >>
rect 245 205 246 206 
<< m1 >>
rect 246 205 247 206 
<< m1 >>
rect 247 205 248 206 
<< m1 >>
rect 248 205 249 206 
<< m1 >>
rect 249 205 250 206 
<< m1 >>
rect 250 205 251 206 
<< m1 >>
rect 251 205 252 206 
<< m1 >>
rect 252 205 253 206 
<< m1 >>
rect 253 205 254 206 
<< m2 >>
rect 253 205 254 206 
<< m1 >>
rect 254 205 255 206 
<< m1 >>
rect 255 205 256 206 
<< m1 >>
rect 256 205 257 206 
<< m1 >>
rect 257 205 258 206 
<< m1 >>
rect 258 205 259 206 
<< m1 >>
rect 260 205 261 206 
<< m1 >>
rect 262 205 263 206 
<< m2 >>
rect 262 205 263 206 
<< m1 >>
rect 268 205 269 206 
<< m1 >>
rect 272 205 273 206 
<< m1 >>
rect 298 205 299 206 
<< m1 >>
rect 300 205 301 206 
<< m1 >>
rect 301 205 302 206 
<< m1 >>
rect 302 205 303 206 
<< m2 >>
rect 302 205 303 206 
<< m1 >>
rect 303 205 304 206 
<< m1 >>
rect 304 205 305 206 
<< m1 >>
rect 305 205 306 206 
<< m1 >>
rect 306 205 307 206 
<< m1 >>
rect 307 205 308 206 
<< m1 >>
rect 308 205 309 206 
<< m1 >>
rect 309 205 310 206 
<< m1 >>
rect 310 205 311 206 
<< m1 >>
rect 311 205 312 206 
<< m1 >>
rect 312 205 313 206 
<< m1 >>
rect 313 205 314 206 
<< m1 >>
rect 314 205 315 206 
<< m1 >>
rect 315 205 316 206 
<< m1 >>
rect 316 205 317 206 
<< m1 >>
rect 317 205 318 206 
<< m1 >>
rect 318 205 319 206 
<< m1 >>
rect 319 205 320 206 
<< m1 >>
rect 320 205 321 206 
<< m2 >>
rect 320 205 321 206 
<< m2 >>
rect 323 205 324 206 
<< m1 >>
rect 327 205 328 206 
<< m1 >>
rect 343 205 344 206 
<< m2 >>
rect 343 205 344 206 
<< m1 >>
rect 345 205 346 206 
<< m1 >>
rect 10 206 11 207 
<< m1 >>
rect 19 206 20 207 
<< m1 >>
rect 21 206 22 207 
<< m2 >>
rect 27 206 28 207 
<< m1 >>
rect 28 206 29 207 
<< m1 >>
rect 37 206 38 207 
<< m2 >>
rect 38 206 39 207 
<< m1 >>
rect 44 206 45 207 
<< m1 >>
rect 46 206 47 207 
<< m1 >>
rect 56 206 57 207 
<< m1 >>
rect 58 206 59 207 
<< m1 >>
rect 62 206 63 207 
<< m1 >>
rect 64 206 65 207 
<< m2 >>
rect 79 206 80 207 
<< m1 >>
rect 80 206 81 207 
<< m1 >>
rect 82 206 83 207 
<< m1 >>
rect 100 206 101 207 
<< m1 >>
rect 118 206 119 207 
<< m1 >>
rect 130 206 131 207 
<< m1 >>
rect 132 206 133 207 
<< m1 >>
rect 136 206 137 207 
<< m1 >>
rect 145 206 146 207 
<< m1 >>
rect 149 206 150 207 
<< m2 >>
rect 149 206 150 207 
<< m2c >>
rect 149 206 150 207 
<< m1 >>
rect 149 206 150 207 
<< m2 >>
rect 149 206 150 207 
<< m1 >>
rect 154 206 155 207 
<< m2 >>
rect 154 206 155 207 
<< m2c >>
rect 154 206 155 207 
<< m1 >>
rect 154 206 155 207 
<< m2 >>
rect 154 206 155 207 
<< m1 >>
rect 163 206 164 207 
<< m1 >>
rect 165 206 166 207 
<< m1 >>
rect 167 206 168 207 
<< m1 >>
rect 172 206 173 207 
<< m2 >>
rect 172 206 173 207 
<< m2c >>
rect 172 206 173 207 
<< m1 >>
rect 172 206 173 207 
<< m2 >>
rect 172 206 173 207 
<< m1 >>
rect 177 206 178 207 
<< m2 >>
rect 177 206 178 207 
<< m2c >>
rect 177 206 178 207 
<< m1 >>
rect 177 206 178 207 
<< m2 >>
rect 177 206 178 207 
<< m1 >>
rect 178 206 179 207 
<< m1 >>
rect 181 206 182 207 
<< m2 >>
rect 181 206 182 207 
<< m2c >>
rect 181 206 182 207 
<< m1 >>
rect 181 206 182 207 
<< m2 >>
rect 181 206 182 207 
<< m1 >>
rect 183 206 184 207 
<< m1 >>
rect 186 206 187 207 
<< m1 >>
rect 188 206 189 207 
<< m1 >>
rect 190 206 191 207 
<< m1 >>
rect 194 206 195 207 
<< m1 >>
rect 199 206 200 207 
<< m1 >>
rect 201 206 202 207 
<< m1 >>
rect 218 206 219 207 
<< m2 >>
rect 225 206 226 207 
<< m1 >>
rect 226 206 227 207 
<< m1 >>
rect 235 206 236 207 
<< m1 >>
rect 237 206 238 207 
<< m1 >>
rect 241 206 242 207 
<< m1 >>
rect 243 206 244 207 
<< m2 >>
rect 253 206 254 207 
<< m1 >>
rect 258 206 259 207 
<< m1 >>
rect 260 206 261 207 
<< m1 >>
rect 262 206 263 207 
<< m2 >>
rect 262 206 263 207 
<< m1 >>
rect 268 206 269 207 
<< m1 >>
rect 272 206 273 207 
<< m1 >>
rect 298 206 299 207 
<< m1 >>
rect 300 206 301 207 
<< m2 >>
rect 302 206 303 207 
<< m1 >>
rect 320 206 321 207 
<< m2 >>
rect 320 206 321 207 
<< m1 >>
rect 321 206 322 207 
<< m1 >>
rect 322 206 323 207 
<< m1 >>
rect 323 206 324 207 
<< m2 >>
rect 323 206 324 207 
<< m1 >>
rect 324 206 325 207 
<< m1 >>
rect 325 206 326 207 
<< m2 >>
rect 325 206 326 207 
<< m2c >>
rect 325 206 326 207 
<< m1 >>
rect 325 206 326 207 
<< m2 >>
rect 325 206 326 207 
<< m2 >>
rect 326 206 327 207 
<< m1 >>
rect 327 206 328 207 
<< m2 >>
rect 327 206 328 207 
<< m2 >>
rect 328 206 329 207 
<< m1 >>
rect 329 206 330 207 
<< m2 >>
rect 329 206 330 207 
<< m2c >>
rect 329 206 330 207 
<< m1 >>
rect 329 206 330 207 
<< m2 >>
rect 329 206 330 207 
<< m1 >>
rect 343 206 344 207 
<< m2 >>
rect 343 206 344 207 
<< m1 >>
rect 345 206 346 207 
<< m1 >>
rect 10 207 11 208 
<< m1 >>
rect 13 207 14 208 
<< m1 >>
rect 14 207 15 208 
<< m1 >>
rect 15 207 16 208 
<< m1 >>
rect 16 207 17 208 
<< m1 >>
rect 17 207 18 208 
<< m2 >>
rect 17 207 18 208 
<< m2c >>
rect 17 207 18 208 
<< m1 >>
rect 17 207 18 208 
<< m2 >>
rect 17 207 18 208 
<< m2 >>
rect 18 207 19 208 
<< m1 >>
rect 19 207 20 208 
<< m2 >>
rect 19 207 20 208 
<< m2 >>
rect 20 207 21 208 
<< m1 >>
rect 21 207 22 208 
<< m2 >>
rect 21 207 22 208 
<< m2c >>
rect 21 207 22 208 
<< m1 >>
rect 21 207 22 208 
<< m2 >>
rect 21 207 22 208 
<< m2 >>
rect 27 207 28 208 
<< m1 >>
rect 28 207 29 208 
<< m1 >>
rect 37 207 38 208 
<< m2 >>
rect 38 207 39 208 
<< m1 >>
rect 44 207 45 208 
<< m1 >>
rect 46 207 47 208 
<< m1 >>
rect 56 207 57 208 
<< m1 >>
rect 58 207 59 208 
<< m1 >>
rect 62 207 63 208 
<< m1 >>
rect 64 207 65 208 
<< m2 >>
rect 79 207 80 208 
<< m1 >>
rect 80 207 81 208 
<< m1 >>
rect 82 207 83 208 
<< m1 >>
rect 100 207 101 208 
<< m1 >>
rect 118 207 119 208 
<< m1 >>
rect 130 207 131 208 
<< m1 >>
rect 132 207 133 208 
<< m1 >>
rect 136 207 137 208 
<< m1 >>
rect 145 207 146 208 
<< m1 >>
rect 149 207 150 208 
<< m1 >>
rect 154 207 155 208 
<< m1 >>
rect 163 207 164 208 
<< m1 >>
rect 165 207 166 208 
<< m1 >>
rect 167 207 168 208 
<< m1 >>
rect 172 207 173 208 
<< m1 >>
rect 178 207 179 208 
<< m1 >>
rect 181 207 182 208 
<< m1 >>
rect 183 207 184 208 
<< m1 >>
rect 186 207 187 208 
<< m1 >>
rect 188 207 189 208 
<< m1 >>
rect 190 207 191 208 
<< m1 >>
rect 194 207 195 208 
<< m1 >>
rect 199 207 200 208 
<< m1 >>
rect 201 207 202 208 
<< m1 >>
rect 218 207 219 208 
<< m2 >>
rect 225 207 226 208 
<< m1 >>
rect 226 207 227 208 
<< m1 >>
rect 235 207 236 208 
<< m1 >>
rect 237 207 238 208 
<< m1 >>
rect 241 207 242 208 
<< m1 >>
rect 243 207 244 208 
<< m1 >>
rect 253 207 254 208 
<< m2 >>
rect 253 207 254 208 
<< m2c >>
rect 253 207 254 208 
<< m1 >>
rect 253 207 254 208 
<< m2 >>
rect 253 207 254 208 
<< m1 >>
rect 256 207 257 208 
<< m2 >>
rect 256 207 257 208 
<< m2c >>
rect 256 207 257 208 
<< m1 >>
rect 256 207 257 208 
<< m2 >>
rect 256 207 257 208 
<< m2 >>
rect 257 207 258 208 
<< m1 >>
rect 258 207 259 208 
<< m2 >>
rect 258 207 259 208 
<< m2 >>
rect 259 207 260 208 
<< m1 >>
rect 260 207 261 208 
<< m2 >>
rect 260 207 261 208 
<< m2 >>
rect 261 207 262 208 
<< m1 >>
rect 262 207 263 208 
<< m2 >>
rect 262 207 263 208 
<< m1 >>
rect 268 207 269 208 
<< m1 >>
rect 269 207 270 208 
<< m1 >>
rect 270 207 271 208 
<< m1 >>
rect 272 207 273 208 
<< m1 >>
rect 298 207 299 208 
<< m1 >>
rect 300 207 301 208 
<< m1 >>
rect 302 207 303 208 
<< m2 >>
rect 302 207 303 208 
<< m2c >>
rect 302 207 303 208 
<< m1 >>
rect 302 207 303 208 
<< m2 >>
rect 302 207 303 208 
<< m1 >>
rect 303 207 304 208 
<< m1 >>
rect 304 207 305 208 
<< m1 >>
rect 305 207 306 208 
<< m1 >>
rect 306 207 307 208 
<< m1 >>
rect 307 207 308 208 
<< m2 >>
rect 320 207 321 208 
<< m2 >>
rect 323 207 324 208 
<< m1 >>
rect 327 207 328 208 
<< m1 >>
rect 329 207 330 208 
<< m1 >>
rect 343 207 344 208 
<< m2 >>
rect 343 207 344 208 
<< m1 >>
rect 345 207 346 208 
<< m1 >>
rect 10 208 11 209 
<< m1 >>
rect 13 208 14 209 
<< m1 >>
rect 19 208 20 209 
<< m2 >>
rect 27 208 28 209 
<< m1 >>
rect 28 208 29 209 
<< m1 >>
rect 37 208 38 209 
<< m2 >>
rect 38 208 39 209 
<< m1 >>
rect 44 208 45 209 
<< m1 >>
rect 46 208 47 209 
<< m1 >>
rect 56 208 57 209 
<< m1 >>
rect 58 208 59 209 
<< m1 >>
rect 62 208 63 209 
<< m1 >>
rect 64 208 65 209 
<< m2 >>
rect 79 208 80 209 
<< m1 >>
rect 80 208 81 209 
<< m1 >>
rect 82 208 83 209 
<< m1 >>
rect 100 208 101 209 
<< m1 >>
rect 118 208 119 209 
<< m1 >>
rect 130 208 131 209 
<< m1 >>
rect 132 208 133 209 
<< m1 >>
rect 136 208 137 209 
<< m1 >>
rect 145 208 146 209 
<< m1 >>
rect 149 208 150 209 
<< m1 >>
rect 154 208 155 209 
<< m1 >>
rect 163 208 164 209 
<< m1 >>
rect 165 208 166 209 
<< m1 >>
rect 167 208 168 209 
<< m1 >>
rect 172 208 173 209 
<< m1 >>
rect 178 208 179 209 
<< m1 >>
rect 181 208 182 209 
<< m1 >>
rect 183 208 184 209 
<< m1 >>
rect 186 208 187 209 
<< m1 >>
rect 188 208 189 209 
<< m1 >>
rect 190 208 191 209 
<< m1 >>
rect 193 208 194 209 
<< m1 >>
rect 194 208 195 209 
<< m1 >>
rect 199 208 200 209 
<< m1 >>
rect 201 208 202 209 
<< m1 >>
rect 218 208 219 209 
<< m2 >>
rect 225 208 226 209 
<< m1 >>
rect 226 208 227 209 
<< m1 >>
rect 235 208 236 209 
<< m1 >>
rect 237 208 238 209 
<< m1 >>
rect 241 208 242 209 
<< m1 >>
rect 243 208 244 209 
<< m1 >>
rect 253 208 254 209 
<< m1 >>
rect 256 208 257 209 
<< m1 >>
rect 258 208 259 209 
<< m1 >>
rect 260 208 261 209 
<< m1 >>
rect 262 208 263 209 
<< m1 >>
rect 270 208 271 209 
<< m2 >>
rect 270 208 271 209 
<< m2c >>
rect 270 208 271 209 
<< m1 >>
rect 270 208 271 209 
<< m2 >>
rect 270 208 271 209 
<< m2 >>
rect 271 208 272 209 
<< m1 >>
rect 272 208 273 209 
<< m2 >>
rect 272 208 273 209 
<< m2 >>
rect 273 208 274 209 
<< m2 >>
rect 297 208 298 209 
<< m1 >>
rect 298 208 299 209 
<< m2 >>
rect 298 208 299 209 
<< m2 >>
rect 299 208 300 209 
<< m1 >>
rect 300 208 301 209 
<< m2 >>
rect 300 208 301 209 
<< m2c >>
rect 300 208 301 209 
<< m1 >>
rect 300 208 301 209 
<< m2 >>
rect 300 208 301 209 
<< m1 >>
rect 307 208 308 209 
<< m1 >>
rect 320 208 321 209 
<< m2 >>
rect 320 208 321 209 
<< m2c >>
rect 320 208 321 209 
<< m1 >>
rect 320 208 321 209 
<< m2 >>
rect 320 208 321 209 
<< m1 >>
rect 321 208 322 209 
<< m1 >>
rect 322 208 323 209 
<< m2 >>
rect 323 208 324 209 
<< m1 >>
rect 324 208 325 209 
<< m2 >>
rect 324 208 325 209 
<< m2c >>
rect 324 208 325 209 
<< m1 >>
rect 324 208 325 209 
<< m2 >>
rect 324 208 325 209 
<< m1 >>
rect 325 208 326 209 
<< m1 >>
rect 327 208 328 209 
<< m1 >>
rect 329 208 330 209 
<< m1 >>
rect 343 208 344 209 
<< m2 >>
rect 343 208 344 209 
<< m1 >>
rect 345 208 346 209 
<< m1 >>
rect 10 209 11 210 
<< m1 >>
rect 13 209 14 210 
<< m1 >>
rect 19 209 20 210 
<< m2 >>
rect 27 209 28 210 
<< m1 >>
rect 28 209 29 210 
<< m1 >>
rect 37 209 38 210 
<< m2 >>
rect 38 209 39 210 
<< m1 >>
rect 44 209 45 210 
<< m1 >>
rect 46 209 47 210 
<< m1 >>
rect 56 209 57 210 
<< m1 >>
rect 58 209 59 210 
<< m1 >>
rect 62 209 63 210 
<< m1 >>
rect 64 209 65 210 
<< m2 >>
rect 79 209 80 210 
<< m1 >>
rect 80 209 81 210 
<< m1 >>
rect 82 209 83 210 
<< m1 >>
rect 100 209 101 210 
<< m1 >>
rect 118 209 119 210 
<< m1 >>
rect 130 209 131 210 
<< m1 >>
rect 132 209 133 210 
<< m1 >>
rect 136 209 137 210 
<< m1 >>
rect 145 209 146 210 
<< m1 >>
rect 149 209 150 210 
<< m1 >>
rect 154 209 155 210 
<< m1 >>
rect 163 209 164 210 
<< m1 >>
rect 165 209 166 210 
<< m1 >>
rect 167 209 168 210 
<< m1 >>
rect 172 209 173 210 
<< m1 >>
rect 178 209 179 210 
<< m1 >>
rect 181 209 182 210 
<< m1 >>
rect 183 209 184 210 
<< m1 >>
rect 186 209 187 210 
<< m1 >>
rect 188 209 189 210 
<< m1 >>
rect 190 209 191 210 
<< m1 >>
rect 193 209 194 210 
<< m1 >>
rect 199 209 200 210 
<< m1 >>
rect 201 209 202 210 
<< m1 >>
rect 218 209 219 210 
<< m2 >>
rect 225 209 226 210 
<< m1 >>
rect 226 209 227 210 
<< m1 >>
rect 235 209 236 210 
<< m1 >>
rect 237 209 238 210 
<< m1 >>
rect 241 209 242 210 
<< m1 >>
rect 243 209 244 210 
<< m1 >>
rect 253 209 254 210 
<< m1 >>
rect 256 209 257 210 
<< m1 >>
rect 258 209 259 210 
<< m1 >>
rect 260 209 261 210 
<< m1 >>
rect 262 209 263 210 
<< m1 >>
rect 272 209 273 210 
<< m2 >>
rect 273 209 274 210 
<< m2 >>
rect 297 209 298 210 
<< m1 >>
rect 298 209 299 210 
<< m1 >>
rect 307 209 308 210 
<< m1 >>
rect 322 209 323 210 
<< m1 >>
rect 325 209 326 210 
<< m1 >>
rect 327 209 328 210 
<< m1 >>
rect 329 209 330 210 
<< m1 >>
rect 343 209 344 210 
<< m2 >>
rect 343 209 344 210 
<< m1 >>
rect 345 209 346 210 
<< m1 >>
rect 10 210 11 211 
<< pdiffusion >>
rect 12 210 13 211 
<< m1 >>
rect 13 210 14 211 
<< pdiffusion >>
rect 13 210 14 211 
<< pdiffusion >>
rect 14 210 15 211 
<< pdiffusion >>
rect 15 210 16 211 
<< pdiffusion >>
rect 16 210 17 211 
<< pdiffusion >>
rect 17 210 18 211 
<< m1 >>
rect 19 210 20 211 
<< m2 >>
rect 27 210 28 211 
<< m1 >>
rect 28 210 29 211 
<< pdiffusion >>
rect 30 210 31 211 
<< pdiffusion >>
rect 31 210 32 211 
<< pdiffusion >>
rect 32 210 33 211 
<< pdiffusion >>
rect 33 210 34 211 
<< pdiffusion >>
rect 34 210 35 211 
<< pdiffusion >>
rect 35 210 36 211 
<< m1 >>
rect 37 210 38 211 
<< m2 >>
rect 38 210 39 211 
<< m1 >>
rect 44 210 45 211 
<< m1 >>
rect 46 210 47 211 
<< pdiffusion >>
rect 48 210 49 211 
<< pdiffusion >>
rect 49 210 50 211 
<< pdiffusion >>
rect 50 210 51 211 
<< pdiffusion >>
rect 51 210 52 211 
<< pdiffusion >>
rect 52 210 53 211 
<< pdiffusion >>
rect 53 210 54 211 
<< m1 >>
rect 56 210 57 211 
<< m1 >>
rect 58 210 59 211 
<< m1 >>
rect 62 210 63 211 
<< m1 >>
rect 64 210 65 211 
<< pdiffusion >>
rect 66 210 67 211 
<< pdiffusion >>
rect 67 210 68 211 
<< pdiffusion >>
rect 68 210 69 211 
<< pdiffusion >>
rect 69 210 70 211 
<< pdiffusion >>
rect 70 210 71 211 
<< pdiffusion >>
rect 71 210 72 211 
<< m2 >>
rect 79 210 80 211 
<< m1 >>
rect 80 210 81 211 
<< m1 >>
rect 82 210 83 211 
<< pdiffusion >>
rect 84 210 85 211 
<< pdiffusion >>
rect 85 210 86 211 
<< pdiffusion >>
rect 86 210 87 211 
<< pdiffusion >>
rect 87 210 88 211 
<< pdiffusion >>
rect 88 210 89 211 
<< pdiffusion >>
rect 89 210 90 211 
<< m1 >>
rect 100 210 101 211 
<< pdiffusion >>
rect 102 210 103 211 
<< pdiffusion >>
rect 103 210 104 211 
<< pdiffusion >>
rect 104 210 105 211 
<< pdiffusion >>
rect 105 210 106 211 
<< pdiffusion >>
rect 106 210 107 211 
<< pdiffusion >>
rect 107 210 108 211 
<< m1 >>
rect 118 210 119 211 
<< pdiffusion >>
rect 120 210 121 211 
<< pdiffusion >>
rect 121 210 122 211 
<< pdiffusion >>
rect 122 210 123 211 
<< pdiffusion >>
rect 123 210 124 211 
<< pdiffusion >>
rect 124 210 125 211 
<< pdiffusion >>
rect 125 210 126 211 
<< m1 >>
rect 130 210 131 211 
<< m1 >>
rect 132 210 133 211 
<< m1 >>
rect 136 210 137 211 
<< pdiffusion >>
rect 138 210 139 211 
<< pdiffusion >>
rect 139 210 140 211 
<< pdiffusion >>
rect 140 210 141 211 
<< pdiffusion >>
rect 141 210 142 211 
<< pdiffusion >>
rect 142 210 143 211 
<< pdiffusion >>
rect 143 210 144 211 
<< m1 >>
rect 145 210 146 211 
<< m1 >>
rect 149 210 150 211 
<< m1 >>
rect 154 210 155 211 
<< pdiffusion >>
rect 156 210 157 211 
<< pdiffusion >>
rect 157 210 158 211 
<< pdiffusion >>
rect 158 210 159 211 
<< pdiffusion >>
rect 159 210 160 211 
<< pdiffusion >>
rect 160 210 161 211 
<< pdiffusion >>
rect 161 210 162 211 
<< m1 >>
rect 163 210 164 211 
<< m1 >>
rect 165 210 166 211 
<< m1 >>
rect 167 210 168 211 
<< m1 >>
rect 172 210 173 211 
<< pdiffusion >>
rect 174 210 175 211 
<< pdiffusion >>
rect 175 210 176 211 
<< pdiffusion >>
rect 176 210 177 211 
<< pdiffusion >>
rect 177 210 178 211 
<< m1 >>
rect 178 210 179 211 
<< pdiffusion >>
rect 178 210 179 211 
<< pdiffusion >>
rect 179 210 180 211 
<< m1 >>
rect 181 210 182 211 
<< m1 >>
rect 183 210 184 211 
<< m1 >>
rect 186 210 187 211 
<< m1 >>
rect 188 210 189 211 
<< m1 >>
rect 190 210 191 211 
<< pdiffusion >>
rect 192 210 193 211 
<< m1 >>
rect 193 210 194 211 
<< pdiffusion >>
rect 193 210 194 211 
<< pdiffusion >>
rect 194 210 195 211 
<< pdiffusion >>
rect 195 210 196 211 
<< pdiffusion >>
rect 196 210 197 211 
<< pdiffusion >>
rect 197 210 198 211 
<< m1 >>
rect 199 210 200 211 
<< m1 >>
rect 201 210 202 211 
<< pdiffusion >>
rect 210 210 211 211 
<< pdiffusion >>
rect 211 210 212 211 
<< pdiffusion >>
rect 212 210 213 211 
<< pdiffusion >>
rect 213 210 214 211 
<< pdiffusion >>
rect 214 210 215 211 
<< pdiffusion >>
rect 215 210 216 211 
<< m1 >>
rect 218 210 219 211 
<< m2 >>
rect 225 210 226 211 
<< m1 >>
rect 226 210 227 211 
<< pdiffusion >>
rect 228 210 229 211 
<< pdiffusion >>
rect 229 210 230 211 
<< pdiffusion >>
rect 230 210 231 211 
<< pdiffusion >>
rect 231 210 232 211 
<< pdiffusion >>
rect 232 210 233 211 
<< pdiffusion >>
rect 233 210 234 211 
<< m1 >>
rect 235 210 236 211 
<< m1 >>
rect 237 210 238 211 
<< m1 >>
rect 241 210 242 211 
<< m1 >>
rect 243 210 244 211 
<< pdiffusion >>
rect 246 210 247 211 
<< pdiffusion >>
rect 247 210 248 211 
<< pdiffusion >>
rect 248 210 249 211 
<< pdiffusion >>
rect 249 210 250 211 
<< pdiffusion >>
rect 250 210 251 211 
<< pdiffusion >>
rect 251 210 252 211 
<< m1 >>
rect 253 210 254 211 
<< m1 >>
rect 256 210 257 211 
<< m1 >>
rect 258 210 259 211 
<< m1 >>
rect 260 210 261 211 
<< m1 >>
rect 262 210 263 211 
<< pdiffusion >>
rect 264 210 265 211 
<< pdiffusion >>
rect 265 210 266 211 
<< pdiffusion >>
rect 266 210 267 211 
<< pdiffusion >>
rect 267 210 268 211 
<< pdiffusion >>
rect 268 210 269 211 
<< pdiffusion >>
rect 269 210 270 211 
<< m1 >>
rect 272 210 273 211 
<< m2 >>
rect 273 210 274 211 
<< pdiffusion >>
rect 282 210 283 211 
<< pdiffusion >>
rect 283 210 284 211 
<< pdiffusion >>
rect 284 210 285 211 
<< pdiffusion >>
rect 285 210 286 211 
<< pdiffusion >>
rect 286 210 287 211 
<< pdiffusion >>
rect 287 210 288 211 
<< m2 >>
rect 297 210 298 211 
<< m1 >>
rect 298 210 299 211 
<< pdiffusion >>
rect 300 210 301 211 
<< pdiffusion >>
rect 301 210 302 211 
<< pdiffusion >>
rect 302 210 303 211 
<< pdiffusion >>
rect 303 210 304 211 
<< pdiffusion >>
rect 304 210 305 211 
<< pdiffusion >>
rect 305 210 306 211 
<< m1 >>
rect 307 210 308 211 
<< pdiffusion >>
rect 318 210 319 211 
<< pdiffusion >>
rect 319 210 320 211 
<< pdiffusion >>
rect 320 210 321 211 
<< pdiffusion >>
rect 321 210 322 211 
<< m1 >>
rect 322 210 323 211 
<< pdiffusion >>
rect 322 210 323 211 
<< pdiffusion >>
rect 323 210 324 211 
<< m1 >>
rect 325 210 326 211 
<< m1 >>
rect 327 210 328 211 
<< m1 >>
rect 329 210 330 211 
<< pdiffusion >>
rect 336 210 337 211 
<< pdiffusion >>
rect 337 210 338 211 
<< pdiffusion >>
rect 338 210 339 211 
<< pdiffusion >>
rect 339 210 340 211 
<< pdiffusion >>
rect 340 210 341 211 
<< pdiffusion >>
rect 341 210 342 211 
<< m1 >>
rect 343 210 344 211 
<< m2 >>
rect 343 210 344 211 
<< m1 >>
rect 345 210 346 211 
<< m1 >>
rect 10 211 11 212 
<< pdiffusion >>
rect 12 211 13 212 
<< pdiffusion >>
rect 13 211 14 212 
<< pdiffusion >>
rect 14 211 15 212 
<< pdiffusion >>
rect 15 211 16 212 
<< pdiffusion >>
rect 16 211 17 212 
<< pdiffusion >>
rect 17 211 18 212 
<< m1 >>
rect 19 211 20 212 
<< m2 >>
rect 27 211 28 212 
<< m1 >>
rect 28 211 29 212 
<< pdiffusion >>
rect 30 211 31 212 
<< pdiffusion >>
rect 31 211 32 212 
<< pdiffusion >>
rect 32 211 33 212 
<< pdiffusion >>
rect 33 211 34 212 
<< pdiffusion >>
rect 34 211 35 212 
<< pdiffusion >>
rect 35 211 36 212 
<< m1 >>
rect 37 211 38 212 
<< m2 >>
rect 38 211 39 212 
<< m1 >>
rect 44 211 45 212 
<< m1 >>
rect 46 211 47 212 
<< pdiffusion >>
rect 48 211 49 212 
<< pdiffusion >>
rect 49 211 50 212 
<< pdiffusion >>
rect 50 211 51 212 
<< pdiffusion >>
rect 51 211 52 212 
<< pdiffusion >>
rect 52 211 53 212 
<< pdiffusion >>
rect 53 211 54 212 
<< m1 >>
rect 56 211 57 212 
<< m1 >>
rect 58 211 59 212 
<< m1 >>
rect 62 211 63 212 
<< m1 >>
rect 64 211 65 212 
<< pdiffusion >>
rect 66 211 67 212 
<< pdiffusion >>
rect 67 211 68 212 
<< pdiffusion >>
rect 68 211 69 212 
<< pdiffusion >>
rect 69 211 70 212 
<< pdiffusion >>
rect 70 211 71 212 
<< pdiffusion >>
rect 71 211 72 212 
<< m2 >>
rect 79 211 80 212 
<< m1 >>
rect 80 211 81 212 
<< m1 >>
rect 82 211 83 212 
<< pdiffusion >>
rect 84 211 85 212 
<< pdiffusion >>
rect 85 211 86 212 
<< pdiffusion >>
rect 86 211 87 212 
<< pdiffusion >>
rect 87 211 88 212 
<< pdiffusion >>
rect 88 211 89 212 
<< pdiffusion >>
rect 89 211 90 212 
<< m1 >>
rect 100 211 101 212 
<< pdiffusion >>
rect 102 211 103 212 
<< pdiffusion >>
rect 103 211 104 212 
<< pdiffusion >>
rect 104 211 105 212 
<< pdiffusion >>
rect 105 211 106 212 
<< pdiffusion >>
rect 106 211 107 212 
<< pdiffusion >>
rect 107 211 108 212 
<< m1 >>
rect 118 211 119 212 
<< pdiffusion >>
rect 120 211 121 212 
<< pdiffusion >>
rect 121 211 122 212 
<< pdiffusion >>
rect 122 211 123 212 
<< pdiffusion >>
rect 123 211 124 212 
<< pdiffusion >>
rect 124 211 125 212 
<< pdiffusion >>
rect 125 211 126 212 
<< m1 >>
rect 130 211 131 212 
<< m1 >>
rect 132 211 133 212 
<< m1 >>
rect 136 211 137 212 
<< pdiffusion >>
rect 138 211 139 212 
<< pdiffusion >>
rect 139 211 140 212 
<< pdiffusion >>
rect 140 211 141 212 
<< pdiffusion >>
rect 141 211 142 212 
<< pdiffusion >>
rect 142 211 143 212 
<< pdiffusion >>
rect 143 211 144 212 
<< m1 >>
rect 145 211 146 212 
<< m1 >>
rect 149 211 150 212 
<< m1 >>
rect 154 211 155 212 
<< pdiffusion >>
rect 156 211 157 212 
<< pdiffusion >>
rect 157 211 158 212 
<< pdiffusion >>
rect 158 211 159 212 
<< pdiffusion >>
rect 159 211 160 212 
<< pdiffusion >>
rect 160 211 161 212 
<< pdiffusion >>
rect 161 211 162 212 
<< m1 >>
rect 163 211 164 212 
<< m1 >>
rect 165 211 166 212 
<< m1 >>
rect 167 211 168 212 
<< m1 >>
rect 172 211 173 212 
<< pdiffusion >>
rect 174 211 175 212 
<< pdiffusion >>
rect 175 211 176 212 
<< pdiffusion >>
rect 176 211 177 212 
<< pdiffusion >>
rect 177 211 178 212 
<< pdiffusion >>
rect 178 211 179 212 
<< pdiffusion >>
rect 179 211 180 212 
<< m1 >>
rect 181 211 182 212 
<< m1 >>
rect 183 211 184 212 
<< m1 >>
rect 186 211 187 212 
<< m1 >>
rect 188 211 189 212 
<< m1 >>
rect 190 211 191 212 
<< pdiffusion >>
rect 192 211 193 212 
<< pdiffusion >>
rect 193 211 194 212 
<< pdiffusion >>
rect 194 211 195 212 
<< pdiffusion >>
rect 195 211 196 212 
<< pdiffusion >>
rect 196 211 197 212 
<< pdiffusion >>
rect 197 211 198 212 
<< m1 >>
rect 199 211 200 212 
<< m1 >>
rect 201 211 202 212 
<< pdiffusion >>
rect 210 211 211 212 
<< pdiffusion >>
rect 211 211 212 212 
<< pdiffusion >>
rect 212 211 213 212 
<< pdiffusion >>
rect 213 211 214 212 
<< pdiffusion >>
rect 214 211 215 212 
<< pdiffusion >>
rect 215 211 216 212 
<< m1 >>
rect 218 211 219 212 
<< m2 >>
rect 225 211 226 212 
<< m1 >>
rect 226 211 227 212 
<< pdiffusion >>
rect 228 211 229 212 
<< pdiffusion >>
rect 229 211 230 212 
<< pdiffusion >>
rect 230 211 231 212 
<< pdiffusion >>
rect 231 211 232 212 
<< pdiffusion >>
rect 232 211 233 212 
<< pdiffusion >>
rect 233 211 234 212 
<< m1 >>
rect 235 211 236 212 
<< m1 >>
rect 237 211 238 212 
<< m1 >>
rect 241 211 242 212 
<< m1 >>
rect 243 211 244 212 
<< pdiffusion >>
rect 246 211 247 212 
<< pdiffusion >>
rect 247 211 248 212 
<< pdiffusion >>
rect 248 211 249 212 
<< pdiffusion >>
rect 249 211 250 212 
<< pdiffusion >>
rect 250 211 251 212 
<< pdiffusion >>
rect 251 211 252 212 
<< m1 >>
rect 253 211 254 212 
<< m1 >>
rect 256 211 257 212 
<< m1 >>
rect 258 211 259 212 
<< m1 >>
rect 260 211 261 212 
<< m1 >>
rect 262 211 263 212 
<< pdiffusion >>
rect 264 211 265 212 
<< pdiffusion >>
rect 265 211 266 212 
<< pdiffusion >>
rect 266 211 267 212 
<< pdiffusion >>
rect 267 211 268 212 
<< pdiffusion >>
rect 268 211 269 212 
<< pdiffusion >>
rect 269 211 270 212 
<< m1 >>
rect 272 211 273 212 
<< m2 >>
rect 273 211 274 212 
<< pdiffusion >>
rect 282 211 283 212 
<< pdiffusion >>
rect 283 211 284 212 
<< pdiffusion >>
rect 284 211 285 212 
<< pdiffusion >>
rect 285 211 286 212 
<< pdiffusion >>
rect 286 211 287 212 
<< pdiffusion >>
rect 287 211 288 212 
<< m2 >>
rect 297 211 298 212 
<< m1 >>
rect 298 211 299 212 
<< pdiffusion >>
rect 300 211 301 212 
<< pdiffusion >>
rect 301 211 302 212 
<< pdiffusion >>
rect 302 211 303 212 
<< pdiffusion >>
rect 303 211 304 212 
<< pdiffusion >>
rect 304 211 305 212 
<< pdiffusion >>
rect 305 211 306 212 
<< m1 >>
rect 307 211 308 212 
<< pdiffusion >>
rect 318 211 319 212 
<< pdiffusion >>
rect 319 211 320 212 
<< pdiffusion >>
rect 320 211 321 212 
<< pdiffusion >>
rect 321 211 322 212 
<< pdiffusion >>
rect 322 211 323 212 
<< pdiffusion >>
rect 323 211 324 212 
<< m1 >>
rect 325 211 326 212 
<< m1 >>
rect 327 211 328 212 
<< m1 >>
rect 329 211 330 212 
<< pdiffusion >>
rect 336 211 337 212 
<< pdiffusion >>
rect 337 211 338 212 
<< pdiffusion >>
rect 338 211 339 212 
<< pdiffusion >>
rect 339 211 340 212 
<< pdiffusion >>
rect 340 211 341 212 
<< pdiffusion >>
rect 341 211 342 212 
<< m1 >>
rect 343 211 344 212 
<< m2 >>
rect 343 211 344 212 
<< m1 >>
rect 345 211 346 212 
<< m1 >>
rect 10 212 11 213 
<< pdiffusion >>
rect 12 212 13 213 
<< pdiffusion >>
rect 13 212 14 213 
<< pdiffusion >>
rect 14 212 15 213 
<< pdiffusion >>
rect 15 212 16 213 
<< pdiffusion >>
rect 16 212 17 213 
<< pdiffusion >>
rect 17 212 18 213 
<< m1 >>
rect 19 212 20 213 
<< m2 >>
rect 27 212 28 213 
<< m1 >>
rect 28 212 29 213 
<< pdiffusion >>
rect 30 212 31 213 
<< pdiffusion >>
rect 31 212 32 213 
<< pdiffusion >>
rect 32 212 33 213 
<< pdiffusion >>
rect 33 212 34 213 
<< pdiffusion >>
rect 34 212 35 213 
<< pdiffusion >>
rect 35 212 36 213 
<< m1 >>
rect 37 212 38 213 
<< m2 >>
rect 38 212 39 213 
<< m1 >>
rect 44 212 45 213 
<< m1 >>
rect 46 212 47 213 
<< pdiffusion >>
rect 48 212 49 213 
<< pdiffusion >>
rect 49 212 50 213 
<< pdiffusion >>
rect 50 212 51 213 
<< pdiffusion >>
rect 51 212 52 213 
<< pdiffusion >>
rect 52 212 53 213 
<< pdiffusion >>
rect 53 212 54 213 
<< m1 >>
rect 56 212 57 213 
<< m1 >>
rect 58 212 59 213 
<< m1 >>
rect 62 212 63 213 
<< m1 >>
rect 64 212 65 213 
<< pdiffusion >>
rect 66 212 67 213 
<< pdiffusion >>
rect 67 212 68 213 
<< pdiffusion >>
rect 68 212 69 213 
<< pdiffusion >>
rect 69 212 70 213 
<< pdiffusion >>
rect 70 212 71 213 
<< pdiffusion >>
rect 71 212 72 213 
<< m2 >>
rect 79 212 80 213 
<< m1 >>
rect 80 212 81 213 
<< m1 >>
rect 82 212 83 213 
<< pdiffusion >>
rect 84 212 85 213 
<< pdiffusion >>
rect 85 212 86 213 
<< pdiffusion >>
rect 86 212 87 213 
<< pdiffusion >>
rect 87 212 88 213 
<< pdiffusion >>
rect 88 212 89 213 
<< pdiffusion >>
rect 89 212 90 213 
<< m1 >>
rect 100 212 101 213 
<< pdiffusion >>
rect 102 212 103 213 
<< pdiffusion >>
rect 103 212 104 213 
<< pdiffusion >>
rect 104 212 105 213 
<< pdiffusion >>
rect 105 212 106 213 
<< pdiffusion >>
rect 106 212 107 213 
<< pdiffusion >>
rect 107 212 108 213 
<< m1 >>
rect 118 212 119 213 
<< pdiffusion >>
rect 120 212 121 213 
<< pdiffusion >>
rect 121 212 122 213 
<< pdiffusion >>
rect 122 212 123 213 
<< pdiffusion >>
rect 123 212 124 213 
<< pdiffusion >>
rect 124 212 125 213 
<< pdiffusion >>
rect 125 212 126 213 
<< m1 >>
rect 130 212 131 213 
<< m1 >>
rect 132 212 133 213 
<< m1 >>
rect 136 212 137 213 
<< pdiffusion >>
rect 138 212 139 213 
<< pdiffusion >>
rect 139 212 140 213 
<< pdiffusion >>
rect 140 212 141 213 
<< pdiffusion >>
rect 141 212 142 213 
<< pdiffusion >>
rect 142 212 143 213 
<< pdiffusion >>
rect 143 212 144 213 
<< m1 >>
rect 145 212 146 213 
<< m1 >>
rect 149 212 150 213 
<< m1 >>
rect 154 212 155 213 
<< pdiffusion >>
rect 156 212 157 213 
<< pdiffusion >>
rect 157 212 158 213 
<< pdiffusion >>
rect 158 212 159 213 
<< pdiffusion >>
rect 159 212 160 213 
<< pdiffusion >>
rect 160 212 161 213 
<< pdiffusion >>
rect 161 212 162 213 
<< m1 >>
rect 163 212 164 213 
<< m1 >>
rect 165 212 166 213 
<< m1 >>
rect 167 212 168 213 
<< m1 >>
rect 172 212 173 213 
<< pdiffusion >>
rect 174 212 175 213 
<< pdiffusion >>
rect 175 212 176 213 
<< pdiffusion >>
rect 176 212 177 213 
<< pdiffusion >>
rect 177 212 178 213 
<< pdiffusion >>
rect 178 212 179 213 
<< pdiffusion >>
rect 179 212 180 213 
<< m1 >>
rect 181 212 182 213 
<< m1 >>
rect 183 212 184 213 
<< m1 >>
rect 186 212 187 213 
<< m1 >>
rect 188 212 189 213 
<< m1 >>
rect 190 212 191 213 
<< pdiffusion >>
rect 192 212 193 213 
<< pdiffusion >>
rect 193 212 194 213 
<< pdiffusion >>
rect 194 212 195 213 
<< pdiffusion >>
rect 195 212 196 213 
<< pdiffusion >>
rect 196 212 197 213 
<< pdiffusion >>
rect 197 212 198 213 
<< m1 >>
rect 199 212 200 213 
<< m1 >>
rect 201 212 202 213 
<< pdiffusion >>
rect 210 212 211 213 
<< pdiffusion >>
rect 211 212 212 213 
<< pdiffusion >>
rect 212 212 213 213 
<< pdiffusion >>
rect 213 212 214 213 
<< pdiffusion >>
rect 214 212 215 213 
<< pdiffusion >>
rect 215 212 216 213 
<< m1 >>
rect 218 212 219 213 
<< m2 >>
rect 225 212 226 213 
<< m1 >>
rect 226 212 227 213 
<< pdiffusion >>
rect 228 212 229 213 
<< pdiffusion >>
rect 229 212 230 213 
<< pdiffusion >>
rect 230 212 231 213 
<< pdiffusion >>
rect 231 212 232 213 
<< pdiffusion >>
rect 232 212 233 213 
<< pdiffusion >>
rect 233 212 234 213 
<< m1 >>
rect 235 212 236 213 
<< m1 >>
rect 237 212 238 213 
<< m1 >>
rect 241 212 242 213 
<< m1 >>
rect 243 212 244 213 
<< pdiffusion >>
rect 246 212 247 213 
<< pdiffusion >>
rect 247 212 248 213 
<< pdiffusion >>
rect 248 212 249 213 
<< pdiffusion >>
rect 249 212 250 213 
<< pdiffusion >>
rect 250 212 251 213 
<< pdiffusion >>
rect 251 212 252 213 
<< m1 >>
rect 253 212 254 213 
<< m1 >>
rect 256 212 257 213 
<< m1 >>
rect 258 212 259 213 
<< m1 >>
rect 260 212 261 213 
<< m1 >>
rect 262 212 263 213 
<< pdiffusion >>
rect 264 212 265 213 
<< pdiffusion >>
rect 265 212 266 213 
<< pdiffusion >>
rect 266 212 267 213 
<< pdiffusion >>
rect 267 212 268 213 
<< pdiffusion >>
rect 268 212 269 213 
<< pdiffusion >>
rect 269 212 270 213 
<< m1 >>
rect 272 212 273 213 
<< m2 >>
rect 273 212 274 213 
<< pdiffusion >>
rect 282 212 283 213 
<< pdiffusion >>
rect 283 212 284 213 
<< pdiffusion >>
rect 284 212 285 213 
<< pdiffusion >>
rect 285 212 286 213 
<< pdiffusion >>
rect 286 212 287 213 
<< pdiffusion >>
rect 287 212 288 213 
<< m2 >>
rect 297 212 298 213 
<< m1 >>
rect 298 212 299 213 
<< pdiffusion >>
rect 300 212 301 213 
<< pdiffusion >>
rect 301 212 302 213 
<< pdiffusion >>
rect 302 212 303 213 
<< pdiffusion >>
rect 303 212 304 213 
<< pdiffusion >>
rect 304 212 305 213 
<< pdiffusion >>
rect 305 212 306 213 
<< m1 >>
rect 307 212 308 213 
<< pdiffusion >>
rect 318 212 319 213 
<< pdiffusion >>
rect 319 212 320 213 
<< pdiffusion >>
rect 320 212 321 213 
<< pdiffusion >>
rect 321 212 322 213 
<< pdiffusion >>
rect 322 212 323 213 
<< pdiffusion >>
rect 323 212 324 213 
<< m1 >>
rect 325 212 326 213 
<< m1 >>
rect 327 212 328 213 
<< m1 >>
rect 329 212 330 213 
<< pdiffusion >>
rect 336 212 337 213 
<< pdiffusion >>
rect 337 212 338 213 
<< pdiffusion >>
rect 338 212 339 213 
<< pdiffusion >>
rect 339 212 340 213 
<< pdiffusion >>
rect 340 212 341 213 
<< pdiffusion >>
rect 341 212 342 213 
<< m1 >>
rect 343 212 344 213 
<< m2 >>
rect 343 212 344 213 
<< m1 >>
rect 345 212 346 213 
<< m1 >>
rect 10 213 11 214 
<< pdiffusion >>
rect 12 213 13 214 
<< pdiffusion >>
rect 13 213 14 214 
<< pdiffusion >>
rect 14 213 15 214 
<< pdiffusion >>
rect 15 213 16 214 
<< pdiffusion >>
rect 16 213 17 214 
<< pdiffusion >>
rect 17 213 18 214 
<< m1 >>
rect 19 213 20 214 
<< m2 >>
rect 27 213 28 214 
<< m1 >>
rect 28 213 29 214 
<< pdiffusion >>
rect 30 213 31 214 
<< pdiffusion >>
rect 31 213 32 214 
<< pdiffusion >>
rect 32 213 33 214 
<< pdiffusion >>
rect 33 213 34 214 
<< pdiffusion >>
rect 34 213 35 214 
<< pdiffusion >>
rect 35 213 36 214 
<< m1 >>
rect 37 213 38 214 
<< m2 >>
rect 38 213 39 214 
<< m1 >>
rect 44 213 45 214 
<< m1 >>
rect 46 213 47 214 
<< pdiffusion >>
rect 48 213 49 214 
<< pdiffusion >>
rect 49 213 50 214 
<< pdiffusion >>
rect 50 213 51 214 
<< pdiffusion >>
rect 51 213 52 214 
<< pdiffusion >>
rect 52 213 53 214 
<< pdiffusion >>
rect 53 213 54 214 
<< m1 >>
rect 56 213 57 214 
<< m1 >>
rect 58 213 59 214 
<< m1 >>
rect 62 213 63 214 
<< m1 >>
rect 64 213 65 214 
<< pdiffusion >>
rect 66 213 67 214 
<< pdiffusion >>
rect 67 213 68 214 
<< pdiffusion >>
rect 68 213 69 214 
<< pdiffusion >>
rect 69 213 70 214 
<< pdiffusion >>
rect 70 213 71 214 
<< pdiffusion >>
rect 71 213 72 214 
<< m2 >>
rect 79 213 80 214 
<< m1 >>
rect 80 213 81 214 
<< m1 >>
rect 82 213 83 214 
<< pdiffusion >>
rect 84 213 85 214 
<< pdiffusion >>
rect 85 213 86 214 
<< pdiffusion >>
rect 86 213 87 214 
<< pdiffusion >>
rect 87 213 88 214 
<< pdiffusion >>
rect 88 213 89 214 
<< pdiffusion >>
rect 89 213 90 214 
<< m1 >>
rect 100 213 101 214 
<< pdiffusion >>
rect 102 213 103 214 
<< pdiffusion >>
rect 103 213 104 214 
<< pdiffusion >>
rect 104 213 105 214 
<< pdiffusion >>
rect 105 213 106 214 
<< pdiffusion >>
rect 106 213 107 214 
<< pdiffusion >>
rect 107 213 108 214 
<< m1 >>
rect 118 213 119 214 
<< pdiffusion >>
rect 120 213 121 214 
<< pdiffusion >>
rect 121 213 122 214 
<< pdiffusion >>
rect 122 213 123 214 
<< pdiffusion >>
rect 123 213 124 214 
<< pdiffusion >>
rect 124 213 125 214 
<< pdiffusion >>
rect 125 213 126 214 
<< m1 >>
rect 130 213 131 214 
<< m1 >>
rect 132 213 133 214 
<< m1 >>
rect 136 213 137 214 
<< pdiffusion >>
rect 138 213 139 214 
<< pdiffusion >>
rect 139 213 140 214 
<< pdiffusion >>
rect 140 213 141 214 
<< pdiffusion >>
rect 141 213 142 214 
<< pdiffusion >>
rect 142 213 143 214 
<< pdiffusion >>
rect 143 213 144 214 
<< m1 >>
rect 145 213 146 214 
<< m1 >>
rect 149 213 150 214 
<< m1 >>
rect 154 213 155 214 
<< pdiffusion >>
rect 156 213 157 214 
<< pdiffusion >>
rect 157 213 158 214 
<< pdiffusion >>
rect 158 213 159 214 
<< pdiffusion >>
rect 159 213 160 214 
<< pdiffusion >>
rect 160 213 161 214 
<< pdiffusion >>
rect 161 213 162 214 
<< m1 >>
rect 163 213 164 214 
<< m1 >>
rect 165 213 166 214 
<< m1 >>
rect 167 213 168 214 
<< m1 >>
rect 172 213 173 214 
<< pdiffusion >>
rect 174 213 175 214 
<< pdiffusion >>
rect 175 213 176 214 
<< pdiffusion >>
rect 176 213 177 214 
<< pdiffusion >>
rect 177 213 178 214 
<< pdiffusion >>
rect 178 213 179 214 
<< pdiffusion >>
rect 179 213 180 214 
<< m1 >>
rect 181 213 182 214 
<< m1 >>
rect 183 213 184 214 
<< m1 >>
rect 186 213 187 214 
<< m1 >>
rect 188 213 189 214 
<< m1 >>
rect 190 213 191 214 
<< pdiffusion >>
rect 192 213 193 214 
<< pdiffusion >>
rect 193 213 194 214 
<< pdiffusion >>
rect 194 213 195 214 
<< pdiffusion >>
rect 195 213 196 214 
<< pdiffusion >>
rect 196 213 197 214 
<< pdiffusion >>
rect 197 213 198 214 
<< m1 >>
rect 199 213 200 214 
<< m1 >>
rect 201 213 202 214 
<< pdiffusion >>
rect 210 213 211 214 
<< pdiffusion >>
rect 211 213 212 214 
<< pdiffusion >>
rect 212 213 213 214 
<< pdiffusion >>
rect 213 213 214 214 
<< pdiffusion >>
rect 214 213 215 214 
<< pdiffusion >>
rect 215 213 216 214 
<< m1 >>
rect 218 213 219 214 
<< m2 >>
rect 225 213 226 214 
<< m1 >>
rect 226 213 227 214 
<< pdiffusion >>
rect 228 213 229 214 
<< pdiffusion >>
rect 229 213 230 214 
<< pdiffusion >>
rect 230 213 231 214 
<< pdiffusion >>
rect 231 213 232 214 
<< pdiffusion >>
rect 232 213 233 214 
<< pdiffusion >>
rect 233 213 234 214 
<< m1 >>
rect 235 213 236 214 
<< m1 >>
rect 237 213 238 214 
<< m1 >>
rect 241 213 242 214 
<< m1 >>
rect 243 213 244 214 
<< pdiffusion >>
rect 246 213 247 214 
<< pdiffusion >>
rect 247 213 248 214 
<< pdiffusion >>
rect 248 213 249 214 
<< pdiffusion >>
rect 249 213 250 214 
<< pdiffusion >>
rect 250 213 251 214 
<< pdiffusion >>
rect 251 213 252 214 
<< m1 >>
rect 253 213 254 214 
<< m1 >>
rect 256 213 257 214 
<< m1 >>
rect 258 213 259 214 
<< m1 >>
rect 260 213 261 214 
<< m1 >>
rect 262 213 263 214 
<< pdiffusion >>
rect 264 213 265 214 
<< pdiffusion >>
rect 265 213 266 214 
<< pdiffusion >>
rect 266 213 267 214 
<< pdiffusion >>
rect 267 213 268 214 
<< pdiffusion >>
rect 268 213 269 214 
<< pdiffusion >>
rect 269 213 270 214 
<< m1 >>
rect 272 213 273 214 
<< m2 >>
rect 273 213 274 214 
<< pdiffusion >>
rect 282 213 283 214 
<< pdiffusion >>
rect 283 213 284 214 
<< pdiffusion >>
rect 284 213 285 214 
<< pdiffusion >>
rect 285 213 286 214 
<< pdiffusion >>
rect 286 213 287 214 
<< pdiffusion >>
rect 287 213 288 214 
<< m2 >>
rect 297 213 298 214 
<< m1 >>
rect 298 213 299 214 
<< pdiffusion >>
rect 300 213 301 214 
<< pdiffusion >>
rect 301 213 302 214 
<< pdiffusion >>
rect 302 213 303 214 
<< pdiffusion >>
rect 303 213 304 214 
<< pdiffusion >>
rect 304 213 305 214 
<< pdiffusion >>
rect 305 213 306 214 
<< m1 >>
rect 307 213 308 214 
<< pdiffusion >>
rect 318 213 319 214 
<< pdiffusion >>
rect 319 213 320 214 
<< pdiffusion >>
rect 320 213 321 214 
<< pdiffusion >>
rect 321 213 322 214 
<< pdiffusion >>
rect 322 213 323 214 
<< pdiffusion >>
rect 323 213 324 214 
<< m1 >>
rect 325 213 326 214 
<< m1 >>
rect 327 213 328 214 
<< m1 >>
rect 329 213 330 214 
<< pdiffusion >>
rect 336 213 337 214 
<< pdiffusion >>
rect 337 213 338 214 
<< pdiffusion >>
rect 338 213 339 214 
<< pdiffusion >>
rect 339 213 340 214 
<< pdiffusion >>
rect 340 213 341 214 
<< pdiffusion >>
rect 341 213 342 214 
<< m1 >>
rect 343 213 344 214 
<< m2 >>
rect 343 213 344 214 
<< m1 >>
rect 345 213 346 214 
<< m1 >>
rect 10 214 11 215 
<< pdiffusion >>
rect 12 214 13 215 
<< pdiffusion >>
rect 13 214 14 215 
<< pdiffusion >>
rect 14 214 15 215 
<< pdiffusion >>
rect 15 214 16 215 
<< pdiffusion >>
rect 16 214 17 215 
<< pdiffusion >>
rect 17 214 18 215 
<< m1 >>
rect 19 214 20 215 
<< m2 >>
rect 27 214 28 215 
<< m1 >>
rect 28 214 29 215 
<< pdiffusion >>
rect 30 214 31 215 
<< pdiffusion >>
rect 31 214 32 215 
<< pdiffusion >>
rect 32 214 33 215 
<< pdiffusion >>
rect 33 214 34 215 
<< pdiffusion >>
rect 34 214 35 215 
<< pdiffusion >>
rect 35 214 36 215 
<< m1 >>
rect 37 214 38 215 
<< m2 >>
rect 38 214 39 215 
<< m1 >>
rect 44 214 45 215 
<< m1 >>
rect 46 214 47 215 
<< pdiffusion >>
rect 48 214 49 215 
<< pdiffusion >>
rect 49 214 50 215 
<< pdiffusion >>
rect 50 214 51 215 
<< pdiffusion >>
rect 51 214 52 215 
<< pdiffusion >>
rect 52 214 53 215 
<< pdiffusion >>
rect 53 214 54 215 
<< m1 >>
rect 56 214 57 215 
<< m1 >>
rect 58 214 59 215 
<< m1 >>
rect 62 214 63 215 
<< m1 >>
rect 64 214 65 215 
<< pdiffusion >>
rect 66 214 67 215 
<< pdiffusion >>
rect 67 214 68 215 
<< pdiffusion >>
rect 68 214 69 215 
<< pdiffusion >>
rect 69 214 70 215 
<< pdiffusion >>
rect 70 214 71 215 
<< pdiffusion >>
rect 71 214 72 215 
<< m2 >>
rect 79 214 80 215 
<< m1 >>
rect 80 214 81 215 
<< m1 >>
rect 82 214 83 215 
<< pdiffusion >>
rect 84 214 85 215 
<< pdiffusion >>
rect 85 214 86 215 
<< pdiffusion >>
rect 86 214 87 215 
<< pdiffusion >>
rect 87 214 88 215 
<< pdiffusion >>
rect 88 214 89 215 
<< pdiffusion >>
rect 89 214 90 215 
<< m1 >>
rect 100 214 101 215 
<< pdiffusion >>
rect 102 214 103 215 
<< pdiffusion >>
rect 103 214 104 215 
<< pdiffusion >>
rect 104 214 105 215 
<< pdiffusion >>
rect 105 214 106 215 
<< pdiffusion >>
rect 106 214 107 215 
<< pdiffusion >>
rect 107 214 108 215 
<< m1 >>
rect 118 214 119 215 
<< pdiffusion >>
rect 120 214 121 215 
<< pdiffusion >>
rect 121 214 122 215 
<< pdiffusion >>
rect 122 214 123 215 
<< pdiffusion >>
rect 123 214 124 215 
<< pdiffusion >>
rect 124 214 125 215 
<< pdiffusion >>
rect 125 214 126 215 
<< m1 >>
rect 130 214 131 215 
<< m1 >>
rect 132 214 133 215 
<< m1 >>
rect 136 214 137 215 
<< pdiffusion >>
rect 138 214 139 215 
<< pdiffusion >>
rect 139 214 140 215 
<< pdiffusion >>
rect 140 214 141 215 
<< pdiffusion >>
rect 141 214 142 215 
<< pdiffusion >>
rect 142 214 143 215 
<< pdiffusion >>
rect 143 214 144 215 
<< m1 >>
rect 145 214 146 215 
<< m1 >>
rect 149 214 150 215 
<< m1 >>
rect 154 214 155 215 
<< pdiffusion >>
rect 156 214 157 215 
<< pdiffusion >>
rect 157 214 158 215 
<< pdiffusion >>
rect 158 214 159 215 
<< pdiffusion >>
rect 159 214 160 215 
<< pdiffusion >>
rect 160 214 161 215 
<< pdiffusion >>
rect 161 214 162 215 
<< m1 >>
rect 163 214 164 215 
<< m1 >>
rect 165 214 166 215 
<< m1 >>
rect 167 214 168 215 
<< m1 >>
rect 172 214 173 215 
<< pdiffusion >>
rect 174 214 175 215 
<< pdiffusion >>
rect 175 214 176 215 
<< pdiffusion >>
rect 176 214 177 215 
<< pdiffusion >>
rect 177 214 178 215 
<< pdiffusion >>
rect 178 214 179 215 
<< pdiffusion >>
rect 179 214 180 215 
<< m1 >>
rect 181 214 182 215 
<< m1 >>
rect 183 214 184 215 
<< m1 >>
rect 186 214 187 215 
<< m1 >>
rect 188 214 189 215 
<< m1 >>
rect 190 214 191 215 
<< pdiffusion >>
rect 192 214 193 215 
<< pdiffusion >>
rect 193 214 194 215 
<< pdiffusion >>
rect 194 214 195 215 
<< pdiffusion >>
rect 195 214 196 215 
<< pdiffusion >>
rect 196 214 197 215 
<< pdiffusion >>
rect 197 214 198 215 
<< m1 >>
rect 199 214 200 215 
<< m1 >>
rect 201 214 202 215 
<< pdiffusion >>
rect 210 214 211 215 
<< pdiffusion >>
rect 211 214 212 215 
<< pdiffusion >>
rect 212 214 213 215 
<< pdiffusion >>
rect 213 214 214 215 
<< pdiffusion >>
rect 214 214 215 215 
<< pdiffusion >>
rect 215 214 216 215 
<< m1 >>
rect 218 214 219 215 
<< m2 >>
rect 225 214 226 215 
<< m1 >>
rect 226 214 227 215 
<< pdiffusion >>
rect 228 214 229 215 
<< pdiffusion >>
rect 229 214 230 215 
<< pdiffusion >>
rect 230 214 231 215 
<< pdiffusion >>
rect 231 214 232 215 
<< pdiffusion >>
rect 232 214 233 215 
<< pdiffusion >>
rect 233 214 234 215 
<< m1 >>
rect 235 214 236 215 
<< m1 >>
rect 237 214 238 215 
<< m1 >>
rect 241 214 242 215 
<< m1 >>
rect 243 214 244 215 
<< pdiffusion >>
rect 246 214 247 215 
<< pdiffusion >>
rect 247 214 248 215 
<< pdiffusion >>
rect 248 214 249 215 
<< pdiffusion >>
rect 249 214 250 215 
<< pdiffusion >>
rect 250 214 251 215 
<< pdiffusion >>
rect 251 214 252 215 
<< m1 >>
rect 253 214 254 215 
<< m1 >>
rect 256 214 257 215 
<< m1 >>
rect 258 214 259 215 
<< m1 >>
rect 260 214 261 215 
<< m1 >>
rect 262 214 263 215 
<< pdiffusion >>
rect 264 214 265 215 
<< pdiffusion >>
rect 265 214 266 215 
<< pdiffusion >>
rect 266 214 267 215 
<< pdiffusion >>
rect 267 214 268 215 
<< pdiffusion >>
rect 268 214 269 215 
<< pdiffusion >>
rect 269 214 270 215 
<< m1 >>
rect 272 214 273 215 
<< m2 >>
rect 273 214 274 215 
<< pdiffusion >>
rect 282 214 283 215 
<< pdiffusion >>
rect 283 214 284 215 
<< pdiffusion >>
rect 284 214 285 215 
<< pdiffusion >>
rect 285 214 286 215 
<< pdiffusion >>
rect 286 214 287 215 
<< pdiffusion >>
rect 287 214 288 215 
<< m2 >>
rect 297 214 298 215 
<< m1 >>
rect 298 214 299 215 
<< pdiffusion >>
rect 300 214 301 215 
<< pdiffusion >>
rect 301 214 302 215 
<< pdiffusion >>
rect 302 214 303 215 
<< pdiffusion >>
rect 303 214 304 215 
<< pdiffusion >>
rect 304 214 305 215 
<< pdiffusion >>
rect 305 214 306 215 
<< m1 >>
rect 307 214 308 215 
<< pdiffusion >>
rect 318 214 319 215 
<< pdiffusion >>
rect 319 214 320 215 
<< pdiffusion >>
rect 320 214 321 215 
<< pdiffusion >>
rect 321 214 322 215 
<< pdiffusion >>
rect 322 214 323 215 
<< pdiffusion >>
rect 323 214 324 215 
<< m1 >>
rect 325 214 326 215 
<< m1 >>
rect 327 214 328 215 
<< m1 >>
rect 329 214 330 215 
<< pdiffusion >>
rect 336 214 337 215 
<< pdiffusion >>
rect 337 214 338 215 
<< pdiffusion >>
rect 338 214 339 215 
<< pdiffusion >>
rect 339 214 340 215 
<< pdiffusion >>
rect 340 214 341 215 
<< pdiffusion >>
rect 341 214 342 215 
<< m1 >>
rect 343 214 344 215 
<< m2 >>
rect 343 214 344 215 
<< m1 >>
rect 345 214 346 215 
<< m1 >>
rect 10 215 11 216 
<< pdiffusion >>
rect 12 215 13 216 
<< m1 >>
rect 13 215 14 216 
<< pdiffusion >>
rect 13 215 14 216 
<< pdiffusion >>
rect 14 215 15 216 
<< pdiffusion >>
rect 15 215 16 216 
<< pdiffusion >>
rect 16 215 17 216 
<< pdiffusion >>
rect 17 215 18 216 
<< m1 >>
rect 19 215 20 216 
<< m2 >>
rect 27 215 28 216 
<< m1 >>
rect 28 215 29 216 
<< pdiffusion >>
rect 30 215 31 216 
<< pdiffusion >>
rect 31 215 32 216 
<< pdiffusion >>
rect 32 215 33 216 
<< pdiffusion >>
rect 33 215 34 216 
<< pdiffusion >>
rect 34 215 35 216 
<< pdiffusion >>
rect 35 215 36 216 
<< m1 >>
rect 37 215 38 216 
<< m2 >>
rect 38 215 39 216 
<< m1 >>
rect 44 215 45 216 
<< m1 >>
rect 46 215 47 216 
<< pdiffusion >>
rect 48 215 49 216 
<< pdiffusion >>
rect 49 215 50 216 
<< pdiffusion >>
rect 50 215 51 216 
<< pdiffusion >>
rect 51 215 52 216 
<< pdiffusion >>
rect 52 215 53 216 
<< pdiffusion >>
rect 53 215 54 216 
<< m1 >>
rect 56 215 57 216 
<< m1 >>
rect 58 215 59 216 
<< m1 >>
rect 62 215 63 216 
<< m1 >>
rect 64 215 65 216 
<< pdiffusion >>
rect 66 215 67 216 
<< pdiffusion >>
rect 67 215 68 216 
<< pdiffusion >>
rect 68 215 69 216 
<< pdiffusion >>
rect 69 215 70 216 
<< m1 >>
rect 70 215 71 216 
<< pdiffusion >>
rect 70 215 71 216 
<< pdiffusion >>
rect 71 215 72 216 
<< m2 >>
rect 79 215 80 216 
<< m1 >>
rect 80 215 81 216 
<< m1 >>
rect 82 215 83 216 
<< pdiffusion >>
rect 84 215 85 216 
<< pdiffusion >>
rect 85 215 86 216 
<< pdiffusion >>
rect 86 215 87 216 
<< pdiffusion >>
rect 87 215 88 216 
<< pdiffusion >>
rect 88 215 89 216 
<< pdiffusion >>
rect 89 215 90 216 
<< m1 >>
rect 100 215 101 216 
<< pdiffusion >>
rect 102 215 103 216 
<< pdiffusion >>
rect 103 215 104 216 
<< pdiffusion >>
rect 104 215 105 216 
<< pdiffusion >>
rect 105 215 106 216 
<< m1 >>
rect 106 215 107 216 
<< pdiffusion >>
rect 106 215 107 216 
<< pdiffusion >>
rect 107 215 108 216 
<< m1 >>
rect 118 215 119 216 
<< pdiffusion >>
rect 120 215 121 216 
<< pdiffusion >>
rect 121 215 122 216 
<< pdiffusion >>
rect 122 215 123 216 
<< pdiffusion >>
rect 123 215 124 216 
<< pdiffusion >>
rect 124 215 125 216 
<< pdiffusion >>
rect 125 215 126 216 
<< m1 >>
rect 130 215 131 216 
<< m1 >>
rect 132 215 133 216 
<< m1 >>
rect 136 215 137 216 
<< pdiffusion >>
rect 138 215 139 216 
<< pdiffusion >>
rect 139 215 140 216 
<< pdiffusion >>
rect 140 215 141 216 
<< pdiffusion >>
rect 141 215 142 216 
<< pdiffusion >>
rect 142 215 143 216 
<< pdiffusion >>
rect 143 215 144 216 
<< m1 >>
rect 145 215 146 216 
<< m1 >>
rect 149 215 150 216 
<< m1 >>
rect 154 215 155 216 
<< pdiffusion >>
rect 156 215 157 216 
<< pdiffusion >>
rect 157 215 158 216 
<< pdiffusion >>
rect 158 215 159 216 
<< pdiffusion >>
rect 159 215 160 216 
<< pdiffusion >>
rect 160 215 161 216 
<< pdiffusion >>
rect 161 215 162 216 
<< m1 >>
rect 163 215 164 216 
<< m1 >>
rect 165 215 166 216 
<< m1 >>
rect 167 215 168 216 
<< m1 >>
rect 172 215 173 216 
<< pdiffusion >>
rect 174 215 175 216 
<< pdiffusion >>
rect 175 215 176 216 
<< pdiffusion >>
rect 176 215 177 216 
<< pdiffusion >>
rect 177 215 178 216 
<< pdiffusion >>
rect 178 215 179 216 
<< pdiffusion >>
rect 179 215 180 216 
<< m1 >>
rect 181 215 182 216 
<< m1 >>
rect 183 215 184 216 
<< m1 >>
rect 186 215 187 216 
<< m1 >>
rect 188 215 189 216 
<< m1 >>
rect 190 215 191 216 
<< pdiffusion >>
rect 192 215 193 216 
<< pdiffusion >>
rect 193 215 194 216 
<< pdiffusion >>
rect 194 215 195 216 
<< pdiffusion >>
rect 195 215 196 216 
<< m1 >>
rect 196 215 197 216 
<< pdiffusion >>
rect 196 215 197 216 
<< pdiffusion >>
rect 197 215 198 216 
<< m1 >>
rect 199 215 200 216 
<< m1 >>
rect 201 215 202 216 
<< pdiffusion >>
rect 210 215 211 216 
<< m1 >>
rect 211 215 212 216 
<< pdiffusion >>
rect 211 215 212 216 
<< pdiffusion >>
rect 212 215 213 216 
<< pdiffusion >>
rect 213 215 214 216 
<< m1 >>
rect 214 215 215 216 
<< pdiffusion >>
rect 214 215 215 216 
<< pdiffusion >>
rect 215 215 216 216 
<< m1 >>
rect 218 215 219 216 
<< m2 >>
rect 225 215 226 216 
<< m1 >>
rect 226 215 227 216 
<< pdiffusion >>
rect 228 215 229 216 
<< pdiffusion >>
rect 229 215 230 216 
<< pdiffusion >>
rect 230 215 231 216 
<< pdiffusion >>
rect 231 215 232 216 
<< pdiffusion >>
rect 232 215 233 216 
<< pdiffusion >>
rect 233 215 234 216 
<< m1 >>
rect 235 215 236 216 
<< m1 >>
rect 237 215 238 216 
<< m1 >>
rect 241 215 242 216 
<< m1 >>
rect 243 215 244 216 
<< pdiffusion >>
rect 246 215 247 216 
<< pdiffusion >>
rect 247 215 248 216 
<< pdiffusion >>
rect 248 215 249 216 
<< pdiffusion >>
rect 249 215 250 216 
<< m1 >>
rect 250 215 251 216 
<< pdiffusion >>
rect 250 215 251 216 
<< pdiffusion >>
rect 251 215 252 216 
<< m1 >>
rect 253 215 254 216 
<< m2 >>
rect 253 215 254 216 
<< m2c >>
rect 253 215 254 216 
<< m1 >>
rect 253 215 254 216 
<< m2 >>
rect 253 215 254 216 
<< m1 >>
rect 256 215 257 216 
<< m1 >>
rect 258 215 259 216 
<< m1 >>
rect 260 215 261 216 
<< m1 >>
rect 262 215 263 216 
<< pdiffusion >>
rect 264 215 265 216 
<< pdiffusion >>
rect 265 215 266 216 
<< pdiffusion >>
rect 266 215 267 216 
<< pdiffusion >>
rect 267 215 268 216 
<< pdiffusion >>
rect 268 215 269 216 
<< pdiffusion >>
rect 269 215 270 216 
<< m1 >>
rect 272 215 273 216 
<< m2 >>
rect 273 215 274 216 
<< pdiffusion >>
rect 282 215 283 216 
<< pdiffusion >>
rect 283 215 284 216 
<< pdiffusion >>
rect 284 215 285 216 
<< pdiffusion >>
rect 285 215 286 216 
<< m1 >>
rect 286 215 287 216 
<< pdiffusion >>
rect 286 215 287 216 
<< pdiffusion >>
rect 287 215 288 216 
<< m2 >>
rect 297 215 298 216 
<< m1 >>
rect 298 215 299 216 
<< pdiffusion >>
rect 300 215 301 216 
<< m1 >>
rect 301 215 302 216 
<< pdiffusion >>
rect 301 215 302 216 
<< pdiffusion >>
rect 302 215 303 216 
<< pdiffusion >>
rect 303 215 304 216 
<< pdiffusion >>
rect 304 215 305 216 
<< pdiffusion >>
rect 305 215 306 216 
<< m1 >>
rect 307 215 308 216 
<< pdiffusion >>
rect 318 215 319 216 
<< pdiffusion >>
rect 319 215 320 216 
<< pdiffusion >>
rect 320 215 321 216 
<< pdiffusion >>
rect 321 215 322 216 
<< m1 >>
rect 322 215 323 216 
<< pdiffusion >>
rect 322 215 323 216 
<< pdiffusion >>
rect 323 215 324 216 
<< m1 >>
rect 325 215 326 216 
<< m1 >>
rect 327 215 328 216 
<< m1 >>
rect 329 215 330 216 
<< pdiffusion >>
rect 336 215 337 216 
<< pdiffusion >>
rect 337 215 338 216 
<< pdiffusion >>
rect 338 215 339 216 
<< pdiffusion >>
rect 339 215 340 216 
<< pdiffusion >>
rect 340 215 341 216 
<< pdiffusion >>
rect 341 215 342 216 
<< m1 >>
rect 343 215 344 216 
<< m2 >>
rect 343 215 344 216 
<< m1 >>
rect 345 215 346 216 
<< m1 >>
rect 10 216 11 217 
<< m1 >>
rect 13 216 14 217 
<< m1 >>
rect 19 216 20 217 
<< m2 >>
rect 27 216 28 217 
<< m1 >>
rect 28 216 29 217 
<< m1 >>
rect 37 216 38 217 
<< m2 >>
rect 38 216 39 217 
<< m1 >>
rect 44 216 45 217 
<< m1 >>
rect 46 216 47 217 
<< m1 >>
rect 56 216 57 217 
<< m1 >>
rect 58 216 59 217 
<< m1 >>
rect 62 216 63 217 
<< m1 >>
rect 64 216 65 217 
<< m1 >>
rect 70 216 71 217 
<< m2 >>
rect 79 216 80 217 
<< m1 >>
rect 80 216 81 217 
<< m1 >>
rect 82 216 83 217 
<< m1 >>
rect 100 216 101 217 
<< m1 >>
rect 106 216 107 217 
<< m1 >>
rect 118 216 119 217 
<< m1 >>
rect 130 216 131 217 
<< m1 >>
rect 132 216 133 217 
<< m1 >>
rect 136 216 137 217 
<< m1 >>
rect 145 216 146 217 
<< m1 >>
rect 149 216 150 217 
<< m1 >>
rect 154 216 155 217 
<< m1 >>
rect 163 216 164 217 
<< m1 >>
rect 165 216 166 217 
<< m1 >>
rect 167 216 168 217 
<< m1 >>
rect 172 216 173 217 
<< m1 >>
rect 181 216 182 217 
<< m1 >>
rect 183 216 184 217 
<< m1 >>
rect 186 216 187 217 
<< m1 >>
rect 188 216 189 217 
<< m1 >>
rect 190 216 191 217 
<< m1 >>
rect 196 216 197 217 
<< m1 >>
rect 199 216 200 217 
<< m1 >>
rect 201 216 202 217 
<< m1 >>
rect 211 216 212 217 
<< m1 >>
rect 214 216 215 217 
<< m2 >>
rect 214 216 215 217 
<< m2c >>
rect 214 216 215 217 
<< m1 >>
rect 214 216 215 217 
<< m2 >>
rect 214 216 215 217 
<< m1 >>
rect 218 216 219 217 
<< m2 >>
rect 225 216 226 217 
<< m1 >>
rect 226 216 227 217 
<< m1 >>
rect 235 216 236 217 
<< m1 >>
rect 237 216 238 217 
<< m1 >>
rect 241 216 242 217 
<< m1 >>
rect 243 216 244 217 
<< m1 >>
rect 250 216 251 217 
<< m2 >>
rect 253 216 254 217 
<< m1 >>
rect 256 216 257 217 
<< m1 >>
rect 258 216 259 217 
<< m1 >>
rect 260 216 261 217 
<< m1 >>
rect 262 216 263 217 
<< m1 >>
rect 272 216 273 217 
<< m2 >>
rect 273 216 274 217 
<< m1 >>
rect 286 216 287 217 
<< m2 >>
rect 297 216 298 217 
<< m1 >>
rect 298 216 299 217 
<< m1 >>
rect 301 216 302 217 
<< m1 >>
rect 307 216 308 217 
<< m1 >>
rect 322 216 323 217 
<< m1 >>
rect 325 216 326 217 
<< m1 >>
rect 327 216 328 217 
<< m1 >>
rect 329 216 330 217 
<< m1 >>
rect 343 216 344 217 
<< m2 >>
rect 343 216 344 217 
<< m1 >>
rect 345 216 346 217 
<< m1 >>
rect 10 217 11 218 
<< m1 >>
rect 13 217 14 218 
<< m1 >>
rect 19 217 20 218 
<< m2 >>
rect 27 217 28 218 
<< m1 >>
rect 28 217 29 218 
<< m1 >>
rect 29 217 30 218 
<< m1 >>
rect 35 217 36 218 
<< m2 >>
rect 35 217 36 218 
<< m2c >>
rect 35 217 36 218 
<< m1 >>
rect 35 217 36 218 
<< m2 >>
rect 35 217 36 218 
<< m2 >>
rect 36 217 37 218 
<< m1 >>
rect 37 217 38 218 
<< m2 >>
rect 37 217 38 218 
<< m2 >>
rect 38 217 39 218 
<< m1 >>
rect 44 217 45 218 
<< m1 >>
rect 46 217 47 218 
<< m1 >>
rect 56 217 57 218 
<< m1 >>
rect 58 217 59 218 
<< m1 >>
rect 62 217 63 218 
<< m1 >>
rect 64 217 65 218 
<< m1 >>
rect 70 217 71 218 
<< m2 >>
rect 79 217 80 218 
<< m1 >>
rect 80 217 81 218 
<< m2 >>
rect 80 217 81 218 
<< m2 >>
rect 81 217 82 218 
<< m1 >>
rect 82 217 83 218 
<< m2 >>
rect 82 217 83 218 
<< m2 >>
rect 83 217 84 218 
<< m1 >>
rect 84 217 85 218 
<< m2 >>
rect 84 217 85 218 
<< m2c >>
rect 84 217 85 218 
<< m1 >>
rect 84 217 85 218 
<< m2 >>
rect 84 217 85 218 
<< m1 >>
rect 100 217 101 218 
<< m1 >>
rect 106 217 107 218 
<< m1 >>
rect 118 217 119 218 
<< m1 >>
rect 130 217 131 218 
<< m1 >>
rect 132 217 133 218 
<< m1 >>
rect 136 217 137 218 
<< m1 >>
rect 145 217 146 218 
<< m1 >>
rect 149 217 150 218 
<< m1 >>
rect 154 217 155 218 
<< m1 >>
rect 163 217 164 218 
<< m1 >>
rect 165 217 166 218 
<< m1 >>
rect 167 217 168 218 
<< m1 >>
rect 172 217 173 218 
<< m1 >>
rect 181 217 182 218 
<< m1 >>
rect 183 217 184 218 
<< m1 >>
rect 186 217 187 218 
<< m1 >>
rect 188 217 189 218 
<< m1 >>
rect 190 217 191 218 
<< m1 >>
rect 196 217 197 218 
<< m1 >>
rect 199 217 200 218 
<< m1 >>
rect 201 217 202 218 
<< m1 >>
rect 211 217 212 218 
<< m2 >>
rect 214 217 215 218 
<< m1 >>
rect 218 217 219 218 
<< m2 >>
rect 225 217 226 218 
<< m1 >>
rect 226 217 227 218 
<< m2 >>
rect 226 217 227 218 
<< m2 >>
rect 227 217 228 218 
<< m1 >>
rect 228 217 229 218 
<< m2 >>
rect 228 217 229 218 
<< m2c >>
rect 228 217 229 218 
<< m1 >>
rect 228 217 229 218 
<< m2 >>
rect 228 217 229 218 
<< m1 >>
rect 235 217 236 218 
<< m1 >>
rect 237 217 238 218 
<< m1 >>
rect 241 217 242 218 
<< m1 >>
rect 243 217 244 218 
<< m1 >>
rect 250 217 251 218 
<< m1 >>
rect 251 217 252 218 
<< m1 >>
rect 252 217 253 218 
<< m1 >>
rect 253 217 254 218 
<< m2 >>
rect 253 217 254 218 
<< m1 >>
rect 254 217 255 218 
<< m1 >>
rect 255 217 256 218 
<< m1 >>
rect 256 217 257 218 
<< m1 >>
rect 258 217 259 218 
<< m1 >>
rect 260 217 261 218 
<< m1 >>
rect 262 217 263 218 
<< m1 >>
rect 272 217 273 218 
<< m2 >>
rect 273 217 274 218 
<< m1 >>
rect 286 217 287 218 
<< m1 >>
rect 287 217 288 218 
<< m1 >>
rect 288 217 289 218 
<< m1 >>
rect 289 217 290 218 
<< m1 >>
rect 290 217 291 218 
<< m1 >>
rect 291 217 292 218 
<< m1 >>
rect 292 217 293 218 
<< m1 >>
rect 293 217 294 218 
<< m1 >>
rect 294 217 295 218 
<< m1 >>
rect 295 217 296 218 
<< m1 >>
rect 296 217 297 218 
<< m2 >>
rect 296 217 297 218 
<< m2c >>
rect 296 217 297 218 
<< m1 >>
rect 296 217 297 218 
<< m2 >>
rect 296 217 297 218 
<< m2 >>
rect 297 217 298 218 
<< m1 >>
rect 298 217 299 218 
<< m1 >>
rect 301 217 302 218 
<< m1 >>
rect 302 217 303 218 
<< m1 >>
rect 305 217 306 218 
<< m2 >>
rect 305 217 306 218 
<< m2c >>
rect 305 217 306 218 
<< m1 >>
rect 305 217 306 218 
<< m2 >>
rect 305 217 306 218 
<< m2 >>
rect 306 217 307 218 
<< m1 >>
rect 307 217 308 218 
<< m2 >>
rect 307 217 308 218 
<< m2 >>
rect 308 217 309 218 
<< m1 >>
rect 309 217 310 218 
<< m2 >>
rect 309 217 310 218 
<< m2c >>
rect 309 217 310 218 
<< m1 >>
rect 309 217 310 218 
<< m2 >>
rect 309 217 310 218 
<< m1 >>
rect 310 217 311 218 
<< m1 >>
rect 311 217 312 218 
<< m1 >>
rect 312 217 313 218 
<< m1 >>
rect 313 217 314 218 
<< m1 >>
rect 314 217 315 218 
<< m1 >>
rect 315 217 316 218 
<< m1 >>
rect 316 217 317 218 
<< m1 >>
rect 317 217 318 218 
<< m1 >>
rect 318 217 319 218 
<< m1 >>
rect 322 217 323 218 
<< m1 >>
rect 325 217 326 218 
<< m1 >>
rect 327 217 328 218 
<< m1 >>
rect 329 217 330 218 
<< m1 >>
rect 343 217 344 218 
<< m2 >>
rect 343 217 344 218 
<< m1 >>
rect 345 217 346 218 
<< m1 >>
rect 10 218 11 219 
<< m1 >>
rect 13 218 14 219 
<< m1 >>
rect 14 218 15 219 
<< m1 >>
rect 15 218 16 219 
<< m1 >>
rect 16 218 17 219 
<< m1 >>
rect 17 218 18 219 
<< m1 >>
rect 18 218 19 219 
<< m1 >>
rect 19 218 20 219 
<< m2 >>
rect 27 218 28 219 
<< m1 >>
rect 29 218 30 219 
<< m2 >>
rect 29 218 30 219 
<< m2c >>
rect 29 218 30 219 
<< m1 >>
rect 29 218 30 219 
<< m2 >>
rect 29 218 30 219 
<< m1 >>
rect 35 218 36 219 
<< m1 >>
rect 37 218 38 219 
<< m1 >>
rect 44 218 45 219 
<< m1 >>
rect 46 218 47 219 
<< m1 >>
rect 56 218 57 219 
<< m1 >>
rect 58 218 59 219 
<< m1 >>
rect 62 218 63 219 
<< m1 >>
rect 64 218 65 219 
<< m1 >>
rect 70 218 71 219 
<< m1 >>
rect 80 218 81 219 
<< m1 >>
rect 82 218 83 219 
<< m1 >>
rect 84 218 85 219 
<< m1 >>
rect 100 218 101 219 
<< m2 >>
rect 100 218 101 219 
<< m2c >>
rect 100 218 101 219 
<< m1 >>
rect 100 218 101 219 
<< m2 >>
rect 100 218 101 219 
<< m1 >>
rect 106 218 107 219 
<< m1 >>
rect 118 218 119 219 
<< m1 >>
rect 130 218 131 219 
<< m1 >>
rect 132 218 133 219 
<< m1 >>
rect 136 218 137 219 
<< m1 >>
rect 140 218 141 219 
<< m2 >>
rect 140 218 141 219 
<< m2c >>
rect 140 218 141 219 
<< m1 >>
rect 140 218 141 219 
<< m2 >>
rect 140 218 141 219 
<< m1 >>
rect 141 218 142 219 
<< m1 >>
rect 142 218 143 219 
<< m1 >>
rect 143 218 144 219 
<< m2 >>
rect 143 218 144 219 
<< m2c >>
rect 143 218 144 219 
<< m1 >>
rect 143 218 144 219 
<< m2 >>
rect 143 218 144 219 
<< m2 >>
rect 144 218 145 219 
<< m1 >>
rect 145 218 146 219 
<< m2 >>
rect 145 218 146 219 
<< m2 >>
rect 146 218 147 219 
<< m1 >>
rect 147 218 148 219 
<< m2 >>
rect 147 218 148 219 
<< m2c >>
rect 147 218 148 219 
<< m1 >>
rect 147 218 148 219 
<< m2 >>
rect 147 218 148 219 
<< m1 >>
rect 148 218 149 219 
<< m1 >>
rect 149 218 150 219 
<< m1 >>
rect 154 218 155 219 
<< m2 >>
rect 154 218 155 219 
<< m2c >>
rect 154 218 155 219 
<< m1 >>
rect 154 218 155 219 
<< m2 >>
rect 154 218 155 219 
<< m1 >>
rect 163 218 164 219 
<< m1 >>
rect 165 218 166 219 
<< m1 >>
rect 167 218 168 219 
<< m1 >>
rect 172 218 173 219 
<< m2 >>
rect 172 218 173 219 
<< m2c >>
rect 172 218 173 219 
<< m1 >>
rect 172 218 173 219 
<< m2 >>
rect 172 218 173 219 
<< m1 >>
rect 181 218 182 219 
<< m2 >>
rect 181 218 182 219 
<< m2c >>
rect 181 218 182 219 
<< m1 >>
rect 181 218 182 219 
<< m2 >>
rect 181 218 182 219 
<< m1 >>
rect 183 218 184 219 
<< m2 >>
rect 183 218 184 219 
<< m2c >>
rect 183 218 184 219 
<< m1 >>
rect 183 218 184 219 
<< m2 >>
rect 183 218 184 219 
<< m1 >>
rect 186 218 187 219 
<< m2 >>
rect 186 218 187 219 
<< m2c >>
rect 186 218 187 219 
<< m1 >>
rect 186 218 187 219 
<< m2 >>
rect 186 218 187 219 
<< m1 >>
rect 188 218 189 219 
<< m2 >>
rect 188 218 189 219 
<< m2c >>
rect 188 218 189 219 
<< m1 >>
rect 188 218 189 219 
<< m2 >>
rect 188 218 189 219 
<< m1 >>
rect 190 218 191 219 
<< m2 >>
rect 190 218 191 219 
<< m2c >>
rect 190 218 191 219 
<< m1 >>
rect 190 218 191 219 
<< m2 >>
rect 190 218 191 219 
<< m1 >>
rect 196 218 197 219 
<< m1 >>
rect 199 218 200 219 
<< m1 >>
rect 201 218 202 219 
<< m1 >>
rect 211 218 212 219 
<< m1 >>
rect 212 218 213 219 
<< m1 >>
rect 213 218 214 219 
<< m1 >>
rect 214 218 215 219 
<< m2 >>
rect 214 218 215 219 
<< m1 >>
rect 215 218 216 219 
<< m1 >>
rect 216 218 217 219 
<< m1 >>
rect 218 218 219 219 
<< m1 >>
rect 226 218 227 219 
<< m1 >>
rect 228 218 229 219 
<< m1 >>
rect 235 218 236 219 
<< m1 >>
rect 237 218 238 219 
<< m1 >>
rect 241 218 242 219 
<< m1 >>
rect 243 218 244 219 
<< m2 >>
rect 253 218 254 219 
<< m1 >>
rect 258 218 259 219 
<< m1 >>
rect 260 218 261 219 
<< m1 >>
rect 262 218 263 219 
<< m1 >>
rect 272 218 273 219 
<< m2 >>
rect 273 218 274 219 
<< m1 >>
rect 298 218 299 219 
<< m1 >>
rect 302 218 303 219 
<< m1 >>
rect 303 218 304 219 
<< m1 >>
rect 304 218 305 219 
<< m1 >>
rect 305 218 306 219 
<< m1 >>
rect 307 218 308 219 
<< m1 >>
rect 318 218 319 219 
<< m1 >>
rect 322 218 323 219 
<< m1 >>
rect 325 218 326 219 
<< m1 >>
rect 327 218 328 219 
<< m1 >>
rect 329 218 330 219 
<< m1 >>
rect 343 218 344 219 
<< m2 >>
rect 343 218 344 219 
<< m1 >>
rect 345 218 346 219 
<< m1 >>
rect 10 219 11 220 
<< m1 >>
rect 27 219 28 220 
<< m2 >>
rect 27 219 28 220 
<< m2c >>
rect 27 219 28 220 
<< m1 >>
rect 27 219 28 220 
<< m2 >>
rect 27 219 28 220 
<< m2 >>
rect 29 219 30 220 
<< m1 >>
rect 35 219 36 220 
<< m1 >>
rect 37 219 38 220 
<< m1 >>
rect 44 219 45 220 
<< m1 >>
rect 46 219 47 220 
<< m1 >>
rect 56 219 57 220 
<< m1 >>
rect 58 219 59 220 
<< m1 >>
rect 62 219 63 220 
<< m1 >>
rect 64 219 65 220 
<< m1 >>
rect 70 219 71 220 
<< m1 >>
rect 80 219 81 220 
<< m1 >>
rect 82 219 83 220 
<< m1 >>
rect 84 219 85 220 
<< m2 >>
rect 100 219 101 220 
<< m1 >>
rect 106 219 107 220 
<< m1 >>
rect 118 219 119 220 
<< m1 >>
rect 130 219 131 220 
<< m1 >>
rect 132 219 133 220 
<< m1 >>
rect 136 219 137 220 
<< m2 >>
rect 140 219 141 220 
<< m1 >>
rect 145 219 146 220 
<< m2 >>
rect 154 219 155 220 
<< m1 >>
rect 163 219 164 220 
<< m1 >>
rect 165 219 166 220 
<< m1 >>
rect 167 219 168 220 
<< m2 >>
rect 172 219 173 220 
<< m2 >>
rect 181 219 182 220 
<< m2 >>
rect 183 219 184 220 
<< m2 >>
rect 186 219 187 220 
<< m2 >>
rect 188 219 189 220 
<< m2 >>
rect 190 219 191 220 
<< m1 >>
rect 196 219 197 220 
<< m1 >>
rect 199 219 200 220 
<< m1 >>
rect 201 219 202 220 
<< m2 >>
rect 212 219 213 220 
<< m2 >>
rect 213 219 214 220 
<< m2 >>
rect 214 219 215 220 
<< m1 >>
rect 216 219 217 220 
<< m1 >>
rect 218 219 219 220 
<< m1 >>
rect 226 219 227 220 
<< m1 >>
rect 228 219 229 220 
<< m1 >>
rect 235 219 236 220 
<< m1 >>
rect 237 219 238 220 
<< m1 >>
rect 241 219 242 220 
<< m1 >>
rect 243 219 244 220 
<< m1 >>
rect 253 219 254 220 
<< m2 >>
rect 253 219 254 220 
<< m2c >>
rect 253 219 254 220 
<< m1 >>
rect 253 219 254 220 
<< m2 >>
rect 253 219 254 220 
<< m1 >>
rect 258 219 259 220 
<< m2 >>
rect 258 219 259 220 
<< m2c >>
rect 258 219 259 220 
<< m1 >>
rect 258 219 259 220 
<< m2 >>
rect 258 219 259 220 
<< m2 >>
rect 259 219 260 220 
<< m1 >>
rect 260 219 261 220 
<< m2 >>
rect 260 219 261 220 
<< m2 >>
rect 261 219 262 220 
<< m1 >>
rect 262 219 263 220 
<< m2 >>
rect 262 219 263 220 
<< m2 >>
rect 263 219 264 220 
<< m1 >>
rect 264 219 265 220 
<< m2 >>
rect 264 219 265 220 
<< m2c >>
rect 264 219 265 220 
<< m1 >>
rect 264 219 265 220 
<< m2 >>
rect 264 219 265 220 
<< m1 >>
rect 272 219 273 220 
<< m2 >>
rect 273 219 274 220 
<< m1 >>
rect 274 219 275 220 
<< m2 >>
rect 274 219 275 220 
<< m2c >>
rect 274 219 275 220 
<< m1 >>
rect 274 219 275 220 
<< m2 >>
rect 274 219 275 220 
<< m1 >>
rect 275 219 276 220 
<< m1 >>
rect 276 219 277 220 
<< m1 >>
rect 277 219 278 220 
<< m1 >>
rect 278 219 279 220 
<< m1 >>
rect 279 219 280 220 
<< m1 >>
rect 280 219 281 220 
<< m1 >>
rect 281 219 282 220 
<< m1 >>
rect 282 219 283 220 
<< m2 >>
rect 282 219 283 220 
<< m2c >>
rect 282 219 283 220 
<< m1 >>
rect 282 219 283 220 
<< m2 >>
rect 282 219 283 220 
<< m1 >>
rect 298 219 299 220 
<< m1 >>
rect 299 219 300 220 
<< m1 >>
rect 300 219 301 220 
<< m2 >>
rect 300 219 301 220 
<< m2c >>
rect 300 219 301 220 
<< m1 >>
rect 300 219 301 220 
<< m2 >>
rect 300 219 301 220 
<< m1 >>
rect 307 219 308 220 
<< m2 >>
rect 307 219 308 220 
<< m2c >>
rect 307 219 308 220 
<< m1 >>
rect 307 219 308 220 
<< m2 >>
rect 307 219 308 220 
<< m1 >>
rect 318 219 319 220 
<< m1 >>
rect 322 219 323 220 
<< m1 >>
rect 325 219 326 220 
<< m1 >>
rect 327 219 328 220 
<< m1 >>
rect 329 219 330 220 
<< m1 >>
rect 343 219 344 220 
<< m2 >>
rect 343 219 344 220 
<< m1 >>
rect 345 219 346 220 
<< m1 >>
rect 10 220 11 221 
<< m1 >>
rect 27 220 28 221 
<< m2 >>
rect 29 220 30 221 
<< m1 >>
rect 30 220 31 221 
<< m2 >>
rect 30 220 31 221 
<< m1 >>
rect 31 220 32 221 
<< m2 >>
rect 31 220 32 221 
<< m1 >>
rect 32 220 33 221 
<< m2 >>
rect 32 220 33 221 
<< m1 >>
rect 33 220 34 221 
<< m2 >>
rect 33 220 34 221 
<< m1 >>
rect 34 220 35 221 
<< m2 >>
rect 34 220 35 221 
<< m1 >>
rect 35 220 36 221 
<< m2 >>
rect 35 220 36 221 
<< m2 >>
rect 36 220 37 221 
<< m1 >>
rect 37 220 38 221 
<< m2 >>
rect 37 220 38 221 
<< m2 >>
rect 38 220 39 221 
<< m1 >>
rect 39 220 40 221 
<< m2 >>
rect 39 220 40 221 
<< m2c >>
rect 39 220 40 221 
<< m1 >>
rect 39 220 40 221 
<< m2 >>
rect 39 220 40 221 
<< m1 >>
rect 40 220 41 221 
<< m1 >>
rect 41 220 42 221 
<< m1 >>
rect 42 220 43 221 
<< m2 >>
rect 42 220 43 221 
<< m2c >>
rect 42 220 43 221 
<< m1 >>
rect 42 220 43 221 
<< m2 >>
rect 42 220 43 221 
<< m2 >>
rect 43 220 44 221 
<< m1 >>
rect 44 220 45 221 
<< m1 >>
rect 46 220 47 221 
<< m1 >>
rect 56 220 57 221 
<< m1 >>
rect 58 220 59 221 
<< m1 >>
rect 60 220 61 221 
<< m2 >>
rect 60 220 61 221 
<< m2c >>
rect 60 220 61 221 
<< m1 >>
rect 60 220 61 221 
<< m2 >>
rect 60 220 61 221 
<< m2 >>
rect 61 220 62 221 
<< m1 >>
rect 62 220 63 221 
<< m2 >>
rect 62 220 63 221 
<< m2 >>
rect 63 220 64 221 
<< m1 >>
rect 64 220 65 221 
<< m2 >>
rect 64 220 65 221 
<< m2 >>
rect 65 220 66 221 
<< m1 >>
rect 66 220 67 221 
<< m2 >>
rect 66 220 67 221 
<< m2c >>
rect 66 220 67 221 
<< m1 >>
rect 66 220 67 221 
<< m2 >>
rect 66 220 67 221 
<< m1 >>
rect 67 220 68 221 
<< m1 >>
rect 68 220 69 221 
<< m1 >>
rect 69 220 70 221 
<< m1 >>
rect 70 220 71 221 
<< m1 >>
rect 76 220 77 221 
<< m1 >>
rect 77 220 78 221 
<< m1 >>
rect 78 220 79 221 
<< m2 >>
rect 78 220 79 221 
<< m2c >>
rect 78 220 79 221 
<< m1 >>
rect 78 220 79 221 
<< m2 >>
rect 78 220 79 221 
<< m2 >>
rect 79 220 80 221 
<< m1 >>
rect 80 220 81 221 
<< m2 >>
rect 80 220 81 221 
<< m2 >>
rect 81 220 82 221 
<< m1 >>
rect 82 220 83 221 
<< m2 >>
rect 82 220 83 221 
<< m2 >>
rect 83 220 84 221 
<< m1 >>
rect 84 220 85 221 
<< m2 >>
rect 84 220 85 221 
<< m1 >>
rect 85 220 86 221 
<< m2 >>
rect 85 220 86 221 
<< m1 >>
rect 86 220 87 221 
<< m2 >>
rect 86 220 87 221 
<< m1 >>
rect 87 220 88 221 
<< m2 >>
rect 87 220 88 221 
<< m1 >>
rect 88 220 89 221 
<< m2 >>
rect 88 220 89 221 
<< m1 >>
rect 89 220 90 221 
<< m2 >>
rect 89 220 90 221 
<< m1 >>
rect 90 220 91 221 
<< m2 >>
rect 90 220 91 221 
<< m1 >>
rect 91 220 92 221 
<< m2 >>
rect 91 220 92 221 
<< m1 >>
rect 92 220 93 221 
<< m2 >>
rect 92 220 93 221 
<< m1 >>
rect 93 220 94 221 
<< m2 >>
rect 93 220 94 221 
<< m1 >>
rect 94 220 95 221 
<< m2 >>
rect 94 220 95 221 
<< m1 >>
rect 95 220 96 221 
<< m2 >>
rect 95 220 96 221 
<< m1 >>
rect 96 220 97 221 
<< m2 >>
rect 96 220 97 221 
<< m1 >>
rect 97 220 98 221 
<< m2 >>
rect 97 220 98 221 
<< m1 >>
rect 98 220 99 221 
<< m2 >>
rect 98 220 99 221 
<< m1 >>
rect 99 220 100 221 
<< m2 >>
rect 99 220 100 221 
<< m1 >>
rect 100 220 101 221 
<< m2 >>
rect 100 220 101 221 
<< m1 >>
rect 101 220 102 221 
<< m1 >>
rect 102 220 103 221 
<< m1 >>
rect 103 220 104 221 
<< m1 >>
rect 104 220 105 221 
<< m1 >>
rect 105 220 106 221 
<< m1 >>
rect 106 220 107 221 
<< m1 >>
rect 118 220 119 221 
<< m1 >>
rect 130 220 131 221 
<< m1 >>
rect 132 220 133 221 
<< m2 >>
rect 132 220 133 221 
<< m2 >>
rect 133 220 134 221 
<< m1 >>
rect 134 220 135 221 
<< m2 >>
rect 134 220 135 221 
<< m2c >>
rect 134 220 135 221 
<< m1 >>
rect 134 220 135 221 
<< m2 >>
rect 134 220 135 221 
<< m2 >>
rect 135 220 136 221 
<< m1 >>
rect 136 220 137 221 
<< m2 >>
rect 136 220 137 221 
<< m2 >>
rect 137 220 138 221 
<< m1 >>
rect 138 220 139 221 
<< m2 >>
rect 138 220 139 221 
<< m2c >>
rect 138 220 139 221 
<< m1 >>
rect 138 220 139 221 
<< m2 >>
rect 138 220 139 221 
<< m1 >>
rect 139 220 140 221 
<< m1 >>
rect 140 220 141 221 
<< m2 >>
rect 140 220 141 221 
<< m1 >>
rect 141 220 142 221 
<< m1 >>
rect 142 220 143 221 
<< m1 >>
rect 143 220 144 221 
<< m2 >>
rect 143 220 144 221 
<< m2c >>
rect 143 220 144 221 
<< m1 >>
rect 143 220 144 221 
<< m2 >>
rect 143 220 144 221 
<< m2 >>
rect 144 220 145 221 
<< m1 >>
rect 145 220 146 221 
<< m2 >>
rect 145 220 146 221 
<< m2 >>
rect 146 220 147 221 
<< m1 >>
rect 147 220 148 221 
<< m2 >>
rect 147 220 148 221 
<< m2c >>
rect 147 220 148 221 
<< m1 >>
rect 147 220 148 221 
<< m2 >>
rect 147 220 148 221 
<< m1 >>
rect 148 220 149 221 
<< m1 >>
rect 149 220 150 221 
<< m1 >>
rect 150 220 151 221 
<< m1 >>
rect 151 220 152 221 
<< m1 >>
rect 152 220 153 221 
<< m1 >>
rect 153 220 154 221 
<< m1 >>
rect 154 220 155 221 
<< m2 >>
rect 154 220 155 221 
<< m1 >>
rect 155 220 156 221 
<< m1 >>
rect 156 220 157 221 
<< m1 >>
rect 157 220 158 221 
<< m1 >>
rect 158 220 159 221 
<< m1 >>
rect 159 220 160 221 
<< m1 >>
rect 160 220 161 221 
<< m1 >>
rect 161 220 162 221 
<< m2 >>
rect 161 220 162 221 
<< m2c >>
rect 161 220 162 221 
<< m1 >>
rect 161 220 162 221 
<< m2 >>
rect 161 220 162 221 
<< m2 >>
rect 162 220 163 221 
<< m1 >>
rect 163 220 164 221 
<< m2 >>
rect 163 220 164 221 
<< m2 >>
rect 164 220 165 221 
<< m1 >>
rect 165 220 166 221 
<< m2 >>
rect 165 220 166 221 
<< m2 >>
rect 166 220 167 221 
<< m1 >>
rect 167 220 168 221 
<< m2 >>
rect 167 220 168 221 
<< m2 >>
rect 168 220 169 221 
<< m1 >>
rect 169 220 170 221 
<< m2 >>
rect 169 220 170 221 
<< m2c >>
rect 169 220 170 221 
<< m1 >>
rect 169 220 170 221 
<< m2 >>
rect 169 220 170 221 
<< m1 >>
rect 170 220 171 221 
<< m1 >>
rect 171 220 172 221 
<< m1 >>
rect 172 220 173 221 
<< m2 >>
rect 172 220 173 221 
<< m1 >>
rect 173 220 174 221 
<< m1 >>
rect 174 220 175 221 
<< m1 >>
rect 175 220 176 221 
<< m1 >>
rect 176 220 177 221 
<< m1 >>
rect 177 220 178 221 
<< m1 >>
rect 178 220 179 221 
<< m1 >>
rect 179 220 180 221 
<< m1 >>
rect 180 220 181 221 
<< m1 >>
rect 181 220 182 221 
<< m2 >>
rect 181 220 182 221 
<< m1 >>
rect 182 220 183 221 
<< m1 >>
rect 183 220 184 221 
<< m2 >>
rect 183 220 184 221 
<< m1 >>
rect 184 220 185 221 
<< m1 >>
rect 185 220 186 221 
<< m1 >>
rect 186 220 187 221 
<< m2 >>
rect 186 220 187 221 
<< m1 >>
rect 187 220 188 221 
<< m1 >>
rect 188 220 189 221 
<< m2 >>
rect 188 220 189 221 
<< m1 >>
rect 189 220 190 221 
<< m1 >>
rect 190 220 191 221 
<< m2 >>
rect 190 220 191 221 
<< m1 >>
rect 191 220 192 221 
<< m1 >>
rect 192 220 193 221 
<< m1 >>
rect 193 220 194 221 
<< m1 >>
rect 194 220 195 221 
<< m1 >>
rect 195 220 196 221 
<< m1 >>
rect 196 220 197 221 
<< m1 >>
rect 199 220 200 221 
<< m1 >>
rect 201 220 202 221 
<< m1 >>
rect 202 220 203 221 
<< m1 >>
rect 203 220 204 221 
<< m1 >>
rect 204 220 205 221 
<< m1 >>
rect 205 220 206 221 
<< m1 >>
rect 206 220 207 221 
<< m1 >>
rect 207 220 208 221 
<< m1 >>
rect 208 220 209 221 
<< m1 >>
rect 209 220 210 221 
<< m1 >>
rect 210 220 211 221 
<< m1 >>
rect 211 220 212 221 
<< m1 >>
rect 212 220 213 221 
<< m2 >>
rect 212 220 213 221 
<< m2c >>
rect 212 220 213 221 
<< m1 >>
rect 212 220 213 221 
<< m2 >>
rect 212 220 213 221 
<< m1 >>
rect 216 220 217 221 
<< m1 >>
rect 218 220 219 221 
<< m1 >>
rect 226 220 227 221 
<< m1 >>
rect 228 220 229 221 
<< m1 >>
rect 235 220 236 221 
<< m1 >>
rect 237 220 238 221 
<< m1 >>
rect 241 220 242 221 
<< m1 >>
rect 243 220 244 221 
<< m1 >>
rect 253 220 254 221 
<< m1 >>
rect 260 220 261 221 
<< m1 >>
rect 262 220 263 221 
<< m2 >>
rect 264 220 265 221 
<< m1 >>
rect 272 220 273 221 
<< m2 >>
rect 282 220 283 221 
<< m2 >>
rect 300 220 301 221 
<< m2 >>
rect 307 220 308 221 
<< m1 >>
rect 318 220 319 221 
<< m1 >>
rect 319 220 320 221 
<< m1 >>
rect 320 220 321 221 
<< m2 >>
rect 320 220 321 221 
<< m2c >>
rect 320 220 321 221 
<< m1 >>
rect 320 220 321 221 
<< m2 >>
rect 320 220 321 221 
<< m2 >>
rect 321 220 322 221 
<< m1 >>
rect 322 220 323 221 
<< m1 >>
rect 325 220 326 221 
<< m1 >>
rect 327 220 328 221 
<< m1 >>
rect 329 220 330 221 
<< m1 >>
rect 343 220 344 221 
<< m2 >>
rect 343 220 344 221 
<< m1 >>
rect 345 220 346 221 
<< m1 >>
rect 10 221 11 222 
<< m1 >>
rect 27 221 28 222 
<< m1 >>
rect 30 221 31 222 
<< m1 >>
rect 37 221 38 222 
<< m2 >>
rect 43 221 44 222 
<< m1 >>
rect 44 221 45 222 
<< m1 >>
rect 46 221 47 222 
<< m1 >>
rect 56 221 57 222 
<< m1 >>
rect 58 221 59 222 
<< m1 >>
rect 60 221 61 222 
<< m1 >>
rect 62 221 63 222 
<< m1 >>
rect 64 221 65 222 
<< m1 >>
rect 76 221 77 222 
<< m1 >>
rect 80 221 81 222 
<< m1 >>
rect 82 221 83 222 
<< m1 >>
rect 118 221 119 222 
<< m1 >>
rect 130 221 131 222 
<< m1 >>
rect 132 221 133 222 
<< m2 >>
rect 132 221 133 222 
<< m1 >>
rect 136 221 137 222 
<< m2 >>
rect 140 221 141 222 
<< m1 >>
rect 145 221 146 222 
<< m2 >>
rect 154 221 155 222 
<< m1 >>
rect 163 221 164 222 
<< m1 >>
rect 165 221 166 222 
<< m1 >>
rect 167 221 168 222 
<< m2 >>
rect 172 221 173 222 
<< m2 >>
rect 181 221 182 222 
<< m2 >>
rect 183 221 184 222 
<< m2 >>
rect 186 221 187 222 
<< m2 >>
rect 188 221 189 222 
<< m2 >>
rect 190 221 191 222 
<< m1 >>
rect 199 221 200 222 
<< m1 >>
rect 216 221 217 222 
<< m2 >>
rect 216 221 217 222 
<< m2c >>
rect 216 221 217 222 
<< m1 >>
rect 216 221 217 222 
<< m2 >>
rect 216 221 217 222 
<< m1 >>
rect 218 221 219 222 
<< m2 >>
rect 218 221 219 222 
<< m2c >>
rect 218 221 219 222 
<< m1 >>
rect 218 221 219 222 
<< m2 >>
rect 218 221 219 222 
<< m1 >>
rect 226 221 227 222 
<< m2 >>
rect 226 221 227 222 
<< m2c >>
rect 226 221 227 222 
<< m1 >>
rect 226 221 227 222 
<< m2 >>
rect 226 221 227 222 
<< m1 >>
rect 228 221 229 222 
<< m2 >>
rect 228 221 229 222 
<< m2c >>
rect 228 221 229 222 
<< m1 >>
rect 228 221 229 222 
<< m2 >>
rect 228 221 229 222 
<< m1 >>
rect 235 221 236 222 
<< m1 >>
rect 237 221 238 222 
<< m1 >>
rect 241 221 242 222 
<< m2 >>
rect 241 221 242 222 
<< m2c >>
rect 241 221 242 222 
<< m1 >>
rect 241 221 242 222 
<< m2 >>
rect 241 221 242 222 
<< m1 >>
rect 243 221 244 222 
<< m2 >>
rect 243 221 244 222 
<< m2c >>
rect 243 221 244 222 
<< m1 >>
rect 243 221 244 222 
<< m2 >>
rect 243 221 244 222 
<< m1 >>
rect 253 221 254 222 
<< m2 >>
rect 253 221 254 222 
<< m2c >>
rect 253 221 254 222 
<< m1 >>
rect 253 221 254 222 
<< m2 >>
rect 253 221 254 222 
<< m1 >>
rect 260 221 261 222 
<< m2 >>
rect 260 221 261 222 
<< m2c >>
rect 260 221 261 222 
<< m1 >>
rect 260 221 261 222 
<< m2 >>
rect 260 221 261 222 
<< m2 >>
rect 261 221 262 222 
<< m1 >>
rect 262 221 263 222 
<< m2 >>
rect 262 221 263 222 
<< m1 >>
rect 263 221 264 222 
<< m1 >>
rect 264 221 265 222 
<< m2 >>
rect 264 221 265 222 
<< m1 >>
rect 265 221 266 222 
<< m2 >>
rect 265 221 266 222 
<< m1 >>
rect 266 221 267 222 
<< m2 >>
rect 266 221 267 222 
<< m1 >>
rect 267 221 268 222 
<< m2 >>
rect 267 221 268 222 
<< m1 >>
rect 268 221 269 222 
<< m2 >>
rect 268 221 269 222 
<< m1 >>
rect 269 221 270 222 
<< m2 >>
rect 269 221 270 222 
<< m1 >>
rect 270 221 271 222 
<< m2 >>
rect 270 221 271 222 
<< m2 >>
rect 271 221 272 222 
<< m1 >>
rect 272 221 273 222 
<< m2 >>
rect 272 221 273 222 
<< m2 >>
rect 273 221 274 222 
<< m1 >>
rect 274 221 275 222 
<< m2 >>
rect 274 221 275 222 
<< m2c >>
rect 274 221 275 222 
<< m1 >>
rect 274 221 275 222 
<< m2 >>
rect 274 221 275 222 
<< m1 >>
rect 275 221 276 222 
<< m1 >>
rect 276 221 277 222 
<< m1 >>
rect 277 221 278 222 
<< m1 >>
rect 278 221 279 222 
<< m1 >>
rect 279 221 280 222 
<< m1 >>
rect 280 221 281 222 
<< m1 >>
rect 281 221 282 222 
<< m1 >>
rect 282 221 283 222 
<< m2 >>
rect 282 221 283 222 
<< m1 >>
rect 283 221 284 222 
<< m1 >>
rect 284 221 285 222 
<< m1 >>
rect 285 221 286 222 
<< m1 >>
rect 286 221 287 222 
<< m1 >>
rect 287 221 288 222 
<< m1 >>
rect 288 221 289 222 
<< m1 >>
rect 289 221 290 222 
<< m1 >>
rect 290 221 291 222 
<< m1 >>
rect 291 221 292 222 
<< m1 >>
rect 292 221 293 222 
<< m1 >>
rect 293 221 294 222 
<< m1 >>
rect 294 221 295 222 
<< m1 >>
rect 295 221 296 222 
<< m1 >>
rect 296 221 297 222 
<< m1 >>
rect 297 221 298 222 
<< m1 >>
rect 298 221 299 222 
<< m1 >>
rect 299 221 300 222 
<< m1 >>
rect 300 221 301 222 
<< m2 >>
rect 300 221 301 222 
<< m1 >>
rect 301 221 302 222 
<< m1 >>
rect 302 221 303 222 
<< m1 >>
rect 303 221 304 222 
<< m1 >>
rect 304 221 305 222 
<< m1 >>
rect 305 221 306 222 
<< m1 >>
rect 306 221 307 222 
<< m1 >>
rect 307 221 308 222 
<< m2 >>
rect 307 221 308 222 
<< m1 >>
rect 308 221 309 222 
<< m1 >>
rect 309 221 310 222 
<< m1 >>
rect 310 221 311 222 
<< m1 >>
rect 311 221 312 222 
<< m1 >>
rect 312 221 313 222 
<< m1 >>
rect 313 221 314 222 
<< m1 >>
rect 314 221 315 222 
<< m1 >>
rect 315 221 316 222 
<< m1 >>
rect 316 221 317 222 
<< m2 >>
rect 316 221 317 222 
<< m2c >>
rect 316 221 317 222 
<< m1 >>
rect 316 221 317 222 
<< m2 >>
rect 316 221 317 222 
<< m2 >>
rect 321 221 322 222 
<< m1 >>
rect 322 221 323 222 
<< m1 >>
rect 325 221 326 222 
<< m1 >>
rect 327 221 328 222 
<< m1 >>
rect 329 221 330 222 
<< m1 >>
rect 343 221 344 222 
<< m2 >>
rect 343 221 344 222 
<< m1 >>
rect 345 221 346 222 
<< m1 >>
rect 10 222 11 223 
<< m1 >>
rect 27 222 28 223 
<< m1 >>
rect 28 222 29 223 
<< m2 >>
rect 28 222 29 223 
<< m2c >>
rect 28 222 29 223 
<< m1 >>
rect 28 222 29 223 
<< m2 >>
rect 28 222 29 223 
<< m2 >>
rect 29 222 30 223 
<< m1 >>
rect 30 222 31 223 
<< m2 >>
rect 30 222 31 223 
<< m2 >>
rect 31 222 32 223 
<< m1 >>
rect 32 222 33 223 
<< m2 >>
rect 32 222 33 223 
<< m2c >>
rect 32 222 33 223 
<< m1 >>
rect 32 222 33 223 
<< m2 >>
rect 32 222 33 223 
<< m1 >>
rect 33 222 34 223 
<< m1 >>
rect 34 222 35 223 
<< m1 >>
rect 35 222 36 223 
<< m2 >>
rect 35 222 36 223 
<< m2c >>
rect 35 222 36 223 
<< m1 >>
rect 35 222 36 223 
<< m2 >>
rect 35 222 36 223 
<< m2 >>
rect 36 222 37 223 
<< m1 >>
rect 37 222 38 223 
<< m2 >>
rect 37 222 38 223 
<< m2 >>
rect 38 222 39 223 
<< m1 >>
rect 39 222 40 223 
<< m2 >>
rect 39 222 40 223 
<< m2c >>
rect 39 222 40 223 
<< m1 >>
rect 39 222 40 223 
<< m2 >>
rect 39 222 40 223 
<< m2 >>
rect 43 222 44 223 
<< m1 >>
rect 44 222 45 223 
<< m1 >>
rect 46 222 47 223 
<< m2 >>
rect 46 222 47 223 
<< m2 >>
rect 47 222 48 223 
<< m1 >>
rect 48 222 49 223 
<< m2 >>
rect 48 222 49 223 
<< m2c >>
rect 48 222 49 223 
<< m1 >>
rect 48 222 49 223 
<< m2 >>
rect 48 222 49 223 
<< m1 >>
rect 49 222 50 223 
<< m1 >>
rect 50 222 51 223 
<< m1 >>
rect 51 222 52 223 
<< m1 >>
rect 52 222 53 223 
<< m1 >>
rect 53 222 54 223 
<< m1 >>
rect 54 222 55 223 
<< m2 >>
rect 54 222 55 223 
<< m2c >>
rect 54 222 55 223 
<< m1 >>
rect 54 222 55 223 
<< m2 >>
rect 54 222 55 223 
<< m2 >>
rect 55 222 56 223 
<< m1 >>
rect 56 222 57 223 
<< m2 >>
rect 56 222 57 223 
<< m2 >>
rect 57 222 58 223 
<< m1 >>
rect 58 222 59 223 
<< m2 >>
rect 58 222 59 223 
<< m2 >>
rect 59 222 60 223 
<< m1 >>
rect 60 222 61 223 
<< m2 >>
rect 60 222 61 223 
<< m2 >>
rect 61 222 62 223 
<< m1 >>
rect 62 222 63 223 
<< m2 >>
rect 62 222 63 223 
<< m2 >>
rect 63 222 64 223 
<< m1 >>
rect 64 222 65 223 
<< m2 >>
rect 64 222 65 223 
<< m2 >>
rect 65 222 66 223 
<< m1 >>
rect 66 222 67 223 
<< m2 >>
rect 66 222 67 223 
<< m2c >>
rect 66 222 67 223 
<< m1 >>
rect 66 222 67 223 
<< m2 >>
rect 66 222 67 223 
<< m1 >>
rect 67 222 68 223 
<< m1 >>
rect 68 222 69 223 
<< m1 >>
rect 69 222 70 223 
<< m1 >>
rect 70 222 71 223 
<< m1 >>
rect 71 222 72 223 
<< m1 >>
rect 72 222 73 223 
<< m1 >>
rect 73 222 74 223 
<< m1 >>
rect 74 222 75 223 
<< m1 >>
rect 75 222 76 223 
<< m1 >>
rect 76 222 77 223 
<< m1 >>
rect 80 222 81 223 
<< m1 >>
rect 82 222 83 223 
<< m1 >>
rect 118 222 119 223 
<< m1 >>
rect 130 222 131 223 
<< m1 >>
rect 132 222 133 223 
<< m2 >>
rect 132 222 133 223 
<< m1 >>
rect 136 222 137 223 
<< m1 >>
rect 140 222 141 223 
<< m2 >>
rect 140 222 141 223 
<< m2c >>
rect 140 222 141 223 
<< m1 >>
rect 140 222 141 223 
<< m2 >>
rect 140 222 141 223 
<< m1 >>
rect 145 222 146 223 
<< m1 >>
rect 154 222 155 223 
<< m2 >>
rect 154 222 155 223 
<< m2c >>
rect 154 222 155 223 
<< m1 >>
rect 154 222 155 223 
<< m2 >>
rect 154 222 155 223 
<< m1 >>
rect 163 222 164 223 
<< m1 >>
rect 165 222 166 223 
<< m1 >>
rect 167 222 168 223 
<< m2 >>
rect 168 222 169 223 
<< m1 >>
rect 169 222 170 223 
<< m2 >>
rect 169 222 170 223 
<< m2c >>
rect 169 222 170 223 
<< m1 >>
rect 169 222 170 223 
<< m2 >>
rect 169 222 170 223 
<< m1 >>
rect 170 222 171 223 
<< m1 >>
rect 171 222 172 223 
<< m1 >>
rect 172 222 173 223 
<< m2 >>
rect 172 222 173 223 
<< m2c >>
rect 172 222 173 223 
<< m1 >>
rect 172 222 173 223 
<< m2 >>
rect 172 222 173 223 
<< m1 >>
rect 181 222 182 223 
<< m2 >>
rect 181 222 182 223 
<< m2c >>
rect 181 222 182 223 
<< m1 >>
rect 181 222 182 223 
<< m2 >>
rect 181 222 182 223 
<< m1 >>
rect 183 222 184 223 
<< m2 >>
rect 183 222 184 223 
<< m2c >>
rect 183 222 184 223 
<< m1 >>
rect 183 222 184 223 
<< m2 >>
rect 183 222 184 223 
<< m1 >>
rect 186 222 187 223 
<< m2 >>
rect 186 222 187 223 
<< m2c >>
rect 186 222 187 223 
<< m1 >>
rect 186 222 187 223 
<< m2 >>
rect 186 222 187 223 
<< m1 >>
rect 188 222 189 223 
<< m2 >>
rect 188 222 189 223 
<< m2c >>
rect 188 222 189 223 
<< m1 >>
rect 188 222 189 223 
<< m2 >>
rect 188 222 189 223 
<< m1 >>
rect 190 222 191 223 
<< m2 >>
rect 190 222 191 223 
<< m2c >>
rect 190 222 191 223 
<< m1 >>
rect 190 222 191 223 
<< m2 >>
rect 190 222 191 223 
<< m1 >>
rect 199 222 200 223 
<< m2 >>
rect 216 222 217 223 
<< m2 >>
rect 218 222 219 223 
<< m2 >>
rect 219 222 220 223 
<< m2 >>
rect 220 222 221 223 
<< m2 >>
rect 221 222 222 223 
<< m2 >>
rect 226 222 227 223 
<< m2 >>
rect 228 222 229 223 
<< m2 >>
rect 229 222 230 223 
<< m2 >>
rect 230 222 231 223 
<< m1 >>
rect 235 222 236 223 
<< m1 >>
rect 237 222 238 223 
<< m2 >>
rect 241 222 242 223 
<< m2 >>
rect 243 222 244 223 
<< m2 >>
rect 253 222 254 223 
<< m2 >>
rect 262 222 263 223 
<< m1 >>
rect 270 222 271 223 
<< m1 >>
rect 272 222 273 223 
<< m2 >>
rect 282 222 283 223 
<< m2 >>
rect 300 222 301 223 
<< m2 >>
rect 307 222 308 223 
<< m2 >>
rect 316 222 317 223 
<< m2 >>
rect 321 222 322 223 
<< m1 >>
rect 322 222 323 223 
<< m1 >>
rect 325 222 326 223 
<< m1 >>
rect 327 222 328 223 
<< m1 >>
rect 329 222 330 223 
<< m1 >>
rect 343 222 344 223 
<< m2 >>
rect 343 222 344 223 
<< m1 >>
rect 345 222 346 223 
<< m1 >>
rect 10 223 11 224 
<< m1 >>
rect 30 223 31 224 
<< m1 >>
rect 37 223 38 224 
<< m1 >>
rect 39 223 40 224 
<< m2 >>
rect 43 223 44 224 
<< m1 >>
rect 44 223 45 224 
<< m1 >>
rect 46 223 47 224 
<< m2 >>
rect 46 223 47 224 
<< m1 >>
rect 56 223 57 224 
<< m1 >>
rect 58 223 59 224 
<< m1 >>
rect 60 223 61 224 
<< m1 >>
rect 62 223 63 224 
<< m1 >>
rect 64 223 65 224 
<< m1 >>
rect 78 223 79 224 
<< m2 >>
rect 78 223 79 224 
<< m2c >>
rect 78 223 79 224 
<< m1 >>
rect 78 223 79 224 
<< m2 >>
rect 78 223 79 224 
<< m2 >>
rect 79 223 80 224 
<< m1 >>
rect 80 223 81 224 
<< m2 >>
rect 80 223 81 224 
<< m2 >>
rect 81 223 82 224 
<< m1 >>
rect 82 223 83 224 
<< m2 >>
rect 82 223 83 224 
<< m2 >>
rect 83 223 84 224 
<< m1 >>
rect 84 223 85 224 
<< m2 >>
rect 84 223 85 224 
<< m2c >>
rect 84 223 85 224 
<< m1 >>
rect 84 223 85 224 
<< m2 >>
rect 84 223 85 224 
<< m1 >>
rect 85 223 86 224 
<< m1 >>
rect 86 223 87 224 
<< m1 >>
rect 87 223 88 224 
<< m1 >>
rect 88 223 89 224 
<< m1 >>
rect 118 223 119 224 
<< m1 >>
rect 130 223 131 224 
<< m1 >>
rect 132 223 133 224 
<< m2 >>
rect 132 223 133 224 
<< m1 >>
rect 136 223 137 224 
<< m1 >>
rect 140 223 141 224 
<< m1 >>
rect 145 223 146 224 
<< m1 >>
rect 154 223 155 224 
<< m1 >>
rect 163 223 164 224 
<< m1 >>
rect 165 223 166 224 
<< m1 >>
rect 167 223 168 224 
<< m2 >>
rect 168 223 169 224 
<< m1 >>
rect 181 223 182 224 
<< m1 >>
rect 183 223 184 224 
<< m1 >>
rect 186 223 187 224 
<< m1 >>
rect 188 223 189 224 
<< m1 >>
rect 190 223 191 224 
<< m1 >>
rect 199 223 200 224 
<< m2 >>
rect 216 223 217 224 
<< m1 >>
rect 217 223 218 224 
<< m1 >>
rect 218 223 219 224 
<< m1 >>
rect 219 223 220 224 
<< m1 >>
rect 220 223 221 224 
<< m1 >>
rect 221 223 222 224 
<< m2 >>
rect 221 223 222 224 
<< m1 >>
rect 222 223 223 224 
<< m1 >>
rect 223 223 224 224 
<< m1 >>
rect 224 223 225 224 
<< m1 >>
rect 225 223 226 224 
<< m1 >>
rect 226 223 227 224 
<< m2 >>
rect 226 223 227 224 
<< m1 >>
rect 227 223 228 224 
<< m1 >>
rect 228 223 229 224 
<< m1 >>
rect 229 223 230 224 
<< m1 >>
rect 230 223 231 224 
<< m2 >>
rect 230 223 231 224 
<< m1 >>
rect 231 223 232 224 
<< m1 >>
rect 232 223 233 224 
<< m1 >>
rect 233 223 234 224 
<< m2 >>
rect 233 223 234 224 
<< m2c >>
rect 233 223 234 224 
<< m1 >>
rect 233 223 234 224 
<< m2 >>
rect 233 223 234 224 
<< m2 >>
rect 234 223 235 224 
<< m1 >>
rect 235 223 236 224 
<< m2 >>
rect 235 223 236 224 
<< m2 >>
rect 236 223 237 224 
<< m1 >>
rect 237 223 238 224 
<< m2 >>
rect 237 223 238 224 
<< m2 >>
rect 238 223 239 224 
<< m1 >>
rect 239 223 240 224 
<< m2 >>
rect 239 223 240 224 
<< m2c >>
rect 239 223 240 224 
<< m1 >>
rect 239 223 240 224 
<< m2 >>
rect 239 223 240 224 
<< m1 >>
rect 240 223 241 224 
<< m1 >>
rect 241 223 242 224 
<< m2 >>
rect 241 223 242 224 
<< m1 >>
rect 242 223 243 224 
<< m1 >>
rect 243 223 244 224 
<< m2 >>
rect 243 223 244 224 
<< m1 >>
rect 244 223 245 224 
<< m1 >>
rect 245 223 246 224 
<< m1 >>
rect 246 223 247 224 
<< m1 >>
rect 247 223 248 224 
<< m1 >>
rect 248 223 249 224 
<< m1 >>
rect 249 223 250 224 
<< m1 >>
rect 250 223 251 224 
<< m1 >>
rect 251 223 252 224 
<< m1 >>
rect 252 223 253 224 
<< m1 >>
rect 253 223 254 224 
<< m2 >>
rect 253 223 254 224 
<< m1 >>
rect 254 223 255 224 
<< m1 >>
rect 255 223 256 224 
<< m1 >>
rect 256 223 257 224 
<< m1 >>
rect 257 223 258 224 
<< m1 >>
rect 258 223 259 224 
<< m1 >>
rect 259 223 260 224 
<< m1 >>
rect 260 223 261 224 
<< m1 >>
rect 261 223 262 224 
<< m1 >>
rect 262 223 263 224 
<< m2 >>
rect 262 223 263 224 
<< m1 >>
rect 263 223 264 224 
<< m1 >>
rect 264 223 265 224 
<< m2 >>
rect 264 223 265 224 
<< m1 >>
rect 265 223 266 224 
<< m2 >>
rect 265 223 266 224 
<< m1 >>
rect 266 223 267 224 
<< m2 >>
rect 266 223 267 224 
<< m1 >>
rect 267 223 268 224 
<< m2 >>
rect 267 223 268 224 
<< m1 >>
rect 268 223 269 224 
<< m2 >>
rect 268 223 269 224 
<< m2 >>
rect 269 223 270 224 
<< m1 >>
rect 270 223 271 224 
<< m2 >>
rect 270 223 271 224 
<< m2 >>
rect 271 223 272 224 
<< m1 >>
rect 272 223 273 224 
<< m2 >>
rect 272 223 273 224 
<< m2 >>
rect 273 223 274 224 
<< m1 >>
rect 282 223 283 224 
<< m2 >>
rect 282 223 283 224 
<< m1 >>
rect 283 223 284 224 
<< m2 >>
rect 283 223 284 224 
<< m1 >>
rect 284 223 285 224 
<< m2 >>
rect 284 223 285 224 
<< m1 >>
rect 285 223 286 224 
<< m2 >>
rect 285 223 286 224 
<< m1 >>
rect 286 223 287 224 
<< m2 >>
rect 286 223 287 224 
<< m1 >>
rect 287 223 288 224 
<< m2 >>
rect 287 223 288 224 
<< m1 >>
rect 288 223 289 224 
<< m2 >>
rect 288 223 289 224 
<< m1 >>
rect 289 223 290 224 
<< m2 >>
rect 289 223 290 224 
<< m1 >>
rect 290 223 291 224 
<< m2 >>
rect 290 223 291 224 
<< m1 >>
rect 291 223 292 224 
<< m2 >>
rect 291 223 292 224 
<< m1 >>
rect 292 223 293 224 
<< m2 >>
rect 292 223 293 224 
<< m1 >>
rect 293 223 294 224 
<< m2 >>
rect 293 223 294 224 
<< m1 >>
rect 294 223 295 224 
<< m2 >>
rect 294 223 295 224 
<< m1 >>
rect 295 223 296 224 
<< m2 >>
rect 295 223 296 224 
<< m1 >>
rect 296 223 297 224 
<< m2 >>
rect 296 223 297 224 
<< m1 >>
rect 297 223 298 224 
<< m2 >>
rect 297 223 298 224 
<< m1 >>
rect 298 223 299 224 
<< m2 >>
rect 298 223 299 224 
<< m1 >>
rect 299 223 300 224 
<< m1 >>
rect 300 223 301 224 
<< m2 >>
rect 300 223 301 224 
<< m1 >>
rect 301 223 302 224 
<< m2 >>
rect 301 223 302 224 
<< m1 >>
rect 302 223 303 224 
<< m2 >>
rect 302 223 303 224 
<< m1 >>
rect 303 223 304 224 
<< m2 >>
rect 303 223 304 224 
<< m1 >>
rect 304 223 305 224 
<< m2 >>
rect 304 223 305 224 
<< m1 >>
rect 305 223 306 224 
<< m1 >>
rect 306 223 307 224 
<< m1 >>
rect 307 223 308 224 
<< m2 >>
rect 307 223 308 224 
<< m1 >>
rect 308 223 309 224 
<< m1 >>
rect 309 223 310 224 
<< m1 >>
rect 310 223 311 224 
<< m1 >>
rect 311 223 312 224 
<< m1 >>
rect 312 223 313 224 
<< m1 >>
rect 313 223 314 224 
<< m1 >>
rect 314 223 315 224 
<< m1 >>
rect 315 223 316 224 
<< m1 >>
rect 316 223 317 224 
<< m2 >>
rect 316 223 317 224 
<< m1 >>
rect 317 223 318 224 
<< m1 >>
rect 318 223 319 224 
<< m1 >>
rect 319 223 320 224 
<< m1 >>
rect 320 223 321 224 
<< m1 >>
rect 321 223 322 224 
<< m2 >>
rect 321 223 322 224 
<< m1 >>
rect 322 223 323 224 
<< m1 >>
rect 325 223 326 224 
<< m1 >>
rect 327 223 328 224 
<< m1 >>
rect 329 223 330 224 
<< m1 >>
rect 331 223 332 224 
<< m1 >>
rect 332 223 333 224 
<< m1 >>
rect 333 223 334 224 
<< m1 >>
rect 334 223 335 224 
<< m1 >>
rect 335 223 336 224 
<< m1 >>
rect 336 223 337 224 
<< m1 >>
rect 337 223 338 224 
<< m1 >>
rect 338 223 339 224 
<< m1 >>
rect 339 223 340 224 
<< m1 >>
rect 340 223 341 224 
<< m1 >>
rect 341 223 342 224 
<< m1 >>
rect 342 223 343 224 
<< m1 >>
rect 343 223 344 224 
<< m2 >>
rect 343 223 344 224 
<< m1 >>
rect 345 223 346 224 
<< m1 >>
rect 10 224 11 225 
<< m2 >>
rect 28 224 29 225 
<< m2 >>
rect 29 224 30 225 
<< m1 >>
rect 30 224 31 225 
<< m2 >>
rect 30 224 31 225 
<< m2c >>
rect 30 224 31 225 
<< m1 >>
rect 30 224 31 225 
<< m2 >>
rect 30 224 31 225 
<< m1 >>
rect 37 224 38 225 
<< m1 >>
rect 39 224 40 225 
<< m2 >>
rect 43 224 44 225 
<< m1 >>
rect 44 224 45 225 
<< m1 >>
rect 46 224 47 225 
<< m2 >>
rect 46 224 47 225 
<< m1 >>
rect 56 224 57 225 
<< m1 >>
rect 58 224 59 225 
<< m1 >>
rect 60 224 61 225 
<< m1 >>
rect 62 224 63 225 
<< m1 >>
rect 64 224 65 225 
<< m1 >>
rect 78 224 79 225 
<< m1 >>
rect 80 224 81 225 
<< m1 >>
rect 82 224 83 225 
<< m1 >>
rect 88 224 89 225 
<< m1 >>
rect 118 224 119 225 
<< m1 >>
rect 130 224 131 225 
<< m1 >>
rect 132 224 133 225 
<< m2 >>
rect 132 224 133 225 
<< m1 >>
rect 136 224 137 225 
<< m1 >>
rect 140 224 141 225 
<< m1 >>
rect 145 224 146 225 
<< m1 >>
rect 154 224 155 225 
<< m1 >>
rect 163 224 164 225 
<< m1 >>
rect 165 224 166 225 
<< m1 >>
rect 167 224 168 225 
<< m2 >>
rect 168 224 169 225 
<< m1 >>
rect 181 224 182 225 
<< m1 >>
rect 183 224 184 225 
<< m1 >>
rect 186 224 187 225 
<< m1 >>
rect 188 224 189 225 
<< m1 >>
rect 190 224 191 225 
<< m1 >>
rect 199 224 200 225 
<< m2 >>
rect 216 224 217 225 
<< m1 >>
rect 217 224 218 225 
<< m2 >>
rect 221 224 222 225 
<< m2 >>
rect 226 224 227 225 
<< m2 >>
rect 230 224 231 225 
<< m1 >>
rect 235 224 236 225 
<< m1 >>
rect 237 224 238 225 
<< m2 >>
rect 241 224 242 225 
<< m2 >>
rect 243 224 244 225 
<< m2 >>
rect 253 224 254 225 
<< m2 >>
rect 262 224 263 225 
<< m2 >>
rect 264 224 265 225 
<< m1 >>
rect 268 224 269 225 
<< m1 >>
rect 270 224 271 225 
<< m1 >>
rect 272 224 273 225 
<< m2 >>
rect 273 224 274 225 
<< m1 >>
rect 274 224 275 225 
<< m2 >>
rect 274 224 275 225 
<< m2c >>
rect 274 224 275 225 
<< m1 >>
rect 274 224 275 225 
<< m2 >>
rect 274 224 275 225 
<< m1 >>
rect 275 224 276 225 
<< m1 >>
rect 276 224 277 225 
<< m1 >>
rect 277 224 278 225 
<< m1 >>
rect 278 224 279 225 
<< m1 >>
rect 279 224 280 225 
<< m1 >>
rect 280 224 281 225 
<< m1 >>
rect 282 224 283 225 
<< m2 >>
rect 298 224 299 225 
<< m2 >>
rect 304 224 305 225 
<< m2 >>
rect 307 224 308 225 
<< m2 >>
rect 316 224 317 225 
<< m2 >>
rect 321 224 322 225 
<< m1 >>
rect 325 224 326 225 
<< m1 >>
rect 327 224 328 225 
<< m1 >>
rect 329 224 330 225 
<< m1 >>
rect 331 224 332 225 
<< m2 >>
rect 343 224 344 225 
<< m1 >>
rect 345 224 346 225 
<< m1 >>
rect 10 225 11 226 
<< m1 >>
rect 13 225 14 226 
<< m1 >>
rect 14 225 15 226 
<< m1 >>
rect 15 225 16 226 
<< m1 >>
rect 16 225 17 226 
<< m1 >>
rect 17 225 18 226 
<< m1 >>
rect 18 225 19 226 
<< m1 >>
rect 19 225 20 226 
<< m1 >>
rect 20 225 21 226 
<< m1 >>
rect 21 225 22 226 
<< m1 >>
rect 22 225 23 226 
<< m1 >>
rect 23 225 24 226 
<< m1 >>
rect 24 225 25 226 
<< m1 >>
rect 25 225 26 226 
<< m1 >>
rect 26 225 27 226 
<< m1 >>
rect 27 225 28 226 
<< m1 >>
rect 28 225 29 226 
<< m2 >>
rect 28 225 29 226 
<< m1 >>
rect 37 225 38 226 
<< m1 >>
rect 39 225 40 226 
<< m2 >>
rect 43 225 44 226 
<< m1 >>
rect 44 225 45 226 
<< m1 >>
rect 46 225 47 226 
<< m2 >>
rect 46 225 47 226 
<< m1 >>
rect 56 225 57 226 
<< m1 >>
rect 58 225 59 226 
<< m1 >>
rect 60 225 61 226 
<< m1 >>
rect 62 225 63 226 
<< m1 >>
rect 64 225 65 226 
<< m1 >>
rect 78 225 79 226 
<< m1 >>
rect 80 225 81 226 
<< m1 >>
rect 82 225 83 226 
<< m1 >>
rect 88 225 89 226 
<< m1 >>
rect 118 225 119 226 
<< m1 >>
rect 130 225 131 226 
<< m1 >>
rect 132 225 133 226 
<< m2 >>
rect 132 225 133 226 
<< m1 >>
rect 136 225 137 226 
<< m1 >>
rect 140 225 141 226 
<< m1 >>
rect 145 225 146 226 
<< m1 >>
rect 154 225 155 226 
<< m1 >>
rect 163 225 164 226 
<< m1 >>
rect 165 225 166 226 
<< m1 >>
rect 167 225 168 226 
<< m2 >>
rect 168 225 169 226 
<< m1 >>
rect 181 225 182 226 
<< m1 >>
rect 183 225 184 226 
<< m1 >>
rect 186 225 187 226 
<< m1 >>
rect 188 225 189 226 
<< m1 >>
rect 190 225 191 226 
<< m1 >>
rect 193 225 194 226 
<< m1 >>
rect 194 225 195 226 
<< m1 >>
rect 195 225 196 226 
<< m1 >>
rect 196 225 197 226 
<< m1 >>
rect 197 225 198 226 
<< m1 >>
rect 198 225 199 226 
<< m1 >>
rect 199 225 200 226 
<< m2 >>
rect 216 225 217 226 
<< m1 >>
rect 217 225 218 226 
<< m2 >>
rect 217 225 218 226 
<< m2 >>
rect 218 225 219 226 
<< m1 >>
rect 219 225 220 226 
<< m2 >>
rect 219 225 220 226 
<< m2c >>
rect 219 225 220 226 
<< m1 >>
rect 219 225 220 226 
<< m2 >>
rect 219 225 220 226 
<< m1 >>
rect 221 225 222 226 
<< m2 >>
rect 221 225 222 226 
<< m2c >>
rect 221 225 222 226 
<< m1 >>
rect 221 225 222 226 
<< m2 >>
rect 221 225 222 226 
<< m1 >>
rect 226 225 227 226 
<< m2 >>
rect 226 225 227 226 
<< m2c >>
rect 226 225 227 226 
<< m1 >>
rect 226 225 227 226 
<< m2 >>
rect 226 225 227 226 
<< m1 >>
rect 230 225 231 226 
<< m2 >>
rect 230 225 231 226 
<< m2c >>
rect 230 225 231 226 
<< m1 >>
rect 230 225 231 226 
<< m2 >>
rect 230 225 231 226 
<< m1 >>
rect 231 225 232 226 
<< m1 >>
rect 232 225 233 226 
<< m1 >>
rect 233 225 234 226 
<< m2 >>
rect 233 225 234 226 
<< m2c >>
rect 233 225 234 226 
<< m1 >>
rect 233 225 234 226 
<< m2 >>
rect 233 225 234 226 
<< m2 >>
rect 234 225 235 226 
<< m1 >>
rect 235 225 236 226 
<< m2 >>
rect 235 225 236 226 
<< m2 >>
rect 236 225 237 226 
<< m1 >>
rect 237 225 238 226 
<< m2 >>
rect 237 225 238 226 
<< m2 >>
rect 238 225 239 226 
<< m1 >>
rect 239 225 240 226 
<< m2 >>
rect 239 225 240 226 
<< m2c >>
rect 239 225 240 226 
<< m1 >>
rect 239 225 240 226 
<< m2 >>
rect 239 225 240 226 
<< m1 >>
rect 240 225 241 226 
<< m1 >>
rect 241 225 242 226 
<< m2 >>
rect 241 225 242 226 
<< m1 >>
rect 242 225 243 226 
<< m1 >>
rect 243 225 244 226 
<< m2 >>
rect 243 225 244 226 
<< m1 >>
rect 244 225 245 226 
<< m1 >>
rect 245 225 246 226 
<< m1 >>
rect 246 225 247 226 
<< m1 >>
rect 247 225 248 226 
<< m1 >>
rect 250 225 251 226 
<< m1 >>
rect 251 225 252 226 
<< m1 >>
rect 252 225 253 226 
<< m1 >>
rect 253 225 254 226 
<< m2 >>
rect 253 225 254 226 
<< m1 >>
rect 254 225 255 226 
<< m1 >>
rect 255 225 256 226 
<< m1 >>
rect 256 225 257 226 
<< m1 >>
rect 257 225 258 226 
<< m1 >>
rect 258 225 259 226 
<< m1 >>
rect 259 225 260 226 
<< m1 >>
rect 260 225 261 226 
<< m1 >>
rect 261 225 262 226 
<< m1 >>
rect 262 225 263 226 
<< m2 >>
rect 262 225 263 226 
<< m1 >>
rect 263 225 264 226 
<< m1 >>
rect 264 225 265 226 
<< m2 >>
rect 264 225 265 226 
<< m2c >>
rect 264 225 265 226 
<< m1 >>
rect 264 225 265 226 
<< m2 >>
rect 264 225 265 226 
<< m1 >>
rect 268 225 269 226 
<< m1 >>
rect 270 225 271 226 
<< m1 >>
rect 272 225 273 226 
<< m1 >>
rect 280 225 281 226 
<< m1 >>
rect 282 225 283 226 
<< m1 >>
rect 298 225 299 226 
<< m2 >>
rect 298 225 299 226 
<< m2c >>
rect 298 225 299 226 
<< m1 >>
rect 298 225 299 226 
<< m2 >>
rect 298 225 299 226 
<< m1 >>
rect 304 225 305 226 
<< m2 >>
rect 304 225 305 226 
<< m2c >>
rect 304 225 305 226 
<< m1 >>
rect 304 225 305 226 
<< m2 >>
rect 304 225 305 226 
<< m1 >>
rect 307 225 308 226 
<< m2 >>
rect 307 225 308 226 
<< m2c >>
rect 307 225 308 226 
<< m1 >>
rect 307 225 308 226 
<< m2 >>
rect 307 225 308 226 
<< m1 >>
rect 316 225 317 226 
<< m2 >>
rect 316 225 317 226 
<< m2c >>
rect 316 225 317 226 
<< m1 >>
rect 316 225 317 226 
<< m2 >>
rect 316 225 317 226 
<< m2 >>
rect 321 225 322 226 
<< m2 >>
rect 322 225 323 226 
<< m2 >>
rect 323 225 324 226 
<< m2 >>
rect 324 225 325 226 
<< m1 >>
rect 325 225 326 226 
<< m2 >>
rect 325 225 326 226 
<< m2 >>
rect 326 225 327 226 
<< m1 >>
rect 327 225 328 226 
<< m2 >>
rect 327 225 328 226 
<< m2 >>
rect 328 225 329 226 
<< m1 >>
rect 329 225 330 226 
<< m2 >>
rect 329 225 330 226 
<< m2 >>
rect 330 225 331 226 
<< m1 >>
rect 331 225 332 226 
<< m2 >>
rect 331 225 332 226 
<< m2 >>
rect 332 225 333 226 
<< m1 >>
rect 333 225 334 226 
<< m2 >>
rect 333 225 334 226 
<< m2c >>
rect 333 225 334 226 
<< m1 >>
rect 333 225 334 226 
<< m2 >>
rect 333 225 334 226 
<< m1 >>
rect 343 225 344 226 
<< m2 >>
rect 343 225 344 226 
<< m2c >>
rect 343 225 344 226 
<< m1 >>
rect 343 225 344 226 
<< m2 >>
rect 343 225 344 226 
<< m1 >>
rect 345 225 346 226 
<< m1 >>
rect 10 226 11 227 
<< m1 >>
rect 13 226 14 227 
<< m1 >>
rect 28 226 29 227 
<< m2 >>
rect 28 226 29 227 
<< m1 >>
rect 37 226 38 227 
<< m1 >>
rect 39 226 40 227 
<< m2 >>
rect 43 226 44 227 
<< m1 >>
rect 44 226 45 227 
<< m1 >>
rect 46 226 47 227 
<< m2 >>
rect 46 226 47 227 
<< m1 >>
rect 56 226 57 227 
<< m1 >>
rect 58 226 59 227 
<< m1 >>
rect 60 226 61 227 
<< m1 >>
rect 62 226 63 227 
<< m1 >>
rect 64 226 65 227 
<< m1 >>
rect 78 226 79 227 
<< m1 >>
rect 80 226 81 227 
<< m1 >>
rect 82 226 83 227 
<< m1 >>
rect 88 226 89 227 
<< m1 >>
rect 118 226 119 227 
<< m1 >>
rect 130 226 131 227 
<< m1 >>
rect 132 226 133 227 
<< m2 >>
rect 132 226 133 227 
<< m1 >>
rect 136 226 137 227 
<< m1 >>
rect 139 226 140 227 
<< m1 >>
rect 140 226 141 227 
<< m1 >>
rect 145 226 146 227 
<< m1 >>
rect 154 226 155 227 
<< m1 >>
rect 163 226 164 227 
<< m1 >>
rect 165 226 166 227 
<< m1 >>
rect 167 226 168 227 
<< m2 >>
rect 168 226 169 227 
<< m1 >>
rect 178 226 179 227 
<< m1 >>
rect 179 226 180 227 
<< m2 >>
rect 179 226 180 227 
<< m2c >>
rect 179 226 180 227 
<< m1 >>
rect 179 226 180 227 
<< m2 >>
rect 179 226 180 227 
<< m2 >>
rect 180 226 181 227 
<< m1 >>
rect 181 226 182 227 
<< m2 >>
rect 181 226 182 227 
<< m2 >>
rect 182 226 183 227 
<< m1 >>
rect 183 226 184 227 
<< m2 >>
rect 183 226 184 227 
<< m2c >>
rect 183 226 184 227 
<< m1 >>
rect 183 226 184 227 
<< m2 >>
rect 183 226 184 227 
<< m1 >>
rect 186 226 187 227 
<< m1 >>
rect 188 226 189 227 
<< m1 >>
rect 190 226 191 227 
<< m1 >>
rect 193 226 194 227 
<< m1 >>
rect 217 226 218 227 
<< m1 >>
rect 219 226 220 227 
<< m2 >>
rect 221 226 222 227 
<< m1 >>
rect 226 226 227 227 
<< m1 >>
rect 235 226 236 227 
<< m1 >>
rect 237 226 238 227 
<< m2 >>
rect 241 226 242 227 
<< m2 >>
rect 243 226 244 227 
<< m1 >>
rect 247 226 248 227 
<< m1 >>
rect 250 226 251 227 
<< m2 >>
rect 253 226 254 227 
<< m2 >>
rect 262 226 263 227 
<< m1 >>
rect 268 226 269 227 
<< m1 >>
rect 270 226 271 227 
<< m2 >>
rect 270 226 271 227 
<< m2c >>
rect 270 226 271 227 
<< m1 >>
rect 270 226 271 227 
<< m2 >>
rect 270 226 271 227 
<< m2 >>
rect 271 226 272 227 
<< m1 >>
rect 272 226 273 227 
<< m2 >>
rect 272 226 273 227 
<< m2 >>
rect 273 226 274 227 
<< m2 >>
rect 279 226 280 227 
<< m1 >>
rect 280 226 281 227 
<< m2 >>
rect 280 226 281 227 
<< m2 >>
rect 281 226 282 227 
<< m1 >>
rect 282 226 283 227 
<< m2 >>
rect 282 226 283 227 
<< m2c >>
rect 282 226 283 227 
<< m1 >>
rect 282 226 283 227 
<< m2 >>
rect 282 226 283 227 
<< m1 >>
rect 298 226 299 227 
<< m1 >>
rect 304 226 305 227 
<< m1 >>
rect 307 226 308 227 
<< m1 >>
rect 316 226 317 227 
<< m1 >>
rect 322 226 323 227 
<< m1 >>
rect 323 226 324 227 
<< m1 >>
rect 324 226 325 227 
<< m1 >>
rect 325 226 326 227 
<< m1 >>
rect 327 226 328 227 
<< m1 >>
rect 329 226 330 227 
<< m1 >>
rect 331 226 332 227 
<< m1 >>
rect 333 226 334 227 
<< m1 >>
rect 343 226 344 227 
<< m1 >>
rect 345 226 346 227 
<< m1 >>
rect 10 227 11 228 
<< m1 >>
rect 13 227 14 228 
<< m1 >>
rect 28 227 29 228 
<< m2 >>
rect 28 227 29 228 
<< m1 >>
rect 37 227 38 228 
<< m1 >>
rect 39 227 40 228 
<< m2 >>
rect 43 227 44 228 
<< m1 >>
rect 44 227 45 228 
<< m1 >>
rect 46 227 47 228 
<< m2 >>
rect 46 227 47 228 
<< m1 >>
rect 56 227 57 228 
<< m1 >>
rect 58 227 59 228 
<< m1 >>
rect 60 227 61 228 
<< m1 >>
rect 62 227 63 228 
<< m1 >>
rect 64 227 65 228 
<< m1 >>
rect 78 227 79 228 
<< m1 >>
rect 80 227 81 228 
<< m1 >>
rect 82 227 83 228 
<< m1 >>
rect 88 227 89 228 
<< m1 >>
rect 118 227 119 228 
<< m1 >>
rect 130 227 131 228 
<< m1 >>
rect 132 227 133 228 
<< m2 >>
rect 132 227 133 228 
<< m1 >>
rect 136 227 137 228 
<< m1 >>
rect 139 227 140 228 
<< m1 >>
rect 145 227 146 228 
<< m1 >>
rect 154 227 155 228 
<< m1 >>
rect 163 227 164 228 
<< m1 >>
rect 165 227 166 228 
<< m1 >>
rect 167 227 168 228 
<< m2 >>
rect 168 227 169 228 
<< m1 >>
rect 178 227 179 228 
<< m1 >>
rect 181 227 182 228 
<< m1 >>
rect 186 227 187 228 
<< m1 >>
rect 188 227 189 228 
<< m1 >>
rect 190 227 191 228 
<< m1 >>
rect 193 227 194 228 
<< m1 >>
rect 217 227 218 228 
<< m1 >>
rect 219 227 220 228 
<< m1 >>
rect 220 227 221 228 
<< m1 >>
rect 221 227 222 228 
<< m2 >>
rect 221 227 222 228 
<< m1 >>
rect 222 227 223 228 
<< m1 >>
rect 223 227 224 228 
<< m1 >>
rect 224 227 225 228 
<< m2 >>
rect 224 227 225 228 
<< m2c >>
rect 224 227 225 228 
<< m1 >>
rect 224 227 225 228 
<< m2 >>
rect 224 227 225 228 
<< m2 >>
rect 225 227 226 228 
<< m1 >>
rect 226 227 227 228 
<< m1 >>
rect 235 227 236 228 
<< m1 >>
rect 237 227 238 228 
<< m1 >>
rect 241 227 242 228 
<< m2 >>
rect 241 227 242 228 
<< m2c >>
rect 241 227 242 228 
<< m1 >>
rect 241 227 242 228 
<< m2 >>
rect 241 227 242 228 
<< m1 >>
rect 243 227 244 228 
<< m2 >>
rect 243 227 244 228 
<< m2c >>
rect 243 227 244 228 
<< m1 >>
rect 243 227 244 228 
<< m2 >>
rect 243 227 244 228 
<< m1 >>
rect 247 227 248 228 
<< m1 >>
rect 250 227 251 228 
<< m1 >>
rect 253 227 254 228 
<< m2 >>
rect 253 227 254 228 
<< m2c >>
rect 253 227 254 228 
<< m1 >>
rect 253 227 254 228 
<< m2 >>
rect 253 227 254 228 
<< m1 >>
rect 262 227 263 228 
<< m2 >>
rect 262 227 263 228 
<< m2c >>
rect 262 227 263 228 
<< m1 >>
rect 262 227 263 228 
<< m2 >>
rect 262 227 263 228 
<< m1 >>
rect 268 227 269 228 
<< m1 >>
rect 272 227 273 228 
<< m2 >>
rect 273 227 274 228 
<< m2 >>
rect 279 227 280 228 
<< m1 >>
rect 280 227 281 228 
<< m1 >>
rect 298 227 299 228 
<< m1 >>
rect 304 227 305 228 
<< m1 >>
rect 307 227 308 228 
<< m1 >>
rect 316 227 317 228 
<< m1 >>
rect 322 227 323 228 
<< m1 >>
rect 327 227 328 228 
<< m1 >>
rect 329 227 330 228 
<< m1 >>
rect 331 227 332 228 
<< m1 >>
rect 333 227 334 228 
<< m1 >>
rect 343 227 344 228 
<< m1 >>
rect 345 227 346 228 
<< m1 >>
rect 10 228 11 229 
<< pdiffusion >>
rect 12 228 13 229 
<< m1 >>
rect 13 228 14 229 
<< pdiffusion >>
rect 13 228 14 229 
<< pdiffusion >>
rect 14 228 15 229 
<< pdiffusion >>
rect 15 228 16 229 
<< pdiffusion >>
rect 16 228 17 229 
<< pdiffusion >>
rect 17 228 18 229 
<< m1 >>
rect 28 228 29 229 
<< m2 >>
rect 28 228 29 229 
<< pdiffusion >>
rect 30 228 31 229 
<< pdiffusion >>
rect 31 228 32 229 
<< pdiffusion >>
rect 32 228 33 229 
<< pdiffusion >>
rect 33 228 34 229 
<< pdiffusion >>
rect 34 228 35 229 
<< pdiffusion >>
rect 35 228 36 229 
<< m1 >>
rect 37 228 38 229 
<< m1 >>
rect 39 228 40 229 
<< m2 >>
rect 43 228 44 229 
<< m1 >>
rect 44 228 45 229 
<< m1 >>
rect 46 228 47 229 
<< m2 >>
rect 46 228 47 229 
<< pdiffusion >>
rect 48 228 49 229 
<< pdiffusion >>
rect 49 228 50 229 
<< pdiffusion >>
rect 50 228 51 229 
<< pdiffusion >>
rect 51 228 52 229 
<< pdiffusion >>
rect 52 228 53 229 
<< pdiffusion >>
rect 53 228 54 229 
<< m1 >>
rect 56 228 57 229 
<< m1 >>
rect 58 228 59 229 
<< m1 >>
rect 60 228 61 229 
<< m1 >>
rect 62 228 63 229 
<< m1 >>
rect 64 228 65 229 
<< pdiffusion >>
rect 66 228 67 229 
<< pdiffusion >>
rect 67 228 68 229 
<< pdiffusion >>
rect 68 228 69 229 
<< pdiffusion >>
rect 69 228 70 229 
<< pdiffusion >>
rect 70 228 71 229 
<< pdiffusion >>
rect 71 228 72 229 
<< m1 >>
rect 78 228 79 229 
<< m1 >>
rect 80 228 81 229 
<< m1 >>
rect 82 228 83 229 
<< pdiffusion >>
rect 84 228 85 229 
<< pdiffusion >>
rect 85 228 86 229 
<< pdiffusion >>
rect 86 228 87 229 
<< pdiffusion >>
rect 87 228 88 229 
<< m1 >>
rect 88 228 89 229 
<< pdiffusion >>
rect 88 228 89 229 
<< pdiffusion >>
rect 89 228 90 229 
<< pdiffusion >>
rect 102 228 103 229 
<< pdiffusion >>
rect 103 228 104 229 
<< pdiffusion >>
rect 104 228 105 229 
<< pdiffusion >>
rect 105 228 106 229 
<< pdiffusion >>
rect 106 228 107 229 
<< pdiffusion >>
rect 107 228 108 229 
<< m1 >>
rect 118 228 119 229 
<< pdiffusion >>
rect 120 228 121 229 
<< pdiffusion >>
rect 121 228 122 229 
<< pdiffusion >>
rect 122 228 123 229 
<< pdiffusion >>
rect 123 228 124 229 
<< pdiffusion >>
rect 124 228 125 229 
<< pdiffusion >>
rect 125 228 126 229 
<< m1 >>
rect 130 228 131 229 
<< m1 >>
rect 132 228 133 229 
<< m2 >>
rect 132 228 133 229 
<< m1 >>
rect 136 228 137 229 
<< pdiffusion >>
rect 138 228 139 229 
<< m1 >>
rect 139 228 140 229 
<< pdiffusion >>
rect 139 228 140 229 
<< pdiffusion >>
rect 140 228 141 229 
<< pdiffusion >>
rect 141 228 142 229 
<< pdiffusion >>
rect 142 228 143 229 
<< pdiffusion >>
rect 143 228 144 229 
<< m1 >>
rect 145 228 146 229 
<< m1 >>
rect 154 228 155 229 
<< pdiffusion >>
rect 156 228 157 229 
<< pdiffusion >>
rect 157 228 158 229 
<< pdiffusion >>
rect 158 228 159 229 
<< pdiffusion >>
rect 159 228 160 229 
<< pdiffusion >>
rect 160 228 161 229 
<< pdiffusion >>
rect 161 228 162 229 
<< m1 >>
rect 163 228 164 229 
<< m1 >>
rect 165 228 166 229 
<< m1 >>
rect 167 228 168 229 
<< m2 >>
rect 168 228 169 229 
<< pdiffusion >>
rect 174 228 175 229 
<< pdiffusion >>
rect 175 228 176 229 
<< pdiffusion >>
rect 176 228 177 229 
<< pdiffusion >>
rect 177 228 178 229 
<< m1 >>
rect 178 228 179 229 
<< pdiffusion >>
rect 178 228 179 229 
<< pdiffusion >>
rect 179 228 180 229 
<< m1 >>
rect 181 228 182 229 
<< m1 >>
rect 186 228 187 229 
<< m1 >>
rect 188 228 189 229 
<< m1 >>
rect 190 228 191 229 
<< pdiffusion >>
rect 192 228 193 229 
<< m1 >>
rect 193 228 194 229 
<< pdiffusion >>
rect 193 228 194 229 
<< pdiffusion >>
rect 194 228 195 229 
<< pdiffusion >>
rect 195 228 196 229 
<< pdiffusion >>
rect 196 228 197 229 
<< pdiffusion >>
rect 197 228 198 229 
<< pdiffusion >>
rect 210 228 211 229 
<< pdiffusion >>
rect 211 228 212 229 
<< pdiffusion >>
rect 212 228 213 229 
<< pdiffusion >>
rect 213 228 214 229 
<< pdiffusion >>
rect 214 228 215 229 
<< pdiffusion >>
rect 215 228 216 229 
<< m1 >>
rect 217 228 218 229 
<< m2 >>
rect 221 228 222 229 
<< m2 >>
rect 225 228 226 229 
<< m1 >>
rect 226 228 227 229 
<< pdiffusion >>
rect 228 228 229 229 
<< pdiffusion >>
rect 229 228 230 229 
<< pdiffusion >>
rect 230 228 231 229 
<< pdiffusion >>
rect 231 228 232 229 
<< pdiffusion >>
rect 232 228 233 229 
<< pdiffusion >>
rect 233 228 234 229 
<< m1 >>
rect 235 228 236 229 
<< m1 >>
rect 237 228 238 229 
<< m1 >>
rect 241 228 242 229 
<< m1 >>
rect 243 228 244 229 
<< pdiffusion >>
rect 246 228 247 229 
<< m1 >>
rect 247 228 248 229 
<< pdiffusion >>
rect 247 228 248 229 
<< pdiffusion >>
rect 248 228 249 229 
<< pdiffusion >>
rect 249 228 250 229 
<< m1 >>
rect 250 228 251 229 
<< pdiffusion >>
rect 250 228 251 229 
<< pdiffusion >>
rect 251 228 252 229 
<< m1 >>
rect 253 228 254 229 
<< m1 >>
rect 262 228 263 229 
<< pdiffusion >>
rect 264 228 265 229 
<< pdiffusion >>
rect 265 228 266 229 
<< pdiffusion >>
rect 266 228 267 229 
<< pdiffusion >>
rect 267 228 268 229 
<< m1 >>
rect 268 228 269 229 
<< pdiffusion >>
rect 268 228 269 229 
<< pdiffusion >>
rect 269 228 270 229 
<< m1 >>
rect 272 228 273 229 
<< m2 >>
rect 273 228 274 229 
<< m2 >>
rect 279 228 280 229 
<< m1 >>
rect 280 228 281 229 
<< pdiffusion >>
rect 282 228 283 229 
<< pdiffusion >>
rect 283 228 284 229 
<< pdiffusion >>
rect 284 228 285 229 
<< pdiffusion >>
rect 285 228 286 229 
<< pdiffusion >>
rect 286 228 287 229 
<< pdiffusion >>
rect 287 228 288 229 
<< m1 >>
rect 298 228 299 229 
<< pdiffusion >>
rect 300 228 301 229 
<< pdiffusion >>
rect 301 228 302 229 
<< pdiffusion >>
rect 302 228 303 229 
<< pdiffusion >>
rect 303 228 304 229 
<< m1 >>
rect 304 228 305 229 
<< pdiffusion >>
rect 304 228 305 229 
<< pdiffusion >>
rect 305 228 306 229 
<< m1 >>
rect 307 228 308 229 
<< m1 >>
rect 316 228 317 229 
<< pdiffusion >>
rect 318 228 319 229 
<< pdiffusion >>
rect 319 228 320 229 
<< pdiffusion >>
rect 320 228 321 229 
<< pdiffusion >>
rect 321 228 322 229 
<< m1 >>
rect 322 228 323 229 
<< pdiffusion >>
rect 322 228 323 229 
<< pdiffusion >>
rect 323 228 324 229 
<< m1 >>
rect 327 228 328 229 
<< m1 >>
rect 329 228 330 229 
<< m1 >>
rect 331 228 332 229 
<< m1 >>
rect 333 228 334 229 
<< pdiffusion >>
rect 336 228 337 229 
<< pdiffusion >>
rect 337 228 338 229 
<< pdiffusion >>
rect 338 228 339 229 
<< pdiffusion >>
rect 339 228 340 229 
<< pdiffusion >>
rect 340 228 341 229 
<< pdiffusion >>
rect 341 228 342 229 
<< m1 >>
rect 343 228 344 229 
<< m1 >>
rect 345 228 346 229 
<< m1 >>
rect 10 229 11 230 
<< pdiffusion >>
rect 12 229 13 230 
<< pdiffusion >>
rect 13 229 14 230 
<< pdiffusion >>
rect 14 229 15 230 
<< pdiffusion >>
rect 15 229 16 230 
<< pdiffusion >>
rect 16 229 17 230 
<< pdiffusion >>
rect 17 229 18 230 
<< m1 >>
rect 28 229 29 230 
<< m2 >>
rect 28 229 29 230 
<< pdiffusion >>
rect 30 229 31 230 
<< pdiffusion >>
rect 31 229 32 230 
<< pdiffusion >>
rect 32 229 33 230 
<< pdiffusion >>
rect 33 229 34 230 
<< pdiffusion >>
rect 34 229 35 230 
<< pdiffusion >>
rect 35 229 36 230 
<< m1 >>
rect 37 229 38 230 
<< m1 >>
rect 39 229 40 230 
<< m2 >>
rect 43 229 44 230 
<< m1 >>
rect 44 229 45 230 
<< m1 >>
rect 46 229 47 230 
<< m2 >>
rect 46 229 47 230 
<< pdiffusion >>
rect 48 229 49 230 
<< pdiffusion >>
rect 49 229 50 230 
<< pdiffusion >>
rect 50 229 51 230 
<< pdiffusion >>
rect 51 229 52 230 
<< pdiffusion >>
rect 52 229 53 230 
<< pdiffusion >>
rect 53 229 54 230 
<< m1 >>
rect 56 229 57 230 
<< m1 >>
rect 58 229 59 230 
<< m1 >>
rect 60 229 61 230 
<< m1 >>
rect 62 229 63 230 
<< m1 >>
rect 64 229 65 230 
<< pdiffusion >>
rect 66 229 67 230 
<< pdiffusion >>
rect 67 229 68 230 
<< pdiffusion >>
rect 68 229 69 230 
<< pdiffusion >>
rect 69 229 70 230 
<< pdiffusion >>
rect 70 229 71 230 
<< pdiffusion >>
rect 71 229 72 230 
<< m1 >>
rect 78 229 79 230 
<< m1 >>
rect 80 229 81 230 
<< m1 >>
rect 82 229 83 230 
<< pdiffusion >>
rect 84 229 85 230 
<< pdiffusion >>
rect 85 229 86 230 
<< pdiffusion >>
rect 86 229 87 230 
<< pdiffusion >>
rect 87 229 88 230 
<< pdiffusion >>
rect 88 229 89 230 
<< pdiffusion >>
rect 89 229 90 230 
<< pdiffusion >>
rect 102 229 103 230 
<< pdiffusion >>
rect 103 229 104 230 
<< pdiffusion >>
rect 104 229 105 230 
<< pdiffusion >>
rect 105 229 106 230 
<< pdiffusion >>
rect 106 229 107 230 
<< pdiffusion >>
rect 107 229 108 230 
<< m1 >>
rect 118 229 119 230 
<< pdiffusion >>
rect 120 229 121 230 
<< pdiffusion >>
rect 121 229 122 230 
<< pdiffusion >>
rect 122 229 123 230 
<< pdiffusion >>
rect 123 229 124 230 
<< pdiffusion >>
rect 124 229 125 230 
<< pdiffusion >>
rect 125 229 126 230 
<< m1 >>
rect 130 229 131 230 
<< m1 >>
rect 132 229 133 230 
<< m2 >>
rect 132 229 133 230 
<< m1 >>
rect 136 229 137 230 
<< pdiffusion >>
rect 138 229 139 230 
<< pdiffusion >>
rect 139 229 140 230 
<< pdiffusion >>
rect 140 229 141 230 
<< pdiffusion >>
rect 141 229 142 230 
<< pdiffusion >>
rect 142 229 143 230 
<< pdiffusion >>
rect 143 229 144 230 
<< m1 >>
rect 145 229 146 230 
<< m1 >>
rect 154 229 155 230 
<< pdiffusion >>
rect 156 229 157 230 
<< pdiffusion >>
rect 157 229 158 230 
<< pdiffusion >>
rect 158 229 159 230 
<< pdiffusion >>
rect 159 229 160 230 
<< pdiffusion >>
rect 160 229 161 230 
<< pdiffusion >>
rect 161 229 162 230 
<< m1 >>
rect 163 229 164 230 
<< m1 >>
rect 165 229 166 230 
<< m1 >>
rect 167 229 168 230 
<< m2 >>
rect 168 229 169 230 
<< pdiffusion >>
rect 174 229 175 230 
<< pdiffusion >>
rect 175 229 176 230 
<< pdiffusion >>
rect 176 229 177 230 
<< pdiffusion >>
rect 177 229 178 230 
<< pdiffusion >>
rect 178 229 179 230 
<< pdiffusion >>
rect 179 229 180 230 
<< m1 >>
rect 181 229 182 230 
<< m1 >>
rect 186 229 187 230 
<< m1 >>
rect 188 229 189 230 
<< m1 >>
rect 190 229 191 230 
<< pdiffusion >>
rect 192 229 193 230 
<< pdiffusion >>
rect 193 229 194 230 
<< pdiffusion >>
rect 194 229 195 230 
<< pdiffusion >>
rect 195 229 196 230 
<< pdiffusion >>
rect 196 229 197 230 
<< pdiffusion >>
rect 197 229 198 230 
<< pdiffusion >>
rect 210 229 211 230 
<< pdiffusion >>
rect 211 229 212 230 
<< pdiffusion >>
rect 212 229 213 230 
<< pdiffusion >>
rect 213 229 214 230 
<< pdiffusion >>
rect 214 229 215 230 
<< pdiffusion >>
rect 215 229 216 230 
<< m1 >>
rect 217 229 218 230 
<< m1 >>
rect 221 229 222 230 
<< m2 >>
rect 221 229 222 230 
<< m2c >>
rect 221 229 222 230 
<< m1 >>
rect 221 229 222 230 
<< m2 >>
rect 221 229 222 230 
<< m2 >>
rect 225 229 226 230 
<< m1 >>
rect 226 229 227 230 
<< pdiffusion >>
rect 228 229 229 230 
<< pdiffusion >>
rect 229 229 230 230 
<< pdiffusion >>
rect 230 229 231 230 
<< pdiffusion >>
rect 231 229 232 230 
<< pdiffusion >>
rect 232 229 233 230 
<< pdiffusion >>
rect 233 229 234 230 
<< m1 >>
rect 235 229 236 230 
<< m1 >>
rect 237 229 238 230 
<< m1 >>
rect 241 229 242 230 
<< m1 >>
rect 243 229 244 230 
<< pdiffusion >>
rect 246 229 247 230 
<< pdiffusion >>
rect 247 229 248 230 
<< pdiffusion >>
rect 248 229 249 230 
<< pdiffusion >>
rect 249 229 250 230 
<< pdiffusion >>
rect 250 229 251 230 
<< pdiffusion >>
rect 251 229 252 230 
<< m1 >>
rect 253 229 254 230 
<< m1 >>
rect 262 229 263 230 
<< pdiffusion >>
rect 264 229 265 230 
<< pdiffusion >>
rect 265 229 266 230 
<< pdiffusion >>
rect 266 229 267 230 
<< pdiffusion >>
rect 267 229 268 230 
<< pdiffusion >>
rect 268 229 269 230 
<< pdiffusion >>
rect 269 229 270 230 
<< m1 >>
rect 272 229 273 230 
<< m2 >>
rect 273 229 274 230 
<< m2 >>
rect 279 229 280 230 
<< m1 >>
rect 280 229 281 230 
<< pdiffusion >>
rect 282 229 283 230 
<< pdiffusion >>
rect 283 229 284 230 
<< pdiffusion >>
rect 284 229 285 230 
<< pdiffusion >>
rect 285 229 286 230 
<< pdiffusion >>
rect 286 229 287 230 
<< pdiffusion >>
rect 287 229 288 230 
<< m1 >>
rect 298 229 299 230 
<< pdiffusion >>
rect 300 229 301 230 
<< pdiffusion >>
rect 301 229 302 230 
<< pdiffusion >>
rect 302 229 303 230 
<< pdiffusion >>
rect 303 229 304 230 
<< pdiffusion >>
rect 304 229 305 230 
<< pdiffusion >>
rect 305 229 306 230 
<< m1 >>
rect 307 229 308 230 
<< m1 >>
rect 316 229 317 230 
<< pdiffusion >>
rect 318 229 319 230 
<< pdiffusion >>
rect 319 229 320 230 
<< pdiffusion >>
rect 320 229 321 230 
<< pdiffusion >>
rect 321 229 322 230 
<< pdiffusion >>
rect 322 229 323 230 
<< pdiffusion >>
rect 323 229 324 230 
<< m1 >>
rect 327 229 328 230 
<< m1 >>
rect 329 229 330 230 
<< m1 >>
rect 331 229 332 230 
<< m1 >>
rect 333 229 334 230 
<< pdiffusion >>
rect 336 229 337 230 
<< pdiffusion >>
rect 337 229 338 230 
<< pdiffusion >>
rect 338 229 339 230 
<< pdiffusion >>
rect 339 229 340 230 
<< pdiffusion >>
rect 340 229 341 230 
<< pdiffusion >>
rect 341 229 342 230 
<< m1 >>
rect 343 229 344 230 
<< m1 >>
rect 345 229 346 230 
<< m1 >>
rect 10 230 11 231 
<< pdiffusion >>
rect 12 230 13 231 
<< pdiffusion >>
rect 13 230 14 231 
<< pdiffusion >>
rect 14 230 15 231 
<< pdiffusion >>
rect 15 230 16 231 
<< pdiffusion >>
rect 16 230 17 231 
<< pdiffusion >>
rect 17 230 18 231 
<< m1 >>
rect 28 230 29 231 
<< m2 >>
rect 28 230 29 231 
<< pdiffusion >>
rect 30 230 31 231 
<< pdiffusion >>
rect 31 230 32 231 
<< pdiffusion >>
rect 32 230 33 231 
<< pdiffusion >>
rect 33 230 34 231 
<< pdiffusion >>
rect 34 230 35 231 
<< pdiffusion >>
rect 35 230 36 231 
<< m1 >>
rect 37 230 38 231 
<< m1 >>
rect 39 230 40 231 
<< m2 >>
rect 43 230 44 231 
<< m1 >>
rect 44 230 45 231 
<< m1 >>
rect 46 230 47 231 
<< m2 >>
rect 46 230 47 231 
<< pdiffusion >>
rect 48 230 49 231 
<< pdiffusion >>
rect 49 230 50 231 
<< pdiffusion >>
rect 50 230 51 231 
<< pdiffusion >>
rect 51 230 52 231 
<< pdiffusion >>
rect 52 230 53 231 
<< pdiffusion >>
rect 53 230 54 231 
<< m1 >>
rect 56 230 57 231 
<< m1 >>
rect 58 230 59 231 
<< m1 >>
rect 60 230 61 231 
<< m1 >>
rect 62 230 63 231 
<< m1 >>
rect 64 230 65 231 
<< pdiffusion >>
rect 66 230 67 231 
<< pdiffusion >>
rect 67 230 68 231 
<< pdiffusion >>
rect 68 230 69 231 
<< pdiffusion >>
rect 69 230 70 231 
<< pdiffusion >>
rect 70 230 71 231 
<< pdiffusion >>
rect 71 230 72 231 
<< m1 >>
rect 78 230 79 231 
<< m1 >>
rect 80 230 81 231 
<< m1 >>
rect 82 230 83 231 
<< pdiffusion >>
rect 84 230 85 231 
<< pdiffusion >>
rect 85 230 86 231 
<< pdiffusion >>
rect 86 230 87 231 
<< pdiffusion >>
rect 87 230 88 231 
<< pdiffusion >>
rect 88 230 89 231 
<< pdiffusion >>
rect 89 230 90 231 
<< pdiffusion >>
rect 102 230 103 231 
<< pdiffusion >>
rect 103 230 104 231 
<< pdiffusion >>
rect 104 230 105 231 
<< pdiffusion >>
rect 105 230 106 231 
<< pdiffusion >>
rect 106 230 107 231 
<< pdiffusion >>
rect 107 230 108 231 
<< m1 >>
rect 118 230 119 231 
<< pdiffusion >>
rect 120 230 121 231 
<< pdiffusion >>
rect 121 230 122 231 
<< pdiffusion >>
rect 122 230 123 231 
<< pdiffusion >>
rect 123 230 124 231 
<< pdiffusion >>
rect 124 230 125 231 
<< pdiffusion >>
rect 125 230 126 231 
<< m1 >>
rect 130 230 131 231 
<< m1 >>
rect 132 230 133 231 
<< m2 >>
rect 132 230 133 231 
<< m1 >>
rect 136 230 137 231 
<< pdiffusion >>
rect 138 230 139 231 
<< pdiffusion >>
rect 139 230 140 231 
<< pdiffusion >>
rect 140 230 141 231 
<< pdiffusion >>
rect 141 230 142 231 
<< pdiffusion >>
rect 142 230 143 231 
<< pdiffusion >>
rect 143 230 144 231 
<< m1 >>
rect 145 230 146 231 
<< m1 >>
rect 154 230 155 231 
<< pdiffusion >>
rect 156 230 157 231 
<< pdiffusion >>
rect 157 230 158 231 
<< pdiffusion >>
rect 158 230 159 231 
<< pdiffusion >>
rect 159 230 160 231 
<< pdiffusion >>
rect 160 230 161 231 
<< pdiffusion >>
rect 161 230 162 231 
<< m1 >>
rect 163 230 164 231 
<< m1 >>
rect 165 230 166 231 
<< m1 >>
rect 167 230 168 231 
<< m2 >>
rect 168 230 169 231 
<< pdiffusion >>
rect 174 230 175 231 
<< pdiffusion >>
rect 175 230 176 231 
<< pdiffusion >>
rect 176 230 177 231 
<< pdiffusion >>
rect 177 230 178 231 
<< pdiffusion >>
rect 178 230 179 231 
<< pdiffusion >>
rect 179 230 180 231 
<< m1 >>
rect 181 230 182 231 
<< m1 >>
rect 186 230 187 231 
<< m1 >>
rect 188 230 189 231 
<< m1 >>
rect 190 230 191 231 
<< pdiffusion >>
rect 192 230 193 231 
<< pdiffusion >>
rect 193 230 194 231 
<< pdiffusion >>
rect 194 230 195 231 
<< pdiffusion >>
rect 195 230 196 231 
<< pdiffusion >>
rect 196 230 197 231 
<< pdiffusion >>
rect 197 230 198 231 
<< pdiffusion >>
rect 210 230 211 231 
<< pdiffusion >>
rect 211 230 212 231 
<< pdiffusion >>
rect 212 230 213 231 
<< pdiffusion >>
rect 213 230 214 231 
<< pdiffusion >>
rect 214 230 215 231 
<< pdiffusion >>
rect 215 230 216 231 
<< m1 >>
rect 217 230 218 231 
<< m1 >>
rect 221 230 222 231 
<< m2 >>
rect 225 230 226 231 
<< m1 >>
rect 226 230 227 231 
<< pdiffusion >>
rect 228 230 229 231 
<< pdiffusion >>
rect 229 230 230 231 
<< pdiffusion >>
rect 230 230 231 231 
<< pdiffusion >>
rect 231 230 232 231 
<< pdiffusion >>
rect 232 230 233 231 
<< pdiffusion >>
rect 233 230 234 231 
<< m1 >>
rect 235 230 236 231 
<< m1 >>
rect 237 230 238 231 
<< m1 >>
rect 241 230 242 231 
<< m1 >>
rect 243 230 244 231 
<< pdiffusion >>
rect 246 230 247 231 
<< pdiffusion >>
rect 247 230 248 231 
<< pdiffusion >>
rect 248 230 249 231 
<< pdiffusion >>
rect 249 230 250 231 
<< pdiffusion >>
rect 250 230 251 231 
<< pdiffusion >>
rect 251 230 252 231 
<< m1 >>
rect 253 230 254 231 
<< m1 >>
rect 262 230 263 231 
<< pdiffusion >>
rect 264 230 265 231 
<< pdiffusion >>
rect 265 230 266 231 
<< pdiffusion >>
rect 266 230 267 231 
<< pdiffusion >>
rect 267 230 268 231 
<< pdiffusion >>
rect 268 230 269 231 
<< pdiffusion >>
rect 269 230 270 231 
<< m1 >>
rect 272 230 273 231 
<< m2 >>
rect 273 230 274 231 
<< m2 >>
rect 279 230 280 231 
<< m1 >>
rect 280 230 281 231 
<< pdiffusion >>
rect 282 230 283 231 
<< pdiffusion >>
rect 283 230 284 231 
<< pdiffusion >>
rect 284 230 285 231 
<< pdiffusion >>
rect 285 230 286 231 
<< pdiffusion >>
rect 286 230 287 231 
<< pdiffusion >>
rect 287 230 288 231 
<< m1 >>
rect 298 230 299 231 
<< pdiffusion >>
rect 300 230 301 231 
<< pdiffusion >>
rect 301 230 302 231 
<< pdiffusion >>
rect 302 230 303 231 
<< pdiffusion >>
rect 303 230 304 231 
<< pdiffusion >>
rect 304 230 305 231 
<< pdiffusion >>
rect 305 230 306 231 
<< m1 >>
rect 307 230 308 231 
<< m1 >>
rect 316 230 317 231 
<< pdiffusion >>
rect 318 230 319 231 
<< pdiffusion >>
rect 319 230 320 231 
<< pdiffusion >>
rect 320 230 321 231 
<< pdiffusion >>
rect 321 230 322 231 
<< pdiffusion >>
rect 322 230 323 231 
<< pdiffusion >>
rect 323 230 324 231 
<< m1 >>
rect 327 230 328 231 
<< m1 >>
rect 329 230 330 231 
<< m1 >>
rect 331 230 332 231 
<< m1 >>
rect 333 230 334 231 
<< pdiffusion >>
rect 336 230 337 231 
<< pdiffusion >>
rect 337 230 338 231 
<< pdiffusion >>
rect 338 230 339 231 
<< pdiffusion >>
rect 339 230 340 231 
<< pdiffusion >>
rect 340 230 341 231 
<< pdiffusion >>
rect 341 230 342 231 
<< m1 >>
rect 343 230 344 231 
<< m1 >>
rect 345 230 346 231 
<< m1 >>
rect 10 231 11 232 
<< pdiffusion >>
rect 12 231 13 232 
<< pdiffusion >>
rect 13 231 14 232 
<< pdiffusion >>
rect 14 231 15 232 
<< pdiffusion >>
rect 15 231 16 232 
<< pdiffusion >>
rect 16 231 17 232 
<< pdiffusion >>
rect 17 231 18 232 
<< m1 >>
rect 28 231 29 232 
<< m2 >>
rect 28 231 29 232 
<< pdiffusion >>
rect 30 231 31 232 
<< pdiffusion >>
rect 31 231 32 232 
<< pdiffusion >>
rect 32 231 33 232 
<< pdiffusion >>
rect 33 231 34 232 
<< pdiffusion >>
rect 34 231 35 232 
<< pdiffusion >>
rect 35 231 36 232 
<< m1 >>
rect 37 231 38 232 
<< m1 >>
rect 39 231 40 232 
<< m2 >>
rect 43 231 44 232 
<< m1 >>
rect 44 231 45 232 
<< m1 >>
rect 46 231 47 232 
<< m2 >>
rect 46 231 47 232 
<< pdiffusion >>
rect 48 231 49 232 
<< pdiffusion >>
rect 49 231 50 232 
<< pdiffusion >>
rect 50 231 51 232 
<< pdiffusion >>
rect 51 231 52 232 
<< pdiffusion >>
rect 52 231 53 232 
<< pdiffusion >>
rect 53 231 54 232 
<< m1 >>
rect 56 231 57 232 
<< m1 >>
rect 58 231 59 232 
<< m1 >>
rect 60 231 61 232 
<< m1 >>
rect 62 231 63 232 
<< m1 >>
rect 64 231 65 232 
<< pdiffusion >>
rect 66 231 67 232 
<< pdiffusion >>
rect 67 231 68 232 
<< pdiffusion >>
rect 68 231 69 232 
<< pdiffusion >>
rect 69 231 70 232 
<< pdiffusion >>
rect 70 231 71 232 
<< pdiffusion >>
rect 71 231 72 232 
<< m1 >>
rect 78 231 79 232 
<< m1 >>
rect 80 231 81 232 
<< m1 >>
rect 82 231 83 232 
<< pdiffusion >>
rect 84 231 85 232 
<< pdiffusion >>
rect 85 231 86 232 
<< pdiffusion >>
rect 86 231 87 232 
<< pdiffusion >>
rect 87 231 88 232 
<< pdiffusion >>
rect 88 231 89 232 
<< pdiffusion >>
rect 89 231 90 232 
<< pdiffusion >>
rect 102 231 103 232 
<< pdiffusion >>
rect 103 231 104 232 
<< pdiffusion >>
rect 104 231 105 232 
<< pdiffusion >>
rect 105 231 106 232 
<< pdiffusion >>
rect 106 231 107 232 
<< pdiffusion >>
rect 107 231 108 232 
<< m1 >>
rect 118 231 119 232 
<< pdiffusion >>
rect 120 231 121 232 
<< pdiffusion >>
rect 121 231 122 232 
<< pdiffusion >>
rect 122 231 123 232 
<< pdiffusion >>
rect 123 231 124 232 
<< pdiffusion >>
rect 124 231 125 232 
<< pdiffusion >>
rect 125 231 126 232 
<< m1 >>
rect 130 231 131 232 
<< m1 >>
rect 132 231 133 232 
<< m2 >>
rect 132 231 133 232 
<< m1 >>
rect 136 231 137 232 
<< pdiffusion >>
rect 138 231 139 232 
<< pdiffusion >>
rect 139 231 140 232 
<< pdiffusion >>
rect 140 231 141 232 
<< pdiffusion >>
rect 141 231 142 232 
<< pdiffusion >>
rect 142 231 143 232 
<< pdiffusion >>
rect 143 231 144 232 
<< m1 >>
rect 145 231 146 232 
<< m1 >>
rect 154 231 155 232 
<< pdiffusion >>
rect 156 231 157 232 
<< pdiffusion >>
rect 157 231 158 232 
<< pdiffusion >>
rect 158 231 159 232 
<< pdiffusion >>
rect 159 231 160 232 
<< pdiffusion >>
rect 160 231 161 232 
<< pdiffusion >>
rect 161 231 162 232 
<< m1 >>
rect 163 231 164 232 
<< m1 >>
rect 165 231 166 232 
<< m1 >>
rect 167 231 168 232 
<< m2 >>
rect 168 231 169 232 
<< pdiffusion >>
rect 174 231 175 232 
<< pdiffusion >>
rect 175 231 176 232 
<< pdiffusion >>
rect 176 231 177 232 
<< pdiffusion >>
rect 177 231 178 232 
<< pdiffusion >>
rect 178 231 179 232 
<< pdiffusion >>
rect 179 231 180 232 
<< m1 >>
rect 181 231 182 232 
<< m1 >>
rect 186 231 187 232 
<< m1 >>
rect 188 231 189 232 
<< m1 >>
rect 190 231 191 232 
<< pdiffusion >>
rect 192 231 193 232 
<< pdiffusion >>
rect 193 231 194 232 
<< pdiffusion >>
rect 194 231 195 232 
<< pdiffusion >>
rect 195 231 196 232 
<< pdiffusion >>
rect 196 231 197 232 
<< pdiffusion >>
rect 197 231 198 232 
<< pdiffusion >>
rect 210 231 211 232 
<< pdiffusion >>
rect 211 231 212 232 
<< pdiffusion >>
rect 212 231 213 232 
<< pdiffusion >>
rect 213 231 214 232 
<< pdiffusion >>
rect 214 231 215 232 
<< pdiffusion >>
rect 215 231 216 232 
<< m1 >>
rect 217 231 218 232 
<< m1 >>
rect 221 231 222 232 
<< m2 >>
rect 225 231 226 232 
<< m1 >>
rect 226 231 227 232 
<< pdiffusion >>
rect 228 231 229 232 
<< pdiffusion >>
rect 229 231 230 232 
<< pdiffusion >>
rect 230 231 231 232 
<< pdiffusion >>
rect 231 231 232 232 
<< pdiffusion >>
rect 232 231 233 232 
<< pdiffusion >>
rect 233 231 234 232 
<< m1 >>
rect 235 231 236 232 
<< m1 >>
rect 237 231 238 232 
<< m1 >>
rect 241 231 242 232 
<< m1 >>
rect 243 231 244 232 
<< pdiffusion >>
rect 246 231 247 232 
<< pdiffusion >>
rect 247 231 248 232 
<< pdiffusion >>
rect 248 231 249 232 
<< pdiffusion >>
rect 249 231 250 232 
<< pdiffusion >>
rect 250 231 251 232 
<< pdiffusion >>
rect 251 231 252 232 
<< m1 >>
rect 253 231 254 232 
<< m1 >>
rect 262 231 263 232 
<< pdiffusion >>
rect 264 231 265 232 
<< pdiffusion >>
rect 265 231 266 232 
<< pdiffusion >>
rect 266 231 267 232 
<< pdiffusion >>
rect 267 231 268 232 
<< pdiffusion >>
rect 268 231 269 232 
<< pdiffusion >>
rect 269 231 270 232 
<< m1 >>
rect 272 231 273 232 
<< m2 >>
rect 273 231 274 232 
<< m2 >>
rect 279 231 280 232 
<< m1 >>
rect 280 231 281 232 
<< pdiffusion >>
rect 282 231 283 232 
<< pdiffusion >>
rect 283 231 284 232 
<< pdiffusion >>
rect 284 231 285 232 
<< pdiffusion >>
rect 285 231 286 232 
<< pdiffusion >>
rect 286 231 287 232 
<< pdiffusion >>
rect 287 231 288 232 
<< m1 >>
rect 298 231 299 232 
<< pdiffusion >>
rect 300 231 301 232 
<< pdiffusion >>
rect 301 231 302 232 
<< pdiffusion >>
rect 302 231 303 232 
<< pdiffusion >>
rect 303 231 304 232 
<< pdiffusion >>
rect 304 231 305 232 
<< pdiffusion >>
rect 305 231 306 232 
<< m1 >>
rect 307 231 308 232 
<< m1 >>
rect 316 231 317 232 
<< pdiffusion >>
rect 318 231 319 232 
<< pdiffusion >>
rect 319 231 320 232 
<< pdiffusion >>
rect 320 231 321 232 
<< pdiffusion >>
rect 321 231 322 232 
<< pdiffusion >>
rect 322 231 323 232 
<< pdiffusion >>
rect 323 231 324 232 
<< m1 >>
rect 327 231 328 232 
<< m1 >>
rect 329 231 330 232 
<< m1 >>
rect 331 231 332 232 
<< m1 >>
rect 333 231 334 232 
<< pdiffusion >>
rect 336 231 337 232 
<< pdiffusion >>
rect 337 231 338 232 
<< pdiffusion >>
rect 338 231 339 232 
<< pdiffusion >>
rect 339 231 340 232 
<< pdiffusion >>
rect 340 231 341 232 
<< pdiffusion >>
rect 341 231 342 232 
<< m1 >>
rect 343 231 344 232 
<< m1 >>
rect 345 231 346 232 
<< m1 >>
rect 10 232 11 233 
<< pdiffusion >>
rect 12 232 13 233 
<< pdiffusion >>
rect 13 232 14 233 
<< pdiffusion >>
rect 14 232 15 233 
<< pdiffusion >>
rect 15 232 16 233 
<< pdiffusion >>
rect 16 232 17 233 
<< pdiffusion >>
rect 17 232 18 233 
<< m1 >>
rect 28 232 29 233 
<< m2 >>
rect 28 232 29 233 
<< pdiffusion >>
rect 30 232 31 233 
<< pdiffusion >>
rect 31 232 32 233 
<< pdiffusion >>
rect 32 232 33 233 
<< pdiffusion >>
rect 33 232 34 233 
<< pdiffusion >>
rect 34 232 35 233 
<< pdiffusion >>
rect 35 232 36 233 
<< m1 >>
rect 37 232 38 233 
<< m1 >>
rect 39 232 40 233 
<< m2 >>
rect 43 232 44 233 
<< m1 >>
rect 44 232 45 233 
<< m1 >>
rect 46 232 47 233 
<< m2 >>
rect 46 232 47 233 
<< pdiffusion >>
rect 48 232 49 233 
<< pdiffusion >>
rect 49 232 50 233 
<< pdiffusion >>
rect 50 232 51 233 
<< pdiffusion >>
rect 51 232 52 233 
<< pdiffusion >>
rect 52 232 53 233 
<< pdiffusion >>
rect 53 232 54 233 
<< m1 >>
rect 56 232 57 233 
<< m1 >>
rect 58 232 59 233 
<< m1 >>
rect 60 232 61 233 
<< m1 >>
rect 62 232 63 233 
<< m1 >>
rect 64 232 65 233 
<< pdiffusion >>
rect 66 232 67 233 
<< pdiffusion >>
rect 67 232 68 233 
<< pdiffusion >>
rect 68 232 69 233 
<< pdiffusion >>
rect 69 232 70 233 
<< pdiffusion >>
rect 70 232 71 233 
<< pdiffusion >>
rect 71 232 72 233 
<< m1 >>
rect 78 232 79 233 
<< m1 >>
rect 80 232 81 233 
<< m1 >>
rect 82 232 83 233 
<< pdiffusion >>
rect 84 232 85 233 
<< pdiffusion >>
rect 85 232 86 233 
<< pdiffusion >>
rect 86 232 87 233 
<< pdiffusion >>
rect 87 232 88 233 
<< pdiffusion >>
rect 88 232 89 233 
<< pdiffusion >>
rect 89 232 90 233 
<< pdiffusion >>
rect 102 232 103 233 
<< pdiffusion >>
rect 103 232 104 233 
<< pdiffusion >>
rect 104 232 105 233 
<< pdiffusion >>
rect 105 232 106 233 
<< pdiffusion >>
rect 106 232 107 233 
<< pdiffusion >>
rect 107 232 108 233 
<< m1 >>
rect 118 232 119 233 
<< pdiffusion >>
rect 120 232 121 233 
<< pdiffusion >>
rect 121 232 122 233 
<< pdiffusion >>
rect 122 232 123 233 
<< pdiffusion >>
rect 123 232 124 233 
<< pdiffusion >>
rect 124 232 125 233 
<< pdiffusion >>
rect 125 232 126 233 
<< m1 >>
rect 130 232 131 233 
<< m1 >>
rect 132 232 133 233 
<< m2 >>
rect 132 232 133 233 
<< m1 >>
rect 136 232 137 233 
<< pdiffusion >>
rect 138 232 139 233 
<< pdiffusion >>
rect 139 232 140 233 
<< pdiffusion >>
rect 140 232 141 233 
<< pdiffusion >>
rect 141 232 142 233 
<< pdiffusion >>
rect 142 232 143 233 
<< pdiffusion >>
rect 143 232 144 233 
<< m1 >>
rect 145 232 146 233 
<< m1 >>
rect 154 232 155 233 
<< pdiffusion >>
rect 156 232 157 233 
<< pdiffusion >>
rect 157 232 158 233 
<< pdiffusion >>
rect 158 232 159 233 
<< pdiffusion >>
rect 159 232 160 233 
<< pdiffusion >>
rect 160 232 161 233 
<< pdiffusion >>
rect 161 232 162 233 
<< m1 >>
rect 163 232 164 233 
<< m1 >>
rect 165 232 166 233 
<< m1 >>
rect 167 232 168 233 
<< m2 >>
rect 168 232 169 233 
<< pdiffusion >>
rect 174 232 175 233 
<< pdiffusion >>
rect 175 232 176 233 
<< pdiffusion >>
rect 176 232 177 233 
<< pdiffusion >>
rect 177 232 178 233 
<< pdiffusion >>
rect 178 232 179 233 
<< pdiffusion >>
rect 179 232 180 233 
<< m1 >>
rect 181 232 182 233 
<< m1 >>
rect 186 232 187 233 
<< m1 >>
rect 188 232 189 233 
<< m1 >>
rect 190 232 191 233 
<< pdiffusion >>
rect 192 232 193 233 
<< pdiffusion >>
rect 193 232 194 233 
<< pdiffusion >>
rect 194 232 195 233 
<< pdiffusion >>
rect 195 232 196 233 
<< pdiffusion >>
rect 196 232 197 233 
<< pdiffusion >>
rect 197 232 198 233 
<< pdiffusion >>
rect 210 232 211 233 
<< pdiffusion >>
rect 211 232 212 233 
<< pdiffusion >>
rect 212 232 213 233 
<< pdiffusion >>
rect 213 232 214 233 
<< pdiffusion >>
rect 214 232 215 233 
<< pdiffusion >>
rect 215 232 216 233 
<< m1 >>
rect 217 232 218 233 
<< m1 >>
rect 221 232 222 233 
<< m2 >>
rect 225 232 226 233 
<< m1 >>
rect 226 232 227 233 
<< pdiffusion >>
rect 228 232 229 233 
<< pdiffusion >>
rect 229 232 230 233 
<< pdiffusion >>
rect 230 232 231 233 
<< pdiffusion >>
rect 231 232 232 233 
<< pdiffusion >>
rect 232 232 233 233 
<< pdiffusion >>
rect 233 232 234 233 
<< m1 >>
rect 235 232 236 233 
<< m1 >>
rect 237 232 238 233 
<< m1 >>
rect 241 232 242 233 
<< m1 >>
rect 243 232 244 233 
<< pdiffusion >>
rect 246 232 247 233 
<< pdiffusion >>
rect 247 232 248 233 
<< pdiffusion >>
rect 248 232 249 233 
<< pdiffusion >>
rect 249 232 250 233 
<< pdiffusion >>
rect 250 232 251 233 
<< pdiffusion >>
rect 251 232 252 233 
<< m1 >>
rect 253 232 254 233 
<< m1 >>
rect 262 232 263 233 
<< pdiffusion >>
rect 264 232 265 233 
<< pdiffusion >>
rect 265 232 266 233 
<< pdiffusion >>
rect 266 232 267 233 
<< pdiffusion >>
rect 267 232 268 233 
<< pdiffusion >>
rect 268 232 269 233 
<< pdiffusion >>
rect 269 232 270 233 
<< m1 >>
rect 272 232 273 233 
<< m2 >>
rect 273 232 274 233 
<< m2 >>
rect 279 232 280 233 
<< m1 >>
rect 280 232 281 233 
<< pdiffusion >>
rect 282 232 283 233 
<< pdiffusion >>
rect 283 232 284 233 
<< pdiffusion >>
rect 284 232 285 233 
<< pdiffusion >>
rect 285 232 286 233 
<< pdiffusion >>
rect 286 232 287 233 
<< pdiffusion >>
rect 287 232 288 233 
<< m1 >>
rect 298 232 299 233 
<< pdiffusion >>
rect 300 232 301 233 
<< pdiffusion >>
rect 301 232 302 233 
<< pdiffusion >>
rect 302 232 303 233 
<< pdiffusion >>
rect 303 232 304 233 
<< pdiffusion >>
rect 304 232 305 233 
<< pdiffusion >>
rect 305 232 306 233 
<< m1 >>
rect 307 232 308 233 
<< m1 >>
rect 316 232 317 233 
<< pdiffusion >>
rect 318 232 319 233 
<< pdiffusion >>
rect 319 232 320 233 
<< pdiffusion >>
rect 320 232 321 233 
<< pdiffusion >>
rect 321 232 322 233 
<< pdiffusion >>
rect 322 232 323 233 
<< pdiffusion >>
rect 323 232 324 233 
<< m1 >>
rect 327 232 328 233 
<< m1 >>
rect 329 232 330 233 
<< m1 >>
rect 331 232 332 233 
<< m1 >>
rect 333 232 334 233 
<< pdiffusion >>
rect 336 232 337 233 
<< pdiffusion >>
rect 337 232 338 233 
<< pdiffusion >>
rect 338 232 339 233 
<< pdiffusion >>
rect 339 232 340 233 
<< pdiffusion >>
rect 340 232 341 233 
<< pdiffusion >>
rect 341 232 342 233 
<< m1 >>
rect 343 232 344 233 
<< m1 >>
rect 345 232 346 233 
<< m1 >>
rect 10 233 11 234 
<< pdiffusion >>
rect 12 233 13 234 
<< pdiffusion >>
rect 13 233 14 234 
<< pdiffusion >>
rect 14 233 15 234 
<< pdiffusion >>
rect 15 233 16 234 
<< pdiffusion >>
rect 16 233 17 234 
<< pdiffusion >>
rect 17 233 18 234 
<< m1 >>
rect 28 233 29 234 
<< m2 >>
rect 28 233 29 234 
<< pdiffusion >>
rect 30 233 31 234 
<< pdiffusion >>
rect 31 233 32 234 
<< pdiffusion >>
rect 32 233 33 234 
<< pdiffusion >>
rect 33 233 34 234 
<< pdiffusion >>
rect 34 233 35 234 
<< pdiffusion >>
rect 35 233 36 234 
<< m1 >>
rect 37 233 38 234 
<< m1 >>
rect 39 233 40 234 
<< m2 >>
rect 43 233 44 234 
<< m1 >>
rect 44 233 45 234 
<< m1 >>
rect 46 233 47 234 
<< m2 >>
rect 46 233 47 234 
<< pdiffusion >>
rect 48 233 49 234 
<< pdiffusion >>
rect 49 233 50 234 
<< pdiffusion >>
rect 50 233 51 234 
<< pdiffusion >>
rect 51 233 52 234 
<< pdiffusion >>
rect 52 233 53 234 
<< pdiffusion >>
rect 53 233 54 234 
<< m1 >>
rect 56 233 57 234 
<< m1 >>
rect 58 233 59 234 
<< m1 >>
rect 60 233 61 234 
<< m1 >>
rect 62 233 63 234 
<< m1 >>
rect 64 233 65 234 
<< pdiffusion >>
rect 66 233 67 234 
<< pdiffusion >>
rect 67 233 68 234 
<< pdiffusion >>
rect 68 233 69 234 
<< pdiffusion >>
rect 69 233 70 234 
<< pdiffusion >>
rect 70 233 71 234 
<< pdiffusion >>
rect 71 233 72 234 
<< m1 >>
rect 78 233 79 234 
<< m1 >>
rect 80 233 81 234 
<< m1 >>
rect 82 233 83 234 
<< pdiffusion >>
rect 84 233 85 234 
<< pdiffusion >>
rect 85 233 86 234 
<< pdiffusion >>
rect 86 233 87 234 
<< pdiffusion >>
rect 87 233 88 234 
<< pdiffusion >>
rect 88 233 89 234 
<< pdiffusion >>
rect 89 233 90 234 
<< pdiffusion >>
rect 102 233 103 234 
<< pdiffusion >>
rect 103 233 104 234 
<< pdiffusion >>
rect 104 233 105 234 
<< pdiffusion >>
rect 105 233 106 234 
<< pdiffusion >>
rect 106 233 107 234 
<< pdiffusion >>
rect 107 233 108 234 
<< m1 >>
rect 118 233 119 234 
<< pdiffusion >>
rect 120 233 121 234 
<< pdiffusion >>
rect 121 233 122 234 
<< pdiffusion >>
rect 122 233 123 234 
<< pdiffusion >>
rect 123 233 124 234 
<< pdiffusion >>
rect 124 233 125 234 
<< pdiffusion >>
rect 125 233 126 234 
<< m1 >>
rect 130 233 131 234 
<< m1 >>
rect 132 233 133 234 
<< m2 >>
rect 132 233 133 234 
<< m1 >>
rect 136 233 137 234 
<< pdiffusion >>
rect 138 233 139 234 
<< pdiffusion >>
rect 139 233 140 234 
<< pdiffusion >>
rect 140 233 141 234 
<< pdiffusion >>
rect 141 233 142 234 
<< pdiffusion >>
rect 142 233 143 234 
<< pdiffusion >>
rect 143 233 144 234 
<< m1 >>
rect 145 233 146 234 
<< m1 >>
rect 154 233 155 234 
<< pdiffusion >>
rect 156 233 157 234 
<< pdiffusion >>
rect 157 233 158 234 
<< pdiffusion >>
rect 158 233 159 234 
<< pdiffusion >>
rect 159 233 160 234 
<< m1 >>
rect 160 233 161 234 
<< pdiffusion >>
rect 160 233 161 234 
<< pdiffusion >>
rect 161 233 162 234 
<< m1 >>
rect 163 233 164 234 
<< m1 >>
rect 165 233 166 234 
<< m1 >>
rect 167 233 168 234 
<< m2 >>
rect 168 233 169 234 
<< pdiffusion >>
rect 174 233 175 234 
<< pdiffusion >>
rect 175 233 176 234 
<< pdiffusion >>
rect 176 233 177 234 
<< pdiffusion >>
rect 177 233 178 234 
<< pdiffusion >>
rect 178 233 179 234 
<< pdiffusion >>
rect 179 233 180 234 
<< m1 >>
rect 181 233 182 234 
<< m1 >>
rect 186 233 187 234 
<< m1 >>
rect 188 233 189 234 
<< m1 >>
rect 190 233 191 234 
<< pdiffusion >>
rect 192 233 193 234 
<< pdiffusion >>
rect 193 233 194 234 
<< pdiffusion >>
rect 194 233 195 234 
<< pdiffusion >>
rect 195 233 196 234 
<< pdiffusion >>
rect 196 233 197 234 
<< pdiffusion >>
rect 197 233 198 234 
<< pdiffusion >>
rect 210 233 211 234 
<< pdiffusion >>
rect 211 233 212 234 
<< pdiffusion >>
rect 212 233 213 234 
<< pdiffusion >>
rect 213 233 214 234 
<< m1 >>
rect 214 233 215 234 
<< pdiffusion >>
rect 214 233 215 234 
<< pdiffusion >>
rect 215 233 216 234 
<< m1 >>
rect 217 233 218 234 
<< m1 >>
rect 221 233 222 234 
<< m2 >>
rect 225 233 226 234 
<< m1 >>
rect 226 233 227 234 
<< pdiffusion >>
rect 228 233 229 234 
<< pdiffusion >>
rect 229 233 230 234 
<< pdiffusion >>
rect 230 233 231 234 
<< pdiffusion >>
rect 231 233 232 234 
<< pdiffusion >>
rect 232 233 233 234 
<< pdiffusion >>
rect 233 233 234 234 
<< m1 >>
rect 235 233 236 234 
<< m1 >>
rect 237 233 238 234 
<< m1 >>
rect 241 233 242 234 
<< m1 >>
rect 243 233 244 234 
<< pdiffusion >>
rect 246 233 247 234 
<< pdiffusion >>
rect 247 233 248 234 
<< pdiffusion >>
rect 248 233 249 234 
<< pdiffusion >>
rect 249 233 250 234 
<< pdiffusion >>
rect 250 233 251 234 
<< pdiffusion >>
rect 251 233 252 234 
<< m1 >>
rect 253 233 254 234 
<< m1 >>
rect 262 233 263 234 
<< pdiffusion >>
rect 264 233 265 234 
<< pdiffusion >>
rect 265 233 266 234 
<< pdiffusion >>
rect 266 233 267 234 
<< pdiffusion >>
rect 267 233 268 234 
<< pdiffusion >>
rect 268 233 269 234 
<< pdiffusion >>
rect 269 233 270 234 
<< m1 >>
rect 272 233 273 234 
<< m2 >>
rect 273 233 274 234 
<< m2 >>
rect 279 233 280 234 
<< m1 >>
rect 280 233 281 234 
<< pdiffusion >>
rect 282 233 283 234 
<< pdiffusion >>
rect 283 233 284 234 
<< pdiffusion >>
rect 284 233 285 234 
<< pdiffusion >>
rect 285 233 286 234 
<< pdiffusion >>
rect 286 233 287 234 
<< pdiffusion >>
rect 287 233 288 234 
<< m1 >>
rect 298 233 299 234 
<< pdiffusion >>
rect 300 233 301 234 
<< pdiffusion >>
rect 301 233 302 234 
<< pdiffusion >>
rect 302 233 303 234 
<< pdiffusion >>
rect 303 233 304 234 
<< pdiffusion >>
rect 304 233 305 234 
<< pdiffusion >>
rect 305 233 306 234 
<< m1 >>
rect 307 233 308 234 
<< m1 >>
rect 316 233 317 234 
<< pdiffusion >>
rect 318 233 319 234 
<< m1 >>
rect 319 233 320 234 
<< pdiffusion >>
rect 319 233 320 234 
<< pdiffusion >>
rect 320 233 321 234 
<< pdiffusion >>
rect 321 233 322 234 
<< pdiffusion >>
rect 322 233 323 234 
<< pdiffusion >>
rect 323 233 324 234 
<< m1 >>
rect 327 233 328 234 
<< m1 >>
rect 329 233 330 234 
<< m1 >>
rect 331 233 332 234 
<< m1 >>
rect 333 233 334 234 
<< pdiffusion >>
rect 336 233 337 234 
<< pdiffusion >>
rect 337 233 338 234 
<< pdiffusion >>
rect 338 233 339 234 
<< pdiffusion >>
rect 339 233 340 234 
<< pdiffusion >>
rect 340 233 341 234 
<< pdiffusion >>
rect 341 233 342 234 
<< m1 >>
rect 343 233 344 234 
<< m1 >>
rect 345 233 346 234 
<< m1 >>
rect 10 234 11 235 
<< m1 >>
rect 28 234 29 235 
<< m2 >>
rect 28 234 29 235 
<< m1 >>
rect 37 234 38 235 
<< m1 >>
rect 39 234 40 235 
<< m2 >>
rect 43 234 44 235 
<< m1 >>
rect 44 234 45 235 
<< m1 >>
rect 46 234 47 235 
<< m2 >>
rect 46 234 47 235 
<< m1 >>
rect 56 234 57 235 
<< m1 >>
rect 58 234 59 235 
<< m1 >>
rect 60 234 61 235 
<< m1 >>
rect 62 234 63 235 
<< m1 >>
rect 64 234 65 235 
<< m1 >>
rect 78 234 79 235 
<< m1 >>
rect 80 234 81 235 
<< m1 >>
rect 82 234 83 235 
<< m1 >>
rect 118 234 119 235 
<< m1 >>
rect 130 234 131 235 
<< m1 >>
rect 132 234 133 235 
<< m2 >>
rect 132 234 133 235 
<< m1 >>
rect 136 234 137 235 
<< m1 >>
rect 145 234 146 235 
<< m1 >>
rect 154 234 155 235 
<< m1 >>
rect 160 234 161 235 
<< m1 >>
rect 163 234 164 235 
<< m1 >>
rect 165 234 166 235 
<< m1 >>
rect 167 234 168 235 
<< m2 >>
rect 168 234 169 235 
<< m1 >>
rect 181 234 182 235 
<< m1 >>
rect 186 234 187 235 
<< m1 >>
rect 188 234 189 235 
<< m1 >>
rect 190 234 191 235 
<< m1 >>
rect 214 234 215 235 
<< m1 >>
rect 217 234 218 235 
<< m1 >>
rect 221 234 222 235 
<< m2 >>
rect 225 234 226 235 
<< m1 >>
rect 226 234 227 235 
<< m1 >>
rect 235 234 236 235 
<< m1 >>
rect 237 234 238 235 
<< m1 >>
rect 241 234 242 235 
<< m1 >>
rect 243 234 244 235 
<< m1 >>
rect 253 234 254 235 
<< m1 >>
rect 262 234 263 235 
<< m1 >>
rect 272 234 273 235 
<< m2 >>
rect 273 234 274 235 
<< m2 >>
rect 279 234 280 235 
<< m1 >>
rect 280 234 281 235 
<< m1 >>
rect 298 234 299 235 
<< m1 >>
rect 307 234 308 235 
<< m1 >>
rect 316 234 317 235 
<< m1 >>
rect 319 234 320 235 
<< m1 >>
rect 327 234 328 235 
<< m1 >>
rect 329 234 330 235 
<< m1 >>
rect 331 234 332 235 
<< m1 >>
rect 333 234 334 235 
<< m1 >>
rect 343 234 344 235 
<< m1 >>
rect 345 234 346 235 
<< m1 >>
rect 10 235 11 236 
<< m1 >>
rect 28 235 29 236 
<< m2 >>
rect 28 235 29 236 
<< m1 >>
rect 37 235 38 236 
<< m1 >>
rect 39 235 40 236 
<< m2 >>
rect 43 235 44 236 
<< m1 >>
rect 44 235 45 236 
<< m1 >>
rect 46 235 47 236 
<< m2 >>
rect 46 235 47 236 
<< m1 >>
rect 56 235 57 236 
<< m1 >>
rect 58 235 59 236 
<< m1 >>
rect 60 235 61 236 
<< m1 >>
rect 62 235 63 236 
<< m1 >>
rect 64 235 65 236 
<< m1 >>
rect 78 235 79 236 
<< m1 >>
rect 80 235 81 236 
<< m1 >>
rect 82 235 83 236 
<< m1 >>
rect 118 235 119 236 
<< m1 >>
rect 130 235 131 236 
<< m1 >>
rect 132 235 133 236 
<< m2 >>
rect 132 235 133 236 
<< m1 >>
rect 136 235 137 236 
<< m1 >>
rect 145 235 146 236 
<< m1 >>
rect 154 235 155 236 
<< m1 >>
rect 160 235 161 236 
<< m1 >>
rect 163 235 164 236 
<< m1 >>
rect 165 235 166 236 
<< m1 >>
rect 167 235 168 236 
<< m2 >>
rect 168 235 169 236 
<< m1 >>
rect 181 235 182 236 
<< m1 >>
rect 186 235 187 236 
<< m1 >>
rect 188 235 189 236 
<< m1 >>
rect 190 235 191 236 
<< m1 >>
rect 214 235 215 236 
<< m1 >>
rect 215 235 216 236 
<< m1 >>
rect 216 235 217 236 
<< m1 >>
rect 217 235 218 236 
<< m1 >>
rect 221 235 222 236 
<< m2 >>
rect 225 235 226 236 
<< m1 >>
rect 226 235 227 236 
<< m2 >>
rect 226 235 227 236 
<< m2 >>
rect 227 235 228 236 
<< m1 >>
rect 228 235 229 236 
<< m2 >>
rect 228 235 229 236 
<< m2c >>
rect 228 235 229 236 
<< m1 >>
rect 228 235 229 236 
<< m2 >>
rect 228 235 229 236 
<< m1 >>
rect 235 235 236 236 
<< m1 >>
rect 237 235 238 236 
<< m1 >>
rect 241 235 242 236 
<< m1 >>
rect 243 235 244 236 
<< m1 >>
rect 253 235 254 236 
<< m1 >>
rect 262 235 263 236 
<< m1 >>
rect 272 235 273 236 
<< m2 >>
rect 273 235 274 236 
<< m2 >>
rect 279 235 280 236 
<< m1 >>
rect 280 235 281 236 
<< m1 >>
rect 298 235 299 236 
<< m1 >>
rect 307 235 308 236 
<< m1 >>
rect 316 235 317 236 
<< m1 >>
rect 319 235 320 236 
<< m1 >>
rect 327 235 328 236 
<< m1 >>
rect 329 235 330 236 
<< m1 >>
rect 331 235 332 236 
<< m1 >>
rect 333 235 334 236 
<< m1 >>
rect 343 235 344 236 
<< m1 >>
rect 345 235 346 236 
<< m1 >>
rect 10 236 11 237 
<< m1 >>
rect 28 236 29 237 
<< m2 >>
rect 28 236 29 237 
<< m1 >>
rect 37 236 38 237 
<< m1 >>
rect 39 236 40 237 
<< m2 >>
rect 43 236 44 237 
<< m1 >>
rect 44 236 45 237 
<< m1 >>
rect 46 236 47 237 
<< m2 >>
rect 46 236 47 237 
<< m1 >>
rect 56 236 57 237 
<< m1 >>
rect 58 236 59 237 
<< m1 >>
rect 60 236 61 237 
<< m1 >>
rect 62 236 63 237 
<< m1 >>
rect 64 236 65 237 
<< m1 >>
rect 78 236 79 237 
<< m1 >>
rect 80 236 81 237 
<< m1 >>
rect 82 236 83 237 
<< m1 >>
rect 118 236 119 237 
<< m1 >>
rect 130 236 131 237 
<< m1 >>
rect 132 236 133 237 
<< m2 >>
rect 132 236 133 237 
<< m1 >>
rect 136 236 137 237 
<< m1 >>
rect 145 236 146 237 
<< m1 >>
rect 154 236 155 237 
<< m1 >>
rect 160 236 161 237 
<< m1 >>
rect 163 236 164 237 
<< m1 >>
rect 165 236 166 237 
<< m1 >>
rect 167 236 168 237 
<< m2 >>
rect 168 236 169 237 
<< m1 >>
rect 181 236 182 237 
<< m1 >>
rect 186 236 187 237 
<< m1 >>
rect 188 236 189 237 
<< m1 >>
rect 190 236 191 237 
<< m1 >>
rect 221 236 222 237 
<< m1 >>
rect 226 236 227 237 
<< m1 >>
rect 228 236 229 237 
<< m1 >>
rect 230 236 231 237 
<< m2 >>
rect 230 236 231 237 
<< m2c >>
rect 230 236 231 237 
<< m1 >>
rect 230 236 231 237 
<< m2 >>
rect 230 236 231 237 
<< m1 >>
rect 231 236 232 237 
<< m1 >>
rect 232 236 233 237 
<< m1 >>
rect 233 236 234 237 
<< m2 >>
rect 233 236 234 237 
<< m2c >>
rect 233 236 234 237 
<< m1 >>
rect 233 236 234 237 
<< m2 >>
rect 233 236 234 237 
<< m2 >>
rect 234 236 235 237 
<< m1 >>
rect 235 236 236 237 
<< m2 >>
rect 235 236 236 237 
<< m2 >>
rect 236 236 237 237 
<< m1 >>
rect 237 236 238 237 
<< m2 >>
rect 237 236 238 237 
<< m2 >>
rect 238 236 239 237 
<< m1 >>
rect 239 236 240 237 
<< m2 >>
rect 239 236 240 237 
<< m2c >>
rect 239 236 240 237 
<< m1 >>
rect 239 236 240 237 
<< m2 >>
rect 239 236 240 237 
<< m2 >>
rect 240 236 241 237 
<< m1 >>
rect 241 236 242 237 
<< m2 >>
rect 241 236 242 237 
<< m2 >>
rect 242 236 243 237 
<< m1 >>
rect 243 236 244 237 
<< m2 >>
rect 243 236 244 237 
<< m2 >>
rect 244 236 245 237 
<< m1 >>
rect 245 236 246 237 
<< m2 >>
rect 245 236 246 237 
<< m2c >>
rect 245 236 246 237 
<< m1 >>
rect 245 236 246 237 
<< m2 >>
rect 245 236 246 237 
<< m1 >>
rect 253 236 254 237 
<< m1 >>
rect 262 236 263 237 
<< m1 >>
rect 272 236 273 237 
<< m2 >>
rect 273 236 274 237 
<< m2 >>
rect 279 236 280 237 
<< m1 >>
rect 280 236 281 237 
<< m1 >>
rect 298 236 299 237 
<< m1 >>
rect 307 236 308 237 
<< m1 >>
rect 316 236 317 237 
<< m1 >>
rect 319 236 320 237 
<< m1 >>
rect 320 236 321 237 
<< m1 >>
rect 321 236 322 237 
<< m1 >>
rect 322 236 323 237 
<< m1 >>
rect 323 236 324 237 
<< m1 >>
rect 324 236 325 237 
<< m1 >>
rect 325 236 326 237 
<< m2 >>
rect 325 236 326 237 
<< m2c >>
rect 325 236 326 237 
<< m1 >>
rect 325 236 326 237 
<< m2 >>
rect 325 236 326 237 
<< m2 >>
rect 326 236 327 237 
<< m1 >>
rect 327 236 328 237 
<< m2 >>
rect 327 236 328 237 
<< m2 >>
rect 328 236 329 237 
<< m1 >>
rect 329 236 330 237 
<< m2 >>
rect 329 236 330 237 
<< m2 >>
rect 330 236 331 237 
<< m1 >>
rect 331 236 332 237 
<< m2 >>
rect 331 236 332 237 
<< m2c >>
rect 331 236 332 237 
<< m1 >>
rect 331 236 332 237 
<< m2 >>
rect 331 236 332 237 
<< m1 >>
rect 333 236 334 237 
<< m2 >>
rect 333 236 334 237 
<< m2c >>
rect 333 236 334 237 
<< m1 >>
rect 333 236 334 237 
<< m2 >>
rect 333 236 334 237 
<< m1 >>
rect 343 236 344 237 
<< m1 >>
rect 345 236 346 237 
<< m1 >>
rect 10 237 11 238 
<< m1 >>
rect 28 237 29 238 
<< m2 >>
rect 28 237 29 238 
<< m1 >>
rect 37 237 38 238 
<< m1 >>
rect 39 237 40 238 
<< m2 >>
rect 43 237 44 238 
<< m1 >>
rect 44 237 45 238 
<< m1 >>
rect 46 237 47 238 
<< m2 >>
rect 46 237 47 238 
<< m1 >>
rect 56 237 57 238 
<< m1 >>
rect 58 237 59 238 
<< m1 >>
rect 60 237 61 238 
<< m1 >>
rect 62 237 63 238 
<< m1 >>
rect 64 237 65 238 
<< m1 >>
rect 78 237 79 238 
<< m1 >>
rect 80 237 81 238 
<< m1 >>
rect 82 237 83 238 
<< m1 >>
rect 118 237 119 238 
<< m1 >>
rect 130 237 131 238 
<< m1 >>
rect 132 237 133 238 
<< m2 >>
rect 132 237 133 238 
<< m1 >>
rect 136 237 137 238 
<< m1 >>
rect 145 237 146 238 
<< m1 >>
rect 154 237 155 238 
<< m1 >>
rect 160 237 161 238 
<< m1 >>
rect 163 237 164 238 
<< m1 >>
rect 165 237 166 238 
<< m1 >>
rect 167 237 168 238 
<< m2 >>
rect 168 237 169 238 
<< m1 >>
rect 181 237 182 238 
<< m1 >>
rect 183 237 184 238 
<< m1 >>
rect 184 237 185 238 
<< m2 >>
rect 184 237 185 238 
<< m2c >>
rect 184 237 185 238 
<< m1 >>
rect 184 237 185 238 
<< m2 >>
rect 184 237 185 238 
<< m2 >>
rect 185 237 186 238 
<< m1 >>
rect 186 237 187 238 
<< m2 >>
rect 186 237 187 238 
<< m2 >>
rect 187 237 188 238 
<< m1 >>
rect 188 237 189 238 
<< m2 >>
rect 188 237 189 238 
<< m2 >>
rect 189 237 190 238 
<< m1 >>
rect 190 237 191 238 
<< m2 >>
rect 190 237 191 238 
<< m2 >>
rect 191 237 192 238 
<< m1 >>
rect 192 237 193 238 
<< m2 >>
rect 192 237 193 238 
<< m2c >>
rect 192 237 193 238 
<< m1 >>
rect 192 237 193 238 
<< m2 >>
rect 192 237 193 238 
<< m1 >>
rect 221 237 222 238 
<< m1 >>
rect 222 237 223 238 
<< m1 >>
rect 223 237 224 238 
<< m1 >>
rect 224 237 225 238 
<< m2 >>
rect 224 237 225 238 
<< m2c >>
rect 224 237 225 238 
<< m1 >>
rect 224 237 225 238 
<< m2 >>
rect 224 237 225 238 
<< m2 >>
rect 225 237 226 238 
<< m1 >>
rect 226 237 227 238 
<< m1 >>
rect 228 237 229 238 
<< m2 >>
rect 230 237 231 238 
<< m1 >>
rect 235 237 236 238 
<< m1 >>
rect 237 237 238 238 
<< m1 >>
rect 241 237 242 238 
<< m1 >>
rect 243 237 244 238 
<< m1 >>
rect 245 237 246 238 
<< m1 >>
rect 253 237 254 238 
<< m1 >>
rect 262 237 263 238 
<< m1 >>
rect 272 237 273 238 
<< m2 >>
rect 273 237 274 238 
<< m2 >>
rect 279 237 280 238 
<< m1 >>
rect 280 237 281 238 
<< m1 >>
rect 298 237 299 238 
<< m1 >>
rect 307 237 308 238 
<< m1 >>
rect 316 237 317 238 
<< m1 >>
rect 327 237 328 238 
<< m1 >>
rect 329 237 330 238 
<< m2 >>
rect 333 237 334 238 
<< m1 >>
rect 343 237 344 238 
<< m1 >>
rect 345 237 346 238 
<< m1 >>
rect 10 238 11 239 
<< m1 >>
rect 28 238 29 239 
<< m2 >>
rect 28 238 29 239 
<< m1 >>
rect 37 238 38 239 
<< m1 >>
rect 39 238 40 239 
<< m2 >>
rect 43 238 44 239 
<< m1 >>
rect 44 238 45 239 
<< m1 >>
rect 46 238 47 239 
<< m2 >>
rect 46 238 47 239 
<< m1 >>
rect 56 238 57 239 
<< m1 >>
rect 58 238 59 239 
<< m1 >>
rect 60 238 61 239 
<< m1 >>
rect 62 238 63 239 
<< m1 >>
rect 64 238 65 239 
<< m1 >>
rect 78 238 79 239 
<< m1 >>
rect 80 238 81 239 
<< m1 >>
rect 82 238 83 239 
<< m1 >>
rect 118 238 119 239 
<< m1 >>
rect 130 238 131 239 
<< m1 >>
rect 132 238 133 239 
<< m2 >>
rect 132 238 133 239 
<< m1 >>
rect 136 238 137 239 
<< m1 >>
rect 145 238 146 239 
<< m1 >>
rect 154 238 155 239 
<< m1 >>
rect 160 238 161 239 
<< m1 >>
rect 163 238 164 239 
<< m1 >>
rect 165 238 166 239 
<< m1 >>
rect 167 238 168 239 
<< m2 >>
rect 168 238 169 239 
<< m1 >>
rect 181 238 182 239 
<< m1 >>
rect 183 238 184 239 
<< m1 >>
rect 186 238 187 239 
<< m1 >>
rect 188 238 189 239 
<< m1 >>
rect 190 238 191 239 
<< m1 >>
rect 192 238 193 239 
<< m2 >>
rect 225 238 226 239 
<< m1 >>
rect 226 238 227 239 
<< m2 >>
rect 226 238 227 239 
<< m2 >>
rect 227 238 228 239 
<< m1 >>
rect 228 238 229 239 
<< m2 >>
rect 228 238 229 239 
<< m1 >>
rect 229 238 230 239 
<< m2 >>
rect 229 238 230 239 
<< m1 >>
rect 230 238 231 239 
<< m2 >>
rect 230 238 231 239 
<< m1 >>
rect 231 238 232 239 
<< m1 >>
rect 232 238 233 239 
<< m1 >>
rect 233 238 234 239 
<< m2 >>
rect 233 238 234 239 
<< m2c >>
rect 233 238 234 239 
<< m1 >>
rect 233 238 234 239 
<< m2 >>
rect 233 238 234 239 
<< m2 >>
rect 234 238 235 239 
<< m1 >>
rect 235 238 236 239 
<< m2 >>
rect 235 238 236 239 
<< m2 >>
rect 236 238 237 239 
<< m1 >>
rect 237 238 238 239 
<< m2 >>
rect 237 238 238 239 
<< m2 >>
rect 238 238 239 239 
<< m1 >>
rect 239 238 240 239 
<< m2 >>
rect 239 238 240 239 
<< m2c >>
rect 239 238 240 239 
<< m1 >>
rect 239 238 240 239 
<< m2 >>
rect 239 238 240 239 
<< m1 >>
rect 241 238 242 239 
<< m1 >>
rect 243 238 244 239 
<< m1 >>
rect 245 238 246 239 
<< m1 >>
rect 246 238 247 239 
<< m1 >>
rect 247 238 248 239 
<< m1 >>
rect 248 238 249 239 
<< m1 >>
rect 249 238 250 239 
<< m1 >>
rect 250 238 251 239 
<< m1 >>
rect 251 238 252 239 
<< m1 >>
rect 252 238 253 239 
<< m1 >>
rect 253 238 254 239 
<< m1 >>
rect 262 238 263 239 
<< m1 >>
rect 272 238 273 239 
<< m2 >>
rect 273 238 274 239 
<< m2 >>
rect 279 238 280 239 
<< m1 >>
rect 280 238 281 239 
<< m1 >>
rect 294 238 295 239 
<< m1 >>
rect 295 238 296 239 
<< m1 >>
rect 296 238 297 239 
<< m2 >>
rect 296 238 297 239 
<< m2c >>
rect 296 238 297 239 
<< m1 >>
rect 296 238 297 239 
<< m2 >>
rect 296 238 297 239 
<< m2 >>
rect 297 238 298 239 
<< m1 >>
rect 298 238 299 239 
<< m2 >>
rect 298 238 299 239 
<< m2 >>
rect 299 238 300 239 
<< m1 >>
rect 300 238 301 239 
<< m2 >>
rect 300 238 301 239 
<< m2c >>
rect 300 238 301 239 
<< m1 >>
rect 300 238 301 239 
<< m2 >>
rect 300 238 301 239 
<< m1 >>
rect 301 238 302 239 
<< m1 >>
rect 302 238 303 239 
<< m1 >>
rect 303 238 304 239 
<< m1 >>
rect 304 238 305 239 
<< m1 >>
rect 305 238 306 239 
<< m1 >>
rect 306 238 307 239 
<< m1 >>
rect 307 238 308 239 
<< m1 >>
rect 316 238 317 239 
<< m1 >>
rect 327 238 328 239 
<< m1 >>
rect 329 238 330 239 
<< m2 >>
rect 330 238 331 239 
<< m1 >>
rect 331 238 332 239 
<< m2 >>
rect 331 238 332 239 
<< m2c >>
rect 331 238 332 239 
<< m1 >>
rect 331 238 332 239 
<< m2 >>
rect 331 238 332 239 
<< m1 >>
rect 332 238 333 239 
<< m1 >>
rect 333 238 334 239 
<< m2 >>
rect 333 238 334 239 
<< m1 >>
rect 334 238 335 239 
<< m2 >>
rect 334 238 335 239 
<< m1 >>
rect 335 238 336 239 
<< m2 >>
rect 335 238 336 239 
<< m1 >>
rect 336 238 337 239 
<< m2 >>
rect 336 238 337 239 
<< m1 >>
rect 337 238 338 239 
<< m2 >>
rect 337 238 338 239 
<< m1 >>
rect 338 238 339 239 
<< m2 >>
rect 338 238 339 239 
<< m1 >>
rect 339 238 340 239 
<< m2 >>
rect 339 238 340 239 
<< m1 >>
rect 340 238 341 239 
<< m2 >>
rect 340 238 341 239 
<< m1 >>
rect 341 238 342 239 
<< m2 >>
rect 341 238 342 239 
<< m1 >>
rect 342 238 343 239 
<< m2 >>
rect 342 238 343 239 
<< m1 >>
rect 343 238 344 239 
<< m2 >>
rect 343 238 344 239 
<< m2 >>
rect 344 238 345 239 
<< m1 >>
rect 345 238 346 239 
<< m2 >>
rect 345 238 346 239 
<< m2c >>
rect 345 238 346 239 
<< m1 >>
rect 345 238 346 239 
<< m2 >>
rect 345 238 346 239 
<< m1 >>
rect 10 239 11 240 
<< m1 >>
rect 28 239 29 240 
<< m2 >>
rect 28 239 29 240 
<< m1 >>
rect 37 239 38 240 
<< m1 >>
rect 39 239 40 240 
<< m2 >>
rect 43 239 44 240 
<< m1 >>
rect 44 239 45 240 
<< m1 >>
rect 46 239 47 240 
<< m2 >>
rect 46 239 47 240 
<< m1 >>
rect 56 239 57 240 
<< m2 >>
rect 56 239 57 240 
<< m2c >>
rect 56 239 57 240 
<< m1 >>
rect 56 239 57 240 
<< m2 >>
rect 56 239 57 240 
<< m1 >>
rect 58 239 59 240 
<< m2 >>
rect 58 239 59 240 
<< m2c >>
rect 58 239 59 240 
<< m1 >>
rect 58 239 59 240 
<< m2 >>
rect 58 239 59 240 
<< m1 >>
rect 60 239 61 240 
<< m2 >>
rect 60 239 61 240 
<< m2c >>
rect 60 239 61 240 
<< m1 >>
rect 60 239 61 240 
<< m2 >>
rect 60 239 61 240 
<< m1 >>
rect 62 239 63 240 
<< m2 >>
rect 62 239 63 240 
<< m2c >>
rect 62 239 63 240 
<< m1 >>
rect 62 239 63 240 
<< m2 >>
rect 62 239 63 240 
<< m1 >>
rect 64 239 65 240 
<< m2 >>
rect 64 239 65 240 
<< m2c >>
rect 64 239 65 240 
<< m1 >>
rect 64 239 65 240 
<< m2 >>
rect 64 239 65 240 
<< m1 >>
rect 78 239 79 240 
<< m2 >>
rect 78 239 79 240 
<< m2c >>
rect 78 239 79 240 
<< m1 >>
rect 78 239 79 240 
<< m2 >>
rect 78 239 79 240 
<< m1 >>
rect 80 239 81 240 
<< m2 >>
rect 80 239 81 240 
<< m2c >>
rect 80 239 81 240 
<< m1 >>
rect 80 239 81 240 
<< m2 >>
rect 80 239 81 240 
<< m2 >>
rect 81 239 82 240 
<< m1 >>
rect 82 239 83 240 
<< m2 >>
rect 82 239 83 240 
<< m1 >>
rect 83 239 84 240 
<< m2 >>
rect 83 239 84 240 
<< m1 >>
rect 84 239 85 240 
<< m2 >>
rect 84 239 85 240 
<< m1 >>
rect 85 239 86 240 
<< m2 >>
rect 85 239 86 240 
<< m1 >>
rect 86 239 87 240 
<< m2 >>
rect 86 239 87 240 
<< m1 >>
rect 87 239 88 240 
<< m2 >>
rect 87 239 88 240 
<< m1 >>
rect 88 239 89 240 
<< m2 >>
rect 88 239 89 240 
<< m1 >>
rect 89 239 90 240 
<< m2 >>
rect 89 239 90 240 
<< m1 >>
rect 90 239 91 240 
<< m2 >>
rect 90 239 91 240 
<< m1 >>
rect 91 239 92 240 
<< m2 >>
rect 91 239 92 240 
<< m1 >>
rect 92 239 93 240 
<< m2 >>
rect 92 239 93 240 
<< m1 >>
rect 93 239 94 240 
<< m2 >>
rect 93 239 94 240 
<< m1 >>
rect 94 239 95 240 
<< m2 >>
rect 94 239 95 240 
<< m1 >>
rect 95 239 96 240 
<< m2 >>
rect 95 239 96 240 
<< m1 >>
rect 96 239 97 240 
<< m2 >>
rect 96 239 97 240 
<< m1 >>
rect 97 239 98 240 
<< m2 >>
rect 97 239 98 240 
<< m1 >>
rect 98 239 99 240 
<< m2 >>
rect 98 239 99 240 
<< m1 >>
rect 99 239 100 240 
<< m2 >>
rect 99 239 100 240 
<< m1 >>
rect 100 239 101 240 
<< m2 >>
rect 100 239 101 240 
<< m1 >>
rect 101 239 102 240 
<< m2 >>
rect 101 239 102 240 
<< m1 >>
rect 102 239 103 240 
<< m2 >>
rect 102 239 103 240 
<< m1 >>
rect 103 239 104 240 
<< m2 >>
rect 103 239 104 240 
<< m1 >>
rect 104 239 105 240 
<< m2 >>
rect 104 239 105 240 
<< m1 >>
rect 105 239 106 240 
<< m2 >>
rect 105 239 106 240 
<< m1 >>
rect 106 239 107 240 
<< m2 >>
rect 106 239 107 240 
<< m1 >>
rect 107 239 108 240 
<< m2 >>
rect 107 239 108 240 
<< m1 >>
rect 108 239 109 240 
<< m2 >>
rect 108 239 109 240 
<< m1 >>
rect 109 239 110 240 
<< m2 >>
rect 109 239 110 240 
<< m1 >>
rect 110 239 111 240 
<< m2 >>
rect 110 239 111 240 
<< m1 >>
rect 111 239 112 240 
<< m2 >>
rect 111 239 112 240 
<< m1 >>
rect 112 239 113 240 
<< m2 >>
rect 112 239 113 240 
<< m1 >>
rect 113 239 114 240 
<< m2 >>
rect 113 239 114 240 
<< m1 >>
rect 114 239 115 240 
<< m2 >>
rect 114 239 115 240 
<< m1 >>
rect 115 239 116 240 
<< m1 >>
rect 116 239 117 240 
<< m2 >>
rect 116 239 117 240 
<< m2c >>
rect 116 239 117 240 
<< m1 >>
rect 116 239 117 240 
<< m2 >>
rect 116 239 117 240 
<< m2 >>
rect 117 239 118 240 
<< m1 >>
rect 118 239 119 240 
<< m2 >>
rect 118 239 119 240 
<< m1 >>
rect 119 239 120 240 
<< m1 >>
rect 120 239 121 240 
<< m1 >>
rect 121 239 122 240 
<< m1 >>
rect 122 239 123 240 
<< m1 >>
rect 123 239 124 240 
<< m1 >>
rect 124 239 125 240 
<< m1 >>
rect 125 239 126 240 
<< m1 >>
rect 126 239 127 240 
<< m1 >>
rect 127 239 128 240 
<< m1 >>
rect 128 239 129 240 
<< m2 >>
rect 128 239 129 240 
<< m2c >>
rect 128 239 129 240 
<< m1 >>
rect 128 239 129 240 
<< m2 >>
rect 128 239 129 240 
<< m1 >>
rect 130 239 131 240 
<< m2 >>
rect 130 239 131 240 
<< m2c >>
rect 130 239 131 240 
<< m1 >>
rect 130 239 131 240 
<< m2 >>
rect 130 239 131 240 
<< m1 >>
rect 132 239 133 240 
<< m2 >>
rect 132 239 133 240 
<< m1 >>
rect 133 239 134 240 
<< m1 >>
rect 134 239 135 240 
<< m2 >>
rect 134 239 135 240 
<< m2c >>
rect 134 239 135 240 
<< m1 >>
rect 134 239 135 240 
<< m2 >>
rect 134 239 135 240 
<< m1 >>
rect 136 239 137 240 
<< m2 >>
rect 136 239 137 240 
<< m2c >>
rect 136 239 137 240 
<< m1 >>
rect 136 239 137 240 
<< m2 >>
rect 136 239 137 240 
<< m1 >>
rect 145 239 146 240 
<< m1 >>
rect 154 239 155 240 
<< m2 >>
rect 154 239 155 240 
<< m2c >>
rect 154 239 155 240 
<< m1 >>
rect 154 239 155 240 
<< m2 >>
rect 154 239 155 240 
<< m1 >>
rect 160 239 161 240 
<< m2 >>
rect 160 239 161 240 
<< m2c >>
rect 160 239 161 240 
<< m1 >>
rect 160 239 161 240 
<< m2 >>
rect 160 239 161 240 
<< m1 >>
rect 163 239 164 240 
<< m1 >>
rect 165 239 166 240 
<< m1 >>
rect 167 239 168 240 
<< m2 >>
rect 168 239 169 240 
<< m1 >>
rect 181 239 182 240 
<< m2 >>
rect 181 239 182 240 
<< m2c >>
rect 181 239 182 240 
<< m1 >>
rect 181 239 182 240 
<< m2 >>
rect 181 239 182 240 
<< m1 >>
rect 183 239 184 240 
<< m2 >>
rect 183 239 184 240 
<< m2c >>
rect 183 239 184 240 
<< m1 >>
rect 183 239 184 240 
<< m2 >>
rect 183 239 184 240 
<< m1 >>
rect 186 239 187 240 
<< m2 >>
rect 186 239 187 240 
<< m2c >>
rect 186 239 187 240 
<< m1 >>
rect 186 239 187 240 
<< m2 >>
rect 186 239 187 240 
<< m1 >>
rect 188 239 189 240 
<< m2 >>
rect 188 239 189 240 
<< m2c >>
rect 188 239 189 240 
<< m1 >>
rect 188 239 189 240 
<< m2 >>
rect 188 239 189 240 
<< m1 >>
rect 190 239 191 240 
<< m2 >>
rect 190 239 191 240 
<< m2c >>
rect 190 239 191 240 
<< m1 >>
rect 190 239 191 240 
<< m2 >>
rect 190 239 191 240 
<< m1 >>
rect 192 239 193 240 
<< m2 >>
rect 192 239 193 240 
<< m2c >>
rect 192 239 193 240 
<< m1 >>
rect 192 239 193 240 
<< m2 >>
rect 192 239 193 240 
<< m1 >>
rect 226 239 227 240 
<< m1 >>
rect 235 239 236 240 
<< m1 >>
rect 237 239 238 240 
<< m1 >>
rect 239 239 240 240 
<< m1 >>
rect 241 239 242 240 
<< m1 >>
rect 243 239 244 240 
<< m1 >>
rect 262 239 263 240 
<< m1 >>
rect 272 239 273 240 
<< m2 >>
rect 273 239 274 240 
<< m2 >>
rect 279 239 280 240 
<< m1 >>
rect 280 239 281 240 
<< m1 >>
rect 294 239 295 240 
<< m1 >>
rect 298 239 299 240 
<< m1 >>
rect 316 239 317 240 
<< m1 >>
rect 327 239 328 240 
<< m1 >>
rect 329 239 330 240 
<< m2 >>
rect 330 239 331 240 
<< m1 >>
rect 10 240 11 241 
<< m1 >>
rect 28 240 29 241 
<< m2 >>
rect 28 240 29 241 
<< m1 >>
rect 37 240 38 241 
<< m1 >>
rect 39 240 40 241 
<< m2 >>
rect 43 240 44 241 
<< m1 >>
rect 44 240 45 241 
<< m1 >>
rect 46 240 47 241 
<< m2 >>
rect 46 240 47 241 
<< m2 >>
rect 56 240 57 241 
<< m2 >>
rect 58 240 59 241 
<< m2 >>
rect 60 240 61 241 
<< m2 >>
rect 62 240 63 241 
<< m2 >>
rect 64 240 65 241 
<< m2 >>
rect 65 240 66 241 
<< m2 >>
rect 66 240 67 241 
<< m2 >>
rect 67 240 68 241 
<< m2 >>
rect 68 240 69 241 
<< m2 >>
rect 74 240 75 241 
<< m2 >>
rect 75 240 76 241 
<< m2 >>
rect 76 240 77 241 
<< m2 >>
rect 77 240 78 241 
<< m2 >>
rect 78 240 79 241 
<< m2 >>
rect 114 240 115 241 
<< m2 >>
rect 118 240 119 241 
<< m2 >>
rect 128 240 129 241 
<< m2 >>
rect 130 240 131 241 
<< m2 >>
rect 132 240 133 241 
<< m2 >>
rect 134 240 135 241 
<< m2 >>
rect 136 240 137 241 
<< m1 >>
rect 145 240 146 241 
<< m2 >>
rect 154 240 155 241 
<< m2 >>
rect 156 240 157 241 
<< m2 >>
rect 157 240 158 241 
<< m2 >>
rect 158 240 159 241 
<< m2 >>
rect 159 240 160 241 
<< m2 >>
rect 160 240 161 241 
<< m1 >>
rect 163 240 164 241 
<< m1 >>
rect 165 240 166 241 
<< m1 >>
rect 167 240 168 241 
<< m2 >>
rect 168 240 169 241 
<< m2 >>
rect 181 240 182 241 
<< m2 >>
rect 183 240 184 241 
<< m2 >>
rect 186 240 187 241 
<< m2 >>
rect 188 240 189 241 
<< m2 >>
rect 190 240 191 241 
<< m2 >>
rect 192 240 193 241 
<< m2 >>
rect 193 240 194 241 
<< m2 >>
rect 194 240 195 241 
<< m1 >>
rect 226 240 227 241 
<< m1 >>
rect 235 240 236 241 
<< m1 >>
rect 237 240 238 241 
<< m1 >>
rect 239 240 240 241 
<< m1 >>
rect 241 240 242 241 
<< m1 >>
rect 243 240 244 241 
<< m1 >>
rect 262 240 263 241 
<< m1 >>
rect 272 240 273 241 
<< m2 >>
rect 273 240 274 241 
<< m2 >>
rect 279 240 280 241 
<< m1 >>
rect 280 240 281 241 
<< m1 >>
rect 294 240 295 241 
<< m1 >>
rect 298 240 299 241 
<< m1 >>
rect 316 240 317 241 
<< m1 >>
rect 327 240 328 241 
<< m1 >>
rect 329 240 330 241 
<< m2 >>
rect 330 240 331 241 
<< m1 >>
rect 10 241 11 242 
<< m1 >>
rect 28 241 29 242 
<< m2 >>
rect 28 241 29 242 
<< m1 >>
rect 37 241 38 242 
<< m1 >>
rect 39 241 40 242 
<< m2 >>
rect 43 241 44 242 
<< m1 >>
rect 44 241 45 242 
<< m1 >>
rect 46 241 47 242 
<< m2 >>
rect 46 241 47 242 
<< m1 >>
rect 49 241 50 242 
<< m1 >>
rect 50 241 51 242 
<< m1 >>
rect 51 241 52 242 
<< m1 >>
rect 52 241 53 242 
<< m1 >>
rect 53 241 54 242 
<< m1 >>
rect 54 241 55 242 
<< m1 >>
rect 55 241 56 242 
<< m1 >>
rect 56 241 57 242 
<< m2 >>
rect 56 241 57 242 
<< m1 >>
rect 57 241 58 242 
<< m1 >>
rect 58 241 59 242 
<< m2 >>
rect 58 241 59 242 
<< m1 >>
rect 59 241 60 242 
<< m1 >>
rect 60 241 61 242 
<< m2 >>
rect 60 241 61 242 
<< m1 >>
rect 61 241 62 242 
<< m1 >>
rect 62 241 63 242 
<< m2 >>
rect 62 241 63 242 
<< m1 >>
rect 63 241 64 242 
<< m1 >>
rect 64 241 65 242 
<< m1 >>
rect 65 241 66 242 
<< m1 >>
rect 66 241 67 242 
<< m1 >>
rect 67 241 68 242 
<< m1 >>
rect 68 241 69 242 
<< m2 >>
rect 68 241 69 242 
<< m1 >>
rect 69 241 70 242 
<< m1 >>
rect 70 241 71 242 
<< m1 >>
rect 71 241 72 242 
<< m1 >>
rect 72 241 73 242 
<< m1 >>
rect 73 241 74 242 
<< m1 >>
rect 74 241 75 242 
<< m2 >>
rect 74 241 75 242 
<< m1 >>
rect 75 241 76 242 
<< m1 >>
rect 76 241 77 242 
<< m1 >>
rect 77 241 78 242 
<< m1 >>
rect 78 241 79 242 
<< m1 >>
rect 79 241 80 242 
<< m1 >>
rect 80 241 81 242 
<< m1 >>
rect 81 241 82 242 
<< m1 >>
rect 82 241 83 242 
<< m1 >>
rect 83 241 84 242 
<< m1 >>
rect 84 241 85 242 
<< m1 >>
rect 85 241 86 242 
<< m1 >>
rect 86 241 87 242 
<< m1 >>
rect 87 241 88 242 
<< m1 >>
rect 88 241 89 242 
<< m1 >>
rect 89 241 90 242 
<< m1 >>
rect 90 241 91 242 
<< m1 >>
rect 91 241 92 242 
<< m1 >>
rect 92 241 93 242 
<< m1 >>
rect 93 241 94 242 
<< m1 >>
rect 94 241 95 242 
<< m1 >>
rect 95 241 96 242 
<< m1 >>
rect 96 241 97 242 
<< m1 >>
rect 97 241 98 242 
<< m1 >>
rect 98 241 99 242 
<< m1 >>
rect 99 241 100 242 
<< m1 >>
rect 100 241 101 242 
<< m1 >>
rect 101 241 102 242 
<< m1 >>
rect 102 241 103 242 
<< m1 >>
rect 103 241 104 242 
<< m1 >>
rect 104 241 105 242 
<< m1 >>
rect 105 241 106 242 
<< m1 >>
rect 106 241 107 242 
<< m1 >>
rect 107 241 108 242 
<< m1 >>
rect 108 241 109 242 
<< m1 >>
rect 109 241 110 242 
<< m1 >>
rect 110 241 111 242 
<< m1 >>
rect 111 241 112 242 
<< m1 >>
rect 112 241 113 242 
<< m1 >>
rect 113 241 114 242 
<< m1 >>
rect 114 241 115 242 
<< m2 >>
rect 114 241 115 242 
<< m1 >>
rect 115 241 116 242 
<< m1 >>
rect 116 241 117 242 
<< m1 >>
rect 117 241 118 242 
<< m1 >>
rect 118 241 119 242 
<< m2 >>
rect 118 241 119 242 
<< m1 >>
rect 119 241 120 242 
<< m1 >>
rect 120 241 121 242 
<< m1 >>
rect 121 241 122 242 
<< m1 >>
rect 122 241 123 242 
<< m1 >>
rect 123 241 124 242 
<< m1 >>
rect 124 241 125 242 
<< m1 >>
rect 125 241 126 242 
<< m1 >>
rect 126 241 127 242 
<< m1 >>
rect 127 241 128 242 
<< m1 >>
rect 128 241 129 242 
<< m2 >>
rect 128 241 129 242 
<< m1 >>
rect 129 241 130 242 
<< m1 >>
rect 130 241 131 242 
<< m2 >>
rect 130 241 131 242 
<< m1 >>
rect 131 241 132 242 
<< m1 >>
rect 132 241 133 242 
<< m2 >>
rect 132 241 133 242 
<< m1 >>
rect 133 241 134 242 
<< m1 >>
rect 134 241 135 242 
<< m2 >>
rect 134 241 135 242 
<< m1 >>
rect 135 241 136 242 
<< m1 >>
rect 136 241 137 242 
<< m2 >>
rect 136 241 137 242 
<< m1 >>
rect 137 241 138 242 
<< m1 >>
rect 138 241 139 242 
<< m1 >>
rect 139 241 140 242 
<< m1 >>
rect 140 241 141 242 
<< m1 >>
rect 141 241 142 242 
<< m1 >>
rect 142 241 143 242 
<< m1 >>
rect 143 241 144 242 
<< m2 >>
rect 143 241 144 242 
<< m2c >>
rect 143 241 144 242 
<< m1 >>
rect 143 241 144 242 
<< m2 >>
rect 143 241 144 242 
<< m2 >>
rect 144 241 145 242 
<< m1 >>
rect 145 241 146 242 
<< m2 >>
rect 145 241 146 242 
<< m2 >>
rect 146 241 147 242 
<< m1 >>
rect 147 241 148 242 
<< m2 >>
rect 147 241 148 242 
<< m2c >>
rect 147 241 148 242 
<< m1 >>
rect 147 241 148 242 
<< m2 >>
rect 147 241 148 242 
<< m1 >>
rect 148 241 149 242 
<< m1 >>
rect 149 241 150 242 
<< m1 >>
rect 150 241 151 242 
<< m1 >>
rect 151 241 152 242 
<< m1 >>
rect 152 241 153 242 
<< m1 >>
rect 153 241 154 242 
<< m1 >>
rect 154 241 155 242 
<< m2 >>
rect 154 241 155 242 
<< m1 >>
rect 155 241 156 242 
<< m1 >>
rect 156 241 157 242 
<< m2 >>
rect 156 241 157 242 
<< m1 >>
rect 157 241 158 242 
<< m1 >>
rect 158 241 159 242 
<< m1 >>
rect 159 241 160 242 
<< m1 >>
rect 160 241 161 242 
<< m1 >>
rect 161 241 162 242 
<< m1 >>
rect 162 241 163 242 
<< m1 >>
rect 163 241 164 242 
<< m1 >>
rect 165 241 166 242 
<< m1 >>
rect 167 241 168 242 
<< m2 >>
rect 168 241 169 242 
<< m1 >>
rect 171 241 172 242 
<< m1 >>
rect 172 241 173 242 
<< m1 >>
rect 173 241 174 242 
<< m1 >>
rect 174 241 175 242 
<< m1 >>
rect 175 241 176 242 
<< m1 >>
rect 176 241 177 242 
<< m1 >>
rect 177 241 178 242 
<< m1 >>
rect 178 241 179 242 
<< m1 >>
rect 179 241 180 242 
<< m1 >>
rect 180 241 181 242 
<< m1 >>
rect 181 241 182 242 
<< m2 >>
rect 181 241 182 242 
<< m1 >>
rect 182 241 183 242 
<< m1 >>
rect 183 241 184 242 
<< m2 >>
rect 183 241 184 242 
<< m1 >>
rect 184 241 185 242 
<< m1 >>
rect 185 241 186 242 
<< m1 >>
rect 186 241 187 242 
<< m2 >>
rect 186 241 187 242 
<< m1 >>
rect 187 241 188 242 
<< m1 >>
rect 188 241 189 242 
<< m2 >>
rect 188 241 189 242 
<< m1 >>
rect 189 241 190 242 
<< m1 >>
rect 190 241 191 242 
<< m2 >>
rect 190 241 191 242 
<< m1 >>
rect 191 241 192 242 
<< m1 >>
rect 192 241 193 242 
<< m1 >>
rect 193 241 194 242 
<< m1 >>
rect 194 241 195 242 
<< m2 >>
rect 194 241 195 242 
<< m1 >>
rect 195 241 196 242 
<< m1 >>
rect 196 241 197 242 
<< m1 >>
rect 197 241 198 242 
<< m1 >>
rect 198 241 199 242 
<< m1 >>
rect 199 241 200 242 
<< m1 >>
rect 200 241 201 242 
<< m1 >>
rect 201 241 202 242 
<< m1 >>
rect 202 241 203 242 
<< m1 >>
rect 203 241 204 242 
<< m1 >>
rect 204 241 205 242 
<< m1 >>
rect 205 241 206 242 
<< m1 >>
rect 206 241 207 242 
<< m1 >>
rect 207 241 208 242 
<< m1 >>
rect 208 241 209 242 
<< m1 >>
rect 209 241 210 242 
<< m1 >>
rect 210 241 211 242 
<< m1 >>
rect 211 241 212 242 
<< m1 >>
rect 212 241 213 242 
<< m1 >>
rect 213 241 214 242 
<< m1 >>
rect 214 241 215 242 
<< m1 >>
rect 215 241 216 242 
<< m1 >>
rect 216 241 217 242 
<< m1 >>
rect 217 241 218 242 
<< m1 >>
rect 218 241 219 242 
<< m1 >>
rect 219 241 220 242 
<< m1 >>
rect 220 241 221 242 
<< m1 >>
rect 221 241 222 242 
<< m1 >>
rect 222 241 223 242 
<< m1 >>
rect 223 241 224 242 
<< m1 >>
rect 224 241 225 242 
<< m2 >>
rect 224 241 225 242 
<< m2c >>
rect 224 241 225 242 
<< m1 >>
rect 224 241 225 242 
<< m2 >>
rect 224 241 225 242 
<< m2 >>
rect 225 241 226 242 
<< m1 >>
rect 226 241 227 242 
<< m2 >>
rect 226 241 227 242 
<< m2 >>
rect 227 241 228 242 
<< m1 >>
rect 228 241 229 242 
<< m2 >>
rect 228 241 229 242 
<< m2c >>
rect 228 241 229 242 
<< m1 >>
rect 228 241 229 242 
<< m2 >>
rect 228 241 229 242 
<< m1 >>
rect 229 241 230 242 
<< m1 >>
rect 230 241 231 242 
<< m1 >>
rect 231 241 232 242 
<< m1 >>
rect 232 241 233 242 
<< m1 >>
rect 233 241 234 242 
<< m2 >>
rect 233 241 234 242 
<< m2c >>
rect 233 241 234 242 
<< m1 >>
rect 233 241 234 242 
<< m2 >>
rect 233 241 234 242 
<< m2 >>
rect 234 241 235 242 
<< m1 >>
rect 235 241 236 242 
<< m2 >>
rect 235 241 236 242 
<< m2 >>
rect 236 241 237 242 
<< m1 >>
rect 237 241 238 242 
<< m2 >>
rect 237 241 238 242 
<< m2 >>
rect 238 241 239 242 
<< m1 >>
rect 239 241 240 242 
<< m2 >>
rect 239 241 240 242 
<< m2 >>
rect 240 241 241 242 
<< m1 >>
rect 241 241 242 242 
<< m2 >>
rect 241 241 242 242 
<< m2c >>
rect 241 241 242 242 
<< m1 >>
rect 241 241 242 242 
<< m2 >>
rect 241 241 242 242 
<< m1 >>
rect 243 241 244 242 
<< m1 >>
rect 262 241 263 242 
<< m1 >>
rect 272 241 273 242 
<< m2 >>
rect 273 241 274 242 
<< m2 >>
rect 279 241 280 242 
<< m1 >>
rect 280 241 281 242 
<< m1 >>
rect 294 241 295 242 
<< m1 >>
rect 298 241 299 242 
<< m1 >>
rect 316 241 317 242 
<< m1 >>
rect 317 241 318 242 
<< m1 >>
rect 318 241 319 242 
<< m1 >>
rect 319 241 320 242 
<< m1 >>
rect 320 241 321 242 
<< m1 >>
rect 321 241 322 242 
<< m1 >>
rect 322 241 323 242 
<< m1 >>
rect 327 241 328 242 
<< m1 >>
rect 329 241 330 242 
<< m2 >>
rect 330 241 331 242 
<< m1 >>
rect 10 242 11 243 
<< m1 >>
rect 28 242 29 243 
<< m2 >>
rect 28 242 29 243 
<< m1 >>
rect 37 242 38 243 
<< m1 >>
rect 39 242 40 243 
<< m2 >>
rect 43 242 44 243 
<< m1 >>
rect 44 242 45 243 
<< m1 >>
rect 46 242 47 243 
<< m2 >>
rect 46 242 47 243 
<< m1 >>
rect 49 242 50 243 
<< m2 >>
rect 56 242 57 243 
<< m2 >>
rect 58 242 59 243 
<< m2 >>
rect 60 242 61 243 
<< m2 >>
rect 62 242 63 243 
<< m2 >>
rect 63 242 64 243 
<< m2 >>
rect 64 242 65 243 
<< m2 >>
rect 68 242 69 243 
<< m2 >>
rect 74 242 75 243 
<< m2 >>
rect 114 242 115 243 
<< m2 >>
rect 115 242 116 243 
<< m2 >>
rect 116 242 117 243 
<< m2 >>
rect 118 242 119 243 
<< m2 >>
rect 128 242 129 243 
<< m2 >>
rect 130 242 131 243 
<< m2 >>
rect 132 242 133 243 
<< m2 >>
rect 134 242 135 243 
<< m2 >>
rect 136 242 137 243 
<< m1 >>
rect 145 242 146 243 
<< m2 >>
rect 154 242 155 243 
<< m2 >>
rect 156 242 157 243 
<< m1 >>
rect 165 242 166 243 
<< m1 >>
rect 167 242 168 243 
<< m2 >>
rect 168 242 169 243 
<< m1 >>
rect 171 242 172 243 
<< m2 >>
rect 181 242 182 243 
<< m2 >>
rect 183 242 184 243 
<< m2 >>
rect 186 242 187 243 
<< m2 >>
rect 188 242 189 243 
<< m2 >>
rect 190 242 191 243 
<< m2 >>
rect 194 242 195 243 
<< m1 >>
rect 226 242 227 243 
<< m1 >>
rect 235 242 236 243 
<< m1 >>
rect 237 242 238 243 
<< m1 >>
rect 239 242 240 243 
<< m1 >>
rect 243 242 244 243 
<< m1 >>
rect 262 242 263 243 
<< m1 >>
rect 272 242 273 243 
<< m2 >>
rect 273 242 274 243 
<< m2 >>
rect 279 242 280 243 
<< m1 >>
rect 280 242 281 243 
<< m1 >>
rect 294 242 295 243 
<< m1 >>
rect 298 242 299 243 
<< m1 >>
rect 322 242 323 243 
<< m1 >>
rect 327 242 328 243 
<< m1 >>
rect 329 242 330 243 
<< m2 >>
rect 330 242 331 243 
<< m1 >>
rect 10 243 11 244 
<< m1 >>
rect 28 243 29 244 
<< m2 >>
rect 28 243 29 244 
<< m1 >>
rect 37 243 38 244 
<< m1 >>
rect 39 243 40 244 
<< m2 >>
rect 43 243 44 244 
<< m1 >>
rect 44 243 45 244 
<< m1 >>
rect 46 243 47 244 
<< m2 >>
rect 46 243 47 244 
<< m1 >>
rect 49 243 50 244 
<< m1 >>
rect 56 243 57 244 
<< m2 >>
rect 56 243 57 244 
<< m2c >>
rect 56 243 57 244 
<< m1 >>
rect 56 243 57 244 
<< m2 >>
rect 56 243 57 244 
<< m1 >>
rect 58 243 59 244 
<< m2 >>
rect 58 243 59 244 
<< m2c >>
rect 58 243 59 244 
<< m1 >>
rect 58 243 59 244 
<< m2 >>
rect 58 243 59 244 
<< m1 >>
rect 60 243 61 244 
<< m2 >>
rect 60 243 61 244 
<< m2c >>
rect 60 243 61 244 
<< m1 >>
rect 60 243 61 244 
<< m2 >>
rect 60 243 61 244 
<< m1 >>
rect 64 243 65 244 
<< m2 >>
rect 64 243 65 244 
<< m2c >>
rect 64 243 65 244 
<< m1 >>
rect 64 243 65 244 
<< m2 >>
rect 64 243 65 244 
<< m1 >>
rect 68 243 69 244 
<< m2 >>
rect 68 243 69 244 
<< m2c >>
rect 68 243 69 244 
<< m1 >>
rect 68 243 69 244 
<< m2 >>
rect 68 243 69 244 
<< m1 >>
rect 69 243 70 244 
<< m1 >>
rect 70 243 71 244 
<< m1 >>
rect 71 243 72 244 
<< m1 >>
rect 72 243 73 244 
<< m1 >>
rect 73 243 74 244 
<< m2 >>
rect 74 243 75 244 
<< m1 >>
rect 85 243 86 244 
<< m1 >>
rect 86 243 87 244 
<< m1 >>
rect 87 243 88 244 
<< m1 >>
rect 88 243 89 244 
<< m1 >>
rect 89 243 90 244 
<< m1 >>
rect 90 243 91 244 
<< m1 >>
rect 91 243 92 244 
<< m1 >>
rect 92 243 93 244 
<< m1 >>
rect 93 243 94 244 
<< m1 >>
rect 94 243 95 244 
<< m1 >>
rect 95 243 96 244 
<< m1 >>
rect 96 243 97 244 
<< m1 >>
rect 97 243 98 244 
<< m1 >>
rect 98 243 99 244 
<< m1 >>
rect 99 243 100 244 
<< m1 >>
rect 100 243 101 244 
<< m1 >>
rect 116 243 117 244 
<< m2 >>
rect 116 243 117 244 
<< m2c >>
rect 116 243 117 244 
<< m1 >>
rect 116 243 117 244 
<< m2 >>
rect 116 243 117 244 
<< m1 >>
rect 118 243 119 244 
<< m2 >>
rect 118 243 119 244 
<< m2c >>
rect 118 243 119 244 
<< m1 >>
rect 118 243 119 244 
<< m2 >>
rect 118 243 119 244 
<< m1 >>
rect 128 243 129 244 
<< m2 >>
rect 128 243 129 244 
<< m2c >>
rect 128 243 129 244 
<< m1 >>
rect 128 243 129 244 
<< m2 >>
rect 128 243 129 244 
<< m1 >>
rect 130 243 131 244 
<< m2 >>
rect 130 243 131 244 
<< m2c >>
rect 130 243 131 244 
<< m1 >>
rect 130 243 131 244 
<< m2 >>
rect 130 243 131 244 
<< m1 >>
rect 132 243 133 244 
<< m2 >>
rect 132 243 133 244 
<< m2c >>
rect 132 243 133 244 
<< m1 >>
rect 132 243 133 244 
<< m2 >>
rect 132 243 133 244 
<< m1 >>
rect 134 243 135 244 
<< m2 >>
rect 134 243 135 244 
<< m2c >>
rect 134 243 135 244 
<< m1 >>
rect 134 243 135 244 
<< m2 >>
rect 134 243 135 244 
<< m1 >>
rect 136 243 137 244 
<< m2 >>
rect 136 243 137 244 
<< m2c >>
rect 136 243 137 244 
<< m1 >>
rect 136 243 137 244 
<< m2 >>
rect 136 243 137 244 
<< m1 >>
rect 139 243 140 244 
<< m1 >>
rect 140 243 141 244 
<< m1 >>
rect 141 243 142 244 
<< m1 >>
rect 142 243 143 244 
<< m1 >>
rect 143 243 144 244 
<< m2 >>
rect 143 243 144 244 
<< m2c >>
rect 143 243 144 244 
<< m1 >>
rect 143 243 144 244 
<< m2 >>
rect 143 243 144 244 
<< m2 >>
rect 144 243 145 244 
<< m1 >>
rect 145 243 146 244 
<< m2 >>
rect 145 243 146 244 
<< m1 >>
rect 154 243 155 244 
<< m2 >>
rect 154 243 155 244 
<< m1 >>
rect 155 243 156 244 
<< m1 >>
rect 156 243 157 244 
<< m2 >>
rect 156 243 157 244 
<< m2c >>
rect 156 243 157 244 
<< m1 >>
rect 156 243 157 244 
<< m2 >>
rect 156 243 157 244 
<< m1 >>
rect 163 243 164 244 
<< m2 >>
rect 163 243 164 244 
<< m2c >>
rect 163 243 164 244 
<< m1 >>
rect 163 243 164 244 
<< m2 >>
rect 163 243 164 244 
<< m2 >>
rect 164 243 165 244 
<< m1 >>
rect 165 243 166 244 
<< m2 >>
rect 165 243 166 244 
<< m2 >>
rect 166 243 167 244 
<< m1 >>
rect 167 243 168 244 
<< m2 >>
rect 167 243 168 244 
<< m2 >>
rect 168 243 169 244 
<< m1 >>
rect 171 243 172 244 
<< m1 >>
rect 181 243 182 244 
<< m2 >>
rect 181 243 182 244 
<< m2c >>
rect 181 243 182 244 
<< m1 >>
rect 181 243 182 244 
<< m2 >>
rect 181 243 182 244 
<< m1 >>
rect 183 243 184 244 
<< m2 >>
rect 183 243 184 244 
<< m2c >>
rect 183 243 184 244 
<< m1 >>
rect 183 243 184 244 
<< m2 >>
rect 183 243 184 244 
<< m1 >>
rect 186 243 187 244 
<< m2 >>
rect 186 243 187 244 
<< m2c >>
rect 186 243 187 244 
<< m1 >>
rect 186 243 187 244 
<< m2 >>
rect 186 243 187 244 
<< m1 >>
rect 188 243 189 244 
<< m2 >>
rect 188 243 189 244 
<< m2c >>
rect 188 243 189 244 
<< m1 >>
rect 188 243 189 244 
<< m2 >>
rect 188 243 189 244 
<< m1 >>
rect 190 243 191 244 
<< m2 >>
rect 190 243 191 244 
<< m2c >>
rect 190 243 191 244 
<< m1 >>
rect 190 243 191 244 
<< m2 >>
rect 190 243 191 244 
<< m1 >>
rect 194 243 195 244 
<< m2 >>
rect 194 243 195 244 
<< m2c >>
rect 194 243 195 244 
<< m1 >>
rect 194 243 195 244 
<< m2 >>
rect 194 243 195 244 
<< m1 >>
rect 195 243 196 244 
<< m1 >>
rect 196 243 197 244 
<< m1 >>
rect 197 243 198 244 
<< m1 >>
rect 198 243 199 244 
<< m1 >>
rect 199 243 200 244 
<< m1 >>
rect 226 243 227 244 
<< m1 >>
rect 235 243 236 244 
<< m1 >>
rect 237 243 238 244 
<< m1 >>
rect 239 243 240 244 
<< m1 >>
rect 243 243 244 244 
<< m1 >>
rect 262 243 263 244 
<< m1 >>
rect 272 243 273 244 
<< m2 >>
rect 273 243 274 244 
<< m2 >>
rect 279 243 280 244 
<< m1 >>
rect 280 243 281 244 
<< m1 >>
rect 294 243 295 244 
<< m1 >>
rect 298 243 299 244 
<< m1 >>
rect 322 243 323 244 
<< m1 >>
rect 327 243 328 244 
<< m1 >>
rect 329 243 330 244 
<< m2 >>
rect 330 243 331 244 
<< m1 >>
rect 10 244 11 245 
<< m1 >>
rect 28 244 29 245 
<< m2 >>
rect 28 244 29 245 
<< m1 >>
rect 34 244 35 245 
<< m1 >>
rect 35 244 36 245 
<< m2 >>
rect 35 244 36 245 
<< m2c >>
rect 35 244 36 245 
<< m1 >>
rect 35 244 36 245 
<< m2 >>
rect 35 244 36 245 
<< m2 >>
rect 36 244 37 245 
<< m1 >>
rect 37 244 38 245 
<< m2 >>
rect 37 244 38 245 
<< m1 >>
rect 39 244 40 245 
<< m2 >>
rect 43 244 44 245 
<< m1 >>
rect 44 244 45 245 
<< m1 >>
rect 46 244 47 245 
<< m2 >>
rect 46 244 47 245 
<< m1 >>
rect 49 244 50 245 
<< m1 >>
rect 56 244 57 245 
<< m1 >>
rect 58 244 59 245 
<< m1 >>
rect 60 244 61 245 
<< m1 >>
rect 64 244 65 245 
<< m1 >>
rect 73 244 74 245 
<< m2 >>
rect 74 244 75 245 
<< m1 >>
rect 85 244 86 245 
<< m1 >>
rect 100 244 101 245 
<< m1 >>
rect 116 244 117 245 
<< m1 >>
rect 118 244 119 245 
<< m1 >>
rect 128 244 129 245 
<< m1 >>
rect 130 244 131 245 
<< m1 >>
rect 132 244 133 245 
<< m1 >>
rect 134 244 135 245 
<< m1 >>
rect 136 244 137 245 
<< m1 >>
rect 139 244 140 245 
<< m1 >>
rect 145 244 146 245 
<< m2 >>
rect 145 244 146 245 
<< m1 >>
rect 154 244 155 245 
<< m2 >>
rect 154 244 155 245 
<< m1 >>
rect 163 244 164 245 
<< m1 >>
rect 165 244 166 245 
<< m1 >>
rect 167 244 168 245 
<< m1 >>
rect 171 244 172 245 
<< m1 >>
rect 181 244 182 245 
<< m1 >>
rect 183 244 184 245 
<< m1 >>
rect 186 244 187 245 
<< m1 >>
rect 188 244 189 245 
<< m1 >>
rect 190 244 191 245 
<< m1 >>
rect 199 244 200 245 
<< m1 >>
rect 226 244 227 245 
<< m1 >>
rect 235 244 236 245 
<< m1 >>
rect 237 244 238 245 
<< m1 >>
rect 239 244 240 245 
<< m1 >>
rect 243 244 244 245 
<< m1 >>
rect 262 244 263 245 
<< m1 >>
rect 272 244 273 245 
<< m2 >>
rect 273 244 274 245 
<< m2 >>
rect 279 244 280 245 
<< m1 >>
rect 280 244 281 245 
<< m1 >>
rect 294 244 295 245 
<< m1 >>
rect 298 244 299 245 
<< m1 >>
rect 322 244 323 245 
<< m1 >>
rect 327 244 328 245 
<< m1 >>
rect 329 244 330 245 
<< m2 >>
rect 330 244 331 245 
<< m1 >>
rect 10 245 11 246 
<< m1 >>
rect 28 245 29 246 
<< m2 >>
rect 28 245 29 246 
<< m1 >>
rect 34 245 35 246 
<< m1 >>
rect 37 245 38 246 
<< m2 >>
rect 37 245 38 246 
<< m1 >>
rect 39 245 40 246 
<< m2 >>
rect 43 245 44 246 
<< m1 >>
rect 44 245 45 246 
<< m1 >>
rect 46 245 47 246 
<< m2 >>
rect 46 245 47 246 
<< m1 >>
rect 49 245 50 246 
<< m1 >>
rect 56 245 57 246 
<< m1 >>
rect 58 245 59 246 
<< m1 >>
rect 60 245 61 246 
<< m1 >>
rect 64 245 65 246 
<< m1 >>
rect 73 245 74 246 
<< m2 >>
rect 74 245 75 246 
<< m1 >>
rect 85 245 86 246 
<< m1 >>
rect 100 245 101 246 
<< m1 >>
rect 116 245 117 246 
<< m1 >>
rect 118 245 119 246 
<< m1 >>
rect 128 245 129 246 
<< m1 >>
rect 130 245 131 246 
<< m1 >>
rect 132 245 133 246 
<< m1 >>
rect 134 245 135 246 
<< m1 >>
rect 136 245 137 246 
<< m1 >>
rect 139 245 140 246 
<< m1 >>
rect 145 245 146 246 
<< m2 >>
rect 145 245 146 246 
<< m1 >>
rect 154 245 155 246 
<< m2 >>
rect 154 245 155 246 
<< m1 >>
rect 163 245 164 246 
<< m1 >>
rect 165 245 166 246 
<< m1 >>
rect 167 245 168 246 
<< m1 >>
rect 171 245 172 246 
<< m1 >>
rect 181 245 182 246 
<< m1 >>
rect 183 245 184 246 
<< m1 >>
rect 186 245 187 246 
<< m1 >>
rect 188 245 189 246 
<< m1 >>
rect 190 245 191 246 
<< m1 >>
rect 199 245 200 246 
<< m1 >>
rect 226 245 227 246 
<< m1 >>
rect 235 245 236 246 
<< m1 >>
rect 237 245 238 246 
<< m1 >>
rect 239 245 240 246 
<< m1 >>
rect 243 245 244 246 
<< m1 >>
rect 262 245 263 246 
<< m1 >>
rect 272 245 273 246 
<< m2 >>
rect 273 245 274 246 
<< m2 >>
rect 279 245 280 246 
<< m1 >>
rect 280 245 281 246 
<< m1 >>
rect 294 245 295 246 
<< m1 >>
rect 298 245 299 246 
<< m1 >>
rect 322 245 323 246 
<< m1 >>
rect 327 245 328 246 
<< m1 >>
rect 329 245 330 246 
<< m2 >>
rect 330 245 331 246 
<< m1 >>
rect 10 246 11 247 
<< pdiffusion >>
rect 12 246 13 247 
<< pdiffusion >>
rect 13 246 14 247 
<< pdiffusion >>
rect 14 246 15 247 
<< pdiffusion >>
rect 15 246 16 247 
<< pdiffusion >>
rect 16 246 17 247 
<< pdiffusion >>
rect 17 246 18 247 
<< m1 >>
rect 28 246 29 247 
<< m2 >>
rect 28 246 29 247 
<< pdiffusion >>
rect 30 246 31 247 
<< pdiffusion >>
rect 31 246 32 247 
<< pdiffusion >>
rect 32 246 33 247 
<< pdiffusion >>
rect 33 246 34 247 
<< m1 >>
rect 34 246 35 247 
<< pdiffusion >>
rect 34 246 35 247 
<< pdiffusion >>
rect 35 246 36 247 
<< m1 >>
rect 37 246 38 247 
<< m2 >>
rect 37 246 38 247 
<< m1 >>
rect 39 246 40 247 
<< m2 >>
rect 43 246 44 247 
<< m1 >>
rect 44 246 45 247 
<< m1 >>
rect 46 246 47 247 
<< m2 >>
rect 46 246 47 247 
<< pdiffusion >>
rect 48 246 49 247 
<< m1 >>
rect 49 246 50 247 
<< pdiffusion >>
rect 49 246 50 247 
<< pdiffusion >>
rect 50 246 51 247 
<< pdiffusion >>
rect 51 246 52 247 
<< pdiffusion >>
rect 52 246 53 247 
<< pdiffusion >>
rect 53 246 54 247 
<< m1 >>
rect 56 246 57 247 
<< m1 >>
rect 58 246 59 247 
<< m1 >>
rect 60 246 61 247 
<< m1 >>
rect 64 246 65 247 
<< pdiffusion >>
rect 66 246 67 247 
<< pdiffusion >>
rect 67 246 68 247 
<< pdiffusion >>
rect 68 246 69 247 
<< pdiffusion >>
rect 69 246 70 247 
<< pdiffusion >>
rect 70 246 71 247 
<< pdiffusion >>
rect 71 246 72 247 
<< m1 >>
rect 73 246 74 247 
<< m2 >>
rect 74 246 75 247 
<< pdiffusion >>
rect 84 246 85 247 
<< m1 >>
rect 85 246 86 247 
<< pdiffusion >>
rect 85 246 86 247 
<< pdiffusion >>
rect 86 246 87 247 
<< pdiffusion >>
rect 87 246 88 247 
<< pdiffusion >>
rect 88 246 89 247 
<< pdiffusion >>
rect 89 246 90 247 
<< m1 >>
rect 100 246 101 247 
<< pdiffusion >>
rect 102 246 103 247 
<< pdiffusion >>
rect 103 246 104 247 
<< pdiffusion >>
rect 104 246 105 247 
<< pdiffusion >>
rect 105 246 106 247 
<< pdiffusion >>
rect 106 246 107 247 
<< pdiffusion >>
rect 107 246 108 247 
<< m1 >>
rect 116 246 117 247 
<< m1 >>
rect 118 246 119 247 
<< pdiffusion >>
rect 120 246 121 247 
<< pdiffusion >>
rect 121 246 122 247 
<< pdiffusion >>
rect 122 246 123 247 
<< pdiffusion >>
rect 123 246 124 247 
<< pdiffusion >>
rect 124 246 125 247 
<< pdiffusion >>
rect 125 246 126 247 
<< m1 >>
rect 128 246 129 247 
<< m1 >>
rect 130 246 131 247 
<< m1 >>
rect 132 246 133 247 
<< m1 >>
rect 134 246 135 247 
<< m1 >>
rect 136 246 137 247 
<< pdiffusion >>
rect 138 246 139 247 
<< m1 >>
rect 139 246 140 247 
<< pdiffusion >>
rect 139 246 140 247 
<< pdiffusion >>
rect 140 246 141 247 
<< pdiffusion >>
rect 141 246 142 247 
<< pdiffusion >>
rect 142 246 143 247 
<< pdiffusion >>
rect 143 246 144 247 
<< m1 >>
rect 145 246 146 247 
<< m2 >>
rect 145 246 146 247 
<< m1 >>
rect 154 246 155 247 
<< m2 >>
rect 154 246 155 247 
<< pdiffusion >>
rect 156 246 157 247 
<< pdiffusion >>
rect 157 246 158 247 
<< pdiffusion >>
rect 158 246 159 247 
<< pdiffusion >>
rect 159 246 160 247 
<< pdiffusion >>
rect 160 246 161 247 
<< pdiffusion >>
rect 161 246 162 247 
<< m1 >>
rect 163 246 164 247 
<< m1 >>
rect 165 246 166 247 
<< m1 >>
rect 167 246 168 247 
<< m1 >>
rect 171 246 172 247 
<< pdiffusion >>
rect 174 246 175 247 
<< pdiffusion >>
rect 175 246 176 247 
<< pdiffusion >>
rect 176 246 177 247 
<< pdiffusion >>
rect 177 246 178 247 
<< pdiffusion >>
rect 178 246 179 247 
<< pdiffusion >>
rect 179 246 180 247 
<< m1 >>
rect 181 246 182 247 
<< m1 >>
rect 183 246 184 247 
<< m1 >>
rect 186 246 187 247 
<< m1 >>
rect 188 246 189 247 
<< m1 >>
rect 190 246 191 247 
<< pdiffusion >>
rect 192 246 193 247 
<< pdiffusion >>
rect 193 246 194 247 
<< pdiffusion >>
rect 194 246 195 247 
<< pdiffusion >>
rect 195 246 196 247 
<< pdiffusion >>
rect 196 246 197 247 
<< pdiffusion >>
rect 197 246 198 247 
<< m1 >>
rect 199 246 200 247 
<< pdiffusion >>
rect 210 246 211 247 
<< pdiffusion >>
rect 211 246 212 247 
<< pdiffusion >>
rect 212 246 213 247 
<< pdiffusion >>
rect 213 246 214 247 
<< pdiffusion >>
rect 214 246 215 247 
<< pdiffusion >>
rect 215 246 216 247 
<< m1 >>
rect 226 246 227 247 
<< pdiffusion >>
rect 228 246 229 247 
<< pdiffusion >>
rect 229 246 230 247 
<< pdiffusion >>
rect 230 246 231 247 
<< pdiffusion >>
rect 231 246 232 247 
<< pdiffusion >>
rect 232 246 233 247 
<< pdiffusion >>
rect 233 246 234 247 
<< m1 >>
rect 235 246 236 247 
<< m1 >>
rect 237 246 238 247 
<< m1 >>
rect 239 246 240 247 
<< m1 >>
rect 243 246 244 247 
<< pdiffusion >>
rect 246 246 247 247 
<< pdiffusion >>
rect 247 246 248 247 
<< pdiffusion >>
rect 248 246 249 247 
<< pdiffusion >>
rect 249 246 250 247 
<< pdiffusion >>
rect 250 246 251 247 
<< pdiffusion >>
rect 251 246 252 247 
<< m1 >>
rect 262 246 263 247 
<< pdiffusion >>
rect 264 246 265 247 
<< pdiffusion >>
rect 265 246 266 247 
<< pdiffusion >>
rect 266 246 267 247 
<< pdiffusion >>
rect 267 246 268 247 
<< pdiffusion >>
rect 268 246 269 247 
<< pdiffusion >>
rect 269 246 270 247 
<< m1 >>
rect 272 246 273 247 
<< m2 >>
rect 273 246 274 247 
<< m2 >>
rect 279 246 280 247 
<< m1 >>
rect 280 246 281 247 
<< pdiffusion >>
rect 282 246 283 247 
<< pdiffusion >>
rect 283 246 284 247 
<< pdiffusion >>
rect 284 246 285 247 
<< pdiffusion >>
rect 285 246 286 247 
<< pdiffusion >>
rect 286 246 287 247 
<< pdiffusion >>
rect 287 246 288 247 
<< m1 >>
rect 294 246 295 247 
<< m1 >>
rect 298 246 299 247 
<< pdiffusion >>
rect 300 246 301 247 
<< pdiffusion >>
rect 301 246 302 247 
<< pdiffusion >>
rect 302 246 303 247 
<< pdiffusion >>
rect 303 246 304 247 
<< pdiffusion >>
rect 304 246 305 247 
<< pdiffusion >>
rect 305 246 306 247 
<< pdiffusion >>
rect 318 246 319 247 
<< pdiffusion >>
rect 319 246 320 247 
<< pdiffusion >>
rect 320 246 321 247 
<< pdiffusion >>
rect 321 246 322 247 
<< m1 >>
rect 322 246 323 247 
<< pdiffusion >>
rect 322 246 323 247 
<< pdiffusion >>
rect 323 246 324 247 
<< m1 >>
rect 327 246 328 247 
<< m1 >>
rect 329 246 330 247 
<< m2 >>
rect 330 246 331 247 
<< pdiffusion >>
rect 336 246 337 247 
<< pdiffusion >>
rect 337 246 338 247 
<< pdiffusion >>
rect 338 246 339 247 
<< pdiffusion >>
rect 339 246 340 247 
<< pdiffusion >>
rect 340 246 341 247 
<< pdiffusion >>
rect 341 246 342 247 
<< m1 >>
rect 10 247 11 248 
<< pdiffusion >>
rect 12 247 13 248 
<< pdiffusion >>
rect 13 247 14 248 
<< pdiffusion >>
rect 14 247 15 248 
<< pdiffusion >>
rect 15 247 16 248 
<< pdiffusion >>
rect 16 247 17 248 
<< pdiffusion >>
rect 17 247 18 248 
<< m1 >>
rect 28 247 29 248 
<< m2 >>
rect 28 247 29 248 
<< pdiffusion >>
rect 30 247 31 248 
<< pdiffusion >>
rect 31 247 32 248 
<< pdiffusion >>
rect 32 247 33 248 
<< pdiffusion >>
rect 33 247 34 248 
<< pdiffusion >>
rect 34 247 35 248 
<< pdiffusion >>
rect 35 247 36 248 
<< m1 >>
rect 37 247 38 248 
<< m2 >>
rect 37 247 38 248 
<< m1 >>
rect 39 247 40 248 
<< m2 >>
rect 43 247 44 248 
<< m1 >>
rect 44 247 45 248 
<< m1 >>
rect 46 247 47 248 
<< m2 >>
rect 46 247 47 248 
<< pdiffusion >>
rect 48 247 49 248 
<< pdiffusion >>
rect 49 247 50 248 
<< pdiffusion >>
rect 50 247 51 248 
<< pdiffusion >>
rect 51 247 52 248 
<< pdiffusion >>
rect 52 247 53 248 
<< pdiffusion >>
rect 53 247 54 248 
<< m1 >>
rect 56 247 57 248 
<< m1 >>
rect 58 247 59 248 
<< m1 >>
rect 60 247 61 248 
<< m1 >>
rect 64 247 65 248 
<< pdiffusion >>
rect 66 247 67 248 
<< pdiffusion >>
rect 67 247 68 248 
<< pdiffusion >>
rect 68 247 69 248 
<< pdiffusion >>
rect 69 247 70 248 
<< pdiffusion >>
rect 70 247 71 248 
<< pdiffusion >>
rect 71 247 72 248 
<< m1 >>
rect 73 247 74 248 
<< m2 >>
rect 74 247 75 248 
<< pdiffusion >>
rect 84 247 85 248 
<< pdiffusion >>
rect 85 247 86 248 
<< pdiffusion >>
rect 86 247 87 248 
<< pdiffusion >>
rect 87 247 88 248 
<< pdiffusion >>
rect 88 247 89 248 
<< pdiffusion >>
rect 89 247 90 248 
<< m1 >>
rect 100 247 101 248 
<< pdiffusion >>
rect 102 247 103 248 
<< pdiffusion >>
rect 103 247 104 248 
<< pdiffusion >>
rect 104 247 105 248 
<< pdiffusion >>
rect 105 247 106 248 
<< pdiffusion >>
rect 106 247 107 248 
<< pdiffusion >>
rect 107 247 108 248 
<< m1 >>
rect 116 247 117 248 
<< m1 >>
rect 118 247 119 248 
<< pdiffusion >>
rect 120 247 121 248 
<< pdiffusion >>
rect 121 247 122 248 
<< pdiffusion >>
rect 122 247 123 248 
<< pdiffusion >>
rect 123 247 124 248 
<< pdiffusion >>
rect 124 247 125 248 
<< pdiffusion >>
rect 125 247 126 248 
<< m1 >>
rect 128 247 129 248 
<< m1 >>
rect 130 247 131 248 
<< m1 >>
rect 132 247 133 248 
<< m1 >>
rect 134 247 135 248 
<< m1 >>
rect 136 247 137 248 
<< pdiffusion >>
rect 138 247 139 248 
<< pdiffusion >>
rect 139 247 140 248 
<< pdiffusion >>
rect 140 247 141 248 
<< pdiffusion >>
rect 141 247 142 248 
<< pdiffusion >>
rect 142 247 143 248 
<< pdiffusion >>
rect 143 247 144 248 
<< m1 >>
rect 145 247 146 248 
<< m2 >>
rect 145 247 146 248 
<< m1 >>
rect 154 247 155 248 
<< m2 >>
rect 154 247 155 248 
<< pdiffusion >>
rect 156 247 157 248 
<< pdiffusion >>
rect 157 247 158 248 
<< pdiffusion >>
rect 158 247 159 248 
<< pdiffusion >>
rect 159 247 160 248 
<< pdiffusion >>
rect 160 247 161 248 
<< pdiffusion >>
rect 161 247 162 248 
<< m1 >>
rect 163 247 164 248 
<< m1 >>
rect 165 247 166 248 
<< m1 >>
rect 167 247 168 248 
<< m1 >>
rect 171 247 172 248 
<< pdiffusion >>
rect 174 247 175 248 
<< pdiffusion >>
rect 175 247 176 248 
<< pdiffusion >>
rect 176 247 177 248 
<< pdiffusion >>
rect 177 247 178 248 
<< pdiffusion >>
rect 178 247 179 248 
<< pdiffusion >>
rect 179 247 180 248 
<< m1 >>
rect 181 247 182 248 
<< m1 >>
rect 183 247 184 248 
<< m1 >>
rect 186 247 187 248 
<< m1 >>
rect 188 247 189 248 
<< m1 >>
rect 190 247 191 248 
<< pdiffusion >>
rect 192 247 193 248 
<< pdiffusion >>
rect 193 247 194 248 
<< pdiffusion >>
rect 194 247 195 248 
<< pdiffusion >>
rect 195 247 196 248 
<< pdiffusion >>
rect 196 247 197 248 
<< pdiffusion >>
rect 197 247 198 248 
<< m1 >>
rect 199 247 200 248 
<< pdiffusion >>
rect 210 247 211 248 
<< pdiffusion >>
rect 211 247 212 248 
<< pdiffusion >>
rect 212 247 213 248 
<< pdiffusion >>
rect 213 247 214 248 
<< pdiffusion >>
rect 214 247 215 248 
<< pdiffusion >>
rect 215 247 216 248 
<< m1 >>
rect 226 247 227 248 
<< pdiffusion >>
rect 228 247 229 248 
<< pdiffusion >>
rect 229 247 230 248 
<< pdiffusion >>
rect 230 247 231 248 
<< pdiffusion >>
rect 231 247 232 248 
<< pdiffusion >>
rect 232 247 233 248 
<< pdiffusion >>
rect 233 247 234 248 
<< m1 >>
rect 235 247 236 248 
<< m1 >>
rect 237 247 238 248 
<< m1 >>
rect 239 247 240 248 
<< m1 >>
rect 243 247 244 248 
<< pdiffusion >>
rect 246 247 247 248 
<< pdiffusion >>
rect 247 247 248 248 
<< pdiffusion >>
rect 248 247 249 248 
<< pdiffusion >>
rect 249 247 250 248 
<< pdiffusion >>
rect 250 247 251 248 
<< pdiffusion >>
rect 251 247 252 248 
<< m1 >>
rect 262 247 263 248 
<< pdiffusion >>
rect 264 247 265 248 
<< pdiffusion >>
rect 265 247 266 248 
<< pdiffusion >>
rect 266 247 267 248 
<< pdiffusion >>
rect 267 247 268 248 
<< pdiffusion >>
rect 268 247 269 248 
<< pdiffusion >>
rect 269 247 270 248 
<< m1 >>
rect 272 247 273 248 
<< m2 >>
rect 273 247 274 248 
<< m2 >>
rect 279 247 280 248 
<< m1 >>
rect 280 247 281 248 
<< pdiffusion >>
rect 282 247 283 248 
<< pdiffusion >>
rect 283 247 284 248 
<< pdiffusion >>
rect 284 247 285 248 
<< pdiffusion >>
rect 285 247 286 248 
<< pdiffusion >>
rect 286 247 287 248 
<< pdiffusion >>
rect 287 247 288 248 
<< m1 >>
rect 294 247 295 248 
<< m1 >>
rect 298 247 299 248 
<< pdiffusion >>
rect 300 247 301 248 
<< pdiffusion >>
rect 301 247 302 248 
<< pdiffusion >>
rect 302 247 303 248 
<< pdiffusion >>
rect 303 247 304 248 
<< pdiffusion >>
rect 304 247 305 248 
<< pdiffusion >>
rect 305 247 306 248 
<< pdiffusion >>
rect 318 247 319 248 
<< pdiffusion >>
rect 319 247 320 248 
<< pdiffusion >>
rect 320 247 321 248 
<< pdiffusion >>
rect 321 247 322 248 
<< pdiffusion >>
rect 322 247 323 248 
<< pdiffusion >>
rect 323 247 324 248 
<< m1 >>
rect 327 247 328 248 
<< m1 >>
rect 329 247 330 248 
<< m2 >>
rect 330 247 331 248 
<< pdiffusion >>
rect 336 247 337 248 
<< pdiffusion >>
rect 337 247 338 248 
<< pdiffusion >>
rect 338 247 339 248 
<< pdiffusion >>
rect 339 247 340 248 
<< pdiffusion >>
rect 340 247 341 248 
<< pdiffusion >>
rect 341 247 342 248 
<< m1 >>
rect 10 248 11 249 
<< pdiffusion >>
rect 12 248 13 249 
<< pdiffusion >>
rect 13 248 14 249 
<< pdiffusion >>
rect 14 248 15 249 
<< pdiffusion >>
rect 15 248 16 249 
<< pdiffusion >>
rect 16 248 17 249 
<< pdiffusion >>
rect 17 248 18 249 
<< m1 >>
rect 28 248 29 249 
<< m2 >>
rect 28 248 29 249 
<< pdiffusion >>
rect 30 248 31 249 
<< pdiffusion >>
rect 31 248 32 249 
<< pdiffusion >>
rect 32 248 33 249 
<< pdiffusion >>
rect 33 248 34 249 
<< pdiffusion >>
rect 34 248 35 249 
<< pdiffusion >>
rect 35 248 36 249 
<< m1 >>
rect 37 248 38 249 
<< m2 >>
rect 37 248 38 249 
<< m1 >>
rect 39 248 40 249 
<< m2 >>
rect 43 248 44 249 
<< m1 >>
rect 44 248 45 249 
<< m1 >>
rect 46 248 47 249 
<< m2 >>
rect 46 248 47 249 
<< pdiffusion >>
rect 48 248 49 249 
<< pdiffusion >>
rect 49 248 50 249 
<< pdiffusion >>
rect 50 248 51 249 
<< pdiffusion >>
rect 51 248 52 249 
<< pdiffusion >>
rect 52 248 53 249 
<< pdiffusion >>
rect 53 248 54 249 
<< m1 >>
rect 56 248 57 249 
<< m1 >>
rect 58 248 59 249 
<< m1 >>
rect 60 248 61 249 
<< m1 >>
rect 64 248 65 249 
<< pdiffusion >>
rect 66 248 67 249 
<< pdiffusion >>
rect 67 248 68 249 
<< pdiffusion >>
rect 68 248 69 249 
<< pdiffusion >>
rect 69 248 70 249 
<< pdiffusion >>
rect 70 248 71 249 
<< pdiffusion >>
rect 71 248 72 249 
<< m1 >>
rect 73 248 74 249 
<< m2 >>
rect 74 248 75 249 
<< pdiffusion >>
rect 84 248 85 249 
<< pdiffusion >>
rect 85 248 86 249 
<< pdiffusion >>
rect 86 248 87 249 
<< pdiffusion >>
rect 87 248 88 249 
<< pdiffusion >>
rect 88 248 89 249 
<< pdiffusion >>
rect 89 248 90 249 
<< m1 >>
rect 100 248 101 249 
<< pdiffusion >>
rect 102 248 103 249 
<< pdiffusion >>
rect 103 248 104 249 
<< pdiffusion >>
rect 104 248 105 249 
<< pdiffusion >>
rect 105 248 106 249 
<< pdiffusion >>
rect 106 248 107 249 
<< pdiffusion >>
rect 107 248 108 249 
<< m1 >>
rect 116 248 117 249 
<< m1 >>
rect 118 248 119 249 
<< pdiffusion >>
rect 120 248 121 249 
<< pdiffusion >>
rect 121 248 122 249 
<< pdiffusion >>
rect 122 248 123 249 
<< pdiffusion >>
rect 123 248 124 249 
<< pdiffusion >>
rect 124 248 125 249 
<< pdiffusion >>
rect 125 248 126 249 
<< m1 >>
rect 128 248 129 249 
<< m1 >>
rect 130 248 131 249 
<< m1 >>
rect 132 248 133 249 
<< m1 >>
rect 134 248 135 249 
<< m1 >>
rect 136 248 137 249 
<< pdiffusion >>
rect 138 248 139 249 
<< pdiffusion >>
rect 139 248 140 249 
<< pdiffusion >>
rect 140 248 141 249 
<< pdiffusion >>
rect 141 248 142 249 
<< pdiffusion >>
rect 142 248 143 249 
<< pdiffusion >>
rect 143 248 144 249 
<< m1 >>
rect 145 248 146 249 
<< m2 >>
rect 145 248 146 249 
<< m1 >>
rect 154 248 155 249 
<< m2 >>
rect 154 248 155 249 
<< pdiffusion >>
rect 156 248 157 249 
<< pdiffusion >>
rect 157 248 158 249 
<< pdiffusion >>
rect 158 248 159 249 
<< pdiffusion >>
rect 159 248 160 249 
<< pdiffusion >>
rect 160 248 161 249 
<< pdiffusion >>
rect 161 248 162 249 
<< m1 >>
rect 163 248 164 249 
<< m1 >>
rect 165 248 166 249 
<< m1 >>
rect 167 248 168 249 
<< m1 >>
rect 171 248 172 249 
<< pdiffusion >>
rect 174 248 175 249 
<< pdiffusion >>
rect 175 248 176 249 
<< pdiffusion >>
rect 176 248 177 249 
<< pdiffusion >>
rect 177 248 178 249 
<< pdiffusion >>
rect 178 248 179 249 
<< pdiffusion >>
rect 179 248 180 249 
<< m1 >>
rect 181 248 182 249 
<< m1 >>
rect 183 248 184 249 
<< m1 >>
rect 186 248 187 249 
<< m1 >>
rect 188 248 189 249 
<< m1 >>
rect 190 248 191 249 
<< pdiffusion >>
rect 192 248 193 249 
<< pdiffusion >>
rect 193 248 194 249 
<< pdiffusion >>
rect 194 248 195 249 
<< pdiffusion >>
rect 195 248 196 249 
<< pdiffusion >>
rect 196 248 197 249 
<< pdiffusion >>
rect 197 248 198 249 
<< m1 >>
rect 199 248 200 249 
<< pdiffusion >>
rect 210 248 211 249 
<< pdiffusion >>
rect 211 248 212 249 
<< pdiffusion >>
rect 212 248 213 249 
<< pdiffusion >>
rect 213 248 214 249 
<< pdiffusion >>
rect 214 248 215 249 
<< pdiffusion >>
rect 215 248 216 249 
<< m1 >>
rect 226 248 227 249 
<< pdiffusion >>
rect 228 248 229 249 
<< pdiffusion >>
rect 229 248 230 249 
<< pdiffusion >>
rect 230 248 231 249 
<< pdiffusion >>
rect 231 248 232 249 
<< pdiffusion >>
rect 232 248 233 249 
<< pdiffusion >>
rect 233 248 234 249 
<< m1 >>
rect 235 248 236 249 
<< m1 >>
rect 237 248 238 249 
<< m1 >>
rect 239 248 240 249 
<< m1 >>
rect 243 248 244 249 
<< pdiffusion >>
rect 246 248 247 249 
<< pdiffusion >>
rect 247 248 248 249 
<< pdiffusion >>
rect 248 248 249 249 
<< pdiffusion >>
rect 249 248 250 249 
<< pdiffusion >>
rect 250 248 251 249 
<< pdiffusion >>
rect 251 248 252 249 
<< m1 >>
rect 262 248 263 249 
<< pdiffusion >>
rect 264 248 265 249 
<< pdiffusion >>
rect 265 248 266 249 
<< pdiffusion >>
rect 266 248 267 249 
<< pdiffusion >>
rect 267 248 268 249 
<< pdiffusion >>
rect 268 248 269 249 
<< pdiffusion >>
rect 269 248 270 249 
<< m1 >>
rect 272 248 273 249 
<< m2 >>
rect 273 248 274 249 
<< m2 >>
rect 279 248 280 249 
<< m1 >>
rect 280 248 281 249 
<< pdiffusion >>
rect 282 248 283 249 
<< pdiffusion >>
rect 283 248 284 249 
<< pdiffusion >>
rect 284 248 285 249 
<< pdiffusion >>
rect 285 248 286 249 
<< pdiffusion >>
rect 286 248 287 249 
<< pdiffusion >>
rect 287 248 288 249 
<< m1 >>
rect 294 248 295 249 
<< m1 >>
rect 298 248 299 249 
<< pdiffusion >>
rect 300 248 301 249 
<< pdiffusion >>
rect 301 248 302 249 
<< pdiffusion >>
rect 302 248 303 249 
<< pdiffusion >>
rect 303 248 304 249 
<< pdiffusion >>
rect 304 248 305 249 
<< pdiffusion >>
rect 305 248 306 249 
<< pdiffusion >>
rect 318 248 319 249 
<< pdiffusion >>
rect 319 248 320 249 
<< pdiffusion >>
rect 320 248 321 249 
<< pdiffusion >>
rect 321 248 322 249 
<< pdiffusion >>
rect 322 248 323 249 
<< pdiffusion >>
rect 323 248 324 249 
<< m1 >>
rect 327 248 328 249 
<< m1 >>
rect 329 248 330 249 
<< m2 >>
rect 330 248 331 249 
<< pdiffusion >>
rect 336 248 337 249 
<< pdiffusion >>
rect 337 248 338 249 
<< pdiffusion >>
rect 338 248 339 249 
<< pdiffusion >>
rect 339 248 340 249 
<< pdiffusion >>
rect 340 248 341 249 
<< pdiffusion >>
rect 341 248 342 249 
<< m1 >>
rect 10 249 11 250 
<< pdiffusion >>
rect 12 249 13 250 
<< pdiffusion >>
rect 13 249 14 250 
<< pdiffusion >>
rect 14 249 15 250 
<< pdiffusion >>
rect 15 249 16 250 
<< pdiffusion >>
rect 16 249 17 250 
<< pdiffusion >>
rect 17 249 18 250 
<< m1 >>
rect 28 249 29 250 
<< m2 >>
rect 28 249 29 250 
<< pdiffusion >>
rect 30 249 31 250 
<< pdiffusion >>
rect 31 249 32 250 
<< pdiffusion >>
rect 32 249 33 250 
<< pdiffusion >>
rect 33 249 34 250 
<< pdiffusion >>
rect 34 249 35 250 
<< pdiffusion >>
rect 35 249 36 250 
<< m1 >>
rect 37 249 38 250 
<< m2 >>
rect 37 249 38 250 
<< m1 >>
rect 39 249 40 250 
<< m2 >>
rect 43 249 44 250 
<< m1 >>
rect 44 249 45 250 
<< m1 >>
rect 46 249 47 250 
<< m2 >>
rect 46 249 47 250 
<< pdiffusion >>
rect 48 249 49 250 
<< pdiffusion >>
rect 49 249 50 250 
<< pdiffusion >>
rect 50 249 51 250 
<< pdiffusion >>
rect 51 249 52 250 
<< pdiffusion >>
rect 52 249 53 250 
<< pdiffusion >>
rect 53 249 54 250 
<< m1 >>
rect 56 249 57 250 
<< m1 >>
rect 58 249 59 250 
<< m1 >>
rect 60 249 61 250 
<< m1 >>
rect 64 249 65 250 
<< pdiffusion >>
rect 66 249 67 250 
<< pdiffusion >>
rect 67 249 68 250 
<< pdiffusion >>
rect 68 249 69 250 
<< pdiffusion >>
rect 69 249 70 250 
<< pdiffusion >>
rect 70 249 71 250 
<< pdiffusion >>
rect 71 249 72 250 
<< m1 >>
rect 73 249 74 250 
<< m2 >>
rect 74 249 75 250 
<< pdiffusion >>
rect 84 249 85 250 
<< pdiffusion >>
rect 85 249 86 250 
<< pdiffusion >>
rect 86 249 87 250 
<< pdiffusion >>
rect 87 249 88 250 
<< pdiffusion >>
rect 88 249 89 250 
<< pdiffusion >>
rect 89 249 90 250 
<< m1 >>
rect 100 249 101 250 
<< pdiffusion >>
rect 102 249 103 250 
<< pdiffusion >>
rect 103 249 104 250 
<< pdiffusion >>
rect 104 249 105 250 
<< pdiffusion >>
rect 105 249 106 250 
<< pdiffusion >>
rect 106 249 107 250 
<< pdiffusion >>
rect 107 249 108 250 
<< m1 >>
rect 116 249 117 250 
<< m1 >>
rect 118 249 119 250 
<< pdiffusion >>
rect 120 249 121 250 
<< pdiffusion >>
rect 121 249 122 250 
<< pdiffusion >>
rect 122 249 123 250 
<< pdiffusion >>
rect 123 249 124 250 
<< pdiffusion >>
rect 124 249 125 250 
<< pdiffusion >>
rect 125 249 126 250 
<< m1 >>
rect 128 249 129 250 
<< m1 >>
rect 130 249 131 250 
<< m1 >>
rect 132 249 133 250 
<< m1 >>
rect 134 249 135 250 
<< m1 >>
rect 136 249 137 250 
<< pdiffusion >>
rect 138 249 139 250 
<< pdiffusion >>
rect 139 249 140 250 
<< pdiffusion >>
rect 140 249 141 250 
<< pdiffusion >>
rect 141 249 142 250 
<< pdiffusion >>
rect 142 249 143 250 
<< pdiffusion >>
rect 143 249 144 250 
<< m1 >>
rect 145 249 146 250 
<< m2 >>
rect 145 249 146 250 
<< m1 >>
rect 154 249 155 250 
<< m2 >>
rect 154 249 155 250 
<< pdiffusion >>
rect 156 249 157 250 
<< pdiffusion >>
rect 157 249 158 250 
<< pdiffusion >>
rect 158 249 159 250 
<< pdiffusion >>
rect 159 249 160 250 
<< pdiffusion >>
rect 160 249 161 250 
<< pdiffusion >>
rect 161 249 162 250 
<< m1 >>
rect 163 249 164 250 
<< m1 >>
rect 165 249 166 250 
<< m1 >>
rect 167 249 168 250 
<< m1 >>
rect 171 249 172 250 
<< pdiffusion >>
rect 174 249 175 250 
<< pdiffusion >>
rect 175 249 176 250 
<< pdiffusion >>
rect 176 249 177 250 
<< pdiffusion >>
rect 177 249 178 250 
<< pdiffusion >>
rect 178 249 179 250 
<< pdiffusion >>
rect 179 249 180 250 
<< m1 >>
rect 181 249 182 250 
<< m1 >>
rect 183 249 184 250 
<< m1 >>
rect 186 249 187 250 
<< m1 >>
rect 188 249 189 250 
<< m1 >>
rect 190 249 191 250 
<< pdiffusion >>
rect 192 249 193 250 
<< pdiffusion >>
rect 193 249 194 250 
<< pdiffusion >>
rect 194 249 195 250 
<< pdiffusion >>
rect 195 249 196 250 
<< pdiffusion >>
rect 196 249 197 250 
<< pdiffusion >>
rect 197 249 198 250 
<< m1 >>
rect 199 249 200 250 
<< pdiffusion >>
rect 210 249 211 250 
<< pdiffusion >>
rect 211 249 212 250 
<< pdiffusion >>
rect 212 249 213 250 
<< pdiffusion >>
rect 213 249 214 250 
<< pdiffusion >>
rect 214 249 215 250 
<< pdiffusion >>
rect 215 249 216 250 
<< m1 >>
rect 226 249 227 250 
<< pdiffusion >>
rect 228 249 229 250 
<< pdiffusion >>
rect 229 249 230 250 
<< pdiffusion >>
rect 230 249 231 250 
<< pdiffusion >>
rect 231 249 232 250 
<< pdiffusion >>
rect 232 249 233 250 
<< pdiffusion >>
rect 233 249 234 250 
<< m1 >>
rect 235 249 236 250 
<< m1 >>
rect 237 249 238 250 
<< m1 >>
rect 239 249 240 250 
<< m1 >>
rect 243 249 244 250 
<< pdiffusion >>
rect 246 249 247 250 
<< pdiffusion >>
rect 247 249 248 250 
<< pdiffusion >>
rect 248 249 249 250 
<< pdiffusion >>
rect 249 249 250 250 
<< pdiffusion >>
rect 250 249 251 250 
<< pdiffusion >>
rect 251 249 252 250 
<< m1 >>
rect 262 249 263 250 
<< pdiffusion >>
rect 264 249 265 250 
<< pdiffusion >>
rect 265 249 266 250 
<< pdiffusion >>
rect 266 249 267 250 
<< pdiffusion >>
rect 267 249 268 250 
<< pdiffusion >>
rect 268 249 269 250 
<< pdiffusion >>
rect 269 249 270 250 
<< m1 >>
rect 272 249 273 250 
<< m2 >>
rect 273 249 274 250 
<< m2 >>
rect 279 249 280 250 
<< m1 >>
rect 280 249 281 250 
<< pdiffusion >>
rect 282 249 283 250 
<< pdiffusion >>
rect 283 249 284 250 
<< pdiffusion >>
rect 284 249 285 250 
<< pdiffusion >>
rect 285 249 286 250 
<< pdiffusion >>
rect 286 249 287 250 
<< pdiffusion >>
rect 287 249 288 250 
<< m1 >>
rect 294 249 295 250 
<< m1 >>
rect 298 249 299 250 
<< pdiffusion >>
rect 300 249 301 250 
<< pdiffusion >>
rect 301 249 302 250 
<< pdiffusion >>
rect 302 249 303 250 
<< pdiffusion >>
rect 303 249 304 250 
<< pdiffusion >>
rect 304 249 305 250 
<< pdiffusion >>
rect 305 249 306 250 
<< pdiffusion >>
rect 318 249 319 250 
<< pdiffusion >>
rect 319 249 320 250 
<< pdiffusion >>
rect 320 249 321 250 
<< pdiffusion >>
rect 321 249 322 250 
<< pdiffusion >>
rect 322 249 323 250 
<< pdiffusion >>
rect 323 249 324 250 
<< m1 >>
rect 327 249 328 250 
<< m1 >>
rect 329 249 330 250 
<< m2 >>
rect 330 249 331 250 
<< pdiffusion >>
rect 336 249 337 250 
<< pdiffusion >>
rect 337 249 338 250 
<< pdiffusion >>
rect 338 249 339 250 
<< pdiffusion >>
rect 339 249 340 250 
<< pdiffusion >>
rect 340 249 341 250 
<< pdiffusion >>
rect 341 249 342 250 
<< m1 >>
rect 10 250 11 251 
<< pdiffusion >>
rect 12 250 13 251 
<< pdiffusion >>
rect 13 250 14 251 
<< pdiffusion >>
rect 14 250 15 251 
<< pdiffusion >>
rect 15 250 16 251 
<< pdiffusion >>
rect 16 250 17 251 
<< pdiffusion >>
rect 17 250 18 251 
<< m1 >>
rect 28 250 29 251 
<< m2 >>
rect 28 250 29 251 
<< pdiffusion >>
rect 30 250 31 251 
<< pdiffusion >>
rect 31 250 32 251 
<< pdiffusion >>
rect 32 250 33 251 
<< pdiffusion >>
rect 33 250 34 251 
<< pdiffusion >>
rect 34 250 35 251 
<< pdiffusion >>
rect 35 250 36 251 
<< m1 >>
rect 37 250 38 251 
<< m2 >>
rect 37 250 38 251 
<< m1 >>
rect 39 250 40 251 
<< m2 >>
rect 43 250 44 251 
<< m1 >>
rect 44 250 45 251 
<< m1 >>
rect 46 250 47 251 
<< m2 >>
rect 46 250 47 251 
<< pdiffusion >>
rect 48 250 49 251 
<< pdiffusion >>
rect 49 250 50 251 
<< pdiffusion >>
rect 50 250 51 251 
<< pdiffusion >>
rect 51 250 52 251 
<< pdiffusion >>
rect 52 250 53 251 
<< pdiffusion >>
rect 53 250 54 251 
<< m1 >>
rect 56 250 57 251 
<< m1 >>
rect 58 250 59 251 
<< m1 >>
rect 60 250 61 251 
<< m1 >>
rect 64 250 65 251 
<< pdiffusion >>
rect 66 250 67 251 
<< pdiffusion >>
rect 67 250 68 251 
<< pdiffusion >>
rect 68 250 69 251 
<< pdiffusion >>
rect 69 250 70 251 
<< pdiffusion >>
rect 70 250 71 251 
<< pdiffusion >>
rect 71 250 72 251 
<< m1 >>
rect 73 250 74 251 
<< m2 >>
rect 74 250 75 251 
<< pdiffusion >>
rect 84 250 85 251 
<< pdiffusion >>
rect 85 250 86 251 
<< pdiffusion >>
rect 86 250 87 251 
<< pdiffusion >>
rect 87 250 88 251 
<< pdiffusion >>
rect 88 250 89 251 
<< pdiffusion >>
rect 89 250 90 251 
<< m1 >>
rect 100 250 101 251 
<< pdiffusion >>
rect 102 250 103 251 
<< pdiffusion >>
rect 103 250 104 251 
<< pdiffusion >>
rect 104 250 105 251 
<< pdiffusion >>
rect 105 250 106 251 
<< pdiffusion >>
rect 106 250 107 251 
<< pdiffusion >>
rect 107 250 108 251 
<< m1 >>
rect 116 250 117 251 
<< m1 >>
rect 118 250 119 251 
<< pdiffusion >>
rect 120 250 121 251 
<< pdiffusion >>
rect 121 250 122 251 
<< pdiffusion >>
rect 122 250 123 251 
<< pdiffusion >>
rect 123 250 124 251 
<< pdiffusion >>
rect 124 250 125 251 
<< pdiffusion >>
rect 125 250 126 251 
<< m1 >>
rect 128 250 129 251 
<< m1 >>
rect 130 250 131 251 
<< m1 >>
rect 132 250 133 251 
<< m1 >>
rect 134 250 135 251 
<< m1 >>
rect 136 250 137 251 
<< pdiffusion >>
rect 138 250 139 251 
<< pdiffusion >>
rect 139 250 140 251 
<< pdiffusion >>
rect 140 250 141 251 
<< pdiffusion >>
rect 141 250 142 251 
<< pdiffusion >>
rect 142 250 143 251 
<< pdiffusion >>
rect 143 250 144 251 
<< m1 >>
rect 145 250 146 251 
<< m2 >>
rect 145 250 146 251 
<< m1 >>
rect 154 250 155 251 
<< m2 >>
rect 154 250 155 251 
<< pdiffusion >>
rect 156 250 157 251 
<< pdiffusion >>
rect 157 250 158 251 
<< pdiffusion >>
rect 158 250 159 251 
<< pdiffusion >>
rect 159 250 160 251 
<< pdiffusion >>
rect 160 250 161 251 
<< pdiffusion >>
rect 161 250 162 251 
<< m1 >>
rect 163 250 164 251 
<< m1 >>
rect 165 250 166 251 
<< m1 >>
rect 167 250 168 251 
<< m1 >>
rect 171 250 172 251 
<< pdiffusion >>
rect 174 250 175 251 
<< pdiffusion >>
rect 175 250 176 251 
<< pdiffusion >>
rect 176 250 177 251 
<< pdiffusion >>
rect 177 250 178 251 
<< pdiffusion >>
rect 178 250 179 251 
<< pdiffusion >>
rect 179 250 180 251 
<< m1 >>
rect 181 250 182 251 
<< m1 >>
rect 183 250 184 251 
<< m1 >>
rect 186 250 187 251 
<< m1 >>
rect 188 250 189 251 
<< m1 >>
rect 190 250 191 251 
<< pdiffusion >>
rect 192 250 193 251 
<< pdiffusion >>
rect 193 250 194 251 
<< pdiffusion >>
rect 194 250 195 251 
<< pdiffusion >>
rect 195 250 196 251 
<< pdiffusion >>
rect 196 250 197 251 
<< pdiffusion >>
rect 197 250 198 251 
<< m1 >>
rect 199 250 200 251 
<< pdiffusion >>
rect 210 250 211 251 
<< pdiffusion >>
rect 211 250 212 251 
<< pdiffusion >>
rect 212 250 213 251 
<< pdiffusion >>
rect 213 250 214 251 
<< pdiffusion >>
rect 214 250 215 251 
<< pdiffusion >>
rect 215 250 216 251 
<< m1 >>
rect 226 250 227 251 
<< pdiffusion >>
rect 228 250 229 251 
<< pdiffusion >>
rect 229 250 230 251 
<< pdiffusion >>
rect 230 250 231 251 
<< pdiffusion >>
rect 231 250 232 251 
<< pdiffusion >>
rect 232 250 233 251 
<< pdiffusion >>
rect 233 250 234 251 
<< m1 >>
rect 235 250 236 251 
<< m1 >>
rect 237 250 238 251 
<< m1 >>
rect 239 250 240 251 
<< m1 >>
rect 243 250 244 251 
<< pdiffusion >>
rect 246 250 247 251 
<< pdiffusion >>
rect 247 250 248 251 
<< pdiffusion >>
rect 248 250 249 251 
<< pdiffusion >>
rect 249 250 250 251 
<< pdiffusion >>
rect 250 250 251 251 
<< pdiffusion >>
rect 251 250 252 251 
<< m1 >>
rect 262 250 263 251 
<< pdiffusion >>
rect 264 250 265 251 
<< pdiffusion >>
rect 265 250 266 251 
<< pdiffusion >>
rect 266 250 267 251 
<< pdiffusion >>
rect 267 250 268 251 
<< pdiffusion >>
rect 268 250 269 251 
<< pdiffusion >>
rect 269 250 270 251 
<< m1 >>
rect 272 250 273 251 
<< m2 >>
rect 273 250 274 251 
<< m2 >>
rect 279 250 280 251 
<< m1 >>
rect 280 250 281 251 
<< pdiffusion >>
rect 282 250 283 251 
<< pdiffusion >>
rect 283 250 284 251 
<< pdiffusion >>
rect 284 250 285 251 
<< pdiffusion >>
rect 285 250 286 251 
<< pdiffusion >>
rect 286 250 287 251 
<< pdiffusion >>
rect 287 250 288 251 
<< m1 >>
rect 294 250 295 251 
<< m1 >>
rect 298 250 299 251 
<< pdiffusion >>
rect 300 250 301 251 
<< pdiffusion >>
rect 301 250 302 251 
<< pdiffusion >>
rect 302 250 303 251 
<< pdiffusion >>
rect 303 250 304 251 
<< pdiffusion >>
rect 304 250 305 251 
<< pdiffusion >>
rect 305 250 306 251 
<< pdiffusion >>
rect 318 250 319 251 
<< pdiffusion >>
rect 319 250 320 251 
<< pdiffusion >>
rect 320 250 321 251 
<< pdiffusion >>
rect 321 250 322 251 
<< pdiffusion >>
rect 322 250 323 251 
<< pdiffusion >>
rect 323 250 324 251 
<< m1 >>
rect 327 250 328 251 
<< m1 >>
rect 329 250 330 251 
<< m2 >>
rect 330 250 331 251 
<< pdiffusion >>
rect 336 250 337 251 
<< pdiffusion >>
rect 337 250 338 251 
<< pdiffusion >>
rect 338 250 339 251 
<< pdiffusion >>
rect 339 250 340 251 
<< pdiffusion >>
rect 340 250 341 251 
<< pdiffusion >>
rect 341 250 342 251 
<< m1 >>
rect 10 251 11 252 
<< pdiffusion >>
rect 12 251 13 252 
<< pdiffusion >>
rect 13 251 14 252 
<< pdiffusion >>
rect 14 251 15 252 
<< pdiffusion >>
rect 15 251 16 252 
<< pdiffusion >>
rect 16 251 17 252 
<< pdiffusion >>
rect 17 251 18 252 
<< m1 >>
rect 28 251 29 252 
<< m2 >>
rect 28 251 29 252 
<< pdiffusion >>
rect 30 251 31 252 
<< pdiffusion >>
rect 31 251 32 252 
<< pdiffusion >>
rect 32 251 33 252 
<< pdiffusion >>
rect 33 251 34 252 
<< pdiffusion >>
rect 34 251 35 252 
<< pdiffusion >>
rect 35 251 36 252 
<< m1 >>
rect 37 251 38 252 
<< m2 >>
rect 37 251 38 252 
<< m1 >>
rect 39 251 40 252 
<< m2 >>
rect 43 251 44 252 
<< m1 >>
rect 44 251 45 252 
<< m1 >>
rect 46 251 47 252 
<< m2 >>
rect 46 251 47 252 
<< pdiffusion >>
rect 48 251 49 252 
<< m1 >>
rect 49 251 50 252 
<< pdiffusion >>
rect 49 251 50 252 
<< pdiffusion >>
rect 50 251 51 252 
<< pdiffusion >>
rect 51 251 52 252 
<< pdiffusion >>
rect 52 251 53 252 
<< pdiffusion >>
rect 53 251 54 252 
<< m1 >>
rect 56 251 57 252 
<< m1 >>
rect 58 251 59 252 
<< m1 >>
rect 60 251 61 252 
<< m1 >>
rect 64 251 65 252 
<< pdiffusion >>
rect 66 251 67 252 
<< pdiffusion >>
rect 67 251 68 252 
<< pdiffusion >>
rect 68 251 69 252 
<< pdiffusion >>
rect 69 251 70 252 
<< pdiffusion >>
rect 70 251 71 252 
<< pdiffusion >>
rect 71 251 72 252 
<< m1 >>
rect 73 251 74 252 
<< m2 >>
rect 74 251 75 252 
<< pdiffusion >>
rect 84 251 85 252 
<< pdiffusion >>
rect 85 251 86 252 
<< pdiffusion >>
rect 86 251 87 252 
<< pdiffusion >>
rect 87 251 88 252 
<< pdiffusion >>
rect 88 251 89 252 
<< pdiffusion >>
rect 89 251 90 252 
<< m1 >>
rect 100 251 101 252 
<< pdiffusion >>
rect 102 251 103 252 
<< pdiffusion >>
rect 103 251 104 252 
<< pdiffusion >>
rect 104 251 105 252 
<< pdiffusion >>
rect 105 251 106 252 
<< pdiffusion >>
rect 106 251 107 252 
<< pdiffusion >>
rect 107 251 108 252 
<< m1 >>
rect 116 251 117 252 
<< m1 >>
rect 118 251 119 252 
<< pdiffusion >>
rect 120 251 121 252 
<< m1 >>
rect 121 251 122 252 
<< pdiffusion >>
rect 121 251 122 252 
<< pdiffusion >>
rect 122 251 123 252 
<< pdiffusion >>
rect 123 251 124 252 
<< pdiffusion >>
rect 124 251 125 252 
<< pdiffusion >>
rect 125 251 126 252 
<< m1 >>
rect 128 251 129 252 
<< m1 >>
rect 130 251 131 252 
<< m1 >>
rect 132 251 133 252 
<< m1 >>
rect 134 251 135 252 
<< m1 >>
rect 136 251 137 252 
<< pdiffusion >>
rect 138 251 139 252 
<< pdiffusion >>
rect 139 251 140 252 
<< pdiffusion >>
rect 140 251 141 252 
<< pdiffusion >>
rect 141 251 142 252 
<< m1 >>
rect 142 251 143 252 
<< pdiffusion >>
rect 142 251 143 252 
<< pdiffusion >>
rect 143 251 144 252 
<< m1 >>
rect 145 251 146 252 
<< m2 >>
rect 145 251 146 252 
<< m1 >>
rect 154 251 155 252 
<< m2 >>
rect 154 251 155 252 
<< pdiffusion >>
rect 156 251 157 252 
<< pdiffusion >>
rect 157 251 158 252 
<< pdiffusion >>
rect 158 251 159 252 
<< pdiffusion >>
rect 159 251 160 252 
<< pdiffusion >>
rect 160 251 161 252 
<< pdiffusion >>
rect 161 251 162 252 
<< m1 >>
rect 163 251 164 252 
<< m1 >>
rect 165 251 166 252 
<< m1 >>
rect 167 251 168 252 
<< m1 >>
rect 171 251 172 252 
<< pdiffusion >>
rect 174 251 175 252 
<< pdiffusion >>
rect 175 251 176 252 
<< pdiffusion >>
rect 176 251 177 252 
<< pdiffusion >>
rect 177 251 178 252 
<< m1 >>
rect 178 251 179 252 
<< pdiffusion >>
rect 178 251 179 252 
<< pdiffusion >>
rect 179 251 180 252 
<< m1 >>
rect 181 251 182 252 
<< m1 >>
rect 183 251 184 252 
<< m1 >>
rect 186 251 187 252 
<< m1 >>
rect 188 251 189 252 
<< m1 >>
rect 190 251 191 252 
<< pdiffusion >>
rect 192 251 193 252 
<< pdiffusion >>
rect 193 251 194 252 
<< pdiffusion >>
rect 194 251 195 252 
<< pdiffusion >>
rect 195 251 196 252 
<< pdiffusion >>
rect 196 251 197 252 
<< pdiffusion >>
rect 197 251 198 252 
<< m1 >>
rect 199 251 200 252 
<< pdiffusion >>
rect 210 251 211 252 
<< m1 >>
rect 211 251 212 252 
<< pdiffusion >>
rect 211 251 212 252 
<< pdiffusion >>
rect 212 251 213 252 
<< pdiffusion >>
rect 213 251 214 252 
<< pdiffusion >>
rect 214 251 215 252 
<< pdiffusion >>
rect 215 251 216 252 
<< m1 >>
rect 226 251 227 252 
<< pdiffusion >>
rect 228 251 229 252 
<< pdiffusion >>
rect 229 251 230 252 
<< pdiffusion >>
rect 230 251 231 252 
<< pdiffusion >>
rect 231 251 232 252 
<< m1 >>
rect 232 251 233 252 
<< pdiffusion >>
rect 232 251 233 252 
<< pdiffusion >>
rect 233 251 234 252 
<< m1 >>
rect 235 251 236 252 
<< m1 >>
rect 237 251 238 252 
<< m1 >>
rect 239 251 240 252 
<< m1 >>
rect 243 251 244 252 
<< pdiffusion >>
rect 246 251 247 252 
<< m1 >>
rect 247 251 248 252 
<< pdiffusion >>
rect 247 251 248 252 
<< pdiffusion >>
rect 248 251 249 252 
<< pdiffusion >>
rect 249 251 250 252 
<< pdiffusion >>
rect 250 251 251 252 
<< pdiffusion >>
rect 251 251 252 252 
<< m1 >>
rect 262 251 263 252 
<< pdiffusion >>
rect 264 251 265 252 
<< pdiffusion >>
rect 265 251 266 252 
<< pdiffusion >>
rect 266 251 267 252 
<< pdiffusion >>
rect 267 251 268 252 
<< pdiffusion >>
rect 268 251 269 252 
<< pdiffusion >>
rect 269 251 270 252 
<< m1 >>
rect 272 251 273 252 
<< m2 >>
rect 273 251 274 252 
<< m2 >>
rect 279 251 280 252 
<< m1 >>
rect 280 251 281 252 
<< pdiffusion >>
rect 282 251 283 252 
<< m1 >>
rect 283 251 284 252 
<< pdiffusion >>
rect 283 251 284 252 
<< pdiffusion >>
rect 284 251 285 252 
<< pdiffusion >>
rect 285 251 286 252 
<< m1 >>
rect 286 251 287 252 
<< pdiffusion >>
rect 286 251 287 252 
<< pdiffusion >>
rect 287 251 288 252 
<< m1 >>
rect 294 251 295 252 
<< m1 >>
rect 298 251 299 252 
<< pdiffusion >>
rect 300 251 301 252 
<< pdiffusion >>
rect 301 251 302 252 
<< pdiffusion >>
rect 302 251 303 252 
<< pdiffusion >>
rect 303 251 304 252 
<< pdiffusion >>
rect 304 251 305 252 
<< pdiffusion >>
rect 305 251 306 252 
<< pdiffusion >>
rect 318 251 319 252 
<< pdiffusion >>
rect 319 251 320 252 
<< pdiffusion >>
rect 320 251 321 252 
<< pdiffusion >>
rect 321 251 322 252 
<< pdiffusion >>
rect 322 251 323 252 
<< pdiffusion >>
rect 323 251 324 252 
<< m1 >>
rect 327 251 328 252 
<< m1 >>
rect 329 251 330 252 
<< m2 >>
rect 330 251 331 252 
<< pdiffusion >>
rect 336 251 337 252 
<< pdiffusion >>
rect 337 251 338 252 
<< pdiffusion >>
rect 338 251 339 252 
<< pdiffusion >>
rect 339 251 340 252 
<< pdiffusion >>
rect 340 251 341 252 
<< pdiffusion >>
rect 341 251 342 252 
<< m1 >>
rect 10 252 11 253 
<< m1 >>
rect 28 252 29 253 
<< m2 >>
rect 28 252 29 253 
<< m1 >>
rect 37 252 38 253 
<< m2 >>
rect 37 252 38 253 
<< m1 >>
rect 39 252 40 253 
<< m2 >>
rect 43 252 44 253 
<< m1 >>
rect 44 252 45 253 
<< m1 >>
rect 46 252 47 253 
<< m2 >>
rect 46 252 47 253 
<< m1 >>
rect 49 252 50 253 
<< m1 >>
rect 56 252 57 253 
<< m2 >>
rect 56 252 57 253 
<< m2c >>
rect 56 252 57 253 
<< m1 >>
rect 56 252 57 253 
<< m2 >>
rect 56 252 57 253 
<< m1 >>
rect 58 252 59 253 
<< m2 >>
rect 58 252 59 253 
<< m2c >>
rect 58 252 59 253 
<< m1 >>
rect 58 252 59 253 
<< m2 >>
rect 58 252 59 253 
<< m2 >>
rect 59 252 60 253 
<< m1 >>
rect 60 252 61 253 
<< m2 >>
rect 60 252 61 253 
<< m1 >>
rect 64 252 65 253 
<< m1 >>
rect 73 252 74 253 
<< m2 >>
rect 74 252 75 253 
<< m1 >>
rect 100 252 101 253 
<< m1 >>
rect 116 252 117 253 
<< m1 >>
rect 118 252 119 253 
<< m1 >>
rect 121 252 122 253 
<< m1 >>
rect 128 252 129 253 
<< m1 >>
rect 130 252 131 253 
<< m1 >>
rect 132 252 133 253 
<< m1 >>
rect 134 252 135 253 
<< m1 >>
rect 136 252 137 253 
<< m1 >>
rect 142 252 143 253 
<< m1 >>
rect 145 252 146 253 
<< m2 >>
rect 145 252 146 253 
<< m1 >>
rect 154 252 155 253 
<< m2 >>
rect 154 252 155 253 
<< m1 >>
rect 163 252 164 253 
<< m1 >>
rect 165 252 166 253 
<< m1 >>
rect 167 252 168 253 
<< m1 >>
rect 171 252 172 253 
<< m1 >>
rect 178 252 179 253 
<< m1 >>
rect 181 252 182 253 
<< m2 >>
rect 181 252 182 253 
<< m2c >>
rect 181 252 182 253 
<< m1 >>
rect 181 252 182 253 
<< m2 >>
rect 181 252 182 253 
<< m1 >>
rect 183 252 184 253 
<< m2 >>
rect 183 252 184 253 
<< m2c >>
rect 183 252 184 253 
<< m1 >>
rect 183 252 184 253 
<< m2 >>
rect 183 252 184 253 
<< m1 >>
rect 186 252 187 253 
<< m2 >>
rect 186 252 187 253 
<< m2c >>
rect 186 252 187 253 
<< m1 >>
rect 186 252 187 253 
<< m2 >>
rect 186 252 187 253 
<< m1 >>
rect 188 252 189 253 
<< m2 >>
rect 188 252 189 253 
<< m2c >>
rect 188 252 189 253 
<< m1 >>
rect 188 252 189 253 
<< m2 >>
rect 188 252 189 253 
<< m1 >>
rect 190 252 191 253 
<< m2 >>
rect 190 252 191 253 
<< m2c >>
rect 190 252 191 253 
<< m1 >>
rect 190 252 191 253 
<< m2 >>
rect 190 252 191 253 
<< m1 >>
rect 199 252 200 253 
<< m1 >>
rect 211 252 212 253 
<< m1 >>
rect 226 252 227 253 
<< m1 >>
rect 232 252 233 253 
<< m1 >>
rect 235 252 236 253 
<< m1 >>
rect 237 252 238 253 
<< m1 >>
rect 239 252 240 253 
<< m1 >>
rect 243 252 244 253 
<< m1 >>
rect 247 252 248 253 
<< m1 >>
rect 262 252 263 253 
<< m1 >>
rect 272 252 273 253 
<< m2 >>
rect 273 252 274 253 
<< m2 >>
rect 279 252 280 253 
<< m1 >>
rect 280 252 281 253 
<< m1 >>
rect 283 252 284 253 
<< m1 >>
rect 286 252 287 253 
<< m1 >>
rect 294 252 295 253 
<< m1 >>
rect 298 252 299 253 
<< m1 >>
rect 327 252 328 253 
<< m1 >>
rect 329 252 330 253 
<< m2 >>
rect 330 252 331 253 
<< m1 >>
rect 10 253 11 254 
<< m1 >>
rect 28 253 29 254 
<< m2 >>
rect 28 253 29 254 
<< m1 >>
rect 37 253 38 254 
<< m2 >>
rect 37 253 38 254 
<< m1 >>
rect 39 253 40 254 
<< m2 >>
rect 43 253 44 254 
<< m1 >>
rect 44 253 45 254 
<< m1 >>
rect 46 253 47 254 
<< m2 >>
rect 46 253 47 254 
<< m1 >>
rect 49 253 50 254 
<< m2 >>
rect 56 253 57 254 
<< m1 >>
rect 60 253 61 254 
<< m2 >>
rect 60 253 61 254 
<< m1 >>
rect 64 253 65 254 
<< m1 >>
rect 71 253 72 254 
<< m2 >>
rect 71 253 72 254 
<< m2c >>
rect 71 253 72 254 
<< m1 >>
rect 71 253 72 254 
<< m2 >>
rect 71 253 72 254 
<< m2 >>
rect 72 253 73 254 
<< m1 >>
rect 73 253 74 254 
<< m2 >>
rect 73 253 74 254 
<< m2 >>
rect 74 253 75 254 
<< m1 >>
rect 100 253 101 254 
<< m1 >>
rect 114 253 115 254 
<< m2 >>
rect 114 253 115 254 
<< m2c >>
rect 114 253 115 254 
<< m1 >>
rect 114 253 115 254 
<< m2 >>
rect 114 253 115 254 
<< m2 >>
rect 115 253 116 254 
<< m1 >>
rect 116 253 117 254 
<< m2 >>
rect 116 253 117 254 
<< m2 >>
rect 117 253 118 254 
<< m1 >>
rect 118 253 119 254 
<< m2 >>
rect 118 253 119 254 
<< m2 >>
rect 119 253 120 254 
<< m1 >>
rect 120 253 121 254 
<< m2 >>
rect 120 253 121 254 
<< m2c >>
rect 120 253 121 254 
<< m1 >>
rect 120 253 121 254 
<< m2 >>
rect 120 253 121 254 
<< m1 >>
rect 121 253 122 254 
<< m1 >>
rect 128 253 129 254 
<< m1 >>
rect 130 253 131 254 
<< m1 >>
rect 132 253 133 254 
<< m1 >>
rect 134 253 135 254 
<< m1 >>
rect 136 253 137 254 
<< m1 >>
rect 142 253 143 254 
<< m1 >>
rect 143 253 144 254 
<< m1 >>
rect 144 253 145 254 
<< m1 >>
rect 145 253 146 254 
<< m2 >>
rect 145 253 146 254 
<< m1 >>
rect 154 253 155 254 
<< m2 >>
rect 154 253 155 254 
<< m1 >>
rect 163 253 164 254 
<< m1 >>
rect 165 253 166 254 
<< m1 >>
rect 167 253 168 254 
<< m1 >>
rect 171 253 172 254 
<< m1 >>
rect 178 253 179 254 
<< m2 >>
rect 181 253 182 254 
<< m2 >>
rect 183 253 184 254 
<< m2 >>
rect 186 253 187 254 
<< m2 >>
rect 188 253 189 254 
<< m2 >>
rect 190 253 191 254 
<< m1 >>
rect 199 253 200 254 
<< m1 >>
rect 200 253 201 254 
<< m1 >>
rect 201 253 202 254 
<< m1 >>
rect 202 253 203 254 
<< m1 >>
rect 203 253 204 254 
<< m1 >>
rect 204 253 205 254 
<< m1 >>
rect 205 253 206 254 
<< m1 >>
rect 206 253 207 254 
<< m1 >>
rect 207 253 208 254 
<< m1 >>
rect 208 253 209 254 
<< m1 >>
rect 209 253 210 254 
<< m1 >>
rect 210 253 211 254 
<< m1 >>
rect 211 253 212 254 
<< m1 >>
rect 226 253 227 254 
<< m1 >>
rect 232 253 233 254 
<< m1 >>
rect 235 253 236 254 
<< m1 >>
rect 237 253 238 254 
<< m1 >>
rect 239 253 240 254 
<< m1 >>
rect 243 253 244 254 
<< m1 >>
rect 247 253 248 254 
<< m1 >>
rect 262 253 263 254 
<< m1 >>
rect 272 253 273 254 
<< m2 >>
rect 273 253 274 254 
<< m2 >>
rect 279 253 280 254 
<< m1 >>
rect 280 253 281 254 
<< m1 >>
rect 281 253 282 254 
<< m1 >>
rect 282 253 283 254 
<< m1 >>
rect 283 253 284 254 
<< m1 >>
rect 286 253 287 254 
<< m1 >>
rect 294 253 295 254 
<< m1 >>
rect 298 253 299 254 
<< m1 >>
rect 327 253 328 254 
<< m1 >>
rect 329 253 330 254 
<< m2 >>
rect 330 253 331 254 
<< m1 >>
rect 10 254 11 255 
<< m1 >>
rect 28 254 29 255 
<< m2 >>
rect 28 254 29 255 
<< m1 >>
rect 37 254 38 255 
<< m2 >>
rect 37 254 38 255 
<< m1 >>
rect 39 254 40 255 
<< m2 >>
rect 43 254 44 255 
<< m1 >>
rect 44 254 45 255 
<< m1 >>
rect 46 254 47 255 
<< m2 >>
rect 46 254 47 255 
<< m1 >>
rect 49 254 50 255 
<< m1 >>
rect 50 254 51 255 
<< m1 >>
rect 51 254 52 255 
<< m1 >>
rect 52 254 53 255 
<< m1 >>
rect 53 254 54 255 
<< m1 >>
rect 54 254 55 255 
<< m1 >>
rect 55 254 56 255 
<< m1 >>
rect 56 254 57 255 
<< m2 >>
rect 56 254 57 255 
<< m1 >>
rect 57 254 58 255 
<< m1 >>
rect 58 254 59 255 
<< m1 >>
rect 59 254 60 255 
<< m1 >>
rect 60 254 61 255 
<< m2 >>
rect 60 254 61 255 
<< m1 >>
rect 64 254 65 255 
<< m1 >>
rect 71 254 72 255 
<< m1 >>
rect 73 254 74 255 
<< m1 >>
rect 100 254 101 255 
<< m1 >>
rect 101 254 102 255 
<< m1 >>
rect 102 254 103 255 
<< m2 >>
rect 102 254 103 255 
<< m2c >>
rect 102 254 103 255 
<< m1 >>
rect 102 254 103 255 
<< m2 >>
rect 102 254 103 255 
<< m1 >>
rect 114 254 115 255 
<< m1 >>
rect 116 254 117 255 
<< m1 >>
rect 118 254 119 255 
<< m1 >>
rect 128 254 129 255 
<< m1 >>
rect 130 254 131 255 
<< m1 >>
rect 132 254 133 255 
<< m1 >>
rect 134 254 135 255 
<< m1 >>
rect 136 254 137 255 
<< m2 >>
rect 145 254 146 255 
<< m1 >>
rect 154 254 155 255 
<< m2 >>
rect 154 254 155 255 
<< m1 >>
rect 163 254 164 255 
<< m1 >>
rect 165 254 166 255 
<< m1 >>
rect 167 254 168 255 
<< m1 >>
rect 171 254 172 255 
<< m2 >>
rect 171 254 172 255 
<< m2c >>
rect 171 254 172 255 
<< m1 >>
rect 171 254 172 255 
<< m2 >>
rect 171 254 172 255 
<< m1 >>
rect 178 254 179 255 
<< m1 >>
rect 179 254 180 255 
<< m1 >>
rect 180 254 181 255 
<< m1 >>
rect 181 254 182 255 
<< m2 >>
rect 181 254 182 255 
<< m1 >>
rect 182 254 183 255 
<< m1 >>
rect 183 254 184 255 
<< m2 >>
rect 183 254 184 255 
<< m1 >>
rect 184 254 185 255 
<< m1 >>
rect 185 254 186 255 
<< m1 >>
rect 186 254 187 255 
<< m2 >>
rect 186 254 187 255 
<< m1 >>
rect 187 254 188 255 
<< m1 >>
rect 188 254 189 255 
<< m2 >>
rect 188 254 189 255 
<< m1 >>
rect 189 254 190 255 
<< m1 >>
rect 190 254 191 255 
<< m2 >>
rect 190 254 191 255 
<< m1 >>
rect 191 254 192 255 
<< m1 >>
rect 192 254 193 255 
<< m2 >>
rect 192 254 193 255 
<< m2c >>
rect 192 254 193 255 
<< m1 >>
rect 192 254 193 255 
<< m2 >>
rect 192 254 193 255 
<< m1 >>
rect 226 254 227 255 
<< m1 >>
rect 227 254 228 255 
<< m1 >>
rect 228 254 229 255 
<< m2 >>
rect 228 254 229 255 
<< m2c >>
rect 228 254 229 255 
<< m1 >>
rect 228 254 229 255 
<< m2 >>
rect 228 254 229 255 
<< m1 >>
rect 232 254 233 255 
<< m1 >>
rect 235 254 236 255 
<< m1 >>
rect 237 254 238 255 
<< m1 >>
rect 239 254 240 255 
<< m1 >>
rect 243 254 244 255 
<< m1 >>
rect 247 254 248 255 
<< m1 >>
rect 248 254 249 255 
<< m1 >>
rect 249 254 250 255 
<< m1 >>
rect 250 254 251 255 
<< m1 >>
rect 251 254 252 255 
<< m1 >>
rect 252 254 253 255 
<< m1 >>
rect 253 254 254 255 
<< m1 >>
rect 262 254 263 255 
<< m1 >>
rect 272 254 273 255 
<< m2 >>
rect 273 254 274 255 
<< m2 >>
rect 279 254 280 255 
<< m1 >>
rect 286 254 287 255 
<< m1 >>
rect 294 254 295 255 
<< m1 >>
rect 298 254 299 255 
<< m1 >>
rect 327 254 328 255 
<< m1 >>
rect 329 254 330 255 
<< m2 >>
rect 330 254 331 255 
<< m1 >>
rect 10 255 11 256 
<< m1 >>
rect 28 255 29 256 
<< m2 >>
rect 28 255 29 256 
<< m1 >>
rect 37 255 38 256 
<< m2 >>
rect 37 255 38 256 
<< m1 >>
rect 39 255 40 256 
<< m2 >>
rect 43 255 44 256 
<< m1 >>
rect 44 255 45 256 
<< m1 >>
rect 46 255 47 256 
<< m2 >>
rect 46 255 47 256 
<< m2 >>
rect 56 255 57 256 
<< m2 >>
rect 57 255 58 256 
<< m2 >>
rect 60 255 61 256 
<< m1 >>
rect 64 255 65 256 
<< m1 >>
rect 71 255 72 256 
<< m1 >>
rect 73 255 74 256 
<< m2 >>
rect 102 255 103 256 
<< m1 >>
rect 114 255 115 256 
<< m1 >>
rect 116 255 117 256 
<< m1 >>
rect 118 255 119 256 
<< m1 >>
rect 128 255 129 256 
<< m1 >>
rect 130 255 131 256 
<< m1 >>
rect 132 255 133 256 
<< m1 >>
rect 134 255 135 256 
<< m1 >>
rect 136 255 137 256 
<< m2 >>
rect 145 255 146 256 
<< m1 >>
rect 154 255 155 256 
<< m2 >>
rect 154 255 155 256 
<< m1 >>
rect 163 255 164 256 
<< m1 >>
rect 165 255 166 256 
<< m1 >>
rect 167 255 168 256 
<< m2 >>
rect 171 255 172 256 
<< m2 >>
rect 181 255 182 256 
<< m2 >>
rect 183 255 184 256 
<< m2 >>
rect 186 255 187 256 
<< m2 >>
rect 188 255 189 256 
<< m2 >>
rect 190 255 191 256 
<< m2 >>
rect 192 255 193 256 
<< m2 >>
rect 228 255 229 256 
<< m1 >>
rect 232 255 233 256 
<< m1 >>
rect 235 255 236 256 
<< m1 >>
rect 237 255 238 256 
<< m1 >>
rect 239 255 240 256 
<< m1 >>
rect 243 255 244 256 
<< m1 >>
rect 253 255 254 256 
<< m1 >>
rect 262 255 263 256 
<< m1 >>
rect 272 255 273 256 
<< m2 >>
rect 273 255 274 256 
<< m1 >>
rect 279 255 280 256 
<< m2 >>
rect 279 255 280 256 
<< m2c >>
rect 279 255 280 256 
<< m1 >>
rect 279 255 280 256 
<< m2 >>
rect 279 255 280 256 
<< m1 >>
rect 286 255 287 256 
<< m1 >>
rect 294 255 295 256 
<< m2 >>
rect 294 255 295 256 
<< m2c >>
rect 294 255 295 256 
<< m1 >>
rect 294 255 295 256 
<< m2 >>
rect 294 255 295 256 
<< m1 >>
rect 298 255 299 256 
<< m1 >>
rect 327 255 328 256 
<< m1 >>
rect 329 255 330 256 
<< m2 >>
rect 330 255 331 256 
<< m1 >>
rect 10 256 11 257 
<< m1 >>
rect 28 256 29 257 
<< m2 >>
rect 28 256 29 257 
<< m1 >>
rect 37 256 38 257 
<< m2 >>
rect 37 256 38 257 
<< m1 >>
rect 39 256 40 257 
<< m2 >>
rect 43 256 44 257 
<< m1 >>
rect 44 256 45 257 
<< m1 >>
rect 46 256 47 257 
<< m2 >>
rect 46 256 47 257 
<< m2 >>
rect 47 256 48 257 
<< m1 >>
rect 48 256 49 257 
<< m2 >>
rect 48 256 49 257 
<< m2c >>
rect 48 256 49 257 
<< m1 >>
rect 48 256 49 257 
<< m2 >>
rect 48 256 49 257 
<< m1 >>
rect 57 256 58 257 
<< m2 >>
rect 57 256 58 257 
<< m2c >>
rect 57 256 58 257 
<< m1 >>
rect 57 256 58 257 
<< m2 >>
rect 57 256 58 257 
<< m1 >>
rect 60 256 61 257 
<< m2 >>
rect 60 256 61 257 
<< m2c >>
rect 60 256 61 257 
<< m1 >>
rect 60 256 61 257 
<< m2 >>
rect 60 256 61 257 
<< m1 >>
rect 62 256 63 257 
<< m2 >>
rect 62 256 63 257 
<< m2c >>
rect 62 256 63 257 
<< m1 >>
rect 62 256 63 257 
<< m2 >>
rect 62 256 63 257 
<< m2 >>
rect 63 256 64 257 
<< m1 >>
rect 64 256 65 257 
<< m2 >>
rect 64 256 65 257 
<< m2 >>
rect 65 256 66 257 
<< m1 >>
rect 66 256 67 257 
<< m2 >>
rect 66 256 67 257 
<< m2c >>
rect 66 256 67 257 
<< m1 >>
rect 66 256 67 257 
<< m2 >>
rect 66 256 67 257 
<< m1 >>
rect 67 256 68 257 
<< m1 >>
rect 68 256 69 257 
<< m1 >>
rect 69 256 70 257 
<< m1 >>
rect 70 256 71 257 
<< m1 >>
rect 71 256 72 257 
<< m1 >>
rect 73 256 74 257 
<< m2 >>
rect 74 256 75 257 
<< m1 >>
rect 75 256 76 257 
<< m2 >>
rect 75 256 76 257 
<< m2c >>
rect 75 256 76 257 
<< m1 >>
rect 75 256 76 257 
<< m2 >>
rect 75 256 76 257 
<< m1 >>
rect 76 256 77 257 
<< m1 >>
rect 77 256 78 257 
<< m1 >>
rect 78 256 79 257 
<< m1 >>
rect 79 256 80 257 
<< m1 >>
rect 80 256 81 257 
<< m1 >>
rect 81 256 82 257 
<< m1 >>
rect 82 256 83 257 
<< m1 >>
rect 83 256 84 257 
<< m1 >>
rect 84 256 85 257 
<< m1 >>
rect 85 256 86 257 
<< m1 >>
rect 86 256 87 257 
<< m1 >>
rect 87 256 88 257 
<< m1 >>
rect 88 256 89 257 
<< m1 >>
rect 89 256 90 257 
<< m1 >>
rect 90 256 91 257 
<< m1 >>
rect 91 256 92 257 
<< m1 >>
rect 92 256 93 257 
<< m1 >>
rect 93 256 94 257 
<< m1 >>
rect 94 256 95 257 
<< m1 >>
rect 95 256 96 257 
<< m1 >>
rect 96 256 97 257 
<< m1 >>
rect 97 256 98 257 
<< m1 >>
rect 98 256 99 257 
<< m1 >>
rect 99 256 100 257 
<< m1 >>
rect 100 256 101 257 
<< m1 >>
rect 101 256 102 257 
<< m1 >>
rect 102 256 103 257 
<< m2 >>
rect 102 256 103 257 
<< m1 >>
rect 103 256 104 257 
<< m1 >>
rect 104 256 105 257 
<< m1 >>
rect 105 256 106 257 
<< m1 >>
rect 106 256 107 257 
<< m1 >>
rect 107 256 108 257 
<< m1 >>
rect 108 256 109 257 
<< m1 >>
rect 109 256 110 257 
<< m1 >>
rect 110 256 111 257 
<< m1 >>
rect 111 256 112 257 
<< m1 >>
rect 112 256 113 257 
<< m1 >>
rect 113 256 114 257 
<< m1 >>
rect 114 256 115 257 
<< m1 >>
rect 116 256 117 257 
<< m1 >>
rect 118 256 119 257 
<< m1 >>
rect 128 256 129 257 
<< m2 >>
rect 128 256 129 257 
<< m2c >>
rect 128 256 129 257 
<< m1 >>
rect 128 256 129 257 
<< m2 >>
rect 128 256 129 257 
<< m2 >>
rect 129 256 130 257 
<< m1 >>
rect 130 256 131 257 
<< m2 >>
rect 130 256 131 257 
<< m2 >>
rect 131 256 132 257 
<< m1 >>
rect 132 256 133 257 
<< m2 >>
rect 132 256 133 257 
<< m2 >>
rect 133 256 134 257 
<< m1 >>
rect 134 256 135 257 
<< m2 >>
rect 134 256 135 257 
<< m2 >>
rect 135 256 136 257 
<< m1 >>
rect 136 256 137 257 
<< m2 >>
rect 136 256 137 257 
<< m2 >>
rect 137 256 138 257 
<< m1 >>
rect 138 256 139 257 
<< m2 >>
rect 138 256 139 257 
<< m2c >>
rect 138 256 139 257 
<< m1 >>
rect 138 256 139 257 
<< m2 >>
rect 138 256 139 257 
<< m1 >>
rect 139 256 140 257 
<< m1 >>
rect 140 256 141 257 
<< m1 >>
rect 141 256 142 257 
<< m1 >>
rect 142 256 143 257 
<< m1 >>
rect 143 256 144 257 
<< m1 >>
rect 144 256 145 257 
<< m1 >>
rect 145 256 146 257 
<< m2 >>
rect 145 256 146 257 
<< m1 >>
rect 146 256 147 257 
<< m1 >>
rect 147 256 148 257 
<< m1 >>
rect 148 256 149 257 
<< m1 >>
rect 149 256 150 257 
<< m1 >>
rect 150 256 151 257 
<< m1 >>
rect 151 256 152 257 
<< m1 >>
rect 152 256 153 257 
<< m1 >>
rect 153 256 154 257 
<< m1 >>
rect 154 256 155 257 
<< m2 >>
rect 154 256 155 257 
<< m1 >>
rect 163 256 164 257 
<< m1 >>
rect 165 256 166 257 
<< m1 >>
rect 167 256 168 257 
<< m1 >>
rect 168 256 169 257 
<< m1 >>
rect 169 256 170 257 
<< m1 >>
rect 170 256 171 257 
<< m1 >>
rect 171 256 172 257 
<< m2 >>
rect 171 256 172 257 
<< m1 >>
rect 172 256 173 257 
<< m1 >>
rect 173 256 174 257 
<< m1 >>
rect 174 256 175 257 
<< m1 >>
rect 175 256 176 257 
<< m1 >>
rect 176 256 177 257 
<< m1 >>
rect 177 256 178 257 
<< m1 >>
rect 178 256 179 257 
<< m1 >>
rect 179 256 180 257 
<< m1 >>
rect 180 256 181 257 
<< m1 >>
rect 181 256 182 257 
<< m2 >>
rect 181 256 182 257 
<< m1 >>
rect 182 256 183 257 
<< m1 >>
rect 183 256 184 257 
<< m2 >>
rect 183 256 184 257 
<< m1 >>
rect 184 256 185 257 
<< m1 >>
rect 185 256 186 257 
<< m1 >>
rect 186 256 187 257 
<< m2 >>
rect 186 256 187 257 
<< m1 >>
rect 187 256 188 257 
<< m1 >>
rect 188 256 189 257 
<< m2 >>
rect 188 256 189 257 
<< m1 >>
rect 189 256 190 257 
<< m1 >>
rect 190 256 191 257 
<< m2 >>
rect 190 256 191 257 
<< m1 >>
rect 191 256 192 257 
<< m1 >>
rect 192 256 193 257 
<< m2 >>
rect 192 256 193 257 
<< m1 >>
rect 193 256 194 257 
<< m1 >>
rect 194 256 195 257 
<< m1 >>
rect 195 256 196 257 
<< m1 >>
rect 196 256 197 257 
<< m1 >>
rect 197 256 198 257 
<< m1 >>
rect 198 256 199 257 
<< m1 >>
rect 199 256 200 257 
<< m1 >>
rect 200 256 201 257 
<< m1 >>
rect 201 256 202 257 
<< m1 >>
rect 202 256 203 257 
<< m1 >>
rect 203 256 204 257 
<< m1 >>
rect 204 256 205 257 
<< m1 >>
rect 205 256 206 257 
<< m1 >>
rect 206 256 207 257 
<< m1 >>
rect 207 256 208 257 
<< m1 >>
rect 208 256 209 257 
<< m1 >>
rect 209 256 210 257 
<< m1 >>
rect 210 256 211 257 
<< m1 >>
rect 211 256 212 257 
<< m1 >>
rect 212 256 213 257 
<< m1 >>
rect 213 256 214 257 
<< m1 >>
rect 214 256 215 257 
<< m1 >>
rect 215 256 216 257 
<< m1 >>
rect 216 256 217 257 
<< m1 >>
rect 217 256 218 257 
<< m1 >>
rect 218 256 219 257 
<< m1 >>
rect 219 256 220 257 
<< m1 >>
rect 220 256 221 257 
<< m1 >>
rect 221 256 222 257 
<< m1 >>
rect 222 256 223 257 
<< m1 >>
rect 223 256 224 257 
<< m1 >>
rect 224 256 225 257 
<< m1 >>
rect 225 256 226 257 
<< m1 >>
rect 226 256 227 257 
<< m1 >>
rect 227 256 228 257 
<< m1 >>
rect 228 256 229 257 
<< m2 >>
rect 228 256 229 257 
<< m1 >>
rect 229 256 230 257 
<< m1 >>
rect 230 256 231 257 
<< m1 >>
rect 231 256 232 257 
<< m1 >>
rect 232 256 233 257 
<< m1 >>
rect 235 256 236 257 
<< m1 >>
rect 237 256 238 257 
<< m1 >>
rect 239 256 240 257 
<< m1 >>
rect 243 256 244 257 
<< m1 >>
rect 253 256 254 257 
<< m1 >>
rect 262 256 263 257 
<< m1 >>
rect 272 256 273 257 
<< m2 >>
rect 273 256 274 257 
<< m1 >>
rect 279 256 280 257 
<< m1 >>
rect 286 256 287 257 
<< m2 >>
rect 294 256 295 257 
<< m1 >>
rect 298 256 299 257 
<< m2 >>
rect 323 256 324 257 
<< m2 >>
rect 324 256 325 257 
<< m2 >>
rect 325 256 326 257 
<< m2 >>
rect 326 256 327 257 
<< m1 >>
rect 327 256 328 257 
<< m2 >>
rect 327 256 328 257 
<< m2 >>
rect 328 256 329 257 
<< m1 >>
rect 329 256 330 257 
<< m2 >>
rect 329 256 330 257 
<< m2 >>
rect 330 256 331 257 
<< m1 >>
rect 10 257 11 258 
<< m1 >>
rect 28 257 29 258 
<< m2 >>
rect 28 257 29 258 
<< m1 >>
rect 37 257 38 258 
<< m2 >>
rect 37 257 38 258 
<< m1 >>
rect 39 257 40 258 
<< m2 >>
rect 43 257 44 258 
<< m1 >>
rect 44 257 45 258 
<< m1 >>
rect 46 257 47 258 
<< m1 >>
rect 48 257 49 258 
<< m1 >>
rect 57 257 58 258 
<< m1 >>
rect 60 257 61 258 
<< m1 >>
rect 62 257 63 258 
<< m1 >>
rect 64 257 65 258 
<< m1 >>
rect 73 257 74 258 
<< m2 >>
rect 74 257 75 258 
<< m2 >>
rect 102 257 103 258 
<< m2 >>
rect 103 257 104 258 
<< m2 >>
rect 104 257 105 258 
<< m2 >>
rect 105 257 106 258 
<< m2 >>
rect 106 257 107 258 
<< m2 >>
rect 107 257 108 258 
<< m2 >>
rect 108 257 109 258 
<< m2 >>
rect 109 257 110 258 
<< m2 >>
rect 110 257 111 258 
<< m2 >>
rect 111 257 112 258 
<< m2 >>
rect 112 257 113 258 
<< m2 >>
rect 113 257 114 258 
<< m2 >>
rect 114 257 115 258 
<< m2 >>
rect 115 257 116 258 
<< m1 >>
rect 116 257 117 258 
<< m2 >>
rect 116 257 117 258 
<< m2 >>
rect 117 257 118 258 
<< m1 >>
rect 118 257 119 258 
<< m2 >>
rect 118 257 119 258 
<< m1 >>
rect 130 257 131 258 
<< m1 >>
rect 132 257 133 258 
<< m1 >>
rect 134 257 135 258 
<< m1 >>
rect 136 257 137 258 
<< m2 >>
rect 145 257 146 258 
<< m2 >>
rect 154 257 155 258 
<< m1 >>
rect 163 257 164 258 
<< m1 >>
rect 165 257 166 258 
<< m2 >>
rect 171 257 172 258 
<< m2 >>
rect 181 257 182 258 
<< m2 >>
rect 183 257 184 258 
<< m2 >>
rect 186 257 187 258 
<< m2 >>
rect 188 257 189 258 
<< m2 >>
rect 190 257 191 258 
<< m2 >>
rect 192 257 193 258 
<< m2 >>
rect 193 257 194 258 
<< m2 >>
rect 194 257 195 258 
<< m2 >>
rect 195 257 196 258 
<< m2 >>
rect 196 257 197 258 
<< m2 >>
rect 197 257 198 258 
<< m2 >>
rect 198 257 199 258 
<< m2 >>
rect 199 257 200 258 
<< m2 >>
rect 200 257 201 258 
<< m2 >>
rect 201 257 202 258 
<< m2 >>
rect 202 257 203 258 
<< m2 >>
rect 203 257 204 258 
<< m2 >>
rect 204 257 205 258 
<< m2 >>
rect 205 257 206 258 
<< m2 >>
rect 206 257 207 258 
<< m2 >>
rect 207 257 208 258 
<< m2 >>
rect 208 257 209 258 
<< m2 >>
rect 209 257 210 258 
<< m2 >>
rect 210 257 211 258 
<< m2 >>
rect 211 257 212 258 
<< m2 >>
rect 212 257 213 258 
<< m2 >>
rect 213 257 214 258 
<< m2 >>
rect 214 257 215 258 
<< m2 >>
rect 215 257 216 258 
<< m2 >>
rect 216 257 217 258 
<< m2 >>
rect 217 257 218 258 
<< m2 >>
rect 218 257 219 258 
<< m2 >>
rect 219 257 220 258 
<< m2 >>
rect 220 257 221 258 
<< m2 >>
rect 221 257 222 258 
<< m2 >>
rect 222 257 223 258 
<< m2 >>
rect 223 257 224 258 
<< m2 >>
rect 224 257 225 258 
<< m2 >>
rect 225 257 226 258 
<< m2 >>
rect 226 257 227 258 
<< m2 >>
rect 228 257 229 258 
<< m1 >>
rect 235 257 236 258 
<< m1 >>
rect 237 257 238 258 
<< m1 >>
rect 239 257 240 258 
<< m2 >>
rect 239 257 240 258 
<< m2 >>
rect 240 257 241 258 
<< m1 >>
rect 241 257 242 258 
<< m2 >>
rect 241 257 242 258 
<< m2c >>
rect 241 257 242 258 
<< m1 >>
rect 241 257 242 258 
<< m2 >>
rect 241 257 242 258 
<< m2 >>
rect 242 257 243 258 
<< m1 >>
rect 243 257 244 258 
<< m2 >>
rect 243 257 244 258 
<< m2 >>
rect 244 257 245 258 
<< m1 >>
rect 245 257 246 258 
<< m2 >>
rect 245 257 246 258 
<< m2c >>
rect 245 257 246 258 
<< m1 >>
rect 245 257 246 258 
<< m2 >>
rect 245 257 246 258 
<< m1 >>
rect 246 257 247 258 
<< m1 >>
rect 247 257 248 258 
<< m1 >>
rect 248 257 249 258 
<< m1 >>
rect 249 257 250 258 
<< m1 >>
rect 250 257 251 258 
<< m1 >>
rect 251 257 252 258 
<< m2 >>
rect 251 257 252 258 
<< m2c >>
rect 251 257 252 258 
<< m1 >>
rect 251 257 252 258 
<< m2 >>
rect 251 257 252 258 
<< m2 >>
rect 252 257 253 258 
<< m1 >>
rect 253 257 254 258 
<< m2 >>
rect 253 257 254 258 
<< m2 >>
rect 254 257 255 258 
<< m1 >>
rect 262 257 263 258 
<< m1 >>
rect 272 257 273 258 
<< m2 >>
rect 273 257 274 258 
<< m1 >>
rect 276 257 277 258 
<< m2 >>
rect 276 257 277 258 
<< m2c >>
rect 276 257 277 258 
<< m1 >>
rect 276 257 277 258 
<< m2 >>
rect 276 257 277 258 
<< m1 >>
rect 277 257 278 258 
<< m1 >>
rect 278 257 279 258 
<< m1 >>
rect 279 257 280 258 
<< m1 >>
rect 286 257 287 258 
<< m1 >>
rect 287 257 288 258 
<< m1 >>
rect 288 257 289 258 
<< m1 >>
rect 289 257 290 258 
<< m1 >>
rect 290 257 291 258 
<< m1 >>
rect 291 257 292 258 
<< m1 >>
rect 292 257 293 258 
<< m1 >>
rect 293 257 294 258 
<< m1 >>
rect 294 257 295 258 
<< m2 >>
rect 294 257 295 258 
<< m1 >>
rect 295 257 296 258 
<< m1 >>
rect 296 257 297 258 
<< m2 >>
rect 296 257 297 258 
<< m2c >>
rect 296 257 297 258 
<< m1 >>
rect 296 257 297 258 
<< m2 >>
rect 296 257 297 258 
<< m2 >>
rect 297 257 298 258 
<< m1 >>
rect 298 257 299 258 
<< m2 >>
rect 298 257 299 258 
<< m1 >>
rect 299 257 300 258 
<< m2 >>
rect 299 257 300 258 
<< m1 >>
rect 300 257 301 258 
<< m2 >>
rect 300 257 301 258 
<< m1 >>
rect 301 257 302 258 
<< m2 >>
rect 301 257 302 258 
<< m1 >>
rect 302 257 303 258 
<< m2 >>
rect 302 257 303 258 
<< m1 >>
rect 303 257 304 258 
<< m2 >>
rect 303 257 304 258 
<< m1 >>
rect 304 257 305 258 
<< m2 >>
rect 304 257 305 258 
<< m1 >>
rect 305 257 306 258 
<< m2 >>
rect 305 257 306 258 
<< m1 >>
rect 306 257 307 258 
<< m2 >>
rect 306 257 307 258 
<< m1 >>
rect 307 257 308 258 
<< m2 >>
rect 307 257 308 258 
<< m1 >>
rect 308 257 309 258 
<< m2 >>
rect 308 257 309 258 
<< m1 >>
rect 309 257 310 258 
<< m2 >>
rect 309 257 310 258 
<< m1 >>
rect 310 257 311 258 
<< m2 >>
rect 310 257 311 258 
<< m1 >>
rect 311 257 312 258 
<< m2 >>
rect 311 257 312 258 
<< m1 >>
rect 312 257 313 258 
<< m2 >>
rect 312 257 313 258 
<< m1 >>
rect 313 257 314 258 
<< m2 >>
rect 313 257 314 258 
<< m1 >>
rect 314 257 315 258 
<< m2 >>
rect 314 257 315 258 
<< m1 >>
rect 315 257 316 258 
<< m2 >>
rect 315 257 316 258 
<< m1 >>
rect 316 257 317 258 
<< m2 >>
rect 316 257 317 258 
<< m1 >>
rect 317 257 318 258 
<< m1 >>
rect 318 257 319 258 
<< m1 >>
rect 319 257 320 258 
<< m1 >>
rect 320 257 321 258 
<< m1 >>
rect 321 257 322 258 
<< m1 >>
rect 322 257 323 258 
<< m1 >>
rect 323 257 324 258 
<< m2 >>
rect 323 257 324 258 
<< m1 >>
rect 324 257 325 258 
<< m1 >>
rect 325 257 326 258 
<< m1 >>
rect 327 257 328 258 
<< m1 >>
rect 329 257 330 258 
<< m1 >>
rect 10 258 11 259 
<< m1 >>
rect 28 258 29 259 
<< m2 >>
rect 28 258 29 259 
<< m1 >>
rect 37 258 38 259 
<< m2 >>
rect 37 258 38 259 
<< m1 >>
rect 39 258 40 259 
<< m2 >>
rect 43 258 44 259 
<< m1 >>
rect 44 258 45 259 
<< m1 >>
rect 46 258 47 259 
<< m1 >>
rect 48 258 49 259 
<< m1 >>
rect 49 258 50 259 
<< m1 >>
rect 50 258 51 259 
<< m1 >>
rect 51 258 52 259 
<< m1 >>
rect 52 258 53 259 
<< m1 >>
rect 53 258 54 259 
<< m1 >>
rect 54 258 55 259 
<< m1 >>
rect 55 258 56 259 
<< m2 >>
rect 55 258 56 259 
<< m2c >>
rect 55 258 56 259 
<< m1 >>
rect 55 258 56 259 
<< m2 >>
rect 55 258 56 259 
<< m2 >>
rect 56 258 57 259 
<< m1 >>
rect 57 258 58 259 
<< m2 >>
rect 57 258 58 259 
<< m2 >>
rect 58 258 59 259 
<< m2 >>
rect 59 258 60 259 
<< m1 >>
rect 60 258 61 259 
<< m2 >>
rect 60 258 61 259 
<< m2 >>
rect 61 258 62 259 
<< m1 >>
rect 62 258 63 259 
<< m2 >>
rect 62 258 63 259 
<< m2 >>
rect 63 258 64 259 
<< m1 >>
rect 64 258 65 259 
<< m2 >>
rect 64 258 65 259 
<< m2 >>
rect 65 258 66 259 
<< m1 >>
rect 66 258 67 259 
<< m2 >>
rect 66 258 67 259 
<< m2c >>
rect 66 258 67 259 
<< m1 >>
rect 66 258 67 259 
<< m2 >>
rect 66 258 67 259 
<< m1 >>
rect 67 258 68 259 
<< m1 >>
rect 68 258 69 259 
<< m1 >>
rect 69 258 70 259 
<< m1 >>
rect 70 258 71 259 
<< m1 >>
rect 73 258 74 259 
<< m2 >>
rect 74 258 75 259 
<< m1 >>
rect 116 258 117 259 
<< m1 >>
rect 118 258 119 259 
<< m2 >>
rect 118 258 119 259 
<< m1 >>
rect 119 258 120 259 
<< m1 >>
rect 120 258 121 259 
<< m1 >>
rect 121 258 122 259 
<< m1 >>
rect 122 258 123 259 
<< m1 >>
rect 123 258 124 259 
<< m1 >>
rect 124 258 125 259 
<< m1 >>
rect 125 258 126 259 
<< m1 >>
rect 126 258 127 259 
<< m1 >>
rect 127 258 128 259 
<< m1 >>
rect 128 258 129 259 
<< m2 >>
rect 128 258 129 259 
<< m2c >>
rect 128 258 129 259 
<< m1 >>
rect 128 258 129 259 
<< m2 >>
rect 128 258 129 259 
<< m2 >>
rect 129 258 130 259 
<< m1 >>
rect 130 258 131 259 
<< m2 >>
rect 130 258 131 259 
<< m2 >>
rect 131 258 132 259 
<< m1 >>
rect 132 258 133 259 
<< m2 >>
rect 132 258 133 259 
<< m2 >>
rect 133 258 134 259 
<< m1 >>
rect 134 258 135 259 
<< m2 >>
rect 134 258 135 259 
<< m2 >>
rect 135 258 136 259 
<< m1 >>
rect 136 258 137 259 
<< m2 >>
rect 136 258 137 259 
<< m2 >>
rect 137 258 138 259 
<< m1 >>
rect 138 258 139 259 
<< m2 >>
rect 138 258 139 259 
<< m2c >>
rect 138 258 139 259 
<< m1 >>
rect 138 258 139 259 
<< m2 >>
rect 138 258 139 259 
<< m1 >>
rect 139 258 140 259 
<< m1 >>
rect 140 258 141 259 
<< m2 >>
rect 140 258 141 259 
<< m2c >>
rect 140 258 141 259 
<< m1 >>
rect 140 258 141 259 
<< m2 >>
rect 140 258 141 259 
<< m2 >>
rect 141 258 142 259 
<< m1 >>
rect 142 258 143 259 
<< m2 >>
rect 142 258 143 259 
<< m1 >>
rect 143 258 144 259 
<< m2 >>
rect 143 258 144 259 
<< m1 >>
rect 144 258 145 259 
<< m2 >>
rect 144 258 145 259 
<< m1 >>
rect 145 258 146 259 
<< m2 >>
rect 145 258 146 259 
<< m1 >>
rect 146 258 147 259 
<< m1 >>
rect 147 258 148 259 
<< m1 >>
rect 148 258 149 259 
<< m1 >>
rect 149 258 150 259 
<< m1 >>
rect 150 258 151 259 
<< m1 >>
rect 151 258 152 259 
<< m1 >>
rect 152 258 153 259 
<< m1 >>
rect 153 258 154 259 
<< m1 >>
rect 154 258 155 259 
<< m2 >>
rect 154 258 155 259 
<< m1 >>
rect 155 258 156 259 
<< m1 >>
rect 156 258 157 259 
<< m1 >>
rect 157 258 158 259 
<< m1 >>
rect 158 258 159 259 
<< m1 >>
rect 159 258 160 259 
<< m1 >>
rect 160 258 161 259 
<< m1 >>
rect 161 258 162 259 
<< m1 >>
rect 162 258 163 259 
<< m1 >>
rect 163 258 164 259 
<< m1 >>
rect 165 258 166 259 
<< m1 >>
rect 171 258 172 259 
<< m2 >>
rect 171 258 172 259 
<< m2c >>
rect 171 258 172 259 
<< m1 >>
rect 171 258 172 259 
<< m2 >>
rect 171 258 172 259 
<< m1 >>
rect 181 258 182 259 
<< m2 >>
rect 181 258 182 259 
<< m2c >>
rect 181 258 182 259 
<< m1 >>
rect 181 258 182 259 
<< m2 >>
rect 181 258 182 259 
<< m1 >>
rect 183 258 184 259 
<< m2 >>
rect 183 258 184 259 
<< m2c >>
rect 183 258 184 259 
<< m1 >>
rect 183 258 184 259 
<< m2 >>
rect 183 258 184 259 
<< m1 >>
rect 186 258 187 259 
<< m2 >>
rect 186 258 187 259 
<< m2c >>
rect 186 258 187 259 
<< m1 >>
rect 186 258 187 259 
<< m2 >>
rect 186 258 187 259 
<< m1 >>
rect 188 258 189 259 
<< m2 >>
rect 188 258 189 259 
<< m2c >>
rect 188 258 189 259 
<< m1 >>
rect 188 258 189 259 
<< m2 >>
rect 188 258 189 259 
<< m1 >>
rect 190 258 191 259 
<< m2 >>
rect 190 258 191 259 
<< m2c >>
rect 190 258 191 259 
<< m1 >>
rect 190 258 191 259 
<< m2 >>
rect 190 258 191 259 
<< m1 >>
rect 226 258 227 259 
<< m2 >>
rect 226 258 227 259 
<< m2c >>
rect 226 258 227 259 
<< m1 >>
rect 226 258 227 259 
<< m2 >>
rect 226 258 227 259 
<< m1 >>
rect 228 258 229 259 
<< m2 >>
rect 228 258 229 259 
<< m2c >>
rect 228 258 229 259 
<< m1 >>
rect 228 258 229 259 
<< m2 >>
rect 228 258 229 259 
<< m1 >>
rect 235 258 236 259 
<< m1 >>
rect 237 258 238 259 
<< m1 >>
rect 239 258 240 259 
<< m2 >>
rect 239 258 240 259 
<< m1 >>
rect 243 258 244 259 
<< m1 >>
rect 253 258 254 259 
<< m2 >>
rect 254 258 255 259 
<< m1 >>
rect 262 258 263 259 
<< m1 >>
rect 272 258 273 259 
<< m2 >>
rect 273 258 274 259 
<< m2 >>
rect 276 258 277 259 
<< m2 >>
rect 294 258 295 259 
<< m2 >>
rect 316 258 317 259 
<< m2 >>
rect 323 258 324 259 
<< m1 >>
rect 325 258 326 259 
<< m1 >>
rect 327 258 328 259 
<< m1 >>
rect 329 258 330 259 
<< m1 >>
rect 10 259 11 260 
<< m1 >>
rect 28 259 29 260 
<< m2 >>
rect 28 259 29 260 
<< m1 >>
rect 37 259 38 260 
<< m2 >>
rect 37 259 38 260 
<< m1 >>
rect 39 259 40 260 
<< m2 >>
rect 43 259 44 260 
<< m1 >>
rect 44 259 45 260 
<< m1 >>
rect 46 259 47 260 
<< m1 >>
rect 57 259 58 260 
<< m1 >>
rect 60 259 61 260 
<< m1 >>
rect 62 259 63 260 
<< m1 >>
rect 64 259 65 260 
<< m1 >>
rect 70 259 71 260 
<< m1 >>
rect 73 259 74 260 
<< m2 >>
rect 74 259 75 260 
<< m1 >>
rect 116 259 117 260 
<< m2 >>
rect 118 259 119 260 
<< m1 >>
rect 130 259 131 260 
<< m1 >>
rect 132 259 133 260 
<< m1 >>
rect 134 259 135 260 
<< m1 >>
rect 136 259 137 260 
<< m1 >>
rect 142 259 143 260 
<< m2 >>
rect 154 259 155 260 
<< m2 >>
rect 155 259 156 260 
<< m2 >>
rect 156 259 157 260 
<< m2 >>
rect 157 259 158 260 
<< m2 >>
rect 158 259 159 260 
<< m2 >>
rect 159 259 160 260 
<< m2 >>
rect 160 259 161 260 
<< m2 >>
rect 161 259 162 260 
<< m2 >>
rect 162 259 163 260 
<< m2 >>
rect 163 259 164 260 
<< m2 >>
rect 164 259 165 260 
<< m1 >>
rect 165 259 166 260 
<< m2 >>
rect 165 259 166 260 
<< m2 >>
rect 166 259 167 260 
<< m1 >>
rect 171 259 172 260 
<< m1 >>
rect 181 259 182 260 
<< m1 >>
rect 183 259 184 260 
<< m1 >>
rect 186 259 187 260 
<< m1 >>
rect 188 259 189 260 
<< m1 >>
rect 190 259 191 260 
<< m1 >>
rect 192 259 193 260 
<< m1 >>
rect 193 259 194 260 
<< m1 >>
rect 194 259 195 260 
<< m1 >>
rect 195 259 196 260 
<< m1 >>
rect 196 259 197 260 
<< m1 >>
rect 197 259 198 260 
<< m1 >>
rect 198 259 199 260 
<< m1 >>
rect 199 259 200 260 
<< m1 >>
rect 200 259 201 260 
<< m1 >>
rect 201 259 202 260 
<< m1 >>
rect 202 259 203 260 
<< m1 >>
rect 203 259 204 260 
<< m1 >>
rect 204 259 205 260 
<< m1 >>
rect 205 259 206 260 
<< m1 >>
rect 206 259 207 260 
<< m1 >>
rect 207 259 208 260 
<< m1 >>
rect 208 259 209 260 
<< m1 >>
rect 209 259 210 260 
<< m1 >>
rect 210 259 211 260 
<< m1 >>
rect 211 259 212 260 
<< m1 >>
rect 212 259 213 260 
<< m1 >>
rect 213 259 214 260 
<< m1 >>
rect 214 259 215 260 
<< m1 >>
rect 215 259 216 260 
<< m1 >>
rect 216 259 217 260 
<< m1 >>
rect 217 259 218 260 
<< m1 >>
rect 218 259 219 260 
<< m1 >>
rect 219 259 220 260 
<< m1 >>
rect 226 259 227 260 
<< m1 >>
rect 228 259 229 260 
<< m1 >>
rect 235 259 236 260 
<< m1 >>
rect 237 259 238 260 
<< m1 >>
rect 239 259 240 260 
<< m2 >>
rect 239 259 240 260 
<< m1 >>
rect 241 259 242 260 
<< m2 >>
rect 241 259 242 260 
<< m2c >>
rect 241 259 242 260 
<< m1 >>
rect 241 259 242 260 
<< m2 >>
rect 241 259 242 260 
<< m2 >>
rect 242 259 243 260 
<< m1 >>
rect 243 259 244 260 
<< m2 >>
rect 243 259 244 260 
<< m2 >>
rect 244 259 245 260 
<< m1 >>
rect 245 259 246 260 
<< m2 >>
rect 245 259 246 260 
<< m2c >>
rect 245 259 246 260 
<< m1 >>
rect 245 259 246 260 
<< m2 >>
rect 245 259 246 260 
<< m1 >>
rect 246 259 247 260 
<< m1 >>
rect 247 259 248 260 
<< m1 >>
rect 248 259 249 260 
<< m1 >>
rect 249 259 250 260 
<< m1 >>
rect 250 259 251 260 
<< m1 >>
rect 251 259 252 260 
<< m1 >>
rect 253 259 254 260 
<< m2 >>
rect 254 259 255 260 
<< m1 >>
rect 255 259 256 260 
<< m2 >>
rect 255 259 256 260 
<< m2c >>
rect 255 259 256 260 
<< m1 >>
rect 255 259 256 260 
<< m2 >>
rect 255 259 256 260 
<< m1 >>
rect 256 259 257 260 
<< m1 >>
rect 257 259 258 260 
<< m1 >>
rect 258 259 259 260 
<< m1 >>
rect 259 259 260 260 
<< m1 >>
rect 260 259 261 260 
<< m2 >>
rect 260 259 261 260 
<< m2c >>
rect 260 259 261 260 
<< m1 >>
rect 260 259 261 260 
<< m2 >>
rect 260 259 261 260 
<< m2 >>
rect 261 259 262 260 
<< m1 >>
rect 262 259 263 260 
<< m2 >>
rect 262 259 263 260 
<< m1 >>
rect 263 259 264 260 
<< m2 >>
rect 263 259 264 260 
<< m1 >>
rect 264 259 265 260 
<< m2 >>
rect 264 259 265 260 
<< m1 >>
rect 265 259 266 260 
<< m2 >>
rect 265 259 266 260 
<< m1 >>
rect 266 259 267 260 
<< m2 >>
rect 266 259 267 260 
<< m1 >>
rect 267 259 268 260 
<< m2 >>
rect 267 259 268 260 
<< m1 >>
rect 268 259 269 260 
<< m2 >>
rect 268 259 269 260 
<< m1 >>
rect 269 259 270 260 
<< m1 >>
rect 270 259 271 260 
<< m1 >>
rect 272 259 273 260 
<< m2 >>
rect 273 259 274 260 
<< m1 >>
rect 274 259 275 260 
<< m2 >>
rect 274 259 275 260 
<< m2c >>
rect 274 259 275 260 
<< m1 >>
rect 274 259 275 260 
<< m2 >>
rect 274 259 275 260 
<< m1 >>
rect 275 259 276 260 
<< m1 >>
rect 276 259 277 260 
<< m2 >>
rect 276 259 277 260 
<< m1 >>
rect 277 259 278 260 
<< m1 >>
rect 278 259 279 260 
<< m1 >>
rect 279 259 280 260 
<< m1 >>
rect 280 259 281 260 
<< m1 >>
rect 281 259 282 260 
<< m1 >>
rect 282 259 283 260 
<< m1 >>
rect 283 259 284 260 
<< m1 >>
rect 284 259 285 260 
<< m1 >>
rect 285 259 286 260 
<< m1 >>
rect 286 259 287 260 
<< m1 >>
rect 287 259 288 260 
<< m1 >>
rect 288 259 289 260 
<< m1 >>
rect 289 259 290 260 
<< m1 >>
rect 290 259 291 260 
<< m1 >>
rect 291 259 292 260 
<< m1 >>
rect 292 259 293 260 
<< m1 >>
rect 293 259 294 260 
<< m1 >>
rect 294 259 295 260 
<< m2 >>
rect 294 259 295 260 
<< m1 >>
rect 295 259 296 260 
<< m1 >>
rect 296 259 297 260 
<< m1 >>
rect 297 259 298 260 
<< m1 >>
rect 298 259 299 260 
<< m1 >>
rect 299 259 300 260 
<< m1 >>
rect 300 259 301 260 
<< m1 >>
rect 301 259 302 260 
<< m1 >>
rect 302 259 303 260 
<< m1 >>
rect 303 259 304 260 
<< m1 >>
rect 304 259 305 260 
<< m1 >>
rect 316 259 317 260 
<< m2 >>
rect 316 259 317 260 
<< m2c >>
rect 316 259 317 260 
<< m1 >>
rect 316 259 317 260 
<< m2 >>
rect 316 259 317 260 
<< m1 >>
rect 318 259 319 260 
<< m1 >>
rect 319 259 320 260 
<< m1 >>
rect 320 259 321 260 
<< m1 >>
rect 321 259 322 260 
<< m1 >>
rect 322 259 323 260 
<< m1 >>
rect 323 259 324 260 
<< m2 >>
rect 323 259 324 260 
<< m2c >>
rect 323 259 324 260 
<< m1 >>
rect 323 259 324 260 
<< m2 >>
rect 323 259 324 260 
<< m1 >>
rect 325 259 326 260 
<< m1 >>
rect 327 259 328 260 
<< m1 >>
rect 329 259 330 260 
<< m1 >>
rect 10 260 11 261 
<< m1 >>
rect 28 260 29 261 
<< m2 >>
rect 28 260 29 261 
<< m1 >>
rect 37 260 38 261 
<< m2 >>
rect 37 260 38 261 
<< m1 >>
rect 39 260 40 261 
<< m2 >>
rect 43 260 44 261 
<< m1 >>
rect 44 260 45 261 
<< m1 >>
rect 46 260 47 261 
<< m1 >>
rect 57 260 58 261 
<< m1 >>
rect 60 260 61 261 
<< m1 >>
rect 62 260 63 261 
<< m1 >>
rect 64 260 65 261 
<< m1 >>
rect 70 260 71 261 
<< m1 >>
rect 73 260 74 261 
<< m2 >>
rect 74 260 75 261 
<< m1 >>
rect 116 260 117 261 
<< m1 >>
rect 118 260 119 261 
<< m2 >>
rect 118 260 119 261 
<< m2c >>
rect 118 260 119 261 
<< m1 >>
rect 118 260 119 261 
<< m2 >>
rect 118 260 119 261 
<< m1 >>
rect 130 260 131 261 
<< m1 >>
rect 132 260 133 261 
<< m1 >>
rect 134 260 135 261 
<< m1 >>
rect 136 260 137 261 
<< m1 >>
rect 142 260 143 261 
<< m1 >>
rect 165 260 166 261 
<< m2 >>
rect 166 260 167 261 
<< m1 >>
rect 171 260 172 261 
<< m1 >>
rect 181 260 182 261 
<< m1 >>
rect 183 260 184 261 
<< m1 >>
rect 186 260 187 261 
<< m2 >>
rect 186 260 187 261 
<< m2c >>
rect 186 260 187 261 
<< m1 >>
rect 186 260 187 261 
<< m2 >>
rect 186 260 187 261 
<< m2 >>
rect 187 260 188 261 
<< m1 >>
rect 188 260 189 261 
<< m2 >>
rect 188 260 189 261 
<< m2 >>
rect 189 260 190 261 
<< m1 >>
rect 190 260 191 261 
<< m2 >>
rect 190 260 191 261 
<< m2 >>
rect 191 260 192 261 
<< m1 >>
rect 192 260 193 261 
<< m2 >>
rect 192 260 193 261 
<< m2c >>
rect 192 260 193 261 
<< m1 >>
rect 192 260 193 261 
<< m2 >>
rect 192 260 193 261 
<< m1 >>
rect 219 260 220 261 
<< m1 >>
rect 226 260 227 261 
<< m1 >>
rect 228 260 229 261 
<< m1 >>
rect 235 260 236 261 
<< m1 >>
rect 237 260 238 261 
<< m1 >>
rect 239 260 240 261 
<< m2 >>
rect 239 260 240 261 
<< m1 >>
rect 241 260 242 261 
<< m1 >>
rect 243 260 244 261 
<< m1 >>
rect 251 260 252 261 
<< m1 >>
rect 253 260 254 261 
<< m2 >>
rect 268 260 269 261 
<< m1 >>
rect 270 260 271 261 
<< m1 >>
rect 272 260 273 261 
<< m2 >>
rect 276 260 277 261 
<< m2 >>
rect 294 260 295 261 
<< m1 >>
rect 304 260 305 261 
<< m1 >>
rect 316 260 317 261 
<< m1 >>
rect 318 260 319 261 
<< m1 >>
rect 325 260 326 261 
<< m2 >>
rect 325 260 326 261 
<< m2c >>
rect 325 260 326 261 
<< m1 >>
rect 325 260 326 261 
<< m2 >>
rect 325 260 326 261 
<< m1 >>
rect 327 260 328 261 
<< m2 >>
rect 327 260 328 261 
<< m2c >>
rect 327 260 328 261 
<< m1 >>
rect 327 260 328 261 
<< m2 >>
rect 327 260 328 261 
<< m1 >>
rect 329 260 330 261 
<< m2 >>
rect 329 260 330 261 
<< m2c >>
rect 329 260 330 261 
<< m1 >>
rect 329 260 330 261 
<< m2 >>
rect 329 260 330 261 
<< m1 >>
rect 10 261 11 262 
<< m1 >>
rect 28 261 29 262 
<< m2 >>
rect 28 261 29 262 
<< m1 >>
rect 37 261 38 262 
<< m2 >>
rect 37 261 38 262 
<< m1 >>
rect 39 261 40 262 
<< m2 >>
rect 43 261 44 262 
<< m1 >>
rect 44 261 45 262 
<< m1 >>
rect 46 261 47 262 
<< m1 >>
rect 57 261 58 262 
<< m1 >>
rect 60 261 61 262 
<< m1 >>
rect 62 261 63 262 
<< m1 >>
rect 64 261 65 262 
<< m1 >>
rect 70 261 71 262 
<< m1 >>
rect 73 261 74 262 
<< m2 >>
rect 74 261 75 262 
<< m1 >>
rect 116 261 117 262 
<< m1 >>
rect 118 261 119 262 
<< m1 >>
rect 130 261 131 262 
<< m1 >>
rect 132 261 133 262 
<< m1 >>
rect 134 261 135 262 
<< m1 >>
rect 136 261 137 262 
<< m1 >>
rect 142 261 143 262 
<< m1 >>
rect 165 261 166 262 
<< m2 >>
rect 166 261 167 262 
<< m1 >>
rect 171 261 172 262 
<< m1 >>
rect 181 261 182 262 
<< m1 >>
rect 183 261 184 262 
<< m1 >>
rect 188 261 189 262 
<< m1 >>
rect 190 261 191 262 
<< m1 >>
rect 219 261 220 262 
<< m1 >>
rect 226 261 227 262 
<< m1 >>
rect 228 261 229 262 
<< m1 >>
rect 235 261 236 262 
<< m1 >>
rect 237 261 238 262 
<< m1 >>
rect 239 261 240 262 
<< m2 >>
rect 239 261 240 262 
<< m1 >>
rect 241 261 242 262 
<< m1 >>
rect 243 261 244 262 
<< m1 >>
rect 251 261 252 262 
<< m1 >>
rect 253 261 254 262 
<< m1 >>
rect 268 261 269 262 
<< m2 >>
rect 268 261 269 262 
<< m2c >>
rect 268 261 269 262 
<< m1 >>
rect 268 261 269 262 
<< m2 >>
rect 268 261 269 262 
<< m1 >>
rect 270 261 271 262 
<< m1 >>
rect 272 261 273 262 
<< m1 >>
rect 276 261 277 262 
<< m2 >>
rect 276 261 277 262 
<< m2c >>
rect 276 261 277 262 
<< m1 >>
rect 276 261 277 262 
<< m2 >>
rect 276 261 277 262 
<< m1 >>
rect 294 261 295 262 
<< m2 >>
rect 294 261 295 262 
<< m2c >>
rect 294 261 295 262 
<< m1 >>
rect 294 261 295 262 
<< m2 >>
rect 294 261 295 262 
<< m1 >>
rect 304 261 305 262 
<< m1 >>
rect 316 261 317 262 
<< m2 >>
rect 316 261 317 262 
<< m2 >>
rect 317 261 318 262 
<< m1 >>
rect 318 261 319 262 
<< m2 >>
rect 318 261 319 262 
<< m2c >>
rect 318 261 319 262 
<< m1 >>
rect 318 261 319 262 
<< m2 >>
rect 318 261 319 262 
<< m2 >>
rect 325 261 326 262 
<< m2 >>
rect 327 261 328 262 
<< m2 >>
rect 329 261 330 262 
<< m1 >>
rect 10 262 11 263 
<< m1 >>
rect 28 262 29 263 
<< m2 >>
rect 28 262 29 263 
<< m1 >>
rect 37 262 38 263 
<< m2 >>
rect 37 262 38 263 
<< m1 >>
rect 39 262 40 263 
<< m2 >>
rect 43 262 44 263 
<< m1 >>
rect 44 262 45 263 
<< m1 >>
rect 46 262 47 263 
<< m1 >>
rect 57 262 58 263 
<< m1 >>
rect 60 262 61 263 
<< m1 >>
rect 62 262 63 263 
<< m1 >>
rect 64 262 65 263 
<< m1 >>
rect 70 262 71 263 
<< m1 >>
rect 73 262 74 263 
<< m2 >>
rect 74 262 75 263 
<< m1 >>
rect 116 262 117 263 
<< m1 >>
rect 118 262 119 263 
<< m1 >>
rect 130 262 131 263 
<< m1 >>
rect 132 262 133 263 
<< m1 >>
rect 134 262 135 263 
<< m1 >>
rect 136 262 137 263 
<< m1 >>
rect 142 262 143 263 
<< m1 >>
rect 165 262 166 263 
<< m2 >>
rect 166 262 167 263 
<< m1 >>
rect 171 262 172 263 
<< m1 >>
rect 181 262 182 263 
<< m1 >>
rect 183 262 184 263 
<< m1 >>
rect 188 262 189 263 
<< m1 >>
rect 190 262 191 263 
<< m1 >>
rect 219 262 220 263 
<< m2 >>
rect 225 262 226 263 
<< m1 >>
rect 226 262 227 263 
<< m2 >>
rect 226 262 227 263 
<< m2 >>
rect 227 262 228 263 
<< m1 >>
rect 228 262 229 263 
<< m2 >>
rect 228 262 229 263 
<< m2c >>
rect 228 262 229 263 
<< m1 >>
rect 228 262 229 263 
<< m2 >>
rect 228 262 229 263 
<< m1 >>
rect 235 262 236 263 
<< m1 >>
rect 237 262 238 263 
<< m1 >>
rect 239 262 240 263 
<< m2 >>
rect 239 262 240 263 
<< m1 >>
rect 241 262 242 263 
<< m1 >>
rect 243 262 244 263 
<< m1 >>
rect 251 262 252 263 
<< m2 >>
rect 251 262 252 263 
<< m2c >>
rect 251 262 252 263 
<< m1 >>
rect 251 262 252 263 
<< m2 >>
rect 251 262 252 263 
<< m2 >>
rect 252 262 253 263 
<< m1 >>
rect 253 262 254 263 
<< m2 >>
rect 253 262 254 263 
<< m1 >>
rect 268 262 269 263 
<< m1 >>
rect 270 262 271 263 
<< m2 >>
rect 270 262 271 263 
<< m2c >>
rect 270 262 271 263 
<< m1 >>
rect 270 262 271 263 
<< m2 >>
rect 270 262 271 263 
<< m2 >>
rect 271 262 272 263 
<< m1 >>
rect 272 262 273 263 
<< m2 >>
rect 272 262 273 263 
<< m2 >>
rect 273 262 274 263 
<< m1 >>
rect 276 262 277 263 
<< m1 >>
rect 286 262 287 263 
<< m1 >>
rect 287 262 288 263 
<< m1 >>
rect 288 262 289 263 
<< m1 >>
rect 289 262 290 263 
<< m1 >>
rect 290 262 291 263 
<< m1 >>
rect 291 262 292 263 
<< m1 >>
rect 292 262 293 263 
<< m1 >>
rect 294 262 295 263 
<< m1 >>
rect 304 262 305 263 
<< m1 >>
rect 316 262 317 263 
<< m2 >>
rect 316 262 317 263 
<< m1 >>
rect 325 262 326 263 
<< m2 >>
rect 325 262 326 263 
<< m1 >>
rect 326 262 327 263 
<< m1 >>
rect 327 262 328 263 
<< m2 >>
rect 327 262 328 263 
<< m1 >>
rect 328 262 329 263 
<< m1 >>
rect 329 262 330 263 
<< m2 >>
rect 329 262 330 263 
<< m1 >>
rect 330 262 331 263 
<< m1 >>
rect 331 262 332 263 
<< m1 >>
rect 332 262 333 263 
<< m1 >>
rect 333 262 334 263 
<< m1 >>
rect 334 262 335 263 
<< m1 >>
rect 335 262 336 263 
<< m1 >>
rect 336 262 337 263 
<< m1 >>
rect 337 262 338 263 
<< m1 >>
rect 10 263 11 264 
<< m1 >>
rect 28 263 29 264 
<< m2 >>
rect 28 263 29 264 
<< m1 >>
rect 37 263 38 264 
<< m2 >>
rect 37 263 38 264 
<< m1 >>
rect 39 263 40 264 
<< m2 >>
rect 43 263 44 264 
<< m1 >>
rect 44 263 45 264 
<< m1 >>
rect 46 263 47 264 
<< m1 >>
rect 57 263 58 264 
<< m1 >>
rect 60 263 61 264 
<< m1 >>
rect 62 263 63 264 
<< m1 >>
rect 64 263 65 264 
<< m1 >>
rect 70 263 71 264 
<< m1 >>
rect 73 263 74 264 
<< m2 >>
rect 74 263 75 264 
<< m1 >>
rect 116 263 117 264 
<< m1 >>
rect 118 263 119 264 
<< m1 >>
rect 130 263 131 264 
<< m1 >>
rect 132 263 133 264 
<< m1 >>
rect 134 263 135 264 
<< m1 >>
rect 136 263 137 264 
<< m1 >>
rect 142 263 143 264 
<< m1 >>
rect 165 263 166 264 
<< m2 >>
rect 166 263 167 264 
<< m1 >>
rect 171 263 172 264 
<< m1 >>
rect 181 263 182 264 
<< m1 >>
rect 183 263 184 264 
<< m1 >>
rect 188 263 189 264 
<< m1 >>
rect 190 263 191 264 
<< m1 >>
rect 219 263 220 264 
<< m2 >>
rect 225 263 226 264 
<< m1 >>
rect 226 263 227 264 
<< m1 >>
rect 235 263 236 264 
<< m1 >>
rect 237 263 238 264 
<< m1 >>
rect 239 263 240 264 
<< m2 >>
rect 239 263 240 264 
<< m1 >>
rect 241 263 242 264 
<< m1 >>
rect 243 263 244 264 
<< m1 >>
rect 253 263 254 264 
<< m2 >>
rect 253 263 254 264 
<< m1 >>
rect 268 263 269 264 
<< m1 >>
rect 272 263 273 264 
<< m2 >>
rect 273 263 274 264 
<< m1 >>
rect 276 263 277 264 
<< m1 >>
rect 286 263 287 264 
<< m1 >>
rect 292 263 293 264 
<< m1 >>
rect 294 263 295 264 
<< m1 >>
rect 304 263 305 264 
<< m1 >>
rect 316 263 317 264 
<< m2 >>
rect 316 263 317 264 
<< m1 >>
rect 325 263 326 264 
<< m2 >>
rect 325 263 326 264 
<< m2 >>
rect 327 263 328 264 
<< m2 >>
rect 329 263 330 264 
<< m1 >>
rect 337 263 338 264 
<< m1 >>
rect 10 264 11 265 
<< pdiffusion >>
rect 12 264 13 265 
<< pdiffusion >>
rect 13 264 14 265 
<< pdiffusion >>
rect 14 264 15 265 
<< pdiffusion >>
rect 15 264 16 265 
<< pdiffusion >>
rect 16 264 17 265 
<< pdiffusion >>
rect 17 264 18 265 
<< m1 >>
rect 28 264 29 265 
<< m2 >>
rect 28 264 29 265 
<< pdiffusion >>
rect 30 264 31 265 
<< pdiffusion >>
rect 31 264 32 265 
<< pdiffusion >>
rect 32 264 33 265 
<< pdiffusion >>
rect 33 264 34 265 
<< pdiffusion >>
rect 34 264 35 265 
<< pdiffusion >>
rect 35 264 36 265 
<< m1 >>
rect 37 264 38 265 
<< m2 >>
rect 37 264 38 265 
<< m1 >>
rect 39 264 40 265 
<< m2 >>
rect 43 264 44 265 
<< m1 >>
rect 44 264 45 265 
<< m1 >>
rect 46 264 47 265 
<< pdiffusion >>
rect 48 264 49 265 
<< pdiffusion >>
rect 49 264 50 265 
<< pdiffusion >>
rect 50 264 51 265 
<< pdiffusion >>
rect 51 264 52 265 
<< pdiffusion >>
rect 52 264 53 265 
<< pdiffusion >>
rect 53 264 54 265 
<< m1 >>
rect 57 264 58 265 
<< m1 >>
rect 60 264 61 265 
<< m1 >>
rect 62 264 63 265 
<< m1 >>
rect 64 264 65 265 
<< pdiffusion >>
rect 66 264 67 265 
<< pdiffusion >>
rect 67 264 68 265 
<< pdiffusion >>
rect 68 264 69 265 
<< pdiffusion >>
rect 69 264 70 265 
<< m1 >>
rect 70 264 71 265 
<< pdiffusion >>
rect 70 264 71 265 
<< pdiffusion >>
rect 71 264 72 265 
<< m1 >>
rect 73 264 74 265 
<< m2 >>
rect 74 264 75 265 
<< pdiffusion >>
rect 84 264 85 265 
<< pdiffusion >>
rect 85 264 86 265 
<< pdiffusion >>
rect 86 264 87 265 
<< pdiffusion >>
rect 87 264 88 265 
<< pdiffusion >>
rect 88 264 89 265 
<< pdiffusion >>
rect 89 264 90 265 
<< pdiffusion >>
rect 102 264 103 265 
<< pdiffusion >>
rect 103 264 104 265 
<< pdiffusion >>
rect 104 264 105 265 
<< pdiffusion >>
rect 105 264 106 265 
<< pdiffusion >>
rect 106 264 107 265 
<< pdiffusion >>
rect 107 264 108 265 
<< m1 >>
rect 116 264 117 265 
<< m1 >>
rect 118 264 119 265 
<< pdiffusion >>
rect 120 264 121 265 
<< pdiffusion >>
rect 121 264 122 265 
<< pdiffusion >>
rect 122 264 123 265 
<< pdiffusion >>
rect 123 264 124 265 
<< pdiffusion >>
rect 124 264 125 265 
<< pdiffusion >>
rect 125 264 126 265 
<< m1 >>
rect 130 264 131 265 
<< m1 >>
rect 132 264 133 265 
<< m1 >>
rect 134 264 135 265 
<< m1 >>
rect 136 264 137 265 
<< pdiffusion >>
rect 138 264 139 265 
<< pdiffusion >>
rect 139 264 140 265 
<< pdiffusion >>
rect 140 264 141 265 
<< pdiffusion >>
rect 141 264 142 265 
<< m1 >>
rect 142 264 143 265 
<< pdiffusion >>
rect 142 264 143 265 
<< pdiffusion >>
rect 143 264 144 265 
<< pdiffusion >>
rect 156 264 157 265 
<< pdiffusion >>
rect 157 264 158 265 
<< pdiffusion >>
rect 158 264 159 265 
<< pdiffusion >>
rect 159 264 160 265 
<< pdiffusion >>
rect 160 264 161 265 
<< pdiffusion >>
rect 161 264 162 265 
<< m1 >>
rect 165 264 166 265 
<< m2 >>
rect 166 264 167 265 
<< m1 >>
rect 171 264 172 265 
<< pdiffusion >>
rect 174 264 175 265 
<< pdiffusion >>
rect 175 264 176 265 
<< pdiffusion >>
rect 176 264 177 265 
<< pdiffusion >>
rect 177 264 178 265 
<< pdiffusion >>
rect 178 264 179 265 
<< pdiffusion >>
rect 179 264 180 265 
<< m1 >>
rect 181 264 182 265 
<< m1 >>
rect 183 264 184 265 
<< m1 >>
rect 188 264 189 265 
<< m1 >>
rect 190 264 191 265 
<< pdiffusion >>
rect 192 264 193 265 
<< pdiffusion >>
rect 193 264 194 265 
<< pdiffusion >>
rect 194 264 195 265 
<< pdiffusion >>
rect 195 264 196 265 
<< pdiffusion >>
rect 196 264 197 265 
<< pdiffusion >>
rect 197 264 198 265 
<< pdiffusion >>
rect 210 264 211 265 
<< pdiffusion >>
rect 211 264 212 265 
<< pdiffusion >>
rect 212 264 213 265 
<< pdiffusion >>
rect 213 264 214 265 
<< pdiffusion >>
rect 214 264 215 265 
<< pdiffusion >>
rect 215 264 216 265 
<< m1 >>
rect 219 264 220 265 
<< m2 >>
rect 225 264 226 265 
<< m1 >>
rect 226 264 227 265 
<< pdiffusion >>
rect 228 264 229 265 
<< pdiffusion >>
rect 229 264 230 265 
<< pdiffusion >>
rect 230 264 231 265 
<< pdiffusion >>
rect 231 264 232 265 
<< pdiffusion >>
rect 232 264 233 265 
<< pdiffusion >>
rect 233 264 234 265 
<< m1 >>
rect 235 264 236 265 
<< m1 >>
rect 237 264 238 265 
<< m1 >>
rect 239 264 240 265 
<< m2 >>
rect 239 264 240 265 
<< m1 >>
rect 241 264 242 265 
<< m1 >>
rect 243 264 244 265 
<< pdiffusion >>
rect 246 264 247 265 
<< pdiffusion >>
rect 247 264 248 265 
<< pdiffusion >>
rect 248 264 249 265 
<< pdiffusion >>
rect 249 264 250 265 
<< pdiffusion >>
rect 250 264 251 265 
<< pdiffusion >>
rect 251 264 252 265 
<< m1 >>
rect 253 264 254 265 
<< m2 >>
rect 253 264 254 265 
<< pdiffusion >>
rect 264 264 265 265 
<< pdiffusion >>
rect 265 264 266 265 
<< pdiffusion >>
rect 266 264 267 265 
<< pdiffusion >>
rect 267 264 268 265 
<< m1 >>
rect 268 264 269 265 
<< pdiffusion >>
rect 268 264 269 265 
<< pdiffusion >>
rect 269 264 270 265 
<< m1 >>
rect 272 264 273 265 
<< m2 >>
rect 273 264 274 265 
<< m1 >>
rect 276 264 277 265 
<< pdiffusion >>
rect 282 264 283 265 
<< pdiffusion >>
rect 283 264 284 265 
<< pdiffusion >>
rect 284 264 285 265 
<< pdiffusion >>
rect 285 264 286 265 
<< m1 >>
rect 286 264 287 265 
<< pdiffusion >>
rect 286 264 287 265 
<< pdiffusion >>
rect 287 264 288 265 
<< m1 >>
rect 292 264 293 265 
<< m1 >>
rect 294 264 295 265 
<< pdiffusion >>
rect 300 264 301 265 
<< pdiffusion >>
rect 301 264 302 265 
<< pdiffusion >>
rect 302 264 303 265 
<< pdiffusion >>
rect 303 264 304 265 
<< m1 >>
rect 304 264 305 265 
<< pdiffusion >>
rect 304 264 305 265 
<< pdiffusion >>
rect 305 264 306 265 
<< m1 >>
rect 316 264 317 265 
<< m2 >>
rect 316 264 317 265 
<< pdiffusion >>
rect 318 264 319 265 
<< pdiffusion >>
rect 319 264 320 265 
<< pdiffusion >>
rect 320 264 321 265 
<< pdiffusion >>
rect 321 264 322 265 
<< pdiffusion >>
rect 322 264 323 265 
<< pdiffusion >>
rect 323 264 324 265 
<< m1 >>
rect 325 264 326 265 
<< m2 >>
rect 325 264 326 265 
<< m1 >>
rect 327 264 328 265 
<< m2 >>
rect 327 264 328 265 
<< m2c >>
rect 327 264 328 265 
<< m1 >>
rect 327 264 328 265 
<< m2 >>
rect 327 264 328 265 
<< m1 >>
rect 329 264 330 265 
<< m2 >>
rect 329 264 330 265 
<< m2c >>
rect 329 264 330 265 
<< m1 >>
rect 329 264 330 265 
<< m2 >>
rect 329 264 330 265 
<< m1 >>
rect 330 264 331 265 
<< m1 >>
rect 331 264 332 265 
<< pdiffusion >>
rect 336 264 337 265 
<< m1 >>
rect 337 264 338 265 
<< pdiffusion >>
rect 337 264 338 265 
<< pdiffusion >>
rect 338 264 339 265 
<< pdiffusion >>
rect 339 264 340 265 
<< pdiffusion >>
rect 340 264 341 265 
<< pdiffusion >>
rect 341 264 342 265 
<< m1 >>
rect 10 265 11 266 
<< pdiffusion >>
rect 12 265 13 266 
<< pdiffusion >>
rect 13 265 14 266 
<< pdiffusion >>
rect 14 265 15 266 
<< pdiffusion >>
rect 15 265 16 266 
<< pdiffusion >>
rect 16 265 17 266 
<< pdiffusion >>
rect 17 265 18 266 
<< m1 >>
rect 28 265 29 266 
<< m2 >>
rect 28 265 29 266 
<< pdiffusion >>
rect 30 265 31 266 
<< pdiffusion >>
rect 31 265 32 266 
<< pdiffusion >>
rect 32 265 33 266 
<< pdiffusion >>
rect 33 265 34 266 
<< pdiffusion >>
rect 34 265 35 266 
<< pdiffusion >>
rect 35 265 36 266 
<< m1 >>
rect 37 265 38 266 
<< m2 >>
rect 37 265 38 266 
<< m1 >>
rect 39 265 40 266 
<< m2 >>
rect 43 265 44 266 
<< m1 >>
rect 44 265 45 266 
<< m1 >>
rect 46 265 47 266 
<< pdiffusion >>
rect 48 265 49 266 
<< pdiffusion >>
rect 49 265 50 266 
<< pdiffusion >>
rect 50 265 51 266 
<< pdiffusion >>
rect 51 265 52 266 
<< pdiffusion >>
rect 52 265 53 266 
<< pdiffusion >>
rect 53 265 54 266 
<< m1 >>
rect 57 265 58 266 
<< m1 >>
rect 60 265 61 266 
<< m1 >>
rect 62 265 63 266 
<< m1 >>
rect 64 265 65 266 
<< pdiffusion >>
rect 66 265 67 266 
<< pdiffusion >>
rect 67 265 68 266 
<< pdiffusion >>
rect 68 265 69 266 
<< pdiffusion >>
rect 69 265 70 266 
<< pdiffusion >>
rect 70 265 71 266 
<< pdiffusion >>
rect 71 265 72 266 
<< m1 >>
rect 73 265 74 266 
<< m2 >>
rect 74 265 75 266 
<< pdiffusion >>
rect 84 265 85 266 
<< pdiffusion >>
rect 85 265 86 266 
<< pdiffusion >>
rect 86 265 87 266 
<< pdiffusion >>
rect 87 265 88 266 
<< pdiffusion >>
rect 88 265 89 266 
<< pdiffusion >>
rect 89 265 90 266 
<< pdiffusion >>
rect 102 265 103 266 
<< pdiffusion >>
rect 103 265 104 266 
<< pdiffusion >>
rect 104 265 105 266 
<< pdiffusion >>
rect 105 265 106 266 
<< pdiffusion >>
rect 106 265 107 266 
<< pdiffusion >>
rect 107 265 108 266 
<< m1 >>
rect 116 265 117 266 
<< m1 >>
rect 118 265 119 266 
<< pdiffusion >>
rect 120 265 121 266 
<< pdiffusion >>
rect 121 265 122 266 
<< pdiffusion >>
rect 122 265 123 266 
<< pdiffusion >>
rect 123 265 124 266 
<< pdiffusion >>
rect 124 265 125 266 
<< pdiffusion >>
rect 125 265 126 266 
<< m1 >>
rect 130 265 131 266 
<< m1 >>
rect 132 265 133 266 
<< m1 >>
rect 134 265 135 266 
<< m1 >>
rect 136 265 137 266 
<< pdiffusion >>
rect 138 265 139 266 
<< pdiffusion >>
rect 139 265 140 266 
<< pdiffusion >>
rect 140 265 141 266 
<< pdiffusion >>
rect 141 265 142 266 
<< pdiffusion >>
rect 142 265 143 266 
<< pdiffusion >>
rect 143 265 144 266 
<< pdiffusion >>
rect 156 265 157 266 
<< pdiffusion >>
rect 157 265 158 266 
<< pdiffusion >>
rect 158 265 159 266 
<< pdiffusion >>
rect 159 265 160 266 
<< pdiffusion >>
rect 160 265 161 266 
<< pdiffusion >>
rect 161 265 162 266 
<< m1 >>
rect 165 265 166 266 
<< m2 >>
rect 166 265 167 266 
<< m1 >>
rect 171 265 172 266 
<< pdiffusion >>
rect 174 265 175 266 
<< pdiffusion >>
rect 175 265 176 266 
<< pdiffusion >>
rect 176 265 177 266 
<< pdiffusion >>
rect 177 265 178 266 
<< pdiffusion >>
rect 178 265 179 266 
<< pdiffusion >>
rect 179 265 180 266 
<< m1 >>
rect 181 265 182 266 
<< m1 >>
rect 183 265 184 266 
<< m1 >>
rect 188 265 189 266 
<< m1 >>
rect 190 265 191 266 
<< pdiffusion >>
rect 192 265 193 266 
<< pdiffusion >>
rect 193 265 194 266 
<< pdiffusion >>
rect 194 265 195 266 
<< pdiffusion >>
rect 195 265 196 266 
<< pdiffusion >>
rect 196 265 197 266 
<< pdiffusion >>
rect 197 265 198 266 
<< pdiffusion >>
rect 210 265 211 266 
<< pdiffusion >>
rect 211 265 212 266 
<< pdiffusion >>
rect 212 265 213 266 
<< pdiffusion >>
rect 213 265 214 266 
<< pdiffusion >>
rect 214 265 215 266 
<< pdiffusion >>
rect 215 265 216 266 
<< m1 >>
rect 219 265 220 266 
<< m2 >>
rect 225 265 226 266 
<< m1 >>
rect 226 265 227 266 
<< pdiffusion >>
rect 228 265 229 266 
<< pdiffusion >>
rect 229 265 230 266 
<< pdiffusion >>
rect 230 265 231 266 
<< pdiffusion >>
rect 231 265 232 266 
<< pdiffusion >>
rect 232 265 233 266 
<< pdiffusion >>
rect 233 265 234 266 
<< m1 >>
rect 235 265 236 266 
<< m1 >>
rect 237 265 238 266 
<< m1 >>
rect 239 265 240 266 
<< m2 >>
rect 239 265 240 266 
<< m1 >>
rect 241 265 242 266 
<< m1 >>
rect 243 265 244 266 
<< pdiffusion >>
rect 246 265 247 266 
<< pdiffusion >>
rect 247 265 248 266 
<< pdiffusion >>
rect 248 265 249 266 
<< pdiffusion >>
rect 249 265 250 266 
<< pdiffusion >>
rect 250 265 251 266 
<< pdiffusion >>
rect 251 265 252 266 
<< m1 >>
rect 253 265 254 266 
<< m2 >>
rect 253 265 254 266 
<< pdiffusion >>
rect 264 265 265 266 
<< pdiffusion >>
rect 265 265 266 266 
<< pdiffusion >>
rect 266 265 267 266 
<< pdiffusion >>
rect 267 265 268 266 
<< pdiffusion >>
rect 268 265 269 266 
<< pdiffusion >>
rect 269 265 270 266 
<< m1 >>
rect 272 265 273 266 
<< m2 >>
rect 273 265 274 266 
<< m1 >>
rect 276 265 277 266 
<< pdiffusion >>
rect 282 265 283 266 
<< pdiffusion >>
rect 283 265 284 266 
<< pdiffusion >>
rect 284 265 285 266 
<< pdiffusion >>
rect 285 265 286 266 
<< pdiffusion >>
rect 286 265 287 266 
<< pdiffusion >>
rect 287 265 288 266 
<< m1 >>
rect 292 265 293 266 
<< m1 >>
rect 294 265 295 266 
<< pdiffusion >>
rect 300 265 301 266 
<< pdiffusion >>
rect 301 265 302 266 
<< pdiffusion >>
rect 302 265 303 266 
<< pdiffusion >>
rect 303 265 304 266 
<< pdiffusion >>
rect 304 265 305 266 
<< pdiffusion >>
rect 305 265 306 266 
<< m1 >>
rect 316 265 317 266 
<< m2 >>
rect 316 265 317 266 
<< pdiffusion >>
rect 318 265 319 266 
<< pdiffusion >>
rect 319 265 320 266 
<< pdiffusion >>
rect 320 265 321 266 
<< pdiffusion >>
rect 321 265 322 266 
<< pdiffusion >>
rect 322 265 323 266 
<< pdiffusion >>
rect 323 265 324 266 
<< m1 >>
rect 325 265 326 266 
<< m2 >>
rect 325 265 326 266 
<< m1 >>
rect 327 265 328 266 
<< m1 >>
rect 331 265 332 266 
<< pdiffusion >>
rect 336 265 337 266 
<< pdiffusion >>
rect 337 265 338 266 
<< pdiffusion >>
rect 338 265 339 266 
<< pdiffusion >>
rect 339 265 340 266 
<< pdiffusion >>
rect 340 265 341 266 
<< pdiffusion >>
rect 341 265 342 266 
<< m1 >>
rect 10 266 11 267 
<< pdiffusion >>
rect 12 266 13 267 
<< pdiffusion >>
rect 13 266 14 267 
<< pdiffusion >>
rect 14 266 15 267 
<< pdiffusion >>
rect 15 266 16 267 
<< pdiffusion >>
rect 16 266 17 267 
<< pdiffusion >>
rect 17 266 18 267 
<< m1 >>
rect 28 266 29 267 
<< m2 >>
rect 28 266 29 267 
<< pdiffusion >>
rect 30 266 31 267 
<< pdiffusion >>
rect 31 266 32 267 
<< pdiffusion >>
rect 32 266 33 267 
<< pdiffusion >>
rect 33 266 34 267 
<< pdiffusion >>
rect 34 266 35 267 
<< pdiffusion >>
rect 35 266 36 267 
<< m1 >>
rect 37 266 38 267 
<< m2 >>
rect 37 266 38 267 
<< m1 >>
rect 39 266 40 267 
<< m2 >>
rect 43 266 44 267 
<< m1 >>
rect 44 266 45 267 
<< m1 >>
rect 46 266 47 267 
<< pdiffusion >>
rect 48 266 49 267 
<< pdiffusion >>
rect 49 266 50 267 
<< pdiffusion >>
rect 50 266 51 267 
<< pdiffusion >>
rect 51 266 52 267 
<< pdiffusion >>
rect 52 266 53 267 
<< pdiffusion >>
rect 53 266 54 267 
<< m1 >>
rect 57 266 58 267 
<< m1 >>
rect 60 266 61 267 
<< m1 >>
rect 62 266 63 267 
<< m1 >>
rect 64 266 65 267 
<< pdiffusion >>
rect 66 266 67 267 
<< pdiffusion >>
rect 67 266 68 267 
<< pdiffusion >>
rect 68 266 69 267 
<< pdiffusion >>
rect 69 266 70 267 
<< pdiffusion >>
rect 70 266 71 267 
<< pdiffusion >>
rect 71 266 72 267 
<< m1 >>
rect 73 266 74 267 
<< m2 >>
rect 74 266 75 267 
<< pdiffusion >>
rect 84 266 85 267 
<< pdiffusion >>
rect 85 266 86 267 
<< pdiffusion >>
rect 86 266 87 267 
<< pdiffusion >>
rect 87 266 88 267 
<< pdiffusion >>
rect 88 266 89 267 
<< pdiffusion >>
rect 89 266 90 267 
<< pdiffusion >>
rect 102 266 103 267 
<< pdiffusion >>
rect 103 266 104 267 
<< pdiffusion >>
rect 104 266 105 267 
<< pdiffusion >>
rect 105 266 106 267 
<< pdiffusion >>
rect 106 266 107 267 
<< pdiffusion >>
rect 107 266 108 267 
<< m1 >>
rect 116 266 117 267 
<< m1 >>
rect 118 266 119 267 
<< pdiffusion >>
rect 120 266 121 267 
<< pdiffusion >>
rect 121 266 122 267 
<< pdiffusion >>
rect 122 266 123 267 
<< pdiffusion >>
rect 123 266 124 267 
<< pdiffusion >>
rect 124 266 125 267 
<< pdiffusion >>
rect 125 266 126 267 
<< m1 >>
rect 130 266 131 267 
<< m1 >>
rect 132 266 133 267 
<< m1 >>
rect 134 266 135 267 
<< m1 >>
rect 136 266 137 267 
<< pdiffusion >>
rect 138 266 139 267 
<< pdiffusion >>
rect 139 266 140 267 
<< pdiffusion >>
rect 140 266 141 267 
<< pdiffusion >>
rect 141 266 142 267 
<< pdiffusion >>
rect 142 266 143 267 
<< pdiffusion >>
rect 143 266 144 267 
<< pdiffusion >>
rect 156 266 157 267 
<< pdiffusion >>
rect 157 266 158 267 
<< pdiffusion >>
rect 158 266 159 267 
<< pdiffusion >>
rect 159 266 160 267 
<< pdiffusion >>
rect 160 266 161 267 
<< pdiffusion >>
rect 161 266 162 267 
<< m1 >>
rect 165 266 166 267 
<< m2 >>
rect 166 266 167 267 
<< m1 >>
rect 171 266 172 267 
<< pdiffusion >>
rect 174 266 175 267 
<< pdiffusion >>
rect 175 266 176 267 
<< pdiffusion >>
rect 176 266 177 267 
<< pdiffusion >>
rect 177 266 178 267 
<< pdiffusion >>
rect 178 266 179 267 
<< pdiffusion >>
rect 179 266 180 267 
<< m1 >>
rect 181 266 182 267 
<< m1 >>
rect 183 266 184 267 
<< m1 >>
rect 188 266 189 267 
<< m1 >>
rect 190 266 191 267 
<< pdiffusion >>
rect 192 266 193 267 
<< pdiffusion >>
rect 193 266 194 267 
<< pdiffusion >>
rect 194 266 195 267 
<< pdiffusion >>
rect 195 266 196 267 
<< pdiffusion >>
rect 196 266 197 267 
<< pdiffusion >>
rect 197 266 198 267 
<< pdiffusion >>
rect 210 266 211 267 
<< pdiffusion >>
rect 211 266 212 267 
<< pdiffusion >>
rect 212 266 213 267 
<< pdiffusion >>
rect 213 266 214 267 
<< pdiffusion >>
rect 214 266 215 267 
<< pdiffusion >>
rect 215 266 216 267 
<< m1 >>
rect 219 266 220 267 
<< m2 >>
rect 225 266 226 267 
<< m1 >>
rect 226 266 227 267 
<< pdiffusion >>
rect 228 266 229 267 
<< pdiffusion >>
rect 229 266 230 267 
<< pdiffusion >>
rect 230 266 231 267 
<< pdiffusion >>
rect 231 266 232 267 
<< pdiffusion >>
rect 232 266 233 267 
<< pdiffusion >>
rect 233 266 234 267 
<< m1 >>
rect 235 266 236 267 
<< m1 >>
rect 237 266 238 267 
<< m1 >>
rect 239 266 240 267 
<< m2 >>
rect 239 266 240 267 
<< m1 >>
rect 241 266 242 267 
<< m1 >>
rect 243 266 244 267 
<< pdiffusion >>
rect 246 266 247 267 
<< pdiffusion >>
rect 247 266 248 267 
<< pdiffusion >>
rect 248 266 249 267 
<< pdiffusion >>
rect 249 266 250 267 
<< pdiffusion >>
rect 250 266 251 267 
<< pdiffusion >>
rect 251 266 252 267 
<< m1 >>
rect 253 266 254 267 
<< m2 >>
rect 253 266 254 267 
<< pdiffusion >>
rect 264 266 265 267 
<< pdiffusion >>
rect 265 266 266 267 
<< pdiffusion >>
rect 266 266 267 267 
<< pdiffusion >>
rect 267 266 268 267 
<< pdiffusion >>
rect 268 266 269 267 
<< pdiffusion >>
rect 269 266 270 267 
<< m1 >>
rect 272 266 273 267 
<< m2 >>
rect 273 266 274 267 
<< m1 >>
rect 276 266 277 267 
<< pdiffusion >>
rect 282 266 283 267 
<< pdiffusion >>
rect 283 266 284 267 
<< pdiffusion >>
rect 284 266 285 267 
<< pdiffusion >>
rect 285 266 286 267 
<< pdiffusion >>
rect 286 266 287 267 
<< pdiffusion >>
rect 287 266 288 267 
<< m1 >>
rect 292 266 293 267 
<< m1 >>
rect 294 266 295 267 
<< pdiffusion >>
rect 300 266 301 267 
<< pdiffusion >>
rect 301 266 302 267 
<< pdiffusion >>
rect 302 266 303 267 
<< pdiffusion >>
rect 303 266 304 267 
<< pdiffusion >>
rect 304 266 305 267 
<< pdiffusion >>
rect 305 266 306 267 
<< m1 >>
rect 316 266 317 267 
<< m2 >>
rect 316 266 317 267 
<< pdiffusion >>
rect 318 266 319 267 
<< pdiffusion >>
rect 319 266 320 267 
<< pdiffusion >>
rect 320 266 321 267 
<< pdiffusion >>
rect 321 266 322 267 
<< pdiffusion >>
rect 322 266 323 267 
<< pdiffusion >>
rect 323 266 324 267 
<< m1 >>
rect 325 266 326 267 
<< m2 >>
rect 325 266 326 267 
<< m1 >>
rect 327 266 328 267 
<< m1 >>
rect 331 266 332 267 
<< pdiffusion >>
rect 336 266 337 267 
<< pdiffusion >>
rect 337 266 338 267 
<< pdiffusion >>
rect 338 266 339 267 
<< pdiffusion >>
rect 339 266 340 267 
<< pdiffusion >>
rect 340 266 341 267 
<< pdiffusion >>
rect 341 266 342 267 
<< m1 >>
rect 10 267 11 268 
<< pdiffusion >>
rect 12 267 13 268 
<< pdiffusion >>
rect 13 267 14 268 
<< pdiffusion >>
rect 14 267 15 268 
<< pdiffusion >>
rect 15 267 16 268 
<< pdiffusion >>
rect 16 267 17 268 
<< pdiffusion >>
rect 17 267 18 268 
<< m1 >>
rect 28 267 29 268 
<< m2 >>
rect 28 267 29 268 
<< pdiffusion >>
rect 30 267 31 268 
<< pdiffusion >>
rect 31 267 32 268 
<< pdiffusion >>
rect 32 267 33 268 
<< pdiffusion >>
rect 33 267 34 268 
<< pdiffusion >>
rect 34 267 35 268 
<< pdiffusion >>
rect 35 267 36 268 
<< m1 >>
rect 37 267 38 268 
<< m2 >>
rect 37 267 38 268 
<< m1 >>
rect 39 267 40 268 
<< m2 >>
rect 43 267 44 268 
<< m1 >>
rect 44 267 45 268 
<< m1 >>
rect 46 267 47 268 
<< pdiffusion >>
rect 48 267 49 268 
<< pdiffusion >>
rect 49 267 50 268 
<< pdiffusion >>
rect 50 267 51 268 
<< pdiffusion >>
rect 51 267 52 268 
<< pdiffusion >>
rect 52 267 53 268 
<< pdiffusion >>
rect 53 267 54 268 
<< m1 >>
rect 57 267 58 268 
<< m1 >>
rect 60 267 61 268 
<< m1 >>
rect 62 267 63 268 
<< m1 >>
rect 64 267 65 268 
<< pdiffusion >>
rect 66 267 67 268 
<< pdiffusion >>
rect 67 267 68 268 
<< pdiffusion >>
rect 68 267 69 268 
<< pdiffusion >>
rect 69 267 70 268 
<< pdiffusion >>
rect 70 267 71 268 
<< pdiffusion >>
rect 71 267 72 268 
<< m1 >>
rect 73 267 74 268 
<< m2 >>
rect 74 267 75 268 
<< pdiffusion >>
rect 84 267 85 268 
<< pdiffusion >>
rect 85 267 86 268 
<< pdiffusion >>
rect 86 267 87 268 
<< pdiffusion >>
rect 87 267 88 268 
<< pdiffusion >>
rect 88 267 89 268 
<< pdiffusion >>
rect 89 267 90 268 
<< pdiffusion >>
rect 102 267 103 268 
<< pdiffusion >>
rect 103 267 104 268 
<< pdiffusion >>
rect 104 267 105 268 
<< pdiffusion >>
rect 105 267 106 268 
<< pdiffusion >>
rect 106 267 107 268 
<< pdiffusion >>
rect 107 267 108 268 
<< m1 >>
rect 116 267 117 268 
<< m1 >>
rect 118 267 119 268 
<< pdiffusion >>
rect 120 267 121 268 
<< pdiffusion >>
rect 121 267 122 268 
<< pdiffusion >>
rect 122 267 123 268 
<< pdiffusion >>
rect 123 267 124 268 
<< pdiffusion >>
rect 124 267 125 268 
<< pdiffusion >>
rect 125 267 126 268 
<< m1 >>
rect 130 267 131 268 
<< m1 >>
rect 132 267 133 268 
<< m1 >>
rect 134 267 135 268 
<< m1 >>
rect 136 267 137 268 
<< pdiffusion >>
rect 138 267 139 268 
<< pdiffusion >>
rect 139 267 140 268 
<< pdiffusion >>
rect 140 267 141 268 
<< pdiffusion >>
rect 141 267 142 268 
<< pdiffusion >>
rect 142 267 143 268 
<< pdiffusion >>
rect 143 267 144 268 
<< pdiffusion >>
rect 156 267 157 268 
<< pdiffusion >>
rect 157 267 158 268 
<< pdiffusion >>
rect 158 267 159 268 
<< pdiffusion >>
rect 159 267 160 268 
<< pdiffusion >>
rect 160 267 161 268 
<< pdiffusion >>
rect 161 267 162 268 
<< m1 >>
rect 165 267 166 268 
<< m2 >>
rect 166 267 167 268 
<< m1 >>
rect 171 267 172 268 
<< pdiffusion >>
rect 174 267 175 268 
<< pdiffusion >>
rect 175 267 176 268 
<< pdiffusion >>
rect 176 267 177 268 
<< pdiffusion >>
rect 177 267 178 268 
<< pdiffusion >>
rect 178 267 179 268 
<< pdiffusion >>
rect 179 267 180 268 
<< m1 >>
rect 181 267 182 268 
<< m1 >>
rect 183 267 184 268 
<< m1 >>
rect 188 267 189 268 
<< m1 >>
rect 190 267 191 268 
<< pdiffusion >>
rect 192 267 193 268 
<< pdiffusion >>
rect 193 267 194 268 
<< pdiffusion >>
rect 194 267 195 268 
<< pdiffusion >>
rect 195 267 196 268 
<< pdiffusion >>
rect 196 267 197 268 
<< pdiffusion >>
rect 197 267 198 268 
<< pdiffusion >>
rect 210 267 211 268 
<< pdiffusion >>
rect 211 267 212 268 
<< pdiffusion >>
rect 212 267 213 268 
<< pdiffusion >>
rect 213 267 214 268 
<< pdiffusion >>
rect 214 267 215 268 
<< pdiffusion >>
rect 215 267 216 268 
<< m1 >>
rect 219 267 220 268 
<< m2 >>
rect 225 267 226 268 
<< m1 >>
rect 226 267 227 268 
<< pdiffusion >>
rect 228 267 229 268 
<< pdiffusion >>
rect 229 267 230 268 
<< pdiffusion >>
rect 230 267 231 268 
<< pdiffusion >>
rect 231 267 232 268 
<< pdiffusion >>
rect 232 267 233 268 
<< pdiffusion >>
rect 233 267 234 268 
<< m1 >>
rect 235 267 236 268 
<< m1 >>
rect 237 267 238 268 
<< m1 >>
rect 239 267 240 268 
<< m2 >>
rect 239 267 240 268 
<< m1 >>
rect 241 267 242 268 
<< m1 >>
rect 243 267 244 268 
<< pdiffusion >>
rect 246 267 247 268 
<< pdiffusion >>
rect 247 267 248 268 
<< pdiffusion >>
rect 248 267 249 268 
<< pdiffusion >>
rect 249 267 250 268 
<< pdiffusion >>
rect 250 267 251 268 
<< pdiffusion >>
rect 251 267 252 268 
<< m1 >>
rect 253 267 254 268 
<< m2 >>
rect 253 267 254 268 
<< pdiffusion >>
rect 264 267 265 268 
<< pdiffusion >>
rect 265 267 266 268 
<< pdiffusion >>
rect 266 267 267 268 
<< pdiffusion >>
rect 267 267 268 268 
<< pdiffusion >>
rect 268 267 269 268 
<< pdiffusion >>
rect 269 267 270 268 
<< m1 >>
rect 272 267 273 268 
<< m2 >>
rect 273 267 274 268 
<< m1 >>
rect 276 267 277 268 
<< pdiffusion >>
rect 282 267 283 268 
<< pdiffusion >>
rect 283 267 284 268 
<< pdiffusion >>
rect 284 267 285 268 
<< pdiffusion >>
rect 285 267 286 268 
<< pdiffusion >>
rect 286 267 287 268 
<< pdiffusion >>
rect 287 267 288 268 
<< m1 >>
rect 292 267 293 268 
<< m1 >>
rect 294 267 295 268 
<< pdiffusion >>
rect 300 267 301 268 
<< pdiffusion >>
rect 301 267 302 268 
<< pdiffusion >>
rect 302 267 303 268 
<< pdiffusion >>
rect 303 267 304 268 
<< pdiffusion >>
rect 304 267 305 268 
<< pdiffusion >>
rect 305 267 306 268 
<< m1 >>
rect 316 267 317 268 
<< m2 >>
rect 316 267 317 268 
<< pdiffusion >>
rect 318 267 319 268 
<< pdiffusion >>
rect 319 267 320 268 
<< pdiffusion >>
rect 320 267 321 268 
<< pdiffusion >>
rect 321 267 322 268 
<< pdiffusion >>
rect 322 267 323 268 
<< pdiffusion >>
rect 323 267 324 268 
<< m1 >>
rect 325 267 326 268 
<< m2 >>
rect 325 267 326 268 
<< m1 >>
rect 327 267 328 268 
<< m1 >>
rect 331 267 332 268 
<< pdiffusion >>
rect 336 267 337 268 
<< pdiffusion >>
rect 337 267 338 268 
<< pdiffusion >>
rect 338 267 339 268 
<< pdiffusion >>
rect 339 267 340 268 
<< pdiffusion >>
rect 340 267 341 268 
<< pdiffusion >>
rect 341 267 342 268 
<< m1 >>
rect 10 268 11 269 
<< pdiffusion >>
rect 12 268 13 269 
<< pdiffusion >>
rect 13 268 14 269 
<< pdiffusion >>
rect 14 268 15 269 
<< pdiffusion >>
rect 15 268 16 269 
<< pdiffusion >>
rect 16 268 17 269 
<< pdiffusion >>
rect 17 268 18 269 
<< m1 >>
rect 28 268 29 269 
<< m2 >>
rect 28 268 29 269 
<< pdiffusion >>
rect 30 268 31 269 
<< pdiffusion >>
rect 31 268 32 269 
<< pdiffusion >>
rect 32 268 33 269 
<< pdiffusion >>
rect 33 268 34 269 
<< pdiffusion >>
rect 34 268 35 269 
<< pdiffusion >>
rect 35 268 36 269 
<< m1 >>
rect 37 268 38 269 
<< m2 >>
rect 37 268 38 269 
<< m1 >>
rect 39 268 40 269 
<< m2 >>
rect 43 268 44 269 
<< m1 >>
rect 44 268 45 269 
<< m1 >>
rect 46 268 47 269 
<< pdiffusion >>
rect 48 268 49 269 
<< pdiffusion >>
rect 49 268 50 269 
<< pdiffusion >>
rect 50 268 51 269 
<< pdiffusion >>
rect 51 268 52 269 
<< pdiffusion >>
rect 52 268 53 269 
<< pdiffusion >>
rect 53 268 54 269 
<< m1 >>
rect 57 268 58 269 
<< m1 >>
rect 60 268 61 269 
<< m1 >>
rect 62 268 63 269 
<< m1 >>
rect 64 268 65 269 
<< pdiffusion >>
rect 66 268 67 269 
<< pdiffusion >>
rect 67 268 68 269 
<< pdiffusion >>
rect 68 268 69 269 
<< pdiffusion >>
rect 69 268 70 269 
<< pdiffusion >>
rect 70 268 71 269 
<< pdiffusion >>
rect 71 268 72 269 
<< m1 >>
rect 73 268 74 269 
<< m2 >>
rect 74 268 75 269 
<< pdiffusion >>
rect 84 268 85 269 
<< pdiffusion >>
rect 85 268 86 269 
<< pdiffusion >>
rect 86 268 87 269 
<< pdiffusion >>
rect 87 268 88 269 
<< pdiffusion >>
rect 88 268 89 269 
<< pdiffusion >>
rect 89 268 90 269 
<< pdiffusion >>
rect 102 268 103 269 
<< pdiffusion >>
rect 103 268 104 269 
<< pdiffusion >>
rect 104 268 105 269 
<< pdiffusion >>
rect 105 268 106 269 
<< pdiffusion >>
rect 106 268 107 269 
<< pdiffusion >>
rect 107 268 108 269 
<< m1 >>
rect 116 268 117 269 
<< m1 >>
rect 118 268 119 269 
<< pdiffusion >>
rect 120 268 121 269 
<< pdiffusion >>
rect 121 268 122 269 
<< pdiffusion >>
rect 122 268 123 269 
<< pdiffusion >>
rect 123 268 124 269 
<< pdiffusion >>
rect 124 268 125 269 
<< pdiffusion >>
rect 125 268 126 269 
<< m1 >>
rect 130 268 131 269 
<< m1 >>
rect 132 268 133 269 
<< m1 >>
rect 134 268 135 269 
<< m1 >>
rect 136 268 137 269 
<< pdiffusion >>
rect 138 268 139 269 
<< pdiffusion >>
rect 139 268 140 269 
<< pdiffusion >>
rect 140 268 141 269 
<< pdiffusion >>
rect 141 268 142 269 
<< pdiffusion >>
rect 142 268 143 269 
<< pdiffusion >>
rect 143 268 144 269 
<< pdiffusion >>
rect 156 268 157 269 
<< pdiffusion >>
rect 157 268 158 269 
<< pdiffusion >>
rect 158 268 159 269 
<< pdiffusion >>
rect 159 268 160 269 
<< pdiffusion >>
rect 160 268 161 269 
<< pdiffusion >>
rect 161 268 162 269 
<< m1 >>
rect 165 268 166 269 
<< m2 >>
rect 166 268 167 269 
<< m1 >>
rect 171 268 172 269 
<< pdiffusion >>
rect 174 268 175 269 
<< pdiffusion >>
rect 175 268 176 269 
<< pdiffusion >>
rect 176 268 177 269 
<< pdiffusion >>
rect 177 268 178 269 
<< pdiffusion >>
rect 178 268 179 269 
<< pdiffusion >>
rect 179 268 180 269 
<< m1 >>
rect 181 268 182 269 
<< m1 >>
rect 183 268 184 269 
<< m1 >>
rect 188 268 189 269 
<< m1 >>
rect 190 268 191 269 
<< pdiffusion >>
rect 192 268 193 269 
<< pdiffusion >>
rect 193 268 194 269 
<< pdiffusion >>
rect 194 268 195 269 
<< pdiffusion >>
rect 195 268 196 269 
<< pdiffusion >>
rect 196 268 197 269 
<< pdiffusion >>
rect 197 268 198 269 
<< pdiffusion >>
rect 210 268 211 269 
<< pdiffusion >>
rect 211 268 212 269 
<< pdiffusion >>
rect 212 268 213 269 
<< pdiffusion >>
rect 213 268 214 269 
<< pdiffusion >>
rect 214 268 215 269 
<< pdiffusion >>
rect 215 268 216 269 
<< m1 >>
rect 219 268 220 269 
<< m2 >>
rect 225 268 226 269 
<< m1 >>
rect 226 268 227 269 
<< pdiffusion >>
rect 228 268 229 269 
<< pdiffusion >>
rect 229 268 230 269 
<< pdiffusion >>
rect 230 268 231 269 
<< pdiffusion >>
rect 231 268 232 269 
<< pdiffusion >>
rect 232 268 233 269 
<< pdiffusion >>
rect 233 268 234 269 
<< m1 >>
rect 235 268 236 269 
<< m1 >>
rect 237 268 238 269 
<< m1 >>
rect 239 268 240 269 
<< m2 >>
rect 239 268 240 269 
<< m1 >>
rect 241 268 242 269 
<< m1 >>
rect 243 268 244 269 
<< pdiffusion >>
rect 246 268 247 269 
<< pdiffusion >>
rect 247 268 248 269 
<< pdiffusion >>
rect 248 268 249 269 
<< pdiffusion >>
rect 249 268 250 269 
<< pdiffusion >>
rect 250 268 251 269 
<< pdiffusion >>
rect 251 268 252 269 
<< m1 >>
rect 253 268 254 269 
<< m2 >>
rect 253 268 254 269 
<< pdiffusion >>
rect 264 268 265 269 
<< pdiffusion >>
rect 265 268 266 269 
<< pdiffusion >>
rect 266 268 267 269 
<< pdiffusion >>
rect 267 268 268 269 
<< pdiffusion >>
rect 268 268 269 269 
<< pdiffusion >>
rect 269 268 270 269 
<< m1 >>
rect 272 268 273 269 
<< m2 >>
rect 273 268 274 269 
<< m1 >>
rect 276 268 277 269 
<< pdiffusion >>
rect 282 268 283 269 
<< pdiffusion >>
rect 283 268 284 269 
<< pdiffusion >>
rect 284 268 285 269 
<< pdiffusion >>
rect 285 268 286 269 
<< pdiffusion >>
rect 286 268 287 269 
<< pdiffusion >>
rect 287 268 288 269 
<< m1 >>
rect 292 268 293 269 
<< m1 >>
rect 294 268 295 269 
<< pdiffusion >>
rect 300 268 301 269 
<< pdiffusion >>
rect 301 268 302 269 
<< pdiffusion >>
rect 302 268 303 269 
<< pdiffusion >>
rect 303 268 304 269 
<< pdiffusion >>
rect 304 268 305 269 
<< pdiffusion >>
rect 305 268 306 269 
<< m1 >>
rect 316 268 317 269 
<< m2 >>
rect 316 268 317 269 
<< pdiffusion >>
rect 318 268 319 269 
<< pdiffusion >>
rect 319 268 320 269 
<< pdiffusion >>
rect 320 268 321 269 
<< pdiffusion >>
rect 321 268 322 269 
<< pdiffusion >>
rect 322 268 323 269 
<< pdiffusion >>
rect 323 268 324 269 
<< m1 >>
rect 325 268 326 269 
<< m2 >>
rect 325 268 326 269 
<< m1 >>
rect 327 268 328 269 
<< m1 >>
rect 331 268 332 269 
<< pdiffusion >>
rect 336 268 337 269 
<< pdiffusion >>
rect 337 268 338 269 
<< pdiffusion >>
rect 338 268 339 269 
<< pdiffusion >>
rect 339 268 340 269 
<< pdiffusion >>
rect 340 268 341 269 
<< pdiffusion >>
rect 341 268 342 269 
<< m1 >>
rect 10 269 11 270 
<< pdiffusion >>
rect 12 269 13 270 
<< pdiffusion >>
rect 13 269 14 270 
<< pdiffusion >>
rect 14 269 15 270 
<< pdiffusion >>
rect 15 269 16 270 
<< pdiffusion >>
rect 16 269 17 270 
<< pdiffusion >>
rect 17 269 18 270 
<< m1 >>
rect 28 269 29 270 
<< m2 >>
rect 28 269 29 270 
<< pdiffusion >>
rect 30 269 31 270 
<< m1 >>
rect 31 269 32 270 
<< pdiffusion >>
rect 31 269 32 270 
<< pdiffusion >>
rect 32 269 33 270 
<< pdiffusion >>
rect 33 269 34 270 
<< pdiffusion >>
rect 34 269 35 270 
<< pdiffusion >>
rect 35 269 36 270 
<< m1 >>
rect 37 269 38 270 
<< m2 >>
rect 37 269 38 270 
<< m1 >>
rect 39 269 40 270 
<< m2 >>
rect 43 269 44 270 
<< m1 >>
rect 44 269 45 270 
<< m1 >>
rect 46 269 47 270 
<< pdiffusion >>
rect 48 269 49 270 
<< m1 >>
rect 49 269 50 270 
<< pdiffusion >>
rect 49 269 50 270 
<< pdiffusion >>
rect 50 269 51 270 
<< pdiffusion >>
rect 51 269 52 270 
<< m1 >>
rect 52 269 53 270 
<< pdiffusion >>
rect 52 269 53 270 
<< pdiffusion >>
rect 53 269 54 270 
<< m1 >>
rect 57 269 58 270 
<< m1 >>
rect 60 269 61 270 
<< m1 >>
rect 62 269 63 270 
<< m1 >>
rect 64 269 65 270 
<< pdiffusion >>
rect 66 269 67 270 
<< pdiffusion >>
rect 67 269 68 270 
<< pdiffusion >>
rect 68 269 69 270 
<< pdiffusion >>
rect 69 269 70 270 
<< pdiffusion >>
rect 70 269 71 270 
<< pdiffusion >>
rect 71 269 72 270 
<< m1 >>
rect 73 269 74 270 
<< m2 >>
rect 74 269 75 270 
<< pdiffusion >>
rect 84 269 85 270 
<< pdiffusion >>
rect 85 269 86 270 
<< pdiffusion >>
rect 86 269 87 270 
<< pdiffusion >>
rect 87 269 88 270 
<< pdiffusion >>
rect 88 269 89 270 
<< pdiffusion >>
rect 89 269 90 270 
<< pdiffusion >>
rect 102 269 103 270 
<< pdiffusion >>
rect 103 269 104 270 
<< pdiffusion >>
rect 104 269 105 270 
<< pdiffusion >>
rect 105 269 106 270 
<< pdiffusion >>
rect 106 269 107 270 
<< pdiffusion >>
rect 107 269 108 270 
<< m1 >>
rect 116 269 117 270 
<< m1 >>
rect 118 269 119 270 
<< pdiffusion >>
rect 120 269 121 270 
<< m1 >>
rect 121 269 122 270 
<< pdiffusion >>
rect 121 269 122 270 
<< pdiffusion >>
rect 122 269 123 270 
<< pdiffusion >>
rect 123 269 124 270 
<< pdiffusion >>
rect 124 269 125 270 
<< pdiffusion >>
rect 125 269 126 270 
<< m1 >>
rect 130 269 131 270 
<< m1 >>
rect 132 269 133 270 
<< m1 >>
rect 134 269 135 270 
<< m1 >>
rect 136 269 137 270 
<< pdiffusion >>
rect 138 269 139 270 
<< pdiffusion >>
rect 139 269 140 270 
<< pdiffusion >>
rect 140 269 141 270 
<< pdiffusion >>
rect 141 269 142 270 
<< pdiffusion >>
rect 142 269 143 270 
<< pdiffusion >>
rect 143 269 144 270 
<< pdiffusion >>
rect 156 269 157 270 
<< pdiffusion >>
rect 157 269 158 270 
<< pdiffusion >>
rect 158 269 159 270 
<< pdiffusion >>
rect 159 269 160 270 
<< pdiffusion >>
rect 160 269 161 270 
<< pdiffusion >>
rect 161 269 162 270 
<< m1 >>
rect 165 269 166 270 
<< m2 >>
rect 166 269 167 270 
<< m1 >>
rect 171 269 172 270 
<< pdiffusion >>
rect 174 269 175 270 
<< pdiffusion >>
rect 175 269 176 270 
<< pdiffusion >>
rect 176 269 177 270 
<< pdiffusion >>
rect 177 269 178 270 
<< pdiffusion >>
rect 178 269 179 270 
<< pdiffusion >>
rect 179 269 180 270 
<< m1 >>
rect 181 269 182 270 
<< m1 >>
rect 183 269 184 270 
<< m1 >>
rect 188 269 189 270 
<< m1 >>
rect 190 269 191 270 
<< pdiffusion >>
rect 192 269 193 270 
<< pdiffusion >>
rect 193 269 194 270 
<< pdiffusion >>
rect 194 269 195 270 
<< pdiffusion >>
rect 195 269 196 270 
<< pdiffusion >>
rect 196 269 197 270 
<< pdiffusion >>
rect 197 269 198 270 
<< pdiffusion >>
rect 210 269 211 270 
<< pdiffusion >>
rect 211 269 212 270 
<< pdiffusion >>
rect 212 269 213 270 
<< pdiffusion >>
rect 213 269 214 270 
<< pdiffusion >>
rect 214 269 215 270 
<< pdiffusion >>
rect 215 269 216 270 
<< m1 >>
rect 219 269 220 270 
<< m2 >>
rect 225 269 226 270 
<< m1 >>
rect 226 269 227 270 
<< pdiffusion >>
rect 228 269 229 270 
<< pdiffusion >>
rect 229 269 230 270 
<< pdiffusion >>
rect 230 269 231 270 
<< pdiffusion >>
rect 231 269 232 270 
<< pdiffusion >>
rect 232 269 233 270 
<< pdiffusion >>
rect 233 269 234 270 
<< m1 >>
rect 235 269 236 270 
<< m1 >>
rect 237 269 238 270 
<< m1 >>
rect 239 269 240 270 
<< m2 >>
rect 239 269 240 270 
<< m1 >>
rect 241 269 242 270 
<< m2 >>
rect 241 269 242 270 
<< m2c >>
rect 241 269 242 270 
<< m1 >>
rect 241 269 242 270 
<< m2 >>
rect 241 269 242 270 
<< m1 >>
rect 243 269 244 270 
<< m2 >>
rect 243 269 244 270 
<< m2c >>
rect 243 269 244 270 
<< m1 >>
rect 243 269 244 270 
<< m2 >>
rect 243 269 244 270 
<< pdiffusion >>
rect 246 269 247 270 
<< m1 >>
rect 247 269 248 270 
<< pdiffusion >>
rect 247 269 248 270 
<< pdiffusion >>
rect 248 269 249 270 
<< pdiffusion >>
rect 249 269 250 270 
<< m1 >>
rect 250 269 251 270 
<< pdiffusion >>
rect 250 269 251 270 
<< pdiffusion >>
rect 251 269 252 270 
<< m1 >>
rect 253 269 254 270 
<< m2 >>
rect 253 269 254 270 
<< pdiffusion >>
rect 264 269 265 270 
<< pdiffusion >>
rect 265 269 266 270 
<< pdiffusion >>
rect 266 269 267 270 
<< pdiffusion >>
rect 267 269 268 270 
<< pdiffusion >>
rect 268 269 269 270 
<< pdiffusion >>
rect 269 269 270 270 
<< m1 >>
rect 272 269 273 270 
<< m2 >>
rect 273 269 274 270 
<< m1 >>
rect 276 269 277 270 
<< pdiffusion >>
rect 282 269 283 270 
<< m1 >>
rect 283 269 284 270 
<< pdiffusion >>
rect 283 269 284 270 
<< pdiffusion >>
rect 284 269 285 270 
<< pdiffusion >>
rect 285 269 286 270 
<< pdiffusion >>
rect 286 269 287 270 
<< pdiffusion >>
rect 287 269 288 270 
<< m1 >>
rect 292 269 293 270 
<< m1 >>
rect 294 269 295 270 
<< pdiffusion >>
rect 300 269 301 270 
<< pdiffusion >>
rect 301 269 302 270 
<< pdiffusion >>
rect 302 269 303 270 
<< pdiffusion >>
rect 303 269 304 270 
<< pdiffusion >>
rect 304 269 305 270 
<< pdiffusion >>
rect 305 269 306 270 
<< m1 >>
rect 316 269 317 270 
<< m2 >>
rect 316 269 317 270 
<< pdiffusion >>
rect 318 269 319 270 
<< pdiffusion >>
rect 319 269 320 270 
<< pdiffusion >>
rect 320 269 321 270 
<< pdiffusion >>
rect 321 269 322 270 
<< m1 >>
rect 322 269 323 270 
<< pdiffusion >>
rect 322 269 323 270 
<< pdiffusion >>
rect 323 269 324 270 
<< m1 >>
rect 325 269 326 270 
<< m2 >>
rect 325 269 326 270 
<< m1 >>
rect 327 269 328 270 
<< m1 >>
rect 331 269 332 270 
<< pdiffusion >>
rect 336 269 337 270 
<< pdiffusion >>
rect 337 269 338 270 
<< pdiffusion >>
rect 338 269 339 270 
<< pdiffusion >>
rect 339 269 340 270 
<< pdiffusion >>
rect 340 269 341 270 
<< pdiffusion >>
rect 341 269 342 270 
<< m1 >>
rect 10 270 11 271 
<< m1 >>
rect 28 270 29 271 
<< m2 >>
rect 28 270 29 271 
<< m1 >>
rect 31 270 32 271 
<< m1 >>
rect 37 270 38 271 
<< m2 >>
rect 37 270 38 271 
<< m1 >>
rect 39 270 40 271 
<< m2 >>
rect 43 270 44 271 
<< m1 >>
rect 44 270 45 271 
<< m1 >>
rect 46 270 47 271 
<< m1 >>
rect 49 270 50 271 
<< m1 >>
rect 52 270 53 271 
<< m1 >>
rect 57 270 58 271 
<< m1 >>
rect 60 270 61 271 
<< m1 >>
rect 62 270 63 271 
<< m1 >>
rect 64 270 65 271 
<< m1 >>
rect 73 270 74 271 
<< m2 >>
rect 74 270 75 271 
<< m1 >>
rect 116 270 117 271 
<< m1 >>
rect 118 270 119 271 
<< m1 >>
rect 121 270 122 271 
<< m1 >>
rect 130 270 131 271 
<< m1 >>
rect 132 270 133 271 
<< m1 >>
rect 134 270 135 271 
<< m1 >>
rect 136 270 137 271 
<< m1 >>
rect 165 270 166 271 
<< m2 >>
rect 166 270 167 271 
<< m1 >>
rect 171 270 172 271 
<< m1 >>
rect 181 270 182 271 
<< m1 >>
rect 183 270 184 271 
<< m1 >>
rect 188 270 189 271 
<< m1 >>
rect 190 270 191 271 
<< m1 >>
rect 219 270 220 271 
<< m2 >>
rect 225 270 226 271 
<< m1 >>
rect 226 270 227 271 
<< m1 >>
rect 235 270 236 271 
<< m1 >>
rect 237 270 238 271 
<< m1 >>
rect 239 270 240 271 
<< m2 >>
rect 239 270 240 271 
<< m2 >>
rect 241 270 242 271 
<< m2 >>
rect 243 270 244 271 
<< m1 >>
rect 247 270 248 271 
<< m1 >>
rect 250 270 251 271 
<< m1 >>
rect 253 270 254 271 
<< m2 >>
rect 253 270 254 271 
<< m1 >>
rect 272 270 273 271 
<< m2 >>
rect 273 270 274 271 
<< m1 >>
rect 274 270 275 271 
<< m2 >>
rect 274 270 275 271 
<< m2c >>
rect 274 270 275 271 
<< m1 >>
rect 274 270 275 271 
<< m2 >>
rect 274 270 275 271 
<< m2 >>
rect 275 270 276 271 
<< m1 >>
rect 276 270 277 271 
<< m2 >>
rect 276 270 277 271 
<< m2 >>
rect 277 270 278 271 
<< m1 >>
rect 278 270 279 271 
<< m2 >>
rect 278 270 279 271 
<< m2c >>
rect 278 270 279 271 
<< m1 >>
rect 278 270 279 271 
<< m2 >>
rect 278 270 279 271 
<< m1 >>
rect 283 270 284 271 
<< m1 >>
rect 292 270 293 271 
<< m2 >>
rect 292 270 293 271 
<< m2c >>
rect 292 270 293 271 
<< m1 >>
rect 292 270 293 271 
<< m2 >>
rect 292 270 293 271 
<< m2 >>
rect 293 270 294 271 
<< m1 >>
rect 294 270 295 271 
<< m2 >>
rect 294 270 295 271 
<< m2 >>
rect 295 270 296 271 
<< m1 >>
rect 316 270 317 271 
<< m2 >>
rect 316 270 317 271 
<< m1 >>
rect 322 270 323 271 
<< m1 >>
rect 325 270 326 271 
<< m2 >>
rect 325 270 326 271 
<< m1 >>
rect 327 270 328 271 
<< m1 >>
rect 331 270 332 271 
<< m1 >>
rect 10 271 11 272 
<< m1 >>
rect 28 271 29 272 
<< m2 >>
rect 28 271 29 272 
<< m1 >>
rect 31 271 32 272 
<< m1 >>
rect 35 271 36 272 
<< m2 >>
rect 35 271 36 272 
<< m2c >>
rect 35 271 36 272 
<< m1 >>
rect 35 271 36 272 
<< m2 >>
rect 35 271 36 272 
<< m2 >>
rect 36 271 37 272 
<< m1 >>
rect 37 271 38 272 
<< m2 >>
rect 37 271 38 272 
<< m1 >>
rect 39 271 40 272 
<< m2 >>
rect 43 271 44 272 
<< m1 >>
rect 44 271 45 272 
<< m1 >>
rect 46 271 47 272 
<< m1 >>
rect 47 271 48 272 
<< m1 >>
rect 48 271 49 272 
<< m1 >>
rect 49 271 50 272 
<< m1 >>
rect 52 271 53 272 
<< m1 >>
rect 57 271 58 272 
<< m1 >>
rect 60 271 61 272 
<< m1 >>
rect 62 271 63 272 
<< m1 >>
rect 64 271 65 272 
<< m1 >>
rect 71 271 72 272 
<< m2 >>
rect 71 271 72 272 
<< m2c >>
rect 71 271 72 272 
<< m1 >>
rect 71 271 72 272 
<< m2 >>
rect 71 271 72 272 
<< m2 >>
rect 72 271 73 272 
<< m1 >>
rect 73 271 74 272 
<< m2 >>
rect 73 271 74 272 
<< m2 >>
rect 74 271 75 272 
<< m1 >>
rect 116 271 117 272 
<< m1 >>
rect 118 271 119 272 
<< m1 >>
rect 119 271 120 272 
<< m1 >>
rect 120 271 121 272 
<< m1 >>
rect 121 271 122 272 
<< m1 >>
rect 130 271 131 272 
<< m1 >>
rect 132 271 133 272 
<< m1 >>
rect 134 271 135 272 
<< m1 >>
rect 136 271 137 272 
<< m1 >>
rect 165 271 166 272 
<< m2 >>
rect 166 271 167 272 
<< m1 >>
rect 171 271 172 272 
<< m1 >>
rect 181 271 182 272 
<< m1 >>
rect 183 271 184 272 
<< m1 >>
rect 188 271 189 272 
<< m1 >>
rect 190 271 191 272 
<< m1 >>
rect 219 271 220 272 
<< m2 >>
rect 225 271 226 272 
<< m1 >>
rect 226 271 227 272 
<< m1 >>
rect 235 271 236 272 
<< m1 >>
rect 237 271 238 272 
<< m1 >>
rect 239 271 240 272 
<< m2 >>
rect 239 271 240 272 
<< m1 >>
rect 240 271 241 272 
<< m1 >>
rect 241 271 242 272 
<< m2 >>
rect 241 271 242 272 
<< m1 >>
rect 242 271 243 272 
<< m1 >>
rect 243 271 244 272 
<< m2 >>
rect 243 271 244 272 
<< m1 >>
rect 244 271 245 272 
<< m1 >>
rect 245 271 246 272 
<< m1 >>
rect 246 271 247 272 
<< m1 >>
rect 247 271 248 272 
<< m1 >>
rect 250 271 251 272 
<< m1 >>
rect 251 271 252 272 
<< m2 >>
rect 251 271 252 272 
<< m2c >>
rect 251 271 252 272 
<< m1 >>
rect 251 271 252 272 
<< m2 >>
rect 251 271 252 272 
<< m2 >>
rect 252 271 253 272 
<< m1 >>
rect 253 271 254 272 
<< m2 >>
rect 253 271 254 272 
<< m1 >>
rect 272 271 273 272 
<< m1 >>
rect 276 271 277 272 
<< m1 >>
rect 278 271 279 272 
<< m1 >>
rect 283 271 284 272 
<< m1 >>
rect 294 271 295 272 
<< m2 >>
rect 295 271 296 272 
<< m1 >>
rect 316 271 317 272 
<< m2 >>
rect 316 271 317 272 
<< m1 >>
rect 322 271 323 272 
<< m1 >>
rect 325 271 326 272 
<< m2 >>
rect 325 271 326 272 
<< m1 >>
rect 327 271 328 272 
<< m1 >>
rect 331 271 332 272 
<< m1 >>
rect 10 272 11 273 
<< m1 >>
rect 28 272 29 273 
<< m2 >>
rect 28 272 29 273 
<< m1 >>
rect 31 272 32 273 
<< m1 >>
rect 32 272 33 273 
<< m1 >>
rect 33 272 34 273 
<< m1 >>
rect 34 272 35 273 
<< m1 >>
rect 35 272 36 273 
<< m1 >>
rect 37 272 38 273 
<< m1 >>
rect 39 272 40 273 
<< m2 >>
rect 43 272 44 273 
<< m1 >>
rect 44 272 45 273 
<< m1 >>
rect 52 272 53 273 
<< m1 >>
rect 57 272 58 273 
<< m1 >>
rect 60 272 61 273 
<< m1 >>
rect 62 272 63 273 
<< m1 >>
rect 64 272 65 273 
<< m1 >>
rect 69 272 70 273 
<< m1 >>
rect 70 272 71 273 
<< m1 >>
rect 71 272 72 273 
<< m1 >>
rect 73 272 74 273 
<< m1 >>
rect 116 272 117 273 
<< m1 >>
rect 130 272 131 273 
<< m1 >>
rect 132 272 133 273 
<< m1 >>
rect 134 272 135 273 
<< m1 >>
rect 136 272 137 273 
<< m1 >>
rect 165 272 166 273 
<< m2 >>
rect 166 272 167 273 
<< m1 >>
rect 171 272 172 273 
<< m1 >>
rect 181 272 182 273 
<< m1 >>
rect 183 272 184 273 
<< m1 >>
rect 188 272 189 273 
<< m1 >>
rect 190 272 191 273 
<< m1 >>
rect 219 272 220 273 
<< m2 >>
rect 225 272 226 273 
<< m1 >>
rect 226 272 227 273 
<< m2 >>
rect 234 272 235 273 
<< m1 >>
rect 235 272 236 273 
<< m2 >>
rect 235 272 236 273 
<< m2 >>
rect 236 272 237 273 
<< m1 >>
rect 237 272 238 273 
<< m2 >>
rect 237 272 238 273 
<< m2c >>
rect 237 272 238 273 
<< m1 >>
rect 237 272 238 273 
<< m2 >>
rect 237 272 238 273 
<< m2 >>
rect 239 272 240 273 
<< m2 >>
rect 241 272 242 273 
<< m2 >>
rect 243 272 244 273 
<< m1 >>
rect 253 272 254 273 
<< m1 >>
rect 272 272 273 273 
<< m2 >>
rect 272 272 273 273 
<< m2c >>
rect 272 272 273 273 
<< m1 >>
rect 272 272 273 273 
<< m2 >>
rect 272 272 273 273 
<< m1 >>
rect 276 272 277 273 
<< m2 >>
rect 276 272 277 273 
<< m2c >>
rect 276 272 277 273 
<< m1 >>
rect 276 272 277 273 
<< m2 >>
rect 276 272 277 273 
<< m1 >>
rect 278 272 279 273 
<< m2 >>
rect 278 272 279 273 
<< m2c >>
rect 278 272 279 273 
<< m1 >>
rect 278 272 279 273 
<< m2 >>
rect 278 272 279 273 
<< m1 >>
rect 283 272 284 273 
<< m1 >>
rect 284 272 285 273 
<< m1 >>
rect 285 272 286 273 
<< m1 >>
rect 286 272 287 273 
<< m1 >>
rect 287 272 288 273 
<< m1 >>
rect 288 272 289 273 
<< m1 >>
rect 289 272 290 273 
<< m1 >>
rect 290 272 291 273 
<< m1 >>
rect 291 272 292 273 
<< m1 >>
rect 292 272 293 273 
<< m1 >>
rect 293 272 294 273 
<< m1 >>
rect 294 272 295 273 
<< m2 >>
rect 295 272 296 273 
<< m1 >>
rect 316 272 317 273 
<< m2 >>
rect 316 272 317 273 
<< m1 >>
rect 322 272 323 273 
<< m1 >>
rect 325 272 326 273 
<< m2 >>
rect 325 272 326 273 
<< m1 >>
rect 327 272 328 273 
<< m1 >>
rect 331 272 332 273 
<< m1 >>
rect 10 273 11 274 
<< m1 >>
rect 28 273 29 274 
<< m2 >>
rect 28 273 29 274 
<< m1 >>
rect 37 273 38 274 
<< m1 >>
rect 39 273 40 274 
<< m2 >>
rect 43 273 44 274 
<< m1 >>
rect 44 273 45 274 
<< m2 >>
rect 44 273 45 274 
<< m2 >>
rect 45 273 46 274 
<< m1 >>
rect 46 273 47 274 
<< m2 >>
rect 46 273 47 274 
<< m2c >>
rect 46 273 47 274 
<< m1 >>
rect 46 273 47 274 
<< m2 >>
rect 46 273 47 274 
<< m1 >>
rect 52 273 53 274 
<< m1 >>
rect 57 273 58 274 
<< m1 >>
rect 60 273 61 274 
<< m1 >>
rect 62 273 63 274 
<< m1 >>
rect 64 273 65 274 
<< m1 >>
rect 69 273 70 274 
<< m1 >>
rect 73 273 74 274 
<< m1 >>
rect 116 273 117 274 
<< m1 >>
rect 130 273 131 274 
<< m1 >>
rect 132 273 133 274 
<< m1 >>
rect 134 273 135 274 
<< m1 >>
rect 136 273 137 274 
<< m1 >>
rect 165 273 166 274 
<< m2 >>
rect 166 273 167 274 
<< m1 >>
rect 171 273 172 274 
<< m2 >>
rect 180 273 181 274 
<< m1 >>
rect 181 273 182 274 
<< m2 >>
rect 181 273 182 274 
<< m2 >>
rect 182 273 183 274 
<< m1 >>
rect 183 273 184 274 
<< m2 >>
rect 183 273 184 274 
<< m2c >>
rect 183 273 184 274 
<< m1 >>
rect 183 273 184 274 
<< m2 >>
rect 183 273 184 274 
<< m1 >>
rect 188 273 189 274 
<< m1 >>
rect 190 273 191 274 
<< m1 >>
rect 219 273 220 274 
<< m2 >>
rect 225 273 226 274 
<< m1 >>
rect 226 273 227 274 
<< m2 >>
rect 234 273 235 274 
<< m1 >>
rect 235 273 236 274 
<< m2 >>
rect 239 273 240 274 
<< m2 >>
rect 241 273 242 274 
<< m2 >>
rect 243 273 244 274 
<< m1 >>
rect 253 273 254 274 
<< m2 >>
rect 272 273 273 274 
<< m2 >>
rect 276 273 277 274 
<< m2 >>
rect 278 273 279 274 
<< m2 >>
rect 295 273 296 274 
<< m1 >>
rect 296 273 297 274 
<< m2 >>
rect 296 273 297 274 
<< m2c >>
rect 296 273 297 274 
<< m1 >>
rect 296 273 297 274 
<< m2 >>
rect 296 273 297 274 
<< m1 >>
rect 297 273 298 274 
<< m1 >>
rect 298 273 299 274 
<< m1 >>
rect 299 273 300 274 
<< m1 >>
rect 300 273 301 274 
<< m1 >>
rect 316 273 317 274 
<< m2 >>
rect 316 273 317 274 
<< m1 >>
rect 322 273 323 274 
<< m1 >>
rect 325 273 326 274 
<< m2 >>
rect 325 273 326 274 
<< m1 >>
rect 327 273 328 274 
<< m1 >>
rect 331 273 332 274 
<< m1 >>
rect 10 274 11 275 
<< m1 >>
rect 28 274 29 275 
<< m2 >>
rect 28 274 29 275 
<< m1 >>
rect 37 274 38 275 
<< m1 >>
rect 39 274 40 275 
<< m1 >>
rect 44 274 45 275 
<< m1 >>
rect 46 274 47 275 
<< m1 >>
rect 47 274 48 275 
<< m1 >>
rect 48 274 49 275 
<< m1 >>
rect 49 274 50 275 
<< m1 >>
rect 50 274 51 275 
<< m1 >>
rect 51 274 52 275 
<< m1 >>
rect 52 274 53 275 
<< m1 >>
rect 57 274 58 275 
<< m1 >>
rect 60 274 61 275 
<< m1 >>
rect 62 274 63 275 
<< m1 >>
rect 64 274 65 275 
<< m1 >>
rect 69 274 70 275 
<< m1 >>
rect 73 274 74 275 
<< m1 >>
rect 116 274 117 275 
<< m1 >>
rect 130 274 131 275 
<< m1 >>
rect 132 274 133 275 
<< m1 >>
rect 134 274 135 275 
<< m1 >>
rect 136 274 137 275 
<< m1 >>
rect 165 274 166 275 
<< m2 >>
rect 166 274 167 275 
<< m1 >>
rect 171 274 172 275 
<< m2 >>
rect 180 274 181 275 
<< m1 >>
rect 181 274 182 275 
<< m1 >>
rect 188 274 189 275 
<< m1 >>
rect 190 274 191 275 
<< m1 >>
rect 219 274 220 275 
<< m2 >>
rect 225 274 226 275 
<< m1 >>
rect 226 274 227 275 
<< m2 >>
rect 234 274 235 275 
<< m1 >>
rect 235 274 236 275 
<< m1 >>
rect 236 274 237 275 
<< m1 >>
rect 237 274 238 275 
<< m1 >>
rect 238 274 239 275 
<< m1 >>
rect 239 274 240 275 
<< m2 >>
rect 239 274 240 275 
<< m1 >>
rect 240 274 241 275 
<< m1 >>
rect 241 274 242 275 
<< m2 >>
rect 241 274 242 275 
<< m1 >>
rect 242 274 243 275 
<< m1 >>
rect 243 274 244 275 
<< m2 >>
rect 243 274 244 275 
<< m1 >>
rect 244 274 245 275 
<< m2 >>
rect 244 274 245 275 
<< m1 >>
rect 245 274 246 275 
<< m2 >>
rect 245 274 246 275 
<< m1 >>
rect 246 274 247 275 
<< m2 >>
rect 246 274 247 275 
<< m1 >>
rect 247 274 248 275 
<< m2 >>
rect 247 274 248 275 
<< m1 >>
rect 248 274 249 275 
<< m2 >>
rect 248 274 249 275 
<< m1 >>
rect 249 274 250 275 
<< m1 >>
rect 250 274 251 275 
<< m1 >>
rect 251 274 252 275 
<< m2 >>
rect 251 274 252 275 
<< m2c >>
rect 251 274 252 275 
<< m1 >>
rect 251 274 252 275 
<< m2 >>
rect 251 274 252 275 
<< m2 >>
rect 252 274 253 275 
<< m1 >>
rect 253 274 254 275 
<< m2 >>
rect 253 274 254 275 
<< m1 >>
rect 254 274 255 275 
<< m2 >>
rect 254 274 255 275 
<< m1 >>
rect 255 274 256 275 
<< m2 >>
rect 255 274 256 275 
<< m1 >>
rect 256 274 257 275 
<< m2 >>
rect 256 274 257 275 
<< m1 >>
rect 257 274 258 275 
<< m2 >>
rect 257 274 258 275 
<< m1 >>
rect 258 274 259 275 
<< m2 >>
rect 258 274 259 275 
<< m1 >>
rect 259 274 260 275 
<< m2 >>
rect 259 274 260 275 
<< m1 >>
rect 260 274 261 275 
<< m2 >>
rect 260 274 261 275 
<< m1 >>
rect 261 274 262 275 
<< m2 >>
rect 261 274 262 275 
<< m1 >>
rect 262 274 263 275 
<< m2 >>
rect 262 274 263 275 
<< m1 >>
rect 263 274 264 275 
<< m2 >>
rect 263 274 264 275 
<< m1 >>
rect 264 274 265 275 
<< m2 >>
rect 264 274 265 275 
<< m1 >>
rect 265 274 266 275 
<< m2 >>
rect 265 274 266 275 
<< m1 >>
rect 266 274 267 275 
<< m2 >>
rect 266 274 267 275 
<< m1 >>
rect 267 274 268 275 
<< m2 >>
rect 267 274 268 275 
<< m1 >>
rect 268 274 269 275 
<< m2 >>
rect 268 274 269 275 
<< m2 >>
rect 269 274 270 275 
<< m1 >>
rect 270 274 271 275 
<< m2 >>
rect 270 274 271 275 
<< m2c >>
rect 270 274 271 275 
<< m1 >>
rect 270 274 271 275 
<< m2 >>
rect 270 274 271 275 
<< m1 >>
rect 271 274 272 275 
<< m1 >>
rect 272 274 273 275 
<< m2 >>
rect 272 274 273 275 
<< m1 >>
rect 273 274 274 275 
<< m1 >>
rect 274 274 275 275 
<< m1 >>
rect 275 274 276 275 
<< m1 >>
rect 276 274 277 275 
<< m2 >>
rect 276 274 277 275 
<< m1 >>
rect 277 274 278 275 
<< m1 >>
rect 278 274 279 275 
<< m2 >>
rect 278 274 279 275 
<< m1 >>
rect 279 274 280 275 
<< m1 >>
rect 280 274 281 275 
<< m1 >>
rect 281 274 282 275 
<< m1 >>
rect 282 274 283 275 
<< m1 >>
rect 283 274 284 275 
<< m1 >>
rect 284 274 285 275 
<< m1 >>
rect 285 274 286 275 
<< m1 >>
rect 286 274 287 275 
<< m1 >>
rect 300 274 301 275 
<< m1 >>
rect 316 274 317 275 
<< m2 >>
rect 316 274 317 275 
<< m1 >>
rect 317 274 318 275 
<< m1 >>
rect 318 274 319 275 
<< m1 >>
rect 319 274 320 275 
<< m1 >>
rect 320 274 321 275 
<< m1 >>
rect 321 274 322 275 
<< m1 >>
rect 322 274 323 275 
<< m1 >>
rect 325 274 326 275 
<< m2 >>
rect 325 274 326 275 
<< m1 >>
rect 327 274 328 275 
<< m1 >>
rect 331 274 332 275 
<< m1 >>
rect 10 275 11 276 
<< m1 >>
rect 28 275 29 276 
<< m2 >>
rect 28 275 29 276 
<< m1 >>
rect 37 275 38 276 
<< m1 >>
rect 39 275 40 276 
<< m1 >>
rect 40 275 41 276 
<< m1 >>
rect 41 275 42 276 
<< m1 >>
rect 42 275 43 276 
<< m2 >>
rect 42 275 43 276 
<< m2c >>
rect 42 275 43 276 
<< m1 >>
rect 42 275 43 276 
<< m2 >>
rect 42 275 43 276 
<< m2 >>
rect 43 275 44 276 
<< m1 >>
rect 44 275 45 276 
<< m2 >>
rect 44 275 45 276 
<< m2 >>
rect 45 275 46 276 
<< m2 >>
rect 46 275 47 276 
<< m2 >>
rect 47 275 48 276 
<< m2 >>
rect 48 275 49 276 
<< m2 >>
rect 49 275 50 276 
<< m2 >>
rect 50 275 51 276 
<< m2 >>
rect 51 275 52 276 
<< m2 >>
rect 52 275 53 276 
<< m2 >>
rect 53 275 54 276 
<< m1 >>
rect 54 275 55 276 
<< m2 >>
rect 54 275 55 276 
<< m2c >>
rect 54 275 55 276 
<< m1 >>
rect 54 275 55 276 
<< m2 >>
rect 54 275 55 276 
<< m1 >>
rect 55 275 56 276 
<< m1 >>
rect 57 275 58 276 
<< m1 >>
rect 60 275 61 276 
<< m1 >>
rect 62 275 63 276 
<< m1 >>
rect 64 275 65 276 
<< m1 >>
rect 69 275 70 276 
<< m2 >>
rect 69 275 70 276 
<< m2c >>
rect 69 275 70 276 
<< m1 >>
rect 69 275 70 276 
<< m2 >>
rect 69 275 70 276 
<< m1 >>
rect 73 275 74 276 
<< m1 >>
rect 116 275 117 276 
<< m1 >>
rect 117 275 118 276 
<< m1 >>
rect 118 275 119 276 
<< m1 >>
rect 119 275 120 276 
<< m1 >>
rect 120 275 121 276 
<< m1 >>
rect 121 275 122 276 
<< m1 >>
rect 122 275 123 276 
<< m1 >>
rect 123 275 124 276 
<< m1 >>
rect 124 275 125 276 
<< m1 >>
rect 125 275 126 276 
<< m1 >>
rect 126 275 127 276 
<< m1 >>
rect 127 275 128 276 
<< m1 >>
rect 128 275 129 276 
<< m2 >>
rect 128 275 129 276 
<< m2c >>
rect 128 275 129 276 
<< m1 >>
rect 128 275 129 276 
<< m2 >>
rect 128 275 129 276 
<< m2 >>
rect 129 275 130 276 
<< m1 >>
rect 130 275 131 276 
<< m2 >>
rect 130 275 131 276 
<< m2 >>
rect 131 275 132 276 
<< m1 >>
rect 132 275 133 276 
<< m2 >>
rect 132 275 133 276 
<< m2 >>
rect 133 275 134 276 
<< m1 >>
rect 134 275 135 276 
<< m2 >>
rect 134 275 135 276 
<< m2 >>
rect 135 275 136 276 
<< m1 >>
rect 136 275 137 276 
<< m2 >>
rect 136 275 137 276 
<< m2 >>
rect 137 275 138 276 
<< m1 >>
rect 138 275 139 276 
<< m2 >>
rect 138 275 139 276 
<< m2c >>
rect 138 275 139 276 
<< m1 >>
rect 138 275 139 276 
<< m2 >>
rect 138 275 139 276 
<< m1 >>
rect 139 275 140 276 
<< m1 >>
rect 140 275 141 276 
<< m1 >>
rect 141 275 142 276 
<< m1 >>
rect 142 275 143 276 
<< m2 >>
rect 142 275 143 276 
<< m2c >>
rect 142 275 143 276 
<< m1 >>
rect 142 275 143 276 
<< m2 >>
rect 142 275 143 276 
<< m1 >>
rect 165 275 166 276 
<< m2 >>
rect 166 275 167 276 
<< m1 >>
rect 171 275 172 276 
<< m2 >>
rect 180 275 181 276 
<< m1 >>
rect 181 275 182 276 
<< m1 >>
rect 183 275 184 276 
<< m1 >>
rect 184 275 185 276 
<< m1 >>
rect 185 275 186 276 
<< m1 >>
rect 186 275 187 276 
<< m2 >>
rect 186 275 187 276 
<< m2c >>
rect 186 275 187 276 
<< m1 >>
rect 186 275 187 276 
<< m2 >>
rect 186 275 187 276 
<< m2 >>
rect 187 275 188 276 
<< m1 >>
rect 188 275 189 276 
<< m2 >>
rect 188 275 189 276 
<< m2 >>
rect 189 275 190 276 
<< m1 >>
rect 190 275 191 276 
<< m2 >>
rect 190 275 191 276 
<< m2 >>
rect 191 275 192 276 
<< m1 >>
rect 192 275 193 276 
<< m2 >>
rect 192 275 193 276 
<< m2c >>
rect 192 275 193 276 
<< m1 >>
rect 192 275 193 276 
<< m2 >>
rect 192 275 193 276 
<< m1 >>
rect 193 275 194 276 
<< m1 >>
rect 194 275 195 276 
<< m2 >>
rect 194 275 195 276 
<< m2c >>
rect 194 275 195 276 
<< m1 >>
rect 194 275 195 276 
<< m2 >>
rect 194 275 195 276 
<< m1 >>
rect 219 275 220 276 
<< m2 >>
rect 219 275 220 276 
<< m2c >>
rect 219 275 220 276 
<< m1 >>
rect 219 275 220 276 
<< m2 >>
rect 219 275 220 276 
<< m2 >>
rect 225 275 226 276 
<< m1 >>
rect 226 275 227 276 
<< m1 >>
rect 227 275 228 276 
<< m1 >>
rect 228 275 229 276 
<< m1 >>
rect 229 275 230 276 
<< m1 >>
rect 230 275 231 276 
<< m1 >>
rect 231 275 232 276 
<< m1 >>
rect 232 275 233 276 
<< m2 >>
rect 232 275 233 276 
<< m2c >>
rect 232 275 233 276 
<< m1 >>
rect 232 275 233 276 
<< m2 >>
rect 232 275 233 276 
<< m2 >>
rect 234 275 235 276 
<< m2 >>
rect 239 275 240 276 
<< m2 >>
rect 241 275 242 276 
<< m2 >>
rect 248 275 249 276 
<< m1 >>
rect 268 275 269 276 
<< m2 >>
rect 272 275 273 276 
<< m2 >>
rect 276 275 277 276 
<< m2 >>
rect 278 275 279 276 
<< m1 >>
rect 286 275 287 276 
<< m1 >>
rect 300 275 301 276 
<< m1 >>
rect 301 275 302 276 
<< m1 >>
rect 302 275 303 276 
<< m1 >>
rect 303 275 304 276 
<< m1 >>
rect 304 275 305 276 
<< m1 >>
rect 305 275 306 276 
<< m1 >>
rect 306 275 307 276 
<< m1 >>
rect 307 275 308 276 
<< m1 >>
rect 308 275 309 276 
<< m1 >>
rect 309 275 310 276 
<< m1 >>
rect 310 275 311 276 
<< m1 >>
rect 311 275 312 276 
<< m1 >>
rect 312 275 313 276 
<< m1 >>
rect 313 275 314 276 
<< m1 >>
rect 314 275 315 276 
<< m2 >>
rect 314 275 315 276 
<< m2c >>
rect 314 275 315 276 
<< m1 >>
rect 314 275 315 276 
<< m2 >>
rect 314 275 315 276 
<< m2 >>
rect 316 275 317 276 
<< m1 >>
rect 325 275 326 276 
<< m2 >>
rect 325 275 326 276 
<< m1 >>
rect 327 275 328 276 
<< m1 >>
rect 331 275 332 276 
<< m1 >>
rect 10 276 11 277 
<< m1 >>
rect 28 276 29 277 
<< m2 >>
rect 28 276 29 277 
<< m1 >>
rect 37 276 38 277 
<< m1 >>
rect 44 276 45 277 
<< m1 >>
rect 55 276 56 277 
<< m1 >>
rect 57 276 58 277 
<< m1 >>
rect 60 276 61 277 
<< m1 >>
rect 62 276 63 277 
<< m1 >>
rect 64 276 65 277 
<< m2 >>
rect 66 276 67 277 
<< m2 >>
rect 67 276 68 277 
<< m2 >>
rect 68 276 69 277 
<< m2 >>
rect 69 276 70 277 
<< m1 >>
rect 73 276 74 277 
<< m1 >>
rect 130 276 131 277 
<< m1 >>
rect 132 276 133 277 
<< m1 >>
rect 134 276 135 277 
<< m1 >>
rect 136 276 137 277 
<< m2 >>
rect 142 276 143 277 
<< m1 >>
rect 165 276 166 277 
<< m2 >>
rect 166 276 167 277 
<< m1 >>
rect 171 276 172 277 
<< m2 >>
rect 180 276 181 277 
<< m1 >>
rect 181 276 182 277 
<< m1 >>
rect 183 276 184 277 
<< m1 >>
rect 188 276 189 277 
<< m1 >>
rect 190 276 191 277 
<< m2 >>
rect 194 276 195 277 
<< m2 >>
rect 195 276 196 277 
<< m2 >>
rect 196 276 197 277 
<< m2 >>
rect 197 276 198 277 
<< m2 >>
rect 198 276 199 277 
<< m2 >>
rect 199 276 200 277 
<< m2 >>
rect 200 276 201 277 
<< m2 >>
rect 201 276 202 277 
<< m2 >>
rect 202 276 203 277 
<< m2 >>
rect 203 276 204 277 
<< m2 >>
rect 204 276 205 277 
<< m2 >>
rect 205 276 206 277 
<< m2 >>
rect 206 276 207 277 
<< m2 >>
rect 207 276 208 277 
<< m2 >>
rect 208 276 209 277 
<< m2 >>
rect 209 276 210 277 
<< m2 >>
rect 210 276 211 277 
<< m2 >>
rect 211 276 212 277 
<< m2 >>
rect 212 276 213 277 
<< m2 >>
rect 213 276 214 277 
<< m2 >>
rect 214 276 215 277 
<< m2 >>
rect 215 276 216 277 
<< m2 >>
rect 216 276 217 277 
<< m2 >>
rect 217 276 218 277 
<< m2 >>
rect 219 276 220 277 
<< m2 >>
rect 225 276 226 277 
<< m2 >>
rect 232 276 233 277 
<< m1 >>
rect 234 276 235 277 
<< m2 >>
rect 234 276 235 277 
<< m2c >>
rect 234 276 235 277 
<< m1 >>
rect 234 276 235 277 
<< m2 >>
rect 234 276 235 277 
<< m2 >>
rect 239 276 240 277 
<< m2 >>
rect 241 276 242 277 
<< m2 >>
rect 248 276 249 277 
<< m1 >>
rect 268 276 269 277 
<< m1 >>
rect 272 276 273 277 
<< m2 >>
rect 272 276 273 277 
<< m2c >>
rect 272 276 273 277 
<< m1 >>
rect 272 276 273 277 
<< m2 >>
rect 272 276 273 277 
<< m2 >>
rect 276 276 277 277 
<< m2 >>
rect 278 276 279 277 
<< m1 >>
rect 286 276 287 277 
<< m2 >>
rect 314 276 315 277 
<< m2 >>
rect 316 276 317 277 
<< m1 >>
rect 325 276 326 277 
<< m2 >>
rect 325 276 326 277 
<< m1 >>
rect 327 276 328 277 
<< m1 >>
rect 331 276 332 277 
<< m1 >>
rect 10 277 11 278 
<< m1 >>
rect 28 277 29 278 
<< m2 >>
rect 28 277 29 278 
<< m1 >>
rect 37 277 38 278 
<< m1 >>
rect 44 277 45 278 
<< m1 >>
rect 55 277 56 278 
<< m1 >>
rect 57 277 58 278 
<< m1 >>
rect 60 277 61 278 
<< m1 >>
rect 62 277 63 278 
<< m1 >>
rect 64 277 65 278 
<< m1 >>
rect 65 277 66 278 
<< m1 >>
rect 66 277 67 278 
<< m2 >>
rect 66 277 67 278 
<< m1 >>
rect 67 277 68 278 
<< m1 >>
rect 68 277 69 278 
<< m1 >>
rect 69 277 70 278 
<< m1 >>
rect 70 277 71 278 
<< m1 >>
rect 71 277 72 278 
<< m2 >>
rect 71 277 72 278 
<< m2c >>
rect 71 277 72 278 
<< m1 >>
rect 71 277 72 278 
<< m2 >>
rect 71 277 72 278 
<< m2 >>
rect 72 277 73 278 
<< m1 >>
rect 73 277 74 278 
<< m2 >>
rect 73 277 74 278 
<< m2 >>
rect 74 277 75 278 
<< m1 >>
rect 75 277 76 278 
<< m2 >>
rect 75 277 76 278 
<< m2c >>
rect 75 277 76 278 
<< m1 >>
rect 75 277 76 278 
<< m2 >>
rect 75 277 76 278 
<< m1 >>
rect 76 277 77 278 
<< m1 >>
rect 77 277 78 278 
<< m1 >>
rect 78 277 79 278 
<< m1 >>
rect 79 277 80 278 
<< m1 >>
rect 80 277 81 278 
<< m1 >>
rect 81 277 82 278 
<< m1 >>
rect 82 277 83 278 
<< m1 >>
rect 83 277 84 278 
<< m1 >>
rect 84 277 85 278 
<< m1 >>
rect 85 277 86 278 
<< m1 >>
rect 86 277 87 278 
<< m1 >>
rect 87 277 88 278 
<< m1 >>
rect 88 277 89 278 
<< m1 >>
rect 89 277 90 278 
<< m1 >>
rect 90 277 91 278 
<< m1 >>
rect 91 277 92 278 
<< m1 >>
rect 92 277 93 278 
<< m1 >>
rect 93 277 94 278 
<< m1 >>
rect 94 277 95 278 
<< m1 >>
rect 95 277 96 278 
<< m1 >>
rect 96 277 97 278 
<< m1 >>
rect 97 277 98 278 
<< m1 >>
rect 98 277 99 278 
<< m1 >>
rect 99 277 100 278 
<< m1 >>
rect 100 277 101 278 
<< m1 >>
rect 101 277 102 278 
<< m1 >>
rect 102 277 103 278 
<< m1 >>
rect 103 277 104 278 
<< m1 >>
rect 104 277 105 278 
<< m1 >>
rect 105 277 106 278 
<< m1 >>
rect 106 277 107 278 
<< m1 >>
rect 107 277 108 278 
<< m1 >>
rect 108 277 109 278 
<< m1 >>
rect 109 277 110 278 
<< m1 >>
rect 110 277 111 278 
<< m1 >>
rect 111 277 112 278 
<< m1 >>
rect 112 277 113 278 
<< m1 >>
rect 113 277 114 278 
<< m1 >>
rect 114 277 115 278 
<< m1 >>
rect 115 277 116 278 
<< m1 >>
rect 116 277 117 278 
<< m1 >>
rect 117 277 118 278 
<< m1 >>
rect 118 277 119 278 
<< m1 >>
rect 130 277 131 278 
<< m2 >>
rect 130 277 131 278 
<< m2c >>
rect 130 277 131 278 
<< m1 >>
rect 130 277 131 278 
<< m2 >>
rect 130 277 131 278 
<< m2 >>
rect 131 277 132 278 
<< m1 >>
rect 132 277 133 278 
<< m2 >>
rect 132 277 133 278 
<< m2 >>
rect 133 277 134 278 
<< m1 >>
rect 134 277 135 278 
<< m2 >>
rect 134 277 135 278 
<< m2 >>
rect 135 277 136 278 
<< m1 >>
rect 136 277 137 278 
<< m2 >>
rect 136 277 137 278 
<< m2 >>
rect 137 277 138 278 
<< m1 >>
rect 138 277 139 278 
<< m2 >>
rect 138 277 139 278 
<< m2c >>
rect 138 277 139 278 
<< m1 >>
rect 138 277 139 278 
<< m2 >>
rect 138 277 139 278 
<< m1 >>
rect 139 277 140 278 
<< m1 >>
rect 140 277 141 278 
<< m1 >>
rect 141 277 142 278 
<< m1 >>
rect 142 277 143 278 
<< m2 >>
rect 142 277 143 278 
<< m1 >>
rect 143 277 144 278 
<< m1 >>
rect 144 277 145 278 
<< m1 >>
rect 145 277 146 278 
<< m1 >>
rect 146 277 147 278 
<< m1 >>
rect 147 277 148 278 
<< m1 >>
rect 148 277 149 278 
<< m1 >>
rect 149 277 150 278 
<< m1 >>
rect 150 277 151 278 
<< m1 >>
rect 151 277 152 278 
<< m1 >>
rect 152 277 153 278 
<< m1 >>
rect 153 277 154 278 
<< m1 >>
rect 154 277 155 278 
<< m1 >>
rect 155 277 156 278 
<< m1 >>
rect 156 277 157 278 
<< m1 >>
rect 157 277 158 278 
<< m1 >>
rect 158 277 159 278 
<< m1 >>
rect 159 277 160 278 
<< m1 >>
rect 160 277 161 278 
<< m1 >>
rect 161 277 162 278 
<< m1 >>
rect 162 277 163 278 
<< m1 >>
rect 163 277 164 278 
<< m1 >>
rect 165 277 166 278 
<< m2 >>
rect 166 277 167 278 
<< m1 >>
rect 171 277 172 278 
<< m1 >>
rect 173 277 174 278 
<< m1 >>
rect 174 277 175 278 
<< m1 >>
rect 175 277 176 278 
<< m1 >>
rect 176 277 177 278 
<< m1 >>
rect 177 277 178 278 
<< m1 >>
rect 178 277 179 278 
<< m1 >>
rect 179 277 180 278 
<< m2 >>
rect 179 277 180 278 
<< m2c >>
rect 179 277 180 278 
<< m1 >>
rect 179 277 180 278 
<< m2 >>
rect 179 277 180 278 
<< m2 >>
rect 180 277 181 278 
<< m1 >>
rect 181 277 182 278 
<< m1 >>
rect 183 277 184 278 
<< m1 >>
rect 188 277 189 278 
<< m2 >>
rect 188 277 189 278 
<< m2c >>
rect 188 277 189 278 
<< m1 >>
rect 188 277 189 278 
<< m2 >>
rect 188 277 189 278 
<< m2 >>
rect 189 277 190 278 
<< m1 >>
rect 190 277 191 278 
<< m2 >>
rect 190 277 191 278 
<< m2 >>
rect 191 277 192 278 
<< m1 >>
rect 192 277 193 278 
<< m2 >>
rect 192 277 193 278 
<< m2c >>
rect 192 277 193 278 
<< m1 >>
rect 192 277 193 278 
<< m2 >>
rect 192 277 193 278 
<< m1 >>
rect 193 277 194 278 
<< m1 >>
rect 194 277 195 278 
<< m1 >>
rect 195 277 196 278 
<< m1 >>
rect 196 277 197 278 
<< m1 >>
rect 197 277 198 278 
<< m1 >>
rect 199 277 200 278 
<< m1 >>
rect 200 277 201 278 
<< m1 >>
rect 201 277 202 278 
<< m1 >>
rect 202 277 203 278 
<< m1 >>
rect 203 277 204 278 
<< m1 >>
rect 204 277 205 278 
<< m1 >>
rect 205 277 206 278 
<< m1 >>
rect 206 277 207 278 
<< m1 >>
rect 207 277 208 278 
<< m1 >>
rect 208 277 209 278 
<< m1 >>
rect 209 277 210 278 
<< m1 >>
rect 210 277 211 278 
<< m1 >>
rect 211 277 212 278 
<< m1 >>
rect 212 277 213 278 
<< m1 >>
rect 213 277 214 278 
<< m1 >>
rect 214 277 215 278 
<< m1 >>
rect 215 277 216 278 
<< m1 >>
rect 216 277 217 278 
<< m1 >>
rect 217 277 218 278 
<< m2 >>
rect 217 277 218 278 
<< m1 >>
rect 218 277 219 278 
<< m1 >>
rect 219 277 220 278 
<< m2 >>
rect 219 277 220 278 
<< m1 >>
rect 220 277 221 278 
<< m1 >>
rect 221 277 222 278 
<< m1 >>
rect 222 277 223 278 
<< m1 >>
rect 223 277 224 278 
<< m1 >>
rect 224 277 225 278 
<< m1 >>
rect 225 277 226 278 
<< m2 >>
rect 225 277 226 278 
<< m1 >>
rect 226 277 227 278 
<< m1 >>
rect 227 277 228 278 
<< m1 >>
rect 228 277 229 278 
<< m1 >>
rect 229 277 230 278 
<< m1 >>
rect 230 277 231 278 
<< m1 >>
rect 231 277 232 278 
<< m1 >>
rect 232 277 233 278 
<< m2 >>
rect 232 277 233 278 
<< m1 >>
rect 233 277 234 278 
<< m1 >>
rect 234 277 235 278 
<< m1 >>
rect 237 277 238 278 
<< m1 >>
rect 238 277 239 278 
<< m1 >>
rect 239 277 240 278 
<< m2 >>
rect 239 277 240 278 
<< m1 >>
rect 240 277 241 278 
<< m1 >>
rect 241 277 242 278 
<< m2 >>
rect 241 277 242 278 
<< m1 >>
rect 242 277 243 278 
<< m1 >>
rect 243 277 244 278 
<< m1 >>
rect 244 277 245 278 
<< m1 >>
rect 245 277 246 278 
<< m1 >>
rect 246 277 247 278 
<< m1 >>
rect 247 277 248 278 
<< m1 >>
rect 248 277 249 278 
<< m2 >>
rect 248 277 249 278 
<< m1 >>
rect 249 277 250 278 
<< m1 >>
rect 250 277 251 278 
<< m1 >>
rect 251 277 252 278 
<< m1 >>
rect 252 277 253 278 
<< m1 >>
rect 253 277 254 278 
<< m1 >>
rect 254 277 255 278 
<< m1 >>
rect 255 277 256 278 
<< m1 >>
rect 256 277 257 278 
<< m1 >>
rect 257 277 258 278 
<< m1 >>
rect 258 277 259 278 
<< m1 >>
rect 259 277 260 278 
<< m1 >>
rect 260 277 261 278 
<< m1 >>
rect 261 277 262 278 
<< m1 >>
rect 262 277 263 278 
<< m1 >>
rect 263 277 264 278 
<< m1 >>
rect 264 277 265 278 
<< m1 >>
rect 265 277 266 278 
<< m1 >>
rect 266 277 267 278 
<< m2 >>
rect 266 277 267 278 
<< m2c >>
rect 266 277 267 278 
<< m1 >>
rect 266 277 267 278 
<< m2 >>
rect 266 277 267 278 
<< m2 >>
rect 267 277 268 278 
<< m1 >>
rect 268 277 269 278 
<< m2 >>
rect 268 277 269 278 
<< m2 >>
rect 269 277 270 278 
<< m1 >>
rect 270 277 271 278 
<< m2 >>
rect 270 277 271 278 
<< m2c >>
rect 270 277 271 278 
<< m1 >>
rect 270 277 271 278 
<< m2 >>
rect 270 277 271 278 
<< m1 >>
rect 272 277 273 278 
<< m1 >>
rect 274 277 275 278 
<< m1 >>
rect 275 277 276 278 
<< m1 >>
rect 276 277 277 278 
<< m2 >>
rect 276 277 277 278 
<< m1 >>
rect 277 277 278 278 
<< m1 >>
rect 278 277 279 278 
<< m2 >>
rect 278 277 279 278 
<< m1 >>
rect 279 277 280 278 
<< m1 >>
rect 280 277 281 278 
<< m1 >>
rect 281 277 282 278 
<< m1 >>
rect 282 277 283 278 
<< m1 >>
rect 283 277 284 278 
<< m1 >>
rect 284 277 285 278 
<< m2 >>
rect 284 277 285 278 
<< m2c >>
rect 284 277 285 278 
<< m1 >>
rect 284 277 285 278 
<< m2 >>
rect 284 277 285 278 
<< m2 >>
rect 285 277 286 278 
<< m1 >>
rect 286 277 287 278 
<< m2 >>
rect 286 277 287 278 
<< m2 >>
rect 287 277 288 278 
<< m1 >>
rect 288 277 289 278 
<< m2 >>
rect 288 277 289 278 
<< m2c >>
rect 288 277 289 278 
<< m1 >>
rect 288 277 289 278 
<< m2 >>
rect 288 277 289 278 
<< m1 >>
rect 289 277 290 278 
<< m1 >>
rect 290 277 291 278 
<< m1 >>
rect 291 277 292 278 
<< m1 >>
rect 292 277 293 278 
<< m1 >>
rect 293 277 294 278 
<< m1 >>
rect 294 277 295 278 
<< m1 >>
rect 295 277 296 278 
<< m1 >>
rect 296 277 297 278 
<< m1 >>
rect 297 277 298 278 
<< m1 >>
rect 298 277 299 278 
<< m1 >>
rect 299 277 300 278 
<< m1 >>
rect 300 277 301 278 
<< m1 >>
rect 301 277 302 278 
<< m1 >>
rect 302 277 303 278 
<< m1 >>
rect 303 277 304 278 
<< m1 >>
rect 304 277 305 278 
<< m1 >>
rect 305 277 306 278 
<< m1 >>
rect 306 277 307 278 
<< m1 >>
rect 307 277 308 278 
<< m1 >>
rect 308 277 309 278 
<< m1 >>
rect 309 277 310 278 
<< m1 >>
rect 310 277 311 278 
<< m1 >>
rect 311 277 312 278 
<< m1 >>
rect 312 277 313 278 
<< m1 >>
rect 313 277 314 278 
<< m1 >>
rect 314 277 315 278 
<< m2 >>
rect 314 277 315 278 
<< m1 >>
rect 315 277 316 278 
<< m1 >>
rect 316 277 317 278 
<< m2 >>
rect 316 277 317 278 
<< m1 >>
rect 317 277 318 278 
<< m1 >>
rect 318 277 319 278 
<< m1 >>
rect 319 277 320 278 
<< m1 >>
rect 320 277 321 278 
<< m1 >>
rect 321 277 322 278 
<< m1 >>
rect 322 277 323 278 
<< m1 >>
rect 323 277 324 278 
<< m1 >>
rect 324 277 325 278 
<< m1 >>
rect 325 277 326 278 
<< m2 >>
rect 325 277 326 278 
<< m1 >>
rect 327 277 328 278 
<< m1 >>
rect 331 277 332 278 
<< m1 >>
rect 10 278 11 279 
<< m1 >>
rect 28 278 29 279 
<< m2 >>
rect 28 278 29 279 
<< m1 >>
rect 37 278 38 279 
<< m1 >>
rect 44 278 45 279 
<< m1 >>
rect 55 278 56 279 
<< m1 >>
rect 57 278 58 279 
<< m1 >>
rect 60 278 61 279 
<< m1 >>
rect 62 278 63 279 
<< m2 >>
rect 66 278 67 279 
<< m1 >>
rect 73 278 74 279 
<< m1 >>
rect 118 278 119 279 
<< m1 >>
rect 132 278 133 279 
<< m1 >>
rect 134 278 135 279 
<< m1 >>
rect 136 278 137 279 
<< m2 >>
rect 142 278 143 279 
<< m1 >>
rect 163 278 164 279 
<< m1 >>
rect 165 278 166 279 
<< m2 >>
rect 166 278 167 279 
<< m1 >>
rect 171 278 172 279 
<< m1 >>
rect 173 278 174 279 
<< m1 >>
rect 181 278 182 279 
<< m1 >>
rect 183 278 184 279 
<< m1 >>
rect 190 278 191 279 
<< m1 >>
rect 197 278 198 279 
<< m1 >>
rect 199 278 200 279 
<< m2 >>
rect 217 278 218 279 
<< m2 >>
rect 219 278 220 279 
<< m2 >>
rect 225 278 226 279 
<< m2 >>
rect 232 278 233 279 
<< m2 >>
rect 233 278 234 279 
<< m2 >>
rect 234 278 235 279 
<< m2 >>
rect 235 278 236 279 
<< m1 >>
rect 237 278 238 279 
<< m2 >>
rect 239 278 240 279 
<< m2 >>
rect 241 278 242 279 
<< m2 >>
rect 248 278 249 279 
<< m1 >>
rect 268 278 269 279 
<< m1 >>
rect 270 278 271 279 
<< m2 >>
rect 270 278 271 279 
<< m2 >>
rect 271 278 272 279 
<< m1 >>
rect 272 278 273 279 
<< m2 >>
rect 272 278 273 279 
<< m2 >>
rect 273 278 274 279 
<< m1 >>
rect 274 278 275 279 
<< m2 >>
rect 274 278 275 279 
<< m2c >>
rect 274 278 275 279 
<< m1 >>
rect 274 278 275 279 
<< m2 >>
rect 274 278 275 279 
<< m2 >>
rect 276 278 277 279 
<< m2 >>
rect 278 278 279 279 
<< m1 >>
rect 286 278 287 279 
<< m2 >>
rect 314 278 315 279 
<< m2 >>
rect 316 278 317 279 
<< m2 >>
rect 325 278 326 279 
<< m1 >>
rect 327 278 328 279 
<< m1 >>
rect 331 278 332 279 
<< m1 >>
rect 10 279 11 280 
<< m1 >>
rect 28 279 29 280 
<< m2 >>
rect 28 279 29 280 
<< m1 >>
rect 37 279 38 280 
<< m1 >>
rect 44 279 45 280 
<< m1 >>
rect 55 279 56 280 
<< m1 >>
rect 57 279 58 280 
<< m1 >>
rect 60 279 61 280 
<< m1 >>
rect 62 279 63 280 
<< m1 >>
rect 64 279 65 280 
<< m1 >>
rect 65 279 66 280 
<< m1 >>
rect 66 279 67 280 
<< m2 >>
rect 66 279 67 280 
<< m2c >>
rect 66 279 67 280 
<< m1 >>
rect 66 279 67 280 
<< m2 >>
rect 66 279 67 280 
<< m1 >>
rect 73 279 74 280 
<< m1 >>
rect 118 279 119 280 
<< m1 >>
rect 132 279 133 280 
<< m1 >>
rect 134 279 135 280 
<< m1 >>
rect 136 279 137 280 
<< m1 >>
rect 142 279 143 280 
<< m2 >>
rect 142 279 143 280 
<< m2c >>
rect 142 279 143 280 
<< m1 >>
rect 142 279 143 280 
<< m2 >>
rect 142 279 143 280 
<< m1 >>
rect 163 279 164 280 
<< m1 >>
rect 165 279 166 280 
<< m2 >>
rect 166 279 167 280 
<< m1 >>
rect 171 279 172 280 
<< m1 >>
rect 173 279 174 280 
<< m1 >>
rect 181 279 182 280 
<< m1 >>
rect 183 279 184 280 
<< m1 >>
rect 190 279 191 280 
<< m1 >>
rect 197 279 198 280 
<< m1 >>
rect 199 279 200 280 
<< m2 >>
rect 217 279 218 280 
<< m2 >>
rect 219 279 220 280 
<< m2 >>
rect 225 279 226 280 
<< m1 >>
rect 235 279 236 280 
<< m2 >>
rect 235 279 236 280 
<< m2c >>
rect 235 279 236 280 
<< m1 >>
rect 235 279 236 280 
<< m2 >>
rect 235 279 236 280 
<< m1 >>
rect 237 279 238 280 
<< m1 >>
rect 239 279 240 280 
<< m2 >>
rect 239 279 240 280 
<< m2c >>
rect 239 279 240 280 
<< m1 >>
rect 239 279 240 280 
<< m2 >>
rect 239 279 240 280 
<< m1 >>
rect 241 279 242 280 
<< m2 >>
rect 241 279 242 280 
<< m2c >>
rect 241 279 242 280 
<< m1 >>
rect 241 279 242 280 
<< m2 >>
rect 241 279 242 280 
<< m1 >>
rect 248 279 249 280 
<< m2 >>
rect 248 279 249 280 
<< m2c >>
rect 248 279 249 280 
<< m1 >>
rect 248 279 249 280 
<< m2 >>
rect 248 279 249 280 
<< m1 >>
rect 249 279 250 280 
<< m1 >>
rect 250 279 251 280 
<< m1 >>
rect 268 279 269 280 
<< m1 >>
rect 272 279 273 280 
<< m1 >>
rect 276 279 277 280 
<< m2 >>
rect 276 279 277 280 
<< m2c >>
rect 276 279 277 280 
<< m1 >>
rect 276 279 277 280 
<< m2 >>
rect 276 279 277 280 
<< m1 >>
rect 278 279 279 280 
<< m2 >>
rect 278 279 279 280 
<< m2c >>
rect 278 279 279 280 
<< m1 >>
rect 278 279 279 280 
<< m2 >>
rect 278 279 279 280 
<< m1 >>
rect 286 279 287 280 
<< m1 >>
rect 314 279 315 280 
<< m2 >>
rect 314 279 315 280 
<< m2c >>
rect 314 279 315 280 
<< m1 >>
rect 314 279 315 280 
<< m2 >>
rect 314 279 315 280 
<< m1 >>
rect 316 279 317 280 
<< m2 >>
rect 316 279 317 280 
<< m2c >>
rect 316 279 317 280 
<< m1 >>
rect 316 279 317 280 
<< m2 >>
rect 316 279 317 280 
<< m1 >>
rect 325 279 326 280 
<< m2 >>
rect 325 279 326 280 
<< m2c >>
rect 325 279 326 280 
<< m1 >>
rect 325 279 326 280 
<< m2 >>
rect 325 279 326 280 
<< m1 >>
rect 327 279 328 280 
<< m1 >>
rect 331 279 332 280 
<< m1 >>
rect 10 280 11 281 
<< m1 >>
rect 28 280 29 281 
<< m2 >>
rect 28 280 29 281 
<< m1 >>
rect 37 280 38 281 
<< m1 >>
rect 44 280 45 281 
<< m1 >>
rect 55 280 56 281 
<< m1 >>
rect 57 280 58 281 
<< m1 >>
rect 60 280 61 281 
<< m1 >>
rect 62 280 63 281 
<< m1 >>
rect 64 280 65 281 
<< m1 >>
rect 73 280 74 281 
<< m1 >>
rect 118 280 119 281 
<< m1 >>
rect 132 280 133 281 
<< m1 >>
rect 134 280 135 281 
<< m1 >>
rect 136 280 137 281 
<< m1 >>
rect 142 280 143 281 
<< m1 >>
rect 163 280 164 281 
<< m1 >>
rect 165 280 166 281 
<< m2 >>
rect 166 280 167 281 
<< m1 >>
rect 171 280 172 281 
<< m2 >>
rect 172 280 173 281 
<< m1 >>
rect 173 280 174 281 
<< m2 >>
rect 173 280 174 281 
<< m2c >>
rect 173 280 174 281 
<< m1 >>
rect 173 280 174 281 
<< m2 >>
rect 173 280 174 281 
<< m1 >>
rect 181 280 182 281 
<< m1 >>
rect 183 280 184 281 
<< m1 >>
rect 190 280 191 281 
<< m1 >>
rect 197 280 198 281 
<< m2 >>
rect 197 280 198 281 
<< m2c >>
rect 197 280 198 281 
<< m1 >>
rect 197 280 198 281 
<< m2 >>
rect 197 280 198 281 
<< m2 >>
rect 198 280 199 281 
<< m1 >>
rect 199 280 200 281 
<< m2 >>
rect 199 280 200 281 
<< m2 >>
rect 200 280 201 281 
<< m1 >>
rect 214 280 215 281 
<< m1 >>
rect 215 280 216 281 
<< m1 >>
rect 216 280 217 281 
<< m1 >>
rect 217 280 218 281 
<< m2 >>
rect 217 280 218 281 
<< m1 >>
rect 218 280 219 281 
<< m1 >>
rect 219 280 220 281 
<< m2 >>
rect 219 280 220 281 
<< m1 >>
rect 220 280 221 281 
<< m1 >>
rect 221 280 222 281 
<< m1 >>
rect 222 280 223 281 
<< m1 >>
rect 223 280 224 281 
<< m1 >>
rect 224 280 225 281 
<< m2 >>
rect 224 280 225 281 
<< m2c >>
rect 224 280 225 281 
<< m1 >>
rect 224 280 225 281 
<< m2 >>
rect 224 280 225 281 
<< m2 >>
rect 225 280 226 281 
<< m1 >>
rect 226 280 227 281 
<< m1 >>
rect 227 280 228 281 
<< m1 >>
rect 228 280 229 281 
<< m1 >>
rect 229 280 230 281 
<< m1 >>
rect 235 280 236 281 
<< m1 >>
rect 237 280 238 281 
<< m1 >>
rect 239 280 240 281 
<< m1 >>
rect 241 280 242 281 
<< m1 >>
rect 250 280 251 281 
<< m1 >>
rect 268 280 269 281 
<< m1 >>
rect 272 280 273 281 
<< m1 >>
rect 276 280 277 281 
<< m1 >>
rect 278 280 279 281 
<< m1 >>
rect 286 280 287 281 
<< m1 >>
rect 314 280 315 281 
<< m1 >>
rect 316 280 317 281 
<< m1 >>
rect 325 280 326 281 
<< m1 >>
rect 327 280 328 281 
<< m1 >>
rect 331 280 332 281 
<< m1 >>
rect 10 281 11 282 
<< m1 >>
rect 28 281 29 282 
<< m2 >>
rect 28 281 29 282 
<< m1 >>
rect 37 281 38 282 
<< m1 >>
rect 44 281 45 282 
<< m1 >>
rect 55 281 56 282 
<< m1 >>
rect 57 281 58 282 
<< m1 >>
rect 60 281 61 282 
<< m1 >>
rect 62 281 63 282 
<< m1 >>
rect 64 281 65 282 
<< m1 >>
rect 73 281 74 282 
<< m1 >>
rect 118 281 119 282 
<< m1 >>
rect 132 281 133 282 
<< m1 >>
rect 134 281 135 282 
<< m1 >>
rect 136 281 137 282 
<< m1 >>
rect 142 281 143 282 
<< m1 >>
rect 163 281 164 282 
<< m1 >>
rect 165 281 166 282 
<< m2 >>
rect 166 281 167 282 
<< m1 >>
rect 171 281 172 282 
<< m2 >>
rect 172 281 173 282 
<< m1 >>
rect 181 281 182 282 
<< m1 >>
rect 183 281 184 282 
<< m1 >>
rect 190 281 191 282 
<< m1 >>
rect 199 281 200 282 
<< m2 >>
rect 200 281 201 282 
<< m1 >>
rect 214 281 215 282 
<< m2 >>
rect 217 281 218 282 
<< m2 >>
rect 219 281 220 282 
<< m1 >>
rect 226 281 227 282 
<< m1 >>
rect 229 281 230 282 
<< m1 >>
rect 235 281 236 282 
<< m1 >>
rect 237 281 238 282 
<< m1 >>
rect 239 281 240 282 
<< m1 >>
rect 241 281 242 282 
<< m1 >>
rect 250 281 251 282 
<< m1 >>
rect 268 281 269 282 
<< m1 >>
rect 272 281 273 282 
<< m1 >>
rect 276 281 277 282 
<< m1 >>
rect 278 281 279 282 
<< m1 >>
rect 286 281 287 282 
<< m1 >>
rect 314 281 315 282 
<< m1 >>
rect 316 281 317 282 
<< m1 >>
rect 325 281 326 282 
<< m1 >>
rect 327 281 328 282 
<< m1 >>
rect 331 281 332 282 
<< m1 >>
rect 10 282 11 283 
<< pdiffusion >>
rect 12 282 13 283 
<< pdiffusion >>
rect 13 282 14 283 
<< pdiffusion >>
rect 14 282 15 283 
<< pdiffusion >>
rect 15 282 16 283 
<< pdiffusion >>
rect 16 282 17 283 
<< pdiffusion >>
rect 17 282 18 283 
<< m1 >>
rect 28 282 29 283 
<< m2 >>
rect 28 282 29 283 
<< pdiffusion >>
rect 30 282 31 283 
<< pdiffusion >>
rect 31 282 32 283 
<< pdiffusion >>
rect 32 282 33 283 
<< pdiffusion >>
rect 33 282 34 283 
<< pdiffusion >>
rect 34 282 35 283 
<< pdiffusion >>
rect 35 282 36 283 
<< m1 >>
rect 37 282 38 283 
<< m1 >>
rect 44 282 45 283 
<< pdiffusion >>
rect 48 282 49 283 
<< pdiffusion >>
rect 49 282 50 283 
<< pdiffusion >>
rect 50 282 51 283 
<< pdiffusion >>
rect 51 282 52 283 
<< pdiffusion >>
rect 52 282 53 283 
<< pdiffusion >>
rect 53 282 54 283 
<< m1 >>
rect 55 282 56 283 
<< m1 >>
rect 57 282 58 283 
<< m1 >>
rect 60 282 61 283 
<< m1 >>
rect 62 282 63 283 
<< m1 >>
rect 64 282 65 283 
<< pdiffusion >>
rect 66 282 67 283 
<< pdiffusion >>
rect 67 282 68 283 
<< pdiffusion >>
rect 68 282 69 283 
<< pdiffusion >>
rect 69 282 70 283 
<< pdiffusion >>
rect 70 282 71 283 
<< pdiffusion >>
rect 71 282 72 283 
<< m1 >>
rect 73 282 74 283 
<< pdiffusion >>
rect 84 282 85 283 
<< pdiffusion >>
rect 85 282 86 283 
<< pdiffusion >>
rect 86 282 87 283 
<< pdiffusion >>
rect 87 282 88 283 
<< pdiffusion >>
rect 88 282 89 283 
<< pdiffusion >>
rect 89 282 90 283 
<< pdiffusion >>
rect 102 282 103 283 
<< pdiffusion >>
rect 103 282 104 283 
<< pdiffusion >>
rect 104 282 105 283 
<< pdiffusion >>
rect 105 282 106 283 
<< pdiffusion >>
rect 106 282 107 283 
<< pdiffusion >>
rect 107 282 108 283 
<< m1 >>
rect 118 282 119 283 
<< pdiffusion >>
rect 120 282 121 283 
<< pdiffusion >>
rect 121 282 122 283 
<< pdiffusion >>
rect 122 282 123 283 
<< pdiffusion >>
rect 123 282 124 283 
<< pdiffusion >>
rect 124 282 125 283 
<< pdiffusion >>
rect 125 282 126 283 
<< m1 >>
rect 132 282 133 283 
<< m1 >>
rect 134 282 135 283 
<< m1 >>
rect 136 282 137 283 
<< pdiffusion >>
rect 138 282 139 283 
<< pdiffusion >>
rect 139 282 140 283 
<< pdiffusion >>
rect 140 282 141 283 
<< pdiffusion >>
rect 141 282 142 283 
<< m1 >>
rect 142 282 143 283 
<< pdiffusion >>
rect 142 282 143 283 
<< pdiffusion >>
rect 143 282 144 283 
<< pdiffusion >>
rect 156 282 157 283 
<< pdiffusion >>
rect 157 282 158 283 
<< pdiffusion >>
rect 158 282 159 283 
<< pdiffusion >>
rect 159 282 160 283 
<< pdiffusion >>
rect 160 282 161 283 
<< pdiffusion >>
rect 161 282 162 283 
<< m1 >>
rect 163 282 164 283 
<< m1 >>
rect 165 282 166 283 
<< m2 >>
rect 166 282 167 283 
<< m1 >>
rect 171 282 172 283 
<< m2 >>
rect 172 282 173 283 
<< pdiffusion >>
rect 174 282 175 283 
<< pdiffusion >>
rect 175 282 176 283 
<< pdiffusion >>
rect 176 282 177 283 
<< pdiffusion >>
rect 177 282 178 283 
<< pdiffusion >>
rect 178 282 179 283 
<< pdiffusion >>
rect 179 282 180 283 
<< m1 >>
rect 181 282 182 283 
<< m1 >>
rect 183 282 184 283 
<< m1 >>
rect 190 282 191 283 
<< pdiffusion >>
rect 192 282 193 283 
<< pdiffusion >>
rect 193 282 194 283 
<< pdiffusion >>
rect 194 282 195 283 
<< pdiffusion >>
rect 195 282 196 283 
<< pdiffusion >>
rect 196 282 197 283 
<< pdiffusion >>
rect 197 282 198 283 
<< m1 >>
rect 199 282 200 283 
<< m2 >>
rect 200 282 201 283 
<< pdiffusion >>
rect 210 282 211 283 
<< pdiffusion >>
rect 211 282 212 283 
<< pdiffusion >>
rect 212 282 213 283 
<< pdiffusion >>
rect 213 282 214 283 
<< m1 >>
rect 214 282 215 283 
<< pdiffusion >>
rect 214 282 215 283 
<< pdiffusion >>
rect 215 282 216 283 
<< m1 >>
rect 217 282 218 283 
<< m2 >>
rect 217 282 218 283 
<< m2c >>
rect 217 282 218 283 
<< m1 >>
rect 217 282 218 283 
<< m2 >>
rect 217 282 218 283 
<< m1 >>
rect 219 282 220 283 
<< m2 >>
rect 219 282 220 283 
<< m2c >>
rect 219 282 220 283 
<< m1 >>
rect 219 282 220 283 
<< m2 >>
rect 219 282 220 283 
<< m1 >>
rect 220 282 221 283 
<< m1 >>
rect 221 282 222 283 
<< m1 >>
rect 222 282 223 283 
<< m1 >>
rect 223 282 224 283 
<< m1 >>
rect 226 282 227 283 
<< pdiffusion >>
rect 228 282 229 283 
<< m1 >>
rect 229 282 230 283 
<< pdiffusion >>
rect 229 282 230 283 
<< pdiffusion >>
rect 230 282 231 283 
<< pdiffusion >>
rect 231 282 232 283 
<< pdiffusion >>
rect 232 282 233 283 
<< pdiffusion >>
rect 233 282 234 283 
<< m1 >>
rect 235 282 236 283 
<< m1 >>
rect 237 282 238 283 
<< m1 >>
rect 239 282 240 283 
<< m1 >>
rect 241 282 242 283 
<< pdiffusion >>
rect 246 282 247 283 
<< pdiffusion >>
rect 247 282 248 283 
<< pdiffusion >>
rect 248 282 249 283 
<< pdiffusion >>
rect 249 282 250 283 
<< m1 >>
rect 250 282 251 283 
<< pdiffusion >>
rect 250 282 251 283 
<< pdiffusion >>
rect 251 282 252 283 
<< pdiffusion >>
rect 264 282 265 283 
<< pdiffusion >>
rect 265 282 266 283 
<< pdiffusion >>
rect 266 282 267 283 
<< pdiffusion >>
rect 267 282 268 283 
<< m1 >>
rect 268 282 269 283 
<< pdiffusion >>
rect 268 282 269 283 
<< pdiffusion >>
rect 269 282 270 283 
<< m1 >>
rect 272 282 273 283 
<< m1 >>
rect 276 282 277 283 
<< m1 >>
rect 278 282 279 283 
<< pdiffusion >>
rect 282 282 283 283 
<< pdiffusion >>
rect 283 282 284 283 
<< pdiffusion >>
rect 284 282 285 283 
<< pdiffusion >>
rect 285 282 286 283 
<< m1 >>
rect 286 282 287 283 
<< pdiffusion >>
rect 286 282 287 283 
<< pdiffusion >>
rect 287 282 288 283 
<< pdiffusion >>
rect 300 282 301 283 
<< pdiffusion >>
rect 301 282 302 283 
<< pdiffusion >>
rect 302 282 303 283 
<< pdiffusion >>
rect 303 282 304 283 
<< pdiffusion >>
rect 304 282 305 283 
<< pdiffusion >>
rect 305 282 306 283 
<< m1 >>
rect 314 282 315 283 
<< m1 >>
rect 316 282 317 283 
<< pdiffusion >>
rect 318 282 319 283 
<< pdiffusion >>
rect 319 282 320 283 
<< pdiffusion >>
rect 320 282 321 283 
<< pdiffusion >>
rect 321 282 322 283 
<< pdiffusion >>
rect 322 282 323 283 
<< pdiffusion >>
rect 323 282 324 283 
<< m1 >>
rect 325 282 326 283 
<< m1 >>
rect 327 282 328 283 
<< m1 >>
rect 331 282 332 283 
<< pdiffusion >>
rect 336 282 337 283 
<< pdiffusion >>
rect 337 282 338 283 
<< pdiffusion >>
rect 338 282 339 283 
<< pdiffusion >>
rect 339 282 340 283 
<< pdiffusion >>
rect 340 282 341 283 
<< pdiffusion >>
rect 341 282 342 283 
<< m1 >>
rect 10 283 11 284 
<< pdiffusion >>
rect 12 283 13 284 
<< pdiffusion >>
rect 13 283 14 284 
<< pdiffusion >>
rect 14 283 15 284 
<< pdiffusion >>
rect 15 283 16 284 
<< pdiffusion >>
rect 16 283 17 284 
<< pdiffusion >>
rect 17 283 18 284 
<< m1 >>
rect 28 283 29 284 
<< m2 >>
rect 28 283 29 284 
<< pdiffusion >>
rect 30 283 31 284 
<< pdiffusion >>
rect 31 283 32 284 
<< pdiffusion >>
rect 32 283 33 284 
<< pdiffusion >>
rect 33 283 34 284 
<< pdiffusion >>
rect 34 283 35 284 
<< pdiffusion >>
rect 35 283 36 284 
<< m1 >>
rect 37 283 38 284 
<< m1 >>
rect 44 283 45 284 
<< pdiffusion >>
rect 48 283 49 284 
<< pdiffusion >>
rect 49 283 50 284 
<< pdiffusion >>
rect 50 283 51 284 
<< pdiffusion >>
rect 51 283 52 284 
<< pdiffusion >>
rect 52 283 53 284 
<< pdiffusion >>
rect 53 283 54 284 
<< m1 >>
rect 55 283 56 284 
<< m1 >>
rect 57 283 58 284 
<< m1 >>
rect 60 283 61 284 
<< m1 >>
rect 62 283 63 284 
<< m1 >>
rect 64 283 65 284 
<< pdiffusion >>
rect 66 283 67 284 
<< pdiffusion >>
rect 67 283 68 284 
<< pdiffusion >>
rect 68 283 69 284 
<< pdiffusion >>
rect 69 283 70 284 
<< pdiffusion >>
rect 70 283 71 284 
<< pdiffusion >>
rect 71 283 72 284 
<< m1 >>
rect 73 283 74 284 
<< pdiffusion >>
rect 84 283 85 284 
<< pdiffusion >>
rect 85 283 86 284 
<< pdiffusion >>
rect 86 283 87 284 
<< pdiffusion >>
rect 87 283 88 284 
<< pdiffusion >>
rect 88 283 89 284 
<< pdiffusion >>
rect 89 283 90 284 
<< pdiffusion >>
rect 102 283 103 284 
<< pdiffusion >>
rect 103 283 104 284 
<< pdiffusion >>
rect 104 283 105 284 
<< pdiffusion >>
rect 105 283 106 284 
<< pdiffusion >>
rect 106 283 107 284 
<< pdiffusion >>
rect 107 283 108 284 
<< m1 >>
rect 118 283 119 284 
<< pdiffusion >>
rect 120 283 121 284 
<< pdiffusion >>
rect 121 283 122 284 
<< pdiffusion >>
rect 122 283 123 284 
<< pdiffusion >>
rect 123 283 124 284 
<< pdiffusion >>
rect 124 283 125 284 
<< pdiffusion >>
rect 125 283 126 284 
<< m1 >>
rect 132 283 133 284 
<< m1 >>
rect 134 283 135 284 
<< m1 >>
rect 136 283 137 284 
<< pdiffusion >>
rect 138 283 139 284 
<< pdiffusion >>
rect 139 283 140 284 
<< pdiffusion >>
rect 140 283 141 284 
<< pdiffusion >>
rect 141 283 142 284 
<< pdiffusion >>
rect 142 283 143 284 
<< pdiffusion >>
rect 143 283 144 284 
<< pdiffusion >>
rect 156 283 157 284 
<< pdiffusion >>
rect 157 283 158 284 
<< pdiffusion >>
rect 158 283 159 284 
<< pdiffusion >>
rect 159 283 160 284 
<< pdiffusion >>
rect 160 283 161 284 
<< pdiffusion >>
rect 161 283 162 284 
<< m1 >>
rect 163 283 164 284 
<< m1 >>
rect 165 283 166 284 
<< m2 >>
rect 166 283 167 284 
<< m1 >>
rect 171 283 172 284 
<< m2 >>
rect 172 283 173 284 
<< pdiffusion >>
rect 174 283 175 284 
<< pdiffusion >>
rect 175 283 176 284 
<< pdiffusion >>
rect 176 283 177 284 
<< pdiffusion >>
rect 177 283 178 284 
<< pdiffusion >>
rect 178 283 179 284 
<< pdiffusion >>
rect 179 283 180 284 
<< m1 >>
rect 181 283 182 284 
<< m1 >>
rect 183 283 184 284 
<< m1 >>
rect 190 283 191 284 
<< pdiffusion >>
rect 192 283 193 284 
<< pdiffusion >>
rect 193 283 194 284 
<< pdiffusion >>
rect 194 283 195 284 
<< pdiffusion >>
rect 195 283 196 284 
<< pdiffusion >>
rect 196 283 197 284 
<< pdiffusion >>
rect 197 283 198 284 
<< m1 >>
rect 199 283 200 284 
<< m2 >>
rect 200 283 201 284 
<< pdiffusion >>
rect 210 283 211 284 
<< pdiffusion >>
rect 211 283 212 284 
<< pdiffusion >>
rect 212 283 213 284 
<< pdiffusion >>
rect 213 283 214 284 
<< pdiffusion >>
rect 214 283 215 284 
<< pdiffusion >>
rect 215 283 216 284 
<< m1 >>
rect 217 283 218 284 
<< m1 >>
rect 223 283 224 284 
<< m1 >>
rect 226 283 227 284 
<< pdiffusion >>
rect 228 283 229 284 
<< pdiffusion >>
rect 229 283 230 284 
<< pdiffusion >>
rect 230 283 231 284 
<< pdiffusion >>
rect 231 283 232 284 
<< pdiffusion >>
rect 232 283 233 284 
<< pdiffusion >>
rect 233 283 234 284 
<< m1 >>
rect 235 283 236 284 
<< m1 >>
rect 237 283 238 284 
<< m1 >>
rect 239 283 240 284 
<< m1 >>
rect 241 283 242 284 
<< pdiffusion >>
rect 246 283 247 284 
<< pdiffusion >>
rect 247 283 248 284 
<< pdiffusion >>
rect 248 283 249 284 
<< pdiffusion >>
rect 249 283 250 284 
<< pdiffusion >>
rect 250 283 251 284 
<< pdiffusion >>
rect 251 283 252 284 
<< pdiffusion >>
rect 264 283 265 284 
<< pdiffusion >>
rect 265 283 266 284 
<< pdiffusion >>
rect 266 283 267 284 
<< pdiffusion >>
rect 267 283 268 284 
<< pdiffusion >>
rect 268 283 269 284 
<< pdiffusion >>
rect 269 283 270 284 
<< m1 >>
rect 272 283 273 284 
<< m1 >>
rect 276 283 277 284 
<< m1 >>
rect 278 283 279 284 
<< pdiffusion >>
rect 282 283 283 284 
<< pdiffusion >>
rect 283 283 284 284 
<< pdiffusion >>
rect 284 283 285 284 
<< pdiffusion >>
rect 285 283 286 284 
<< pdiffusion >>
rect 286 283 287 284 
<< pdiffusion >>
rect 287 283 288 284 
<< pdiffusion >>
rect 300 283 301 284 
<< pdiffusion >>
rect 301 283 302 284 
<< pdiffusion >>
rect 302 283 303 284 
<< pdiffusion >>
rect 303 283 304 284 
<< pdiffusion >>
rect 304 283 305 284 
<< pdiffusion >>
rect 305 283 306 284 
<< m1 >>
rect 314 283 315 284 
<< m1 >>
rect 316 283 317 284 
<< pdiffusion >>
rect 318 283 319 284 
<< pdiffusion >>
rect 319 283 320 284 
<< pdiffusion >>
rect 320 283 321 284 
<< pdiffusion >>
rect 321 283 322 284 
<< pdiffusion >>
rect 322 283 323 284 
<< pdiffusion >>
rect 323 283 324 284 
<< m1 >>
rect 325 283 326 284 
<< m1 >>
rect 327 283 328 284 
<< m1 >>
rect 331 283 332 284 
<< pdiffusion >>
rect 336 283 337 284 
<< pdiffusion >>
rect 337 283 338 284 
<< pdiffusion >>
rect 338 283 339 284 
<< pdiffusion >>
rect 339 283 340 284 
<< pdiffusion >>
rect 340 283 341 284 
<< pdiffusion >>
rect 341 283 342 284 
<< m1 >>
rect 10 284 11 285 
<< pdiffusion >>
rect 12 284 13 285 
<< pdiffusion >>
rect 13 284 14 285 
<< pdiffusion >>
rect 14 284 15 285 
<< pdiffusion >>
rect 15 284 16 285 
<< pdiffusion >>
rect 16 284 17 285 
<< pdiffusion >>
rect 17 284 18 285 
<< m1 >>
rect 28 284 29 285 
<< m2 >>
rect 28 284 29 285 
<< pdiffusion >>
rect 30 284 31 285 
<< pdiffusion >>
rect 31 284 32 285 
<< pdiffusion >>
rect 32 284 33 285 
<< pdiffusion >>
rect 33 284 34 285 
<< pdiffusion >>
rect 34 284 35 285 
<< pdiffusion >>
rect 35 284 36 285 
<< m1 >>
rect 37 284 38 285 
<< m1 >>
rect 44 284 45 285 
<< pdiffusion >>
rect 48 284 49 285 
<< pdiffusion >>
rect 49 284 50 285 
<< pdiffusion >>
rect 50 284 51 285 
<< pdiffusion >>
rect 51 284 52 285 
<< pdiffusion >>
rect 52 284 53 285 
<< pdiffusion >>
rect 53 284 54 285 
<< m1 >>
rect 55 284 56 285 
<< m1 >>
rect 57 284 58 285 
<< m1 >>
rect 60 284 61 285 
<< m1 >>
rect 62 284 63 285 
<< m1 >>
rect 64 284 65 285 
<< pdiffusion >>
rect 66 284 67 285 
<< pdiffusion >>
rect 67 284 68 285 
<< pdiffusion >>
rect 68 284 69 285 
<< pdiffusion >>
rect 69 284 70 285 
<< pdiffusion >>
rect 70 284 71 285 
<< pdiffusion >>
rect 71 284 72 285 
<< m1 >>
rect 73 284 74 285 
<< pdiffusion >>
rect 84 284 85 285 
<< pdiffusion >>
rect 85 284 86 285 
<< pdiffusion >>
rect 86 284 87 285 
<< pdiffusion >>
rect 87 284 88 285 
<< pdiffusion >>
rect 88 284 89 285 
<< pdiffusion >>
rect 89 284 90 285 
<< pdiffusion >>
rect 102 284 103 285 
<< pdiffusion >>
rect 103 284 104 285 
<< pdiffusion >>
rect 104 284 105 285 
<< pdiffusion >>
rect 105 284 106 285 
<< pdiffusion >>
rect 106 284 107 285 
<< pdiffusion >>
rect 107 284 108 285 
<< m1 >>
rect 118 284 119 285 
<< pdiffusion >>
rect 120 284 121 285 
<< pdiffusion >>
rect 121 284 122 285 
<< pdiffusion >>
rect 122 284 123 285 
<< pdiffusion >>
rect 123 284 124 285 
<< pdiffusion >>
rect 124 284 125 285 
<< pdiffusion >>
rect 125 284 126 285 
<< m1 >>
rect 132 284 133 285 
<< m1 >>
rect 134 284 135 285 
<< m1 >>
rect 136 284 137 285 
<< pdiffusion >>
rect 138 284 139 285 
<< pdiffusion >>
rect 139 284 140 285 
<< pdiffusion >>
rect 140 284 141 285 
<< pdiffusion >>
rect 141 284 142 285 
<< pdiffusion >>
rect 142 284 143 285 
<< pdiffusion >>
rect 143 284 144 285 
<< pdiffusion >>
rect 156 284 157 285 
<< pdiffusion >>
rect 157 284 158 285 
<< pdiffusion >>
rect 158 284 159 285 
<< pdiffusion >>
rect 159 284 160 285 
<< pdiffusion >>
rect 160 284 161 285 
<< pdiffusion >>
rect 161 284 162 285 
<< m1 >>
rect 163 284 164 285 
<< m1 >>
rect 165 284 166 285 
<< m2 >>
rect 166 284 167 285 
<< m1 >>
rect 171 284 172 285 
<< m2 >>
rect 172 284 173 285 
<< pdiffusion >>
rect 174 284 175 285 
<< pdiffusion >>
rect 175 284 176 285 
<< pdiffusion >>
rect 176 284 177 285 
<< pdiffusion >>
rect 177 284 178 285 
<< pdiffusion >>
rect 178 284 179 285 
<< pdiffusion >>
rect 179 284 180 285 
<< m1 >>
rect 181 284 182 285 
<< m1 >>
rect 183 284 184 285 
<< m1 >>
rect 190 284 191 285 
<< pdiffusion >>
rect 192 284 193 285 
<< pdiffusion >>
rect 193 284 194 285 
<< pdiffusion >>
rect 194 284 195 285 
<< pdiffusion >>
rect 195 284 196 285 
<< pdiffusion >>
rect 196 284 197 285 
<< pdiffusion >>
rect 197 284 198 285 
<< m1 >>
rect 199 284 200 285 
<< m2 >>
rect 200 284 201 285 
<< pdiffusion >>
rect 210 284 211 285 
<< pdiffusion >>
rect 211 284 212 285 
<< pdiffusion >>
rect 212 284 213 285 
<< pdiffusion >>
rect 213 284 214 285 
<< pdiffusion >>
rect 214 284 215 285 
<< pdiffusion >>
rect 215 284 216 285 
<< m1 >>
rect 217 284 218 285 
<< m1 >>
rect 223 284 224 285 
<< m1 >>
rect 226 284 227 285 
<< pdiffusion >>
rect 228 284 229 285 
<< pdiffusion >>
rect 229 284 230 285 
<< pdiffusion >>
rect 230 284 231 285 
<< pdiffusion >>
rect 231 284 232 285 
<< pdiffusion >>
rect 232 284 233 285 
<< pdiffusion >>
rect 233 284 234 285 
<< m1 >>
rect 235 284 236 285 
<< m1 >>
rect 237 284 238 285 
<< m1 >>
rect 239 284 240 285 
<< m1 >>
rect 241 284 242 285 
<< pdiffusion >>
rect 246 284 247 285 
<< pdiffusion >>
rect 247 284 248 285 
<< pdiffusion >>
rect 248 284 249 285 
<< pdiffusion >>
rect 249 284 250 285 
<< pdiffusion >>
rect 250 284 251 285 
<< pdiffusion >>
rect 251 284 252 285 
<< pdiffusion >>
rect 264 284 265 285 
<< pdiffusion >>
rect 265 284 266 285 
<< pdiffusion >>
rect 266 284 267 285 
<< pdiffusion >>
rect 267 284 268 285 
<< pdiffusion >>
rect 268 284 269 285 
<< pdiffusion >>
rect 269 284 270 285 
<< m1 >>
rect 272 284 273 285 
<< m1 >>
rect 276 284 277 285 
<< m1 >>
rect 278 284 279 285 
<< pdiffusion >>
rect 282 284 283 285 
<< pdiffusion >>
rect 283 284 284 285 
<< pdiffusion >>
rect 284 284 285 285 
<< pdiffusion >>
rect 285 284 286 285 
<< pdiffusion >>
rect 286 284 287 285 
<< pdiffusion >>
rect 287 284 288 285 
<< pdiffusion >>
rect 300 284 301 285 
<< pdiffusion >>
rect 301 284 302 285 
<< pdiffusion >>
rect 302 284 303 285 
<< pdiffusion >>
rect 303 284 304 285 
<< pdiffusion >>
rect 304 284 305 285 
<< pdiffusion >>
rect 305 284 306 285 
<< m1 >>
rect 314 284 315 285 
<< m1 >>
rect 316 284 317 285 
<< pdiffusion >>
rect 318 284 319 285 
<< pdiffusion >>
rect 319 284 320 285 
<< pdiffusion >>
rect 320 284 321 285 
<< pdiffusion >>
rect 321 284 322 285 
<< pdiffusion >>
rect 322 284 323 285 
<< pdiffusion >>
rect 323 284 324 285 
<< m1 >>
rect 325 284 326 285 
<< m1 >>
rect 327 284 328 285 
<< m1 >>
rect 331 284 332 285 
<< pdiffusion >>
rect 336 284 337 285 
<< pdiffusion >>
rect 337 284 338 285 
<< pdiffusion >>
rect 338 284 339 285 
<< pdiffusion >>
rect 339 284 340 285 
<< pdiffusion >>
rect 340 284 341 285 
<< pdiffusion >>
rect 341 284 342 285 
<< m1 >>
rect 10 285 11 286 
<< pdiffusion >>
rect 12 285 13 286 
<< pdiffusion >>
rect 13 285 14 286 
<< pdiffusion >>
rect 14 285 15 286 
<< pdiffusion >>
rect 15 285 16 286 
<< pdiffusion >>
rect 16 285 17 286 
<< pdiffusion >>
rect 17 285 18 286 
<< m1 >>
rect 28 285 29 286 
<< m2 >>
rect 28 285 29 286 
<< pdiffusion >>
rect 30 285 31 286 
<< pdiffusion >>
rect 31 285 32 286 
<< pdiffusion >>
rect 32 285 33 286 
<< pdiffusion >>
rect 33 285 34 286 
<< pdiffusion >>
rect 34 285 35 286 
<< pdiffusion >>
rect 35 285 36 286 
<< m1 >>
rect 37 285 38 286 
<< m1 >>
rect 44 285 45 286 
<< pdiffusion >>
rect 48 285 49 286 
<< pdiffusion >>
rect 49 285 50 286 
<< pdiffusion >>
rect 50 285 51 286 
<< pdiffusion >>
rect 51 285 52 286 
<< pdiffusion >>
rect 52 285 53 286 
<< pdiffusion >>
rect 53 285 54 286 
<< m1 >>
rect 55 285 56 286 
<< m1 >>
rect 57 285 58 286 
<< m1 >>
rect 60 285 61 286 
<< m1 >>
rect 62 285 63 286 
<< m1 >>
rect 64 285 65 286 
<< pdiffusion >>
rect 66 285 67 286 
<< pdiffusion >>
rect 67 285 68 286 
<< pdiffusion >>
rect 68 285 69 286 
<< pdiffusion >>
rect 69 285 70 286 
<< pdiffusion >>
rect 70 285 71 286 
<< pdiffusion >>
rect 71 285 72 286 
<< m1 >>
rect 73 285 74 286 
<< pdiffusion >>
rect 84 285 85 286 
<< pdiffusion >>
rect 85 285 86 286 
<< pdiffusion >>
rect 86 285 87 286 
<< pdiffusion >>
rect 87 285 88 286 
<< pdiffusion >>
rect 88 285 89 286 
<< pdiffusion >>
rect 89 285 90 286 
<< pdiffusion >>
rect 102 285 103 286 
<< pdiffusion >>
rect 103 285 104 286 
<< pdiffusion >>
rect 104 285 105 286 
<< pdiffusion >>
rect 105 285 106 286 
<< pdiffusion >>
rect 106 285 107 286 
<< pdiffusion >>
rect 107 285 108 286 
<< m1 >>
rect 118 285 119 286 
<< pdiffusion >>
rect 120 285 121 286 
<< pdiffusion >>
rect 121 285 122 286 
<< pdiffusion >>
rect 122 285 123 286 
<< pdiffusion >>
rect 123 285 124 286 
<< pdiffusion >>
rect 124 285 125 286 
<< pdiffusion >>
rect 125 285 126 286 
<< m1 >>
rect 132 285 133 286 
<< m1 >>
rect 134 285 135 286 
<< m1 >>
rect 136 285 137 286 
<< pdiffusion >>
rect 138 285 139 286 
<< pdiffusion >>
rect 139 285 140 286 
<< pdiffusion >>
rect 140 285 141 286 
<< pdiffusion >>
rect 141 285 142 286 
<< pdiffusion >>
rect 142 285 143 286 
<< pdiffusion >>
rect 143 285 144 286 
<< pdiffusion >>
rect 156 285 157 286 
<< pdiffusion >>
rect 157 285 158 286 
<< pdiffusion >>
rect 158 285 159 286 
<< pdiffusion >>
rect 159 285 160 286 
<< pdiffusion >>
rect 160 285 161 286 
<< pdiffusion >>
rect 161 285 162 286 
<< m1 >>
rect 163 285 164 286 
<< m1 >>
rect 165 285 166 286 
<< m2 >>
rect 166 285 167 286 
<< m1 >>
rect 171 285 172 286 
<< m2 >>
rect 172 285 173 286 
<< pdiffusion >>
rect 174 285 175 286 
<< pdiffusion >>
rect 175 285 176 286 
<< pdiffusion >>
rect 176 285 177 286 
<< pdiffusion >>
rect 177 285 178 286 
<< pdiffusion >>
rect 178 285 179 286 
<< pdiffusion >>
rect 179 285 180 286 
<< m1 >>
rect 181 285 182 286 
<< m1 >>
rect 183 285 184 286 
<< m1 >>
rect 190 285 191 286 
<< pdiffusion >>
rect 192 285 193 286 
<< pdiffusion >>
rect 193 285 194 286 
<< pdiffusion >>
rect 194 285 195 286 
<< pdiffusion >>
rect 195 285 196 286 
<< pdiffusion >>
rect 196 285 197 286 
<< pdiffusion >>
rect 197 285 198 286 
<< m1 >>
rect 199 285 200 286 
<< m2 >>
rect 200 285 201 286 
<< pdiffusion >>
rect 210 285 211 286 
<< pdiffusion >>
rect 211 285 212 286 
<< pdiffusion >>
rect 212 285 213 286 
<< pdiffusion >>
rect 213 285 214 286 
<< pdiffusion >>
rect 214 285 215 286 
<< pdiffusion >>
rect 215 285 216 286 
<< m1 >>
rect 217 285 218 286 
<< m1 >>
rect 223 285 224 286 
<< m1 >>
rect 226 285 227 286 
<< pdiffusion >>
rect 228 285 229 286 
<< pdiffusion >>
rect 229 285 230 286 
<< pdiffusion >>
rect 230 285 231 286 
<< pdiffusion >>
rect 231 285 232 286 
<< pdiffusion >>
rect 232 285 233 286 
<< pdiffusion >>
rect 233 285 234 286 
<< m1 >>
rect 235 285 236 286 
<< m1 >>
rect 237 285 238 286 
<< m1 >>
rect 239 285 240 286 
<< m1 >>
rect 241 285 242 286 
<< pdiffusion >>
rect 246 285 247 286 
<< pdiffusion >>
rect 247 285 248 286 
<< pdiffusion >>
rect 248 285 249 286 
<< pdiffusion >>
rect 249 285 250 286 
<< pdiffusion >>
rect 250 285 251 286 
<< pdiffusion >>
rect 251 285 252 286 
<< pdiffusion >>
rect 264 285 265 286 
<< pdiffusion >>
rect 265 285 266 286 
<< pdiffusion >>
rect 266 285 267 286 
<< pdiffusion >>
rect 267 285 268 286 
<< pdiffusion >>
rect 268 285 269 286 
<< pdiffusion >>
rect 269 285 270 286 
<< m1 >>
rect 272 285 273 286 
<< m1 >>
rect 276 285 277 286 
<< m1 >>
rect 278 285 279 286 
<< pdiffusion >>
rect 282 285 283 286 
<< pdiffusion >>
rect 283 285 284 286 
<< pdiffusion >>
rect 284 285 285 286 
<< pdiffusion >>
rect 285 285 286 286 
<< pdiffusion >>
rect 286 285 287 286 
<< pdiffusion >>
rect 287 285 288 286 
<< pdiffusion >>
rect 300 285 301 286 
<< pdiffusion >>
rect 301 285 302 286 
<< pdiffusion >>
rect 302 285 303 286 
<< pdiffusion >>
rect 303 285 304 286 
<< pdiffusion >>
rect 304 285 305 286 
<< pdiffusion >>
rect 305 285 306 286 
<< m1 >>
rect 314 285 315 286 
<< m1 >>
rect 316 285 317 286 
<< pdiffusion >>
rect 318 285 319 286 
<< pdiffusion >>
rect 319 285 320 286 
<< pdiffusion >>
rect 320 285 321 286 
<< pdiffusion >>
rect 321 285 322 286 
<< pdiffusion >>
rect 322 285 323 286 
<< pdiffusion >>
rect 323 285 324 286 
<< m1 >>
rect 325 285 326 286 
<< m1 >>
rect 327 285 328 286 
<< m1 >>
rect 331 285 332 286 
<< pdiffusion >>
rect 336 285 337 286 
<< pdiffusion >>
rect 337 285 338 286 
<< pdiffusion >>
rect 338 285 339 286 
<< pdiffusion >>
rect 339 285 340 286 
<< pdiffusion >>
rect 340 285 341 286 
<< pdiffusion >>
rect 341 285 342 286 
<< m1 >>
rect 10 286 11 287 
<< pdiffusion >>
rect 12 286 13 287 
<< pdiffusion >>
rect 13 286 14 287 
<< pdiffusion >>
rect 14 286 15 287 
<< pdiffusion >>
rect 15 286 16 287 
<< pdiffusion >>
rect 16 286 17 287 
<< pdiffusion >>
rect 17 286 18 287 
<< m1 >>
rect 28 286 29 287 
<< m2 >>
rect 28 286 29 287 
<< pdiffusion >>
rect 30 286 31 287 
<< pdiffusion >>
rect 31 286 32 287 
<< pdiffusion >>
rect 32 286 33 287 
<< pdiffusion >>
rect 33 286 34 287 
<< pdiffusion >>
rect 34 286 35 287 
<< pdiffusion >>
rect 35 286 36 287 
<< m1 >>
rect 37 286 38 287 
<< m1 >>
rect 44 286 45 287 
<< pdiffusion >>
rect 48 286 49 287 
<< pdiffusion >>
rect 49 286 50 287 
<< pdiffusion >>
rect 50 286 51 287 
<< pdiffusion >>
rect 51 286 52 287 
<< pdiffusion >>
rect 52 286 53 287 
<< pdiffusion >>
rect 53 286 54 287 
<< m1 >>
rect 55 286 56 287 
<< m1 >>
rect 57 286 58 287 
<< m1 >>
rect 60 286 61 287 
<< m1 >>
rect 62 286 63 287 
<< m1 >>
rect 64 286 65 287 
<< pdiffusion >>
rect 66 286 67 287 
<< pdiffusion >>
rect 67 286 68 287 
<< pdiffusion >>
rect 68 286 69 287 
<< pdiffusion >>
rect 69 286 70 287 
<< pdiffusion >>
rect 70 286 71 287 
<< pdiffusion >>
rect 71 286 72 287 
<< m1 >>
rect 73 286 74 287 
<< pdiffusion >>
rect 84 286 85 287 
<< pdiffusion >>
rect 85 286 86 287 
<< pdiffusion >>
rect 86 286 87 287 
<< pdiffusion >>
rect 87 286 88 287 
<< pdiffusion >>
rect 88 286 89 287 
<< pdiffusion >>
rect 89 286 90 287 
<< pdiffusion >>
rect 102 286 103 287 
<< pdiffusion >>
rect 103 286 104 287 
<< pdiffusion >>
rect 104 286 105 287 
<< pdiffusion >>
rect 105 286 106 287 
<< pdiffusion >>
rect 106 286 107 287 
<< pdiffusion >>
rect 107 286 108 287 
<< m1 >>
rect 118 286 119 287 
<< pdiffusion >>
rect 120 286 121 287 
<< pdiffusion >>
rect 121 286 122 287 
<< pdiffusion >>
rect 122 286 123 287 
<< pdiffusion >>
rect 123 286 124 287 
<< pdiffusion >>
rect 124 286 125 287 
<< pdiffusion >>
rect 125 286 126 287 
<< m1 >>
rect 132 286 133 287 
<< m1 >>
rect 134 286 135 287 
<< m1 >>
rect 136 286 137 287 
<< pdiffusion >>
rect 138 286 139 287 
<< pdiffusion >>
rect 139 286 140 287 
<< pdiffusion >>
rect 140 286 141 287 
<< pdiffusion >>
rect 141 286 142 287 
<< pdiffusion >>
rect 142 286 143 287 
<< pdiffusion >>
rect 143 286 144 287 
<< pdiffusion >>
rect 156 286 157 287 
<< pdiffusion >>
rect 157 286 158 287 
<< pdiffusion >>
rect 158 286 159 287 
<< pdiffusion >>
rect 159 286 160 287 
<< pdiffusion >>
rect 160 286 161 287 
<< pdiffusion >>
rect 161 286 162 287 
<< m1 >>
rect 163 286 164 287 
<< m1 >>
rect 165 286 166 287 
<< m2 >>
rect 166 286 167 287 
<< m1 >>
rect 171 286 172 287 
<< m2 >>
rect 172 286 173 287 
<< pdiffusion >>
rect 174 286 175 287 
<< pdiffusion >>
rect 175 286 176 287 
<< pdiffusion >>
rect 176 286 177 287 
<< pdiffusion >>
rect 177 286 178 287 
<< pdiffusion >>
rect 178 286 179 287 
<< pdiffusion >>
rect 179 286 180 287 
<< m1 >>
rect 181 286 182 287 
<< m1 >>
rect 183 286 184 287 
<< m1 >>
rect 190 286 191 287 
<< pdiffusion >>
rect 192 286 193 287 
<< pdiffusion >>
rect 193 286 194 287 
<< pdiffusion >>
rect 194 286 195 287 
<< pdiffusion >>
rect 195 286 196 287 
<< pdiffusion >>
rect 196 286 197 287 
<< pdiffusion >>
rect 197 286 198 287 
<< m1 >>
rect 199 286 200 287 
<< m2 >>
rect 200 286 201 287 
<< pdiffusion >>
rect 210 286 211 287 
<< pdiffusion >>
rect 211 286 212 287 
<< pdiffusion >>
rect 212 286 213 287 
<< pdiffusion >>
rect 213 286 214 287 
<< pdiffusion >>
rect 214 286 215 287 
<< pdiffusion >>
rect 215 286 216 287 
<< m1 >>
rect 217 286 218 287 
<< m1 >>
rect 223 286 224 287 
<< m1 >>
rect 226 286 227 287 
<< pdiffusion >>
rect 228 286 229 287 
<< pdiffusion >>
rect 229 286 230 287 
<< pdiffusion >>
rect 230 286 231 287 
<< pdiffusion >>
rect 231 286 232 287 
<< pdiffusion >>
rect 232 286 233 287 
<< pdiffusion >>
rect 233 286 234 287 
<< m1 >>
rect 235 286 236 287 
<< m1 >>
rect 237 286 238 287 
<< m1 >>
rect 239 286 240 287 
<< m1 >>
rect 241 286 242 287 
<< pdiffusion >>
rect 246 286 247 287 
<< pdiffusion >>
rect 247 286 248 287 
<< pdiffusion >>
rect 248 286 249 287 
<< pdiffusion >>
rect 249 286 250 287 
<< pdiffusion >>
rect 250 286 251 287 
<< pdiffusion >>
rect 251 286 252 287 
<< pdiffusion >>
rect 264 286 265 287 
<< pdiffusion >>
rect 265 286 266 287 
<< pdiffusion >>
rect 266 286 267 287 
<< pdiffusion >>
rect 267 286 268 287 
<< pdiffusion >>
rect 268 286 269 287 
<< pdiffusion >>
rect 269 286 270 287 
<< m1 >>
rect 272 286 273 287 
<< m1 >>
rect 276 286 277 287 
<< m1 >>
rect 278 286 279 287 
<< pdiffusion >>
rect 282 286 283 287 
<< pdiffusion >>
rect 283 286 284 287 
<< pdiffusion >>
rect 284 286 285 287 
<< pdiffusion >>
rect 285 286 286 287 
<< pdiffusion >>
rect 286 286 287 287 
<< pdiffusion >>
rect 287 286 288 287 
<< pdiffusion >>
rect 300 286 301 287 
<< pdiffusion >>
rect 301 286 302 287 
<< pdiffusion >>
rect 302 286 303 287 
<< pdiffusion >>
rect 303 286 304 287 
<< pdiffusion >>
rect 304 286 305 287 
<< pdiffusion >>
rect 305 286 306 287 
<< m1 >>
rect 314 286 315 287 
<< m1 >>
rect 316 286 317 287 
<< pdiffusion >>
rect 318 286 319 287 
<< pdiffusion >>
rect 319 286 320 287 
<< pdiffusion >>
rect 320 286 321 287 
<< pdiffusion >>
rect 321 286 322 287 
<< pdiffusion >>
rect 322 286 323 287 
<< pdiffusion >>
rect 323 286 324 287 
<< m1 >>
rect 325 286 326 287 
<< m1 >>
rect 327 286 328 287 
<< m1 >>
rect 331 286 332 287 
<< pdiffusion >>
rect 336 286 337 287 
<< pdiffusion >>
rect 337 286 338 287 
<< pdiffusion >>
rect 338 286 339 287 
<< pdiffusion >>
rect 339 286 340 287 
<< pdiffusion >>
rect 340 286 341 287 
<< pdiffusion >>
rect 341 286 342 287 
<< m1 >>
rect 10 287 11 288 
<< pdiffusion >>
rect 12 287 13 288 
<< pdiffusion >>
rect 13 287 14 288 
<< pdiffusion >>
rect 14 287 15 288 
<< pdiffusion >>
rect 15 287 16 288 
<< pdiffusion >>
rect 16 287 17 288 
<< pdiffusion >>
rect 17 287 18 288 
<< m1 >>
rect 28 287 29 288 
<< m2 >>
rect 28 287 29 288 
<< pdiffusion >>
rect 30 287 31 288 
<< pdiffusion >>
rect 31 287 32 288 
<< pdiffusion >>
rect 32 287 33 288 
<< pdiffusion >>
rect 33 287 34 288 
<< pdiffusion >>
rect 34 287 35 288 
<< pdiffusion >>
rect 35 287 36 288 
<< m1 >>
rect 37 287 38 288 
<< m1 >>
rect 44 287 45 288 
<< pdiffusion >>
rect 48 287 49 288 
<< pdiffusion >>
rect 49 287 50 288 
<< pdiffusion >>
rect 50 287 51 288 
<< pdiffusion >>
rect 51 287 52 288 
<< pdiffusion >>
rect 52 287 53 288 
<< pdiffusion >>
rect 53 287 54 288 
<< m1 >>
rect 55 287 56 288 
<< m1 >>
rect 57 287 58 288 
<< m1 >>
rect 60 287 61 288 
<< m1 >>
rect 62 287 63 288 
<< m1 >>
rect 64 287 65 288 
<< pdiffusion >>
rect 66 287 67 288 
<< m1 >>
rect 67 287 68 288 
<< pdiffusion >>
rect 67 287 68 288 
<< pdiffusion >>
rect 68 287 69 288 
<< pdiffusion >>
rect 69 287 70 288 
<< pdiffusion >>
rect 70 287 71 288 
<< pdiffusion >>
rect 71 287 72 288 
<< m1 >>
rect 73 287 74 288 
<< pdiffusion >>
rect 84 287 85 288 
<< pdiffusion >>
rect 85 287 86 288 
<< pdiffusion >>
rect 86 287 87 288 
<< pdiffusion >>
rect 87 287 88 288 
<< pdiffusion >>
rect 88 287 89 288 
<< pdiffusion >>
rect 89 287 90 288 
<< pdiffusion >>
rect 102 287 103 288 
<< pdiffusion >>
rect 103 287 104 288 
<< pdiffusion >>
rect 104 287 105 288 
<< pdiffusion >>
rect 105 287 106 288 
<< pdiffusion >>
rect 106 287 107 288 
<< pdiffusion >>
rect 107 287 108 288 
<< m1 >>
rect 118 287 119 288 
<< pdiffusion >>
rect 120 287 121 288 
<< m1 >>
rect 121 287 122 288 
<< pdiffusion >>
rect 121 287 122 288 
<< pdiffusion >>
rect 122 287 123 288 
<< pdiffusion >>
rect 123 287 124 288 
<< pdiffusion >>
rect 124 287 125 288 
<< pdiffusion >>
rect 125 287 126 288 
<< m1 >>
rect 132 287 133 288 
<< m1 >>
rect 134 287 135 288 
<< m1 >>
rect 136 287 137 288 
<< pdiffusion >>
rect 138 287 139 288 
<< pdiffusion >>
rect 139 287 140 288 
<< pdiffusion >>
rect 140 287 141 288 
<< pdiffusion >>
rect 141 287 142 288 
<< pdiffusion >>
rect 142 287 143 288 
<< pdiffusion >>
rect 143 287 144 288 
<< pdiffusion >>
rect 156 287 157 288 
<< pdiffusion >>
rect 157 287 158 288 
<< pdiffusion >>
rect 158 287 159 288 
<< pdiffusion >>
rect 159 287 160 288 
<< pdiffusion >>
rect 160 287 161 288 
<< pdiffusion >>
rect 161 287 162 288 
<< m1 >>
rect 163 287 164 288 
<< m1 >>
rect 165 287 166 288 
<< m2 >>
rect 166 287 167 288 
<< m1 >>
rect 171 287 172 288 
<< m2 >>
rect 172 287 173 288 
<< pdiffusion >>
rect 174 287 175 288 
<< m1 >>
rect 175 287 176 288 
<< pdiffusion >>
rect 175 287 176 288 
<< pdiffusion >>
rect 176 287 177 288 
<< pdiffusion >>
rect 177 287 178 288 
<< m1 >>
rect 178 287 179 288 
<< pdiffusion >>
rect 178 287 179 288 
<< pdiffusion >>
rect 179 287 180 288 
<< m1 >>
rect 181 287 182 288 
<< m1 >>
rect 183 287 184 288 
<< m1 >>
rect 190 287 191 288 
<< pdiffusion >>
rect 192 287 193 288 
<< pdiffusion >>
rect 193 287 194 288 
<< pdiffusion >>
rect 194 287 195 288 
<< pdiffusion >>
rect 195 287 196 288 
<< pdiffusion >>
rect 196 287 197 288 
<< pdiffusion >>
rect 197 287 198 288 
<< m1 >>
rect 199 287 200 288 
<< m2 >>
rect 200 287 201 288 
<< pdiffusion >>
rect 210 287 211 288 
<< pdiffusion >>
rect 211 287 212 288 
<< pdiffusion >>
rect 212 287 213 288 
<< pdiffusion >>
rect 213 287 214 288 
<< m1 >>
rect 214 287 215 288 
<< pdiffusion >>
rect 214 287 215 288 
<< pdiffusion >>
rect 215 287 216 288 
<< m1 >>
rect 217 287 218 288 
<< m1 >>
rect 223 287 224 288 
<< m1 >>
rect 226 287 227 288 
<< pdiffusion >>
rect 228 287 229 288 
<< pdiffusion >>
rect 229 287 230 288 
<< pdiffusion >>
rect 230 287 231 288 
<< pdiffusion >>
rect 231 287 232 288 
<< m1 >>
rect 232 287 233 288 
<< pdiffusion >>
rect 232 287 233 288 
<< pdiffusion >>
rect 233 287 234 288 
<< m1 >>
rect 235 287 236 288 
<< m1 >>
rect 237 287 238 288 
<< m1 >>
rect 239 287 240 288 
<< m1 >>
rect 241 287 242 288 
<< pdiffusion >>
rect 246 287 247 288 
<< pdiffusion >>
rect 247 287 248 288 
<< pdiffusion >>
rect 248 287 249 288 
<< pdiffusion >>
rect 249 287 250 288 
<< pdiffusion >>
rect 250 287 251 288 
<< pdiffusion >>
rect 251 287 252 288 
<< pdiffusion >>
rect 264 287 265 288 
<< pdiffusion >>
rect 265 287 266 288 
<< pdiffusion >>
rect 266 287 267 288 
<< pdiffusion >>
rect 267 287 268 288 
<< pdiffusion >>
rect 268 287 269 288 
<< pdiffusion >>
rect 269 287 270 288 
<< m1 >>
rect 272 287 273 288 
<< m1 >>
rect 276 287 277 288 
<< m1 >>
rect 278 287 279 288 
<< pdiffusion >>
rect 282 287 283 288 
<< pdiffusion >>
rect 283 287 284 288 
<< pdiffusion >>
rect 284 287 285 288 
<< pdiffusion >>
rect 285 287 286 288 
<< pdiffusion >>
rect 286 287 287 288 
<< pdiffusion >>
rect 287 287 288 288 
<< pdiffusion >>
rect 300 287 301 288 
<< pdiffusion >>
rect 301 287 302 288 
<< pdiffusion >>
rect 302 287 303 288 
<< pdiffusion >>
rect 303 287 304 288 
<< m1 >>
rect 304 287 305 288 
<< pdiffusion >>
rect 304 287 305 288 
<< pdiffusion >>
rect 305 287 306 288 
<< m1 >>
rect 314 287 315 288 
<< m2 >>
rect 314 287 315 288 
<< m2c >>
rect 314 287 315 288 
<< m1 >>
rect 314 287 315 288 
<< m2 >>
rect 314 287 315 288 
<< m2 >>
rect 315 287 316 288 
<< m1 >>
rect 316 287 317 288 
<< m2 >>
rect 316 287 317 288 
<< pdiffusion >>
rect 318 287 319 288 
<< pdiffusion >>
rect 319 287 320 288 
<< pdiffusion >>
rect 320 287 321 288 
<< pdiffusion >>
rect 321 287 322 288 
<< pdiffusion >>
rect 322 287 323 288 
<< pdiffusion >>
rect 323 287 324 288 
<< m1 >>
rect 325 287 326 288 
<< m1 >>
rect 327 287 328 288 
<< m1 >>
rect 331 287 332 288 
<< pdiffusion >>
rect 336 287 337 288 
<< pdiffusion >>
rect 337 287 338 288 
<< pdiffusion >>
rect 338 287 339 288 
<< pdiffusion >>
rect 339 287 340 288 
<< m1 >>
rect 340 287 341 288 
<< pdiffusion >>
rect 340 287 341 288 
<< pdiffusion >>
rect 341 287 342 288 
<< m1 >>
rect 10 288 11 289 
<< m1 >>
rect 28 288 29 289 
<< m2 >>
rect 28 288 29 289 
<< m1 >>
rect 37 288 38 289 
<< m1 >>
rect 44 288 45 289 
<< m1 >>
rect 55 288 56 289 
<< m1 >>
rect 57 288 58 289 
<< m1 >>
rect 60 288 61 289 
<< m1 >>
rect 62 288 63 289 
<< m1 >>
rect 64 288 65 289 
<< m1 >>
rect 67 288 68 289 
<< m1 >>
rect 73 288 74 289 
<< m1 >>
rect 118 288 119 289 
<< m1 >>
rect 121 288 122 289 
<< m1 >>
rect 132 288 133 289 
<< m1 >>
rect 134 288 135 289 
<< m1 >>
rect 136 288 137 289 
<< m1 >>
rect 163 288 164 289 
<< m1 >>
rect 165 288 166 289 
<< m2 >>
rect 166 288 167 289 
<< m1 >>
rect 171 288 172 289 
<< m2 >>
rect 172 288 173 289 
<< m1 >>
rect 175 288 176 289 
<< m1 >>
rect 178 288 179 289 
<< m1 >>
rect 181 288 182 289 
<< m1 >>
rect 183 288 184 289 
<< m1 >>
rect 190 288 191 289 
<< m1 >>
rect 199 288 200 289 
<< m2 >>
rect 200 288 201 289 
<< m1 >>
rect 214 288 215 289 
<< m1 >>
rect 217 288 218 289 
<< m1 >>
rect 223 288 224 289 
<< m1 >>
rect 226 288 227 289 
<< m1 >>
rect 232 288 233 289 
<< m1 >>
rect 235 288 236 289 
<< m1 >>
rect 237 288 238 289 
<< m1 >>
rect 239 288 240 289 
<< m1 >>
rect 241 288 242 289 
<< m1 >>
rect 272 288 273 289 
<< m1 >>
rect 276 288 277 289 
<< m1 >>
rect 278 288 279 289 
<< m1 >>
rect 304 288 305 289 
<< m1 >>
rect 316 288 317 289 
<< m2 >>
rect 316 288 317 289 
<< m1 >>
rect 325 288 326 289 
<< m1 >>
rect 327 288 328 289 
<< m1 >>
rect 331 288 332 289 
<< m1 >>
rect 340 288 341 289 
<< m1 >>
rect 10 289 11 290 
<< m1 >>
rect 28 289 29 290 
<< m2 >>
rect 28 289 29 290 
<< m1 >>
rect 37 289 38 290 
<< m1 >>
rect 44 289 45 290 
<< m1 >>
rect 55 289 56 290 
<< m1 >>
rect 57 289 58 290 
<< m1 >>
rect 60 289 61 290 
<< m1 >>
rect 62 289 63 290 
<< m1 >>
rect 64 289 65 290 
<< m1 >>
rect 67 289 68 290 
<< m1 >>
rect 73 289 74 290 
<< m1 >>
rect 118 289 119 290 
<< m1 >>
rect 119 289 120 290 
<< m1 >>
rect 120 289 121 290 
<< m1 >>
rect 121 289 122 290 
<< m1 >>
rect 132 289 133 290 
<< m1 >>
rect 134 289 135 290 
<< m1 >>
rect 136 289 137 290 
<< m1 >>
rect 163 289 164 290 
<< m1 >>
rect 165 289 166 290 
<< m2 >>
rect 166 289 167 290 
<< m1 >>
rect 171 289 172 290 
<< m2 >>
rect 172 289 173 290 
<< m1 >>
rect 173 289 174 290 
<< m2 >>
rect 173 289 174 290 
<< m2c >>
rect 173 289 174 290 
<< m1 >>
rect 173 289 174 290 
<< m2 >>
rect 173 289 174 290 
<< m1 >>
rect 174 289 175 290 
<< m1 >>
rect 175 289 176 290 
<< m1 >>
rect 178 289 179 290 
<< m1 >>
rect 179 289 180 290 
<< m2 >>
rect 179 289 180 290 
<< m2c >>
rect 179 289 180 290 
<< m1 >>
rect 179 289 180 290 
<< m2 >>
rect 179 289 180 290 
<< m2 >>
rect 180 289 181 290 
<< m1 >>
rect 181 289 182 290 
<< m2 >>
rect 181 289 182 290 
<< m2 >>
rect 182 289 183 290 
<< m1 >>
rect 183 289 184 290 
<< m2 >>
rect 183 289 184 290 
<< m2c >>
rect 183 289 184 290 
<< m1 >>
rect 183 289 184 290 
<< m2 >>
rect 183 289 184 290 
<< m1 >>
rect 190 289 191 290 
<< m1 >>
rect 199 289 200 290 
<< m2 >>
rect 200 289 201 290 
<< m1 >>
rect 214 289 215 290 
<< m1 >>
rect 217 289 218 290 
<< m1 >>
rect 223 289 224 290 
<< m1 >>
rect 226 289 227 290 
<< m1 >>
rect 232 289 233 290 
<< m1 >>
rect 233 289 234 290 
<< m1 >>
rect 234 289 235 290 
<< m1 >>
rect 235 289 236 290 
<< m1 >>
rect 237 289 238 290 
<< m1 >>
rect 239 289 240 290 
<< m1 >>
rect 241 289 242 290 
<< m1 >>
rect 272 289 273 290 
<< m1 >>
rect 276 289 277 290 
<< m1 >>
rect 278 289 279 290 
<< m1 >>
rect 304 289 305 290 
<< m1 >>
rect 305 289 306 290 
<< m1 >>
rect 306 289 307 290 
<< m1 >>
rect 307 289 308 290 
<< m1 >>
rect 308 289 309 290 
<< m1 >>
rect 309 289 310 290 
<< m1 >>
rect 310 289 311 290 
<< m1 >>
rect 311 289 312 290 
<< m1 >>
rect 312 289 313 290 
<< m1 >>
rect 313 289 314 290 
<< m1 >>
rect 314 289 315 290 
<< m1 >>
rect 315 289 316 290 
<< m1 >>
rect 316 289 317 290 
<< m2 >>
rect 316 289 317 290 
<< m1 >>
rect 325 289 326 290 
<< m1 >>
rect 327 289 328 290 
<< m1 >>
rect 331 289 332 290 
<< m1 >>
rect 340 289 341 290 
<< m1 >>
rect 10 290 11 291 
<< m1 >>
rect 28 290 29 291 
<< m2 >>
rect 28 290 29 291 
<< m1 >>
rect 29 290 30 291 
<< m1 >>
rect 30 290 31 291 
<< m2 >>
rect 30 290 31 291 
<< m2c >>
rect 30 290 31 291 
<< m1 >>
rect 30 290 31 291 
<< m2 >>
rect 30 290 31 291 
<< m1 >>
rect 37 290 38 291 
<< m2 >>
rect 37 290 38 291 
<< m2c >>
rect 37 290 38 291 
<< m1 >>
rect 37 290 38 291 
<< m2 >>
rect 37 290 38 291 
<< m1 >>
rect 44 290 45 291 
<< m1 >>
rect 45 290 46 291 
<< m1 >>
rect 46 290 47 291 
<< m2 >>
rect 46 290 47 291 
<< m2c >>
rect 46 290 47 291 
<< m1 >>
rect 46 290 47 291 
<< m2 >>
rect 46 290 47 291 
<< m1 >>
rect 55 290 56 291 
<< m2 >>
rect 55 290 56 291 
<< m2c >>
rect 55 290 56 291 
<< m1 >>
rect 55 290 56 291 
<< m2 >>
rect 55 290 56 291 
<< m1 >>
rect 57 290 58 291 
<< m2 >>
rect 57 290 58 291 
<< m2c >>
rect 57 290 58 291 
<< m1 >>
rect 57 290 58 291 
<< m2 >>
rect 57 290 58 291 
<< m1 >>
rect 60 290 61 291 
<< m2 >>
rect 60 290 61 291 
<< m2c >>
rect 60 290 61 291 
<< m1 >>
rect 60 290 61 291 
<< m2 >>
rect 60 290 61 291 
<< m1 >>
rect 62 290 63 291 
<< m2 >>
rect 62 290 63 291 
<< m2c >>
rect 62 290 63 291 
<< m1 >>
rect 62 290 63 291 
<< m2 >>
rect 62 290 63 291 
<< m1 >>
rect 64 290 65 291 
<< m2 >>
rect 64 290 65 291 
<< m2c >>
rect 64 290 65 291 
<< m1 >>
rect 64 290 65 291 
<< m2 >>
rect 64 290 65 291 
<< m1 >>
rect 67 290 68 291 
<< m2 >>
rect 67 290 68 291 
<< m2c >>
rect 67 290 68 291 
<< m1 >>
rect 67 290 68 291 
<< m2 >>
rect 67 290 68 291 
<< m1 >>
rect 73 290 74 291 
<< m2 >>
rect 73 290 74 291 
<< m2c >>
rect 73 290 74 291 
<< m1 >>
rect 73 290 74 291 
<< m2 >>
rect 73 290 74 291 
<< m1 >>
rect 132 290 133 291 
<< m2 >>
rect 132 290 133 291 
<< m2c >>
rect 132 290 133 291 
<< m1 >>
rect 132 290 133 291 
<< m2 >>
rect 132 290 133 291 
<< m1 >>
rect 134 290 135 291 
<< m2 >>
rect 134 290 135 291 
<< m2c >>
rect 134 290 135 291 
<< m1 >>
rect 134 290 135 291 
<< m2 >>
rect 134 290 135 291 
<< m2 >>
rect 135 290 136 291 
<< m1 >>
rect 136 290 137 291 
<< m2 >>
rect 136 290 137 291 
<< m2 >>
rect 137 290 138 291 
<< m1 >>
rect 163 290 164 291 
<< m1 >>
rect 165 290 166 291 
<< m2 >>
rect 166 290 167 291 
<< m1 >>
rect 171 290 172 291 
<< m1 >>
rect 181 290 182 291 
<< m1 >>
rect 190 290 191 291 
<< m1 >>
rect 199 290 200 291 
<< m2 >>
rect 200 290 201 291 
<< m1 >>
rect 214 290 215 291 
<< m1 >>
rect 217 290 218 291 
<< m2 >>
rect 217 290 218 291 
<< m2c >>
rect 217 290 218 291 
<< m1 >>
rect 217 290 218 291 
<< m2 >>
rect 217 290 218 291 
<< m1 >>
rect 223 290 224 291 
<< m2 >>
rect 223 290 224 291 
<< m2c >>
rect 223 290 224 291 
<< m1 >>
rect 223 290 224 291 
<< m2 >>
rect 223 290 224 291 
<< m1 >>
rect 226 290 227 291 
<< m2 >>
rect 226 290 227 291 
<< m2c >>
rect 226 290 227 291 
<< m1 >>
rect 226 290 227 291 
<< m2 >>
rect 226 290 227 291 
<< m2 >>
rect 231 290 232 291 
<< m2 >>
rect 232 290 233 291 
<< m2 >>
rect 233 290 234 291 
<< m2 >>
rect 234 290 235 291 
<< m2 >>
rect 235 290 236 291 
<< m2 >>
rect 236 290 237 291 
<< m1 >>
rect 237 290 238 291 
<< m2 >>
rect 237 290 238 291 
<< m2c >>
rect 237 290 238 291 
<< m1 >>
rect 237 290 238 291 
<< m2 >>
rect 237 290 238 291 
<< m1 >>
rect 239 290 240 291 
<< m2 >>
rect 239 290 240 291 
<< m2c >>
rect 239 290 240 291 
<< m1 >>
rect 239 290 240 291 
<< m2 >>
rect 239 290 240 291 
<< m1 >>
rect 241 290 242 291 
<< m2 >>
rect 241 290 242 291 
<< m2c >>
rect 241 290 242 291 
<< m1 >>
rect 241 290 242 291 
<< m2 >>
rect 241 290 242 291 
<< m1 >>
rect 271 290 272 291 
<< m2 >>
rect 271 290 272 291 
<< m2c >>
rect 271 290 272 291 
<< m1 >>
rect 271 290 272 291 
<< m2 >>
rect 271 290 272 291 
<< m1 >>
rect 272 290 273 291 
<< m1 >>
rect 276 290 277 291 
<< m1 >>
rect 278 290 279 291 
<< m2 >>
rect 316 290 317 291 
<< m2 >>
rect 317 290 318 291 
<< m1 >>
rect 318 290 319 291 
<< m2 >>
rect 318 290 319 291 
<< m2c >>
rect 318 290 319 291 
<< m1 >>
rect 318 290 319 291 
<< m2 >>
rect 318 290 319 291 
<< m1 >>
rect 325 290 326 291 
<< m1 >>
rect 327 290 328 291 
<< m1 >>
rect 331 290 332 291 
<< m1 >>
rect 340 290 341 291 
<< m1 >>
rect 10 291 11 292 
<< m2 >>
rect 28 291 29 292 
<< m2 >>
rect 30 291 31 292 
<< m2 >>
rect 37 291 38 292 
<< m2 >>
rect 46 291 47 292 
<< m2 >>
rect 55 291 56 292 
<< m2 >>
rect 57 291 58 292 
<< m2 >>
rect 60 291 61 292 
<< m2 >>
rect 62 291 63 292 
<< m2 >>
rect 64 291 65 292 
<< m2 >>
rect 67 291 68 292 
<< m2 >>
rect 68 291 69 292 
<< m2 >>
rect 73 291 74 292 
<< m2 >>
rect 74 291 75 292 
<< m2 >>
rect 75 291 76 292 
<< m2 >>
rect 76 291 77 292 
<< m2 >>
rect 77 291 78 292 
<< m2 >>
rect 78 291 79 292 
<< m2 >>
rect 79 291 80 292 
<< m2 >>
rect 80 291 81 292 
<< m2 >>
rect 81 291 82 292 
<< m2 >>
rect 132 291 133 292 
<< m1 >>
rect 136 291 137 292 
<< m2 >>
rect 137 291 138 292 
<< m1 >>
rect 163 291 164 292 
<< m1 >>
rect 165 291 166 292 
<< m2 >>
rect 166 291 167 292 
<< m1 >>
rect 167 291 168 292 
<< m2 >>
rect 167 291 168 292 
<< m2c >>
rect 167 291 168 292 
<< m1 >>
rect 167 291 168 292 
<< m2 >>
rect 167 291 168 292 
<< m1 >>
rect 168 291 169 292 
<< m1 >>
rect 169 291 170 292 
<< m2 >>
rect 169 291 170 292 
<< m2c >>
rect 169 291 170 292 
<< m1 >>
rect 169 291 170 292 
<< m2 >>
rect 169 291 170 292 
<< m1 >>
rect 171 291 172 292 
<< m2 >>
rect 171 291 172 292 
<< m2c >>
rect 171 291 172 292 
<< m1 >>
rect 171 291 172 292 
<< m2 >>
rect 171 291 172 292 
<< m1 >>
rect 181 291 182 292 
<< m2 >>
rect 181 291 182 292 
<< m2c >>
rect 181 291 182 292 
<< m1 >>
rect 181 291 182 292 
<< m2 >>
rect 181 291 182 292 
<< m1 >>
rect 190 291 191 292 
<< m1 >>
rect 191 291 192 292 
<< m1 >>
rect 192 291 193 292 
<< m2 >>
rect 192 291 193 292 
<< m2c >>
rect 192 291 193 292 
<< m1 >>
rect 192 291 193 292 
<< m2 >>
rect 192 291 193 292 
<< m1 >>
rect 199 291 200 292 
<< m2 >>
rect 200 291 201 292 
<< m1 >>
rect 201 291 202 292 
<< m2 >>
rect 201 291 202 292 
<< m2c >>
rect 201 291 202 292 
<< m1 >>
rect 201 291 202 292 
<< m2 >>
rect 201 291 202 292 
<< m1 >>
rect 202 291 203 292 
<< m1 >>
rect 203 291 204 292 
<< m1 >>
rect 204 291 205 292 
<< m1 >>
rect 205 291 206 292 
<< m1 >>
rect 206 291 207 292 
<< m1 >>
rect 207 291 208 292 
<< m1 >>
rect 208 291 209 292 
<< m1 >>
rect 209 291 210 292 
<< m1 >>
rect 210 291 211 292 
<< m2 >>
rect 210 291 211 292 
<< m2c >>
rect 210 291 211 292 
<< m1 >>
rect 210 291 211 292 
<< m2 >>
rect 210 291 211 292 
<< m1 >>
rect 214 291 215 292 
<< m2 >>
rect 217 291 218 292 
<< m2 >>
rect 218 291 219 292 
<< m2 >>
rect 219 291 220 292 
<< m2 >>
rect 220 291 221 292 
<< m2 >>
rect 221 291 222 292 
<< m2 >>
rect 223 291 224 292 
<< m2 >>
rect 226 291 227 292 
<< m2 >>
rect 231 291 232 292 
<< m2 >>
rect 239 291 240 292 
<< m2 >>
rect 241 291 242 292 
<< m2 >>
rect 271 291 272 292 
<< m1 >>
rect 276 291 277 292 
<< m1 >>
rect 278 291 279 292 
<< m1 >>
rect 318 291 319 292 
<< m1 >>
rect 325 291 326 292 
<< m1 >>
rect 327 291 328 292 
<< m1 >>
rect 331 291 332 292 
<< m1 >>
rect 340 291 341 292 
<< m1 >>
rect 10 292 11 293 
<< m1 >>
rect 13 292 14 293 
<< m1 >>
rect 14 292 15 293 
<< m1 >>
rect 15 292 16 293 
<< m1 >>
rect 16 292 17 293 
<< m1 >>
rect 17 292 18 293 
<< m1 >>
rect 18 292 19 293 
<< m1 >>
rect 19 292 20 293 
<< m1 >>
rect 20 292 21 293 
<< m1 >>
rect 21 292 22 293 
<< m1 >>
rect 22 292 23 293 
<< m1 >>
rect 23 292 24 293 
<< m1 >>
rect 24 292 25 293 
<< m1 >>
rect 25 292 26 293 
<< m1 >>
rect 26 292 27 293 
<< m1 >>
rect 27 292 28 293 
<< m1 >>
rect 28 292 29 293 
<< m2 >>
rect 28 292 29 293 
<< m1 >>
rect 29 292 30 293 
<< m1 >>
rect 30 292 31 293 
<< m2 >>
rect 30 292 31 293 
<< m1 >>
rect 31 292 32 293 
<< m1 >>
rect 32 292 33 293 
<< m1 >>
rect 33 292 34 293 
<< m1 >>
rect 34 292 35 293 
<< m1 >>
rect 35 292 36 293 
<< m1 >>
rect 36 292 37 293 
<< m1 >>
rect 37 292 38 293 
<< m2 >>
rect 37 292 38 293 
<< m1 >>
rect 38 292 39 293 
<< m1 >>
rect 39 292 40 293 
<< m1 >>
rect 40 292 41 293 
<< m1 >>
rect 41 292 42 293 
<< m1 >>
rect 42 292 43 293 
<< m1 >>
rect 43 292 44 293 
<< m1 >>
rect 44 292 45 293 
<< m1 >>
rect 45 292 46 293 
<< m1 >>
rect 46 292 47 293 
<< m2 >>
rect 46 292 47 293 
<< m1 >>
rect 47 292 48 293 
<< m1 >>
rect 48 292 49 293 
<< m1 >>
rect 49 292 50 293 
<< m1 >>
rect 50 292 51 293 
<< m1 >>
rect 51 292 52 293 
<< m1 >>
rect 52 292 53 293 
<< m1 >>
rect 53 292 54 293 
<< m1 >>
rect 54 292 55 293 
<< m1 >>
rect 55 292 56 293 
<< m2 >>
rect 55 292 56 293 
<< m1 >>
rect 56 292 57 293 
<< m1 >>
rect 57 292 58 293 
<< m2 >>
rect 57 292 58 293 
<< m1 >>
rect 58 292 59 293 
<< m1 >>
rect 59 292 60 293 
<< m1 >>
rect 60 292 61 293 
<< m2 >>
rect 60 292 61 293 
<< m1 >>
rect 61 292 62 293 
<< m1 >>
rect 62 292 63 293 
<< m2 >>
rect 62 292 63 293 
<< m1 >>
rect 63 292 64 293 
<< m1 >>
rect 64 292 65 293 
<< m2 >>
rect 64 292 65 293 
<< m1 >>
rect 65 292 66 293 
<< m1 >>
rect 66 292 67 293 
<< m1 >>
rect 67 292 68 293 
<< m1 >>
rect 68 292 69 293 
<< m2 >>
rect 68 292 69 293 
<< m1 >>
rect 69 292 70 293 
<< m1 >>
rect 70 292 71 293 
<< m1 >>
rect 71 292 72 293 
<< m1 >>
rect 72 292 73 293 
<< m1 >>
rect 73 292 74 293 
<< m1 >>
rect 74 292 75 293 
<< m1 >>
rect 75 292 76 293 
<< m1 >>
rect 76 292 77 293 
<< m1 >>
rect 77 292 78 293 
<< m1 >>
rect 78 292 79 293 
<< m1 >>
rect 79 292 80 293 
<< m1 >>
rect 80 292 81 293 
<< m1 >>
rect 81 292 82 293 
<< m2 >>
rect 81 292 82 293 
<< m1 >>
rect 82 292 83 293 
<< m1 >>
rect 83 292 84 293 
<< m1 >>
rect 84 292 85 293 
<< m2 >>
rect 84 292 85 293 
<< m1 >>
rect 85 292 86 293 
<< m2 >>
rect 85 292 86 293 
<< m1 >>
rect 86 292 87 293 
<< m2 >>
rect 86 292 87 293 
<< m1 >>
rect 87 292 88 293 
<< m2 >>
rect 87 292 88 293 
<< m1 >>
rect 88 292 89 293 
<< m2 >>
rect 88 292 89 293 
<< m1 >>
rect 89 292 90 293 
<< m2 >>
rect 89 292 90 293 
<< m1 >>
rect 90 292 91 293 
<< m2 >>
rect 90 292 91 293 
<< m1 >>
rect 91 292 92 293 
<< m2 >>
rect 91 292 92 293 
<< m1 >>
rect 92 292 93 293 
<< m2 >>
rect 92 292 93 293 
<< m1 >>
rect 93 292 94 293 
<< m2 >>
rect 93 292 94 293 
<< m1 >>
rect 94 292 95 293 
<< m2 >>
rect 94 292 95 293 
<< m1 >>
rect 95 292 96 293 
<< m2 >>
rect 95 292 96 293 
<< m1 >>
rect 96 292 97 293 
<< m2 >>
rect 96 292 97 293 
<< m1 >>
rect 97 292 98 293 
<< m2 >>
rect 97 292 98 293 
<< m1 >>
rect 98 292 99 293 
<< m2 >>
rect 98 292 99 293 
<< m1 >>
rect 99 292 100 293 
<< m2 >>
rect 99 292 100 293 
<< m1 >>
rect 100 292 101 293 
<< m2 >>
rect 100 292 101 293 
<< m1 >>
rect 101 292 102 293 
<< m2 >>
rect 101 292 102 293 
<< m1 >>
rect 102 292 103 293 
<< m2 >>
rect 102 292 103 293 
<< m1 >>
rect 103 292 104 293 
<< m2 >>
rect 103 292 104 293 
<< m1 >>
rect 104 292 105 293 
<< m2 >>
rect 104 292 105 293 
<< m1 >>
rect 105 292 106 293 
<< m2 >>
rect 105 292 106 293 
<< m1 >>
rect 106 292 107 293 
<< m2 >>
rect 106 292 107 293 
<< m1 >>
rect 107 292 108 293 
<< m2 >>
rect 107 292 108 293 
<< m1 >>
rect 108 292 109 293 
<< m2 >>
rect 108 292 109 293 
<< m1 >>
rect 109 292 110 293 
<< m2 >>
rect 109 292 110 293 
<< m1 >>
rect 110 292 111 293 
<< m2 >>
rect 110 292 111 293 
<< m1 >>
rect 111 292 112 293 
<< m2 >>
rect 111 292 112 293 
<< m1 >>
rect 112 292 113 293 
<< m2 >>
rect 112 292 113 293 
<< m1 >>
rect 113 292 114 293 
<< m2 >>
rect 113 292 114 293 
<< m1 >>
rect 114 292 115 293 
<< m2 >>
rect 114 292 115 293 
<< m1 >>
rect 115 292 116 293 
<< m2 >>
rect 115 292 116 293 
<< m1 >>
rect 116 292 117 293 
<< m2 >>
rect 116 292 117 293 
<< m1 >>
rect 117 292 118 293 
<< m2 >>
rect 117 292 118 293 
<< m1 >>
rect 118 292 119 293 
<< m2 >>
rect 118 292 119 293 
<< m1 >>
rect 119 292 120 293 
<< m2 >>
rect 119 292 120 293 
<< m1 >>
rect 120 292 121 293 
<< m2 >>
rect 120 292 121 293 
<< m1 >>
rect 121 292 122 293 
<< m2 >>
rect 121 292 122 293 
<< m1 >>
rect 122 292 123 293 
<< m2 >>
rect 122 292 123 293 
<< m1 >>
rect 123 292 124 293 
<< m2 >>
rect 123 292 124 293 
<< m1 >>
rect 124 292 125 293 
<< m2 >>
rect 124 292 125 293 
<< m1 >>
rect 125 292 126 293 
<< m2 >>
rect 125 292 126 293 
<< m1 >>
rect 126 292 127 293 
<< m2 >>
rect 126 292 127 293 
<< m1 >>
rect 127 292 128 293 
<< m2 >>
rect 127 292 128 293 
<< m1 >>
rect 128 292 129 293 
<< m2 >>
rect 128 292 129 293 
<< m1 >>
rect 129 292 130 293 
<< m2 >>
rect 129 292 130 293 
<< m1 >>
rect 130 292 131 293 
<< m2 >>
rect 130 292 131 293 
<< m1 >>
rect 131 292 132 293 
<< m2 >>
rect 131 292 132 293 
<< m1 >>
rect 132 292 133 293 
<< m2 >>
rect 132 292 133 293 
<< m1 >>
rect 133 292 134 293 
<< m1 >>
rect 134 292 135 293 
<< m1 >>
rect 135 292 136 293 
<< m1 >>
rect 136 292 137 293 
<< m2 >>
rect 137 292 138 293 
<< m1 >>
rect 163 292 164 293 
<< m1 >>
rect 165 292 166 293 
<< m2 >>
rect 169 292 170 293 
<< m2 >>
rect 171 292 172 293 
<< m2 >>
rect 181 292 182 293 
<< m2 >>
rect 192 292 193 293 
<< m1 >>
rect 199 292 200 293 
<< m2 >>
rect 210 292 211 293 
<< m1 >>
rect 214 292 215 293 
<< m1 >>
rect 215 292 216 293 
<< m1 >>
rect 216 292 217 293 
<< m1 >>
rect 217 292 218 293 
<< m1 >>
rect 218 292 219 293 
<< m1 >>
rect 219 292 220 293 
<< m1 >>
rect 220 292 221 293 
<< m1 >>
rect 221 292 222 293 
<< m2 >>
rect 221 292 222 293 
<< m1 >>
rect 222 292 223 293 
<< m1 >>
rect 223 292 224 293 
<< m2 >>
rect 223 292 224 293 
<< m1 >>
rect 224 292 225 293 
<< m1 >>
rect 225 292 226 293 
<< m1 >>
rect 226 292 227 293 
<< m2 >>
rect 226 292 227 293 
<< m1 >>
rect 227 292 228 293 
<< m1 >>
rect 228 292 229 293 
<< m1 >>
rect 229 292 230 293 
<< m1 >>
rect 230 292 231 293 
<< m1 >>
rect 231 292 232 293 
<< m2 >>
rect 231 292 232 293 
<< m1 >>
rect 232 292 233 293 
<< m1 >>
rect 233 292 234 293 
<< m1 >>
rect 234 292 235 293 
<< m1 >>
rect 235 292 236 293 
<< m1 >>
rect 236 292 237 293 
<< m1 >>
rect 237 292 238 293 
<< m1 >>
rect 238 292 239 293 
<< m1 >>
rect 239 292 240 293 
<< m2 >>
rect 239 292 240 293 
<< m1 >>
rect 240 292 241 293 
<< m1 >>
rect 241 292 242 293 
<< m2 >>
rect 241 292 242 293 
<< m1 >>
rect 242 292 243 293 
<< m2 >>
rect 242 292 243 293 
<< m1 >>
rect 243 292 244 293 
<< m2 >>
rect 243 292 244 293 
<< m1 >>
rect 244 292 245 293 
<< m2 >>
rect 244 292 245 293 
<< m1 >>
rect 245 292 246 293 
<< m2 >>
rect 245 292 246 293 
<< m1 >>
rect 246 292 247 293 
<< m2 >>
rect 246 292 247 293 
<< m1 >>
rect 247 292 248 293 
<< m2 >>
rect 247 292 248 293 
<< m1 >>
rect 248 292 249 293 
<< m2 >>
rect 248 292 249 293 
<< m1 >>
rect 249 292 250 293 
<< m1 >>
rect 250 292 251 293 
<< m1 >>
rect 251 292 252 293 
<< m1 >>
rect 252 292 253 293 
<< m1 >>
rect 253 292 254 293 
<< m1 >>
rect 254 292 255 293 
<< m1 >>
rect 255 292 256 293 
<< m1 >>
rect 256 292 257 293 
<< m1 >>
rect 257 292 258 293 
<< m1 >>
rect 258 292 259 293 
<< m1 >>
rect 259 292 260 293 
<< m1 >>
rect 260 292 261 293 
<< m1 >>
rect 261 292 262 293 
<< m1 >>
rect 262 292 263 293 
<< m1 >>
rect 263 292 264 293 
<< m1 >>
rect 264 292 265 293 
<< m1 >>
rect 265 292 266 293 
<< m1 >>
rect 266 292 267 293 
<< m1 >>
rect 267 292 268 293 
<< m1 >>
rect 268 292 269 293 
<< m1 >>
rect 269 292 270 293 
<< m1 >>
rect 270 292 271 293 
<< m1 >>
rect 271 292 272 293 
<< m2 >>
rect 271 292 272 293 
<< m1 >>
rect 276 292 277 293 
<< m1 >>
rect 278 292 279 293 
<< m1 >>
rect 318 292 319 293 
<< m1 >>
rect 325 292 326 293 
<< m1 >>
rect 327 292 328 293 
<< m1 >>
rect 331 292 332 293 
<< m1 >>
rect 334 292 335 293 
<< m1 >>
rect 335 292 336 293 
<< m1 >>
rect 336 292 337 293 
<< m1 >>
rect 337 292 338 293 
<< m1 >>
rect 338 292 339 293 
<< m1 >>
rect 339 292 340 293 
<< m1 >>
rect 340 292 341 293 
<< m1 >>
rect 10 293 11 294 
<< m1 >>
rect 13 293 14 294 
<< m2 >>
rect 28 293 29 294 
<< m2 >>
rect 30 293 31 294 
<< m2 >>
rect 31 293 32 294 
<< m2 >>
rect 32 293 33 294 
<< m2 >>
rect 33 293 34 294 
<< m2 >>
rect 34 293 35 294 
<< m2 >>
rect 35 293 36 294 
<< m2 >>
rect 37 293 38 294 
<< m2 >>
rect 46 293 47 294 
<< m2 >>
rect 55 293 56 294 
<< m2 >>
rect 57 293 58 294 
<< m2 >>
rect 60 293 61 294 
<< m2 >>
rect 62 293 63 294 
<< m2 >>
rect 64 293 65 294 
<< m2 >>
rect 68 293 69 294 
<< m2 >>
rect 81 293 82 294 
<< m2 >>
rect 84 293 85 294 
<< m2 >>
rect 137 293 138 294 
<< m1 >>
rect 163 293 164 294 
<< m2 >>
rect 163 293 164 294 
<< m2c >>
rect 163 293 164 294 
<< m1 >>
rect 163 293 164 294 
<< m2 >>
rect 163 293 164 294 
<< m2 >>
rect 164 293 165 294 
<< m1 >>
rect 165 293 166 294 
<< m2 >>
rect 165 293 166 294 
<< m2 >>
rect 166 293 167 294 
<< m1 >>
rect 167 293 168 294 
<< m2 >>
rect 167 293 168 294 
<< m2c >>
rect 167 293 168 294 
<< m1 >>
rect 167 293 168 294 
<< m2 >>
rect 167 293 168 294 
<< m1 >>
rect 168 293 169 294 
<< m1 >>
rect 169 293 170 294 
<< m2 >>
rect 169 293 170 294 
<< m1 >>
rect 170 293 171 294 
<< m1 >>
rect 171 293 172 294 
<< m2 >>
rect 171 293 172 294 
<< m1 >>
rect 172 293 173 294 
<< m1 >>
rect 173 293 174 294 
<< m1 >>
rect 174 293 175 294 
<< m1 >>
rect 175 293 176 294 
<< m1 >>
rect 176 293 177 294 
<< m1 >>
rect 177 293 178 294 
<< m1 >>
rect 178 293 179 294 
<< m1 >>
rect 179 293 180 294 
<< m1 >>
rect 180 293 181 294 
<< m1 >>
rect 181 293 182 294 
<< m2 >>
rect 181 293 182 294 
<< m1 >>
rect 182 293 183 294 
<< m1 >>
rect 183 293 184 294 
<< m1 >>
rect 184 293 185 294 
<< m1 >>
rect 185 293 186 294 
<< m1 >>
rect 186 293 187 294 
<< m1 >>
rect 187 293 188 294 
<< m1 >>
rect 188 293 189 294 
<< m1 >>
rect 189 293 190 294 
<< m1 >>
rect 190 293 191 294 
<< m1 >>
rect 191 293 192 294 
<< m1 >>
rect 192 293 193 294 
<< m2 >>
rect 192 293 193 294 
<< m1 >>
rect 193 293 194 294 
<< m2 >>
rect 193 293 194 294 
<< m1 >>
rect 194 293 195 294 
<< m2 >>
rect 194 293 195 294 
<< m1 >>
rect 195 293 196 294 
<< m2 >>
rect 195 293 196 294 
<< m1 >>
rect 196 293 197 294 
<< m2 >>
rect 196 293 197 294 
<< m1 >>
rect 197 293 198 294 
<< m2 >>
rect 197 293 198 294 
<< m2 >>
rect 198 293 199 294 
<< m1 >>
rect 199 293 200 294 
<< m2 >>
rect 199 293 200 294 
<< m2 >>
rect 200 293 201 294 
<< m1 >>
rect 201 293 202 294 
<< m2 >>
rect 201 293 202 294 
<< m2c >>
rect 201 293 202 294 
<< m1 >>
rect 201 293 202 294 
<< m2 >>
rect 201 293 202 294 
<< m1 >>
rect 202 293 203 294 
<< m1 >>
rect 203 293 204 294 
<< m1 >>
rect 204 293 205 294 
<< m1 >>
rect 205 293 206 294 
<< m1 >>
rect 206 293 207 294 
<< m1 >>
rect 207 293 208 294 
<< m1 >>
rect 208 293 209 294 
<< m1 >>
rect 209 293 210 294 
<< m1 >>
rect 210 293 211 294 
<< m2 >>
rect 210 293 211 294 
<< m1 >>
rect 211 293 212 294 
<< m1 >>
rect 212 293 213 294 
<< m2 >>
rect 212 293 213 294 
<< m2c >>
rect 212 293 213 294 
<< m1 >>
rect 212 293 213 294 
<< m2 >>
rect 212 293 213 294 
<< m2 >>
rect 213 293 214 294 
<< m2 >>
rect 214 293 215 294 
<< m2 >>
rect 215 293 216 294 
<< m2 >>
rect 216 293 217 294 
<< m2 >>
rect 217 293 218 294 
<< m2 >>
rect 218 293 219 294 
<< m2 >>
rect 219 293 220 294 
<< m2 >>
rect 221 293 222 294 
<< m2 >>
rect 223 293 224 294 
<< m2 >>
rect 226 293 227 294 
<< m2 >>
rect 231 293 232 294 
<< m2 >>
rect 239 293 240 294 
<< m2 >>
rect 248 293 249 294 
<< m1 >>
rect 271 293 272 294 
<< m2 >>
rect 271 293 272 294 
<< m1 >>
rect 276 293 277 294 
<< m1 >>
rect 278 293 279 294 
<< m1 >>
rect 318 293 319 294 
<< m1 >>
rect 325 293 326 294 
<< m1 >>
rect 327 293 328 294 
<< m1 >>
rect 331 293 332 294 
<< m1 >>
rect 334 293 335 294 
<< m1 >>
rect 10 294 11 295 
<< m1 >>
rect 13 294 14 295 
<< m1 >>
rect 28 294 29 295 
<< m2 >>
rect 28 294 29 295 
<< m2c >>
rect 28 294 29 295 
<< m1 >>
rect 28 294 29 295 
<< m2 >>
rect 28 294 29 295 
<< m1 >>
rect 35 294 36 295 
<< m2 >>
rect 35 294 36 295 
<< m2c >>
rect 35 294 36 295 
<< m1 >>
rect 35 294 36 295 
<< m2 >>
rect 35 294 36 295 
<< m1 >>
rect 37 294 38 295 
<< m2 >>
rect 37 294 38 295 
<< m2c >>
rect 37 294 38 295 
<< m1 >>
rect 37 294 38 295 
<< m2 >>
rect 37 294 38 295 
<< m1 >>
rect 46 294 47 295 
<< m2 >>
rect 46 294 47 295 
<< m2c >>
rect 46 294 47 295 
<< m1 >>
rect 46 294 47 295 
<< m2 >>
rect 46 294 47 295 
<< m2 >>
rect 55 294 56 295 
<< m2 >>
rect 57 294 58 295 
<< m2 >>
rect 60 294 61 295 
<< m2 >>
rect 62 294 63 295 
<< m2 >>
rect 64 294 65 295 
<< m2 >>
rect 68 294 69 295 
<< m2 >>
rect 81 294 82 295 
<< m2 >>
rect 84 294 85 295 
<< m2 >>
rect 137 294 138 295 
<< m1 >>
rect 165 294 166 295 
<< m2 >>
rect 169 294 170 295 
<< m2 >>
rect 171 294 172 295 
<< m2 >>
rect 181 294 182 295 
<< m1 >>
rect 197 294 198 295 
<< m1 >>
rect 199 294 200 295 
<< m2 >>
rect 210 294 211 295 
<< m1 >>
rect 219 294 220 295 
<< m2 >>
rect 219 294 220 295 
<< m2c >>
rect 219 294 220 295 
<< m1 >>
rect 219 294 220 295 
<< m2 >>
rect 219 294 220 295 
<< m1 >>
rect 221 294 222 295 
<< m2 >>
rect 221 294 222 295 
<< m2c >>
rect 221 294 222 295 
<< m1 >>
rect 221 294 222 295 
<< m2 >>
rect 221 294 222 295 
<< m1 >>
rect 223 294 224 295 
<< m2 >>
rect 223 294 224 295 
<< m2c >>
rect 223 294 224 295 
<< m1 >>
rect 223 294 224 295 
<< m2 >>
rect 223 294 224 295 
<< m1 >>
rect 226 294 227 295 
<< m2 >>
rect 226 294 227 295 
<< m2c >>
rect 226 294 227 295 
<< m1 >>
rect 226 294 227 295 
<< m2 >>
rect 226 294 227 295 
<< m1 >>
rect 227 294 228 295 
<< m1 >>
rect 228 294 229 295 
<< m1 >>
rect 229 294 230 295 
<< m1 >>
rect 230 294 231 295 
<< m1 >>
rect 231 294 232 295 
<< m2 >>
rect 231 294 232 295 
<< m1 >>
rect 232 294 233 295 
<< m1 >>
rect 233 294 234 295 
<< m1 >>
rect 234 294 235 295 
<< m1 >>
rect 235 294 236 295 
<< m1 >>
rect 236 294 237 295 
<< m1 >>
rect 237 294 238 295 
<< m1 >>
rect 238 294 239 295 
<< m1 >>
rect 239 294 240 295 
<< m2 >>
rect 239 294 240 295 
<< m1 >>
rect 240 294 241 295 
<< m1 >>
rect 241 294 242 295 
<< m1 >>
rect 242 294 243 295 
<< m1 >>
rect 243 294 244 295 
<< m1 >>
rect 244 294 245 295 
<< m1 >>
rect 245 294 246 295 
<< m1 >>
rect 246 294 247 295 
<< m1 >>
rect 247 294 248 295 
<< m1 >>
rect 248 294 249 295 
<< m2 >>
rect 248 294 249 295 
<< m1 >>
rect 249 294 250 295 
<< m1 >>
rect 250 294 251 295 
<< m1 >>
rect 251 294 252 295 
<< m1 >>
rect 252 294 253 295 
<< m1 >>
rect 253 294 254 295 
<< m1 >>
rect 254 294 255 295 
<< m1 >>
rect 255 294 256 295 
<< m1 >>
rect 256 294 257 295 
<< m1 >>
rect 257 294 258 295 
<< m1 >>
rect 258 294 259 295 
<< m1 >>
rect 259 294 260 295 
<< m1 >>
rect 260 294 261 295 
<< m1 >>
rect 261 294 262 295 
<< m1 >>
rect 262 294 263 295 
<< m1 >>
rect 263 294 264 295 
<< m1 >>
rect 264 294 265 295 
<< m1 >>
rect 265 294 266 295 
<< m1 >>
rect 271 294 272 295 
<< m2 >>
rect 271 294 272 295 
<< m1 >>
rect 276 294 277 295 
<< m1 >>
rect 278 294 279 295 
<< m1 >>
rect 318 294 319 295 
<< m1 >>
rect 325 294 326 295 
<< m1 >>
rect 327 294 328 295 
<< m1 >>
rect 331 294 332 295 
<< m1 >>
rect 334 294 335 295 
<< m1 >>
rect 10 295 11 296 
<< m1 >>
rect 13 295 14 296 
<< m1 >>
rect 28 295 29 296 
<< m1 >>
rect 35 295 36 296 
<< m1 >>
rect 37 295 38 296 
<< m1 >>
rect 46 295 47 296 
<< m1 >>
rect 55 295 56 296 
<< m2 >>
rect 55 295 56 296 
<< m1 >>
rect 56 295 57 296 
<< m1 >>
rect 57 295 58 296 
<< m2 >>
rect 57 295 58 296 
<< m1 >>
rect 58 295 59 296 
<< m1 >>
rect 59 295 60 296 
<< m1 >>
rect 60 295 61 296 
<< m2 >>
rect 60 295 61 296 
<< m1 >>
rect 61 295 62 296 
<< m1 >>
rect 62 295 63 296 
<< m2 >>
rect 62 295 63 296 
<< m1 >>
rect 63 295 64 296 
<< m1 >>
rect 64 295 65 296 
<< m2 >>
rect 64 295 65 296 
<< m1 >>
rect 65 295 66 296 
<< m1 >>
rect 66 295 67 296 
<< m1 >>
rect 67 295 68 296 
<< m1 >>
rect 68 295 69 296 
<< m2 >>
rect 68 295 69 296 
<< m1 >>
rect 69 295 70 296 
<< m1 >>
rect 70 295 71 296 
<< m1 >>
rect 71 295 72 296 
<< m1 >>
rect 72 295 73 296 
<< m1 >>
rect 73 295 74 296 
<< m1 >>
rect 74 295 75 296 
<< m1 >>
rect 75 295 76 296 
<< m1 >>
rect 76 295 77 296 
<< m1 >>
rect 77 295 78 296 
<< m1 >>
rect 78 295 79 296 
<< m1 >>
rect 79 295 80 296 
<< m1 >>
rect 80 295 81 296 
<< m1 >>
rect 81 295 82 296 
<< m2 >>
rect 81 295 82 296 
<< m1 >>
rect 82 295 83 296 
<< m1 >>
rect 83 295 84 296 
<< m1 >>
rect 84 295 85 296 
<< m2 >>
rect 84 295 85 296 
<< m1 >>
rect 85 295 86 296 
<< m1 >>
rect 86 295 87 296 
<< m1 >>
rect 87 295 88 296 
<< m1 >>
rect 88 295 89 296 
<< m1 >>
rect 89 295 90 296 
<< m1 >>
rect 90 295 91 296 
<< m1 >>
rect 91 295 92 296 
<< m1 >>
rect 92 295 93 296 
<< m1 >>
rect 93 295 94 296 
<< m1 >>
rect 94 295 95 296 
<< m1 >>
rect 95 295 96 296 
<< m1 >>
rect 96 295 97 296 
<< m1 >>
rect 97 295 98 296 
<< m1 >>
rect 98 295 99 296 
<< m1 >>
rect 99 295 100 296 
<< m1 >>
rect 100 295 101 296 
<< m1 >>
rect 101 295 102 296 
<< m1 >>
rect 102 295 103 296 
<< m1 >>
rect 103 295 104 296 
<< m1 >>
rect 104 295 105 296 
<< m1 >>
rect 105 295 106 296 
<< m1 >>
rect 106 295 107 296 
<< m1 >>
rect 107 295 108 296 
<< m1 >>
rect 108 295 109 296 
<< m1 >>
rect 109 295 110 296 
<< m1 >>
rect 110 295 111 296 
<< m1 >>
rect 111 295 112 296 
<< m1 >>
rect 112 295 113 296 
<< m1 >>
rect 113 295 114 296 
<< m1 >>
rect 114 295 115 296 
<< m1 >>
rect 115 295 116 296 
<< m1 >>
rect 116 295 117 296 
<< m1 >>
rect 117 295 118 296 
<< m1 >>
rect 118 295 119 296 
<< m1 >>
rect 119 295 120 296 
<< m1 >>
rect 120 295 121 296 
<< m1 >>
rect 121 295 122 296 
<< m1 >>
rect 122 295 123 296 
<< m1 >>
rect 123 295 124 296 
<< m1 >>
rect 124 295 125 296 
<< m1 >>
rect 125 295 126 296 
<< m1 >>
rect 126 295 127 296 
<< m1 >>
rect 127 295 128 296 
<< m1 >>
rect 128 295 129 296 
<< m1 >>
rect 129 295 130 296 
<< m1 >>
rect 130 295 131 296 
<< m1 >>
rect 131 295 132 296 
<< m1 >>
rect 132 295 133 296 
<< m1 >>
rect 133 295 134 296 
<< m1 >>
rect 134 295 135 296 
<< m1 >>
rect 135 295 136 296 
<< m1 >>
rect 136 295 137 296 
<< m1 >>
rect 137 295 138 296 
<< m2 >>
rect 137 295 138 296 
<< m1 >>
rect 138 295 139 296 
<< m2 >>
rect 138 295 139 296 
<< m1 >>
rect 139 295 140 296 
<< m2 >>
rect 139 295 140 296 
<< m1 >>
rect 140 295 141 296 
<< m2 >>
rect 140 295 141 296 
<< m1 >>
rect 141 295 142 296 
<< m2 >>
rect 141 295 142 296 
<< m1 >>
rect 142 295 143 296 
<< m2 >>
rect 142 295 143 296 
<< m1 >>
rect 143 295 144 296 
<< m2 >>
rect 143 295 144 296 
<< m1 >>
rect 144 295 145 296 
<< m2 >>
rect 144 295 145 296 
<< m1 >>
rect 145 295 146 296 
<< m2 >>
rect 145 295 146 296 
<< m1 >>
rect 146 295 147 296 
<< m2 >>
rect 146 295 147 296 
<< m1 >>
rect 147 295 148 296 
<< m2 >>
rect 147 295 148 296 
<< m1 >>
rect 148 295 149 296 
<< m2 >>
rect 148 295 149 296 
<< m1 >>
rect 149 295 150 296 
<< m2 >>
rect 149 295 150 296 
<< m1 >>
rect 150 295 151 296 
<< m2 >>
rect 150 295 151 296 
<< m1 >>
rect 151 295 152 296 
<< m2 >>
rect 151 295 152 296 
<< m1 >>
rect 152 295 153 296 
<< m2 >>
rect 152 295 153 296 
<< m1 >>
rect 153 295 154 296 
<< m2 >>
rect 153 295 154 296 
<< m1 >>
rect 154 295 155 296 
<< m2 >>
rect 154 295 155 296 
<< m1 >>
rect 155 295 156 296 
<< m2 >>
rect 155 295 156 296 
<< m1 >>
rect 156 295 157 296 
<< m2 >>
rect 156 295 157 296 
<< m1 >>
rect 157 295 158 296 
<< m2 >>
rect 157 295 158 296 
<< m1 >>
rect 158 295 159 296 
<< m2 >>
rect 158 295 159 296 
<< m1 >>
rect 159 295 160 296 
<< m2 >>
rect 159 295 160 296 
<< m1 >>
rect 160 295 161 296 
<< m2 >>
rect 160 295 161 296 
<< m1 >>
rect 161 295 162 296 
<< m2 >>
rect 161 295 162 296 
<< m1 >>
rect 162 295 163 296 
<< m2 >>
rect 162 295 163 296 
<< m1 >>
rect 163 295 164 296 
<< m2 >>
rect 163 295 164 296 
<< m1 >>
rect 164 295 165 296 
<< m2 >>
rect 164 295 165 296 
<< m1 >>
rect 165 295 166 296 
<< m2 >>
rect 165 295 166 296 
<< m2 >>
rect 166 295 167 296 
<< m2 >>
rect 169 295 170 296 
<< m2 >>
rect 171 295 172 296 
<< m1 >>
rect 181 295 182 296 
<< m2 >>
rect 181 295 182 296 
<< m2c >>
rect 181 295 182 296 
<< m1 >>
rect 181 295 182 296 
<< m2 >>
rect 181 295 182 296 
<< m1 >>
rect 197 295 198 296 
<< m2 >>
rect 197 295 198 296 
<< m2c >>
rect 197 295 198 296 
<< m1 >>
rect 197 295 198 296 
<< m2 >>
rect 197 295 198 296 
<< m2 >>
rect 198 295 199 296 
<< m1 >>
rect 199 295 200 296 
<< m2 >>
rect 199 295 200 296 
<< m2 >>
rect 200 295 201 296 
<< m1 >>
rect 203 295 204 296 
<< m1 >>
rect 204 295 205 296 
<< m1 >>
rect 205 295 206 296 
<< m1 >>
rect 206 295 207 296 
<< m1 >>
rect 207 295 208 296 
<< m1 >>
rect 208 295 209 296 
<< m1 >>
rect 209 295 210 296 
<< m1 >>
rect 210 295 211 296 
<< m2 >>
rect 210 295 211 296 
<< m1 >>
rect 211 295 212 296 
<< m2 >>
rect 211 295 212 296 
<< m1 >>
rect 212 295 213 296 
<< m2 >>
rect 212 295 213 296 
<< m2 >>
rect 213 295 214 296 
<< m2 >>
rect 214 295 215 296 
<< m2 >>
rect 215 295 216 296 
<< m2 >>
rect 216 295 217 296 
<< m2 >>
rect 217 295 218 296 
<< m2 >>
rect 219 295 220 296 
<< m2 >>
rect 221 295 222 296 
<< m2 >>
rect 223 295 224 296 
<< m2 >>
rect 228 295 229 296 
<< m2 >>
rect 229 295 230 296 
<< m2 >>
rect 230 295 231 296 
<< m2 >>
rect 231 295 232 296 
<< m2 >>
rect 239 295 240 296 
<< m2 >>
rect 248 295 249 296 
<< m1 >>
rect 265 295 266 296 
<< m1 >>
rect 271 295 272 296 
<< m2 >>
rect 271 295 272 296 
<< m1 >>
rect 276 295 277 296 
<< m1 >>
rect 278 295 279 296 
<< m1 >>
rect 318 295 319 296 
<< m1 >>
rect 319 295 320 296 
<< m1 >>
rect 320 295 321 296 
<< m1 >>
rect 321 295 322 296 
<< m1 >>
rect 322 295 323 296 
<< m1 >>
rect 323 295 324 296 
<< m1 >>
rect 325 295 326 296 
<< m1 >>
rect 327 295 328 296 
<< m1 >>
rect 331 295 332 296 
<< m1 >>
rect 334 295 335 296 
<< m1 >>
rect 10 296 11 297 
<< m1 >>
rect 13 296 14 297 
<< m1 >>
rect 28 296 29 297 
<< m1 >>
rect 35 296 36 297 
<< m1 >>
rect 37 296 38 297 
<< m1 >>
rect 46 296 47 297 
<< m1 >>
rect 55 296 56 297 
<< m2 >>
rect 55 296 56 297 
<< m2 >>
rect 57 296 58 297 
<< m2 >>
rect 60 296 61 297 
<< m2 >>
rect 62 296 63 297 
<< m2 >>
rect 64 296 65 297 
<< m2 >>
rect 68 296 69 297 
<< m2 >>
rect 81 296 82 297 
<< m2 >>
rect 84 296 85 297 
<< m2 >>
rect 166 296 167 297 
<< m1 >>
rect 167 296 168 297 
<< m2 >>
rect 167 296 168 297 
<< m2c >>
rect 167 296 168 297 
<< m1 >>
rect 167 296 168 297 
<< m2 >>
rect 167 296 168 297 
<< m1 >>
rect 168 296 169 297 
<< m1 >>
rect 169 296 170 297 
<< m2 >>
rect 169 296 170 297 
<< m1 >>
rect 170 296 171 297 
<< m1 >>
rect 171 296 172 297 
<< m2 >>
rect 171 296 172 297 
<< m1 >>
rect 172 296 173 297 
<< m1 >>
rect 181 296 182 297 
<< m1 >>
rect 199 296 200 297 
<< m2 >>
rect 200 296 201 297 
<< m1 >>
rect 203 296 204 297 
<< m2 >>
rect 203 296 204 297 
<< m2c >>
rect 203 296 204 297 
<< m1 >>
rect 203 296 204 297 
<< m2 >>
rect 203 296 204 297 
<< m1 >>
rect 212 296 213 297 
<< m1 >>
rect 213 296 214 297 
<< m1 >>
rect 214 296 215 297 
<< m1 >>
rect 215 296 216 297 
<< m1 >>
rect 216 296 217 297 
<< m1 >>
rect 217 296 218 297 
<< m2 >>
rect 217 296 218 297 
<< m1 >>
rect 218 296 219 297 
<< m1 >>
rect 219 296 220 297 
<< m2 >>
rect 219 296 220 297 
<< m1 >>
rect 220 296 221 297 
<< m1 >>
rect 221 296 222 297 
<< m2 >>
rect 221 296 222 297 
<< m1 >>
rect 222 296 223 297 
<< m1 >>
rect 223 296 224 297 
<< m2 >>
rect 223 296 224 297 
<< m1 >>
rect 224 296 225 297 
<< m1 >>
rect 225 296 226 297 
<< m1 >>
rect 226 296 227 297 
<< m1 >>
rect 227 296 228 297 
<< m1 >>
rect 228 296 229 297 
<< m2 >>
rect 228 296 229 297 
<< m2c >>
rect 228 296 229 297 
<< m1 >>
rect 228 296 229 297 
<< m2 >>
rect 228 296 229 297 
<< m1 >>
rect 239 296 240 297 
<< m2 >>
rect 239 296 240 297 
<< m2c >>
rect 239 296 240 297 
<< m1 >>
rect 239 296 240 297 
<< m2 >>
rect 239 296 240 297 
<< m2 >>
rect 248 296 249 297 
<< m2 >>
rect 249 296 250 297 
<< m2 >>
rect 250 296 251 297 
<< m2 >>
rect 251 296 252 297 
<< m2 >>
rect 252 296 253 297 
<< m2 >>
rect 253 296 254 297 
<< m2 >>
rect 254 296 255 297 
<< m1 >>
rect 255 296 256 297 
<< m2 >>
rect 255 296 256 297 
<< m2c >>
rect 255 296 256 297 
<< m1 >>
rect 255 296 256 297 
<< m2 >>
rect 255 296 256 297 
<< m1 >>
rect 265 296 266 297 
<< m1 >>
rect 271 296 272 297 
<< m2 >>
rect 271 296 272 297 
<< m1 >>
rect 276 296 277 297 
<< m1 >>
rect 278 296 279 297 
<< m1 >>
rect 323 296 324 297 
<< m1 >>
rect 325 296 326 297 
<< m1 >>
rect 327 296 328 297 
<< m1 >>
rect 331 296 332 297 
<< m1 >>
rect 334 296 335 297 
<< m1 >>
rect 10 297 11 298 
<< m1 >>
rect 13 297 14 298 
<< m1 >>
rect 28 297 29 298 
<< m1 >>
rect 35 297 36 298 
<< m1 >>
rect 37 297 38 298 
<< m1 >>
rect 46 297 47 298 
<< m1 >>
rect 55 297 56 298 
<< m2 >>
rect 55 297 56 298 
<< m1 >>
rect 57 297 58 298 
<< m2 >>
rect 57 297 58 298 
<< m2c >>
rect 57 297 58 298 
<< m1 >>
rect 57 297 58 298 
<< m2 >>
rect 57 297 58 298 
<< m1 >>
rect 60 297 61 298 
<< m2 >>
rect 60 297 61 298 
<< m2c >>
rect 60 297 61 298 
<< m1 >>
rect 60 297 61 298 
<< m2 >>
rect 60 297 61 298 
<< m1 >>
rect 62 297 63 298 
<< m2 >>
rect 62 297 63 298 
<< m2c >>
rect 62 297 63 298 
<< m1 >>
rect 62 297 63 298 
<< m2 >>
rect 62 297 63 298 
<< m1 >>
rect 64 297 65 298 
<< m2 >>
rect 64 297 65 298 
<< m2c >>
rect 64 297 65 298 
<< m1 >>
rect 64 297 65 298 
<< m2 >>
rect 64 297 65 298 
<< m1 >>
rect 68 297 69 298 
<< m2 >>
rect 68 297 69 298 
<< m2c >>
rect 68 297 69 298 
<< m1 >>
rect 68 297 69 298 
<< m2 >>
rect 68 297 69 298 
<< m1 >>
rect 69 297 70 298 
<< m1 >>
rect 70 297 71 298 
<< m1 >>
rect 71 297 72 298 
<< m1 >>
rect 72 297 73 298 
<< m1 >>
rect 73 297 74 298 
<< m2 >>
rect 81 297 82 298 
<< m1 >>
rect 82 297 83 298 
<< m1 >>
rect 83 297 84 298 
<< m1 >>
rect 84 297 85 298 
<< m2 >>
rect 84 297 85 298 
<< m2c >>
rect 84 297 85 298 
<< m1 >>
rect 84 297 85 298 
<< m2 >>
rect 84 297 85 298 
<< m1 >>
rect 103 297 104 298 
<< m1 >>
rect 104 297 105 298 
<< m1 >>
rect 105 297 106 298 
<< m1 >>
rect 106 297 107 298 
<< m1 >>
rect 107 297 108 298 
<< m1 >>
rect 108 297 109 298 
<< m1 >>
rect 109 297 110 298 
<< m2 >>
rect 169 297 170 298 
<< m2 >>
rect 171 297 172 298 
<< m1 >>
rect 172 297 173 298 
<< m1 >>
rect 181 297 182 298 
<< m1 >>
rect 193 297 194 298 
<< m1 >>
rect 194 297 195 298 
<< m1 >>
rect 195 297 196 298 
<< m1 >>
rect 196 297 197 298 
<< m1 >>
rect 197 297 198 298 
<< m1 >>
rect 198 297 199 298 
<< m1 >>
rect 199 297 200 298 
<< m2 >>
rect 200 297 201 298 
<< m2 >>
rect 203 297 204 298 
<< m2 >>
rect 217 297 218 298 
<< m2 >>
rect 219 297 220 298 
<< m2 >>
rect 221 297 222 298 
<< m2 >>
rect 223 297 224 298 
<< m1 >>
rect 239 297 240 298 
<< m1 >>
rect 247 297 248 298 
<< m1 >>
rect 248 297 249 298 
<< m1 >>
rect 249 297 250 298 
<< m1 >>
rect 250 297 251 298 
<< m1 >>
rect 251 297 252 298 
<< m1 >>
rect 252 297 253 298 
<< m1 >>
rect 253 297 254 298 
<< m1 >>
rect 255 297 256 298 
<< m1 >>
rect 265 297 266 298 
<< m1 >>
rect 271 297 272 298 
<< m2 >>
rect 271 297 272 298 
<< m1 >>
rect 276 297 277 298 
<< m1 >>
rect 278 297 279 298 
<< m1 >>
rect 323 297 324 298 
<< m1 >>
rect 325 297 326 298 
<< m1 >>
rect 327 297 328 298 
<< m1 >>
rect 331 297 332 298 
<< m1 >>
rect 334 297 335 298 
<< m1 >>
rect 10 298 11 299 
<< m1 >>
rect 13 298 14 299 
<< m1 >>
rect 28 298 29 299 
<< m1 >>
rect 35 298 36 299 
<< m2 >>
rect 35 298 36 299 
<< m2c >>
rect 35 298 36 299 
<< m1 >>
rect 35 298 36 299 
<< m2 >>
rect 35 298 36 299 
<< m2 >>
rect 36 298 37 299 
<< m1 >>
rect 37 298 38 299 
<< m2 >>
rect 37 298 38 299 
<< m2 >>
rect 38 298 39 299 
<< m1 >>
rect 46 298 47 299 
<< m1 >>
rect 55 298 56 299 
<< m2 >>
rect 55 298 56 299 
<< m1 >>
rect 57 298 58 299 
<< m1 >>
rect 60 298 61 299 
<< m1 >>
rect 62 298 63 299 
<< m1 >>
rect 64 298 65 299 
<< m1 >>
rect 73 298 74 299 
<< m2 >>
rect 81 298 82 299 
<< m1 >>
rect 82 298 83 299 
<< m1 >>
rect 103 298 104 299 
<< m1 >>
rect 109 298 110 299 
<< m1 >>
rect 142 298 143 299 
<< m1 >>
rect 143 298 144 299 
<< m1 >>
rect 144 298 145 299 
<< m1 >>
rect 145 298 146 299 
<< m1 >>
rect 169 298 170 299 
<< m2 >>
rect 169 298 170 299 
<< m2c >>
rect 169 298 170 299 
<< m1 >>
rect 169 298 170 299 
<< m2 >>
rect 169 298 170 299 
<< m2 >>
rect 171 298 172 299 
<< m1 >>
rect 172 298 173 299 
<< m1 >>
rect 181 298 182 299 
<< m1 >>
rect 193 298 194 299 
<< m2 >>
rect 200 298 201 299 
<< m1 >>
rect 201 298 202 299 
<< m2 >>
rect 201 298 202 299 
<< m2c >>
rect 201 298 202 299 
<< m1 >>
rect 201 298 202 299 
<< m2 >>
rect 201 298 202 299 
<< m1 >>
rect 202 298 203 299 
<< m1 >>
rect 203 298 204 299 
<< m2 >>
rect 203 298 204 299 
<< m1 >>
rect 204 298 205 299 
<< m1 >>
rect 205 298 206 299 
<< m1 >>
rect 206 298 207 299 
<< m1 >>
rect 207 298 208 299 
<< m1 >>
rect 208 298 209 299 
<< m1 >>
rect 217 298 218 299 
<< m2 >>
rect 217 298 218 299 
<< m2c >>
rect 217 298 218 299 
<< m1 >>
rect 217 298 218 299 
<< m2 >>
rect 217 298 218 299 
<< m1 >>
rect 219 298 220 299 
<< m2 >>
rect 219 298 220 299 
<< m2c >>
rect 219 298 220 299 
<< m1 >>
rect 219 298 220 299 
<< m2 >>
rect 219 298 220 299 
<< m1 >>
rect 221 298 222 299 
<< m2 >>
rect 221 298 222 299 
<< m2c >>
rect 221 298 222 299 
<< m1 >>
rect 221 298 222 299 
<< m2 >>
rect 221 298 222 299 
<< m1 >>
rect 223 298 224 299 
<< m2 >>
rect 223 298 224 299 
<< m2c >>
rect 223 298 224 299 
<< m1 >>
rect 223 298 224 299 
<< m2 >>
rect 223 298 224 299 
<< m1 >>
rect 239 298 240 299 
<< m1 >>
rect 247 298 248 299 
<< m1 >>
rect 253 298 254 299 
<< m1 >>
rect 255 298 256 299 
<< m1 >>
rect 265 298 266 299 
<< m1 >>
rect 271 298 272 299 
<< m2 >>
rect 271 298 272 299 
<< m1 >>
rect 276 298 277 299 
<< m1 >>
rect 278 298 279 299 
<< m1 >>
rect 323 298 324 299 
<< m2 >>
rect 323 298 324 299 
<< m2c >>
rect 323 298 324 299 
<< m1 >>
rect 323 298 324 299 
<< m2 >>
rect 323 298 324 299 
<< m2 >>
rect 324 298 325 299 
<< m1 >>
rect 325 298 326 299 
<< m2 >>
rect 325 298 326 299 
<< m2 >>
rect 326 298 327 299 
<< m1 >>
rect 327 298 328 299 
<< m2 >>
rect 327 298 328 299 
<< m2 >>
rect 328 298 329 299 
<< m1 >>
rect 331 298 332 299 
<< m1 >>
rect 334 298 335 299 
<< m1 >>
rect 10 299 11 300 
<< m1 >>
rect 13 299 14 300 
<< m1 >>
rect 28 299 29 300 
<< m1 >>
rect 37 299 38 300 
<< m2 >>
rect 38 299 39 300 
<< m1 >>
rect 46 299 47 300 
<< m1 >>
rect 55 299 56 300 
<< m2 >>
rect 55 299 56 300 
<< m1 >>
rect 57 299 58 300 
<< m1 >>
rect 60 299 61 300 
<< m1 >>
rect 62 299 63 300 
<< m1 >>
rect 64 299 65 300 
<< m1 >>
rect 73 299 74 300 
<< m2 >>
rect 81 299 82 300 
<< m1 >>
rect 82 299 83 300 
<< m1 >>
rect 103 299 104 300 
<< m1 >>
rect 109 299 110 300 
<< m1 >>
rect 142 299 143 300 
<< m1 >>
rect 145 299 146 300 
<< m1 >>
rect 169 299 170 300 
<< m2 >>
rect 171 299 172 300 
<< m1 >>
rect 172 299 173 300 
<< m1 >>
rect 181 299 182 300 
<< m1 >>
rect 193 299 194 300 
<< m2 >>
rect 203 299 204 300 
<< m1 >>
rect 208 299 209 300 
<< m1 >>
rect 217 299 218 300 
<< m1 >>
rect 219 299 220 300 
<< m1 >>
rect 221 299 222 300 
<< m1 >>
rect 223 299 224 300 
<< m1 >>
rect 239 299 240 300 
<< m1 >>
rect 247 299 248 300 
<< m1 >>
rect 253 299 254 300 
<< m1 >>
rect 255 299 256 300 
<< m1 >>
rect 265 299 266 300 
<< m1 >>
rect 271 299 272 300 
<< m2 >>
rect 271 299 272 300 
<< m1 >>
rect 276 299 277 300 
<< m1 >>
rect 278 299 279 300 
<< m1 >>
rect 325 299 326 300 
<< m1 >>
rect 327 299 328 300 
<< m2 >>
rect 328 299 329 300 
<< m1 >>
rect 331 299 332 300 
<< m1 >>
rect 334 299 335 300 
<< m1 >>
rect 10 300 11 301 
<< pdiffusion >>
rect 12 300 13 301 
<< m1 >>
rect 13 300 14 301 
<< pdiffusion >>
rect 13 300 14 301 
<< pdiffusion >>
rect 14 300 15 301 
<< pdiffusion >>
rect 15 300 16 301 
<< pdiffusion >>
rect 16 300 17 301 
<< pdiffusion >>
rect 17 300 18 301 
<< m1 >>
rect 28 300 29 301 
<< pdiffusion >>
rect 30 300 31 301 
<< pdiffusion >>
rect 31 300 32 301 
<< pdiffusion >>
rect 32 300 33 301 
<< pdiffusion >>
rect 33 300 34 301 
<< pdiffusion >>
rect 34 300 35 301 
<< pdiffusion >>
rect 35 300 36 301 
<< m1 >>
rect 37 300 38 301 
<< m2 >>
rect 38 300 39 301 
<< m1 >>
rect 46 300 47 301 
<< pdiffusion >>
rect 48 300 49 301 
<< pdiffusion >>
rect 49 300 50 301 
<< pdiffusion >>
rect 50 300 51 301 
<< pdiffusion >>
rect 51 300 52 301 
<< pdiffusion >>
rect 52 300 53 301 
<< pdiffusion >>
rect 53 300 54 301 
<< m1 >>
rect 55 300 56 301 
<< m2 >>
rect 55 300 56 301 
<< m1 >>
rect 57 300 58 301 
<< m1 >>
rect 60 300 61 301 
<< m1 >>
rect 62 300 63 301 
<< m1 >>
rect 64 300 65 301 
<< pdiffusion >>
rect 66 300 67 301 
<< pdiffusion >>
rect 67 300 68 301 
<< pdiffusion >>
rect 68 300 69 301 
<< pdiffusion >>
rect 69 300 70 301 
<< pdiffusion >>
rect 70 300 71 301 
<< pdiffusion >>
rect 71 300 72 301 
<< m1 >>
rect 73 300 74 301 
<< m2 >>
rect 81 300 82 301 
<< m1 >>
rect 82 300 83 301 
<< pdiffusion >>
rect 84 300 85 301 
<< pdiffusion >>
rect 85 300 86 301 
<< pdiffusion >>
rect 86 300 87 301 
<< pdiffusion >>
rect 87 300 88 301 
<< pdiffusion >>
rect 88 300 89 301 
<< pdiffusion >>
rect 89 300 90 301 
<< pdiffusion >>
rect 102 300 103 301 
<< m1 >>
rect 103 300 104 301 
<< pdiffusion >>
rect 103 300 104 301 
<< pdiffusion >>
rect 104 300 105 301 
<< pdiffusion >>
rect 105 300 106 301 
<< pdiffusion >>
rect 106 300 107 301 
<< pdiffusion >>
rect 107 300 108 301 
<< m1 >>
rect 109 300 110 301 
<< pdiffusion >>
rect 120 300 121 301 
<< pdiffusion >>
rect 121 300 122 301 
<< pdiffusion >>
rect 122 300 123 301 
<< pdiffusion >>
rect 123 300 124 301 
<< pdiffusion >>
rect 124 300 125 301 
<< pdiffusion >>
rect 125 300 126 301 
<< pdiffusion >>
rect 138 300 139 301 
<< pdiffusion >>
rect 139 300 140 301 
<< pdiffusion >>
rect 140 300 141 301 
<< pdiffusion >>
rect 141 300 142 301 
<< m1 >>
rect 142 300 143 301 
<< pdiffusion >>
rect 142 300 143 301 
<< pdiffusion >>
rect 143 300 144 301 
<< m1 >>
rect 145 300 146 301 
<< pdiffusion >>
rect 156 300 157 301 
<< pdiffusion >>
rect 157 300 158 301 
<< pdiffusion >>
rect 158 300 159 301 
<< pdiffusion >>
rect 159 300 160 301 
<< pdiffusion >>
rect 160 300 161 301 
<< pdiffusion >>
rect 161 300 162 301 
<< m1 >>
rect 169 300 170 301 
<< m2 >>
rect 171 300 172 301 
<< m1 >>
rect 172 300 173 301 
<< pdiffusion >>
rect 174 300 175 301 
<< pdiffusion >>
rect 175 300 176 301 
<< pdiffusion >>
rect 176 300 177 301 
<< pdiffusion >>
rect 177 300 178 301 
<< pdiffusion >>
rect 178 300 179 301 
<< pdiffusion >>
rect 179 300 180 301 
<< m1 >>
rect 181 300 182 301 
<< pdiffusion >>
rect 192 300 193 301 
<< m1 >>
rect 193 300 194 301 
<< pdiffusion >>
rect 193 300 194 301 
<< pdiffusion >>
rect 194 300 195 301 
<< pdiffusion >>
rect 195 300 196 301 
<< pdiffusion >>
rect 196 300 197 301 
<< pdiffusion >>
rect 197 300 198 301 
<< m1 >>
rect 203 300 204 301 
<< m2 >>
rect 203 300 204 301 
<< m2c >>
rect 203 300 204 301 
<< m1 >>
rect 203 300 204 301 
<< m2 >>
rect 203 300 204 301 
<< m1 >>
rect 208 300 209 301 
<< pdiffusion >>
rect 210 300 211 301 
<< pdiffusion >>
rect 211 300 212 301 
<< pdiffusion >>
rect 212 300 213 301 
<< pdiffusion >>
rect 213 300 214 301 
<< pdiffusion >>
rect 214 300 215 301 
<< pdiffusion >>
rect 215 300 216 301 
<< m1 >>
rect 217 300 218 301 
<< m1 >>
rect 219 300 220 301 
<< m1 >>
rect 221 300 222 301 
<< m1 >>
rect 223 300 224 301 
<< pdiffusion >>
rect 228 300 229 301 
<< pdiffusion >>
rect 229 300 230 301 
<< pdiffusion >>
rect 230 300 231 301 
<< pdiffusion >>
rect 231 300 232 301 
<< pdiffusion >>
rect 232 300 233 301 
<< pdiffusion >>
rect 233 300 234 301 
<< m1 >>
rect 239 300 240 301 
<< pdiffusion >>
rect 246 300 247 301 
<< m1 >>
rect 247 300 248 301 
<< pdiffusion >>
rect 247 300 248 301 
<< pdiffusion >>
rect 248 300 249 301 
<< pdiffusion >>
rect 249 300 250 301 
<< pdiffusion >>
rect 250 300 251 301 
<< pdiffusion >>
rect 251 300 252 301 
<< m1 >>
rect 253 300 254 301 
<< m1 >>
rect 255 300 256 301 
<< pdiffusion >>
rect 264 300 265 301 
<< m1 >>
rect 265 300 266 301 
<< pdiffusion >>
rect 265 300 266 301 
<< pdiffusion >>
rect 266 300 267 301 
<< pdiffusion >>
rect 267 300 268 301 
<< pdiffusion >>
rect 268 300 269 301 
<< pdiffusion >>
rect 269 300 270 301 
<< m1 >>
rect 271 300 272 301 
<< m2 >>
rect 271 300 272 301 
<< m1 >>
rect 276 300 277 301 
<< m1 >>
rect 278 300 279 301 
<< pdiffusion >>
rect 282 300 283 301 
<< pdiffusion >>
rect 283 300 284 301 
<< pdiffusion >>
rect 284 300 285 301 
<< pdiffusion >>
rect 285 300 286 301 
<< pdiffusion >>
rect 286 300 287 301 
<< pdiffusion >>
rect 287 300 288 301 
<< pdiffusion >>
rect 300 300 301 301 
<< pdiffusion >>
rect 301 300 302 301 
<< pdiffusion >>
rect 302 300 303 301 
<< pdiffusion >>
rect 303 300 304 301 
<< pdiffusion >>
rect 304 300 305 301 
<< pdiffusion >>
rect 305 300 306 301 
<< pdiffusion >>
rect 318 300 319 301 
<< pdiffusion >>
rect 319 300 320 301 
<< pdiffusion >>
rect 320 300 321 301 
<< pdiffusion >>
rect 321 300 322 301 
<< pdiffusion >>
rect 322 300 323 301 
<< pdiffusion >>
rect 323 300 324 301 
<< m1 >>
rect 325 300 326 301 
<< m1 >>
rect 327 300 328 301 
<< m2 >>
rect 328 300 329 301 
<< m1 >>
rect 331 300 332 301 
<< m1 >>
rect 334 300 335 301 
<< pdiffusion >>
rect 336 300 337 301 
<< pdiffusion >>
rect 337 300 338 301 
<< pdiffusion >>
rect 338 300 339 301 
<< pdiffusion >>
rect 339 300 340 301 
<< pdiffusion >>
rect 340 300 341 301 
<< pdiffusion >>
rect 341 300 342 301 
<< m1 >>
rect 10 301 11 302 
<< pdiffusion >>
rect 12 301 13 302 
<< pdiffusion >>
rect 13 301 14 302 
<< pdiffusion >>
rect 14 301 15 302 
<< pdiffusion >>
rect 15 301 16 302 
<< pdiffusion >>
rect 16 301 17 302 
<< pdiffusion >>
rect 17 301 18 302 
<< m1 >>
rect 28 301 29 302 
<< pdiffusion >>
rect 30 301 31 302 
<< pdiffusion >>
rect 31 301 32 302 
<< pdiffusion >>
rect 32 301 33 302 
<< pdiffusion >>
rect 33 301 34 302 
<< pdiffusion >>
rect 34 301 35 302 
<< pdiffusion >>
rect 35 301 36 302 
<< m1 >>
rect 37 301 38 302 
<< m2 >>
rect 38 301 39 302 
<< m1 >>
rect 46 301 47 302 
<< pdiffusion >>
rect 48 301 49 302 
<< pdiffusion >>
rect 49 301 50 302 
<< pdiffusion >>
rect 50 301 51 302 
<< pdiffusion >>
rect 51 301 52 302 
<< pdiffusion >>
rect 52 301 53 302 
<< pdiffusion >>
rect 53 301 54 302 
<< m1 >>
rect 55 301 56 302 
<< m2 >>
rect 55 301 56 302 
<< m1 >>
rect 57 301 58 302 
<< m1 >>
rect 60 301 61 302 
<< m1 >>
rect 62 301 63 302 
<< m1 >>
rect 64 301 65 302 
<< pdiffusion >>
rect 66 301 67 302 
<< pdiffusion >>
rect 67 301 68 302 
<< pdiffusion >>
rect 68 301 69 302 
<< pdiffusion >>
rect 69 301 70 302 
<< pdiffusion >>
rect 70 301 71 302 
<< pdiffusion >>
rect 71 301 72 302 
<< m1 >>
rect 73 301 74 302 
<< m2 >>
rect 81 301 82 302 
<< m1 >>
rect 82 301 83 302 
<< pdiffusion >>
rect 84 301 85 302 
<< pdiffusion >>
rect 85 301 86 302 
<< pdiffusion >>
rect 86 301 87 302 
<< pdiffusion >>
rect 87 301 88 302 
<< pdiffusion >>
rect 88 301 89 302 
<< pdiffusion >>
rect 89 301 90 302 
<< pdiffusion >>
rect 102 301 103 302 
<< pdiffusion >>
rect 103 301 104 302 
<< pdiffusion >>
rect 104 301 105 302 
<< pdiffusion >>
rect 105 301 106 302 
<< pdiffusion >>
rect 106 301 107 302 
<< pdiffusion >>
rect 107 301 108 302 
<< m1 >>
rect 109 301 110 302 
<< pdiffusion >>
rect 120 301 121 302 
<< pdiffusion >>
rect 121 301 122 302 
<< pdiffusion >>
rect 122 301 123 302 
<< pdiffusion >>
rect 123 301 124 302 
<< pdiffusion >>
rect 124 301 125 302 
<< pdiffusion >>
rect 125 301 126 302 
<< pdiffusion >>
rect 138 301 139 302 
<< pdiffusion >>
rect 139 301 140 302 
<< pdiffusion >>
rect 140 301 141 302 
<< pdiffusion >>
rect 141 301 142 302 
<< pdiffusion >>
rect 142 301 143 302 
<< pdiffusion >>
rect 143 301 144 302 
<< m1 >>
rect 145 301 146 302 
<< pdiffusion >>
rect 156 301 157 302 
<< pdiffusion >>
rect 157 301 158 302 
<< pdiffusion >>
rect 158 301 159 302 
<< pdiffusion >>
rect 159 301 160 302 
<< pdiffusion >>
rect 160 301 161 302 
<< pdiffusion >>
rect 161 301 162 302 
<< m1 >>
rect 169 301 170 302 
<< m2 >>
rect 171 301 172 302 
<< m1 >>
rect 172 301 173 302 
<< pdiffusion >>
rect 174 301 175 302 
<< pdiffusion >>
rect 175 301 176 302 
<< pdiffusion >>
rect 176 301 177 302 
<< pdiffusion >>
rect 177 301 178 302 
<< pdiffusion >>
rect 178 301 179 302 
<< pdiffusion >>
rect 179 301 180 302 
<< m1 >>
rect 181 301 182 302 
<< pdiffusion >>
rect 192 301 193 302 
<< pdiffusion >>
rect 193 301 194 302 
<< pdiffusion >>
rect 194 301 195 302 
<< pdiffusion >>
rect 195 301 196 302 
<< pdiffusion >>
rect 196 301 197 302 
<< pdiffusion >>
rect 197 301 198 302 
<< m1 >>
rect 203 301 204 302 
<< m1 >>
rect 208 301 209 302 
<< pdiffusion >>
rect 210 301 211 302 
<< pdiffusion >>
rect 211 301 212 302 
<< pdiffusion >>
rect 212 301 213 302 
<< pdiffusion >>
rect 213 301 214 302 
<< pdiffusion >>
rect 214 301 215 302 
<< pdiffusion >>
rect 215 301 216 302 
<< m1 >>
rect 217 301 218 302 
<< m1 >>
rect 219 301 220 302 
<< m1 >>
rect 221 301 222 302 
<< m1 >>
rect 223 301 224 302 
<< pdiffusion >>
rect 228 301 229 302 
<< pdiffusion >>
rect 229 301 230 302 
<< pdiffusion >>
rect 230 301 231 302 
<< pdiffusion >>
rect 231 301 232 302 
<< pdiffusion >>
rect 232 301 233 302 
<< pdiffusion >>
rect 233 301 234 302 
<< m1 >>
rect 239 301 240 302 
<< pdiffusion >>
rect 246 301 247 302 
<< pdiffusion >>
rect 247 301 248 302 
<< pdiffusion >>
rect 248 301 249 302 
<< pdiffusion >>
rect 249 301 250 302 
<< pdiffusion >>
rect 250 301 251 302 
<< pdiffusion >>
rect 251 301 252 302 
<< m1 >>
rect 253 301 254 302 
<< m1 >>
rect 255 301 256 302 
<< pdiffusion >>
rect 264 301 265 302 
<< pdiffusion >>
rect 265 301 266 302 
<< pdiffusion >>
rect 266 301 267 302 
<< pdiffusion >>
rect 267 301 268 302 
<< pdiffusion >>
rect 268 301 269 302 
<< pdiffusion >>
rect 269 301 270 302 
<< m1 >>
rect 271 301 272 302 
<< m2 >>
rect 271 301 272 302 
<< m1 >>
rect 276 301 277 302 
<< m1 >>
rect 278 301 279 302 
<< pdiffusion >>
rect 282 301 283 302 
<< pdiffusion >>
rect 283 301 284 302 
<< pdiffusion >>
rect 284 301 285 302 
<< pdiffusion >>
rect 285 301 286 302 
<< pdiffusion >>
rect 286 301 287 302 
<< pdiffusion >>
rect 287 301 288 302 
<< pdiffusion >>
rect 300 301 301 302 
<< pdiffusion >>
rect 301 301 302 302 
<< pdiffusion >>
rect 302 301 303 302 
<< pdiffusion >>
rect 303 301 304 302 
<< pdiffusion >>
rect 304 301 305 302 
<< pdiffusion >>
rect 305 301 306 302 
<< pdiffusion >>
rect 318 301 319 302 
<< pdiffusion >>
rect 319 301 320 302 
<< pdiffusion >>
rect 320 301 321 302 
<< pdiffusion >>
rect 321 301 322 302 
<< pdiffusion >>
rect 322 301 323 302 
<< pdiffusion >>
rect 323 301 324 302 
<< m1 >>
rect 325 301 326 302 
<< m1 >>
rect 327 301 328 302 
<< m2 >>
rect 328 301 329 302 
<< m1 >>
rect 331 301 332 302 
<< m1 >>
rect 334 301 335 302 
<< pdiffusion >>
rect 336 301 337 302 
<< pdiffusion >>
rect 337 301 338 302 
<< pdiffusion >>
rect 338 301 339 302 
<< pdiffusion >>
rect 339 301 340 302 
<< pdiffusion >>
rect 340 301 341 302 
<< pdiffusion >>
rect 341 301 342 302 
<< m1 >>
rect 10 302 11 303 
<< pdiffusion >>
rect 12 302 13 303 
<< pdiffusion >>
rect 13 302 14 303 
<< pdiffusion >>
rect 14 302 15 303 
<< pdiffusion >>
rect 15 302 16 303 
<< pdiffusion >>
rect 16 302 17 303 
<< pdiffusion >>
rect 17 302 18 303 
<< m1 >>
rect 28 302 29 303 
<< pdiffusion >>
rect 30 302 31 303 
<< pdiffusion >>
rect 31 302 32 303 
<< pdiffusion >>
rect 32 302 33 303 
<< pdiffusion >>
rect 33 302 34 303 
<< pdiffusion >>
rect 34 302 35 303 
<< pdiffusion >>
rect 35 302 36 303 
<< m1 >>
rect 37 302 38 303 
<< m2 >>
rect 38 302 39 303 
<< m1 >>
rect 46 302 47 303 
<< pdiffusion >>
rect 48 302 49 303 
<< pdiffusion >>
rect 49 302 50 303 
<< pdiffusion >>
rect 50 302 51 303 
<< pdiffusion >>
rect 51 302 52 303 
<< pdiffusion >>
rect 52 302 53 303 
<< pdiffusion >>
rect 53 302 54 303 
<< m1 >>
rect 55 302 56 303 
<< m2 >>
rect 55 302 56 303 
<< m1 >>
rect 57 302 58 303 
<< m1 >>
rect 60 302 61 303 
<< m1 >>
rect 62 302 63 303 
<< m1 >>
rect 64 302 65 303 
<< pdiffusion >>
rect 66 302 67 303 
<< pdiffusion >>
rect 67 302 68 303 
<< pdiffusion >>
rect 68 302 69 303 
<< pdiffusion >>
rect 69 302 70 303 
<< pdiffusion >>
rect 70 302 71 303 
<< pdiffusion >>
rect 71 302 72 303 
<< m1 >>
rect 73 302 74 303 
<< m2 >>
rect 81 302 82 303 
<< m1 >>
rect 82 302 83 303 
<< pdiffusion >>
rect 84 302 85 303 
<< pdiffusion >>
rect 85 302 86 303 
<< pdiffusion >>
rect 86 302 87 303 
<< pdiffusion >>
rect 87 302 88 303 
<< pdiffusion >>
rect 88 302 89 303 
<< pdiffusion >>
rect 89 302 90 303 
<< pdiffusion >>
rect 102 302 103 303 
<< pdiffusion >>
rect 103 302 104 303 
<< pdiffusion >>
rect 104 302 105 303 
<< pdiffusion >>
rect 105 302 106 303 
<< pdiffusion >>
rect 106 302 107 303 
<< pdiffusion >>
rect 107 302 108 303 
<< m1 >>
rect 109 302 110 303 
<< pdiffusion >>
rect 120 302 121 303 
<< pdiffusion >>
rect 121 302 122 303 
<< pdiffusion >>
rect 122 302 123 303 
<< pdiffusion >>
rect 123 302 124 303 
<< pdiffusion >>
rect 124 302 125 303 
<< pdiffusion >>
rect 125 302 126 303 
<< pdiffusion >>
rect 138 302 139 303 
<< pdiffusion >>
rect 139 302 140 303 
<< pdiffusion >>
rect 140 302 141 303 
<< pdiffusion >>
rect 141 302 142 303 
<< pdiffusion >>
rect 142 302 143 303 
<< pdiffusion >>
rect 143 302 144 303 
<< m1 >>
rect 145 302 146 303 
<< pdiffusion >>
rect 156 302 157 303 
<< pdiffusion >>
rect 157 302 158 303 
<< pdiffusion >>
rect 158 302 159 303 
<< pdiffusion >>
rect 159 302 160 303 
<< pdiffusion >>
rect 160 302 161 303 
<< pdiffusion >>
rect 161 302 162 303 
<< m1 >>
rect 169 302 170 303 
<< m2 >>
rect 171 302 172 303 
<< m1 >>
rect 172 302 173 303 
<< pdiffusion >>
rect 174 302 175 303 
<< pdiffusion >>
rect 175 302 176 303 
<< pdiffusion >>
rect 176 302 177 303 
<< pdiffusion >>
rect 177 302 178 303 
<< pdiffusion >>
rect 178 302 179 303 
<< pdiffusion >>
rect 179 302 180 303 
<< m1 >>
rect 181 302 182 303 
<< pdiffusion >>
rect 192 302 193 303 
<< pdiffusion >>
rect 193 302 194 303 
<< pdiffusion >>
rect 194 302 195 303 
<< pdiffusion >>
rect 195 302 196 303 
<< pdiffusion >>
rect 196 302 197 303 
<< pdiffusion >>
rect 197 302 198 303 
<< m1 >>
rect 203 302 204 303 
<< m1 >>
rect 208 302 209 303 
<< pdiffusion >>
rect 210 302 211 303 
<< pdiffusion >>
rect 211 302 212 303 
<< pdiffusion >>
rect 212 302 213 303 
<< pdiffusion >>
rect 213 302 214 303 
<< pdiffusion >>
rect 214 302 215 303 
<< pdiffusion >>
rect 215 302 216 303 
<< m1 >>
rect 217 302 218 303 
<< m1 >>
rect 219 302 220 303 
<< m1 >>
rect 221 302 222 303 
<< m1 >>
rect 223 302 224 303 
<< pdiffusion >>
rect 228 302 229 303 
<< pdiffusion >>
rect 229 302 230 303 
<< pdiffusion >>
rect 230 302 231 303 
<< pdiffusion >>
rect 231 302 232 303 
<< pdiffusion >>
rect 232 302 233 303 
<< pdiffusion >>
rect 233 302 234 303 
<< m1 >>
rect 239 302 240 303 
<< pdiffusion >>
rect 246 302 247 303 
<< pdiffusion >>
rect 247 302 248 303 
<< pdiffusion >>
rect 248 302 249 303 
<< pdiffusion >>
rect 249 302 250 303 
<< pdiffusion >>
rect 250 302 251 303 
<< pdiffusion >>
rect 251 302 252 303 
<< m1 >>
rect 253 302 254 303 
<< m1 >>
rect 255 302 256 303 
<< pdiffusion >>
rect 264 302 265 303 
<< pdiffusion >>
rect 265 302 266 303 
<< pdiffusion >>
rect 266 302 267 303 
<< pdiffusion >>
rect 267 302 268 303 
<< pdiffusion >>
rect 268 302 269 303 
<< pdiffusion >>
rect 269 302 270 303 
<< m1 >>
rect 271 302 272 303 
<< m2 >>
rect 271 302 272 303 
<< m1 >>
rect 276 302 277 303 
<< m1 >>
rect 278 302 279 303 
<< pdiffusion >>
rect 282 302 283 303 
<< pdiffusion >>
rect 283 302 284 303 
<< pdiffusion >>
rect 284 302 285 303 
<< pdiffusion >>
rect 285 302 286 303 
<< pdiffusion >>
rect 286 302 287 303 
<< pdiffusion >>
rect 287 302 288 303 
<< pdiffusion >>
rect 300 302 301 303 
<< pdiffusion >>
rect 301 302 302 303 
<< pdiffusion >>
rect 302 302 303 303 
<< pdiffusion >>
rect 303 302 304 303 
<< pdiffusion >>
rect 304 302 305 303 
<< pdiffusion >>
rect 305 302 306 303 
<< pdiffusion >>
rect 318 302 319 303 
<< pdiffusion >>
rect 319 302 320 303 
<< pdiffusion >>
rect 320 302 321 303 
<< pdiffusion >>
rect 321 302 322 303 
<< pdiffusion >>
rect 322 302 323 303 
<< pdiffusion >>
rect 323 302 324 303 
<< m1 >>
rect 325 302 326 303 
<< m1 >>
rect 327 302 328 303 
<< m2 >>
rect 328 302 329 303 
<< m1 >>
rect 331 302 332 303 
<< m1 >>
rect 334 302 335 303 
<< pdiffusion >>
rect 336 302 337 303 
<< pdiffusion >>
rect 337 302 338 303 
<< pdiffusion >>
rect 338 302 339 303 
<< pdiffusion >>
rect 339 302 340 303 
<< pdiffusion >>
rect 340 302 341 303 
<< pdiffusion >>
rect 341 302 342 303 
<< m1 >>
rect 10 303 11 304 
<< pdiffusion >>
rect 12 303 13 304 
<< pdiffusion >>
rect 13 303 14 304 
<< pdiffusion >>
rect 14 303 15 304 
<< pdiffusion >>
rect 15 303 16 304 
<< pdiffusion >>
rect 16 303 17 304 
<< pdiffusion >>
rect 17 303 18 304 
<< m1 >>
rect 28 303 29 304 
<< pdiffusion >>
rect 30 303 31 304 
<< pdiffusion >>
rect 31 303 32 304 
<< pdiffusion >>
rect 32 303 33 304 
<< pdiffusion >>
rect 33 303 34 304 
<< pdiffusion >>
rect 34 303 35 304 
<< pdiffusion >>
rect 35 303 36 304 
<< m1 >>
rect 37 303 38 304 
<< m2 >>
rect 38 303 39 304 
<< m1 >>
rect 46 303 47 304 
<< pdiffusion >>
rect 48 303 49 304 
<< pdiffusion >>
rect 49 303 50 304 
<< pdiffusion >>
rect 50 303 51 304 
<< pdiffusion >>
rect 51 303 52 304 
<< pdiffusion >>
rect 52 303 53 304 
<< pdiffusion >>
rect 53 303 54 304 
<< m1 >>
rect 55 303 56 304 
<< m2 >>
rect 55 303 56 304 
<< m1 >>
rect 57 303 58 304 
<< m1 >>
rect 60 303 61 304 
<< m1 >>
rect 62 303 63 304 
<< m1 >>
rect 64 303 65 304 
<< pdiffusion >>
rect 66 303 67 304 
<< pdiffusion >>
rect 67 303 68 304 
<< pdiffusion >>
rect 68 303 69 304 
<< pdiffusion >>
rect 69 303 70 304 
<< pdiffusion >>
rect 70 303 71 304 
<< pdiffusion >>
rect 71 303 72 304 
<< m1 >>
rect 73 303 74 304 
<< m2 >>
rect 81 303 82 304 
<< m1 >>
rect 82 303 83 304 
<< pdiffusion >>
rect 84 303 85 304 
<< pdiffusion >>
rect 85 303 86 304 
<< pdiffusion >>
rect 86 303 87 304 
<< pdiffusion >>
rect 87 303 88 304 
<< pdiffusion >>
rect 88 303 89 304 
<< pdiffusion >>
rect 89 303 90 304 
<< pdiffusion >>
rect 102 303 103 304 
<< pdiffusion >>
rect 103 303 104 304 
<< pdiffusion >>
rect 104 303 105 304 
<< pdiffusion >>
rect 105 303 106 304 
<< pdiffusion >>
rect 106 303 107 304 
<< pdiffusion >>
rect 107 303 108 304 
<< m1 >>
rect 109 303 110 304 
<< pdiffusion >>
rect 120 303 121 304 
<< pdiffusion >>
rect 121 303 122 304 
<< pdiffusion >>
rect 122 303 123 304 
<< pdiffusion >>
rect 123 303 124 304 
<< pdiffusion >>
rect 124 303 125 304 
<< pdiffusion >>
rect 125 303 126 304 
<< pdiffusion >>
rect 138 303 139 304 
<< pdiffusion >>
rect 139 303 140 304 
<< pdiffusion >>
rect 140 303 141 304 
<< pdiffusion >>
rect 141 303 142 304 
<< pdiffusion >>
rect 142 303 143 304 
<< pdiffusion >>
rect 143 303 144 304 
<< m1 >>
rect 145 303 146 304 
<< pdiffusion >>
rect 156 303 157 304 
<< pdiffusion >>
rect 157 303 158 304 
<< pdiffusion >>
rect 158 303 159 304 
<< pdiffusion >>
rect 159 303 160 304 
<< pdiffusion >>
rect 160 303 161 304 
<< pdiffusion >>
rect 161 303 162 304 
<< m1 >>
rect 169 303 170 304 
<< m2 >>
rect 171 303 172 304 
<< m1 >>
rect 172 303 173 304 
<< pdiffusion >>
rect 174 303 175 304 
<< pdiffusion >>
rect 175 303 176 304 
<< pdiffusion >>
rect 176 303 177 304 
<< pdiffusion >>
rect 177 303 178 304 
<< pdiffusion >>
rect 178 303 179 304 
<< pdiffusion >>
rect 179 303 180 304 
<< m1 >>
rect 181 303 182 304 
<< pdiffusion >>
rect 192 303 193 304 
<< pdiffusion >>
rect 193 303 194 304 
<< pdiffusion >>
rect 194 303 195 304 
<< pdiffusion >>
rect 195 303 196 304 
<< pdiffusion >>
rect 196 303 197 304 
<< pdiffusion >>
rect 197 303 198 304 
<< m1 >>
rect 203 303 204 304 
<< m1 >>
rect 208 303 209 304 
<< pdiffusion >>
rect 210 303 211 304 
<< pdiffusion >>
rect 211 303 212 304 
<< pdiffusion >>
rect 212 303 213 304 
<< pdiffusion >>
rect 213 303 214 304 
<< pdiffusion >>
rect 214 303 215 304 
<< pdiffusion >>
rect 215 303 216 304 
<< m1 >>
rect 217 303 218 304 
<< m1 >>
rect 219 303 220 304 
<< m1 >>
rect 221 303 222 304 
<< m1 >>
rect 223 303 224 304 
<< pdiffusion >>
rect 228 303 229 304 
<< pdiffusion >>
rect 229 303 230 304 
<< pdiffusion >>
rect 230 303 231 304 
<< pdiffusion >>
rect 231 303 232 304 
<< pdiffusion >>
rect 232 303 233 304 
<< pdiffusion >>
rect 233 303 234 304 
<< m1 >>
rect 239 303 240 304 
<< pdiffusion >>
rect 246 303 247 304 
<< pdiffusion >>
rect 247 303 248 304 
<< pdiffusion >>
rect 248 303 249 304 
<< pdiffusion >>
rect 249 303 250 304 
<< pdiffusion >>
rect 250 303 251 304 
<< pdiffusion >>
rect 251 303 252 304 
<< m1 >>
rect 253 303 254 304 
<< m1 >>
rect 255 303 256 304 
<< pdiffusion >>
rect 264 303 265 304 
<< pdiffusion >>
rect 265 303 266 304 
<< pdiffusion >>
rect 266 303 267 304 
<< pdiffusion >>
rect 267 303 268 304 
<< pdiffusion >>
rect 268 303 269 304 
<< pdiffusion >>
rect 269 303 270 304 
<< m1 >>
rect 271 303 272 304 
<< m2 >>
rect 271 303 272 304 
<< m1 >>
rect 276 303 277 304 
<< m1 >>
rect 278 303 279 304 
<< pdiffusion >>
rect 282 303 283 304 
<< pdiffusion >>
rect 283 303 284 304 
<< pdiffusion >>
rect 284 303 285 304 
<< pdiffusion >>
rect 285 303 286 304 
<< pdiffusion >>
rect 286 303 287 304 
<< pdiffusion >>
rect 287 303 288 304 
<< pdiffusion >>
rect 300 303 301 304 
<< pdiffusion >>
rect 301 303 302 304 
<< pdiffusion >>
rect 302 303 303 304 
<< pdiffusion >>
rect 303 303 304 304 
<< pdiffusion >>
rect 304 303 305 304 
<< pdiffusion >>
rect 305 303 306 304 
<< pdiffusion >>
rect 318 303 319 304 
<< pdiffusion >>
rect 319 303 320 304 
<< pdiffusion >>
rect 320 303 321 304 
<< pdiffusion >>
rect 321 303 322 304 
<< pdiffusion >>
rect 322 303 323 304 
<< pdiffusion >>
rect 323 303 324 304 
<< m1 >>
rect 325 303 326 304 
<< m1 >>
rect 327 303 328 304 
<< m2 >>
rect 328 303 329 304 
<< m1 >>
rect 331 303 332 304 
<< m1 >>
rect 334 303 335 304 
<< pdiffusion >>
rect 336 303 337 304 
<< pdiffusion >>
rect 337 303 338 304 
<< pdiffusion >>
rect 338 303 339 304 
<< pdiffusion >>
rect 339 303 340 304 
<< pdiffusion >>
rect 340 303 341 304 
<< pdiffusion >>
rect 341 303 342 304 
<< m1 >>
rect 10 304 11 305 
<< pdiffusion >>
rect 12 304 13 305 
<< pdiffusion >>
rect 13 304 14 305 
<< pdiffusion >>
rect 14 304 15 305 
<< pdiffusion >>
rect 15 304 16 305 
<< pdiffusion >>
rect 16 304 17 305 
<< pdiffusion >>
rect 17 304 18 305 
<< m1 >>
rect 28 304 29 305 
<< pdiffusion >>
rect 30 304 31 305 
<< pdiffusion >>
rect 31 304 32 305 
<< pdiffusion >>
rect 32 304 33 305 
<< pdiffusion >>
rect 33 304 34 305 
<< pdiffusion >>
rect 34 304 35 305 
<< pdiffusion >>
rect 35 304 36 305 
<< m1 >>
rect 37 304 38 305 
<< m2 >>
rect 38 304 39 305 
<< m1 >>
rect 46 304 47 305 
<< pdiffusion >>
rect 48 304 49 305 
<< pdiffusion >>
rect 49 304 50 305 
<< pdiffusion >>
rect 50 304 51 305 
<< pdiffusion >>
rect 51 304 52 305 
<< pdiffusion >>
rect 52 304 53 305 
<< pdiffusion >>
rect 53 304 54 305 
<< m1 >>
rect 55 304 56 305 
<< m2 >>
rect 55 304 56 305 
<< m1 >>
rect 57 304 58 305 
<< m1 >>
rect 60 304 61 305 
<< m1 >>
rect 62 304 63 305 
<< m1 >>
rect 64 304 65 305 
<< pdiffusion >>
rect 66 304 67 305 
<< pdiffusion >>
rect 67 304 68 305 
<< pdiffusion >>
rect 68 304 69 305 
<< pdiffusion >>
rect 69 304 70 305 
<< pdiffusion >>
rect 70 304 71 305 
<< pdiffusion >>
rect 71 304 72 305 
<< m1 >>
rect 73 304 74 305 
<< m2 >>
rect 81 304 82 305 
<< m1 >>
rect 82 304 83 305 
<< pdiffusion >>
rect 84 304 85 305 
<< pdiffusion >>
rect 85 304 86 305 
<< pdiffusion >>
rect 86 304 87 305 
<< pdiffusion >>
rect 87 304 88 305 
<< pdiffusion >>
rect 88 304 89 305 
<< pdiffusion >>
rect 89 304 90 305 
<< pdiffusion >>
rect 102 304 103 305 
<< pdiffusion >>
rect 103 304 104 305 
<< pdiffusion >>
rect 104 304 105 305 
<< pdiffusion >>
rect 105 304 106 305 
<< pdiffusion >>
rect 106 304 107 305 
<< pdiffusion >>
rect 107 304 108 305 
<< m1 >>
rect 109 304 110 305 
<< pdiffusion >>
rect 120 304 121 305 
<< pdiffusion >>
rect 121 304 122 305 
<< pdiffusion >>
rect 122 304 123 305 
<< pdiffusion >>
rect 123 304 124 305 
<< pdiffusion >>
rect 124 304 125 305 
<< pdiffusion >>
rect 125 304 126 305 
<< pdiffusion >>
rect 138 304 139 305 
<< pdiffusion >>
rect 139 304 140 305 
<< pdiffusion >>
rect 140 304 141 305 
<< pdiffusion >>
rect 141 304 142 305 
<< pdiffusion >>
rect 142 304 143 305 
<< pdiffusion >>
rect 143 304 144 305 
<< m1 >>
rect 145 304 146 305 
<< pdiffusion >>
rect 156 304 157 305 
<< pdiffusion >>
rect 157 304 158 305 
<< pdiffusion >>
rect 158 304 159 305 
<< pdiffusion >>
rect 159 304 160 305 
<< pdiffusion >>
rect 160 304 161 305 
<< pdiffusion >>
rect 161 304 162 305 
<< m1 >>
rect 169 304 170 305 
<< m2 >>
rect 171 304 172 305 
<< m1 >>
rect 172 304 173 305 
<< pdiffusion >>
rect 174 304 175 305 
<< pdiffusion >>
rect 175 304 176 305 
<< pdiffusion >>
rect 176 304 177 305 
<< pdiffusion >>
rect 177 304 178 305 
<< pdiffusion >>
rect 178 304 179 305 
<< pdiffusion >>
rect 179 304 180 305 
<< m1 >>
rect 181 304 182 305 
<< pdiffusion >>
rect 192 304 193 305 
<< pdiffusion >>
rect 193 304 194 305 
<< pdiffusion >>
rect 194 304 195 305 
<< pdiffusion >>
rect 195 304 196 305 
<< pdiffusion >>
rect 196 304 197 305 
<< pdiffusion >>
rect 197 304 198 305 
<< m1 >>
rect 203 304 204 305 
<< m1 >>
rect 208 304 209 305 
<< pdiffusion >>
rect 210 304 211 305 
<< pdiffusion >>
rect 211 304 212 305 
<< pdiffusion >>
rect 212 304 213 305 
<< pdiffusion >>
rect 213 304 214 305 
<< pdiffusion >>
rect 214 304 215 305 
<< pdiffusion >>
rect 215 304 216 305 
<< m1 >>
rect 217 304 218 305 
<< m1 >>
rect 219 304 220 305 
<< m1 >>
rect 221 304 222 305 
<< m1 >>
rect 223 304 224 305 
<< pdiffusion >>
rect 228 304 229 305 
<< pdiffusion >>
rect 229 304 230 305 
<< pdiffusion >>
rect 230 304 231 305 
<< pdiffusion >>
rect 231 304 232 305 
<< pdiffusion >>
rect 232 304 233 305 
<< pdiffusion >>
rect 233 304 234 305 
<< m1 >>
rect 239 304 240 305 
<< pdiffusion >>
rect 246 304 247 305 
<< pdiffusion >>
rect 247 304 248 305 
<< pdiffusion >>
rect 248 304 249 305 
<< pdiffusion >>
rect 249 304 250 305 
<< pdiffusion >>
rect 250 304 251 305 
<< pdiffusion >>
rect 251 304 252 305 
<< m1 >>
rect 253 304 254 305 
<< m1 >>
rect 255 304 256 305 
<< pdiffusion >>
rect 264 304 265 305 
<< pdiffusion >>
rect 265 304 266 305 
<< pdiffusion >>
rect 266 304 267 305 
<< pdiffusion >>
rect 267 304 268 305 
<< pdiffusion >>
rect 268 304 269 305 
<< pdiffusion >>
rect 269 304 270 305 
<< m1 >>
rect 271 304 272 305 
<< m2 >>
rect 271 304 272 305 
<< m1 >>
rect 276 304 277 305 
<< m1 >>
rect 278 304 279 305 
<< pdiffusion >>
rect 282 304 283 305 
<< pdiffusion >>
rect 283 304 284 305 
<< pdiffusion >>
rect 284 304 285 305 
<< pdiffusion >>
rect 285 304 286 305 
<< pdiffusion >>
rect 286 304 287 305 
<< pdiffusion >>
rect 287 304 288 305 
<< pdiffusion >>
rect 300 304 301 305 
<< pdiffusion >>
rect 301 304 302 305 
<< pdiffusion >>
rect 302 304 303 305 
<< pdiffusion >>
rect 303 304 304 305 
<< pdiffusion >>
rect 304 304 305 305 
<< pdiffusion >>
rect 305 304 306 305 
<< pdiffusion >>
rect 318 304 319 305 
<< pdiffusion >>
rect 319 304 320 305 
<< pdiffusion >>
rect 320 304 321 305 
<< pdiffusion >>
rect 321 304 322 305 
<< pdiffusion >>
rect 322 304 323 305 
<< pdiffusion >>
rect 323 304 324 305 
<< m1 >>
rect 325 304 326 305 
<< m1 >>
rect 327 304 328 305 
<< m2 >>
rect 328 304 329 305 
<< m1 >>
rect 331 304 332 305 
<< m1 >>
rect 334 304 335 305 
<< pdiffusion >>
rect 336 304 337 305 
<< pdiffusion >>
rect 337 304 338 305 
<< pdiffusion >>
rect 338 304 339 305 
<< pdiffusion >>
rect 339 304 340 305 
<< pdiffusion >>
rect 340 304 341 305 
<< pdiffusion >>
rect 341 304 342 305 
<< m1 >>
rect 10 305 11 306 
<< pdiffusion >>
rect 12 305 13 306 
<< pdiffusion >>
rect 13 305 14 306 
<< pdiffusion >>
rect 14 305 15 306 
<< pdiffusion >>
rect 15 305 16 306 
<< pdiffusion >>
rect 16 305 17 306 
<< pdiffusion >>
rect 17 305 18 306 
<< m1 >>
rect 28 305 29 306 
<< pdiffusion >>
rect 30 305 31 306 
<< pdiffusion >>
rect 31 305 32 306 
<< pdiffusion >>
rect 32 305 33 306 
<< pdiffusion >>
rect 33 305 34 306 
<< pdiffusion >>
rect 34 305 35 306 
<< pdiffusion >>
rect 35 305 36 306 
<< m1 >>
rect 37 305 38 306 
<< m2 >>
rect 38 305 39 306 
<< m1 >>
rect 46 305 47 306 
<< pdiffusion >>
rect 48 305 49 306 
<< m1 >>
rect 49 305 50 306 
<< pdiffusion >>
rect 49 305 50 306 
<< pdiffusion >>
rect 50 305 51 306 
<< pdiffusion >>
rect 51 305 52 306 
<< pdiffusion >>
rect 52 305 53 306 
<< pdiffusion >>
rect 53 305 54 306 
<< m1 >>
rect 55 305 56 306 
<< m2 >>
rect 55 305 56 306 
<< m1 >>
rect 57 305 58 306 
<< m1 >>
rect 60 305 61 306 
<< m1 >>
rect 62 305 63 306 
<< m1 >>
rect 64 305 65 306 
<< pdiffusion >>
rect 66 305 67 306 
<< pdiffusion >>
rect 67 305 68 306 
<< pdiffusion >>
rect 68 305 69 306 
<< pdiffusion >>
rect 69 305 70 306 
<< pdiffusion >>
rect 70 305 71 306 
<< pdiffusion >>
rect 71 305 72 306 
<< m1 >>
rect 73 305 74 306 
<< m2 >>
rect 81 305 82 306 
<< m1 >>
rect 82 305 83 306 
<< pdiffusion >>
rect 84 305 85 306 
<< pdiffusion >>
rect 85 305 86 306 
<< pdiffusion >>
rect 86 305 87 306 
<< pdiffusion >>
rect 87 305 88 306 
<< pdiffusion >>
rect 88 305 89 306 
<< pdiffusion >>
rect 89 305 90 306 
<< pdiffusion >>
rect 102 305 103 306 
<< pdiffusion >>
rect 103 305 104 306 
<< pdiffusion >>
rect 104 305 105 306 
<< pdiffusion >>
rect 105 305 106 306 
<< pdiffusion >>
rect 106 305 107 306 
<< pdiffusion >>
rect 107 305 108 306 
<< m1 >>
rect 109 305 110 306 
<< pdiffusion >>
rect 120 305 121 306 
<< pdiffusion >>
rect 121 305 122 306 
<< pdiffusion >>
rect 122 305 123 306 
<< pdiffusion >>
rect 123 305 124 306 
<< pdiffusion >>
rect 124 305 125 306 
<< pdiffusion >>
rect 125 305 126 306 
<< pdiffusion >>
rect 138 305 139 306 
<< pdiffusion >>
rect 139 305 140 306 
<< pdiffusion >>
rect 140 305 141 306 
<< pdiffusion >>
rect 141 305 142 306 
<< pdiffusion >>
rect 142 305 143 306 
<< pdiffusion >>
rect 143 305 144 306 
<< m1 >>
rect 145 305 146 306 
<< pdiffusion >>
rect 156 305 157 306 
<< pdiffusion >>
rect 157 305 158 306 
<< pdiffusion >>
rect 158 305 159 306 
<< pdiffusion >>
rect 159 305 160 306 
<< pdiffusion >>
rect 160 305 161 306 
<< pdiffusion >>
rect 161 305 162 306 
<< m1 >>
rect 169 305 170 306 
<< m2 >>
rect 171 305 172 306 
<< m1 >>
rect 172 305 173 306 
<< pdiffusion >>
rect 174 305 175 306 
<< pdiffusion >>
rect 175 305 176 306 
<< pdiffusion >>
rect 176 305 177 306 
<< pdiffusion >>
rect 177 305 178 306 
<< pdiffusion >>
rect 178 305 179 306 
<< pdiffusion >>
rect 179 305 180 306 
<< m1 >>
rect 181 305 182 306 
<< pdiffusion >>
rect 192 305 193 306 
<< pdiffusion >>
rect 193 305 194 306 
<< pdiffusion >>
rect 194 305 195 306 
<< pdiffusion >>
rect 195 305 196 306 
<< pdiffusion >>
rect 196 305 197 306 
<< pdiffusion >>
rect 197 305 198 306 
<< m1 >>
rect 203 305 204 306 
<< m1 >>
rect 208 305 209 306 
<< pdiffusion >>
rect 210 305 211 306 
<< m1 >>
rect 211 305 212 306 
<< pdiffusion >>
rect 211 305 212 306 
<< pdiffusion >>
rect 212 305 213 306 
<< pdiffusion >>
rect 213 305 214 306 
<< m1 >>
rect 214 305 215 306 
<< pdiffusion >>
rect 214 305 215 306 
<< pdiffusion >>
rect 215 305 216 306 
<< m1 >>
rect 217 305 218 306 
<< m1 >>
rect 219 305 220 306 
<< m1 >>
rect 221 305 222 306 
<< m1 >>
rect 223 305 224 306 
<< pdiffusion >>
rect 228 305 229 306 
<< pdiffusion >>
rect 229 305 230 306 
<< pdiffusion >>
rect 230 305 231 306 
<< pdiffusion >>
rect 231 305 232 306 
<< pdiffusion >>
rect 232 305 233 306 
<< pdiffusion >>
rect 233 305 234 306 
<< m1 >>
rect 239 305 240 306 
<< pdiffusion >>
rect 246 305 247 306 
<< pdiffusion >>
rect 247 305 248 306 
<< pdiffusion >>
rect 248 305 249 306 
<< pdiffusion >>
rect 249 305 250 306 
<< pdiffusion >>
rect 250 305 251 306 
<< pdiffusion >>
rect 251 305 252 306 
<< m1 >>
rect 253 305 254 306 
<< m1 >>
rect 255 305 256 306 
<< pdiffusion >>
rect 264 305 265 306 
<< pdiffusion >>
rect 265 305 266 306 
<< pdiffusion >>
rect 266 305 267 306 
<< pdiffusion >>
rect 267 305 268 306 
<< pdiffusion >>
rect 268 305 269 306 
<< pdiffusion >>
rect 269 305 270 306 
<< m1 >>
rect 271 305 272 306 
<< m2 >>
rect 271 305 272 306 
<< m1 >>
rect 273 305 274 306 
<< m2 >>
rect 273 305 274 306 
<< m2c >>
rect 273 305 274 306 
<< m1 >>
rect 273 305 274 306 
<< m2 >>
rect 273 305 274 306 
<< m1 >>
rect 274 305 275 306 
<< m1 >>
rect 275 305 276 306 
<< m2 >>
rect 275 305 276 306 
<< m1 >>
rect 276 305 277 306 
<< m2 >>
rect 276 305 277 306 
<< m2 >>
rect 277 305 278 306 
<< m1 >>
rect 278 305 279 306 
<< m2 >>
rect 278 305 279 306 
<< m2c >>
rect 278 305 279 306 
<< m1 >>
rect 278 305 279 306 
<< m2 >>
rect 278 305 279 306 
<< pdiffusion >>
rect 282 305 283 306 
<< m1 >>
rect 283 305 284 306 
<< pdiffusion >>
rect 283 305 284 306 
<< pdiffusion >>
rect 284 305 285 306 
<< pdiffusion >>
rect 285 305 286 306 
<< m1 >>
rect 286 305 287 306 
<< pdiffusion >>
rect 286 305 287 306 
<< pdiffusion >>
rect 287 305 288 306 
<< pdiffusion >>
rect 300 305 301 306 
<< pdiffusion >>
rect 301 305 302 306 
<< pdiffusion >>
rect 302 305 303 306 
<< pdiffusion >>
rect 303 305 304 306 
<< pdiffusion >>
rect 304 305 305 306 
<< pdiffusion >>
rect 305 305 306 306 
<< pdiffusion >>
rect 318 305 319 306 
<< pdiffusion >>
rect 319 305 320 306 
<< pdiffusion >>
rect 320 305 321 306 
<< pdiffusion >>
rect 321 305 322 306 
<< pdiffusion >>
rect 322 305 323 306 
<< pdiffusion >>
rect 323 305 324 306 
<< m1 >>
rect 325 305 326 306 
<< m1 >>
rect 327 305 328 306 
<< m2 >>
rect 328 305 329 306 
<< m1 >>
rect 331 305 332 306 
<< m1 >>
rect 334 305 335 306 
<< pdiffusion >>
rect 336 305 337 306 
<< pdiffusion >>
rect 337 305 338 306 
<< pdiffusion >>
rect 338 305 339 306 
<< pdiffusion >>
rect 339 305 340 306 
<< pdiffusion >>
rect 340 305 341 306 
<< pdiffusion >>
rect 341 305 342 306 
<< m1 >>
rect 10 306 11 307 
<< m1 >>
rect 28 306 29 307 
<< m1 >>
rect 37 306 38 307 
<< m2 >>
rect 38 306 39 307 
<< m1 >>
rect 46 306 47 307 
<< m1 >>
rect 49 306 50 307 
<< m1 >>
rect 55 306 56 307 
<< m2 >>
rect 55 306 56 307 
<< m1 >>
rect 57 306 58 307 
<< m1 >>
rect 60 306 61 307 
<< m1 >>
rect 62 306 63 307 
<< m1 >>
rect 64 306 65 307 
<< m1 >>
rect 73 306 74 307 
<< m2 >>
rect 81 306 82 307 
<< m1 >>
rect 82 306 83 307 
<< m1 >>
rect 109 306 110 307 
<< m1 >>
rect 145 306 146 307 
<< m1 >>
rect 169 306 170 307 
<< m2 >>
rect 171 306 172 307 
<< m1 >>
rect 172 306 173 307 
<< m1 >>
rect 181 306 182 307 
<< m1 >>
rect 203 306 204 307 
<< m1 >>
rect 208 306 209 307 
<< m1 >>
rect 211 306 212 307 
<< m1 >>
rect 214 306 215 307 
<< m1 >>
rect 217 306 218 307 
<< m1 >>
rect 219 306 220 307 
<< m1 >>
rect 221 306 222 307 
<< m1 >>
rect 223 306 224 307 
<< m1 >>
rect 239 306 240 307 
<< m1 >>
rect 253 306 254 307 
<< m1 >>
rect 255 306 256 307 
<< m1 >>
rect 271 306 272 307 
<< m2 >>
rect 271 306 272 307 
<< m2 >>
rect 273 306 274 307 
<< m2 >>
rect 275 306 276 307 
<< m1 >>
rect 283 306 284 307 
<< m1 >>
rect 286 306 287 307 
<< m1 >>
rect 325 306 326 307 
<< m1 >>
rect 327 306 328 307 
<< m2 >>
rect 328 306 329 307 
<< m1 >>
rect 331 306 332 307 
<< m1 >>
rect 334 306 335 307 
<< m1 >>
rect 10 307 11 308 
<< m1 >>
rect 28 307 29 308 
<< m1 >>
rect 37 307 38 308 
<< m2 >>
rect 38 307 39 308 
<< m1 >>
rect 46 307 47 308 
<< m1 >>
rect 49 307 50 308 
<< m1 >>
rect 55 307 56 308 
<< m2 >>
rect 55 307 56 308 
<< m2 >>
rect 56 307 57 308 
<< m1 >>
rect 57 307 58 308 
<< m2 >>
rect 57 307 58 308 
<< m2 >>
rect 58 307 59 308 
<< m2 >>
rect 59 307 60 308 
<< m1 >>
rect 60 307 61 308 
<< m2 >>
rect 60 307 61 308 
<< m2 >>
rect 61 307 62 308 
<< m1 >>
rect 62 307 63 308 
<< m2 >>
rect 62 307 63 308 
<< m2 >>
rect 63 307 64 308 
<< m1 >>
rect 64 307 65 308 
<< m2 >>
rect 64 307 65 308 
<< m2 >>
rect 65 307 66 308 
<< m1 >>
rect 66 307 67 308 
<< m2 >>
rect 66 307 67 308 
<< m2c >>
rect 66 307 67 308 
<< m1 >>
rect 66 307 67 308 
<< m2 >>
rect 66 307 67 308 
<< m1 >>
rect 71 307 72 308 
<< m2 >>
rect 71 307 72 308 
<< m2c >>
rect 71 307 72 308 
<< m1 >>
rect 71 307 72 308 
<< m2 >>
rect 71 307 72 308 
<< m2 >>
rect 72 307 73 308 
<< m1 >>
rect 73 307 74 308 
<< m2 >>
rect 73 307 74 308 
<< m2 >>
rect 74 307 75 308 
<< m1 >>
rect 75 307 76 308 
<< m2 >>
rect 75 307 76 308 
<< m2c >>
rect 75 307 76 308 
<< m1 >>
rect 75 307 76 308 
<< m2 >>
rect 75 307 76 308 
<< m2 >>
rect 81 307 82 308 
<< m1 >>
rect 82 307 83 308 
<< m2 >>
rect 82 307 83 308 
<< m2 >>
rect 83 307 84 308 
<< m1 >>
rect 84 307 85 308 
<< m2 >>
rect 84 307 85 308 
<< m2c >>
rect 84 307 85 308 
<< m1 >>
rect 84 307 85 308 
<< m2 >>
rect 84 307 85 308 
<< m1 >>
rect 109 307 110 308 
<< m1 >>
rect 145 307 146 308 
<< m1 >>
rect 169 307 170 308 
<< m2 >>
rect 171 307 172 308 
<< m1 >>
rect 172 307 173 308 
<< m1 >>
rect 181 307 182 308 
<< m1 >>
rect 203 307 204 308 
<< m1 >>
rect 208 307 209 308 
<< m1 >>
rect 211 307 212 308 
<< m1 >>
rect 214 307 215 308 
<< m1 >>
rect 217 307 218 308 
<< m1 >>
rect 219 307 220 308 
<< m1 >>
rect 221 307 222 308 
<< m1 >>
rect 223 307 224 308 
<< m1 >>
rect 239 307 240 308 
<< m1 >>
rect 253 307 254 308 
<< m1 >>
rect 255 307 256 308 
<< m1 >>
rect 271 307 272 308 
<< m2 >>
rect 271 307 272 308 
<< m1 >>
rect 272 307 273 308 
<< m1 >>
rect 273 307 274 308 
<< m2 >>
rect 273 307 274 308 
<< m1 >>
rect 274 307 275 308 
<< m1 >>
rect 275 307 276 308 
<< m2 >>
rect 275 307 276 308 
<< m1 >>
rect 276 307 277 308 
<< m1 >>
rect 277 307 278 308 
<< m1 >>
rect 278 307 279 308 
<< m1 >>
rect 279 307 280 308 
<< m1 >>
rect 280 307 281 308 
<< m1 >>
rect 281 307 282 308 
<< m1 >>
rect 282 307 283 308 
<< m1 >>
rect 283 307 284 308 
<< m1 >>
rect 286 307 287 308 
<< m1 >>
rect 325 307 326 308 
<< m1 >>
rect 327 307 328 308 
<< m2 >>
rect 328 307 329 308 
<< m1 >>
rect 331 307 332 308 
<< m1 >>
rect 334 307 335 308 
<< m1 >>
rect 10 308 11 309 
<< m1 >>
rect 28 308 29 309 
<< m1 >>
rect 37 308 38 309 
<< m2 >>
rect 38 308 39 309 
<< m1 >>
rect 46 308 47 309 
<< m1 >>
rect 49 308 50 309 
<< m1 >>
rect 50 308 51 309 
<< m1 >>
rect 51 308 52 309 
<< m1 >>
rect 52 308 53 309 
<< m1 >>
rect 53 308 54 309 
<< m1 >>
rect 54 308 55 309 
<< m1 >>
rect 55 308 56 309 
<< m1 >>
rect 57 308 58 309 
<< m1 >>
rect 60 308 61 309 
<< m1 >>
rect 62 308 63 309 
<< m1 >>
rect 64 308 65 309 
<< m1 >>
rect 66 308 67 309 
<< m1 >>
rect 71 308 72 309 
<< m1 >>
rect 73 308 74 309 
<< m1 >>
rect 75 308 76 309 
<< m1 >>
rect 82 308 83 309 
<< m1 >>
rect 84 308 85 309 
<< m1 >>
rect 109 308 110 309 
<< m2 >>
rect 109 308 110 309 
<< m2c >>
rect 109 308 110 309 
<< m1 >>
rect 109 308 110 309 
<< m2 >>
rect 109 308 110 309 
<< m1 >>
rect 145 308 146 309 
<< m1 >>
rect 169 308 170 309 
<< m2 >>
rect 171 308 172 309 
<< m1 >>
rect 172 308 173 309 
<< m1 >>
rect 181 308 182 309 
<< m1 >>
rect 203 308 204 309 
<< m1 >>
rect 208 308 209 309 
<< m1 >>
rect 211 308 212 309 
<< m1 >>
rect 214 308 215 309 
<< m1 >>
rect 217 308 218 309 
<< m1 >>
rect 219 308 220 309 
<< m1 >>
rect 221 308 222 309 
<< m1 >>
rect 223 308 224 309 
<< m2 >>
rect 223 308 224 309 
<< m2c >>
rect 223 308 224 309 
<< m1 >>
rect 223 308 224 309 
<< m2 >>
rect 223 308 224 309 
<< m1 >>
rect 239 308 240 309 
<< m2 >>
rect 239 308 240 309 
<< m2c >>
rect 239 308 240 309 
<< m1 >>
rect 239 308 240 309 
<< m2 >>
rect 239 308 240 309 
<< m1 >>
rect 253 308 254 309 
<< m1 >>
rect 255 308 256 309 
<< m2 >>
rect 271 308 272 309 
<< m2 >>
rect 273 308 274 309 
<< m2 >>
rect 275 308 276 309 
<< m1 >>
rect 286 308 287 309 
<< m1 >>
rect 325 308 326 309 
<< m1 >>
rect 327 308 328 309 
<< m2 >>
rect 328 308 329 309 
<< m1 >>
rect 331 308 332 309 
<< m1 >>
rect 334 308 335 309 
<< m1 >>
rect 10 309 11 310 
<< m1 >>
rect 28 309 29 310 
<< m1 >>
rect 37 309 38 310 
<< m2 >>
rect 38 309 39 310 
<< m1 >>
rect 46 309 47 310 
<< m1 >>
rect 57 309 58 310 
<< m2 >>
rect 57 309 58 310 
<< m2c >>
rect 57 309 58 310 
<< m1 >>
rect 57 309 58 310 
<< m2 >>
rect 57 309 58 310 
<< m1 >>
rect 60 309 61 310 
<< m2 >>
rect 60 309 61 310 
<< m2c >>
rect 60 309 61 310 
<< m1 >>
rect 60 309 61 310 
<< m2 >>
rect 60 309 61 310 
<< m1 >>
rect 62 309 63 310 
<< m2 >>
rect 62 309 63 310 
<< m2c >>
rect 62 309 63 310 
<< m1 >>
rect 62 309 63 310 
<< m2 >>
rect 62 309 63 310 
<< m1 >>
rect 64 309 65 310 
<< m2 >>
rect 64 309 65 310 
<< m2c >>
rect 64 309 65 310 
<< m1 >>
rect 64 309 65 310 
<< m2 >>
rect 64 309 65 310 
<< m1 >>
rect 66 309 67 310 
<< m2 >>
rect 66 309 67 310 
<< m2c >>
rect 66 309 67 310 
<< m1 >>
rect 66 309 67 310 
<< m2 >>
rect 66 309 67 310 
<< m1 >>
rect 68 309 69 310 
<< m2 >>
rect 68 309 69 310 
<< m2c >>
rect 68 309 69 310 
<< m1 >>
rect 68 309 69 310 
<< m2 >>
rect 68 309 69 310 
<< m1 >>
rect 69 309 70 310 
<< m1 >>
rect 70 309 71 310 
<< m1 >>
rect 71 309 72 310 
<< m1 >>
rect 73 309 74 310 
<< m2 >>
rect 73 309 74 310 
<< m2c >>
rect 73 309 74 310 
<< m1 >>
rect 73 309 74 310 
<< m2 >>
rect 73 309 74 310 
<< m1 >>
rect 75 309 76 310 
<< m2 >>
rect 75 309 76 310 
<< m2c >>
rect 75 309 76 310 
<< m1 >>
rect 75 309 76 310 
<< m2 >>
rect 75 309 76 310 
<< m1 >>
rect 82 309 83 310 
<< m1 >>
rect 84 309 85 310 
<< m2 >>
rect 109 309 110 310 
<< m1 >>
rect 145 309 146 310 
<< m2 >>
rect 158 309 159 310 
<< m2 >>
rect 159 309 160 310 
<< m2 >>
rect 160 309 161 310 
<< m2 >>
rect 161 309 162 310 
<< m2 >>
rect 162 309 163 310 
<< m2 >>
rect 163 309 164 310 
<< m2 >>
rect 164 309 165 310 
<< m2 >>
rect 165 309 166 310 
<< m2 >>
rect 166 309 167 310 
<< m2 >>
rect 167 309 168 310 
<< m2 >>
rect 168 309 169 310 
<< m1 >>
rect 169 309 170 310 
<< m2 >>
rect 169 309 170 310 
<< m2 >>
rect 170 309 171 310 
<< m2 >>
rect 171 309 172 310 
<< m1 >>
rect 172 309 173 310 
<< m1 >>
rect 176 309 177 310 
<< m2 >>
rect 176 309 177 310 
<< m2c >>
rect 176 309 177 310 
<< m1 >>
rect 176 309 177 310 
<< m2 >>
rect 176 309 177 310 
<< m1 >>
rect 177 309 178 310 
<< m1 >>
rect 178 309 179 310 
<< m1 >>
rect 179 309 180 310 
<< m1 >>
rect 180 309 181 310 
<< m1 >>
rect 181 309 182 310 
<< m1 >>
rect 203 309 204 310 
<< m2 >>
rect 207 309 208 310 
<< m1 >>
rect 208 309 209 310 
<< m2 >>
rect 208 309 209 310 
<< m2 >>
rect 209 309 210 310 
<< m1 >>
rect 210 309 211 310 
<< m2 >>
rect 210 309 211 310 
<< m2c >>
rect 210 309 211 310 
<< m1 >>
rect 210 309 211 310 
<< m2 >>
rect 210 309 211 310 
<< m1 >>
rect 211 309 212 310 
<< m1 >>
rect 214 309 215 310 
<< m1 >>
rect 217 309 218 310 
<< m1 >>
rect 219 309 220 310 
<< m1 >>
rect 221 309 222 310 
<< m2 >>
rect 223 309 224 310 
<< m2 >>
rect 239 309 240 310 
<< m1 >>
rect 253 309 254 310 
<< m1 >>
rect 255 309 256 310 
<< m1 >>
rect 271 309 272 310 
<< m2 >>
rect 271 309 272 310 
<< m2c >>
rect 271 309 272 310 
<< m1 >>
rect 271 309 272 310 
<< m2 >>
rect 271 309 272 310 
<< m1 >>
rect 273 309 274 310 
<< m2 >>
rect 273 309 274 310 
<< m2c >>
rect 273 309 274 310 
<< m1 >>
rect 273 309 274 310 
<< m2 >>
rect 273 309 274 310 
<< m1 >>
rect 275 309 276 310 
<< m2 >>
rect 275 309 276 310 
<< m2c >>
rect 275 309 276 310 
<< m1 >>
rect 275 309 276 310 
<< m2 >>
rect 275 309 276 310 
<< m1 >>
rect 286 309 287 310 
<< m1 >>
rect 325 309 326 310 
<< m1 >>
rect 327 309 328 310 
<< m2 >>
rect 328 309 329 310 
<< m1 >>
rect 331 309 332 310 
<< m1 >>
rect 334 309 335 310 
<< m1 >>
rect 10 310 11 311 
<< m1 >>
rect 28 310 29 311 
<< m1 >>
rect 37 310 38 311 
<< m2 >>
rect 38 310 39 311 
<< m1 >>
rect 46 310 47 311 
<< m2 >>
rect 57 310 58 311 
<< m2 >>
rect 60 310 61 311 
<< m2 >>
rect 62 310 63 311 
<< m2 >>
rect 64 310 65 311 
<< m2 >>
rect 66 310 67 311 
<< m2 >>
rect 67 310 68 311 
<< m2 >>
rect 68 310 69 311 
<< m2 >>
rect 73 310 74 311 
<< m2 >>
rect 75 310 76 311 
<< m1 >>
rect 82 310 83 311 
<< m1 >>
rect 84 310 85 311 
<< m1 >>
rect 85 310 86 311 
<< m1 >>
rect 86 310 87 311 
<< m1 >>
rect 87 310 88 311 
<< m1 >>
rect 88 310 89 311 
<< m1 >>
rect 89 310 90 311 
<< m1 >>
rect 90 310 91 311 
<< m1 >>
rect 91 310 92 311 
<< m1 >>
rect 92 310 93 311 
<< m1 >>
rect 93 310 94 311 
<< m1 >>
rect 94 310 95 311 
<< m1 >>
rect 95 310 96 311 
<< m1 >>
rect 96 310 97 311 
<< m1 >>
rect 97 310 98 311 
<< m1 >>
rect 98 310 99 311 
<< m1 >>
rect 99 310 100 311 
<< m1 >>
rect 100 310 101 311 
<< m1 >>
rect 101 310 102 311 
<< m1 >>
rect 102 310 103 311 
<< m1 >>
rect 103 310 104 311 
<< m1 >>
rect 104 310 105 311 
<< m1 >>
rect 105 310 106 311 
<< m1 >>
rect 106 310 107 311 
<< m1 >>
rect 107 310 108 311 
<< m1 >>
rect 108 310 109 311 
<< m1 >>
rect 109 310 110 311 
<< m2 >>
rect 109 310 110 311 
<< m1 >>
rect 110 310 111 311 
<< m2 >>
rect 110 310 111 311 
<< m1 >>
rect 111 310 112 311 
<< m2 >>
rect 111 310 112 311 
<< m1 >>
rect 112 310 113 311 
<< m2 >>
rect 112 310 113 311 
<< m1 >>
rect 113 310 114 311 
<< m2 >>
rect 113 310 114 311 
<< m1 >>
rect 114 310 115 311 
<< m2 >>
rect 114 310 115 311 
<< m1 >>
rect 115 310 116 311 
<< m2 >>
rect 115 310 116 311 
<< m1 >>
rect 116 310 117 311 
<< m2 >>
rect 116 310 117 311 
<< m1 >>
rect 117 310 118 311 
<< m2 >>
rect 117 310 118 311 
<< m1 >>
rect 118 310 119 311 
<< m2 >>
rect 118 310 119 311 
<< m1 >>
rect 119 310 120 311 
<< m2 >>
rect 119 310 120 311 
<< m1 >>
rect 120 310 121 311 
<< m2 >>
rect 120 310 121 311 
<< m1 >>
rect 121 310 122 311 
<< m2 >>
rect 121 310 122 311 
<< m1 >>
rect 122 310 123 311 
<< m2 >>
rect 122 310 123 311 
<< m1 >>
rect 123 310 124 311 
<< m2 >>
rect 123 310 124 311 
<< m1 >>
rect 124 310 125 311 
<< m2 >>
rect 124 310 125 311 
<< m1 >>
rect 125 310 126 311 
<< m2 >>
rect 125 310 126 311 
<< m1 >>
rect 126 310 127 311 
<< m2 >>
rect 126 310 127 311 
<< m1 >>
rect 127 310 128 311 
<< m2 >>
rect 127 310 128 311 
<< m1 >>
rect 128 310 129 311 
<< m2 >>
rect 128 310 129 311 
<< m1 >>
rect 129 310 130 311 
<< m2 >>
rect 129 310 130 311 
<< m1 >>
rect 130 310 131 311 
<< m2 >>
rect 130 310 131 311 
<< m1 >>
rect 131 310 132 311 
<< m2 >>
rect 131 310 132 311 
<< m1 >>
rect 132 310 133 311 
<< m2 >>
rect 132 310 133 311 
<< m1 >>
rect 133 310 134 311 
<< m2 >>
rect 133 310 134 311 
<< m1 >>
rect 134 310 135 311 
<< m2 >>
rect 134 310 135 311 
<< m1 >>
rect 135 310 136 311 
<< m2 >>
rect 135 310 136 311 
<< m1 >>
rect 136 310 137 311 
<< m2 >>
rect 136 310 137 311 
<< m1 >>
rect 137 310 138 311 
<< m2 >>
rect 137 310 138 311 
<< m1 >>
rect 138 310 139 311 
<< m2 >>
rect 138 310 139 311 
<< m1 >>
rect 139 310 140 311 
<< m2 >>
rect 139 310 140 311 
<< m1 >>
rect 140 310 141 311 
<< m2 >>
rect 140 310 141 311 
<< m1 >>
rect 141 310 142 311 
<< m2 >>
rect 141 310 142 311 
<< m1 >>
rect 142 310 143 311 
<< m2 >>
rect 142 310 143 311 
<< m1 >>
rect 143 310 144 311 
<< m2 >>
rect 143 310 144 311 
<< m1 >>
rect 144 310 145 311 
<< m2 >>
rect 144 310 145 311 
<< m1 >>
rect 145 310 146 311 
<< m2 >>
rect 145 310 146 311 
<< m2 >>
rect 146 310 147 311 
<< m1 >>
rect 147 310 148 311 
<< m2 >>
rect 147 310 148 311 
<< m2c >>
rect 147 310 148 311 
<< m1 >>
rect 147 310 148 311 
<< m2 >>
rect 147 310 148 311 
<< m1 >>
rect 148 310 149 311 
<< m1 >>
rect 149 310 150 311 
<< m1 >>
rect 150 310 151 311 
<< m1 >>
rect 151 310 152 311 
<< m1 >>
rect 152 310 153 311 
<< m1 >>
rect 153 310 154 311 
<< m1 >>
rect 154 310 155 311 
<< m1 >>
rect 155 310 156 311 
<< m1 >>
rect 156 310 157 311 
<< m1 >>
rect 157 310 158 311 
<< m1 >>
rect 158 310 159 311 
<< m2 >>
rect 158 310 159 311 
<< m1 >>
rect 159 310 160 311 
<< m1 >>
rect 160 310 161 311 
<< m1 >>
rect 161 310 162 311 
<< m1 >>
rect 162 310 163 311 
<< m1 >>
rect 163 310 164 311 
<< m1 >>
rect 164 310 165 311 
<< m1 >>
rect 165 310 166 311 
<< m1 >>
rect 166 310 167 311 
<< m1 >>
rect 167 310 168 311 
<< m1 >>
rect 168 310 169 311 
<< m1 >>
rect 169 310 170 311 
<< m1 >>
rect 172 310 173 311 
<< m2 >>
rect 176 310 177 311 
<< m1 >>
rect 203 310 204 311 
<< m2 >>
rect 207 310 208 311 
<< m1 >>
rect 208 310 209 311 
<< m1 >>
rect 214 310 215 311 
<< m1 >>
rect 217 310 218 311 
<< m1 >>
rect 219 310 220 311 
<< m1 >>
rect 221 310 222 311 
<< m1 >>
rect 222 310 223 311 
<< m1 >>
rect 223 310 224 311 
<< m2 >>
rect 223 310 224 311 
<< m1 >>
rect 224 310 225 311 
<< m1 >>
rect 225 310 226 311 
<< m1 >>
rect 226 310 227 311 
<< m1 >>
rect 227 310 228 311 
<< m1 >>
rect 228 310 229 311 
<< m1 >>
rect 229 310 230 311 
<< m1 >>
rect 230 310 231 311 
<< m1 >>
rect 231 310 232 311 
<< m1 >>
rect 232 310 233 311 
<< m1 >>
rect 233 310 234 311 
<< m1 >>
rect 234 310 235 311 
<< m1 >>
rect 235 310 236 311 
<< m1 >>
rect 236 310 237 311 
<< m1 >>
rect 237 310 238 311 
<< m1 >>
rect 238 310 239 311 
<< m1 >>
rect 239 310 240 311 
<< m2 >>
rect 239 310 240 311 
<< m1 >>
rect 240 310 241 311 
<< m1 >>
rect 241 310 242 311 
<< m1 >>
rect 242 310 243 311 
<< m1 >>
rect 243 310 244 311 
<< m1 >>
rect 244 310 245 311 
<< m1 >>
rect 245 310 246 311 
<< m1 >>
rect 246 310 247 311 
<< m1 >>
rect 247 310 248 311 
<< m1 >>
rect 248 310 249 311 
<< m1 >>
rect 249 310 250 311 
<< m1 >>
rect 250 310 251 311 
<< m1 >>
rect 251 310 252 311 
<< m2 >>
rect 251 310 252 311 
<< m2c >>
rect 251 310 252 311 
<< m1 >>
rect 251 310 252 311 
<< m2 >>
rect 251 310 252 311 
<< m2 >>
rect 252 310 253 311 
<< m1 >>
rect 253 310 254 311 
<< m2 >>
rect 253 310 254 311 
<< m2 >>
rect 254 310 255 311 
<< m1 >>
rect 255 310 256 311 
<< m2 >>
rect 255 310 256 311 
<< m2 >>
rect 256 310 257 311 
<< m2 >>
rect 257 310 258 311 
<< m2 >>
rect 258 310 259 311 
<< m2 >>
rect 259 310 260 311 
<< m2 >>
rect 260 310 261 311 
<< m2 >>
rect 261 310 262 311 
<< m2 >>
rect 262 310 263 311 
<< m2 >>
rect 263 310 264 311 
<< m2 >>
rect 264 310 265 311 
<< m2 >>
rect 265 310 266 311 
<< m2 >>
rect 266 310 267 311 
<< m1 >>
rect 271 310 272 311 
<< m1 >>
rect 273 310 274 311 
<< m1 >>
rect 275 310 276 311 
<< m1 >>
rect 286 310 287 311 
<< m1 >>
rect 325 310 326 311 
<< m1 >>
rect 327 310 328 311 
<< m2 >>
rect 328 310 329 311 
<< m1 >>
rect 331 310 332 311 
<< m1 >>
rect 334 310 335 311 
<< m1 >>
rect 10 311 11 312 
<< m1 >>
rect 28 311 29 312 
<< m1 >>
rect 37 311 38 312 
<< m2 >>
rect 38 311 39 312 
<< m1 >>
rect 46 311 47 312 
<< m1 >>
rect 55 311 56 312 
<< m2 >>
rect 55 311 56 312 
<< m2c >>
rect 55 311 56 312 
<< m1 >>
rect 55 311 56 312 
<< m2 >>
rect 55 311 56 312 
<< m1 >>
rect 56 311 57 312 
<< m1 >>
rect 57 311 58 312 
<< m2 >>
rect 57 311 58 312 
<< m1 >>
rect 58 311 59 312 
<< m1 >>
rect 59 311 60 312 
<< m1 >>
rect 60 311 61 312 
<< m2 >>
rect 60 311 61 312 
<< m1 >>
rect 61 311 62 312 
<< m1 >>
rect 62 311 63 312 
<< m2 >>
rect 62 311 63 312 
<< m1 >>
rect 63 311 64 312 
<< m1 >>
rect 64 311 65 312 
<< m2 >>
rect 64 311 65 312 
<< m1 >>
rect 65 311 66 312 
<< m1 >>
rect 66 311 67 312 
<< m1 >>
rect 67 311 68 312 
<< m1 >>
rect 68 311 69 312 
<< m1 >>
rect 69 311 70 312 
<< m1 >>
rect 70 311 71 312 
<< m1 >>
rect 71 311 72 312 
<< m1 >>
rect 72 311 73 312 
<< m1 >>
rect 73 311 74 312 
<< m2 >>
rect 73 311 74 312 
<< m1 >>
rect 74 311 75 312 
<< m1 >>
rect 75 311 76 312 
<< m2 >>
rect 75 311 76 312 
<< m1 >>
rect 76 311 77 312 
<< m1 >>
rect 77 311 78 312 
<< m1 >>
rect 78 311 79 312 
<< m1 >>
rect 79 311 80 312 
<< m1 >>
rect 80 311 81 312 
<< m2 >>
rect 80 311 81 312 
<< m2c >>
rect 80 311 81 312 
<< m1 >>
rect 80 311 81 312 
<< m2 >>
rect 80 311 81 312 
<< m2 >>
rect 81 311 82 312 
<< m1 >>
rect 82 311 83 312 
<< m2 >>
rect 82 311 83 312 
<< m2 >>
rect 83 311 84 312 
<< m2 >>
rect 84 311 85 312 
<< m2 >>
rect 85 311 86 312 
<< m2 >>
rect 86 311 87 312 
<< m2 >>
rect 158 311 159 312 
<< m2 >>
rect 171 311 172 312 
<< m1 >>
rect 172 311 173 312 
<< m2 >>
rect 172 311 173 312 
<< m2 >>
rect 173 311 174 312 
<< m1 >>
rect 174 311 175 312 
<< m2 >>
rect 174 311 175 312 
<< m2c >>
rect 174 311 175 312 
<< m1 >>
rect 174 311 175 312 
<< m2 >>
rect 174 311 175 312 
<< m1 >>
rect 175 311 176 312 
<< m1 >>
rect 176 311 177 312 
<< m2 >>
rect 176 311 177 312 
<< m1 >>
rect 177 311 178 312 
<< m1 >>
rect 178 311 179 312 
<< m1 >>
rect 179 311 180 312 
<< m1 >>
rect 180 311 181 312 
<< m1 >>
rect 181 311 182 312 
<< m1 >>
rect 182 311 183 312 
<< m1 >>
rect 183 311 184 312 
<< m1 >>
rect 184 311 185 312 
<< m1 >>
rect 185 311 186 312 
<< m1 >>
rect 186 311 187 312 
<< m1 >>
rect 187 311 188 312 
<< m1 >>
rect 188 311 189 312 
<< m1 >>
rect 189 311 190 312 
<< m1 >>
rect 190 311 191 312 
<< m1 >>
rect 191 311 192 312 
<< m1 >>
rect 192 311 193 312 
<< m1 >>
rect 193 311 194 312 
<< m1 >>
rect 194 311 195 312 
<< m1 >>
rect 195 311 196 312 
<< m1 >>
rect 196 311 197 312 
<< m1 >>
rect 197 311 198 312 
<< m1 >>
rect 198 311 199 312 
<< m1 >>
rect 199 311 200 312 
<< m1 >>
rect 200 311 201 312 
<< m1 >>
rect 201 311 202 312 
<< m1 >>
rect 202 311 203 312 
<< m1 >>
rect 203 311 204 312 
<< m2 >>
rect 207 311 208 312 
<< m1 >>
rect 208 311 209 312 
<< m1 >>
rect 209 311 210 312 
<< m1 >>
rect 210 311 211 312 
<< m1 >>
rect 211 311 212 312 
<< m2 >>
rect 211 311 212 312 
<< m2c >>
rect 211 311 212 312 
<< m1 >>
rect 211 311 212 312 
<< m2 >>
rect 211 311 212 312 
<< m1 >>
rect 214 311 215 312 
<< m2 >>
rect 214 311 215 312 
<< m2c >>
rect 214 311 215 312 
<< m1 >>
rect 214 311 215 312 
<< m2 >>
rect 214 311 215 312 
<< m1 >>
rect 217 311 218 312 
<< m2 >>
rect 217 311 218 312 
<< m2c >>
rect 217 311 218 312 
<< m1 >>
rect 217 311 218 312 
<< m2 >>
rect 217 311 218 312 
<< m1 >>
rect 219 311 220 312 
<< m2 >>
rect 219 311 220 312 
<< m2c >>
rect 219 311 220 312 
<< m1 >>
rect 219 311 220 312 
<< m2 >>
rect 219 311 220 312 
<< m2 >>
rect 223 311 224 312 
<< m2 >>
rect 239 311 240 312 
<< m1 >>
rect 253 311 254 312 
<< m1 >>
rect 255 311 256 312 
<< m1 >>
rect 256 311 257 312 
<< m1 >>
rect 257 311 258 312 
<< m1 >>
rect 258 311 259 312 
<< m1 >>
rect 259 311 260 312 
<< m1 >>
rect 260 311 261 312 
<< m1 >>
rect 261 311 262 312 
<< m1 >>
rect 262 311 263 312 
<< m1 >>
rect 263 311 264 312 
<< m1 >>
rect 264 311 265 312 
<< m1 >>
rect 265 311 266 312 
<< m1 >>
rect 266 311 267 312 
<< m2 >>
rect 266 311 267 312 
<< m1 >>
rect 267 311 268 312 
<< m1 >>
rect 268 311 269 312 
<< m1 >>
rect 269 311 270 312 
<< m2 >>
rect 269 311 270 312 
<< m2c >>
rect 269 311 270 312 
<< m1 >>
rect 269 311 270 312 
<< m2 >>
rect 269 311 270 312 
<< m2 >>
rect 270 311 271 312 
<< m1 >>
rect 271 311 272 312 
<< m2 >>
rect 271 311 272 312 
<< m2 >>
rect 272 311 273 312 
<< m1 >>
rect 273 311 274 312 
<< m2 >>
rect 273 311 274 312 
<< m2 >>
rect 274 311 275 312 
<< m1 >>
rect 275 311 276 312 
<< m2 >>
rect 275 311 276 312 
<< m2 >>
rect 276 311 277 312 
<< m1 >>
rect 277 311 278 312 
<< m2 >>
rect 277 311 278 312 
<< m2c >>
rect 277 311 278 312 
<< m1 >>
rect 277 311 278 312 
<< m2 >>
rect 277 311 278 312 
<< m1 >>
rect 278 311 279 312 
<< m1 >>
rect 279 311 280 312 
<< m1 >>
rect 280 311 281 312 
<< m1 >>
rect 281 311 282 312 
<< m1 >>
rect 282 311 283 312 
<< m1 >>
rect 283 311 284 312 
<< m1 >>
rect 284 311 285 312 
<< m1 >>
rect 285 311 286 312 
<< m1 >>
rect 286 311 287 312 
<< m1 >>
rect 325 311 326 312 
<< m1 >>
rect 327 311 328 312 
<< m2 >>
rect 328 311 329 312 
<< m1 >>
rect 329 311 330 312 
<< m2 >>
rect 329 311 330 312 
<< m2c >>
rect 329 311 330 312 
<< m1 >>
rect 329 311 330 312 
<< m2 >>
rect 329 311 330 312 
<< m2 >>
rect 330 311 331 312 
<< m1 >>
rect 331 311 332 312 
<< m2 >>
rect 331 311 332 312 
<< m2 >>
rect 332 311 333 312 
<< m2 >>
rect 333 311 334 312 
<< m1 >>
rect 334 311 335 312 
<< m2 >>
rect 334 311 335 312 
<< m2 >>
rect 335 311 336 312 
<< m1 >>
rect 10 312 11 313 
<< m1 >>
rect 28 312 29 313 
<< m1 >>
rect 37 312 38 313 
<< m2 >>
rect 38 312 39 313 
<< m1 >>
rect 46 312 47 313 
<< m2 >>
rect 55 312 56 313 
<< m2 >>
rect 57 312 58 313 
<< m2 >>
rect 60 312 61 313 
<< m2 >>
rect 62 312 63 313 
<< m2 >>
rect 64 312 65 313 
<< m2 >>
rect 73 312 74 313 
<< m2 >>
rect 75 312 76 313 
<< m1 >>
rect 82 312 83 313 
<< m2 >>
rect 86 312 87 313 
<< m2 >>
rect 87 312 88 313 
<< m2 >>
rect 88 312 89 313 
<< m2 >>
rect 89 312 90 313 
<< m2 >>
rect 90 312 91 313 
<< m2 >>
rect 91 312 92 313 
<< m2 >>
rect 92 312 93 313 
<< m2 >>
rect 93 312 94 313 
<< m2 >>
rect 94 312 95 313 
<< m2 >>
rect 95 312 96 313 
<< m2 >>
rect 96 312 97 313 
<< m2 >>
rect 97 312 98 313 
<< m2 >>
rect 98 312 99 313 
<< m2 >>
rect 99 312 100 313 
<< m2 >>
rect 100 312 101 313 
<< m2 >>
rect 101 312 102 313 
<< m2 >>
rect 102 312 103 313 
<< m2 >>
rect 103 312 104 313 
<< m2 >>
rect 104 312 105 313 
<< m2 >>
rect 105 312 106 313 
<< m2 >>
rect 106 312 107 313 
<< m2 >>
rect 107 312 108 313 
<< m2 >>
rect 108 312 109 313 
<< m2 >>
rect 109 312 110 313 
<< m2 >>
rect 110 312 111 313 
<< m2 >>
rect 111 312 112 313 
<< m2 >>
rect 112 312 113 313 
<< m2 >>
rect 113 312 114 313 
<< m2 >>
rect 114 312 115 313 
<< m2 >>
rect 115 312 116 313 
<< m2 >>
rect 116 312 117 313 
<< m2 >>
rect 117 312 118 313 
<< m2 >>
rect 118 312 119 313 
<< m2 >>
rect 119 312 120 313 
<< m2 >>
rect 120 312 121 313 
<< m2 >>
rect 121 312 122 313 
<< m2 >>
rect 122 312 123 313 
<< m2 >>
rect 123 312 124 313 
<< m2 >>
rect 124 312 125 313 
<< m2 >>
rect 125 312 126 313 
<< m2 >>
rect 126 312 127 313 
<< m2 >>
rect 127 312 128 313 
<< m2 >>
rect 128 312 129 313 
<< m2 >>
rect 129 312 130 313 
<< m2 >>
rect 130 312 131 313 
<< m2 >>
rect 131 312 132 313 
<< m2 >>
rect 132 312 133 313 
<< m2 >>
rect 133 312 134 313 
<< m2 >>
rect 134 312 135 313 
<< m2 >>
rect 135 312 136 313 
<< m2 >>
rect 136 312 137 313 
<< m2 >>
rect 137 312 138 313 
<< m2 >>
rect 138 312 139 313 
<< m2 >>
rect 139 312 140 313 
<< m2 >>
rect 140 312 141 313 
<< m2 >>
rect 141 312 142 313 
<< m2 >>
rect 142 312 143 313 
<< m2 >>
rect 143 312 144 313 
<< m2 >>
rect 144 312 145 313 
<< m2 >>
rect 145 312 146 313 
<< m2 >>
rect 146 312 147 313 
<< m2 >>
rect 147 312 148 313 
<< m2 >>
rect 148 312 149 313 
<< m2 >>
rect 149 312 150 313 
<< m2 >>
rect 150 312 151 313 
<< m2 >>
rect 151 312 152 313 
<< m2 >>
rect 152 312 153 313 
<< m2 >>
rect 153 312 154 313 
<< m2 >>
rect 154 312 155 313 
<< m2 >>
rect 155 312 156 313 
<< m2 >>
rect 156 312 157 313 
<< m2 >>
rect 157 312 158 313 
<< m2 >>
rect 158 312 159 313 
<< m2 >>
rect 171 312 172 313 
<< m1 >>
rect 172 312 173 313 
<< m2 >>
rect 176 312 177 313 
<< m2 >>
rect 207 312 208 313 
<< m2 >>
rect 211 312 212 313 
<< m2 >>
rect 214 312 215 313 
<< m2 >>
rect 217 312 218 313 
<< m2 >>
rect 219 312 220 313 
<< m2 >>
rect 223 312 224 313 
<< m1 >>
rect 239 312 240 313 
<< m2 >>
rect 239 312 240 313 
<< m2c >>
rect 239 312 240 313 
<< m1 >>
rect 239 312 240 313 
<< m2 >>
rect 239 312 240 313 
<< m1 >>
rect 253 312 254 313 
<< m2 >>
rect 266 312 267 313 
<< m1 >>
rect 271 312 272 313 
<< m1 >>
rect 273 312 274 313 
<< m1 >>
rect 275 312 276 313 
<< m1 >>
rect 325 312 326 313 
<< m1 >>
rect 327 312 328 313 
<< m1 >>
rect 331 312 332 313 
<< m1 >>
rect 334 312 335 313 
<< m2 >>
rect 335 312 336 313 
<< m1 >>
rect 10 313 11 314 
<< m1 >>
rect 28 313 29 314 
<< m1 >>
rect 37 313 38 314 
<< m2 >>
rect 38 313 39 314 
<< m1 >>
rect 46 313 47 314 
<< m1 >>
rect 49 313 50 314 
<< m1 >>
rect 50 313 51 314 
<< m1 >>
rect 51 313 52 314 
<< m1 >>
rect 52 313 53 314 
<< m1 >>
rect 53 313 54 314 
<< m1 >>
rect 54 313 55 314 
<< m1 >>
rect 55 313 56 314 
<< m2 >>
rect 55 313 56 314 
<< m1 >>
rect 56 313 57 314 
<< m1 >>
rect 57 313 58 314 
<< m2 >>
rect 57 313 58 314 
<< m1 >>
rect 58 313 59 314 
<< m1 >>
rect 59 313 60 314 
<< m1 >>
rect 60 313 61 314 
<< m2 >>
rect 60 313 61 314 
<< m1 >>
rect 61 313 62 314 
<< m1 >>
rect 62 313 63 314 
<< m2 >>
rect 62 313 63 314 
<< m1 >>
rect 63 313 64 314 
<< m1 >>
rect 64 313 65 314 
<< m2 >>
rect 64 313 65 314 
<< m1 >>
rect 65 313 66 314 
<< m1 >>
rect 66 313 67 314 
<< m1 >>
rect 67 313 68 314 
<< m1 >>
rect 68 313 69 314 
<< m1 >>
rect 69 313 70 314 
<< m1 >>
rect 70 313 71 314 
<< m1 >>
rect 71 313 72 314 
<< m1 >>
rect 72 313 73 314 
<< m1 >>
rect 73 313 74 314 
<< m2 >>
rect 73 313 74 314 
<< m1 >>
rect 74 313 75 314 
<< m1 >>
rect 75 313 76 314 
<< m2 >>
rect 75 313 76 314 
<< m1 >>
rect 76 313 77 314 
<< m1 >>
rect 77 313 78 314 
<< m1 >>
rect 78 313 79 314 
<< m1 >>
rect 79 313 80 314 
<< m1 >>
rect 80 313 81 314 
<< m2 >>
rect 80 313 81 314 
<< m2c >>
rect 80 313 81 314 
<< m1 >>
rect 80 313 81 314 
<< m2 >>
rect 80 313 81 314 
<< m2 >>
rect 81 313 82 314 
<< m1 >>
rect 82 313 83 314 
<< m2 >>
rect 82 313 83 314 
<< m2 >>
rect 83 313 84 314 
<< m1 >>
rect 84 313 85 314 
<< m2 >>
rect 84 313 85 314 
<< m2c >>
rect 84 313 85 314 
<< m1 >>
rect 84 313 85 314 
<< m2 >>
rect 84 313 85 314 
<< m1 >>
rect 85 313 86 314 
<< m1 >>
rect 86 313 87 314 
<< m1 >>
rect 87 313 88 314 
<< m1 >>
rect 88 313 89 314 
<< m1 >>
rect 89 313 90 314 
<< m1 >>
rect 90 313 91 314 
<< m1 >>
rect 91 313 92 314 
<< m1 >>
rect 92 313 93 314 
<< m1 >>
rect 93 313 94 314 
<< m1 >>
rect 94 313 95 314 
<< m1 >>
rect 95 313 96 314 
<< m1 >>
rect 96 313 97 314 
<< m1 >>
rect 97 313 98 314 
<< m1 >>
rect 98 313 99 314 
<< m1 >>
rect 99 313 100 314 
<< m1 >>
rect 100 313 101 314 
<< m1 >>
rect 101 313 102 314 
<< m1 >>
rect 102 313 103 314 
<< m1 >>
rect 103 313 104 314 
<< m1 >>
rect 104 313 105 314 
<< m1 >>
rect 105 313 106 314 
<< m1 >>
rect 106 313 107 314 
<< m1 >>
rect 107 313 108 314 
<< m1 >>
rect 108 313 109 314 
<< m1 >>
rect 109 313 110 314 
<< m1 >>
rect 110 313 111 314 
<< m1 >>
rect 111 313 112 314 
<< m1 >>
rect 112 313 113 314 
<< m1 >>
rect 113 313 114 314 
<< m1 >>
rect 114 313 115 314 
<< m1 >>
rect 115 313 116 314 
<< m1 >>
rect 116 313 117 314 
<< m1 >>
rect 117 313 118 314 
<< m1 >>
rect 118 313 119 314 
<< m1 >>
rect 119 313 120 314 
<< m1 >>
rect 120 313 121 314 
<< m1 >>
rect 121 313 122 314 
<< m1 >>
rect 122 313 123 314 
<< m1 >>
rect 123 313 124 314 
<< m1 >>
rect 124 313 125 314 
<< m1 >>
rect 125 313 126 314 
<< m1 >>
rect 126 313 127 314 
<< m1 >>
rect 127 313 128 314 
<< m1 >>
rect 128 313 129 314 
<< m1 >>
rect 129 313 130 314 
<< m1 >>
rect 130 313 131 314 
<< m1 >>
rect 131 313 132 314 
<< m1 >>
rect 132 313 133 314 
<< m1 >>
rect 133 313 134 314 
<< m1 >>
rect 134 313 135 314 
<< m1 >>
rect 135 313 136 314 
<< m1 >>
rect 136 313 137 314 
<< m1 >>
rect 137 313 138 314 
<< m1 >>
rect 138 313 139 314 
<< m1 >>
rect 139 313 140 314 
<< m1 >>
rect 140 313 141 314 
<< m1 >>
rect 141 313 142 314 
<< m1 >>
rect 142 313 143 314 
<< m1 >>
rect 143 313 144 314 
<< m1 >>
rect 144 313 145 314 
<< m1 >>
rect 145 313 146 314 
<< m1 >>
rect 146 313 147 314 
<< m1 >>
rect 147 313 148 314 
<< m1 >>
rect 148 313 149 314 
<< m1 >>
rect 149 313 150 314 
<< m1 >>
rect 150 313 151 314 
<< m1 >>
rect 151 313 152 314 
<< m1 >>
rect 152 313 153 314 
<< m1 >>
rect 153 313 154 314 
<< m1 >>
rect 154 313 155 314 
<< m1 >>
rect 155 313 156 314 
<< m1 >>
rect 156 313 157 314 
<< m1 >>
rect 157 313 158 314 
<< m1 >>
rect 158 313 159 314 
<< m1 >>
rect 159 313 160 314 
<< m1 >>
rect 160 313 161 314 
<< m1 >>
rect 161 313 162 314 
<< m1 >>
rect 162 313 163 314 
<< m1 >>
rect 163 313 164 314 
<< m1 >>
rect 164 313 165 314 
<< m1 >>
rect 165 313 166 314 
<< m1 >>
rect 166 313 167 314 
<< m1 >>
rect 167 313 168 314 
<< m1 >>
rect 168 313 169 314 
<< m1 >>
rect 169 313 170 314 
<< m1 >>
rect 170 313 171 314 
<< m2 >>
rect 170 313 171 314 
<< m2c >>
rect 170 313 171 314 
<< m1 >>
rect 170 313 171 314 
<< m2 >>
rect 170 313 171 314 
<< m2 >>
rect 171 313 172 314 
<< m1 >>
rect 172 313 173 314 
<< m2 >>
rect 172 313 173 314 
<< m1 >>
rect 173 313 174 314 
<< m2 >>
rect 173 313 174 314 
<< m1 >>
rect 174 313 175 314 
<< m2 >>
rect 174 313 175 314 
<< m1 >>
rect 175 313 176 314 
<< m2 >>
rect 175 313 176 314 
<< m1 >>
rect 176 313 177 314 
<< m2 >>
rect 176 313 177 314 
<< m1 >>
rect 177 313 178 314 
<< m1 >>
rect 178 313 179 314 
<< m1 >>
rect 179 313 180 314 
<< m1 >>
rect 180 313 181 314 
<< m1 >>
rect 181 313 182 314 
<< m1 >>
rect 182 313 183 314 
<< m1 >>
rect 183 313 184 314 
<< m1 >>
rect 184 313 185 314 
<< m1 >>
rect 185 313 186 314 
<< m1 >>
rect 186 313 187 314 
<< m1 >>
rect 187 313 188 314 
<< m1 >>
rect 188 313 189 314 
<< m1 >>
rect 189 313 190 314 
<< m1 >>
rect 190 313 191 314 
<< m1 >>
rect 191 313 192 314 
<< m1 >>
rect 192 313 193 314 
<< m1 >>
rect 193 313 194 314 
<< m1 >>
rect 194 313 195 314 
<< m1 >>
rect 195 313 196 314 
<< m1 >>
rect 196 313 197 314 
<< m1 >>
rect 197 313 198 314 
<< m1 >>
rect 198 313 199 314 
<< m1 >>
rect 199 313 200 314 
<< m1 >>
rect 200 313 201 314 
<< m1 >>
rect 201 313 202 314 
<< m1 >>
rect 202 313 203 314 
<< m1 >>
rect 203 313 204 314 
<< m1 >>
rect 204 313 205 314 
<< m1 >>
rect 205 313 206 314 
<< m1 >>
rect 206 313 207 314 
<< m1 >>
rect 207 313 208 314 
<< m2 >>
rect 207 313 208 314 
<< m1 >>
rect 208 313 209 314 
<< m1 >>
rect 209 313 210 314 
<< m1 >>
rect 210 313 211 314 
<< m1 >>
rect 211 313 212 314 
<< m2 >>
rect 211 313 212 314 
<< m1 >>
rect 212 313 213 314 
<< m1 >>
rect 213 313 214 314 
<< m1 >>
rect 214 313 215 314 
<< m2 >>
rect 214 313 215 314 
<< m1 >>
rect 215 313 216 314 
<< m1 >>
rect 216 313 217 314 
<< m1 >>
rect 217 313 218 314 
<< m2 >>
rect 217 313 218 314 
<< m1 >>
rect 218 313 219 314 
<< m1 >>
rect 219 313 220 314 
<< m2 >>
rect 219 313 220 314 
<< m1 >>
rect 220 313 221 314 
<< m1 >>
rect 221 313 222 314 
<< m1 >>
rect 222 313 223 314 
<< m1 >>
rect 223 313 224 314 
<< m2 >>
rect 223 313 224 314 
<< m1 >>
rect 224 313 225 314 
<< m1 >>
rect 225 313 226 314 
<< m1 >>
rect 226 313 227 314 
<< m1 >>
rect 227 313 228 314 
<< m1 >>
rect 228 313 229 314 
<< m1 >>
rect 229 313 230 314 
<< m1 >>
rect 230 313 231 314 
<< m1 >>
rect 231 313 232 314 
<< m1 >>
rect 232 313 233 314 
<< m1 >>
rect 239 313 240 314 
<< m1 >>
rect 253 313 254 314 
<< m1 >>
rect 255 313 256 314 
<< m1 >>
rect 256 313 257 314 
<< m1 >>
rect 257 313 258 314 
<< m1 >>
rect 258 313 259 314 
<< m1 >>
rect 259 313 260 314 
<< m1 >>
rect 260 313 261 314 
<< m1 >>
rect 261 313 262 314 
<< m1 >>
rect 262 313 263 314 
<< m1 >>
rect 263 313 264 314 
<< m1 >>
rect 264 313 265 314 
<< m1 >>
rect 265 313 266 314 
<< m1 >>
rect 266 313 267 314 
<< m2 >>
rect 266 313 267 314 
<< m1 >>
rect 267 313 268 314 
<< m1 >>
rect 268 313 269 314 
<< m1 >>
rect 269 313 270 314 
<< m2 >>
rect 269 313 270 314 
<< m2c >>
rect 269 313 270 314 
<< m1 >>
rect 269 313 270 314 
<< m2 >>
rect 269 313 270 314 
<< m2 >>
rect 270 313 271 314 
<< m1 >>
rect 271 313 272 314 
<< m2 >>
rect 271 313 272 314 
<< m2 >>
rect 272 313 273 314 
<< m1 >>
rect 273 313 274 314 
<< m2 >>
rect 273 313 274 314 
<< m2c >>
rect 273 313 274 314 
<< m1 >>
rect 273 313 274 314 
<< m2 >>
rect 273 313 274 314 
<< m1 >>
rect 275 313 276 314 
<< m1 >>
rect 307 313 308 314 
<< m1 >>
rect 308 313 309 314 
<< m1 >>
rect 309 313 310 314 
<< m1 >>
rect 310 313 311 314 
<< m1 >>
rect 311 313 312 314 
<< m1 >>
rect 312 313 313 314 
<< m1 >>
rect 313 313 314 314 
<< m1 >>
rect 314 313 315 314 
<< m1 >>
rect 315 313 316 314 
<< m1 >>
rect 316 313 317 314 
<< m1 >>
rect 317 313 318 314 
<< m1 >>
rect 318 313 319 314 
<< m1 >>
rect 319 313 320 314 
<< m1 >>
rect 320 313 321 314 
<< m1 >>
rect 321 313 322 314 
<< m1 >>
rect 322 313 323 314 
<< m1 >>
rect 323 313 324 314 
<< m2 >>
rect 323 313 324 314 
<< m2c >>
rect 323 313 324 314 
<< m1 >>
rect 323 313 324 314 
<< m2 >>
rect 323 313 324 314 
<< m2 >>
rect 324 313 325 314 
<< m1 >>
rect 325 313 326 314 
<< m2 >>
rect 325 313 326 314 
<< m2 >>
rect 326 313 327 314 
<< m1 >>
rect 327 313 328 314 
<< m2 >>
rect 327 313 328 314 
<< m2 >>
rect 328 313 329 314 
<< m1 >>
rect 329 313 330 314 
<< m2 >>
rect 329 313 330 314 
<< m2c >>
rect 329 313 330 314 
<< m1 >>
rect 329 313 330 314 
<< m2 >>
rect 329 313 330 314 
<< m1 >>
rect 331 313 332 314 
<< m1 >>
rect 334 313 335 314 
<< m2 >>
rect 335 313 336 314 
<< m1 >>
rect 336 313 337 314 
<< m2 >>
rect 336 313 337 314 
<< m2c >>
rect 336 313 337 314 
<< m1 >>
rect 336 313 337 314 
<< m2 >>
rect 336 313 337 314 
<< m1 >>
rect 337 313 338 314 
<< m1 >>
rect 338 313 339 314 
<< m1 >>
rect 339 313 340 314 
<< m1 >>
rect 340 313 341 314 
<< m1 >>
rect 341 313 342 314 
<< m1 >>
rect 342 313 343 314 
<< m1 >>
rect 343 313 344 314 
<< m1 >>
rect 10 314 11 315 
<< m1 >>
rect 28 314 29 315 
<< m1 >>
rect 37 314 38 315 
<< m2 >>
rect 38 314 39 315 
<< m1 >>
rect 46 314 47 315 
<< m1 >>
rect 49 314 50 315 
<< m2 >>
rect 55 314 56 315 
<< m2 >>
rect 57 314 58 315 
<< m2 >>
rect 60 314 61 315 
<< m2 >>
rect 62 314 63 315 
<< m2 >>
rect 64 314 65 315 
<< m2 >>
rect 73 314 74 315 
<< m2 >>
rect 75 314 76 315 
<< m1 >>
rect 82 314 83 315 
<< m2 >>
rect 172 314 173 315 
<< m2 >>
rect 199 314 200 315 
<< m2 >>
rect 200 314 201 315 
<< m2 >>
rect 201 314 202 315 
<< m2 >>
rect 202 314 203 315 
<< m2 >>
rect 203 314 204 315 
<< m2 >>
rect 204 314 205 315 
<< m2 >>
rect 205 314 206 315 
<< m2 >>
rect 206 314 207 315 
<< m2 >>
rect 207 314 208 315 
<< m2 >>
rect 211 314 212 315 
<< m2 >>
rect 214 314 215 315 
<< m2 >>
rect 217 314 218 315 
<< m2 >>
rect 219 314 220 315 
<< m2 >>
rect 223 314 224 315 
<< m1 >>
rect 232 314 233 315 
<< m1 >>
rect 239 314 240 315 
<< m1 >>
rect 253 314 254 315 
<< m1 >>
rect 255 314 256 315 
<< m2 >>
rect 266 314 267 315 
<< m1 >>
rect 271 314 272 315 
<< m1 >>
rect 275 314 276 315 
<< m1 >>
rect 307 314 308 315 
<< m1 >>
rect 325 314 326 315 
<< m1 >>
rect 327 314 328 315 
<< m1 >>
rect 329 314 330 315 
<< m1 >>
rect 331 314 332 315 
<< m1 >>
rect 334 314 335 315 
<< m1 >>
rect 343 314 344 315 
<< m1 >>
rect 10 315 11 316 
<< m1 >>
rect 28 315 29 316 
<< m1 >>
rect 37 315 38 316 
<< m2 >>
rect 38 315 39 316 
<< m1 >>
rect 46 315 47 316 
<< m1 >>
rect 49 315 50 316 
<< m1 >>
rect 55 315 56 316 
<< m2 >>
rect 55 315 56 316 
<< m2c >>
rect 55 315 56 316 
<< m1 >>
rect 55 315 56 316 
<< m2 >>
rect 55 315 56 316 
<< m1 >>
rect 57 315 58 316 
<< m2 >>
rect 57 315 58 316 
<< m2c >>
rect 57 315 58 316 
<< m1 >>
rect 57 315 58 316 
<< m2 >>
rect 57 315 58 316 
<< m1 >>
rect 60 315 61 316 
<< m2 >>
rect 60 315 61 316 
<< m2c >>
rect 60 315 61 316 
<< m1 >>
rect 60 315 61 316 
<< m2 >>
rect 60 315 61 316 
<< m1 >>
rect 62 315 63 316 
<< m2 >>
rect 62 315 63 316 
<< m2c >>
rect 62 315 63 316 
<< m1 >>
rect 62 315 63 316 
<< m2 >>
rect 62 315 63 316 
<< m1 >>
rect 64 315 65 316 
<< m2 >>
rect 64 315 65 316 
<< m2c >>
rect 64 315 65 316 
<< m1 >>
rect 64 315 65 316 
<< m2 >>
rect 64 315 65 316 
<< m1 >>
rect 73 315 74 316 
<< m2 >>
rect 73 315 74 316 
<< m2c >>
rect 73 315 74 316 
<< m1 >>
rect 73 315 74 316 
<< m2 >>
rect 73 315 74 316 
<< m1 >>
rect 75 315 76 316 
<< m2 >>
rect 75 315 76 316 
<< m2c >>
rect 75 315 76 316 
<< m1 >>
rect 75 315 76 316 
<< m2 >>
rect 75 315 76 316 
<< m1 >>
rect 82 315 83 316 
<< m1 >>
rect 85 315 86 316 
<< m1 >>
rect 86 315 87 316 
<< m1 >>
rect 87 315 88 316 
<< m1 >>
rect 88 315 89 316 
<< m1 >>
rect 89 315 90 316 
<< m1 >>
rect 90 315 91 316 
<< m1 >>
rect 91 315 92 316 
<< m1 >>
rect 92 315 93 316 
<< m1 >>
rect 93 315 94 316 
<< m1 >>
rect 94 315 95 316 
<< m1 >>
rect 95 315 96 316 
<< m1 >>
rect 96 315 97 316 
<< m1 >>
rect 97 315 98 316 
<< m1 >>
rect 98 315 99 316 
<< m1 >>
rect 99 315 100 316 
<< m1 >>
rect 100 315 101 316 
<< m1 >>
rect 172 315 173 316 
<< m2 >>
rect 172 315 173 316 
<< m2c >>
rect 172 315 173 316 
<< m1 >>
rect 172 315 173 316 
<< m2 >>
rect 172 315 173 316 
<< m1 >>
rect 199 315 200 316 
<< m2 >>
rect 199 315 200 316 
<< m2c >>
rect 199 315 200 316 
<< m1 >>
rect 199 315 200 316 
<< m2 >>
rect 199 315 200 316 
<< m1 >>
rect 211 315 212 316 
<< m2 >>
rect 211 315 212 316 
<< m2c >>
rect 211 315 212 316 
<< m1 >>
rect 211 315 212 316 
<< m2 >>
rect 211 315 212 316 
<< m1 >>
rect 214 315 215 316 
<< m2 >>
rect 214 315 215 316 
<< m2c >>
rect 214 315 215 316 
<< m1 >>
rect 214 315 215 316 
<< m2 >>
rect 214 315 215 316 
<< m1 >>
rect 215 315 216 316 
<< m1 >>
rect 216 315 217 316 
<< m1 >>
rect 217 315 218 316 
<< m2 >>
rect 217 315 218 316 
<< m1 >>
rect 219 315 220 316 
<< m2 >>
rect 219 315 220 316 
<< m2c >>
rect 219 315 220 316 
<< m1 >>
rect 219 315 220 316 
<< m2 >>
rect 219 315 220 316 
<< m1 >>
rect 223 315 224 316 
<< m2 >>
rect 223 315 224 316 
<< m2c >>
rect 223 315 224 316 
<< m1 >>
rect 223 315 224 316 
<< m2 >>
rect 223 315 224 316 
<< m1 >>
rect 232 315 233 316 
<< m1 >>
rect 239 315 240 316 
<< m1 >>
rect 253 315 254 316 
<< m1 >>
rect 255 315 256 316 
<< m1 >>
rect 266 315 267 316 
<< m2 >>
rect 266 315 267 316 
<< m2c >>
rect 266 315 267 316 
<< m1 >>
rect 266 315 267 316 
<< m2 >>
rect 266 315 267 316 
<< m1 >>
rect 267 315 268 316 
<< m1 >>
rect 268 315 269 316 
<< m1 >>
rect 269 315 270 316 
<< m2 >>
rect 269 315 270 316 
<< m2c >>
rect 269 315 270 316 
<< m1 >>
rect 269 315 270 316 
<< m2 >>
rect 269 315 270 316 
<< m2 >>
rect 270 315 271 316 
<< m1 >>
rect 271 315 272 316 
<< m2 >>
rect 271 315 272 316 
<< m2 >>
rect 272 315 273 316 
<< m1 >>
rect 273 315 274 316 
<< m2 >>
rect 273 315 274 316 
<< m2c >>
rect 273 315 274 316 
<< m1 >>
rect 273 315 274 316 
<< m2 >>
rect 273 315 274 316 
<< m2 >>
rect 274 315 275 316 
<< m1 >>
rect 275 315 276 316 
<< m2 >>
rect 275 315 276 316 
<< m1 >>
rect 307 315 308 316 
<< m1 >>
rect 325 315 326 316 
<< m1 >>
rect 327 315 328 316 
<< m1 >>
rect 329 315 330 316 
<< m1 >>
rect 331 315 332 316 
<< m1 >>
rect 334 315 335 316 
<< m1 >>
rect 343 315 344 316 
<< m1 >>
rect 10 316 11 317 
<< m1 >>
rect 28 316 29 317 
<< m1 >>
rect 37 316 38 317 
<< m2 >>
rect 38 316 39 317 
<< m1 >>
rect 46 316 47 317 
<< m1 >>
rect 49 316 50 317 
<< m1 >>
rect 55 316 56 317 
<< m1 >>
rect 57 316 58 317 
<< m1 >>
rect 60 316 61 317 
<< m1 >>
rect 62 316 63 317 
<< m1 >>
rect 64 316 65 317 
<< m1 >>
rect 73 316 74 317 
<< m1 >>
rect 75 316 76 317 
<< m1 >>
rect 82 316 83 317 
<< m1 >>
rect 85 316 86 317 
<< m2 >>
rect 91 316 92 317 
<< m2 >>
rect 92 316 93 317 
<< m2 >>
rect 93 316 94 317 
<< m2 >>
rect 94 316 95 317 
<< m2 >>
rect 95 316 96 317 
<< m2 >>
rect 96 316 97 317 
<< m2 >>
rect 97 316 98 317 
<< m2 >>
rect 98 316 99 317 
<< m2 >>
rect 99 316 100 317 
<< m1 >>
rect 100 316 101 317 
<< m2 >>
rect 100 316 101 317 
<< m2 >>
rect 101 316 102 317 
<< m1 >>
rect 102 316 103 317 
<< m2 >>
rect 102 316 103 317 
<< m2c >>
rect 102 316 103 317 
<< m1 >>
rect 102 316 103 317 
<< m2 >>
rect 102 316 103 317 
<< m1 >>
rect 103 316 104 317 
<< m1 >>
rect 172 316 173 317 
<< m1 >>
rect 199 316 200 317 
<< m1 >>
rect 211 316 212 317 
<< m1 >>
rect 217 316 218 317 
<< m2 >>
rect 217 316 218 317 
<< m1 >>
rect 219 316 220 317 
<< m1 >>
rect 223 316 224 317 
<< m1 >>
rect 232 316 233 317 
<< m1 >>
rect 239 316 240 317 
<< m1 >>
rect 253 316 254 317 
<< m1 >>
rect 255 316 256 317 
<< m1 >>
rect 271 316 272 317 
<< m1 >>
rect 275 316 276 317 
<< m2 >>
rect 275 316 276 317 
<< m1 >>
rect 307 316 308 317 
<< m1 >>
rect 325 316 326 317 
<< m1 >>
rect 327 316 328 317 
<< m1 >>
rect 329 316 330 317 
<< m1 >>
rect 331 316 332 317 
<< m1 >>
rect 334 316 335 317 
<< m1 >>
rect 343 316 344 317 
<< m1 >>
rect 10 317 11 318 
<< m1 >>
rect 28 317 29 318 
<< m1 >>
rect 37 317 38 318 
<< m2 >>
rect 38 317 39 318 
<< m1 >>
rect 46 317 47 318 
<< m1 >>
rect 49 317 50 318 
<< m1 >>
rect 55 317 56 318 
<< m1 >>
rect 57 317 58 318 
<< m1 >>
rect 60 317 61 318 
<< m1 >>
rect 62 317 63 318 
<< m1 >>
rect 64 317 65 318 
<< m1 >>
rect 73 317 74 318 
<< m1 >>
rect 75 317 76 318 
<< m1 >>
rect 82 317 83 318 
<< m1 >>
rect 85 317 86 318 
<< m1 >>
rect 91 317 92 318 
<< m2 >>
rect 91 317 92 318 
<< m2c >>
rect 91 317 92 318 
<< m1 >>
rect 91 317 92 318 
<< m2 >>
rect 91 317 92 318 
<< m1 >>
rect 100 317 101 318 
<< m1 >>
rect 103 317 104 318 
<< m1 >>
rect 172 317 173 318 
<< m1 >>
rect 199 317 200 318 
<< m1 >>
rect 211 317 212 318 
<< m1 >>
rect 217 317 218 318 
<< m2 >>
rect 217 317 218 318 
<< m1 >>
rect 219 317 220 318 
<< m1 >>
rect 223 317 224 318 
<< m1 >>
rect 232 317 233 318 
<< m1 >>
rect 239 317 240 318 
<< m1 >>
rect 253 317 254 318 
<< m1 >>
rect 255 317 256 318 
<< m1 >>
rect 271 317 272 318 
<< m1 >>
rect 275 317 276 318 
<< m2 >>
rect 275 317 276 318 
<< m1 >>
rect 307 317 308 318 
<< m1 >>
rect 325 317 326 318 
<< m1 >>
rect 327 317 328 318 
<< m1 >>
rect 329 317 330 318 
<< m1 >>
rect 331 317 332 318 
<< m1 >>
rect 334 317 335 318 
<< m1 >>
rect 343 317 344 318 
<< m1 >>
rect 10 318 11 319 
<< pdiffusion >>
rect 12 318 13 319 
<< pdiffusion >>
rect 13 318 14 319 
<< pdiffusion >>
rect 14 318 15 319 
<< pdiffusion >>
rect 15 318 16 319 
<< pdiffusion >>
rect 16 318 17 319 
<< pdiffusion >>
rect 17 318 18 319 
<< m1 >>
rect 28 318 29 319 
<< pdiffusion >>
rect 30 318 31 319 
<< pdiffusion >>
rect 31 318 32 319 
<< pdiffusion >>
rect 32 318 33 319 
<< pdiffusion >>
rect 33 318 34 319 
<< pdiffusion >>
rect 34 318 35 319 
<< pdiffusion >>
rect 35 318 36 319 
<< m1 >>
rect 37 318 38 319 
<< m2 >>
rect 38 318 39 319 
<< m1 >>
rect 46 318 47 319 
<< pdiffusion >>
rect 48 318 49 319 
<< m1 >>
rect 49 318 50 319 
<< pdiffusion >>
rect 49 318 50 319 
<< pdiffusion >>
rect 50 318 51 319 
<< pdiffusion >>
rect 51 318 52 319 
<< pdiffusion >>
rect 52 318 53 319 
<< pdiffusion >>
rect 53 318 54 319 
<< m1 >>
rect 55 318 56 319 
<< m1 >>
rect 57 318 58 319 
<< m1 >>
rect 60 318 61 319 
<< m1 >>
rect 62 318 63 319 
<< m1 >>
rect 64 318 65 319 
<< pdiffusion >>
rect 66 318 67 319 
<< pdiffusion >>
rect 67 318 68 319 
<< pdiffusion >>
rect 68 318 69 319 
<< pdiffusion >>
rect 69 318 70 319 
<< pdiffusion >>
rect 70 318 71 319 
<< pdiffusion >>
rect 71 318 72 319 
<< m1 >>
rect 73 318 74 319 
<< m1 >>
rect 75 318 76 319 
<< m1 >>
rect 82 318 83 319 
<< pdiffusion >>
rect 84 318 85 319 
<< m1 >>
rect 85 318 86 319 
<< pdiffusion >>
rect 85 318 86 319 
<< pdiffusion >>
rect 86 318 87 319 
<< pdiffusion >>
rect 87 318 88 319 
<< pdiffusion >>
rect 88 318 89 319 
<< pdiffusion >>
rect 89 318 90 319 
<< m1 >>
rect 91 318 92 319 
<< m1 >>
rect 100 318 101 319 
<< pdiffusion >>
rect 102 318 103 319 
<< m1 >>
rect 103 318 104 319 
<< pdiffusion >>
rect 103 318 104 319 
<< pdiffusion >>
rect 104 318 105 319 
<< pdiffusion >>
rect 105 318 106 319 
<< pdiffusion >>
rect 106 318 107 319 
<< pdiffusion >>
rect 107 318 108 319 
<< pdiffusion >>
rect 120 318 121 319 
<< pdiffusion >>
rect 121 318 122 319 
<< pdiffusion >>
rect 122 318 123 319 
<< pdiffusion >>
rect 123 318 124 319 
<< pdiffusion >>
rect 124 318 125 319 
<< pdiffusion >>
rect 125 318 126 319 
<< pdiffusion >>
rect 138 318 139 319 
<< pdiffusion >>
rect 139 318 140 319 
<< pdiffusion >>
rect 140 318 141 319 
<< pdiffusion >>
rect 141 318 142 319 
<< pdiffusion >>
rect 142 318 143 319 
<< pdiffusion >>
rect 143 318 144 319 
<< pdiffusion >>
rect 156 318 157 319 
<< pdiffusion >>
rect 157 318 158 319 
<< pdiffusion >>
rect 158 318 159 319 
<< pdiffusion >>
rect 159 318 160 319 
<< pdiffusion >>
rect 160 318 161 319 
<< pdiffusion >>
rect 161 318 162 319 
<< m1 >>
rect 172 318 173 319 
<< pdiffusion >>
rect 174 318 175 319 
<< pdiffusion >>
rect 175 318 176 319 
<< pdiffusion >>
rect 176 318 177 319 
<< pdiffusion >>
rect 177 318 178 319 
<< pdiffusion >>
rect 178 318 179 319 
<< pdiffusion >>
rect 179 318 180 319 
<< pdiffusion >>
rect 192 318 193 319 
<< pdiffusion >>
rect 193 318 194 319 
<< pdiffusion >>
rect 194 318 195 319 
<< pdiffusion >>
rect 195 318 196 319 
<< pdiffusion >>
rect 196 318 197 319 
<< pdiffusion >>
rect 197 318 198 319 
<< m1 >>
rect 199 318 200 319 
<< pdiffusion >>
rect 210 318 211 319 
<< m1 >>
rect 211 318 212 319 
<< pdiffusion >>
rect 211 318 212 319 
<< pdiffusion >>
rect 212 318 213 319 
<< pdiffusion >>
rect 213 318 214 319 
<< pdiffusion >>
rect 214 318 215 319 
<< pdiffusion >>
rect 215 318 216 319 
<< m1 >>
rect 217 318 218 319 
<< m2 >>
rect 217 318 218 319 
<< m1 >>
rect 219 318 220 319 
<< m1 >>
rect 223 318 224 319 
<< pdiffusion >>
rect 228 318 229 319 
<< pdiffusion >>
rect 229 318 230 319 
<< pdiffusion >>
rect 230 318 231 319 
<< pdiffusion >>
rect 231 318 232 319 
<< m1 >>
rect 232 318 233 319 
<< pdiffusion >>
rect 232 318 233 319 
<< pdiffusion >>
rect 233 318 234 319 
<< m1 >>
rect 239 318 240 319 
<< pdiffusion >>
rect 246 318 247 319 
<< pdiffusion >>
rect 247 318 248 319 
<< pdiffusion >>
rect 248 318 249 319 
<< pdiffusion >>
rect 249 318 250 319 
<< pdiffusion >>
rect 250 318 251 319 
<< pdiffusion >>
rect 251 318 252 319 
<< m1 >>
rect 253 318 254 319 
<< m1 >>
rect 255 318 256 319 
<< pdiffusion >>
rect 264 318 265 319 
<< pdiffusion >>
rect 265 318 266 319 
<< pdiffusion >>
rect 266 318 267 319 
<< pdiffusion >>
rect 267 318 268 319 
<< pdiffusion >>
rect 268 318 269 319 
<< pdiffusion >>
rect 269 318 270 319 
<< m1 >>
rect 271 318 272 319 
<< m1 >>
rect 275 318 276 319 
<< m2 >>
rect 275 318 276 319 
<< pdiffusion >>
rect 282 318 283 319 
<< pdiffusion >>
rect 283 318 284 319 
<< pdiffusion >>
rect 284 318 285 319 
<< pdiffusion >>
rect 285 318 286 319 
<< pdiffusion >>
rect 286 318 287 319 
<< pdiffusion >>
rect 287 318 288 319 
<< pdiffusion >>
rect 300 318 301 319 
<< pdiffusion >>
rect 301 318 302 319 
<< pdiffusion >>
rect 302 318 303 319 
<< pdiffusion >>
rect 303 318 304 319 
<< pdiffusion >>
rect 304 318 305 319 
<< pdiffusion >>
rect 305 318 306 319 
<< m1 >>
rect 307 318 308 319 
<< pdiffusion >>
rect 318 318 319 319 
<< pdiffusion >>
rect 319 318 320 319 
<< pdiffusion >>
rect 320 318 321 319 
<< pdiffusion >>
rect 321 318 322 319 
<< pdiffusion >>
rect 322 318 323 319 
<< pdiffusion >>
rect 323 318 324 319 
<< m1 >>
rect 325 318 326 319 
<< m1 >>
rect 327 318 328 319 
<< m1 >>
rect 329 318 330 319 
<< m1 >>
rect 331 318 332 319 
<< m1 >>
rect 334 318 335 319 
<< pdiffusion >>
rect 336 318 337 319 
<< pdiffusion >>
rect 337 318 338 319 
<< pdiffusion >>
rect 338 318 339 319 
<< pdiffusion >>
rect 339 318 340 319 
<< pdiffusion >>
rect 340 318 341 319 
<< pdiffusion >>
rect 341 318 342 319 
<< m1 >>
rect 343 318 344 319 
<< m1 >>
rect 10 319 11 320 
<< pdiffusion >>
rect 12 319 13 320 
<< pdiffusion >>
rect 13 319 14 320 
<< pdiffusion >>
rect 14 319 15 320 
<< pdiffusion >>
rect 15 319 16 320 
<< pdiffusion >>
rect 16 319 17 320 
<< pdiffusion >>
rect 17 319 18 320 
<< m1 >>
rect 28 319 29 320 
<< pdiffusion >>
rect 30 319 31 320 
<< pdiffusion >>
rect 31 319 32 320 
<< pdiffusion >>
rect 32 319 33 320 
<< pdiffusion >>
rect 33 319 34 320 
<< pdiffusion >>
rect 34 319 35 320 
<< pdiffusion >>
rect 35 319 36 320 
<< m1 >>
rect 37 319 38 320 
<< m2 >>
rect 38 319 39 320 
<< m1 >>
rect 46 319 47 320 
<< pdiffusion >>
rect 48 319 49 320 
<< pdiffusion >>
rect 49 319 50 320 
<< pdiffusion >>
rect 50 319 51 320 
<< pdiffusion >>
rect 51 319 52 320 
<< pdiffusion >>
rect 52 319 53 320 
<< pdiffusion >>
rect 53 319 54 320 
<< m1 >>
rect 55 319 56 320 
<< m1 >>
rect 57 319 58 320 
<< m1 >>
rect 60 319 61 320 
<< m1 >>
rect 62 319 63 320 
<< m1 >>
rect 64 319 65 320 
<< pdiffusion >>
rect 66 319 67 320 
<< pdiffusion >>
rect 67 319 68 320 
<< pdiffusion >>
rect 68 319 69 320 
<< pdiffusion >>
rect 69 319 70 320 
<< pdiffusion >>
rect 70 319 71 320 
<< pdiffusion >>
rect 71 319 72 320 
<< m1 >>
rect 73 319 74 320 
<< m1 >>
rect 75 319 76 320 
<< m1 >>
rect 82 319 83 320 
<< pdiffusion >>
rect 84 319 85 320 
<< pdiffusion >>
rect 85 319 86 320 
<< pdiffusion >>
rect 86 319 87 320 
<< pdiffusion >>
rect 87 319 88 320 
<< pdiffusion >>
rect 88 319 89 320 
<< pdiffusion >>
rect 89 319 90 320 
<< m1 >>
rect 91 319 92 320 
<< m1 >>
rect 100 319 101 320 
<< pdiffusion >>
rect 102 319 103 320 
<< pdiffusion >>
rect 103 319 104 320 
<< pdiffusion >>
rect 104 319 105 320 
<< pdiffusion >>
rect 105 319 106 320 
<< pdiffusion >>
rect 106 319 107 320 
<< pdiffusion >>
rect 107 319 108 320 
<< pdiffusion >>
rect 120 319 121 320 
<< pdiffusion >>
rect 121 319 122 320 
<< pdiffusion >>
rect 122 319 123 320 
<< pdiffusion >>
rect 123 319 124 320 
<< pdiffusion >>
rect 124 319 125 320 
<< pdiffusion >>
rect 125 319 126 320 
<< pdiffusion >>
rect 138 319 139 320 
<< pdiffusion >>
rect 139 319 140 320 
<< pdiffusion >>
rect 140 319 141 320 
<< pdiffusion >>
rect 141 319 142 320 
<< pdiffusion >>
rect 142 319 143 320 
<< pdiffusion >>
rect 143 319 144 320 
<< pdiffusion >>
rect 156 319 157 320 
<< pdiffusion >>
rect 157 319 158 320 
<< pdiffusion >>
rect 158 319 159 320 
<< pdiffusion >>
rect 159 319 160 320 
<< pdiffusion >>
rect 160 319 161 320 
<< pdiffusion >>
rect 161 319 162 320 
<< m1 >>
rect 172 319 173 320 
<< pdiffusion >>
rect 174 319 175 320 
<< pdiffusion >>
rect 175 319 176 320 
<< pdiffusion >>
rect 176 319 177 320 
<< pdiffusion >>
rect 177 319 178 320 
<< pdiffusion >>
rect 178 319 179 320 
<< pdiffusion >>
rect 179 319 180 320 
<< pdiffusion >>
rect 192 319 193 320 
<< pdiffusion >>
rect 193 319 194 320 
<< pdiffusion >>
rect 194 319 195 320 
<< pdiffusion >>
rect 195 319 196 320 
<< pdiffusion >>
rect 196 319 197 320 
<< pdiffusion >>
rect 197 319 198 320 
<< m1 >>
rect 199 319 200 320 
<< pdiffusion >>
rect 210 319 211 320 
<< pdiffusion >>
rect 211 319 212 320 
<< pdiffusion >>
rect 212 319 213 320 
<< pdiffusion >>
rect 213 319 214 320 
<< pdiffusion >>
rect 214 319 215 320 
<< pdiffusion >>
rect 215 319 216 320 
<< m1 >>
rect 217 319 218 320 
<< m2 >>
rect 217 319 218 320 
<< m1 >>
rect 219 319 220 320 
<< m1 >>
rect 223 319 224 320 
<< pdiffusion >>
rect 228 319 229 320 
<< pdiffusion >>
rect 229 319 230 320 
<< pdiffusion >>
rect 230 319 231 320 
<< pdiffusion >>
rect 231 319 232 320 
<< pdiffusion >>
rect 232 319 233 320 
<< pdiffusion >>
rect 233 319 234 320 
<< m1 >>
rect 239 319 240 320 
<< pdiffusion >>
rect 246 319 247 320 
<< pdiffusion >>
rect 247 319 248 320 
<< pdiffusion >>
rect 248 319 249 320 
<< pdiffusion >>
rect 249 319 250 320 
<< pdiffusion >>
rect 250 319 251 320 
<< pdiffusion >>
rect 251 319 252 320 
<< m1 >>
rect 253 319 254 320 
<< m1 >>
rect 255 319 256 320 
<< pdiffusion >>
rect 264 319 265 320 
<< pdiffusion >>
rect 265 319 266 320 
<< pdiffusion >>
rect 266 319 267 320 
<< pdiffusion >>
rect 267 319 268 320 
<< pdiffusion >>
rect 268 319 269 320 
<< pdiffusion >>
rect 269 319 270 320 
<< m1 >>
rect 271 319 272 320 
<< m1 >>
rect 275 319 276 320 
<< m2 >>
rect 275 319 276 320 
<< pdiffusion >>
rect 282 319 283 320 
<< pdiffusion >>
rect 283 319 284 320 
<< pdiffusion >>
rect 284 319 285 320 
<< pdiffusion >>
rect 285 319 286 320 
<< pdiffusion >>
rect 286 319 287 320 
<< pdiffusion >>
rect 287 319 288 320 
<< pdiffusion >>
rect 300 319 301 320 
<< pdiffusion >>
rect 301 319 302 320 
<< pdiffusion >>
rect 302 319 303 320 
<< pdiffusion >>
rect 303 319 304 320 
<< pdiffusion >>
rect 304 319 305 320 
<< pdiffusion >>
rect 305 319 306 320 
<< m1 >>
rect 307 319 308 320 
<< pdiffusion >>
rect 318 319 319 320 
<< pdiffusion >>
rect 319 319 320 320 
<< pdiffusion >>
rect 320 319 321 320 
<< pdiffusion >>
rect 321 319 322 320 
<< pdiffusion >>
rect 322 319 323 320 
<< pdiffusion >>
rect 323 319 324 320 
<< m1 >>
rect 325 319 326 320 
<< m1 >>
rect 327 319 328 320 
<< m1 >>
rect 329 319 330 320 
<< m1 >>
rect 331 319 332 320 
<< m1 >>
rect 334 319 335 320 
<< pdiffusion >>
rect 336 319 337 320 
<< pdiffusion >>
rect 337 319 338 320 
<< pdiffusion >>
rect 338 319 339 320 
<< pdiffusion >>
rect 339 319 340 320 
<< pdiffusion >>
rect 340 319 341 320 
<< pdiffusion >>
rect 341 319 342 320 
<< m1 >>
rect 343 319 344 320 
<< m1 >>
rect 10 320 11 321 
<< pdiffusion >>
rect 12 320 13 321 
<< pdiffusion >>
rect 13 320 14 321 
<< pdiffusion >>
rect 14 320 15 321 
<< pdiffusion >>
rect 15 320 16 321 
<< pdiffusion >>
rect 16 320 17 321 
<< pdiffusion >>
rect 17 320 18 321 
<< m1 >>
rect 28 320 29 321 
<< pdiffusion >>
rect 30 320 31 321 
<< pdiffusion >>
rect 31 320 32 321 
<< pdiffusion >>
rect 32 320 33 321 
<< pdiffusion >>
rect 33 320 34 321 
<< pdiffusion >>
rect 34 320 35 321 
<< pdiffusion >>
rect 35 320 36 321 
<< m1 >>
rect 37 320 38 321 
<< m2 >>
rect 38 320 39 321 
<< m1 >>
rect 46 320 47 321 
<< pdiffusion >>
rect 48 320 49 321 
<< pdiffusion >>
rect 49 320 50 321 
<< pdiffusion >>
rect 50 320 51 321 
<< pdiffusion >>
rect 51 320 52 321 
<< pdiffusion >>
rect 52 320 53 321 
<< pdiffusion >>
rect 53 320 54 321 
<< m1 >>
rect 55 320 56 321 
<< m1 >>
rect 57 320 58 321 
<< m1 >>
rect 60 320 61 321 
<< m1 >>
rect 62 320 63 321 
<< m1 >>
rect 64 320 65 321 
<< pdiffusion >>
rect 66 320 67 321 
<< pdiffusion >>
rect 67 320 68 321 
<< pdiffusion >>
rect 68 320 69 321 
<< pdiffusion >>
rect 69 320 70 321 
<< pdiffusion >>
rect 70 320 71 321 
<< pdiffusion >>
rect 71 320 72 321 
<< m1 >>
rect 73 320 74 321 
<< m1 >>
rect 75 320 76 321 
<< m1 >>
rect 82 320 83 321 
<< pdiffusion >>
rect 84 320 85 321 
<< pdiffusion >>
rect 85 320 86 321 
<< pdiffusion >>
rect 86 320 87 321 
<< pdiffusion >>
rect 87 320 88 321 
<< pdiffusion >>
rect 88 320 89 321 
<< pdiffusion >>
rect 89 320 90 321 
<< m1 >>
rect 91 320 92 321 
<< m1 >>
rect 100 320 101 321 
<< pdiffusion >>
rect 102 320 103 321 
<< pdiffusion >>
rect 103 320 104 321 
<< pdiffusion >>
rect 104 320 105 321 
<< pdiffusion >>
rect 105 320 106 321 
<< pdiffusion >>
rect 106 320 107 321 
<< pdiffusion >>
rect 107 320 108 321 
<< pdiffusion >>
rect 120 320 121 321 
<< pdiffusion >>
rect 121 320 122 321 
<< pdiffusion >>
rect 122 320 123 321 
<< pdiffusion >>
rect 123 320 124 321 
<< pdiffusion >>
rect 124 320 125 321 
<< pdiffusion >>
rect 125 320 126 321 
<< pdiffusion >>
rect 138 320 139 321 
<< pdiffusion >>
rect 139 320 140 321 
<< pdiffusion >>
rect 140 320 141 321 
<< pdiffusion >>
rect 141 320 142 321 
<< pdiffusion >>
rect 142 320 143 321 
<< pdiffusion >>
rect 143 320 144 321 
<< pdiffusion >>
rect 156 320 157 321 
<< pdiffusion >>
rect 157 320 158 321 
<< pdiffusion >>
rect 158 320 159 321 
<< pdiffusion >>
rect 159 320 160 321 
<< pdiffusion >>
rect 160 320 161 321 
<< pdiffusion >>
rect 161 320 162 321 
<< m1 >>
rect 172 320 173 321 
<< pdiffusion >>
rect 174 320 175 321 
<< pdiffusion >>
rect 175 320 176 321 
<< pdiffusion >>
rect 176 320 177 321 
<< pdiffusion >>
rect 177 320 178 321 
<< pdiffusion >>
rect 178 320 179 321 
<< pdiffusion >>
rect 179 320 180 321 
<< pdiffusion >>
rect 192 320 193 321 
<< pdiffusion >>
rect 193 320 194 321 
<< pdiffusion >>
rect 194 320 195 321 
<< pdiffusion >>
rect 195 320 196 321 
<< pdiffusion >>
rect 196 320 197 321 
<< pdiffusion >>
rect 197 320 198 321 
<< m1 >>
rect 199 320 200 321 
<< pdiffusion >>
rect 210 320 211 321 
<< pdiffusion >>
rect 211 320 212 321 
<< pdiffusion >>
rect 212 320 213 321 
<< pdiffusion >>
rect 213 320 214 321 
<< pdiffusion >>
rect 214 320 215 321 
<< pdiffusion >>
rect 215 320 216 321 
<< m1 >>
rect 217 320 218 321 
<< m2 >>
rect 217 320 218 321 
<< m1 >>
rect 219 320 220 321 
<< m1 >>
rect 223 320 224 321 
<< pdiffusion >>
rect 228 320 229 321 
<< pdiffusion >>
rect 229 320 230 321 
<< pdiffusion >>
rect 230 320 231 321 
<< pdiffusion >>
rect 231 320 232 321 
<< pdiffusion >>
rect 232 320 233 321 
<< pdiffusion >>
rect 233 320 234 321 
<< m1 >>
rect 239 320 240 321 
<< pdiffusion >>
rect 246 320 247 321 
<< pdiffusion >>
rect 247 320 248 321 
<< pdiffusion >>
rect 248 320 249 321 
<< pdiffusion >>
rect 249 320 250 321 
<< pdiffusion >>
rect 250 320 251 321 
<< pdiffusion >>
rect 251 320 252 321 
<< m1 >>
rect 253 320 254 321 
<< m1 >>
rect 255 320 256 321 
<< pdiffusion >>
rect 264 320 265 321 
<< pdiffusion >>
rect 265 320 266 321 
<< pdiffusion >>
rect 266 320 267 321 
<< pdiffusion >>
rect 267 320 268 321 
<< pdiffusion >>
rect 268 320 269 321 
<< pdiffusion >>
rect 269 320 270 321 
<< m1 >>
rect 271 320 272 321 
<< m1 >>
rect 275 320 276 321 
<< m2 >>
rect 275 320 276 321 
<< pdiffusion >>
rect 282 320 283 321 
<< pdiffusion >>
rect 283 320 284 321 
<< pdiffusion >>
rect 284 320 285 321 
<< pdiffusion >>
rect 285 320 286 321 
<< pdiffusion >>
rect 286 320 287 321 
<< pdiffusion >>
rect 287 320 288 321 
<< pdiffusion >>
rect 300 320 301 321 
<< pdiffusion >>
rect 301 320 302 321 
<< pdiffusion >>
rect 302 320 303 321 
<< pdiffusion >>
rect 303 320 304 321 
<< pdiffusion >>
rect 304 320 305 321 
<< pdiffusion >>
rect 305 320 306 321 
<< m1 >>
rect 307 320 308 321 
<< pdiffusion >>
rect 318 320 319 321 
<< pdiffusion >>
rect 319 320 320 321 
<< pdiffusion >>
rect 320 320 321 321 
<< pdiffusion >>
rect 321 320 322 321 
<< pdiffusion >>
rect 322 320 323 321 
<< pdiffusion >>
rect 323 320 324 321 
<< m1 >>
rect 325 320 326 321 
<< m1 >>
rect 327 320 328 321 
<< m1 >>
rect 329 320 330 321 
<< m1 >>
rect 331 320 332 321 
<< m1 >>
rect 334 320 335 321 
<< pdiffusion >>
rect 336 320 337 321 
<< pdiffusion >>
rect 337 320 338 321 
<< pdiffusion >>
rect 338 320 339 321 
<< pdiffusion >>
rect 339 320 340 321 
<< pdiffusion >>
rect 340 320 341 321 
<< pdiffusion >>
rect 341 320 342 321 
<< m1 >>
rect 343 320 344 321 
<< m1 >>
rect 10 321 11 322 
<< pdiffusion >>
rect 12 321 13 322 
<< pdiffusion >>
rect 13 321 14 322 
<< pdiffusion >>
rect 14 321 15 322 
<< pdiffusion >>
rect 15 321 16 322 
<< pdiffusion >>
rect 16 321 17 322 
<< pdiffusion >>
rect 17 321 18 322 
<< m1 >>
rect 28 321 29 322 
<< pdiffusion >>
rect 30 321 31 322 
<< pdiffusion >>
rect 31 321 32 322 
<< pdiffusion >>
rect 32 321 33 322 
<< pdiffusion >>
rect 33 321 34 322 
<< pdiffusion >>
rect 34 321 35 322 
<< pdiffusion >>
rect 35 321 36 322 
<< m1 >>
rect 37 321 38 322 
<< m2 >>
rect 38 321 39 322 
<< m1 >>
rect 46 321 47 322 
<< pdiffusion >>
rect 48 321 49 322 
<< pdiffusion >>
rect 49 321 50 322 
<< pdiffusion >>
rect 50 321 51 322 
<< pdiffusion >>
rect 51 321 52 322 
<< pdiffusion >>
rect 52 321 53 322 
<< pdiffusion >>
rect 53 321 54 322 
<< m1 >>
rect 55 321 56 322 
<< m1 >>
rect 57 321 58 322 
<< m1 >>
rect 60 321 61 322 
<< m1 >>
rect 62 321 63 322 
<< m1 >>
rect 64 321 65 322 
<< pdiffusion >>
rect 66 321 67 322 
<< pdiffusion >>
rect 67 321 68 322 
<< pdiffusion >>
rect 68 321 69 322 
<< pdiffusion >>
rect 69 321 70 322 
<< pdiffusion >>
rect 70 321 71 322 
<< pdiffusion >>
rect 71 321 72 322 
<< m1 >>
rect 73 321 74 322 
<< m1 >>
rect 75 321 76 322 
<< m1 >>
rect 82 321 83 322 
<< pdiffusion >>
rect 84 321 85 322 
<< pdiffusion >>
rect 85 321 86 322 
<< pdiffusion >>
rect 86 321 87 322 
<< pdiffusion >>
rect 87 321 88 322 
<< pdiffusion >>
rect 88 321 89 322 
<< pdiffusion >>
rect 89 321 90 322 
<< m1 >>
rect 91 321 92 322 
<< m1 >>
rect 100 321 101 322 
<< pdiffusion >>
rect 102 321 103 322 
<< pdiffusion >>
rect 103 321 104 322 
<< pdiffusion >>
rect 104 321 105 322 
<< pdiffusion >>
rect 105 321 106 322 
<< pdiffusion >>
rect 106 321 107 322 
<< pdiffusion >>
rect 107 321 108 322 
<< pdiffusion >>
rect 120 321 121 322 
<< pdiffusion >>
rect 121 321 122 322 
<< pdiffusion >>
rect 122 321 123 322 
<< pdiffusion >>
rect 123 321 124 322 
<< pdiffusion >>
rect 124 321 125 322 
<< pdiffusion >>
rect 125 321 126 322 
<< pdiffusion >>
rect 138 321 139 322 
<< pdiffusion >>
rect 139 321 140 322 
<< pdiffusion >>
rect 140 321 141 322 
<< pdiffusion >>
rect 141 321 142 322 
<< pdiffusion >>
rect 142 321 143 322 
<< pdiffusion >>
rect 143 321 144 322 
<< pdiffusion >>
rect 156 321 157 322 
<< pdiffusion >>
rect 157 321 158 322 
<< pdiffusion >>
rect 158 321 159 322 
<< pdiffusion >>
rect 159 321 160 322 
<< pdiffusion >>
rect 160 321 161 322 
<< pdiffusion >>
rect 161 321 162 322 
<< m1 >>
rect 172 321 173 322 
<< pdiffusion >>
rect 174 321 175 322 
<< pdiffusion >>
rect 175 321 176 322 
<< pdiffusion >>
rect 176 321 177 322 
<< pdiffusion >>
rect 177 321 178 322 
<< pdiffusion >>
rect 178 321 179 322 
<< pdiffusion >>
rect 179 321 180 322 
<< pdiffusion >>
rect 192 321 193 322 
<< pdiffusion >>
rect 193 321 194 322 
<< pdiffusion >>
rect 194 321 195 322 
<< pdiffusion >>
rect 195 321 196 322 
<< pdiffusion >>
rect 196 321 197 322 
<< pdiffusion >>
rect 197 321 198 322 
<< m1 >>
rect 199 321 200 322 
<< pdiffusion >>
rect 210 321 211 322 
<< pdiffusion >>
rect 211 321 212 322 
<< pdiffusion >>
rect 212 321 213 322 
<< pdiffusion >>
rect 213 321 214 322 
<< pdiffusion >>
rect 214 321 215 322 
<< pdiffusion >>
rect 215 321 216 322 
<< m1 >>
rect 217 321 218 322 
<< m2 >>
rect 217 321 218 322 
<< m1 >>
rect 219 321 220 322 
<< m1 >>
rect 223 321 224 322 
<< pdiffusion >>
rect 228 321 229 322 
<< pdiffusion >>
rect 229 321 230 322 
<< pdiffusion >>
rect 230 321 231 322 
<< pdiffusion >>
rect 231 321 232 322 
<< pdiffusion >>
rect 232 321 233 322 
<< pdiffusion >>
rect 233 321 234 322 
<< m1 >>
rect 239 321 240 322 
<< pdiffusion >>
rect 246 321 247 322 
<< pdiffusion >>
rect 247 321 248 322 
<< pdiffusion >>
rect 248 321 249 322 
<< pdiffusion >>
rect 249 321 250 322 
<< pdiffusion >>
rect 250 321 251 322 
<< pdiffusion >>
rect 251 321 252 322 
<< m1 >>
rect 253 321 254 322 
<< m1 >>
rect 255 321 256 322 
<< pdiffusion >>
rect 264 321 265 322 
<< pdiffusion >>
rect 265 321 266 322 
<< pdiffusion >>
rect 266 321 267 322 
<< pdiffusion >>
rect 267 321 268 322 
<< pdiffusion >>
rect 268 321 269 322 
<< pdiffusion >>
rect 269 321 270 322 
<< m1 >>
rect 271 321 272 322 
<< m1 >>
rect 275 321 276 322 
<< m2 >>
rect 275 321 276 322 
<< pdiffusion >>
rect 282 321 283 322 
<< pdiffusion >>
rect 283 321 284 322 
<< pdiffusion >>
rect 284 321 285 322 
<< pdiffusion >>
rect 285 321 286 322 
<< pdiffusion >>
rect 286 321 287 322 
<< pdiffusion >>
rect 287 321 288 322 
<< pdiffusion >>
rect 300 321 301 322 
<< pdiffusion >>
rect 301 321 302 322 
<< pdiffusion >>
rect 302 321 303 322 
<< pdiffusion >>
rect 303 321 304 322 
<< pdiffusion >>
rect 304 321 305 322 
<< pdiffusion >>
rect 305 321 306 322 
<< m1 >>
rect 307 321 308 322 
<< pdiffusion >>
rect 318 321 319 322 
<< pdiffusion >>
rect 319 321 320 322 
<< pdiffusion >>
rect 320 321 321 322 
<< pdiffusion >>
rect 321 321 322 322 
<< pdiffusion >>
rect 322 321 323 322 
<< pdiffusion >>
rect 323 321 324 322 
<< m1 >>
rect 325 321 326 322 
<< m1 >>
rect 327 321 328 322 
<< m1 >>
rect 329 321 330 322 
<< m1 >>
rect 331 321 332 322 
<< m1 >>
rect 334 321 335 322 
<< pdiffusion >>
rect 336 321 337 322 
<< pdiffusion >>
rect 337 321 338 322 
<< pdiffusion >>
rect 338 321 339 322 
<< pdiffusion >>
rect 339 321 340 322 
<< pdiffusion >>
rect 340 321 341 322 
<< pdiffusion >>
rect 341 321 342 322 
<< m1 >>
rect 343 321 344 322 
<< m1 >>
rect 10 322 11 323 
<< pdiffusion >>
rect 12 322 13 323 
<< pdiffusion >>
rect 13 322 14 323 
<< pdiffusion >>
rect 14 322 15 323 
<< pdiffusion >>
rect 15 322 16 323 
<< pdiffusion >>
rect 16 322 17 323 
<< pdiffusion >>
rect 17 322 18 323 
<< m1 >>
rect 28 322 29 323 
<< pdiffusion >>
rect 30 322 31 323 
<< pdiffusion >>
rect 31 322 32 323 
<< pdiffusion >>
rect 32 322 33 323 
<< pdiffusion >>
rect 33 322 34 323 
<< pdiffusion >>
rect 34 322 35 323 
<< pdiffusion >>
rect 35 322 36 323 
<< m1 >>
rect 37 322 38 323 
<< m2 >>
rect 38 322 39 323 
<< m1 >>
rect 46 322 47 323 
<< pdiffusion >>
rect 48 322 49 323 
<< pdiffusion >>
rect 49 322 50 323 
<< pdiffusion >>
rect 50 322 51 323 
<< pdiffusion >>
rect 51 322 52 323 
<< pdiffusion >>
rect 52 322 53 323 
<< pdiffusion >>
rect 53 322 54 323 
<< m1 >>
rect 55 322 56 323 
<< m1 >>
rect 57 322 58 323 
<< m1 >>
rect 60 322 61 323 
<< m1 >>
rect 62 322 63 323 
<< m1 >>
rect 64 322 65 323 
<< pdiffusion >>
rect 66 322 67 323 
<< pdiffusion >>
rect 67 322 68 323 
<< pdiffusion >>
rect 68 322 69 323 
<< pdiffusion >>
rect 69 322 70 323 
<< pdiffusion >>
rect 70 322 71 323 
<< pdiffusion >>
rect 71 322 72 323 
<< m1 >>
rect 73 322 74 323 
<< m1 >>
rect 75 322 76 323 
<< m1 >>
rect 82 322 83 323 
<< pdiffusion >>
rect 84 322 85 323 
<< pdiffusion >>
rect 85 322 86 323 
<< pdiffusion >>
rect 86 322 87 323 
<< pdiffusion >>
rect 87 322 88 323 
<< pdiffusion >>
rect 88 322 89 323 
<< pdiffusion >>
rect 89 322 90 323 
<< m1 >>
rect 91 322 92 323 
<< m1 >>
rect 100 322 101 323 
<< pdiffusion >>
rect 102 322 103 323 
<< pdiffusion >>
rect 103 322 104 323 
<< pdiffusion >>
rect 104 322 105 323 
<< pdiffusion >>
rect 105 322 106 323 
<< pdiffusion >>
rect 106 322 107 323 
<< pdiffusion >>
rect 107 322 108 323 
<< pdiffusion >>
rect 120 322 121 323 
<< pdiffusion >>
rect 121 322 122 323 
<< pdiffusion >>
rect 122 322 123 323 
<< pdiffusion >>
rect 123 322 124 323 
<< pdiffusion >>
rect 124 322 125 323 
<< pdiffusion >>
rect 125 322 126 323 
<< pdiffusion >>
rect 138 322 139 323 
<< pdiffusion >>
rect 139 322 140 323 
<< pdiffusion >>
rect 140 322 141 323 
<< pdiffusion >>
rect 141 322 142 323 
<< pdiffusion >>
rect 142 322 143 323 
<< pdiffusion >>
rect 143 322 144 323 
<< pdiffusion >>
rect 156 322 157 323 
<< pdiffusion >>
rect 157 322 158 323 
<< pdiffusion >>
rect 158 322 159 323 
<< pdiffusion >>
rect 159 322 160 323 
<< pdiffusion >>
rect 160 322 161 323 
<< pdiffusion >>
rect 161 322 162 323 
<< m1 >>
rect 172 322 173 323 
<< pdiffusion >>
rect 174 322 175 323 
<< pdiffusion >>
rect 175 322 176 323 
<< pdiffusion >>
rect 176 322 177 323 
<< pdiffusion >>
rect 177 322 178 323 
<< pdiffusion >>
rect 178 322 179 323 
<< pdiffusion >>
rect 179 322 180 323 
<< pdiffusion >>
rect 192 322 193 323 
<< pdiffusion >>
rect 193 322 194 323 
<< pdiffusion >>
rect 194 322 195 323 
<< pdiffusion >>
rect 195 322 196 323 
<< pdiffusion >>
rect 196 322 197 323 
<< pdiffusion >>
rect 197 322 198 323 
<< m1 >>
rect 199 322 200 323 
<< pdiffusion >>
rect 210 322 211 323 
<< pdiffusion >>
rect 211 322 212 323 
<< pdiffusion >>
rect 212 322 213 323 
<< pdiffusion >>
rect 213 322 214 323 
<< pdiffusion >>
rect 214 322 215 323 
<< pdiffusion >>
rect 215 322 216 323 
<< m1 >>
rect 217 322 218 323 
<< m2 >>
rect 217 322 218 323 
<< m1 >>
rect 219 322 220 323 
<< m1 >>
rect 223 322 224 323 
<< pdiffusion >>
rect 228 322 229 323 
<< pdiffusion >>
rect 229 322 230 323 
<< pdiffusion >>
rect 230 322 231 323 
<< pdiffusion >>
rect 231 322 232 323 
<< pdiffusion >>
rect 232 322 233 323 
<< pdiffusion >>
rect 233 322 234 323 
<< m1 >>
rect 239 322 240 323 
<< pdiffusion >>
rect 246 322 247 323 
<< pdiffusion >>
rect 247 322 248 323 
<< pdiffusion >>
rect 248 322 249 323 
<< pdiffusion >>
rect 249 322 250 323 
<< pdiffusion >>
rect 250 322 251 323 
<< pdiffusion >>
rect 251 322 252 323 
<< m1 >>
rect 253 322 254 323 
<< m1 >>
rect 255 322 256 323 
<< pdiffusion >>
rect 264 322 265 323 
<< pdiffusion >>
rect 265 322 266 323 
<< pdiffusion >>
rect 266 322 267 323 
<< pdiffusion >>
rect 267 322 268 323 
<< pdiffusion >>
rect 268 322 269 323 
<< pdiffusion >>
rect 269 322 270 323 
<< m1 >>
rect 271 322 272 323 
<< m1 >>
rect 275 322 276 323 
<< m2 >>
rect 275 322 276 323 
<< pdiffusion >>
rect 282 322 283 323 
<< pdiffusion >>
rect 283 322 284 323 
<< pdiffusion >>
rect 284 322 285 323 
<< pdiffusion >>
rect 285 322 286 323 
<< pdiffusion >>
rect 286 322 287 323 
<< pdiffusion >>
rect 287 322 288 323 
<< pdiffusion >>
rect 300 322 301 323 
<< pdiffusion >>
rect 301 322 302 323 
<< pdiffusion >>
rect 302 322 303 323 
<< pdiffusion >>
rect 303 322 304 323 
<< pdiffusion >>
rect 304 322 305 323 
<< pdiffusion >>
rect 305 322 306 323 
<< m1 >>
rect 307 322 308 323 
<< pdiffusion >>
rect 318 322 319 323 
<< pdiffusion >>
rect 319 322 320 323 
<< pdiffusion >>
rect 320 322 321 323 
<< pdiffusion >>
rect 321 322 322 323 
<< pdiffusion >>
rect 322 322 323 323 
<< pdiffusion >>
rect 323 322 324 323 
<< m1 >>
rect 325 322 326 323 
<< m1 >>
rect 327 322 328 323 
<< m1 >>
rect 329 322 330 323 
<< m1 >>
rect 331 322 332 323 
<< m1 >>
rect 334 322 335 323 
<< pdiffusion >>
rect 336 322 337 323 
<< pdiffusion >>
rect 337 322 338 323 
<< pdiffusion >>
rect 338 322 339 323 
<< pdiffusion >>
rect 339 322 340 323 
<< pdiffusion >>
rect 340 322 341 323 
<< pdiffusion >>
rect 341 322 342 323 
<< m1 >>
rect 343 322 344 323 
<< m1 >>
rect 10 323 11 324 
<< pdiffusion >>
rect 12 323 13 324 
<< pdiffusion >>
rect 13 323 14 324 
<< pdiffusion >>
rect 14 323 15 324 
<< pdiffusion >>
rect 15 323 16 324 
<< pdiffusion >>
rect 16 323 17 324 
<< pdiffusion >>
rect 17 323 18 324 
<< m1 >>
rect 28 323 29 324 
<< pdiffusion >>
rect 30 323 31 324 
<< pdiffusion >>
rect 31 323 32 324 
<< pdiffusion >>
rect 32 323 33 324 
<< pdiffusion >>
rect 33 323 34 324 
<< m1 >>
rect 34 323 35 324 
<< pdiffusion >>
rect 34 323 35 324 
<< pdiffusion >>
rect 35 323 36 324 
<< m1 >>
rect 37 323 38 324 
<< m2 >>
rect 38 323 39 324 
<< m1 >>
rect 46 323 47 324 
<< pdiffusion >>
rect 48 323 49 324 
<< pdiffusion >>
rect 49 323 50 324 
<< pdiffusion >>
rect 50 323 51 324 
<< pdiffusion >>
rect 51 323 52 324 
<< m1 >>
rect 52 323 53 324 
<< pdiffusion >>
rect 52 323 53 324 
<< pdiffusion >>
rect 53 323 54 324 
<< m1 >>
rect 55 323 56 324 
<< m1 >>
rect 57 323 58 324 
<< m1 >>
rect 60 323 61 324 
<< m1 >>
rect 62 323 63 324 
<< m1 >>
rect 64 323 65 324 
<< pdiffusion >>
rect 66 323 67 324 
<< pdiffusion >>
rect 67 323 68 324 
<< pdiffusion >>
rect 68 323 69 324 
<< pdiffusion >>
rect 69 323 70 324 
<< m1 >>
rect 70 323 71 324 
<< pdiffusion >>
rect 70 323 71 324 
<< pdiffusion >>
rect 71 323 72 324 
<< m1 >>
rect 73 323 74 324 
<< m2 >>
rect 73 323 74 324 
<< m2c >>
rect 73 323 74 324 
<< m1 >>
rect 73 323 74 324 
<< m2 >>
rect 73 323 74 324 
<< m1 >>
rect 75 323 76 324 
<< m2 >>
rect 75 323 76 324 
<< m2c >>
rect 75 323 76 324 
<< m1 >>
rect 75 323 76 324 
<< m2 >>
rect 75 323 76 324 
<< m1 >>
rect 82 323 83 324 
<< pdiffusion >>
rect 84 323 85 324 
<< pdiffusion >>
rect 85 323 86 324 
<< pdiffusion >>
rect 86 323 87 324 
<< pdiffusion >>
rect 87 323 88 324 
<< pdiffusion >>
rect 88 323 89 324 
<< pdiffusion >>
rect 89 323 90 324 
<< m1 >>
rect 91 323 92 324 
<< m1 >>
rect 100 323 101 324 
<< pdiffusion >>
rect 102 323 103 324 
<< pdiffusion >>
rect 103 323 104 324 
<< pdiffusion >>
rect 104 323 105 324 
<< pdiffusion >>
rect 105 323 106 324 
<< pdiffusion >>
rect 106 323 107 324 
<< pdiffusion >>
rect 107 323 108 324 
<< pdiffusion >>
rect 120 323 121 324 
<< m1 >>
rect 121 323 122 324 
<< pdiffusion >>
rect 121 323 122 324 
<< pdiffusion >>
rect 122 323 123 324 
<< pdiffusion >>
rect 123 323 124 324 
<< pdiffusion >>
rect 124 323 125 324 
<< pdiffusion >>
rect 125 323 126 324 
<< pdiffusion >>
rect 138 323 139 324 
<< pdiffusion >>
rect 139 323 140 324 
<< pdiffusion >>
rect 140 323 141 324 
<< pdiffusion >>
rect 141 323 142 324 
<< pdiffusion >>
rect 142 323 143 324 
<< pdiffusion >>
rect 143 323 144 324 
<< pdiffusion >>
rect 156 323 157 324 
<< pdiffusion >>
rect 157 323 158 324 
<< pdiffusion >>
rect 158 323 159 324 
<< pdiffusion >>
rect 159 323 160 324 
<< pdiffusion >>
rect 160 323 161 324 
<< pdiffusion >>
rect 161 323 162 324 
<< m1 >>
rect 172 323 173 324 
<< pdiffusion >>
rect 174 323 175 324 
<< pdiffusion >>
rect 175 323 176 324 
<< pdiffusion >>
rect 176 323 177 324 
<< pdiffusion >>
rect 177 323 178 324 
<< pdiffusion >>
rect 178 323 179 324 
<< pdiffusion >>
rect 179 323 180 324 
<< pdiffusion >>
rect 192 323 193 324 
<< pdiffusion >>
rect 193 323 194 324 
<< pdiffusion >>
rect 194 323 195 324 
<< pdiffusion >>
rect 195 323 196 324 
<< pdiffusion >>
rect 196 323 197 324 
<< pdiffusion >>
rect 197 323 198 324 
<< m1 >>
rect 199 323 200 324 
<< pdiffusion >>
rect 210 323 211 324 
<< pdiffusion >>
rect 211 323 212 324 
<< pdiffusion >>
rect 212 323 213 324 
<< pdiffusion >>
rect 213 323 214 324 
<< pdiffusion >>
rect 214 323 215 324 
<< pdiffusion >>
rect 215 323 216 324 
<< m1 >>
rect 217 323 218 324 
<< m2 >>
rect 217 323 218 324 
<< m1 >>
rect 219 323 220 324 
<< m1 >>
rect 223 323 224 324 
<< pdiffusion >>
rect 228 323 229 324 
<< pdiffusion >>
rect 229 323 230 324 
<< pdiffusion >>
rect 230 323 231 324 
<< pdiffusion >>
rect 231 323 232 324 
<< pdiffusion >>
rect 232 323 233 324 
<< pdiffusion >>
rect 233 323 234 324 
<< m1 >>
rect 239 323 240 324 
<< pdiffusion >>
rect 246 323 247 324 
<< pdiffusion >>
rect 247 323 248 324 
<< pdiffusion >>
rect 248 323 249 324 
<< pdiffusion >>
rect 249 323 250 324 
<< pdiffusion >>
rect 250 323 251 324 
<< pdiffusion >>
rect 251 323 252 324 
<< m1 >>
rect 253 323 254 324 
<< m1 >>
rect 255 323 256 324 
<< pdiffusion >>
rect 264 323 265 324 
<< pdiffusion >>
rect 265 323 266 324 
<< pdiffusion >>
rect 266 323 267 324 
<< pdiffusion >>
rect 267 323 268 324 
<< m1 >>
rect 268 323 269 324 
<< pdiffusion >>
rect 268 323 269 324 
<< pdiffusion >>
rect 269 323 270 324 
<< m1 >>
rect 271 323 272 324 
<< m1 >>
rect 275 323 276 324 
<< m2 >>
rect 275 323 276 324 
<< pdiffusion >>
rect 282 323 283 324 
<< pdiffusion >>
rect 283 323 284 324 
<< pdiffusion >>
rect 284 323 285 324 
<< pdiffusion >>
rect 285 323 286 324 
<< pdiffusion >>
rect 286 323 287 324 
<< pdiffusion >>
rect 287 323 288 324 
<< pdiffusion >>
rect 300 323 301 324 
<< m1 >>
rect 301 323 302 324 
<< pdiffusion >>
rect 301 323 302 324 
<< pdiffusion >>
rect 302 323 303 324 
<< pdiffusion >>
rect 303 323 304 324 
<< pdiffusion >>
rect 304 323 305 324 
<< pdiffusion >>
rect 305 323 306 324 
<< m1 >>
rect 307 323 308 324 
<< pdiffusion >>
rect 318 323 319 324 
<< pdiffusion >>
rect 319 323 320 324 
<< pdiffusion >>
rect 320 323 321 324 
<< pdiffusion >>
rect 321 323 322 324 
<< pdiffusion >>
rect 322 323 323 324 
<< pdiffusion >>
rect 323 323 324 324 
<< m1 >>
rect 325 323 326 324 
<< m1 >>
rect 327 323 328 324 
<< m1 >>
rect 329 323 330 324 
<< m1 >>
rect 331 323 332 324 
<< m1 >>
rect 334 323 335 324 
<< pdiffusion >>
rect 336 323 337 324 
<< pdiffusion >>
rect 337 323 338 324 
<< pdiffusion >>
rect 338 323 339 324 
<< pdiffusion >>
rect 339 323 340 324 
<< m1 >>
rect 340 323 341 324 
<< pdiffusion >>
rect 340 323 341 324 
<< pdiffusion >>
rect 341 323 342 324 
<< m1 >>
rect 343 323 344 324 
<< m1 >>
rect 10 324 11 325 
<< m1 >>
rect 28 324 29 325 
<< m1 >>
rect 34 324 35 325 
<< m1 >>
rect 37 324 38 325 
<< m2 >>
rect 38 324 39 325 
<< m1 >>
rect 46 324 47 325 
<< m1 >>
rect 52 324 53 325 
<< m1 >>
rect 55 324 56 325 
<< m1 >>
rect 57 324 58 325 
<< m1 >>
rect 60 324 61 325 
<< m1 >>
rect 62 324 63 325 
<< m1 >>
rect 64 324 65 325 
<< m1 >>
rect 70 324 71 325 
<< m2 >>
rect 73 324 74 325 
<< m2 >>
rect 75 324 76 325 
<< m1 >>
rect 82 324 83 325 
<< m1 >>
rect 91 324 92 325 
<< m1 >>
rect 100 324 101 325 
<< m1 >>
rect 121 324 122 325 
<< m1 >>
rect 172 324 173 325 
<< m1 >>
rect 199 324 200 325 
<< m1 >>
rect 217 324 218 325 
<< m2 >>
rect 217 324 218 325 
<< m2 >>
rect 218 324 219 325 
<< m1 >>
rect 219 324 220 325 
<< m2 >>
rect 219 324 220 325 
<< m2 >>
rect 220 324 221 325 
<< m1 >>
rect 221 324 222 325 
<< m2 >>
rect 221 324 222 325 
<< m2c >>
rect 221 324 222 325 
<< m1 >>
rect 221 324 222 325 
<< m2 >>
rect 221 324 222 325 
<< m1 >>
rect 223 324 224 325 
<< m1 >>
rect 239 324 240 325 
<< m1 >>
rect 253 324 254 325 
<< m1 >>
rect 255 324 256 325 
<< m1 >>
rect 268 324 269 325 
<< m1 >>
rect 271 324 272 325 
<< m1 >>
rect 275 324 276 325 
<< m2 >>
rect 275 324 276 325 
<< m1 >>
rect 301 324 302 325 
<< m1 >>
rect 307 324 308 325 
<< m1 >>
rect 325 324 326 325 
<< m1 >>
rect 327 324 328 325 
<< m1 >>
rect 329 324 330 325 
<< m1 >>
rect 331 324 332 325 
<< m1 >>
rect 334 324 335 325 
<< m1 >>
rect 340 324 341 325 
<< m1 >>
rect 343 324 344 325 
<< m1 >>
rect 10 325 11 326 
<< m1 >>
rect 28 325 29 326 
<< m1 >>
rect 34 325 35 326 
<< m1 >>
rect 37 325 38 326 
<< m2 >>
rect 38 325 39 326 
<< m1 >>
rect 46 325 47 326 
<< m1 >>
rect 52 325 53 326 
<< m1 >>
rect 53 325 54 326 
<< m1 >>
rect 54 325 55 326 
<< m1 >>
rect 55 325 56 326 
<< m1 >>
rect 57 325 58 326 
<< m1 >>
rect 60 325 61 326 
<< m1 >>
rect 62 325 63 326 
<< m1 >>
rect 64 325 65 326 
<< m1 >>
rect 70 325 71 326 
<< m1 >>
rect 71 325 72 326 
<< m1 >>
rect 72 325 73 326 
<< m1 >>
rect 73 325 74 326 
<< m2 >>
rect 73 325 74 326 
<< m1 >>
rect 74 325 75 326 
<< m1 >>
rect 75 325 76 326 
<< m2 >>
rect 75 325 76 326 
<< m1 >>
rect 76 325 77 326 
<< m1 >>
rect 77 325 78 326 
<< m1 >>
rect 78 325 79 326 
<< m1 >>
rect 79 325 80 326 
<< m1 >>
rect 80 325 81 326 
<< m1 >>
rect 81 325 82 326 
<< m1 >>
rect 82 325 83 326 
<< m1 >>
rect 91 325 92 326 
<< m1 >>
rect 100 325 101 326 
<< m1 >>
rect 121 325 122 326 
<< m1 >>
rect 172 325 173 326 
<< m1 >>
rect 199 325 200 326 
<< m1 >>
rect 217 325 218 326 
<< m1 >>
rect 219 325 220 326 
<< m1 >>
rect 221 325 222 326 
<< m1 >>
rect 223 325 224 326 
<< m1 >>
rect 239 325 240 326 
<< m1 >>
rect 253 325 254 326 
<< m1 >>
rect 255 325 256 326 
<< m1 >>
rect 268 325 269 326 
<< m1 >>
rect 271 325 272 326 
<< m1 >>
rect 275 325 276 326 
<< m2 >>
rect 275 325 276 326 
<< m1 >>
rect 301 325 302 326 
<< m1 >>
rect 307 325 308 326 
<< m1 >>
rect 325 325 326 326 
<< m1 >>
rect 327 325 328 326 
<< m1 >>
rect 329 325 330 326 
<< m1 >>
rect 331 325 332 326 
<< m1 >>
rect 334 325 335 326 
<< m1 >>
rect 340 325 341 326 
<< m1 >>
rect 343 325 344 326 
<< m1 >>
rect 10 326 11 327 
<< m1 >>
rect 28 326 29 327 
<< m1 >>
rect 34 326 35 327 
<< m1 >>
rect 37 326 38 327 
<< m2 >>
rect 38 326 39 327 
<< m1 >>
rect 46 326 47 327 
<< m1 >>
rect 47 326 48 327 
<< m1 >>
rect 48 326 49 327 
<< m2 >>
rect 48 326 49 327 
<< m2c >>
rect 48 326 49 327 
<< m1 >>
rect 48 326 49 327 
<< m2 >>
rect 48 326 49 327 
<< m1 >>
rect 57 326 58 327 
<< m1 >>
rect 60 326 61 327 
<< m1 >>
rect 62 326 63 327 
<< m1 >>
rect 64 326 65 327 
<< m2 >>
rect 73 326 74 327 
<< m2 >>
rect 75 326 76 327 
<< m1 >>
rect 86 326 87 327 
<< m2 >>
rect 86 326 87 327 
<< m2c >>
rect 86 326 87 327 
<< m1 >>
rect 86 326 87 327 
<< m2 >>
rect 86 326 87 327 
<< m1 >>
rect 87 326 88 327 
<< m1 >>
rect 88 326 89 327 
<< m1 >>
rect 89 326 90 327 
<< m1 >>
rect 90 326 91 327 
<< m1 >>
rect 91 326 92 327 
<< m1 >>
rect 100 326 101 327 
<< m1 >>
rect 101 326 102 327 
<< m1 >>
rect 102 326 103 327 
<< m2 >>
rect 102 326 103 327 
<< m2c >>
rect 102 326 103 327 
<< m1 >>
rect 102 326 103 327 
<< m2 >>
rect 102 326 103 327 
<< m1 >>
rect 121 326 122 327 
<< m1 >>
rect 158 326 159 327 
<< m2 >>
rect 158 326 159 327 
<< m2c >>
rect 158 326 159 327 
<< m1 >>
rect 158 326 159 327 
<< m2 >>
rect 158 326 159 327 
<< m1 >>
rect 159 326 160 327 
<< m1 >>
rect 160 326 161 327 
<< m1 >>
rect 161 326 162 327 
<< m1 >>
rect 162 326 163 327 
<< m1 >>
rect 163 326 164 327 
<< m1 >>
rect 164 326 165 327 
<< m1 >>
rect 165 326 166 327 
<< m1 >>
rect 166 326 167 327 
<< m1 >>
rect 167 326 168 327 
<< m1 >>
rect 168 326 169 327 
<< m1 >>
rect 169 326 170 327 
<< m1 >>
rect 170 326 171 327 
<< m1 >>
rect 171 326 172 327 
<< m1 >>
rect 172 326 173 327 
<< m1 >>
rect 194 326 195 327 
<< m2 >>
rect 194 326 195 327 
<< m2c >>
rect 194 326 195 327 
<< m1 >>
rect 194 326 195 327 
<< m2 >>
rect 194 326 195 327 
<< m1 >>
rect 195 326 196 327 
<< m1 >>
rect 196 326 197 327 
<< m1 >>
rect 197 326 198 327 
<< m1 >>
rect 198 326 199 327 
<< m1 >>
rect 199 326 200 327 
<< m1 >>
rect 217 326 218 327 
<< m2 >>
rect 217 326 218 327 
<< m2c >>
rect 217 326 218 327 
<< m1 >>
rect 217 326 218 327 
<< m2 >>
rect 217 326 218 327 
<< m1 >>
rect 219 326 220 327 
<< m2 >>
rect 219 326 220 327 
<< m2c >>
rect 219 326 220 327 
<< m1 >>
rect 219 326 220 327 
<< m2 >>
rect 219 326 220 327 
<< m1 >>
rect 221 326 222 327 
<< m2 >>
rect 221 326 222 327 
<< m2c >>
rect 221 326 222 327 
<< m1 >>
rect 221 326 222 327 
<< m2 >>
rect 221 326 222 327 
<< m1 >>
rect 223 326 224 327 
<< m2 >>
rect 223 326 224 327 
<< m2c >>
rect 223 326 224 327 
<< m1 >>
rect 223 326 224 327 
<< m2 >>
rect 223 326 224 327 
<< m1 >>
rect 239 326 240 327 
<< m2 >>
rect 239 326 240 327 
<< m2c >>
rect 239 326 240 327 
<< m1 >>
rect 239 326 240 327 
<< m2 >>
rect 239 326 240 327 
<< m2 >>
rect 252 326 253 327 
<< m1 >>
rect 253 326 254 327 
<< m2 >>
rect 253 326 254 327 
<< m2 >>
rect 254 326 255 327 
<< m1 >>
rect 255 326 256 327 
<< m2 >>
rect 255 326 256 327 
<< m2c >>
rect 255 326 256 327 
<< m1 >>
rect 255 326 256 327 
<< m2 >>
rect 255 326 256 327 
<< m1 >>
rect 268 326 269 327 
<< m2 >>
rect 268 326 269 327 
<< m2c >>
rect 268 326 269 327 
<< m1 >>
rect 268 326 269 327 
<< m2 >>
rect 268 326 269 327 
<< m1 >>
rect 271 326 272 327 
<< m2 >>
rect 271 326 272 327 
<< m2c >>
rect 271 326 272 327 
<< m1 >>
rect 271 326 272 327 
<< m2 >>
rect 271 326 272 327 
<< m1 >>
rect 273 326 274 327 
<< m2 >>
rect 273 326 274 327 
<< m2c >>
rect 273 326 274 327 
<< m1 >>
rect 273 326 274 327 
<< m2 >>
rect 273 326 274 327 
<< m1 >>
rect 274 326 275 327 
<< m1 >>
rect 275 326 276 327 
<< m2 >>
rect 275 326 276 327 
<< m1 >>
rect 301 326 302 327 
<< m1 >>
rect 302 326 303 327 
<< m1 >>
rect 303 326 304 327 
<< m1 >>
rect 304 326 305 327 
<< m1 >>
rect 305 326 306 327 
<< m1 >>
rect 306 326 307 327 
<< m1 >>
rect 307 326 308 327 
<< m1 >>
rect 323 326 324 327 
<< m2 >>
rect 323 326 324 327 
<< m2c >>
rect 323 326 324 327 
<< m1 >>
rect 323 326 324 327 
<< m2 >>
rect 323 326 324 327 
<< m1 >>
rect 324 326 325 327 
<< m1 >>
rect 325 326 326 327 
<< m2 >>
rect 325 326 326 327 
<< m2 >>
rect 326 326 327 327 
<< m1 >>
rect 327 326 328 327 
<< m2 >>
rect 327 326 328 327 
<< m2c >>
rect 327 326 328 327 
<< m1 >>
rect 327 326 328 327 
<< m2 >>
rect 327 326 328 327 
<< m1 >>
rect 329 326 330 327 
<< m2 >>
rect 329 326 330 327 
<< m2c >>
rect 329 326 330 327 
<< m1 >>
rect 329 326 330 327 
<< m2 >>
rect 329 326 330 327 
<< m1 >>
rect 331 326 332 327 
<< m2 >>
rect 331 326 332 327 
<< m2c >>
rect 331 326 332 327 
<< m1 >>
rect 331 326 332 327 
<< m2 >>
rect 331 326 332 327 
<< m1 >>
rect 334 326 335 327 
<< m2 >>
rect 334 326 335 327 
<< m2c >>
rect 334 326 335 327 
<< m1 >>
rect 334 326 335 327 
<< m2 >>
rect 334 326 335 327 
<< m1 >>
rect 340 326 341 327 
<< m2 >>
rect 340 326 341 327 
<< m2c >>
rect 340 326 341 327 
<< m1 >>
rect 340 326 341 327 
<< m2 >>
rect 340 326 341 327 
<< m1 >>
rect 343 326 344 327 
<< m1 >>
rect 10 327 11 328 
<< m1 >>
rect 28 327 29 328 
<< m1 >>
rect 34 327 35 328 
<< m1 >>
rect 37 327 38 328 
<< m2 >>
rect 38 327 39 328 
<< m2 >>
rect 48 327 49 328 
<< m1 >>
rect 57 327 58 328 
<< m1 >>
rect 60 327 61 328 
<< m1 >>
rect 62 327 63 328 
<< m1 >>
rect 64 327 65 328 
<< m2 >>
rect 73 327 74 328 
<< m2 >>
rect 75 327 76 328 
<< m2 >>
rect 86 327 87 328 
<< m2 >>
rect 102 327 103 328 
<< m1 >>
rect 121 327 122 328 
<< m2 >>
rect 158 327 159 328 
<< m2 >>
rect 194 327 195 328 
<< m2 >>
rect 217 327 218 328 
<< m2 >>
rect 219 327 220 328 
<< m2 >>
rect 221 327 222 328 
<< m2 >>
rect 223 327 224 328 
<< m2 >>
rect 239 327 240 328 
<< m2 >>
rect 252 327 253 328 
<< m1 >>
rect 253 327 254 328 
<< m2 >>
rect 268 327 269 328 
<< m2 >>
rect 271 327 272 328 
<< m2 >>
rect 273 327 274 328 
<< m2 >>
rect 275 327 276 328 
<< m2 >>
rect 323 327 324 328 
<< m2 >>
rect 325 327 326 328 
<< m2 >>
rect 329 327 330 328 
<< m2 >>
rect 331 327 332 328 
<< m2 >>
rect 334 327 335 328 
<< m2 >>
rect 340 327 341 328 
<< m1 >>
rect 343 327 344 328 
<< m1 >>
rect 10 328 11 329 
<< m1 >>
rect 26 328 27 329 
<< m2 >>
rect 26 328 27 329 
<< m2c >>
rect 26 328 27 329 
<< m1 >>
rect 26 328 27 329 
<< m2 >>
rect 26 328 27 329 
<< m2 >>
rect 27 328 28 329 
<< m1 >>
rect 28 328 29 329 
<< m2 >>
rect 28 328 29 329 
<< m2 >>
rect 29 328 30 329 
<< m1 >>
rect 30 328 31 329 
<< m2 >>
rect 30 328 31 329 
<< m2c >>
rect 30 328 31 329 
<< m1 >>
rect 30 328 31 329 
<< m2 >>
rect 30 328 31 329 
<< m1 >>
rect 31 328 32 329 
<< m1 >>
rect 32 328 33 329 
<< m1 >>
rect 33 328 34 329 
<< m1 >>
rect 34 328 35 329 
<< m1 >>
rect 37 328 38 329 
<< m1 >>
rect 38 328 39 329 
<< m2 >>
rect 38 328 39 329 
<< m1 >>
rect 39 328 40 329 
<< m1 >>
rect 40 328 41 329 
<< m1 >>
rect 41 328 42 329 
<< m1 >>
rect 42 328 43 329 
<< m1 >>
rect 43 328 44 329 
<< m1 >>
rect 44 328 45 329 
<< m1 >>
rect 45 328 46 329 
<< m1 >>
rect 46 328 47 329 
<< m1 >>
rect 47 328 48 329 
<< m1 >>
rect 48 328 49 329 
<< m2 >>
rect 48 328 49 329 
<< m1 >>
rect 49 328 50 329 
<< m1 >>
rect 52 328 53 329 
<< m1 >>
rect 53 328 54 329 
<< m1 >>
rect 54 328 55 329 
<< m2 >>
rect 54 328 55 329 
<< m2c >>
rect 54 328 55 329 
<< m1 >>
rect 54 328 55 329 
<< m2 >>
rect 54 328 55 329 
<< m2 >>
rect 55 328 56 329 
<< m2 >>
rect 56 328 57 329 
<< m1 >>
rect 57 328 58 329 
<< m2 >>
rect 57 328 58 329 
<< m2 >>
rect 58 328 59 329 
<< m2 >>
rect 59 328 60 329 
<< m1 >>
rect 60 328 61 329 
<< m2 >>
rect 60 328 61 329 
<< m2 >>
rect 61 328 62 329 
<< m1 >>
rect 62 328 63 329 
<< m2 >>
rect 62 328 63 329 
<< m2 >>
rect 63 328 64 329 
<< m1 >>
rect 64 328 65 329 
<< m2 >>
rect 64 328 65 329 
<< m1 >>
rect 65 328 66 329 
<< m2 >>
rect 65 328 66 329 
<< m1 >>
rect 66 328 67 329 
<< m2 >>
rect 66 328 67 329 
<< m1 >>
rect 67 328 68 329 
<< m2 >>
rect 67 328 68 329 
<< m1 >>
rect 68 328 69 329 
<< m2 >>
rect 68 328 69 329 
<< m1 >>
rect 69 328 70 329 
<< m2 >>
rect 69 328 70 329 
<< m1 >>
rect 70 328 71 329 
<< m2 >>
rect 70 328 71 329 
<< m1 >>
rect 71 328 72 329 
<< m2 >>
rect 71 328 72 329 
<< m1 >>
rect 72 328 73 329 
<< m2 >>
rect 72 328 73 329 
<< m1 >>
rect 73 328 74 329 
<< m2 >>
rect 73 328 74 329 
<< m1 >>
rect 74 328 75 329 
<< m1 >>
rect 75 328 76 329 
<< m2 >>
rect 75 328 76 329 
<< m1 >>
rect 76 328 77 329 
<< m2 >>
rect 76 328 77 329 
<< m1 >>
rect 77 328 78 329 
<< m2 >>
rect 77 328 78 329 
<< m1 >>
rect 78 328 79 329 
<< m2 >>
rect 78 328 79 329 
<< m1 >>
rect 79 328 80 329 
<< m2 >>
rect 79 328 80 329 
<< m1 >>
rect 80 328 81 329 
<< m2 >>
rect 80 328 81 329 
<< m1 >>
rect 81 328 82 329 
<< m2 >>
rect 81 328 82 329 
<< m1 >>
rect 82 328 83 329 
<< m2 >>
rect 82 328 83 329 
<< m1 >>
rect 83 328 84 329 
<< m2 >>
rect 83 328 84 329 
<< m1 >>
rect 84 328 85 329 
<< m2 >>
rect 84 328 85 329 
<< m1 >>
rect 85 328 86 329 
<< m2 >>
rect 85 328 86 329 
<< m1 >>
rect 86 328 87 329 
<< m2 >>
rect 86 328 87 329 
<< m1 >>
rect 87 328 88 329 
<< m1 >>
rect 88 328 89 329 
<< m1 >>
rect 89 328 90 329 
<< m1 >>
rect 90 328 91 329 
<< m1 >>
rect 91 328 92 329 
<< m1 >>
rect 92 328 93 329 
<< m1 >>
rect 93 328 94 329 
<< m1 >>
rect 94 328 95 329 
<< m1 >>
rect 95 328 96 329 
<< m1 >>
rect 96 328 97 329 
<< m1 >>
rect 97 328 98 329 
<< m1 >>
rect 98 328 99 329 
<< m1 >>
rect 99 328 100 329 
<< m1 >>
rect 100 328 101 329 
<< m1 >>
rect 101 328 102 329 
<< m1 >>
rect 102 328 103 329 
<< m2 >>
rect 102 328 103 329 
<< m1 >>
rect 103 328 104 329 
<< m1 >>
rect 104 328 105 329 
<< m1 >>
rect 105 328 106 329 
<< m1 >>
rect 106 328 107 329 
<< m1 >>
rect 107 328 108 329 
<< m1 >>
rect 108 328 109 329 
<< m1 >>
rect 109 328 110 329 
<< m1 >>
rect 110 328 111 329 
<< m1 >>
rect 111 328 112 329 
<< m1 >>
rect 112 328 113 329 
<< m1 >>
rect 113 328 114 329 
<< m1 >>
rect 114 328 115 329 
<< m1 >>
rect 115 328 116 329 
<< m1 >>
rect 116 328 117 329 
<< m1 >>
rect 117 328 118 329 
<< m1 >>
rect 118 328 119 329 
<< m1 >>
rect 119 328 120 329 
<< m2 >>
rect 119 328 120 329 
<< m2c >>
rect 119 328 120 329 
<< m1 >>
rect 119 328 120 329 
<< m2 >>
rect 119 328 120 329 
<< m2 >>
rect 120 328 121 329 
<< m1 >>
rect 121 328 122 329 
<< m2 >>
rect 121 328 122 329 
<< m1 >>
rect 122 328 123 329 
<< m2 >>
rect 122 328 123 329 
<< m1 >>
rect 123 328 124 329 
<< m2 >>
rect 123 328 124 329 
<< m1 >>
rect 124 328 125 329 
<< m2 >>
rect 124 328 125 329 
<< m1 >>
rect 125 328 126 329 
<< m2 >>
rect 125 328 126 329 
<< m1 >>
rect 126 328 127 329 
<< m2 >>
rect 126 328 127 329 
<< m1 >>
rect 127 328 128 329 
<< m2 >>
rect 127 328 128 329 
<< m1 >>
rect 128 328 129 329 
<< m2 >>
rect 128 328 129 329 
<< m1 >>
rect 129 328 130 329 
<< m2 >>
rect 129 328 130 329 
<< m1 >>
rect 130 328 131 329 
<< m2 >>
rect 130 328 131 329 
<< m1 >>
rect 131 328 132 329 
<< m2 >>
rect 131 328 132 329 
<< m1 >>
rect 132 328 133 329 
<< m2 >>
rect 132 328 133 329 
<< m1 >>
rect 133 328 134 329 
<< m2 >>
rect 133 328 134 329 
<< m1 >>
rect 134 328 135 329 
<< m2 >>
rect 134 328 135 329 
<< m1 >>
rect 135 328 136 329 
<< m2 >>
rect 135 328 136 329 
<< m1 >>
rect 136 328 137 329 
<< m2 >>
rect 136 328 137 329 
<< m1 >>
rect 137 328 138 329 
<< m2 >>
rect 137 328 138 329 
<< m1 >>
rect 138 328 139 329 
<< m2 >>
rect 138 328 139 329 
<< m1 >>
rect 139 328 140 329 
<< m2 >>
rect 139 328 140 329 
<< m1 >>
rect 140 328 141 329 
<< m2 >>
rect 140 328 141 329 
<< m1 >>
rect 141 328 142 329 
<< m2 >>
rect 141 328 142 329 
<< m1 >>
rect 142 328 143 329 
<< m2 >>
rect 142 328 143 329 
<< m1 >>
rect 143 328 144 329 
<< m2 >>
rect 143 328 144 329 
<< m1 >>
rect 144 328 145 329 
<< m2 >>
rect 144 328 145 329 
<< m1 >>
rect 145 328 146 329 
<< m2 >>
rect 145 328 146 329 
<< m1 >>
rect 146 328 147 329 
<< m2 >>
rect 146 328 147 329 
<< m1 >>
rect 147 328 148 329 
<< m2 >>
rect 147 328 148 329 
<< m1 >>
rect 148 328 149 329 
<< m2 >>
rect 148 328 149 329 
<< m1 >>
rect 149 328 150 329 
<< m2 >>
rect 149 328 150 329 
<< m1 >>
rect 150 328 151 329 
<< m2 >>
rect 150 328 151 329 
<< m1 >>
rect 151 328 152 329 
<< m2 >>
rect 151 328 152 329 
<< m1 >>
rect 152 328 153 329 
<< m2 >>
rect 152 328 153 329 
<< m1 >>
rect 153 328 154 329 
<< m2 >>
rect 153 328 154 329 
<< m1 >>
rect 154 328 155 329 
<< m2 >>
rect 154 328 155 329 
<< m1 >>
rect 155 328 156 329 
<< m2 >>
rect 155 328 156 329 
<< m1 >>
rect 156 328 157 329 
<< m2 >>
rect 156 328 157 329 
<< m1 >>
rect 157 328 158 329 
<< m2 >>
rect 157 328 158 329 
<< m1 >>
rect 158 328 159 329 
<< m2 >>
rect 158 328 159 329 
<< m1 >>
rect 159 328 160 329 
<< m1 >>
rect 160 328 161 329 
<< m1 >>
rect 161 328 162 329 
<< m1 >>
rect 162 328 163 329 
<< m1 >>
rect 163 328 164 329 
<< m1 >>
rect 164 328 165 329 
<< m1 >>
rect 165 328 166 329 
<< m1 >>
rect 166 328 167 329 
<< m1 >>
rect 167 328 168 329 
<< m1 >>
rect 168 328 169 329 
<< m1 >>
rect 169 328 170 329 
<< m1 >>
rect 170 328 171 329 
<< m1 >>
rect 171 328 172 329 
<< m1 >>
rect 172 328 173 329 
<< m1 >>
rect 173 328 174 329 
<< m1 >>
rect 174 328 175 329 
<< m1 >>
rect 175 328 176 329 
<< m1 >>
rect 176 328 177 329 
<< m1 >>
rect 177 328 178 329 
<< m1 >>
rect 178 328 179 329 
<< m1 >>
rect 179 328 180 329 
<< m1 >>
rect 180 328 181 329 
<< m1 >>
rect 181 328 182 329 
<< m1 >>
rect 182 328 183 329 
<< m1 >>
rect 183 328 184 329 
<< m1 >>
rect 184 328 185 329 
<< m1 >>
rect 185 328 186 329 
<< m1 >>
rect 186 328 187 329 
<< m1 >>
rect 187 328 188 329 
<< m1 >>
rect 188 328 189 329 
<< m1 >>
rect 189 328 190 329 
<< m1 >>
rect 190 328 191 329 
<< m1 >>
rect 191 328 192 329 
<< m1 >>
rect 192 328 193 329 
<< m1 >>
rect 193 328 194 329 
<< m1 >>
rect 194 328 195 329 
<< m2 >>
rect 194 328 195 329 
<< m1 >>
rect 195 328 196 329 
<< m1 >>
rect 196 328 197 329 
<< m1 >>
rect 197 328 198 329 
<< m1 >>
rect 198 328 199 329 
<< m1 >>
rect 199 328 200 329 
<< m1 >>
rect 200 328 201 329 
<< m1 >>
rect 201 328 202 329 
<< m1 >>
rect 202 328 203 329 
<< m1 >>
rect 203 328 204 329 
<< m1 >>
rect 204 328 205 329 
<< m1 >>
rect 205 328 206 329 
<< m1 >>
rect 206 328 207 329 
<< m1 >>
rect 207 328 208 329 
<< m1 >>
rect 208 328 209 329 
<< m1 >>
rect 209 328 210 329 
<< m1 >>
rect 210 328 211 329 
<< m1 >>
rect 211 328 212 329 
<< m1 >>
rect 212 328 213 329 
<< m1 >>
rect 213 328 214 329 
<< m1 >>
rect 214 328 215 329 
<< m1 >>
rect 215 328 216 329 
<< m1 >>
rect 216 328 217 329 
<< m1 >>
rect 217 328 218 329 
<< m2 >>
rect 217 328 218 329 
<< m1 >>
rect 218 328 219 329 
<< m1 >>
rect 219 328 220 329 
<< m2 >>
rect 219 328 220 329 
<< m1 >>
rect 220 328 221 329 
<< m1 >>
rect 221 328 222 329 
<< m2 >>
rect 221 328 222 329 
<< m1 >>
rect 222 328 223 329 
<< m1 >>
rect 223 328 224 329 
<< m2 >>
rect 223 328 224 329 
<< m1 >>
rect 224 328 225 329 
<< m1 >>
rect 225 328 226 329 
<< m1 >>
rect 226 328 227 329 
<< m1 >>
rect 227 328 228 329 
<< m1 >>
rect 228 328 229 329 
<< m1 >>
rect 229 328 230 329 
<< m1 >>
rect 230 328 231 329 
<< m1 >>
rect 231 328 232 329 
<< m1 >>
rect 232 328 233 329 
<< m1 >>
rect 233 328 234 329 
<< m1 >>
rect 234 328 235 329 
<< m1 >>
rect 235 328 236 329 
<< m1 >>
rect 236 328 237 329 
<< m1 >>
rect 237 328 238 329 
<< m1 >>
rect 238 328 239 329 
<< m1 >>
rect 239 328 240 329 
<< m2 >>
rect 239 328 240 329 
<< m1 >>
rect 240 328 241 329 
<< m1 >>
rect 241 328 242 329 
<< m1 >>
rect 242 328 243 329 
<< m1 >>
rect 243 328 244 329 
<< m1 >>
rect 244 328 245 329 
<< m1 >>
rect 245 328 246 329 
<< m1 >>
rect 246 328 247 329 
<< m1 >>
rect 247 328 248 329 
<< m1 >>
rect 248 328 249 329 
<< m1 >>
rect 249 328 250 329 
<< m1 >>
rect 250 328 251 329 
<< m1 >>
rect 251 328 252 329 
<< m2 >>
rect 251 328 252 329 
<< m2c >>
rect 251 328 252 329 
<< m1 >>
rect 251 328 252 329 
<< m2 >>
rect 251 328 252 329 
<< m2 >>
rect 252 328 253 329 
<< m1 >>
rect 253 328 254 329 
<< m1 >>
rect 254 328 255 329 
<< m1 >>
rect 255 328 256 329 
<< m1 >>
rect 256 328 257 329 
<< m1 >>
rect 257 328 258 329 
<< m1 >>
rect 258 328 259 329 
<< m1 >>
rect 259 328 260 329 
<< m1 >>
rect 260 328 261 329 
<< m1 >>
rect 261 328 262 329 
<< m1 >>
rect 262 328 263 329 
<< m1 >>
rect 263 328 264 329 
<< m1 >>
rect 264 328 265 329 
<< m1 >>
rect 265 328 266 329 
<< m1 >>
rect 266 328 267 329 
<< m1 >>
rect 267 328 268 329 
<< m1 >>
rect 268 328 269 329 
<< m2 >>
rect 268 328 269 329 
<< m1 >>
rect 269 328 270 329 
<< m1 >>
rect 270 328 271 329 
<< m1 >>
rect 271 328 272 329 
<< m2 >>
rect 271 328 272 329 
<< m1 >>
rect 272 328 273 329 
<< m1 >>
rect 273 328 274 329 
<< m2 >>
rect 273 328 274 329 
<< m1 >>
rect 274 328 275 329 
<< m1 >>
rect 275 328 276 329 
<< m2 >>
rect 275 328 276 329 
<< m1 >>
rect 276 328 277 329 
<< m2 >>
rect 276 328 277 329 
<< m1 >>
rect 277 328 278 329 
<< m2 >>
rect 277 328 278 329 
<< m1 >>
rect 278 328 279 329 
<< m2 >>
rect 278 328 279 329 
<< m1 >>
rect 279 328 280 329 
<< m2 >>
rect 279 328 280 329 
<< m1 >>
rect 280 328 281 329 
<< m2 >>
rect 280 328 281 329 
<< m1 >>
rect 281 328 282 329 
<< m2 >>
rect 281 328 282 329 
<< m1 >>
rect 282 328 283 329 
<< m2 >>
rect 282 328 283 329 
<< m1 >>
rect 283 328 284 329 
<< m2 >>
rect 283 328 284 329 
<< m1 >>
rect 284 328 285 329 
<< m2 >>
rect 284 328 285 329 
<< m1 >>
rect 285 328 286 329 
<< m2 >>
rect 285 328 286 329 
<< m1 >>
rect 286 328 287 329 
<< m2 >>
rect 286 328 287 329 
<< m1 >>
rect 287 328 288 329 
<< m2 >>
rect 287 328 288 329 
<< m1 >>
rect 288 328 289 329 
<< m2 >>
rect 288 328 289 329 
<< m1 >>
rect 289 328 290 329 
<< m2 >>
rect 289 328 290 329 
<< m1 >>
rect 290 328 291 329 
<< m2 >>
rect 290 328 291 329 
<< m1 >>
rect 291 328 292 329 
<< m2 >>
rect 291 328 292 329 
<< m1 >>
rect 292 328 293 329 
<< m2 >>
rect 292 328 293 329 
<< m1 >>
rect 293 328 294 329 
<< m2 >>
rect 293 328 294 329 
<< m1 >>
rect 294 328 295 329 
<< m2 >>
rect 294 328 295 329 
<< m1 >>
rect 295 328 296 329 
<< m2 >>
rect 295 328 296 329 
<< m1 >>
rect 296 328 297 329 
<< m2 >>
rect 296 328 297 329 
<< m1 >>
rect 297 328 298 329 
<< m2 >>
rect 297 328 298 329 
<< m1 >>
rect 298 328 299 329 
<< m2 >>
rect 298 328 299 329 
<< m1 >>
rect 299 328 300 329 
<< m2 >>
rect 299 328 300 329 
<< m1 >>
rect 300 328 301 329 
<< m2 >>
rect 300 328 301 329 
<< m1 >>
rect 301 328 302 329 
<< m2 >>
rect 301 328 302 329 
<< m1 >>
rect 302 328 303 329 
<< m2 >>
rect 302 328 303 329 
<< m1 >>
rect 303 328 304 329 
<< m2 >>
rect 303 328 304 329 
<< m1 >>
rect 304 328 305 329 
<< m2 >>
rect 304 328 305 329 
<< m1 >>
rect 305 328 306 329 
<< m2 >>
rect 305 328 306 329 
<< m1 >>
rect 306 328 307 329 
<< m2 >>
rect 306 328 307 329 
<< m1 >>
rect 307 328 308 329 
<< m2 >>
rect 307 328 308 329 
<< m1 >>
rect 308 328 309 329 
<< m2 >>
rect 308 328 309 329 
<< m1 >>
rect 309 328 310 329 
<< m2 >>
rect 309 328 310 329 
<< m1 >>
rect 310 328 311 329 
<< m2 >>
rect 310 328 311 329 
<< m1 >>
rect 311 328 312 329 
<< m2 >>
rect 311 328 312 329 
<< m1 >>
rect 312 328 313 329 
<< m2 >>
rect 312 328 313 329 
<< m1 >>
rect 313 328 314 329 
<< m2 >>
rect 313 328 314 329 
<< m1 >>
rect 314 328 315 329 
<< m2 >>
rect 314 328 315 329 
<< m1 >>
rect 315 328 316 329 
<< m2 >>
rect 315 328 316 329 
<< m1 >>
rect 316 328 317 329 
<< m2 >>
rect 316 328 317 329 
<< m1 >>
rect 317 328 318 329 
<< m2 >>
rect 317 328 318 329 
<< m1 >>
rect 318 328 319 329 
<< m2 >>
rect 318 328 319 329 
<< m1 >>
rect 319 328 320 329 
<< m2 >>
rect 319 328 320 329 
<< m2 >>
rect 320 328 321 329 
<< m1 >>
rect 321 328 322 329 
<< m2 >>
rect 321 328 322 329 
<< m2c >>
rect 321 328 322 329 
<< m1 >>
rect 321 328 322 329 
<< m2 >>
rect 321 328 322 329 
<< m1 >>
rect 322 328 323 329 
<< m1 >>
rect 323 328 324 329 
<< m2 >>
rect 323 328 324 329 
<< m1 >>
rect 324 328 325 329 
<< m1 >>
rect 325 328 326 329 
<< m2 >>
rect 325 328 326 329 
<< m1 >>
rect 326 328 327 329 
<< m1 >>
rect 327 328 328 329 
<< m1 >>
rect 328 328 329 329 
<< m1 >>
rect 329 328 330 329 
<< m2 >>
rect 329 328 330 329 
<< m1 >>
rect 330 328 331 329 
<< m1 >>
rect 331 328 332 329 
<< m2 >>
rect 331 328 332 329 
<< m1 >>
rect 332 328 333 329 
<< m1 >>
rect 333 328 334 329 
<< m1 >>
rect 334 328 335 329 
<< m2 >>
rect 334 328 335 329 
<< m1 >>
rect 335 328 336 329 
<< m1 >>
rect 336 328 337 329 
<< m1 >>
rect 337 328 338 329 
<< m1 >>
rect 338 328 339 329 
<< m1 >>
rect 339 328 340 329 
<< m1 >>
rect 340 328 341 329 
<< m2 >>
rect 340 328 341 329 
<< m1 >>
rect 343 328 344 329 
<< m1 >>
rect 10 329 11 330 
<< m1 >>
rect 26 329 27 330 
<< m1 >>
rect 28 329 29 330 
<< m2 >>
rect 38 329 39 330 
<< m2 >>
rect 39 329 40 330 
<< m2 >>
rect 40 329 41 330 
<< m2 >>
rect 41 329 42 330 
<< m2 >>
rect 42 329 43 330 
<< m2 >>
rect 43 329 44 330 
<< m2 >>
rect 44 329 45 330 
<< m2 >>
rect 45 329 46 330 
<< m2 >>
rect 46 329 47 330 
<< m2 >>
rect 48 329 49 330 
<< m1 >>
rect 49 329 50 330 
<< m1 >>
rect 52 329 53 330 
<< m1 >>
rect 56 329 57 330 
<< m1 >>
rect 57 329 58 330 
<< m1 >>
rect 60 329 61 330 
<< m1 >>
rect 62 329 63 330 
<< m2 >>
rect 102 329 103 330 
<< m2 >>
rect 103 329 104 330 
<< m2 >>
rect 104 329 105 330 
<< m2 >>
rect 105 329 106 330 
<< m2 >>
rect 106 329 107 330 
<< m2 >>
rect 107 329 108 330 
<< m2 >>
rect 108 329 109 330 
<< m2 >>
rect 109 329 110 330 
<< m2 >>
rect 110 329 111 330 
<< m2 >>
rect 111 329 112 330 
<< m2 >>
rect 112 329 113 330 
<< m2 >>
rect 113 329 114 330 
<< m2 >>
rect 114 329 115 330 
<< m2 >>
rect 115 329 116 330 
<< m2 >>
rect 116 329 117 330 
<< m2 >>
rect 117 329 118 330 
<< m2 >>
rect 194 329 195 330 
<< m2 >>
rect 217 329 218 330 
<< m2 >>
rect 219 329 220 330 
<< m2 >>
rect 221 329 222 330 
<< m2 >>
rect 223 329 224 330 
<< m2 >>
rect 239 329 240 330 
<< m2 >>
rect 268 329 269 330 
<< m2 >>
rect 271 329 272 330 
<< m2 >>
rect 273 329 274 330 
<< m1 >>
rect 319 329 320 330 
<< m2 >>
rect 323 329 324 330 
<< m2 >>
rect 325 329 326 330 
<< m2 >>
rect 329 329 330 330 
<< m2 >>
rect 331 329 332 330 
<< m2 >>
rect 334 329 335 330 
<< m1 >>
rect 340 329 341 330 
<< m2 >>
rect 340 329 341 330 
<< m1 >>
rect 343 329 344 330 
<< m1 >>
rect 10 330 11 331 
<< m1 >>
rect 26 330 27 331 
<< m1 >>
rect 28 330 29 331 
<< m1 >>
rect 46 330 47 331 
<< m2 >>
rect 46 330 47 331 
<< m2c >>
rect 46 330 47 331 
<< m1 >>
rect 46 330 47 331 
<< m2 >>
rect 46 330 47 331 
<< m2 >>
rect 48 330 49 331 
<< m1 >>
rect 49 330 50 331 
<< m1 >>
rect 52 330 53 331 
<< m1 >>
rect 56 330 57 331 
<< m1 >>
rect 60 330 61 331 
<< m1 >>
rect 62 330 63 331 
<< m1 >>
rect 117 330 118 331 
<< m2 >>
rect 117 330 118 331 
<< m2c >>
rect 117 330 118 331 
<< m1 >>
rect 117 330 118 331 
<< m2 >>
rect 117 330 118 331 
<< m1 >>
rect 118 330 119 331 
<< m1 >>
rect 119 330 120 331 
<< m1 >>
rect 120 330 121 331 
<< m1 >>
rect 121 330 122 331 
<< m1 >>
rect 122 330 123 331 
<< m1 >>
rect 123 330 124 331 
<< m1 >>
rect 124 330 125 331 
<< m1 >>
rect 125 330 126 331 
<< m1 >>
rect 126 330 127 331 
<< m1 >>
rect 127 330 128 331 
<< m1 >>
rect 128 330 129 331 
<< m1 >>
rect 129 330 130 331 
<< m1 >>
rect 130 330 131 331 
<< m1 >>
rect 131 330 132 331 
<< m1 >>
rect 132 330 133 331 
<< m1 >>
rect 133 330 134 331 
<< m1 >>
rect 134 330 135 331 
<< m1 >>
rect 135 330 136 331 
<< m1 >>
rect 136 330 137 331 
<< m1 >>
rect 137 330 138 331 
<< m1 >>
rect 138 330 139 331 
<< m1 >>
rect 139 330 140 331 
<< m1 >>
rect 140 330 141 331 
<< m1 >>
rect 141 330 142 331 
<< m1 >>
rect 142 330 143 331 
<< m1 >>
rect 143 330 144 331 
<< m1 >>
rect 144 330 145 331 
<< m1 >>
rect 145 330 146 331 
<< m1 >>
rect 146 330 147 331 
<< m1 >>
rect 147 330 148 331 
<< m1 >>
rect 148 330 149 331 
<< m1 >>
rect 149 330 150 331 
<< m1 >>
rect 150 330 151 331 
<< m1 >>
rect 151 330 152 331 
<< m1 >>
rect 152 330 153 331 
<< m1 >>
rect 153 330 154 331 
<< m1 >>
rect 154 330 155 331 
<< m1 >>
rect 155 330 156 331 
<< m1 >>
rect 156 330 157 331 
<< m1 >>
rect 157 330 158 331 
<< m1 >>
rect 158 330 159 331 
<< m1 >>
rect 159 330 160 331 
<< m1 >>
rect 160 330 161 331 
<< m1 >>
rect 161 330 162 331 
<< m1 >>
rect 162 330 163 331 
<< m1 >>
rect 163 330 164 331 
<< m1 >>
rect 164 330 165 331 
<< m1 >>
rect 165 330 166 331 
<< m1 >>
rect 166 330 167 331 
<< m1 >>
rect 167 330 168 331 
<< m1 >>
rect 168 330 169 331 
<< m1 >>
rect 169 330 170 331 
<< m1 >>
rect 170 330 171 331 
<< m1 >>
rect 171 330 172 331 
<< m1 >>
rect 172 330 173 331 
<< m1 >>
rect 173 330 174 331 
<< m1 >>
rect 174 330 175 331 
<< m1 >>
rect 175 330 176 331 
<< m1 >>
rect 176 330 177 331 
<< m1 >>
rect 177 330 178 331 
<< m1 >>
rect 178 330 179 331 
<< m1 >>
rect 179 330 180 331 
<< m1 >>
rect 180 330 181 331 
<< m1 >>
rect 181 330 182 331 
<< m1 >>
rect 182 330 183 331 
<< m1 >>
rect 183 330 184 331 
<< m1 >>
rect 184 330 185 331 
<< m1 >>
rect 185 330 186 331 
<< m1 >>
rect 186 330 187 331 
<< m1 >>
rect 187 330 188 331 
<< m1 >>
rect 188 330 189 331 
<< m1 >>
rect 189 330 190 331 
<< m1 >>
rect 190 330 191 331 
<< m1 >>
rect 191 330 192 331 
<< m1 >>
rect 192 330 193 331 
<< m1 >>
rect 193 330 194 331 
<< m1 >>
rect 194 330 195 331 
<< m2 >>
rect 194 330 195 331 
<< m1 >>
rect 195 330 196 331 
<< m1 >>
rect 196 330 197 331 
<< m1 >>
rect 197 330 198 331 
<< m1 >>
rect 198 330 199 331 
<< m1 >>
rect 199 330 200 331 
<< m1 >>
rect 200 330 201 331 
<< m1 >>
rect 201 330 202 331 
<< m1 >>
rect 202 330 203 331 
<< m1 >>
rect 203 330 204 331 
<< m1 >>
rect 204 330 205 331 
<< m1 >>
rect 205 330 206 331 
<< m1 >>
rect 206 330 207 331 
<< m1 >>
rect 207 330 208 331 
<< m1 >>
rect 208 330 209 331 
<< m1 >>
rect 209 330 210 331 
<< m1 >>
rect 210 330 211 331 
<< m1 >>
rect 211 330 212 331 
<< m1 >>
rect 212 330 213 331 
<< m1 >>
rect 213 330 214 331 
<< m1 >>
rect 214 330 215 331 
<< m1 >>
rect 215 330 216 331 
<< m1 >>
rect 216 330 217 331 
<< m1 >>
rect 217 330 218 331 
<< m2 >>
rect 217 330 218 331 
<< m2c >>
rect 217 330 218 331 
<< m1 >>
rect 217 330 218 331 
<< m2 >>
rect 217 330 218 331 
<< m1 >>
rect 219 330 220 331 
<< m2 >>
rect 219 330 220 331 
<< m2c >>
rect 219 330 220 331 
<< m1 >>
rect 219 330 220 331 
<< m2 >>
rect 219 330 220 331 
<< m1 >>
rect 221 330 222 331 
<< m2 >>
rect 221 330 222 331 
<< m2c >>
rect 221 330 222 331 
<< m1 >>
rect 221 330 222 331 
<< m2 >>
rect 221 330 222 331 
<< m1 >>
rect 223 330 224 331 
<< m2 >>
rect 223 330 224 331 
<< m2c >>
rect 223 330 224 331 
<< m1 >>
rect 223 330 224 331 
<< m2 >>
rect 223 330 224 331 
<< m1 >>
rect 239 330 240 331 
<< m2 >>
rect 239 330 240 331 
<< m2c >>
rect 239 330 240 331 
<< m1 >>
rect 239 330 240 331 
<< m2 >>
rect 239 330 240 331 
<< m1 >>
rect 268 330 269 331 
<< m2 >>
rect 268 330 269 331 
<< m2c >>
rect 268 330 269 331 
<< m1 >>
rect 268 330 269 331 
<< m2 >>
rect 268 330 269 331 
<< m1 >>
rect 271 330 272 331 
<< m2 >>
rect 271 330 272 331 
<< m2c >>
rect 271 330 272 331 
<< m1 >>
rect 271 330 272 331 
<< m2 >>
rect 271 330 272 331 
<< m1 >>
rect 273 330 274 331 
<< m2 >>
rect 273 330 274 331 
<< m2c >>
rect 273 330 274 331 
<< m1 >>
rect 273 330 274 331 
<< m2 >>
rect 273 330 274 331 
<< m1 >>
rect 319 330 320 331 
<< m1 >>
rect 323 330 324 331 
<< m2 >>
rect 323 330 324 331 
<< m2c >>
rect 323 330 324 331 
<< m1 >>
rect 323 330 324 331 
<< m2 >>
rect 323 330 324 331 
<< m1 >>
rect 325 330 326 331 
<< m2 >>
rect 325 330 326 331 
<< m2c >>
rect 325 330 326 331 
<< m1 >>
rect 325 330 326 331 
<< m2 >>
rect 325 330 326 331 
<< m1 >>
rect 329 330 330 331 
<< m2 >>
rect 329 330 330 331 
<< m2c >>
rect 329 330 330 331 
<< m1 >>
rect 329 330 330 331 
<< m2 >>
rect 329 330 330 331 
<< m1 >>
rect 331 330 332 331 
<< m2 >>
rect 331 330 332 331 
<< m2c >>
rect 331 330 332 331 
<< m1 >>
rect 331 330 332 331 
<< m2 >>
rect 331 330 332 331 
<< m1 >>
rect 334 330 335 331 
<< m2 >>
rect 334 330 335 331 
<< m2c >>
rect 334 330 335 331 
<< m1 >>
rect 334 330 335 331 
<< m2 >>
rect 334 330 335 331 
<< m1 >>
rect 336 330 337 331 
<< m1 >>
rect 337 330 338 331 
<< m1 >>
rect 338 330 339 331 
<< m2 >>
rect 338 330 339 331 
<< m2c >>
rect 338 330 339 331 
<< m1 >>
rect 338 330 339 331 
<< m2 >>
rect 338 330 339 331 
<< m2 >>
rect 339 330 340 331 
<< m1 >>
rect 340 330 341 331 
<< m2 >>
rect 340 330 341 331 
<< m1 >>
rect 343 330 344 331 
<< m1 >>
rect 10 331 11 332 
<< m1 >>
rect 26 331 27 332 
<< m1 >>
rect 28 331 29 332 
<< m1 >>
rect 46 331 47 332 
<< m2 >>
rect 48 331 49 332 
<< m1 >>
rect 49 331 50 332 
<< m1 >>
rect 52 331 53 332 
<< m1 >>
rect 56 331 57 332 
<< m1 >>
rect 58 331 59 332 
<< m2 >>
rect 58 331 59 332 
<< m2c >>
rect 58 331 59 332 
<< m1 >>
rect 58 331 59 332 
<< m2 >>
rect 58 331 59 332 
<< m2 >>
rect 59 331 60 332 
<< m1 >>
rect 60 331 61 332 
<< m2 >>
rect 60 331 61 332 
<< m2 >>
rect 61 331 62 332 
<< m1 >>
rect 62 331 63 332 
<< m2 >>
rect 62 331 63 332 
<< m2 >>
rect 63 331 64 332 
<< m1 >>
rect 64 331 65 332 
<< m2 >>
rect 64 331 65 332 
<< m2c >>
rect 64 331 65 332 
<< m1 >>
rect 64 331 65 332 
<< m2 >>
rect 64 331 65 332 
<< m1 >>
rect 65 331 66 332 
<< m1 >>
rect 66 331 67 332 
<< m1 >>
rect 67 331 68 332 
<< m1 >>
rect 68 331 69 332 
<< m1 >>
rect 69 331 70 332 
<< m1 >>
rect 70 331 71 332 
<< m1 >>
rect 71 331 72 332 
<< m1 >>
rect 72 331 73 332 
<< m1 >>
rect 73 331 74 332 
<< m1 >>
rect 74 331 75 332 
<< m1 >>
rect 75 331 76 332 
<< m1 >>
rect 76 331 77 332 
<< m1 >>
rect 77 331 78 332 
<< m1 >>
rect 78 331 79 332 
<< m1 >>
rect 79 331 80 332 
<< m1 >>
rect 80 331 81 332 
<< m1 >>
rect 81 331 82 332 
<< m1 >>
rect 82 331 83 332 
<< m1 >>
rect 83 331 84 332 
<< m1 >>
rect 84 331 85 332 
<< m1 >>
rect 85 331 86 332 
<< m1 >>
rect 86 331 87 332 
<< m1 >>
rect 87 331 88 332 
<< m1 >>
rect 88 331 89 332 
<< m1 >>
rect 89 331 90 332 
<< m1 >>
rect 90 331 91 332 
<< m1 >>
rect 91 331 92 332 
<< m1 >>
rect 92 331 93 332 
<< m1 >>
rect 93 331 94 332 
<< m1 >>
rect 94 331 95 332 
<< m1 >>
rect 95 331 96 332 
<< m1 >>
rect 96 331 97 332 
<< m1 >>
rect 97 331 98 332 
<< m1 >>
rect 98 331 99 332 
<< m1 >>
rect 99 331 100 332 
<< m1 >>
rect 100 331 101 332 
<< m1 >>
rect 101 331 102 332 
<< m1 >>
rect 102 331 103 332 
<< m1 >>
rect 103 331 104 332 
<< m1 >>
rect 104 331 105 332 
<< m1 >>
rect 105 331 106 332 
<< m1 >>
rect 106 331 107 332 
<< m1 >>
rect 107 331 108 332 
<< m1 >>
rect 108 331 109 332 
<< m1 >>
rect 109 331 110 332 
<< m1 >>
rect 110 331 111 332 
<< m1 >>
rect 111 331 112 332 
<< m1 >>
rect 112 331 113 332 
<< m1 >>
rect 113 331 114 332 
<< m1 >>
rect 114 331 115 332 
<< m1 >>
rect 115 331 116 332 
<< m2 >>
rect 115 331 116 332 
<< m2c >>
rect 115 331 116 332 
<< m1 >>
rect 115 331 116 332 
<< m2 >>
rect 115 331 116 332 
<< m2 >>
rect 119 331 120 332 
<< m2 >>
rect 120 331 121 332 
<< m2 >>
rect 121 331 122 332 
<< m2 >>
rect 122 331 123 332 
<< m2 >>
rect 123 331 124 332 
<< m2 >>
rect 124 331 125 332 
<< m2 >>
rect 125 331 126 332 
<< m2 >>
rect 126 331 127 332 
<< m2 >>
rect 127 331 128 332 
<< m2 >>
rect 128 331 129 332 
<< m2 >>
rect 129 331 130 332 
<< m2 >>
rect 130 331 131 332 
<< m2 >>
rect 131 331 132 332 
<< m2 >>
rect 132 331 133 332 
<< m2 >>
rect 133 331 134 332 
<< m2 >>
rect 134 331 135 332 
<< m2 >>
rect 135 331 136 332 
<< m2 >>
rect 136 331 137 332 
<< m2 >>
rect 137 331 138 332 
<< m2 >>
rect 138 331 139 332 
<< m2 >>
rect 139 331 140 332 
<< m2 >>
rect 140 331 141 332 
<< m2 >>
rect 141 331 142 332 
<< m2 >>
rect 142 331 143 332 
<< m2 >>
rect 143 331 144 332 
<< m2 >>
rect 144 331 145 332 
<< m2 >>
rect 145 331 146 332 
<< m2 >>
rect 146 331 147 332 
<< m2 >>
rect 147 331 148 332 
<< m2 >>
rect 148 331 149 332 
<< m2 >>
rect 149 331 150 332 
<< m2 >>
rect 150 331 151 332 
<< m2 >>
rect 151 331 152 332 
<< m2 >>
rect 152 331 153 332 
<< m2 >>
rect 153 331 154 332 
<< m2 >>
rect 154 331 155 332 
<< m2 >>
rect 155 331 156 332 
<< m2 >>
rect 156 331 157 332 
<< m2 >>
rect 157 331 158 332 
<< m2 >>
rect 158 331 159 332 
<< m2 >>
rect 159 331 160 332 
<< m2 >>
rect 160 331 161 332 
<< m2 >>
rect 161 331 162 332 
<< m2 >>
rect 162 331 163 332 
<< m2 >>
rect 163 331 164 332 
<< m2 >>
rect 164 331 165 332 
<< m2 >>
rect 165 331 166 332 
<< m2 >>
rect 166 331 167 332 
<< m2 >>
rect 167 331 168 332 
<< m2 >>
rect 168 331 169 332 
<< m2 >>
rect 169 331 170 332 
<< m2 >>
rect 170 331 171 332 
<< m2 >>
rect 171 331 172 332 
<< m2 >>
rect 172 331 173 332 
<< m2 >>
rect 173 331 174 332 
<< m2 >>
rect 174 331 175 332 
<< m2 >>
rect 175 331 176 332 
<< m2 >>
rect 176 331 177 332 
<< m2 >>
rect 177 331 178 332 
<< m2 >>
rect 178 331 179 332 
<< m2 >>
rect 179 331 180 332 
<< m2 >>
rect 180 331 181 332 
<< m2 >>
rect 181 331 182 332 
<< m2 >>
rect 182 331 183 332 
<< m2 >>
rect 183 331 184 332 
<< m2 >>
rect 184 331 185 332 
<< m2 >>
rect 185 331 186 332 
<< m2 >>
rect 186 331 187 332 
<< m2 >>
rect 187 331 188 332 
<< m2 >>
rect 188 331 189 332 
<< m2 >>
rect 189 331 190 332 
<< m2 >>
rect 190 331 191 332 
<< m2 >>
rect 191 331 192 332 
<< m2 >>
rect 192 331 193 332 
<< m2 >>
rect 193 331 194 332 
<< m2 >>
rect 194 331 195 332 
<< m1 >>
rect 219 331 220 332 
<< m1 >>
rect 221 331 222 332 
<< m1 >>
rect 223 331 224 332 
<< m1 >>
rect 239 331 240 332 
<< m1 >>
rect 268 331 269 332 
<< m1 >>
rect 271 331 272 332 
<< m1 >>
rect 273 331 274 332 
<< m2 >>
rect 318 331 319 332 
<< m1 >>
rect 319 331 320 332 
<< m2 >>
rect 319 331 320 332 
<< m2 >>
rect 320 331 321 332 
<< m1 >>
rect 321 331 322 332 
<< m2 >>
rect 321 331 322 332 
<< m2c >>
rect 321 331 322 332 
<< m1 >>
rect 321 331 322 332 
<< m2 >>
rect 321 331 322 332 
<< m1 >>
rect 322 331 323 332 
<< m1 >>
rect 323 331 324 332 
<< m1 >>
rect 325 331 326 332 
<< m1 >>
rect 329 331 330 332 
<< m1 >>
rect 331 331 332 332 
<< m1 >>
rect 334 331 335 332 
<< m1 >>
rect 336 331 337 332 
<< m1 >>
rect 340 331 341 332 
<< m1 >>
rect 343 331 344 332 
<< m1 >>
rect 10 332 11 333 
<< m1 >>
rect 26 332 27 333 
<< m1 >>
rect 28 332 29 333 
<< m1 >>
rect 46 332 47 333 
<< m2 >>
rect 48 332 49 333 
<< m1 >>
rect 49 332 50 333 
<< m1 >>
rect 52 332 53 333 
<< m1 >>
rect 56 332 57 333 
<< m1 >>
rect 58 332 59 333 
<< m1 >>
rect 60 332 61 333 
<< m1 >>
rect 62 332 63 333 
<< m2 >>
rect 115 332 116 333 
<< m1 >>
rect 119 332 120 333 
<< m2 >>
rect 119 332 120 333 
<< m2c >>
rect 119 332 120 333 
<< m1 >>
rect 119 332 120 333 
<< m2 >>
rect 119 332 120 333 
<< m1 >>
rect 219 332 220 333 
<< m1 >>
rect 221 332 222 333 
<< m1 >>
rect 223 332 224 333 
<< m1 >>
rect 239 332 240 333 
<< m1 >>
rect 268 332 269 333 
<< m1 >>
rect 269 332 270 333 
<< m2 >>
rect 269 332 270 333 
<< m2c >>
rect 269 332 270 333 
<< m1 >>
rect 269 332 270 333 
<< m2 >>
rect 269 332 270 333 
<< m2 >>
rect 270 332 271 333 
<< m1 >>
rect 271 332 272 333 
<< m2 >>
rect 271 332 272 333 
<< m2 >>
rect 272 332 273 333 
<< m1 >>
rect 273 332 274 333 
<< m2 >>
rect 273 332 274 333 
<< m2c >>
rect 273 332 274 333 
<< m1 >>
rect 273 332 274 333 
<< m2 >>
rect 273 332 274 333 
<< m2 >>
rect 318 332 319 333 
<< m1 >>
rect 319 332 320 333 
<< m1 >>
rect 325 332 326 333 
<< m2 >>
rect 326 332 327 333 
<< m1 >>
rect 327 332 328 333 
<< m2 >>
rect 327 332 328 333 
<< m2c >>
rect 327 332 328 333 
<< m1 >>
rect 327 332 328 333 
<< m2 >>
rect 327 332 328 333 
<< m1 >>
rect 328 332 329 333 
<< m1 >>
rect 329 332 330 333 
<< m1 >>
rect 331 332 332 333 
<< m2 >>
rect 332 332 333 333 
<< m1 >>
rect 333 332 334 333 
<< m2 >>
rect 333 332 334 333 
<< m2c >>
rect 333 332 334 333 
<< m1 >>
rect 333 332 334 333 
<< m2 >>
rect 333 332 334 333 
<< m1 >>
rect 334 332 335 333 
<< m1 >>
rect 336 332 337 333 
<< m1 >>
rect 340 332 341 333 
<< m1 >>
rect 343 332 344 333 
<< m1 >>
rect 10 333 11 334 
<< m1 >>
rect 26 333 27 334 
<< m1 >>
rect 28 333 29 334 
<< m1 >>
rect 46 333 47 334 
<< m2 >>
rect 48 333 49 334 
<< m1 >>
rect 49 333 50 334 
<< m1 >>
rect 52 333 53 334 
<< m1 >>
rect 56 333 57 334 
<< m1 >>
rect 58 333 59 334 
<< m1 >>
rect 60 333 61 334 
<< m1 >>
rect 62 333 63 334 
<< m1 >>
rect 103 333 104 334 
<< m1 >>
rect 104 333 105 334 
<< m1 >>
rect 105 333 106 334 
<< m1 >>
rect 106 333 107 334 
<< m1 >>
rect 107 333 108 334 
<< m1 >>
rect 108 333 109 334 
<< m1 >>
rect 109 333 110 334 
<< m1 >>
rect 110 333 111 334 
<< m1 >>
rect 111 333 112 334 
<< m1 >>
rect 112 333 113 334 
<< m1 >>
rect 113 333 114 334 
<< m1 >>
rect 114 333 115 334 
<< m1 >>
rect 115 333 116 334 
<< m2 >>
rect 115 333 116 334 
<< m1 >>
rect 116 333 117 334 
<< m1 >>
rect 117 333 118 334 
<< m1 >>
rect 118 333 119 334 
<< m1 >>
rect 119 333 120 334 
<< m1 >>
rect 219 333 220 334 
<< m1 >>
rect 221 333 222 334 
<< m1 >>
rect 223 333 224 334 
<< m1 >>
rect 239 333 240 334 
<< m1 >>
rect 271 333 272 334 
<< m2 >>
rect 318 333 319 334 
<< m1 >>
rect 319 333 320 334 
<< m1 >>
rect 325 333 326 334 
<< m2 >>
rect 326 333 327 334 
<< m1 >>
rect 331 333 332 334 
<< m2 >>
rect 332 333 333 334 
<< m1 >>
rect 336 333 337 334 
<< m1 >>
rect 340 333 341 334 
<< m1 >>
rect 343 333 344 334 
<< m1 >>
rect 10 334 11 335 
<< m1 >>
rect 26 334 27 335 
<< m1 >>
rect 28 334 29 335 
<< m1 >>
rect 46 334 47 335 
<< m2 >>
rect 46 334 47 335 
<< m2 >>
rect 47 334 48 335 
<< m2 >>
rect 48 334 49 335 
<< m1 >>
rect 49 334 50 335 
<< m1 >>
rect 52 334 53 335 
<< m1 >>
rect 56 334 57 335 
<< m1 >>
rect 58 334 59 335 
<< m1 >>
rect 60 334 61 335 
<< m1 >>
rect 62 334 63 335 
<< m1 >>
rect 103 334 104 335 
<< m2 >>
rect 115 334 116 335 
<< m2 >>
rect 116 334 117 335 
<< m2 >>
rect 117 334 118 335 
<< m2 >>
rect 118 334 119 335 
<< m1 >>
rect 142 334 143 335 
<< m1 >>
rect 143 334 144 335 
<< m1 >>
rect 144 334 145 335 
<< m1 >>
rect 145 334 146 335 
<< m1 >>
rect 219 334 220 335 
<< m1 >>
rect 221 334 222 335 
<< m1 >>
rect 223 334 224 335 
<< m1 >>
rect 239 334 240 335 
<< m1 >>
rect 271 334 272 335 
<< m1 >>
rect 307 334 308 335 
<< m1 >>
rect 308 334 309 335 
<< m1 >>
rect 309 334 310 335 
<< m1 >>
rect 310 334 311 335 
<< m1 >>
rect 311 334 312 335 
<< m1 >>
rect 312 334 313 335 
<< m1 >>
rect 313 334 314 335 
<< m1 >>
rect 314 334 315 335 
<< m1 >>
rect 315 334 316 335 
<< m1 >>
rect 316 334 317 335 
<< m1 >>
rect 317 334 318 335 
<< m2 >>
rect 317 334 318 335 
<< m2c >>
rect 317 334 318 335 
<< m1 >>
rect 317 334 318 335 
<< m2 >>
rect 317 334 318 335 
<< m2 >>
rect 318 334 319 335 
<< m1 >>
rect 319 334 320 335 
<< m1 >>
rect 325 334 326 335 
<< m2 >>
rect 326 334 327 335 
<< m1 >>
rect 331 334 332 335 
<< m2 >>
rect 332 334 333 335 
<< m1 >>
rect 334 334 335 335 
<< m1 >>
rect 335 334 336 335 
<< m1 >>
rect 336 334 337 335 
<< m1 >>
rect 340 334 341 335 
<< m1 >>
rect 343 334 344 335 
<< m1 >>
rect 10 335 11 336 
<< m1 >>
rect 26 335 27 336 
<< m1 >>
rect 28 335 29 336 
<< m1 >>
rect 46 335 47 336 
<< m2 >>
rect 46 335 47 336 
<< m1 >>
rect 49 335 50 336 
<< m1 >>
rect 52 335 53 336 
<< m1 >>
rect 56 335 57 336 
<< m1 >>
rect 58 335 59 336 
<< m1 >>
rect 60 335 61 336 
<< m1 >>
rect 62 335 63 336 
<< m1 >>
rect 103 335 104 336 
<< m1 >>
rect 118 335 119 336 
<< m2 >>
rect 118 335 119 336 
<< m2c >>
rect 118 335 119 336 
<< m1 >>
rect 118 335 119 336 
<< m2 >>
rect 118 335 119 336 
<< m1 >>
rect 142 335 143 336 
<< m1 >>
rect 145 335 146 336 
<< m1 >>
rect 219 335 220 336 
<< m1 >>
rect 221 335 222 336 
<< m1 >>
rect 223 335 224 336 
<< m1 >>
rect 239 335 240 336 
<< m1 >>
rect 271 335 272 336 
<< m1 >>
rect 307 335 308 336 
<< m1 >>
rect 319 335 320 336 
<< m1 >>
rect 325 335 326 336 
<< m2 >>
rect 326 335 327 336 
<< m1 >>
rect 331 335 332 336 
<< m2 >>
rect 332 335 333 336 
<< m1 >>
rect 334 335 335 336 
<< m1 >>
rect 340 335 341 336 
<< m1 >>
rect 343 335 344 336 
<< m1 >>
rect 10 336 11 337 
<< pdiffusion >>
rect 12 336 13 337 
<< pdiffusion >>
rect 13 336 14 337 
<< pdiffusion >>
rect 14 336 15 337 
<< pdiffusion >>
rect 15 336 16 337 
<< pdiffusion >>
rect 16 336 17 337 
<< pdiffusion >>
rect 17 336 18 337 
<< m1 >>
rect 26 336 27 337 
<< m1 >>
rect 28 336 29 337 
<< pdiffusion >>
rect 30 336 31 337 
<< pdiffusion >>
rect 31 336 32 337 
<< pdiffusion >>
rect 32 336 33 337 
<< pdiffusion >>
rect 33 336 34 337 
<< pdiffusion >>
rect 34 336 35 337 
<< pdiffusion >>
rect 35 336 36 337 
<< m1 >>
rect 46 336 47 337 
<< m2 >>
rect 46 336 47 337 
<< pdiffusion >>
rect 48 336 49 337 
<< m1 >>
rect 49 336 50 337 
<< pdiffusion >>
rect 49 336 50 337 
<< pdiffusion >>
rect 50 336 51 337 
<< pdiffusion >>
rect 51 336 52 337 
<< m1 >>
rect 52 336 53 337 
<< pdiffusion >>
rect 52 336 53 337 
<< pdiffusion >>
rect 53 336 54 337 
<< m1 >>
rect 56 336 57 337 
<< m1 >>
rect 58 336 59 337 
<< m1 >>
rect 60 336 61 337 
<< m1 >>
rect 62 336 63 337 
<< pdiffusion >>
rect 66 336 67 337 
<< pdiffusion >>
rect 67 336 68 337 
<< pdiffusion >>
rect 68 336 69 337 
<< pdiffusion >>
rect 69 336 70 337 
<< pdiffusion >>
rect 70 336 71 337 
<< pdiffusion >>
rect 71 336 72 337 
<< pdiffusion >>
rect 84 336 85 337 
<< pdiffusion >>
rect 85 336 86 337 
<< pdiffusion >>
rect 86 336 87 337 
<< pdiffusion >>
rect 87 336 88 337 
<< pdiffusion >>
rect 88 336 89 337 
<< pdiffusion >>
rect 89 336 90 337 
<< pdiffusion >>
rect 102 336 103 337 
<< m1 >>
rect 103 336 104 337 
<< pdiffusion >>
rect 103 336 104 337 
<< pdiffusion >>
rect 104 336 105 337 
<< pdiffusion >>
rect 105 336 106 337 
<< pdiffusion >>
rect 106 336 107 337 
<< pdiffusion >>
rect 107 336 108 337 
<< m1 >>
rect 118 336 119 337 
<< pdiffusion >>
rect 120 336 121 337 
<< pdiffusion >>
rect 121 336 122 337 
<< pdiffusion >>
rect 122 336 123 337 
<< pdiffusion >>
rect 123 336 124 337 
<< pdiffusion >>
rect 124 336 125 337 
<< pdiffusion >>
rect 125 336 126 337 
<< pdiffusion >>
rect 138 336 139 337 
<< pdiffusion >>
rect 139 336 140 337 
<< pdiffusion >>
rect 140 336 141 337 
<< pdiffusion >>
rect 141 336 142 337 
<< m1 >>
rect 142 336 143 337 
<< pdiffusion >>
rect 142 336 143 337 
<< pdiffusion >>
rect 143 336 144 337 
<< m1 >>
rect 145 336 146 337 
<< pdiffusion >>
rect 156 336 157 337 
<< pdiffusion >>
rect 157 336 158 337 
<< pdiffusion >>
rect 158 336 159 337 
<< pdiffusion >>
rect 159 336 160 337 
<< pdiffusion >>
rect 160 336 161 337 
<< pdiffusion >>
rect 161 336 162 337 
<< pdiffusion >>
rect 174 336 175 337 
<< pdiffusion >>
rect 175 336 176 337 
<< pdiffusion >>
rect 176 336 177 337 
<< pdiffusion >>
rect 177 336 178 337 
<< pdiffusion >>
rect 178 336 179 337 
<< pdiffusion >>
rect 179 336 180 337 
<< pdiffusion >>
rect 192 336 193 337 
<< pdiffusion >>
rect 193 336 194 337 
<< pdiffusion >>
rect 194 336 195 337 
<< pdiffusion >>
rect 195 336 196 337 
<< pdiffusion >>
rect 196 336 197 337 
<< pdiffusion >>
rect 197 336 198 337 
<< pdiffusion >>
rect 210 336 211 337 
<< pdiffusion >>
rect 211 336 212 337 
<< pdiffusion >>
rect 212 336 213 337 
<< pdiffusion >>
rect 213 336 214 337 
<< pdiffusion >>
rect 214 336 215 337 
<< pdiffusion >>
rect 215 336 216 337 
<< m1 >>
rect 219 336 220 337 
<< m1 >>
rect 221 336 222 337 
<< m1 >>
rect 223 336 224 337 
<< pdiffusion >>
rect 228 336 229 337 
<< pdiffusion >>
rect 229 336 230 337 
<< pdiffusion >>
rect 230 336 231 337 
<< pdiffusion >>
rect 231 336 232 337 
<< pdiffusion >>
rect 232 336 233 337 
<< pdiffusion >>
rect 233 336 234 337 
<< m1 >>
rect 239 336 240 337 
<< pdiffusion >>
rect 246 336 247 337 
<< pdiffusion >>
rect 247 336 248 337 
<< pdiffusion >>
rect 248 336 249 337 
<< pdiffusion >>
rect 249 336 250 337 
<< pdiffusion >>
rect 250 336 251 337 
<< pdiffusion >>
rect 251 336 252 337 
<< pdiffusion >>
rect 264 336 265 337 
<< pdiffusion >>
rect 265 336 266 337 
<< pdiffusion >>
rect 266 336 267 337 
<< pdiffusion >>
rect 267 336 268 337 
<< pdiffusion >>
rect 268 336 269 337 
<< pdiffusion >>
rect 269 336 270 337 
<< m1 >>
rect 271 336 272 337 
<< pdiffusion >>
rect 282 336 283 337 
<< pdiffusion >>
rect 283 336 284 337 
<< pdiffusion >>
rect 284 336 285 337 
<< pdiffusion >>
rect 285 336 286 337 
<< pdiffusion >>
rect 286 336 287 337 
<< pdiffusion >>
rect 287 336 288 337 
<< pdiffusion >>
rect 300 336 301 337 
<< pdiffusion >>
rect 301 336 302 337 
<< pdiffusion >>
rect 302 336 303 337 
<< pdiffusion >>
rect 303 336 304 337 
<< pdiffusion >>
rect 304 336 305 337 
<< pdiffusion >>
rect 305 336 306 337 
<< m1 >>
rect 307 336 308 337 
<< pdiffusion >>
rect 318 336 319 337 
<< m1 >>
rect 319 336 320 337 
<< pdiffusion >>
rect 319 336 320 337 
<< pdiffusion >>
rect 320 336 321 337 
<< pdiffusion >>
rect 321 336 322 337 
<< pdiffusion >>
rect 322 336 323 337 
<< pdiffusion >>
rect 323 336 324 337 
<< m1 >>
rect 325 336 326 337 
<< m2 >>
rect 326 336 327 337 
<< m1 >>
rect 331 336 332 337 
<< m2 >>
rect 332 336 333 337 
<< m1 >>
rect 334 336 335 337 
<< pdiffusion >>
rect 336 336 337 337 
<< pdiffusion >>
rect 337 336 338 337 
<< pdiffusion >>
rect 338 336 339 337 
<< pdiffusion >>
rect 339 336 340 337 
<< m1 >>
rect 340 336 341 337 
<< pdiffusion >>
rect 340 336 341 337 
<< pdiffusion >>
rect 341 336 342 337 
<< m1 >>
rect 343 336 344 337 
<< m1 >>
rect 10 337 11 338 
<< pdiffusion >>
rect 12 337 13 338 
<< pdiffusion >>
rect 13 337 14 338 
<< pdiffusion >>
rect 14 337 15 338 
<< pdiffusion >>
rect 15 337 16 338 
<< pdiffusion >>
rect 16 337 17 338 
<< pdiffusion >>
rect 17 337 18 338 
<< m1 >>
rect 26 337 27 338 
<< m1 >>
rect 28 337 29 338 
<< pdiffusion >>
rect 30 337 31 338 
<< pdiffusion >>
rect 31 337 32 338 
<< pdiffusion >>
rect 32 337 33 338 
<< pdiffusion >>
rect 33 337 34 338 
<< pdiffusion >>
rect 34 337 35 338 
<< pdiffusion >>
rect 35 337 36 338 
<< m1 >>
rect 46 337 47 338 
<< m2 >>
rect 46 337 47 338 
<< pdiffusion >>
rect 48 337 49 338 
<< pdiffusion >>
rect 49 337 50 338 
<< pdiffusion >>
rect 50 337 51 338 
<< pdiffusion >>
rect 51 337 52 338 
<< pdiffusion >>
rect 52 337 53 338 
<< pdiffusion >>
rect 53 337 54 338 
<< m1 >>
rect 56 337 57 338 
<< m1 >>
rect 58 337 59 338 
<< m1 >>
rect 60 337 61 338 
<< m1 >>
rect 62 337 63 338 
<< pdiffusion >>
rect 66 337 67 338 
<< pdiffusion >>
rect 67 337 68 338 
<< pdiffusion >>
rect 68 337 69 338 
<< pdiffusion >>
rect 69 337 70 338 
<< pdiffusion >>
rect 70 337 71 338 
<< pdiffusion >>
rect 71 337 72 338 
<< pdiffusion >>
rect 84 337 85 338 
<< pdiffusion >>
rect 85 337 86 338 
<< pdiffusion >>
rect 86 337 87 338 
<< pdiffusion >>
rect 87 337 88 338 
<< pdiffusion >>
rect 88 337 89 338 
<< pdiffusion >>
rect 89 337 90 338 
<< pdiffusion >>
rect 102 337 103 338 
<< pdiffusion >>
rect 103 337 104 338 
<< pdiffusion >>
rect 104 337 105 338 
<< pdiffusion >>
rect 105 337 106 338 
<< pdiffusion >>
rect 106 337 107 338 
<< pdiffusion >>
rect 107 337 108 338 
<< m1 >>
rect 118 337 119 338 
<< pdiffusion >>
rect 120 337 121 338 
<< pdiffusion >>
rect 121 337 122 338 
<< pdiffusion >>
rect 122 337 123 338 
<< pdiffusion >>
rect 123 337 124 338 
<< pdiffusion >>
rect 124 337 125 338 
<< pdiffusion >>
rect 125 337 126 338 
<< pdiffusion >>
rect 138 337 139 338 
<< pdiffusion >>
rect 139 337 140 338 
<< pdiffusion >>
rect 140 337 141 338 
<< pdiffusion >>
rect 141 337 142 338 
<< pdiffusion >>
rect 142 337 143 338 
<< pdiffusion >>
rect 143 337 144 338 
<< m1 >>
rect 145 337 146 338 
<< pdiffusion >>
rect 156 337 157 338 
<< pdiffusion >>
rect 157 337 158 338 
<< pdiffusion >>
rect 158 337 159 338 
<< pdiffusion >>
rect 159 337 160 338 
<< pdiffusion >>
rect 160 337 161 338 
<< pdiffusion >>
rect 161 337 162 338 
<< pdiffusion >>
rect 174 337 175 338 
<< pdiffusion >>
rect 175 337 176 338 
<< pdiffusion >>
rect 176 337 177 338 
<< pdiffusion >>
rect 177 337 178 338 
<< pdiffusion >>
rect 178 337 179 338 
<< pdiffusion >>
rect 179 337 180 338 
<< pdiffusion >>
rect 192 337 193 338 
<< pdiffusion >>
rect 193 337 194 338 
<< pdiffusion >>
rect 194 337 195 338 
<< pdiffusion >>
rect 195 337 196 338 
<< pdiffusion >>
rect 196 337 197 338 
<< pdiffusion >>
rect 197 337 198 338 
<< pdiffusion >>
rect 210 337 211 338 
<< pdiffusion >>
rect 211 337 212 338 
<< pdiffusion >>
rect 212 337 213 338 
<< pdiffusion >>
rect 213 337 214 338 
<< pdiffusion >>
rect 214 337 215 338 
<< pdiffusion >>
rect 215 337 216 338 
<< m1 >>
rect 219 337 220 338 
<< m1 >>
rect 221 337 222 338 
<< m1 >>
rect 223 337 224 338 
<< pdiffusion >>
rect 228 337 229 338 
<< pdiffusion >>
rect 229 337 230 338 
<< pdiffusion >>
rect 230 337 231 338 
<< pdiffusion >>
rect 231 337 232 338 
<< pdiffusion >>
rect 232 337 233 338 
<< pdiffusion >>
rect 233 337 234 338 
<< m1 >>
rect 239 337 240 338 
<< pdiffusion >>
rect 246 337 247 338 
<< pdiffusion >>
rect 247 337 248 338 
<< pdiffusion >>
rect 248 337 249 338 
<< pdiffusion >>
rect 249 337 250 338 
<< pdiffusion >>
rect 250 337 251 338 
<< pdiffusion >>
rect 251 337 252 338 
<< pdiffusion >>
rect 264 337 265 338 
<< pdiffusion >>
rect 265 337 266 338 
<< pdiffusion >>
rect 266 337 267 338 
<< pdiffusion >>
rect 267 337 268 338 
<< pdiffusion >>
rect 268 337 269 338 
<< pdiffusion >>
rect 269 337 270 338 
<< m1 >>
rect 271 337 272 338 
<< pdiffusion >>
rect 282 337 283 338 
<< pdiffusion >>
rect 283 337 284 338 
<< pdiffusion >>
rect 284 337 285 338 
<< pdiffusion >>
rect 285 337 286 338 
<< pdiffusion >>
rect 286 337 287 338 
<< pdiffusion >>
rect 287 337 288 338 
<< pdiffusion >>
rect 300 337 301 338 
<< pdiffusion >>
rect 301 337 302 338 
<< pdiffusion >>
rect 302 337 303 338 
<< pdiffusion >>
rect 303 337 304 338 
<< pdiffusion >>
rect 304 337 305 338 
<< pdiffusion >>
rect 305 337 306 338 
<< m1 >>
rect 307 337 308 338 
<< pdiffusion >>
rect 318 337 319 338 
<< pdiffusion >>
rect 319 337 320 338 
<< pdiffusion >>
rect 320 337 321 338 
<< pdiffusion >>
rect 321 337 322 338 
<< pdiffusion >>
rect 322 337 323 338 
<< pdiffusion >>
rect 323 337 324 338 
<< m1 >>
rect 325 337 326 338 
<< m2 >>
rect 326 337 327 338 
<< m1 >>
rect 331 337 332 338 
<< m2 >>
rect 332 337 333 338 
<< m1 >>
rect 334 337 335 338 
<< pdiffusion >>
rect 336 337 337 338 
<< pdiffusion >>
rect 337 337 338 338 
<< pdiffusion >>
rect 338 337 339 338 
<< pdiffusion >>
rect 339 337 340 338 
<< pdiffusion >>
rect 340 337 341 338 
<< pdiffusion >>
rect 341 337 342 338 
<< m1 >>
rect 343 337 344 338 
<< m1 >>
rect 10 338 11 339 
<< pdiffusion >>
rect 12 338 13 339 
<< pdiffusion >>
rect 13 338 14 339 
<< pdiffusion >>
rect 14 338 15 339 
<< pdiffusion >>
rect 15 338 16 339 
<< pdiffusion >>
rect 16 338 17 339 
<< pdiffusion >>
rect 17 338 18 339 
<< m1 >>
rect 26 338 27 339 
<< m1 >>
rect 28 338 29 339 
<< pdiffusion >>
rect 30 338 31 339 
<< pdiffusion >>
rect 31 338 32 339 
<< pdiffusion >>
rect 32 338 33 339 
<< pdiffusion >>
rect 33 338 34 339 
<< pdiffusion >>
rect 34 338 35 339 
<< pdiffusion >>
rect 35 338 36 339 
<< m1 >>
rect 46 338 47 339 
<< m2 >>
rect 46 338 47 339 
<< pdiffusion >>
rect 48 338 49 339 
<< pdiffusion >>
rect 49 338 50 339 
<< pdiffusion >>
rect 50 338 51 339 
<< pdiffusion >>
rect 51 338 52 339 
<< pdiffusion >>
rect 52 338 53 339 
<< pdiffusion >>
rect 53 338 54 339 
<< m1 >>
rect 56 338 57 339 
<< m1 >>
rect 58 338 59 339 
<< m1 >>
rect 60 338 61 339 
<< m1 >>
rect 62 338 63 339 
<< pdiffusion >>
rect 66 338 67 339 
<< pdiffusion >>
rect 67 338 68 339 
<< pdiffusion >>
rect 68 338 69 339 
<< pdiffusion >>
rect 69 338 70 339 
<< pdiffusion >>
rect 70 338 71 339 
<< pdiffusion >>
rect 71 338 72 339 
<< pdiffusion >>
rect 84 338 85 339 
<< pdiffusion >>
rect 85 338 86 339 
<< pdiffusion >>
rect 86 338 87 339 
<< pdiffusion >>
rect 87 338 88 339 
<< pdiffusion >>
rect 88 338 89 339 
<< pdiffusion >>
rect 89 338 90 339 
<< pdiffusion >>
rect 102 338 103 339 
<< pdiffusion >>
rect 103 338 104 339 
<< pdiffusion >>
rect 104 338 105 339 
<< pdiffusion >>
rect 105 338 106 339 
<< pdiffusion >>
rect 106 338 107 339 
<< pdiffusion >>
rect 107 338 108 339 
<< m1 >>
rect 118 338 119 339 
<< pdiffusion >>
rect 120 338 121 339 
<< pdiffusion >>
rect 121 338 122 339 
<< pdiffusion >>
rect 122 338 123 339 
<< pdiffusion >>
rect 123 338 124 339 
<< pdiffusion >>
rect 124 338 125 339 
<< pdiffusion >>
rect 125 338 126 339 
<< pdiffusion >>
rect 138 338 139 339 
<< pdiffusion >>
rect 139 338 140 339 
<< pdiffusion >>
rect 140 338 141 339 
<< pdiffusion >>
rect 141 338 142 339 
<< pdiffusion >>
rect 142 338 143 339 
<< pdiffusion >>
rect 143 338 144 339 
<< m1 >>
rect 145 338 146 339 
<< pdiffusion >>
rect 156 338 157 339 
<< pdiffusion >>
rect 157 338 158 339 
<< pdiffusion >>
rect 158 338 159 339 
<< pdiffusion >>
rect 159 338 160 339 
<< pdiffusion >>
rect 160 338 161 339 
<< pdiffusion >>
rect 161 338 162 339 
<< pdiffusion >>
rect 174 338 175 339 
<< pdiffusion >>
rect 175 338 176 339 
<< pdiffusion >>
rect 176 338 177 339 
<< pdiffusion >>
rect 177 338 178 339 
<< pdiffusion >>
rect 178 338 179 339 
<< pdiffusion >>
rect 179 338 180 339 
<< pdiffusion >>
rect 192 338 193 339 
<< pdiffusion >>
rect 193 338 194 339 
<< pdiffusion >>
rect 194 338 195 339 
<< pdiffusion >>
rect 195 338 196 339 
<< pdiffusion >>
rect 196 338 197 339 
<< pdiffusion >>
rect 197 338 198 339 
<< pdiffusion >>
rect 210 338 211 339 
<< pdiffusion >>
rect 211 338 212 339 
<< pdiffusion >>
rect 212 338 213 339 
<< pdiffusion >>
rect 213 338 214 339 
<< pdiffusion >>
rect 214 338 215 339 
<< pdiffusion >>
rect 215 338 216 339 
<< m1 >>
rect 219 338 220 339 
<< m1 >>
rect 221 338 222 339 
<< m1 >>
rect 223 338 224 339 
<< pdiffusion >>
rect 228 338 229 339 
<< pdiffusion >>
rect 229 338 230 339 
<< pdiffusion >>
rect 230 338 231 339 
<< pdiffusion >>
rect 231 338 232 339 
<< pdiffusion >>
rect 232 338 233 339 
<< pdiffusion >>
rect 233 338 234 339 
<< m1 >>
rect 239 338 240 339 
<< pdiffusion >>
rect 246 338 247 339 
<< pdiffusion >>
rect 247 338 248 339 
<< pdiffusion >>
rect 248 338 249 339 
<< pdiffusion >>
rect 249 338 250 339 
<< pdiffusion >>
rect 250 338 251 339 
<< pdiffusion >>
rect 251 338 252 339 
<< pdiffusion >>
rect 264 338 265 339 
<< pdiffusion >>
rect 265 338 266 339 
<< pdiffusion >>
rect 266 338 267 339 
<< pdiffusion >>
rect 267 338 268 339 
<< pdiffusion >>
rect 268 338 269 339 
<< pdiffusion >>
rect 269 338 270 339 
<< m1 >>
rect 271 338 272 339 
<< pdiffusion >>
rect 282 338 283 339 
<< pdiffusion >>
rect 283 338 284 339 
<< pdiffusion >>
rect 284 338 285 339 
<< pdiffusion >>
rect 285 338 286 339 
<< pdiffusion >>
rect 286 338 287 339 
<< pdiffusion >>
rect 287 338 288 339 
<< pdiffusion >>
rect 300 338 301 339 
<< pdiffusion >>
rect 301 338 302 339 
<< pdiffusion >>
rect 302 338 303 339 
<< pdiffusion >>
rect 303 338 304 339 
<< pdiffusion >>
rect 304 338 305 339 
<< pdiffusion >>
rect 305 338 306 339 
<< m1 >>
rect 307 338 308 339 
<< pdiffusion >>
rect 318 338 319 339 
<< pdiffusion >>
rect 319 338 320 339 
<< pdiffusion >>
rect 320 338 321 339 
<< pdiffusion >>
rect 321 338 322 339 
<< pdiffusion >>
rect 322 338 323 339 
<< pdiffusion >>
rect 323 338 324 339 
<< m1 >>
rect 325 338 326 339 
<< m2 >>
rect 326 338 327 339 
<< m1 >>
rect 331 338 332 339 
<< m2 >>
rect 332 338 333 339 
<< m1 >>
rect 334 338 335 339 
<< pdiffusion >>
rect 336 338 337 339 
<< pdiffusion >>
rect 337 338 338 339 
<< pdiffusion >>
rect 338 338 339 339 
<< pdiffusion >>
rect 339 338 340 339 
<< pdiffusion >>
rect 340 338 341 339 
<< pdiffusion >>
rect 341 338 342 339 
<< m1 >>
rect 343 338 344 339 
<< m1 >>
rect 10 339 11 340 
<< pdiffusion >>
rect 12 339 13 340 
<< pdiffusion >>
rect 13 339 14 340 
<< pdiffusion >>
rect 14 339 15 340 
<< pdiffusion >>
rect 15 339 16 340 
<< pdiffusion >>
rect 16 339 17 340 
<< pdiffusion >>
rect 17 339 18 340 
<< m1 >>
rect 26 339 27 340 
<< m1 >>
rect 28 339 29 340 
<< pdiffusion >>
rect 30 339 31 340 
<< pdiffusion >>
rect 31 339 32 340 
<< pdiffusion >>
rect 32 339 33 340 
<< pdiffusion >>
rect 33 339 34 340 
<< pdiffusion >>
rect 34 339 35 340 
<< pdiffusion >>
rect 35 339 36 340 
<< m1 >>
rect 46 339 47 340 
<< m2 >>
rect 46 339 47 340 
<< pdiffusion >>
rect 48 339 49 340 
<< pdiffusion >>
rect 49 339 50 340 
<< pdiffusion >>
rect 50 339 51 340 
<< pdiffusion >>
rect 51 339 52 340 
<< pdiffusion >>
rect 52 339 53 340 
<< pdiffusion >>
rect 53 339 54 340 
<< m1 >>
rect 56 339 57 340 
<< m1 >>
rect 58 339 59 340 
<< m1 >>
rect 60 339 61 340 
<< m1 >>
rect 62 339 63 340 
<< pdiffusion >>
rect 66 339 67 340 
<< pdiffusion >>
rect 67 339 68 340 
<< pdiffusion >>
rect 68 339 69 340 
<< pdiffusion >>
rect 69 339 70 340 
<< pdiffusion >>
rect 70 339 71 340 
<< pdiffusion >>
rect 71 339 72 340 
<< pdiffusion >>
rect 84 339 85 340 
<< pdiffusion >>
rect 85 339 86 340 
<< pdiffusion >>
rect 86 339 87 340 
<< pdiffusion >>
rect 87 339 88 340 
<< pdiffusion >>
rect 88 339 89 340 
<< pdiffusion >>
rect 89 339 90 340 
<< pdiffusion >>
rect 102 339 103 340 
<< pdiffusion >>
rect 103 339 104 340 
<< pdiffusion >>
rect 104 339 105 340 
<< pdiffusion >>
rect 105 339 106 340 
<< pdiffusion >>
rect 106 339 107 340 
<< pdiffusion >>
rect 107 339 108 340 
<< m1 >>
rect 118 339 119 340 
<< pdiffusion >>
rect 120 339 121 340 
<< pdiffusion >>
rect 121 339 122 340 
<< pdiffusion >>
rect 122 339 123 340 
<< pdiffusion >>
rect 123 339 124 340 
<< pdiffusion >>
rect 124 339 125 340 
<< pdiffusion >>
rect 125 339 126 340 
<< pdiffusion >>
rect 138 339 139 340 
<< pdiffusion >>
rect 139 339 140 340 
<< pdiffusion >>
rect 140 339 141 340 
<< pdiffusion >>
rect 141 339 142 340 
<< pdiffusion >>
rect 142 339 143 340 
<< pdiffusion >>
rect 143 339 144 340 
<< m1 >>
rect 145 339 146 340 
<< pdiffusion >>
rect 156 339 157 340 
<< pdiffusion >>
rect 157 339 158 340 
<< pdiffusion >>
rect 158 339 159 340 
<< pdiffusion >>
rect 159 339 160 340 
<< pdiffusion >>
rect 160 339 161 340 
<< pdiffusion >>
rect 161 339 162 340 
<< pdiffusion >>
rect 174 339 175 340 
<< pdiffusion >>
rect 175 339 176 340 
<< pdiffusion >>
rect 176 339 177 340 
<< pdiffusion >>
rect 177 339 178 340 
<< pdiffusion >>
rect 178 339 179 340 
<< pdiffusion >>
rect 179 339 180 340 
<< pdiffusion >>
rect 192 339 193 340 
<< pdiffusion >>
rect 193 339 194 340 
<< pdiffusion >>
rect 194 339 195 340 
<< pdiffusion >>
rect 195 339 196 340 
<< pdiffusion >>
rect 196 339 197 340 
<< pdiffusion >>
rect 197 339 198 340 
<< pdiffusion >>
rect 210 339 211 340 
<< pdiffusion >>
rect 211 339 212 340 
<< pdiffusion >>
rect 212 339 213 340 
<< pdiffusion >>
rect 213 339 214 340 
<< pdiffusion >>
rect 214 339 215 340 
<< pdiffusion >>
rect 215 339 216 340 
<< m1 >>
rect 219 339 220 340 
<< m1 >>
rect 221 339 222 340 
<< m1 >>
rect 223 339 224 340 
<< pdiffusion >>
rect 228 339 229 340 
<< pdiffusion >>
rect 229 339 230 340 
<< pdiffusion >>
rect 230 339 231 340 
<< pdiffusion >>
rect 231 339 232 340 
<< pdiffusion >>
rect 232 339 233 340 
<< pdiffusion >>
rect 233 339 234 340 
<< m1 >>
rect 239 339 240 340 
<< pdiffusion >>
rect 246 339 247 340 
<< pdiffusion >>
rect 247 339 248 340 
<< pdiffusion >>
rect 248 339 249 340 
<< pdiffusion >>
rect 249 339 250 340 
<< pdiffusion >>
rect 250 339 251 340 
<< pdiffusion >>
rect 251 339 252 340 
<< pdiffusion >>
rect 264 339 265 340 
<< pdiffusion >>
rect 265 339 266 340 
<< pdiffusion >>
rect 266 339 267 340 
<< pdiffusion >>
rect 267 339 268 340 
<< pdiffusion >>
rect 268 339 269 340 
<< pdiffusion >>
rect 269 339 270 340 
<< m1 >>
rect 271 339 272 340 
<< pdiffusion >>
rect 282 339 283 340 
<< pdiffusion >>
rect 283 339 284 340 
<< pdiffusion >>
rect 284 339 285 340 
<< pdiffusion >>
rect 285 339 286 340 
<< pdiffusion >>
rect 286 339 287 340 
<< pdiffusion >>
rect 287 339 288 340 
<< pdiffusion >>
rect 300 339 301 340 
<< pdiffusion >>
rect 301 339 302 340 
<< pdiffusion >>
rect 302 339 303 340 
<< pdiffusion >>
rect 303 339 304 340 
<< pdiffusion >>
rect 304 339 305 340 
<< pdiffusion >>
rect 305 339 306 340 
<< m1 >>
rect 307 339 308 340 
<< pdiffusion >>
rect 318 339 319 340 
<< pdiffusion >>
rect 319 339 320 340 
<< pdiffusion >>
rect 320 339 321 340 
<< pdiffusion >>
rect 321 339 322 340 
<< pdiffusion >>
rect 322 339 323 340 
<< pdiffusion >>
rect 323 339 324 340 
<< m1 >>
rect 325 339 326 340 
<< m2 >>
rect 326 339 327 340 
<< m1 >>
rect 331 339 332 340 
<< m2 >>
rect 332 339 333 340 
<< m1 >>
rect 334 339 335 340 
<< pdiffusion >>
rect 336 339 337 340 
<< pdiffusion >>
rect 337 339 338 340 
<< pdiffusion >>
rect 338 339 339 340 
<< pdiffusion >>
rect 339 339 340 340 
<< pdiffusion >>
rect 340 339 341 340 
<< pdiffusion >>
rect 341 339 342 340 
<< m1 >>
rect 343 339 344 340 
<< m1 >>
rect 10 340 11 341 
<< pdiffusion >>
rect 12 340 13 341 
<< pdiffusion >>
rect 13 340 14 341 
<< pdiffusion >>
rect 14 340 15 341 
<< pdiffusion >>
rect 15 340 16 341 
<< pdiffusion >>
rect 16 340 17 341 
<< pdiffusion >>
rect 17 340 18 341 
<< m1 >>
rect 26 340 27 341 
<< m1 >>
rect 28 340 29 341 
<< pdiffusion >>
rect 30 340 31 341 
<< pdiffusion >>
rect 31 340 32 341 
<< pdiffusion >>
rect 32 340 33 341 
<< pdiffusion >>
rect 33 340 34 341 
<< pdiffusion >>
rect 34 340 35 341 
<< pdiffusion >>
rect 35 340 36 341 
<< m1 >>
rect 46 340 47 341 
<< m2 >>
rect 46 340 47 341 
<< pdiffusion >>
rect 48 340 49 341 
<< pdiffusion >>
rect 49 340 50 341 
<< pdiffusion >>
rect 50 340 51 341 
<< pdiffusion >>
rect 51 340 52 341 
<< pdiffusion >>
rect 52 340 53 341 
<< pdiffusion >>
rect 53 340 54 341 
<< m1 >>
rect 56 340 57 341 
<< m1 >>
rect 58 340 59 341 
<< m1 >>
rect 60 340 61 341 
<< m1 >>
rect 62 340 63 341 
<< pdiffusion >>
rect 66 340 67 341 
<< pdiffusion >>
rect 67 340 68 341 
<< pdiffusion >>
rect 68 340 69 341 
<< pdiffusion >>
rect 69 340 70 341 
<< pdiffusion >>
rect 70 340 71 341 
<< pdiffusion >>
rect 71 340 72 341 
<< pdiffusion >>
rect 84 340 85 341 
<< pdiffusion >>
rect 85 340 86 341 
<< pdiffusion >>
rect 86 340 87 341 
<< pdiffusion >>
rect 87 340 88 341 
<< pdiffusion >>
rect 88 340 89 341 
<< pdiffusion >>
rect 89 340 90 341 
<< pdiffusion >>
rect 102 340 103 341 
<< pdiffusion >>
rect 103 340 104 341 
<< pdiffusion >>
rect 104 340 105 341 
<< pdiffusion >>
rect 105 340 106 341 
<< pdiffusion >>
rect 106 340 107 341 
<< pdiffusion >>
rect 107 340 108 341 
<< m1 >>
rect 118 340 119 341 
<< pdiffusion >>
rect 120 340 121 341 
<< pdiffusion >>
rect 121 340 122 341 
<< pdiffusion >>
rect 122 340 123 341 
<< pdiffusion >>
rect 123 340 124 341 
<< pdiffusion >>
rect 124 340 125 341 
<< pdiffusion >>
rect 125 340 126 341 
<< pdiffusion >>
rect 138 340 139 341 
<< pdiffusion >>
rect 139 340 140 341 
<< pdiffusion >>
rect 140 340 141 341 
<< pdiffusion >>
rect 141 340 142 341 
<< pdiffusion >>
rect 142 340 143 341 
<< pdiffusion >>
rect 143 340 144 341 
<< m1 >>
rect 145 340 146 341 
<< pdiffusion >>
rect 156 340 157 341 
<< pdiffusion >>
rect 157 340 158 341 
<< pdiffusion >>
rect 158 340 159 341 
<< pdiffusion >>
rect 159 340 160 341 
<< pdiffusion >>
rect 160 340 161 341 
<< pdiffusion >>
rect 161 340 162 341 
<< pdiffusion >>
rect 174 340 175 341 
<< pdiffusion >>
rect 175 340 176 341 
<< pdiffusion >>
rect 176 340 177 341 
<< pdiffusion >>
rect 177 340 178 341 
<< pdiffusion >>
rect 178 340 179 341 
<< pdiffusion >>
rect 179 340 180 341 
<< pdiffusion >>
rect 192 340 193 341 
<< pdiffusion >>
rect 193 340 194 341 
<< pdiffusion >>
rect 194 340 195 341 
<< pdiffusion >>
rect 195 340 196 341 
<< pdiffusion >>
rect 196 340 197 341 
<< pdiffusion >>
rect 197 340 198 341 
<< pdiffusion >>
rect 210 340 211 341 
<< pdiffusion >>
rect 211 340 212 341 
<< pdiffusion >>
rect 212 340 213 341 
<< pdiffusion >>
rect 213 340 214 341 
<< pdiffusion >>
rect 214 340 215 341 
<< pdiffusion >>
rect 215 340 216 341 
<< m1 >>
rect 219 340 220 341 
<< m1 >>
rect 221 340 222 341 
<< m1 >>
rect 223 340 224 341 
<< pdiffusion >>
rect 228 340 229 341 
<< pdiffusion >>
rect 229 340 230 341 
<< pdiffusion >>
rect 230 340 231 341 
<< pdiffusion >>
rect 231 340 232 341 
<< pdiffusion >>
rect 232 340 233 341 
<< pdiffusion >>
rect 233 340 234 341 
<< m1 >>
rect 239 340 240 341 
<< pdiffusion >>
rect 246 340 247 341 
<< pdiffusion >>
rect 247 340 248 341 
<< pdiffusion >>
rect 248 340 249 341 
<< pdiffusion >>
rect 249 340 250 341 
<< pdiffusion >>
rect 250 340 251 341 
<< pdiffusion >>
rect 251 340 252 341 
<< pdiffusion >>
rect 264 340 265 341 
<< pdiffusion >>
rect 265 340 266 341 
<< pdiffusion >>
rect 266 340 267 341 
<< pdiffusion >>
rect 267 340 268 341 
<< pdiffusion >>
rect 268 340 269 341 
<< pdiffusion >>
rect 269 340 270 341 
<< m1 >>
rect 271 340 272 341 
<< pdiffusion >>
rect 282 340 283 341 
<< pdiffusion >>
rect 283 340 284 341 
<< pdiffusion >>
rect 284 340 285 341 
<< pdiffusion >>
rect 285 340 286 341 
<< pdiffusion >>
rect 286 340 287 341 
<< pdiffusion >>
rect 287 340 288 341 
<< pdiffusion >>
rect 300 340 301 341 
<< pdiffusion >>
rect 301 340 302 341 
<< pdiffusion >>
rect 302 340 303 341 
<< pdiffusion >>
rect 303 340 304 341 
<< pdiffusion >>
rect 304 340 305 341 
<< pdiffusion >>
rect 305 340 306 341 
<< m1 >>
rect 307 340 308 341 
<< pdiffusion >>
rect 318 340 319 341 
<< pdiffusion >>
rect 319 340 320 341 
<< pdiffusion >>
rect 320 340 321 341 
<< pdiffusion >>
rect 321 340 322 341 
<< pdiffusion >>
rect 322 340 323 341 
<< pdiffusion >>
rect 323 340 324 341 
<< m1 >>
rect 325 340 326 341 
<< m2 >>
rect 326 340 327 341 
<< m1 >>
rect 331 340 332 341 
<< m2 >>
rect 332 340 333 341 
<< m1 >>
rect 334 340 335 341 
<< pdiffusion >>
rect 336 340 337 341 
<< pdiffusion >>
rect 337 340 338 341 
<< pdiffusion >>
rect 338 340 339 341 
<< pdiffusion >>
rect 339 340 340 341 
<< pdiffusion >>
rect 340 340 341 341 
<< pdiffusion >>
rect 341 340 342 341 
<< m1 >>
rect 343 340 344 341 
<< m1 >>
rect 10 341 11 342 
<< pdiffusion >>
rect 12 341 13 342 
<< pdiffusion >>
rect 13 341 14 342 
<< pdiffusion >>
rect 14 341 15 342 
<< pdiffusion >>
rect 15 341 16 342 
<< m1 >>
rect 16 341 17 342 
<< pdiffusion >>
rect 16 341 17 342 
<< pdiffusion >>
rect 17 341 18 342 
<< m1 >>
rect 26 341 27 342 
<< m1 >>
rect 28 341 29 342 
<< pdiffusion >>
rect 30 341 31 342 
<< pdiffusion >>
rect 31 341 32 342 
<< pdiffusion >>
rect 32 341 33 342 
<< pdiffusion >>
rect 33 341 34 342 
<< pdiffusion >>
rect 34 341 35 342 
<< pdiffusion >>
rect 35 341 36 342 
<< m1 >>
rect 46 341 47 342 
<< m2 >>
rect 46 341 47 342 
<< pdiffusion >>
rect 48 341 49 342 
<< pdiffusion >>
rect 49 341 50 342 
<< pdiffusion >>
rect 50 341 51 342 
<< pdiffusion >>
rect 51 341 52 342 
<< pdiffusion >>
rect 52 341 53 342 
<< pdiffusion >>
rect 53 341 54 342 
<< m1 >>
rect 56 341 57 342 
<< m1 >>
rect 58 341 59 342 
<< m1 >>
rect 60 341 61 342 
<< m1 >>
rect 62 341 63 342 
<< pdiffusion >>
rect 66 341 67 342 
<< pdiffusion >>
rect 67 341 68 342 
<< pdiffusion >>
rect 68 341 69 342 
<< pdiffusion >>
rect 69 341 70 342 
<< pdiffusion >>
rect 70 341 71 342 
<< pdiffusion >>
rect 71 341 72 342 
<< pdiffusion >>
rect 84 341 85 342 
<< pdiffusion >>
rect 85 341 86 342 
<< pdiffusion >>
rect 86 341 87 342 
<< pdiffusion >>
rect 87 341 88 342 
<< pdiffusion >>
rect 88 341 89 342 
<< pdiffusion >>
rect 89 341 90 342 
<< pdiffusion >>
rect 102 341 103 342 
<< pdiffusion >>
rect 103 341 104 342 
<< pdiffusion >>
rect 104 341 105 342 
<< pdiffusion >>
rect 105 341 106 342 
<< pdiffusion >>
rect 106 341 107 342 
<< pdiffusion >>
rect 107 341 108 342 
<< m1 >>
rect 118 341 119 342 
<< pdiffusion >>
rect 120 341 121 342 
<< pdiffusion >>
rect 121 341 122 342 
<< pdiffusion >>
rect 122 341 123 342 
<< pdiffusion >>
rect 123 341 124 342 
<< m1 >>
rect 124 341 125 342 
<< pdiffusion >>
rect 124 341 125 342 
<< pdiffusion >>
rect 125 341 126 342 
<< pdiffusion >>
rect 138 341 139 342 
<< pdiffusion >>
rect 139 341 140 342 
<< pdiffusion >>
rect 140 341 141 342 
<< pdiffusion >>
rect 141 341 142 342 
<< pdiffusion >>
rect 142 341 143 342 
<< pdiffusion >>
rect 143 341 144 342 
<< m1 >>
rect 145 341 146 342 
<< pdiffusion >>
rect 156 341 157 342 
<< pdiffusion >>
rect 157 341 158 342 
<< pdiffusion >>
rect 158 341 159 342 
<< pdiffusion >>
rect 159 341 160 342 
<< pdiffusion >>
rect 160 341 161 342 
<< pdiffusion >>
rect 161 341 162 342 
<< pdiffusion >>
rect 174 341 175 342 
<< pdiffusion >>
rect 175 341 176 342 
<< pdiffusion >>
rect 176 341 177 342 
<< pdiffusion >>
rect 177 341 178 342 
<< pdiffusion >>
rect 178 341 179 342 
<< pdiffusion >>
rect 179 341 180 342 
<< pdiffusion >>
rect 192 341 193 342 
<< pdiffusion >>
rect 193 341 194 342 
<< pdiffusion >>
rect 194 341 195 342 
<< pdiffusion >>
rect 195 341 196 342 
<< pdiffusion >>
rect 196 341 197 342 
<< pdiffusion >>
rect 197 341 198 342 
<< pdiffusion >>
rect 210 341 211 342 
<< pdiffusion >>
rect 211 341 212 342 
<< pdiffusion >>
rect 212 341 213 342 
<< pdiffusion >>
rect 213 341 214 342 
<< pdiffusion >>
rect 214 341 215 342 
<< pdiffusion >>
rect 215 341 216 342 
<< m1 >>
rect 219 341 220 342 
<< m1 >>
rect 221 341 222 342 
<< m1 >>
rect 223 341 224 342 
<< pdiffusion >>
rect 228 341 229 342 
<< pdiffusion >>
rect 229 341 230 342 
<< pdiffusion >>
rect 230 341 231 342 
<< pdiffusion >>
rect 231 341 232 342 
<< pdiffusion >>
rect 232 341 233 342 
<< pdiffusion >>
rect 233 341 234 342 
<< m1 >>
rect 239 341 240 342 
<< pdiffusion >>
rect 246 341 247 342 
<< pdiffusion >>
rect 247 341 248 342 
<< pdiffusion >>
rect 248 341 249 342 
<< pdiffusion >>
rect 249 341 250 342 
<< pdiffusion >>
rect 250 341 251 342 
<< pdiffusion >>
rect 251 341 252 342 
<< pdiffusion >>
rect 264 341 265 342 
<< pdiffusion >>
rect 265 341 266 342 
<< pdiffusion >>
rect 266 341 267 342 
<< pdiffusion >>
rect 267 341 268 342 
<< m1 >>
rect 268 341 269 342 
<< pdiffusion >>
rect 268 341 269 342 
<< pdiffusion >>
rect 269 341 270 342 
<< m1 >>
rect 271 341 272 342 
<< pdiffusion >>
rect 282 341 283 342 
<< pdiffusion >>
rect 283 341 284 342 
<< pdiffusion >>
rect 284 341 285 342 
<< pdiffusion >>
rect 285 341 286 342 
<< pdiffusion >>
rect 286 341 287 342 
<< pdiffusion >>
rect 287 341 288 342 
<< pdiffusion >>
rect 300 341 301 342 
<< pdiffusion >>
rect 301 341 302 342 
<< pdiffusion >>
rect 302 341 303 342 
<< pdiffusion >>
rect 303 341 304 342 
<< m1 >>
rect 304 341 305 342 
<< pdiffusion >>
rect 304 341 305 342 
<< pdiffusion >>
rect 305 341 306 342 
<< m1 >>
rect 307 341 308 342 
<< pdiffusion >>
rect 318 341 319 342 
<< pdiffusion >>
rect 319 341 320 342 
<< pdiffusion >>
rect 320 341 321 342 
<< pdiffusion >>
rect 321 341 322 342 
<< pdiffusion >>
rect 322 341 323 342 
<< pdiffusion >>
rect 323 341 324 342 
<< m1 >>
rect 325 341 326 342 
<< m2 >>
rect 326 341 327 342 
<< m1 >>
rect 331 341 332 342 
<< m2 >>
rect 332 341 333 342 
<< m1 >>
rect 334 341 335 342 
<< pdiffusion >>
rect 336 341 337 342 
<< pdiffusion >>
rect 337 341 338 342 
<< pdiffusion >>
rect 338 341 339 342 
<< pdiffusion >>
rect 339 341 340 342 
<< m1 >>
rect 340 341 341 342 
<< pdiffusion >>
rect 340 341 341 342 
<< pdiffusion >>
rect 341 341 342 342 
<< m1 >>
rect 343 341 344 342 
<< m1 >>
rect 10 342 11 343 
<< m1 >>
rect 16 342 17 343 
<< m1 >>
rect 26 342 27 343 
<< m1 >>
rect 28 342 29 343 
<< m1 >>
rect 46 342 47 343 
<< m2 >>
rect 46 342 47 343 
<< m1 >>
rect 56 342 57 343 
<< m1 >>
rect 58 342 59 343 
<< m1 >>
rect 60 342 61 343 
<< m2 >>
rect 60 342 61 343 
<< m2c >>
rect 60 342 61 343 
<< m1 >>
rect 60 342 61 343 
<< m2 >>
rect 60 342 61 343 
<< m2 >>
rect 61 342 62 343 
<< m1 >>
rect 62 342 63 343 
<< m2 >>
rect 62 342 63 343 
<< m2 >>
rect 63 342 64 343 
<< m1 >>
rect 64 342 65 343 
<< m2 >>
rect 64 342 65 343 
<< m2c >>
rect 64 342 65 343 
<< m1 >>
rect 64 342 65 343 
<< m2 >>
rect 64 342 65 343 
<< m1 >>
rect 118 342 119 343 
<< m1 >>
rect 124 342 125 343 
<< m1 >>
rect 145 342 146 343 
<< m1 >>
rect 219 342 220 343 
<< m1 >>
rect 221 342 222 343 
<< m1 >>
rect 223 342 224 343 
<< m1 >>
rect 239 342 240 343 
<< m1 >>
rect 268 342 269 343 
<< m1 >>
rect 271 342 272 343 
<< m1 >>
rect 304 342 305 343 
<< m1 >>
rect 307 342 308 343 
<< m1 >>
rect 325 342 326 343 
<< m2 >>
rect 326 342 327 343 
<< m1 >>
rect 331 342 332 343 
<< m2 >>
rect 332 342 333 343 
<< m1 >>
rect 334 342 335 343 
<< m1 >>
rect 340 342 341 343 
<< m1 >>
rect 343 342 344 343 
<< m1 >>
rect 10 343 11 344 
<< m1 >>
rect 16 343 17 344 
<< m1 >>
rect 26 343 27 344 
<< m1 >>
rect 28 343 29 344 
<< m1 >>
rect 46 343 47 344 
<< m2 >>
rect 46 343 47 344 
<< m1 >>
rect 56 343 57 344 
<< m1 >>
rect 58 343 59 344 
<< m1 >>
rect 62 343 63 344 
<< m1 >>
rect 64 343 65 344 
<< m1 >>
rect 118 343 119 344 
<< m1 >>
rect 124 343 125 344 
<< m1 >>
rect 145 343 146 344 
<< m1 >>
rect 219 343 220 344 
<< m1 >>
rect 221 343 222 344 
<< m1 >>
rect 223 343 224 344 
<< m1 >>
rect 239 343 240 344 
<< m1 >>
rect 268 343 269 344 
<< m1 >>
rect 269 343 270 344 
<< m1 >>
rect 270 343 271 344 
<< m1 >>
rect 271 343 272 344 
<< m1 >>
rect 304 343 305 344 
<< m1 >>
rect 307 343 308 344 
<< m1 >>
rect 325 343 326 344 
<< m2 >>
rect 326 343 327 344 
<< m1 >>
rect 331 343 332 344 
<< m2 >>
rect 332 343 333 344 
<< m1 >>
rect 334 343 335 344 
<< m1 >>
rect 340 343 341 344 
<< m1 >>
rect 343 343 344 344 
<< m1 >>
rect 10 344 11 345 
<< m1 >>
rect 16 344 17 345 
<< m1 >>
rect 26 344 27 345 
<< m2 >>
rect 26 344 27 345 
<< m2c >>
rect 26 344 27 345 
<< m1 >>
rect 26 344 27 345 
<< m2 >>
rect 26 344 27 345 
<< m1 >>
rect 28 344 29 345 
<< m2 >>
rect 28 344 29 345 
<< m2c >>
rect 28 344 29 345 
<< m1 >>
rect 28 344 29 345 
<< m2 >>
rect 28 344 29 345 
<< m1 >>
rect 46 344 47 345 
<< m2 >>
rect 46 344 47 345 
<< m1 >>
rect 47 344 48 345 
<< m1 >>
rect 48 344 49 345 
<< m2 >>
rect 48 344 49 345 
<< m2c >>
rect 48 344 49 345 
<< m1 >>
rect 48 344 49 345 
<< m2 >>
rect 48 344 49 345 
<< m1 >>
rect 56 344 57 345 
<< m2 >>
rect 56 344 57 345 
<< m2c >>
rect 56 344 57 345 
<< m1 >>
rect 56 344 57 345 
<< m2 >>
rect 56 344 57 345 
<< m1 >>
rect 58 344 59 345 
<< m2 >>
rect 58 344 59 345 
<< m2c >>
rect 58 344 59 345 
<< m1 >>
rect 58 344 59 345 
<< m2 >>
rect 58 344 59 345 
<< m1 >>
rect 62 344 63 345 
<< m2 >>
rect 62 344 63 345 
<< m2c >>
rect 62 344 63 345 
<< m1 >>
rect 62 344 63 345 
<< m2 >>
rect 62 344 63 345 
<< m1 >>
rect 64 344 65 345 
<< m1 >>
rect 65 344 66 345 
<< m1 >>
rect 66 344 67 345 
<< m2 >>
rect 66 344 67 345 
<< m2c >>
rect 66 344 67 345 
<< m1 >>
rect 66 344 67 345 
<< m2 >>
rect 66 344 67 345 
<< m1 >>
rect 118 344 119 345 
<< m1 >>
rect 119 344 120 345 
<< m1 >>
rect 120 344 121 345 
<< m2 >>
rect 120 344 121 345 
<< m2c >>
rect 120 344 121 345 
<< m1 >>
rect 120 344 121 345 
<< m2 >>
rect 120 344 121 345 
<< m1 >>
rect 124 344 125 345 
<< m2 >>
rect 124 344 125 345 
<< m2c >>
rect 124 344 125 345 
<< m1 >>
rect 124 344 125 345 
<< m2 >>
rect 124 344 125 345 
<< m1 >>
rect 145 344 146 345 
<< m2 >>
rect 145 344 146 345 
<< m2c >>
rect 145 344 146 345 
<< m1 >>
rect 145 344 146 345 
<< m2 >>
rect 145 344 146 345 
<< m1 >>
rect 219 344 220 345 
<< m1 >>
rect 221 344 222 345 
<< m1 >>
rect 223 344 224 345 
<< m1 >>
rect 239 344 240 345 
<< m1 >>
rect 304 344 305 345 
<< m1 >>
rect 307 344 308 345 
<< m1 >>
rect 325 344 326 345 
<< m2 >>
rect 326 344 327 345 
<< m1 >>
rect 331 344 332 345 
<< m2 >>
rect 332 344 333 345 
<< m1 >>
rect 334 344 335 345 
<< m1 >>
rect 340 344 341 345 
<< m1 >>
rect 343 344 344 345 
<< m1 >>
rect 10 345 11 346 
<< m1 >>
rect 16 345 17 346 
<< m2 >>
rect 26 345 27 346 
<< m2 >>
rect 28 345 29 346 
<< m2 >>
rect 46 345 47 346 
<< m2 >>
rect 48 345 49 346 
<< m2 >>
rect 56 345 57 346 
<< m2 >>
rect 58 345 59 346 
<< m2 >>
rect 62 345 63 346 
<< m2 >>
rect 66 345 67 346 
<< m2 >>
rect 120 345 121 346 
<< m2 >>
rect 124 345 125 346 
<< m2 >>
rect 145 345 146 346 
<< m1 >>
rect 219 345 220 346 
<< m1 >>
rect 221 345 222 346 
<< m1 >>
rect 223 345 224 346 
<< m1 >>
rect 239 345 240 346 
<< m1 >>
rect 304 345 305 346 
<< m1 >>
rect 307 345 308 346 
<< m1 >>
rect 325 345 326 346 
<< m2 >>
rect 326 345 327 346 
<< m1 >>
rect 331 345 332 346 
<< m2 >>
rect 332 345 333 346 
<< m1 >>
rect 334 345 335 346 
<< m1 >>
rect 340 345 341 346 
<< m1 >>
rect 343 345 344 346 
<< m1 >>
rect 10 346 11 347 
<< m1 >>
rect 16 346 17 347 
<< m1 >>
rect 17 346 18 347 
<< m1 >>
rect 18 346 19 347 
<< m1 >>
rect 19 346 20 347 
<< m1 >>
rect 20 346 21 347 
<< m1 >>
rect 21 346 22 347 
<< m1 >>
rect 22 346 23 347 
<< m1 >>
rect 23 346 24 347 
<< m1 >>
rect 24 346 25 347 
<< m1 >>
rect 25 346 26 347 
<< m1 >>
rect 26 346 27 347 
<< m2 >>
rect 26 346 27 347 
<< m1 >>
rect 27 346 28 347 
<< m1 >>
rect 28 346 29 347 
<< m2 >>
rect 28 346 29 347 
<< m1 >>
rect 29 346 30 347 
<< m1 >>
rect 30 346 31 347 
<< m1 >>
rect 31 346 32 347 
<< m1 >>
rect 32 346 33 347 
<< m1 >>
rect 33 346 34 347 
<< m1 >>
rect 34 346 35 347 
<< m1 >>
rect 35 346 36 347 
<< m1 >>
rect 36 346 37 347 
<< m1 >>
rect 37 346 38 347 
<< m1 >>
rect 38 346 39 347 
<< m1 >>
rect 39 346 40 347 
<< m1 >>
rect 40 346 41 347 
<< m1 >>
rect 41 346 42 347 
<< m1 >>
rect 42 346 43 347 
<< m1 >>
rect 43 346 44 347 
<< m1 >>
rect 44 346 45 347 
<< m1 >>
rect 45 346 46 347 
<< m1 >>
rect 46 346 47 347 
<< m2 >>
rect 46 346 47 347 
<< m1 >>
rect 47 346 48 347 
<< m1 >>
rect 48 346 49 347 
<< m2 >>
rect 48 346 49 347 
<< m1 >>
rect 49 346 50 347 
<< m1 >>
rect 50 346 51 347 
<< m1 >>
rect 51 346 52 347 
<< m1 >>
rect 52 346 53 347 
<< m1 >>
rect 53 346 54 347 
<< m1 >>
rect 54 346 55 347 
<< m1 >>
rect 55 346 56 347 
<< m1 >>
rect 56 346 57 347 
<< m2 >>
rect 56 346 57 347 
<< m1 >>
rect 57 346 58 347 
<< m1 >>
rect 58 346 59 347 
<< m2 >>
rect 58 346 59 347 
<< m1 >>
rect 59 346 60 347 
<< m1 >>
rect 60 346 61 347 
<< m1 >>
rect 61 346 62 347 
<< m1 >>
rect 62 346 63 347 
<< m2 >>
rect 62 346 63 347 
<< m1 >>
rect 63 346 64 347 
<< m1 >>
rect 64 346 65 347 
<< m1 >>
rect 65 346 66 347 
<< m1 >>
rect 66 346 67 347 
<< m2 >>
rect 66 346 67 347 
<< m1 >>
rect 67 346 68 347 
<< m1 >>
rect 68 346 69 347 
<< m1 >>
rect 69 346 70 347 
<< m1 >>
rect 70 346 71 347 
<< m1 >>
rect 71 346 72 347 
<< m1 >>
rect 72 346 73 347 
<< m1 >>
rect 73 346 74 347 
<< m1 >>
rect 74 346 75 347 
<< m1 >>
rect 75 346 76 347 
<< m1 >>
rect 76 346 77 347 
<< m1 >>
rect 77 346 78 347 
<< m1 >>
rect 78 346 79 347 
<< m1 >>
rect 79 346 80 347 
<< m1 >>
rect 80 346 81 347 
<< m1 >>
rect 81 346 82 347 
<< m1 >>
rect 82 346 83 347 
<< m1 >>
rect 83 346 84 347 
<< m1 >>
rect 84 346 85 347 
<< m1 >>
rect 85 346 86 347 
<< m1 >>
rect 86 346 87 347 
<< m1 >>
rect 87 346 88 347 
<< m1 >>
rect 88 346 89 347 
<< m1 >>
rect 89 346 90 347 
<< m1 >>
rect 90 346 91 347 
<< m1 >>
rect 91 346 92 347 
<< m1 >>
rect 92 346 93 347 
<< m1 >>
rect 93 346 94 347 
<< m1 >>
rect 94 346 95 347 
<< m1 >>
rect 95 346 96 347 
<< m1 >>
rect 96 346 97 347 
<< m1 >>
rect 97 346 98 347 
<< m1 >>
rect 98 346 99 347 
<< m1 >>
rect 99 346 100 347 
<< m1 >>
rect 100 346 101 347 
<< m1 >>
rect 101 346 102 347 
<< m1 >>
rect 102 346 103 347 
<< m1 >>
rect 103 346 104 347 
<< m1 >>
rect 104 346 105 347 
<< m1 >>
rect 105 346 106 347 
<< m1 >>
rect 106 346 107 347 
<< m1 >>
rect 107 346 108 347 
<< m1 >>
rect 108 346 109 347 
<< m1 >>
rect 109 346 110 347 
<< m1 >>
rect 110 346 111 347 
<< m1 >>
rect 111 346 112 347 
<< m1 >>
rect 112 346 113 347 
<< m1 >>
rect 113 346 114 347 
<< m1 >>
rect 114 346 115 347 
<< m1 >>
rect 115 346 116 347 
<< m1 >>
rect 116 346 117 347 
<< m1 >>
rect 117 346 118 347 
<< m1 >>
rect 118 346 119 347 
<< m1 >>
rect 119 346 120 347 
<< m1 >>
rect 120 346 121 347 
<< m2 >>
rect 120 346 121 347 
<< m1 >>
rect 121 346 122 347 
<< m2 >>
rect 121 346 122 347 
<< m1 >>
rect 122 346 123 347 
<< m2 >>
rect 122 346 123 347 
<< m1 >>
rect 123 346 124 347 
<< m2 >>
rect 123 346 124 347 
<< m1 >>
rect 124 346 125 347 
<< m2 >>
rect 124 346 125 347 
<< m1 >>
rect 125 346 126 347 
<< m1 >>
rect 126 346 127 347 
<< m1 >>
rect 127 346 128 347 
<< m1 >>
rect 128 346 129 347 
<< m1 >>
rect 129 346 130 347 
<< m1 >>
rect 130 346 131 347 
<< m1 >>
rect 131 346 132 347 
<< m1 >>
rect 132 346 133 347 
<< m1 >>
rect 133 346 134 347 
<< m1 >>
rect 134 346 135 347 
<< m1 >>
rect 135 346 136 347 
<< m1 >>
rect 136 346 137 347 
<< m1 >>
rect 137 346 138 347 
<< m1 >>
rect 138 346 139 347 
<< m1 >>
rect 139 346 140 347 
<< m1 >>
rect 140 346 141 347 
<< m1 >>
rect 141 346 142 347 
<< m1 >>
rect 142 346 143 347 
<< m1 >>
rect 143 346 144 347 
<< m1 >>
rect 144 346 145 347 
<< m1 >>
rect 145 346 146 347 
<< m2 >>
rect 145 346 146 347 
<< m1 >>
rect 146 346 147 347 
<< m2 >>
rect 146 346 147 347 
<< m1 >>
rect 147 346 148 347 
<< m2 >>
rect 147 346 148 347 
<< m1 >>
rect 148 346 149 347 
<< m2 >>
rect 148 346 149 347 
<< m1 >>
rect 149 346 150 347 
<< m2 >>
rect 149 346 150 347 
<< m1 >>
rect 150 346 151 347 
<< m2 >>
rect 150 346 151 347 
<< m1 >>
rect 151 346 152 347 
<< m2 >>
rect 151 346 152 347 
<< m1 >>
rect 152 346 153 347 
<< m2 >>
rect 152 346 153 347 
<< m1 >>
rect 153 346 154 347 
<< m2 >>
rect 153 346 154 347 
<< m1 >>
rect 154 346 155 347 
<< m2 >>
rect 154 346 155 347 
<< m1 >>
rect 155 346 156 347 
<< m2 >>
rect 155 346 156 347 
<< m1 >>
rect 156 346 157 347 
<< m2 >>
rect 156 346 157 347 
<< m1 >>
rect 157 346 158 347 
<< m2 >>
rect 157 346 158 347 
<< m1 >>
rect 158 346 159 347 
<< m2 >>
rect 158 346 159 347 
<< m1 >>
rect 159 346 160 347 
<< m2 >>
rect 159 346 160 347 
<< m1 >>
rect 160 346 161 347 
<< m2 >>
rect 160 346 161 347 
<< m1 >>
rect 161 346 162 347 
<< m2 >>
rect 161 346 162 347 
<< m1 >>
rect 162 346 163 347 
<< m2 >>
rect 162 346 163 347 
<< m1 >>
rect 163 346 164 347 
<< m2 >>
rect 163 346 164 347 
<< m1 >>
rect 164 346 165 347 
<< m2 >>
rect 164 346 165 347 
<< m1 >>
rect 165 346 166 347 
<< m2 >>
rect 165 346 166 347 
<< m1 >>
rect 166 346 167 347 
<< m2 >>
rect 166 346 167 347 
<< m1 >>
rect 167 346 168 347 
<< m2 >>
rect 167 346 168 347 
<< m1 >>
rect 168 346 169 347 
<< m2 >>
rect 168 346 169 347 
<< m1 >>
rect 169 346 170 347 
<< m2 >>
rect 169 346 170 347 
<< m1 >>
rect 170 346 171 347 
<< m2 >>
rect 170 346 171 347 
<< m1 >>
rect 171 346 172 347 
<< m2 >>
rect 171 346 172 347 
<< m1 >>
rect 172 346 173 347 
<< m2 >>
rect 172 346 173 347 
<< m1 >>
rect 173 346 174 347 
<< m2 >>
rect 173 346 174 347 
<< m1 >>
rect 174 346 175 347 
<< m2 >>
rect 174 346 175 347 
<< m1 >>
rect 175 346 176 347 
<< m2 >>
rect 175 346 176 347 
<< m1 >>
rect 176 346 177 347 
<< m2 >>
rect 176 346 177 347 
<< m1 >>
rect 177 346 178 347 
<< m2 >>
rect 177 346 178 347 
<< m1 >>
rect 178 346 179 347 
<< m2 >>
rect 178 346 179 347 
<< m1 >>
rect 179 346 180 347 
<< m2 >>
rect 179 346 180 347 
<< m1 >>
rect 180 346 181 347 
<< m2 >>
rect 180 346 181 347 
<< m1 >>
rect 181 346 182 347 
<< m2 >>
rect 181 346 182 347 
<< m1 >>
rect 182 346 183 347 
<< m2 >>
rect 182 346 183 347 
<< m1 >>
rect 183 346 184 347 
<< m2 >>
rect 183 346 184 347 
<< m1 >>
rect 184 346 185 347 
<< m2 >>
rect 184 346 185 347 
<< m1 >>
rect 185 346 186 347 
<< m2 >>
rect 185 346 186 347 
<< m1 >>
rect 186 346 187 347 
<< m2 >>
rect 186 346 187 347 
<< m1 >>
rect 187 346 188 347 
<< m2 >>
rect 187 346 188 347 
<< m1 >>
rect 188 346 189 347 
<< m2 >>
rect 188 346 189 347 
<< m1 >>
rect 189 346 190 347 
<< m2 >>
rect 189 346 190 347 
<< m1 >>
rect 190 346 191 347 
<< m2 >>
rect 190 346 191 347 
<< m1 >>
rect 191 346 192 347 
<< m2 >>
rect 191 346 192 347 
<< m1 >>
rect 192 346 193 347 
<< m2 >>
rect 192 346 193 347 
<< m1 >>
rect 193 346 194 347 
<< m2 >>
rect 193 346 194 347 
<< m1 >>
rect 194 346 195 347 
<< m2 >>
rect 194 346 195 347 
<< m1 >>
rect 195 346 196 347 
<< m2 >>
rect 195 346 196 347 
<< m1 >>
rect 196 346 197 347 
<< m2 >>
rect 196 346 197 347 
<< m1 >>
rect 197 346 198 347 
<< m2 >>
rect 197 346 198 347 
<< m1 >>
rect 198 346 199 347 
<< m2 >>
rect 198 346 199 347 
<< m1 >>
rect 199 346 200 347 
<< m2 >>
rect 199 346 200 347 
<< m1 >>
rect 200 346 201 347 
<< m2 >>
rect 200 346 201 347 
<< m1 >>
rect 201 346 202 347 
<< m2 >>
rect 201 346 202 347 
<< m1 >>
rect 202 346 203 347 
<< m2 >>
rect 202 346 203 347 
<< m1 >>
rect 203 346 204 347 
<< m2 >>
rect 203 346 204 347 
<< m1 >>
rect 204 346 205 347 
<< m2 >>
rect 204 346 205 347 
<< m1 >>
rect 205 346 206 347 
<< m2 >>
rect 205 346 206 347 
<< m1 >>
rect 206 346 207 347 
<< m2 >>
rect 206 346 207 347 
<< m1 >>
rect 207 346 208 347 
<< m2 >>
rect 207 346 208 347 
<< m1 >>
rect 208 346 209 347 
<< m2 >>
rect 208 346 209 347 
<< m1 >>
rect 209 346 210 347 
<< m2 >>
rect 209 346 210 347 
<< m1 >>
rect 210 346 211 347 
<< m2 >>
rect 210 346 211 347 
<< m1 >>
rect 211 346 212 347 
<< m2 >>
rect 211 346 212 347 
<< m1 >>
rect 212 346 213 347 
<< m2 >>
rect 212 346 213 347 
<< m1 >>
rect 213 346 214 347 
<< m2 >>
rect 213 346 214 347 
<< m1 >>
rect 214 346 215 347 
<< m2 >>
rect 214 346 215 347 
<< m1 >>
rect 215 346 216 347 
<< m2 >>
rect 215 346 216 347 
<< m1 >>
rect 216 346 217 347 
<< m2 >>
rect 216 346 217 347 
<< m1 >>
rect 217 346 218 347 
<< m2 >>
rect 217 346 218 347 
<< m1 >>
rect 218 346 219 347 
<< m2 >>
rect 218 346 219 347 
<< m1 >>
rect 219 346 220 347 
<< m2 >>
rect 219 346 220 347 
<< m2 >>
rect 220 346 221 347 
<< m1 >>
rect 221 346 222 347 
<< m2 >>
rect 221 346 222 347 
<< m2c >>
rect 221 346 222 347 
<< m1 >>
rect 221 346 222 347 
<< m2 >>
rect 221 346 222 347 
<< m1 >>
rect 223 346 224 347 
<< m2 >>
rect 223 346 224 347 
<< m2c >>
rect 223 346 224 347 
<< m1 >>
rect 223 346 224 347 
<< m2 >>
rect 223 346 224 347 
<< m1 >>
rect 239 346 240 347 
<< m1 >>
rect 240 346 241 347 
<< m1 >>
rect 241 346 242 347 
<< m1 >>
rect 242 346 243 347 
<< m1 >>
rect 243 346 244 347 
<< m1 >>
rect 244 346 245 347 
<< m1 >>
rect 245 346 246 347 
<< m1 >>
rect 246 346 247 347 
<< m1 >>
rect 247 346 248 347 
<< m1 >>
rect 248 346 249 347 
<< m1 >>
rect 249 346 250 347 
<< m1 >>
rect 250 346 251 347 
<< m1 >>
rect 251 346 252 347 
<< m1 >>
rect 252 346 253 347 
<< m1 >>
rect 253 346 254 347 
<< m1 >>
rect 254 346 255 347 
<< m1 >>
rect 255 346 256 347 
<< m1 >>
rect 256 346 257 347 
<< m1 >>
rect 257 346 258 347 
<< m1 >>
rect 258 346 259 347 
<< m1 >>
rect 259 346 260 347 
<< m1 >>
rect 260 346 261 347 
<< m1 >>
rect 261 346 262 347 
<< m1 >>
rect 262 346 263 347 
<< m1 >>
rect 263 346 264 347 
<< m1 >>
rect 264 346 265 347 
<< m1 >>
rect 265 346 266 347 
<< m1 >>
rect 266 346 267 347 
<< m1 >>
rect 267 346 268 347 
<< m1 >>
rect 268 346 269 347 
<< m1 >>
rect 269 346 270 347 
<< m1 >>
rect 270 346 271 347 
<< m1 >>
rect 271 346 272 347 
<< m1 >>
rect 272 346 273 347 
<< m1 >>
rect 273 346 274 347 
<< m1 >>
rect 274 346 275 347 
<< m1 >>
rect 275 346 276 347 
<< m1 >>
rect 276 346 277 347 
<< m1 >>
rect 277 346 278 347 
<< m1 >>
rect 278 346 279 347 
<< m1 >>
rect 279 346 280 347 
<< m1 >>
rect 280 346 281 347 
<< m1 >>
rect 281 346 282 347 
<< m1 >>
rect 282 346 283 347 
<< m1 >>
rect 283 346 284 347 
<< m1 >>
rect 284 346 285 347 
<< m1 >>
rect 285 346 286 347 
<< m1 >>
rect 286 346 287 347 
<< m1 >>
rect 287 346 288 347 
<< m1 >>
rect 288 346 289 347 
<< m1 >>
rect 289 346 290 347 
<< m1 >>
rect 290 346 291 347 
<< m1 >>
rect 291 346 292 347 
<< m1 >>
rect 292 346 293 347 
<< m1 >>
rect 293 346 294 347 
<< m1 >>
rect 294 346 295 347 
<< m1 >>
rect 295 346 296 347 
<< m1 >>
rect 296 346 297 347 
<< m1 >>
rect 297 346 298 347 
<< m1 >>
rect 298 346 299 347 
<< m1 >>
rect 299 346 300 347 
<< m1 >>
rect 300 346 301 347 
<< m1 >>
rect 301 346 302 347 
<< m1 >>
rect 302 346 303 347 
<< m2 >>
rect 302 346 303 347 
<< m2c >>
rect 302 346 303 347 
<< m1 >>
rect 302 346 303 347 
<< m2 >>
rect 302 346 303 347 
<< m2 >>
rect 303 346 304 347 
<< m1 >>
rect 304 346 305 347 
<< m2 >>
rect 304 346 305 347 
<< m2 >>
rect 305 346 306 347 
<< m1 >>
rect 306 346 307 347 
<< m2 >>
rect 306 346 307 347 
<< m2c >>
rect 306 346 307 347 
<< m1 >>
rect 306 346 307 347 
<< m2 >>
rect 306 346 307 347 
<< m1 >>
rect 307 346 308 347 
<< m1 >>
rect 325 346 326 347 
<< m2 >>
rect 326 346 327 347 
<< m1 >>
rect 331 346 332 347 
<< m2 >>
rect 332 346 333 347 
<< m1 >>
rect 334 346 335 347 
<< m1 >>
rect 340 346 341 347 
<< m1 >>
rect 343 346 344 347 
<< m1 >>
rect 10 347 11 348 
<< m2 >>
rect 26 347 27 348 
<< m2 >>
rect 28 347 29 348 
<< m2 >>
rect 46 347 47 348 
<< m2 >>
rect 48 347 49 348 
<< m2 >>
rect 49 347 50 348 
<< m2 >>
rect 50 347 51 348 
<< m2 >>
rect 51 347 52 348 
<< m2 >>
rect 52 347 53 348 
<< m2 >>
rect 53 347 54 348 
<< m2 >>
rect 54 347 55 348 
<< m2 >>
rect 56 347 57 348 
<< m2 >>
rect 58 347 59 348 
<< m2 >>
rect 62 347 63 348 
<< m2 >>
rect 66 347 67 348 
<< m2 >>
rect 223 347 224 348 
<< m1 >>
rect 304 347 305 348 
<< m1 >>
rect 325 347 326 348 
<< m2 >>
rect 326 347 327 348 
<< m1 >>
rect 331 347 332 348 
<< m2 >>
rect 332 347 333 348 
<< m1 >>
rect 334 347 335 348 
<< m1 >>
rect 340 347 341 348 
<< m1 >>
rect 343 347 344 348 
<< m1 >>
rect 10 348 11 349 
<< m1 >>
rect 24 348 25 349 
<< m1 >>
rect 25 348 26 349 
<< m1 >>
rect 26 348 27 349 
<< m2 >>
rect 26 348 27 349 
<< m2c >>
rect 26 348 27 349 
<< m1 >>
rect 26 348 27 349 
<< m2 >>
rect 26 348 27 349 
<< m1 >>
rect 28 348 29 349 
<< m2 >>
rect 28 348 29 349 
<< m2c >>
rect 28 348 29 349 
<< m1 >>
rect 28 348 29 349 
<< m2 >>
rect 28 348 29 349 
<< m1 >>
rect 46 348 47 349 
<< m2 >>
rect 46 348 47 349 
<< m2c >>
rect 46 348 47 349 
<< m1 >>
rect 46 348 47 349 
<< m2 >>
rect 46 348 47 349 
<< m1 >>
rect 54 348 55 349 
<< m2 >>
rect 54 348 55 349 
<< m2c >>
rect 54 348 55 349 
<< m1 >>
rect 54 348 55 349 
<< m2 >>
rect 54 348 55 349 
<< m1 >>
rect 56 348 57 349 
<< m2 >>
rect 56 348 57 349 
<< m2c >>
rect 56 348 57 349 
<< m1 >>
rect 56 348 57 349 
<< m2 >>
rect 56 348 57 349 
<< m1 >>
rect 58 348 59 349 
<< m2 >>
rect 58 348 59 349 
<< m2c >>
rect 58 348 59 349 
<< m1 >>
rect 58 348 59 349 
<< m2 >>
rect 58 348 59 349 
<< m1 >>
rect 62 348 63 349 
<< m2 >>
rect 62 348 63 349 
<< m2c >>
rect 62 348 63 349 
<< m1 >>
rect 62 348 63 349 
<< m2 >>
rect 62 348 63 349 
<< m1 >>
rect 63 348 64 349 
<< m1 >>
rect 64 348 65 349 
<< m1 >>
rect 65 348 66 349 
<< m1 >>
rect 66 348 67 349 
<< m2 >>
rect 66 348 67 349 
<< m1 >>
rect 67 348 68 349 
<< m2 >>
rect 67 348 68 349 
<< m1 >>
rect 68 348 69 349 
<< m2 >>
rect 68 348 69 349 
<< m1 >>
rect 69 348 70 349 
<< m2 >>
rect 69 348 70 349 
<< m1 >>
rect 70 348 71 349 
<< m2 >>
rect 70 348 71 349 
<< m1 >>
rect 71 348 72 349 
<< m2 >>
rect 71 348 72 349 
<< m1 >>
rect 72 348 73 349 
<< m2 >>
rect 72 348 73 349 
<< m1 >>
rect 73 348 74 349 
<< m2 >>
rect 73 348 74 349 
<< m1 >>
rect 74 348 75 349 
<< m2 >>
rect 74 348 75 349 
<< m1 >>
rect 75 348 76 349 
<< m2 >>
rect 75 348 76 349 
<< m1 >>
rect 76 348 77 349 
<< m2 >>
rect 76 348 77 349 
<< m1 >>
rect 77 348 78 349 
<< m2 >>
rect 77 348 78 349 
<< m1 >>
rect 78 348 79 349 
<< m2 >>
rect 78 348 79 349 
<< m1 >>
rect 79 348 80 349 
<< m2 >>
rect 79 348 80 349 
<< m1 >>
rect 80 348 81 349 
<< m2 >>
rect 80 348 81 349 
<< m1 >>
rect 81 348 82 349 
<< m2 >>
rect 81 348 82 349 
<< m1 >>
rect 82 348 83 349 
<< m2 >>
rect 82 348 83 349 
<< m1 >>
rect 83 348 84 349 
<< m2 >>
rect 83 348 84 349 
<< m1 >>
rect 84 348 85 349 
<< m2 >>
rect 84 348 85 349 
<< m1 >>
rect 85 348 86 349 
<< m2 >>
rect 85 348 86 349 
<< m1 >>
rect 86 348 87 349 
<< m2 >>
rect 86 348 87 349 
<< m1 >>
rect 87 348 88 349 
<< m2 >>
rect 87 348 88 349 
<< m1 >>
rect 88 348 89 349 
<< m2 >>
rect 88 348 89 349 
<< m1 >>
rect 89 348 90 349 
<< m2 >>
rect 89 348 90 349 
<< m1 >>
rect 90 348 91 349 
<< m2 >>
rect 90 348 91 349 
<< m1 >>
rect 91 348 92 349 
<< m2 >>
rect 91 348 92 349 
<< m1 >>
rect 92 348 93 349 
<< m2 >>
rect 92 348 93 349 
<< m1 >>
rect 93 348 94 349 
<< m2 >>
rect 93 348 94 349 
<< m1 >>
rect 94 348 95 349 
<< m2 >>
rect 94 348 95 349 
<< m1 >>
rect 95 348 96 349 
<< m2 >>
rect 95 348 96 349 
<< m1 >>
rect 96 348 97 349 
<< m2 >>
rect 96 348 97 349 
<< m1 >>
rect 97 348 98 349 
<< m2 >>
rect 97 348 98 349 
<< m1 >>
rect 98 348 99 349 
<< m2 >>
rect 98 348 99 349 
<< m1 >>
rect 99 348 100 349 
<< m2 >>
rect 99 348 100 349 
<< m1 >>
rect 100 348 101 349 
<< m2 >>
rect 100 348 101 349 
<< m1 >>
rect 101 348 102 349 
<< m2 >>
rect 101 348 102 349 
<< m1 >>
rect 102 348 103 349 
<< m2 >>
rect 102 348 103 349 
<< m1 >>
rect 103 348 104 349 
<< m2 >>
rect 103 348 104 349 
<< m1 >>
rect 104 348 105 349 
<< m2 >>
rect 104 348 105 349 
<< m1 >>
rect 105 348 106 349 
<< m2 >>
rect 105 348 106 349 
<< m1 >>
rect 106 348 107 349 
<< m2 >>
rect 106 348 107 349 
<< m1 >>
rect 107 348 108 349 
<< m2 >>
rect 107 348 108 349 
<< m1 >>
rect 108 348 109 349 
<< m2 >>
rect 108 348 109 349 
<< m1 >>
rect 109 348 110 349 
<< m2 >>
rect 109 348 110 349 
<< m1 >>
rect 110 348 111 349 
<< m2 >>
rect 110 348 111 349 
<< m1 >>
rect 111 348 112 349 
<< m2 >>
rect 111 348 112 349 
<< m1 >>
rect 112 348 113 349 
<< m2 >>
rect 112 348 113 349 
<< m1 >>
rect 113 348 114 349 
<< m2 >>
rect 113 348 114 349 
<< m1 >>
rect 114 348 115 349 
<< m2 >>
rect 114 348 115 349 
<< m1 >>
rect 115 348 116 349 
<< m2 >>
rect 115 348 116 349 
<< m1 >>
rect 116 348 117 349 
<< m2 >>
rect 116 348 117 349 
<< m1 >>
rect 117 348 118 349 
<< m2 >>
rect 117 348 118 349 
<< m1 >>
rect 118 348 119 349 
<< m2 >>
rect 118 348 119 349 
<< m1 >>
rect 119 348 120 349 
<< m2 >>
rect 119 348 120 349 
<< m1 >>
rect 120 348 121 349 
<< m2 >>
rect 120 348 121 349 
<< m1 >>
rect 121 348 122 349 
<< m2 >>
rect 121 348 122 349 
<< m1 >>
rect 122 348 123 349 
<< m2 >>
rect 122 348 123 349 
<< m1 >>
rect 123 348 124 349 
<< m2 >>
rect 123 348 124 349 
<< m1 >>
rect 124 348 125 349 
<< m2 >>
rect 124 348 125 349 
<< m1 >>
rect 125 348 126 349 
<< m2 >>
rect 125 348 126 349 
<< m1 >>
rect 126 348 127 349 
<< m2 >>
rect 126 348 127 349 
<< m1 >>
rect 127 348 128 349 
<< m2 >>
rect 127 348 128 349 
<< m1 >>
rect 128 348 129 349 
<< m2 >>
rect 128 348 129 349 
<< m1 >>
rect 129 348 130 349 
<< m2 >>
rect 129 348 130 349 
<< m1 >>
rect 130 348 131 349 
<< m2 >>
rect 130 348 131 349 
<< m1 >>
rect 131 348 132 349 
<< m2 >>
rect 131 348 132 349 
<< m1 >>
rect 132 348 133 349 
<< m2 >>
rect 132 348 133 349 
<< m1 >>
rect 133 348 134 349 
<< m2 >>
rect 133 348 134 349 
<< m1 >>
rect 134 348 135 349 
<< m2 >>
rect 134 348 135 349 
<< m1 >>
rect 135 348 136 349 
<< m2 >>
rect 135 348 136 349 
<< m1 >>
rect 136 348 137 349 
<< m2 >>
rect 136 348 137 349 
<< m1 >>
rect 137 348 138 349 
<< m2 >>
rect 137 348 138 349 
<< m1 >>
rect 138 348 139 349 
<< m2 >>
rect 138 348 139 349 
<< m1 >>
rect 139 348 140 349 
<< m2 >>
rect 139 348 140 349 
<< m1 >>
rect 140 348 141 349 
<< m2 >>
rect 140 348 141 349 
<< m1 >>
rect 141 348 142 349 
<< m2 >>
rect 141 348 142 349 
<< m1 >>
rect 142 348 143 349 
<< m2 >>
rect 142 348 143 349 
<< m1 >>
rect 143 348 144 349 
<< m2 >>
rect 143 348 144 349 
<< m1 >>
rect 144 348 145 349 
<< m2 >>
rect 144 348 145 349 
<< m1 >>
rect 145 348 146 349 
<< m2 >>
rect 145 348 146 349 
<< m1 >>
rect 146 348 147 349 
<< m2 >>
rect 146 348 147 349 
<< m1 >>
rect 147 348 148 349 
<< m2 >>
rect 147 348 148 349 
<< m1 >>
rect 148 348 149 349 
<< m2 >>
rect 148 348 149 349 
<< m1 >>
rect 149 348 150 349 
<< m2 >>
rect 149 348 150 349 
<< m1 >>
rect 150 348 151 349 
<< m2 >>
rect 150 348 151 349 
<< m1 >>
rect 151 348 152 349 
<< m2 >>
rect 151 348 152 349 
<< m1 >>
rect 152 348 153 349 
<< m2 >>
rect 152 348 153 349 
<< m1 >>
rect 153 348 154 349 
<< m2 >>
rect 153 348 154 349 
<< m1 >>
rect 154 348 155 349 
<< m2 >>
rect 154 348 155 349 
<< m1 >>
rect 155 348 156 349 
<< m2 >>
rect 155 348 156 349 
<< m1 >>
rect 156 348 157 349 
<< m2 >>
rect 156 348 157 349 
<< m1 >>
rect 157 348 158 349 
<< m2 >>
rect 157 348 158 349 
<< m1 >>
rect 158 348 159 349 
<< m2 >>
rect 158 348 159 349 
<< m1 >>
rect 159 348 160 349 
<< m2 >>
rect 159 348 160 349 
<< m1 >>
rect 160 348 161 349 
<< m2 >>
rect 160 348 161 349 
<< m1 >>
rect 161 348 162 349 
<< m2 >>
rect 161 348 162 349 
<< m1 >>
rect 162 348 163 349 
<< m2 >>
rect 162 348 163 349 
<< m1 >>
rect 163 348 164 349 
<< m2 >>
rect 163 348 164 349 
<< m1 >>
rect 164 348 165 349 
<< m2 >>
rect 164 348 165 349 
<< m1 >>
rect 165 348 166 349 
<< m2 >>
rect 165 348 166 349 
<< m1 >>
rect 166 348 167 349 
<< m2 >>
rect 166 348 167 349 
<< m1 >>
rect 167 348 168 349 
<< m2 >>
rect 167 348 168 349 
<< m1 >>
rect 168 348 169 349 
<< m2 >>
rect 168 348 169 349 
<< m1 >>
rect 169 348 170 349 
<< m2 >>
rect 169 348 170 349 
<< m1 >>
rect 170 348 171 349 
<< m2 >>
rect 170 348 171 349 
<< m1 >>
rect 171 348 172 349 
<< m2 >>
rect 171 348 172 349 
<< m1 >>
rect 172 348 173 349 
<< m2 >>
rect 172 348 173 349 
<< m1 >>
rect 173 348 174 349 
<< m2 >>
rect 173 348 174 349 
<< m1 >>
rect 174 348 175 349 
<< m2 >>
rect 174 348 175 349 
<< m1 >>
rect 175 348 176 349 
<< m2 >>
rect 175 348 176 349 
<< m1 >>
rect 176 348 177 349 
<< m2 >>
rect 176 348 177 349 
<< m1 >>
rect 177 348 178 349 
<< m2 >>
rect 177 348 178 349 
<< m1 >>
rect 178 348 179 349 
<< m2 >>
rect 178 348 179 349 
<< m1 >>
rect 179 348 180 349 
<< m2 >>
rect 179 348 180 349 
<< m1 >>
rect 180 348 181 349 
<< m2 >>
rect 180 348 181 349 
<< m1 >>
rect 181 348 182 349 
<< m2 >>
rect 181 348 182 349 
<< m1 >>
rect 182 348 183 349 
<< m2 >>
rect 182 348 183 349 
<< m1 >>
rect 183 348 184 349 
<< m2 >>
rect 183 348 184 349 
<< m1 >>
rect 184 348 185 349 
<< m2 >>
rect 184 348 185 349 
<< m1 >>
rect 185 348 186 349 
<< m2 >>
rect 185 348 186 349 
<< m1 >>
rect 186 348 187 349 
<< m2 >>
rect 186 348 187 349 
<< m1 >>
rect 187 348 188 349 
<< m2 >>
rect 187 348 188 349 
<< m1 >>
rect 188 348 189 349 
<< m2 >>
rect 188 348 189 349 
<< m1 >>
rect 189 348 190 349 
<< m2 >>
rect 189 348 190 349 
<< m1 >>
rect 190 348 191 349 
<< m2 >>
rect 190 348 191 349 
<< m1 >>
rect 191 348 192 349 
<< m2 >>
rect 191 348 192 349 
<< m1 >>
rect 192 348 193 349 
<< m2 >>
rect 192 348 193 349 
<< m1 >>
rect 193 348 194 349 
<< m2 >>
rect 193 348 194 349 
<< m1 >>
rect 194 348 195 349 
<< m2 >>
rect 194 348 195 349 
<< m1 >>
rect 195 348 196 349 
<< m2 >>
rect 195 348 196 349 
<< m1 >>
rect 196 348 197 349 
<< m2 >>
rect 196 348 197 349 
<< m1 >>
rect 197 348 198 349 
<< m2 >>
rect 197 348 198 349 
<< m1 >>
rect 198 348 199 349 
<< m2 >>
rect 198 348 199 349 
<< m1 >>
rect 199 348 200 349 
<< m2 >>
rect 199 348 200 349 
<< m1 >>
rect 200 348 201 349 
<< m2 >>
rect 200 348 201 349 
<< m1 >>
rect 201 348 202 349 
<< m2 >>
rect 201 348 202 349 
<< m1 >>
rect 202 348 203 349 
<< m2 >>
rect 202 348 203 349 
<< m1 >>
rect 203 348 204 349 
<< m2 >>
rect 203 348 204 349 
<< m1 >>
rect 204 348 205 349 
<< m2 >>
rect 204 348 205 349 
<< m1 >>
rect 205 348 206 349 
<< m2 >>
rect 205 348 206 349 
<< m1 >>
rect 206 348 207 349 
<< m2 >>
rect 206 348 207 349 
<< m1 >>
rect 207 348 208 349 
<< m2 >>
rect 207 348 208 349 
<< m1 >>
rect 208 348 209 349 
<< m2 >>
rect 208 348 209 349 
<< m1 >>
rect 209 348 210 349 
<< m2 >>
rect 209 348 210 349 
<< m1 >>
rect 210 348 211 349 
<< m2 >>
rect 210 348 211 349 
<< m1 >>
rect 211 348 212 349 
<< m2 >>
rect 211 348 212 349 
<< m1 >>
rect 212 348 213 349 
<< m2 >>
rect 212 348 213 349 
<< m1 >>
rect 213 348 214 349 
<< m2 >>
rect 213 348 214 349 
<< m1 >>
rect 214 348 215 349 
<< m2 >>
rect 214 348 215 349 
<< m1 >>
rect 215 348 216 349 
<< m2 >>
rect 215 348 216 349 
<< m1 >>
rect 216 348 217 349 
<< m2 >>
rect 216 348 217 349 
<< m1 >>
rect 217 348 218 349 
<< m2 >>
rect 217 348 218 349 
<< m1 >>
rect 218 348 219 349 
<< m2 >>
rect 218 348 219 349 
<< m1 >>
rect 219 348 220 349 
<< m2 >>
rect 219 348 220 349 
<< m1 >>
rect 220 348 221 349 
<< m2 >>
rect 220 348 221 349 
<< m1 >>
rect 221 348 222 349 
<< m2 >>
rect 221 348 222 349 
<< m1 >>
rect 222 348 223 349 
<< m2 >>
rect 222 348 223 349 
<< m1 >>
rect 223 348 224 349 
<< m2 >>
rect 223 348 224 349 
<< m1 >>
rect 224 348 225 349 
<< m1 >>
rect 225 348 226 349 
<< m1 >>
rect 226 348 227 349 
<< m1 >>
rect 227 348 228 349 
<< m1 >>
rect 228 348 229 349 
<< m1 >>
rect 229 348 230 349 
<< m1 >>
rect 230 348 231 349 
<< m1 >>
rect 231 348 232 349 
<< m1 >>
rect 232 348 233 349 
<< m1 >>
rect 233 348 234 349 
<< m1 >>
rect 234 348 235 349 
<< m1 >>
rect 235 348 236 349 
<< m1 >>
rect 236 348 237 349 
<< m1 >>
rect 237 348 238 349 
<< m1 >>
rect 238 348 239 349 
<< m1 >>
rect 239 348 240 349 
<< m1 >>
rect 240 348 241 349 
<< m1 >>
rect 241 348 242 349 
<< m1 >>
rect 242 348 243 349 
<< m1 >>
rect 243 348 244 349 
<< m1 >>
rect 244 348 245 349 
<< m1 >>
rect 245 348 246 349 
<< m1 >>
rect 246 348 247 349 
<< m1 >>
rect 247 348 248 349 
<< m1 >>
rect 248 348 249 349 
<< m1 >>
rect 249 348 250 349 
<< m1 >>
rect 250 348 251 349 
<< m1 >>
rect 251 348 252 349 
<< m1 >>
rect 252 348 253 349 
<< m1 >>
rect 253 348 254 349 
<< m1 >>
rect 254 348 255 349 
<< m1 >>
rect 255 348 256 349 
<< m1 >>
rect 256 348 257 349 
<< m1 >>
rect 257 348 258 349 
<< m1 >>
rect 258 348 259 349 
<< m1 >>
rect 259 348 260 349 
<< m1 >>
rect 260 348 261 349 
<< m1 >>
rect 261 348 262 349 
<< m1 >>
rect 262 348 263 349 
<< m1 >>
rect 263 348 264 349 
<< m1 >>
rect 264 348 265 349 
<< m1 >>
rect 265 348 266 349 
<< m1 >>
rect 266 348 267 349 
<< m1 >>
rect 267 348 268 349 
<< m1 >>
rect 268 348 269 349 
<< m1 >>
rect 269 348 270 349 
<< m1 >>
rect 270 348 271 349 
<< m1 >>
rect 271 348 272 349 
<< m1 >>
rect 272 348 273 349 
<< m1 >>
rect 273 348 274 349 
<< m1 >>
rect 274 348 275 349 
<< m1 >>
rect 275 348 276 349 
<< m1 >>
rect 276 348 277 349 
<< m1 >>
rect 277 348 278 349 
<< m1 >>
rect 278 348 279 349 
<< m1 >>
rect 279 348 280 349 
<< m1 >>
rect 280 348 281 349 
<< m1 >>
rect 281 348 282 349 
<< m1 >>
rect 282 348 283 349 
<< m1 >>
rect 283 348 284 349 
<< m1 >>
rect 284 348 285 349 
<< m1 >>
rect 285 348 286 349 
<< m1 >>
rect 286 348 287 349 
<< m1 >>
rect 287 348 288 349 
<< m1 >>
rect 288 348 289 349 
<< m1 >>
rect 289 348 290 349 
<< m1 >>
rect 290 348 291 349 
<< m1 >>
rect 291 348 292 349 
<< m1 >>
rect 292 348 293 349 
<< m1 >>
rect 293 348 294 349 
<< m1 >>
rect 294 348 295 349 
<< m1 >>
rect 295 348 296 349 
<< m1 >>
rect 296 348 297 349 
<< m1 >>
rect 297 348 298 349 
<< m1 >>
rect 298 348 299 349 
<< m1 >>
rect 299 348 300 349 
<< m1 >>
rect 300 348 301 349 
<< m1 >>
rect 301 348 302 349 
<< m1 >>
rect 302 348 303 349 
<< m1 >>
rect 303 348 304 349 
<< m1 >>
rect 304 348 305 349 
<< m1 >>
rect 325 348 326 349 
<< m2 >>
rect 326 348 327 349 
<< m1 >>
rect 331 348 332 349 
<< m2 >>
rect 332 348 333 349 
<< m1 >>
rect 334 348 335 349 
<< m1 >>
rect 340 348 341 349 
<< m1 >>
rect 343 348 344 349 
<< m1 >>
rect 10 349 11 350 
<< m1 >>
rect 24 349 25 350 
<< m1 >>
rect 28 349 29 350 
<< m1 >>
rect 46 349 47 350 
<< m1 >>
rect 54 349 55 350 
<< m1 >>
rect 56 349 57 350 
<< m1 >>
rect 58 349 59 350 
<< m1 >>
rect 325 349 326 350 
<< m2 >>
rect 326 349 327 350 
<< m1 >>
rect 331 349 332 350 
<< m2 >>
rect 332 349 333 350 
<< m1 >>
rect 334 349 335 350 
<< m1 >>
rect 340 349 341 350 
<< m1 >>
rect 343 349 344 350 
<< m1 >>
rect 10 350 11 351 
<< m1 >>
rect 24 350 25 351 
<< m1 >>
rect 28 350 29 351 
<< m1 >>
rect 46 350 47 351 
<< m1 >>
rect 54 350 55 351 
<< m1 >>
rect 56 350 57 351 
<< m2 >>
rect 56 350 57 351 
<< m2c >>
rect 56 350 57 351 
<< m1 >>
rect 56 350 57 351 
<< m2 >>
rect 56 350 57 351 
<< m2 >>
rect 57 350 58 351 
<< m1 >>
rect 58 350 59 351 
<< m2 >>
rect 58 350 59 351 
<< m1 >>
rect 59 350 60 351 
<< m2 >>
rect 59 350 60 351 
<< m1 >>
rect 60 350 61 351 
<< m2 >>
rect 60 350 61 351 
<< m1 >>
rect 61 350 62 351 
<< m2 >>
rect 61 350 62 351 
<< m1 >>
rect 62 350 63 351 
<< m2 >>
rect 62 350 63 351 
<< m1 >>
rect 63 350 64 351 
<< m2 >>
rect 63 350 64 351 
<< m1 >>
rect 64 350 65 351 
<< m2 >>
rect 64 350 65 351 
<< m1 >>
rect 65 350 66 351 
<< m2 >>
rect 65 350 66 351 
<< m1 >>
rect 66 350 67 351 
<< m2 >>
rect 66 350 67 351 
<< m1 >>
rect 67 350 68 351 
<< m2 >>
rect 67 350 68 351 
<< m1 >>
rect 68 350 69 351 
<< m2 >>
rect 68 350 69 351 
<< m1 >>
rect 69 350 70 351 
<< m2 >>
rect 69 350 70 351 
<< m1 >>
rect 70 350 71 351 
<< m2 >>
rect 70 350 71 351 
<< m1 >>
rect 71 350 72 351 
<< m2 >>
rect 71 350 72 351 
<< m1 >>
rect 72 350 73 351 
<< m2 >>
rect 72 350 73 351 
<< m1 >>
rect 73 350 74 351 
<< m2 >>
rect 73 350 74 351 
<< m1 >>
rect 74 350 75 351 
<< m2 >>
rect 74 350 75 351 
<< m1 >>
rect 75 350 76 351 
<< m2 >>
rect 75 350 76 351 
<< m1 >>
rect 76 350 77 351 
<< m2 >>
rect 76 350 77 351 
<< m1 >>
rect 77 350 78 351 
<< m2 >>
rect 77 350 78 351 
<< m1 >>
rect 78 350 79 351 
<< m2 >>
rect 78 350 79 351 
<< m1 >>
rect 79 350 80 351 
<< m2 >>
rect 79 350 80 351 
<< m1 >>
rect 80 350 81 351 
<< m2 >>
rect 80 350 81 351 
<< m1 >>
rect 81 350 82 351 
<< m2 >>
rect 81 350 82 351 
<< m1 >>
rect 82 350 83 351 
<< m2 >>
rect 82 350 83 351 
<< m1 >>
rect 83 350 84 351 
<< m2 >>
rect 83 350 84 351 
<< m1 >>
rect 84 350 85 351 
<< m2 >>
rect 84 350 85 351 
<< m1 >>
rect 85 350 86 351 
<< m2 >>
rect 85 350 86 351 
<< m1 >>
rect 86 350 87 351 
<< m2 >>
rect 86 350 87 351 
<< m1 >>
rect 87 350 88 351 
<< m2 >>
rect 87 350 88 351 
<< m1 >>
rect 88 350 89 351 
<< m2 >>
rect 88 350 89 351 
<< m1 >>
rect 89 350 90 351 
<< m2 >>
rect 89 350 90 351 
<< m1 >>
rect 90 350 91 351 
<< m2 >>
rect 90 350 91 351 
<< m1 >>
rect 91 350 92 351 
<< m2 >>
rect 91 350 92 351 
<< m1 >>
rect 92 350 93 351 
<< m2 >>
rect 92 350 93 351 
<< m1 >>
rect 93 350 94 351 
<< m2 >>
rect 93 350 94 351 
<< m1 >>
rect 94 350 95 351 
<< m2 >>
rect 94 350 95 351 
<< m1 >>
rect 95 350 96 351 
<< m2 >>
rect 95 350 96 351 
<< m1 >>
rect 96 350 97 351 
<< m2 >>
rect 96 350 97 351 
<< m1 >>
rect 97 350 98 351 
<< m2 >>
rect 97 350 98 351 
<< m1 >>
rect 98 350 99 351 
<< m2 >>
rect 98 350 99 351 
<< m1 >>
rect 99 350 100 351 
<< m2 >>
rect 99 350 100 351 
<< m1 >>
rect 100 350 101 351 
<< m2 >>
rect 100 350 101 351 
<< m1 >>
rect 101 350 102 351 
<< m2 >>
rect 101 350 102 351 
<< m1 >>
rect 102 350 103 351 
<< m2 >>
rect 102 350 103 351 
<< m1 >>
rect 103 350 104 351 
<< m2 >>
rect 103 350 104 351 
<< m1 >>
rect 104 350 105 351 
<< m2 >>
rect 104 350 105 351 
<< m1 >>
rect 105 350 106 351 
<< m2 >>
rect 105 350 106 351 
<< m1 >>
rect 106 350 107 351 
<< m2 >>
rect 106 350 107 351 
<< m1 >>
rect 107 350 108 351 
<< m2 >>
rect 107 350 108 351 
<< m1 >>
rect 108 350 109 351 
<< m2 >>
rect 108 350 109 351 
<< m1 >>
rect 109 350 110 351 
<< m2 >>
rect 109 350 110 351 
<< m1 >>
rect 110 350 111 351 
<< m2 >>
rect 110 350 111 351 
<< m1 >>
rect 111 350 112 351 
<< m2 >>
rect 111 350 112 351 
<< m1 >>
rect 112 350 113 351 
<< m2 >>
rect 112 350 113 351 
<< m1 >>
rect 113 350 114 351 
<< m2 >>
rect 113 350 114 351 
<< m1 >>
rect 114 350 115 351 
<< m2 >>
rect 114 350 115 351 
<< m1 >>
rect 115 350 116 351 
<< m2 >>
rect 115 350 116 351 
<< m1 >>
rect 116 350 117 351 
<< m2 >>
rect 116 350 117 351 
<< m1 >>
rect 117 350 118 351 
<< m2 >>
rect 117 350 118 351 
<< m1 >>
rect 118 350 119 351 
<< m2 >>
rect 118 350 119 351 
<< m1 >>
rect 119 350 120 351 
<< m2 >>
rect 119 350 120 351 
<< m1 >>
rect 120 350 121 351 
<< m2 >>
rect 120 350 121 351 
<< m1 >>
rect 121 350 122 351 
<< m2 >>
rect 121 350 122 351 
<< m1 >>
rect 122 350 123 351 
<< m2 >>
rect 122 350 123 351 
<< m1 >>
rect 123 350 124 351 
<< m2 >>
rect 123 350 124 351 
<< m1 >>
rect 124 350 125 351 
<< m2 >>
rect 124 350 125 351 
<< m1 >>
rect 125 350 126 351 
<< m2 >>
rect 125 350 126 351 
<< m1 >>
rect 126 350 127 351 
<< m2 >>
rect 126 350 127 351 
<< m1 >>
rect 127 350 128 351 
<< m2 >>
rect 127 350 128 351 
<< m1 >>
rect 128 350 129 351 
<< m2 >>
rect 128 350 129 351 
<< m1 >>
rect 129 350 130 351 
<< m2 >>
rect 129 350 130 351 
<< m1 >>
rect 130 350 131 351 
<< m2 >>
rect 130 350 131 351 
<< m1 >>
rect 131 350 132 351 
<< m2 >>
rect 131 350 132 351 
<< m1 >>
rect 132 350 133 351 
<< m2 >>
rect 132 350 133 351 
<< m1 >>
rect 133 350 134 351 
<< m2 >>
rect 133 350 134 351 
<< m1 >>
rect 134 350 135 351 
<< m2 >>
rect 134 350 135 351 
<< m1 >>
rect 135 350 136 351 
<< m2 >>
rect 135 350 136 351 
<< m1 >>
rect 136 350 137 351 
<< m2 >>
rect 136 350 137 351 
<< m1 >>
rect 137 350 138 351 
<< m2 >>
rect 137 350 138 351 
<< m1 >>
rect 138 350 139 351 
<< m2 >>
rect 138 350 139 351 
<< m1 >>
rect 139 350 140 351 
<< m2 >>
rect 139 350 140 351 
<< m1 >>
rect 140 350 141 351 
<< m2 >>
rect 140 350 141 351 
<< m1 >>
rect 141 350 142 351 
<< m2 >>
rect 141 350 142 351 
<< m1 >>
rect 142 350 143 351 
<< m2 >>
rect 142 350 143 351 
<< m1 >>
rect 143 350 144 351 
<< m2 >>
rect 143 350 144 351 
<< m1 >>
rect 144 350 145 351 
<< m2 >>
rect 144 350 145 351 
<< m1 >>
rect 145 350 146 351 
<< m2 >>
rect 145 350 146 351 
<< m1 >>
rect 146 350 147 351 
<< m2 >>
rect 146 350 147 351 
<< m1 >>
rect 147 350 148 351 
<< m2 >>
rect 147 350 148 351 
<< m1 >>
rect 148 350 149 351 
<< m2 >>
rect 148 350 149 351 
<< m1 >>
rect 149 350 150 351 
<< m2 >>
rect 149 350 150 351 
<< m1 >>
rect 150 350 151 351 
<< m2 >>
rect 150 350 151 351 
<< m1 >>
rect 151 350 152 351 
<< m2 >>
rect 151 350 152 351 
<< m1 >>
rect 152 350 153 351 
<< m2 >>
rect 152 350 153 351 
<< m1 >>
rect 153 350 154 351 
<< m2 >>
rect 153 350 154 351 
<< m1 >>
rect 154 350 155 351 
<< m2 >>
rect 154 350 155 351 
<< m1 >>
rect 155 350 156 351 
<< m2 >>
rect 155 350 156 351 
<< m1 >>
rect 156 350 157 351 
<< m2 >>
rect 156 350 157 351 
<< m1 >>
rect 157 350 158 351 
<< m2 >>
rect 157 350 158 351 
<< m1 >>
rect 158 350 159 351 
<< m2 >>
rect 158 350 159 351 
<< m1 >>
rect 159 350 160 351 
<< m2 >>
rect 159 350 160 351 
<< m1 >>
rect 160 350 161 351 
<< m2 >>
rect 160 350 161 351 
<< m1 >>
rect 161 350 162 351 
<< m2 >>
rect 161 350 162 351 
<< m1 >>
rect 162 350 163 351 
<< m2 >>
rect 162 350 163 351 
<< m1 >>
rect 163 350 164 351 
<< m2 >>
rect 163 350 164 351 
<< m1 >>
rect 164 350 165 351 
<< m2 >>
rect 164 350 165 351 
<< m1 >>
rect 165 350 166 351 
<< m2 >>
rect 165 350 166 351 
<< m1 >>
rect 166 350 167 351 
<< m2 >>
rect 166 350 167 351 
<< m1 >>
rect 167 350 168 351 
<< m2 >>
rect 167 350 168 351 
<< m1 >>
rect 168 350 169 351 
<< m2 >>
rect 168 350 169 351 
<< m1 >>
rect 169 350 170 351 
<< m2 >>
rect 169 350 170 351 
<< m1 >>
rect 170 350 171 351 
<< m2 >>
rect 170 350 171 351 
<< m1 >>
rect 171 350 172 351 
<< m2 >>
rect 171 350 172 351 
<< m1 >>
rect 172 350 173 351 
<< m2 >>
rect 172 350 173 351 
<< m1 >>
rect 173 350 174 351 
<< m2 >>
rect 173 350 174 351 
<< m1 >>
rect 174 350 175 351 
<< m2 >>
rect 174 350 175 351 
<< m1 >>
rect 175 350 176 351 
<< m2 >>
rect 175 350 176 351 
<< m1 >>
rect 176 350 177 351 
<< m2 >>
rect 176 350 177 351 
<< m1 >>
rect 177 350 178 351 
<< m2 >>
rect 177 350 178 351 
<< m1 >>
rect 178 350 179 351 
<< m2 >>
rect 178 350 179 351 
<< m1 >>
rect 179 350 180 351 
<< m2 >>
rect 179 350 180 351 
<< m1 >>
rect 180 350 181 351 
<< m2 >>
rect 180 350 181 351 
<< m1 >>
rect 181 350 182 351 
<< m2 >>
rect 181 350 182 351 
<< m1 >>
rect 182 350 183 351 
<< m2 >>
rect 182 350 183 351 
<< m1 >>
rect 183 350 184 351 
<< m2 >>
rect 183 350 184 351 
<< m1 >>
rect 184 350 185 351 
<< m2 >>
rect 184 350 185 351 
<< m1 >>
rect 185 350 186 351 
<< m2 >>
rect 185 350 186 351 
<< m1 >>
rect 186 350 187 351 
<< m2 >>
rect 186 350 187 351 
<< m1 >>
rect 187 350 188 351 
<< m2 >>
rect 187 350 188 351 
<< m1 >>
rect 188 350 189 351 
<< m2 >>
rect 188 350 189 351 
<< m1 >>
rect 189 350 190 351 
<< m2 >>
rect 189 350 190 351 
<< m1 >>
rect 190 350 191 351 
<< m2 >>
rect 190 350 191 351 
<< m1 >>
rect 191 350 192 351 
<< m2 >>
rect 191 350 192 351 
<< m1 >>
rect 192 350 193 351 
<< m2 >>
rect 192 350 193 351 
<< m1 >>
rect 193 350 194 351 
<< m2 >>
rect 193 350 194 351 
<< m1 >>
rect 194 350 195 351 
<< m2 >>
rect 194 350 195 351 
<< m1 >>
rect 195 350 196 351 
<< m2 >>
rect 195 350 196 351 
<< m1 >>
rect 196 350 197 351 
<< m2 >>
rect 196 350 197 351 
<< m1 >>
rect 197 350 198 351 
<< m2 >>
rect 197 350 198 351 
<< m1 >>
rect 198 350 199 351 
<< m2 >>
rect 198 350 199 351 
<< m1 >>
rect 199 350 200 351 
<< m2 >>
rect 199 350 200 351 
<< m1 >>
rect 200 350 201 351 
<< m2 >>
rect 200 350 201 351 
<< m1 >>
rect 201 350 202 351 
<< m2 >>
rect 201 350 202 351 
<< m1 >>
rect 202 350 203 351 
<< m2 >>
rect 202 350 203 351 
<< m1 >>
rect 203 350 204 351 
<< m2 >>
rect 203 350 204 351 
<< m1 >>
rect 204 350 205 351 
<< m2 >>
rect 204 350 205 351 
<< m1 >>
rect 205 350 206 351 
<< m2 >>
rect 205 350 206 351 
<< m1 >>
rect 206 350 207 351 
<< m2 >>
rect 206 350 207 351 
<< m1 >>
rect 207 350 208 351 
<< m2 >>
rect 207 350 208 351 
<< m1 >>
rect 208 350 209 351 
<< m2 >>
rect 208 350 209 351 
<< m1 >>
rect 209 350 210 351 
<< m2 >>
rect 209 350 210 351 
<< m1 >>
rect 210 350 211 351 
<< m2 >>
rect 210 350 211 351 
<< m1 >>
rect 211 350 212 351 
<< m2 >>
rect 211 350 212 351 
<< m1 >>
rect 212 350 213 351 
<< m2 >>
rect 212 350 213 351 
<< m1 >>
rect 213 350 214 351 
<< m2 >>
rect 213 350 214 351 
<< m1 >>
rect 214 350 215 351 
<< m2 >>
rect 214 350 215 351 
<< m1 >>
rect 215 350 216 351 
<< m2 >>
rect 215 350 216 351 
<< m1 >>
rect 216 350 217 351 
<< m2 >>
rect 216 350 217 351 
<< m1 >>
rect 217 350 218 351 
<< m2 >>
rect 217 350 218 351 
<< m1 >>
rect 218 350 219 351 
<< m2 >>
rect 218 350 219 351 
<< m1 >>
rect 219 350 220 351 
<< m2 >>
rect 219 350 220 351 
<< m1 >>
rect 220 350 221 351 
<< m2 >>
rect 220 350 221 351 
<< m1 >>
rect 221 350 222 351 
<< m2 >>
rect 221 350 222 351 
<< m1 >>
rect 222 350 223 351 
<< m2 >>
rect 222 350 223 351 
<< m1 >>
rect 223 350 224 351 
<< m2 >>
rect 223 350 224 351 
<< m1 >>
rect 224 350 225 351 
<< m2 >>
rect 224 350 225 351 
<< m1 >>
rect 225 350 226 351 
<< m2 >>
rect 225 350 226 351 
<< m1 >>
rect 226 350 227 351 
<< m2 >>
rect 226 350 227 351 
<< m1 >>
rect 227 350 228 351 
<< m2 >>
rect 227 350 228 351 
<< m1 >>
rect 228 350 229 351 
<< m2 >>
rect 228 350 229 351 
<< m1 >>
rect 229 350 230 351 
<< m2 >>
rect 229 350 230 351 
<< m1 >>
rect 230 350 231 351 
<< m2 >>
rect 230 350 231 351 
<< m1 >>
rect 231 350 232 351 
<< m2 >>
rect 231 350 232 351 
<< m1 >>
rect 232 350 233 351 
<< m2 >>
rect 232 350 233 351 
<< m1 >>
rect 233 350 234 351 
<< m2 >>
rect 233 350 234 351 
<< m1 >>
rect 234 350 235 351 
<< m2 >>
rect 234 350 235 351 
<< m1 >>
rect 235 350 236 351 
<< m2 >>
rect 235 350 236 351 
<< m1 >>
rect 236 350 237 351 
<< m2 >>
rect 236 350 237 351 
<< m1 >>
rect 237 350 238 351 
<< m2 >>
rect 237 350 238 351 
<< m1 >>
rect 238 350 239 351 
<< m2 >>
rect 238 350 239 351 
<< m1 >>
rect 239 350 240 351 
<< m2 >>
rect 239 350 240 351 
<< m1 >>
rect 240 350 241 351 
<< m2 >>
rect 240 350 241 351 
<< m1 >>
rect 241 350 242 351 
<< m2 >>
rect 241 350 242 351 
<< m1 >>
rect 242 350 243 351 
<< m2 >>
rect 242 350 243 351 
<< m1 >>
rect 243 350 244 351 
<< m2 >>
rect 243 350 244 351 
<< m1 >>
rect 244 350 245 351 
<< m2 >>
rect 244 350 245 351 
<< m1 >>
rect 245 350 246 351 
<< m2 >>
rect 245 350 246 351 
<< m1 >>
rect 246 350 247 351 
<< m2 >>
rect 246 350 247 351 
<< m1 >>
rect 247 350 248 351 
<< m2 >>
rect 247 350 248 351 
<< m1 >>
rect 248 350 249 351 
<< m2 >>
rect 248 350 249 351 
<< m1 >>
rect 249 350 250 351 
<< m2 >>
rect 249 350 250 351 
<< m1 >>
rect 250 350 251 351 
<< m2 >>
rect 250 350 251 351 
<< m1 >>
rect 251 350 252 351 
<< m2 >>
rect 251 350 252 351 
<< m1 >>
rect 252 350 253 351 
<< m2 >>
rect 252 350 253 351 
<< m1 >>
rect 253 350 254 351 
<< m2 >>
rect 253 350 254 351 
<< m1 >>
rect 254 350 255 351 
<< m2 >>
rect 254 350 255 351 
<< m1 >>
rect 255 350 256 351 
<< m2 >>
rect 255 350 256 351 
<< m1 >>
rect 256 350 257 351 
<< m2 >>
rect 256 350 257 351 
<< m1 >>
rect 257 350 258 351 
<< m2 >>
rect 257 350 258 351 
<< m1 >>
rect 258 350 259 351 
<< m2 >>
rect 258 350 259 351 
<< m1 >>
rect 259 350 260 351 
<< m2 >>
rect 259 350 260 351 
<< m1 >>
rect 260 350 261 351 
<< m2 >>
rect 260 350 261 351 
<< m1 >>
rect 261 350 262 351 
<< m2 >>
rect 261 350 262 351 
<< m1 >>
rect 262 350 263 351 
<< m2 >>
rect 262 350 263 351 
<< m1 >>
rect 263 350 264 351 
<< m2 >>
rect 263 350 264 351 
<< m1 >>
rect 264 350 265 351 
<< m2 >>
rect 264 350 265 351 
<< m1 >>
rect 265 350 266 351 
<< m2 >>
rect 265 350 266 351 
<< m1 >>
rect 266 350 267 351 
<< m2 >>
rect 266 350 267 351 
<< m1 >>
rect 267 350 268 351 
<< m2 >>
rect 267 350 268 351 
<< m1 >>
rect 268 350 269 351 
<< m2 >>
rect 268 350 269 351 
<< m1 >>
rect 269 350 270 351 
<< m2 >>
rect 269 350 270 351 
<< m1 >>
rect 270 350 271 351 
<< m2 >>
rect 270 350 271 351 
<< m1 >>
rect 271 350 272 351 
<< m2 >>
rect 271 350 272 351 
<< m1 >>
rect 272 350 273 351 
<< m2 >>
rect 272 350 273 351 
<< m1 >>
rect 273 350 274 351 
<< m2 >>
rect 273 350 274 351 
<< m1 >>
rect 274 350 275 351 
<< m2 >>
rect 274 350 275 351 
<< m1 >>
rect 275 350 276 351 
<< m2 >>
rect 275 350 276 351 
<< m1 >>
rect 276 350 277 351 
<< m2 >>
rect 276 350 277 351 
<< m1 >>
rect 277 350 278 351 
<< m2 >>
rect 277 350 278 351 
<< m1 >>
rect 278 350 279 351 
<< m2 >>
rect 278 350 279 351 
<< m1 >>
rect 279 350 280 351 
<< m2 >>
rect 279 350 280 351 
<< m1 >>
rect 280 350 281 351 
<< m2 >>
rect 280 350 281 351 
<< m1 >>
rect 281 350 282 351 
<< m2 >>
rect 281 350 282 351 
<< m1 >>
rect 282 350 283 351 
<< m2 >>
rect 282 350 283 351 
<< m1 >>
rect 283 350 284 351 
<< m2 >>
rect 283 350 284 351 
<< m1 >>
rect 284 350 285 351 
<< m2 >>
rect 284 350 285 351 
<< m1 >>
rect 285 350 286 351 
<< m2 >>
rect 285 350 286 351 
<< m1 >>
rect 286 350 287 351 
<< m2 >>
rect 286 350 287 351 
<< m1 >>
rect 287 350 288 351 
<< m2 >>
rect 287 350 288 351 
<< m1 >>
rect 288 350 289 351 
<< m2 >>
rect 288 350 289 351 
<< m1 >>
rect 289 350 290 351 
<< m2 >>
rect 289 350 290 351 
<< m1 >>
rect 290 350 291 351 
<< m2 >>
rect 290 350 291 351 
<< m1 >>
rect 291 350 292 351 
<< m2 >>
rect 291 350 292 351 
<< m1 >>
rect 292 350 293 351 
<< m2 >>
rect 292 350 293 351 
<< m1 >>
rect 293 350 294 351 
<< m2 >>
rect 293 350 294 351 
<< m1 >>
rect 294 350 295 351 
<< m2 >>
rect 294 350 295 351 
<< m1 >>
rect 295 350 296 351 
<< m2 >>
rect 295 350 296 351 
<< m1 >>
rect 296 350 297 351 
<< m2 >>
rect 296 350 297 351 
<< m1 >>
rect 297 350 298 351 
<< m2 >>
rect 297 350 298 351 
<< m1 >>
rect 298 350 299 351 
<< m2 >>
rect 298 350 299 351 
<< m1 >>
rect 299 350 300 351 
<< m2 >>
rect 299 350 300 351 
<< m1 >>
rect 300 350 301 351 
<< m2 >>
rect 300 350 301 351 
<< m1 >>
rect 301 350 302 351 
<< m2 >>
rect 301 350 302 351 
<< m1 >>
rect 302 350 303 351 
<< m2 >>
rect 302 350 303 351 
<< m1 >>
rect 303 350 304 351 
<< m2 >>
rect 303 350 304 351 
<< m1 >>
rect 304 350 305 351 
<< m2 >>
rect 304 350 305 351 
<< m1 >>
rect 305 350 306 351 
<< m2 >>
rect 305 350 306 351 
<< m1 >>
rect 306 350 307 351 
<< m2 >>
rect 306 350 307 351 
<< m1 >>
rect 307 350 308 351 
<< m2 >>
rect 307 350 308 351 
<< m1 >>
rect 308 350 309 351 
<< m2 >>
rect 308 350 309 351 
<< m1 >>
rect 309 350 310 351 
<< m2 >>
rect 309 350 310 351 
<< m1 >>
rect 310 350 311 351 
<< m2 >>
rect 310 350 311 351 
<< m1 >>
rect 311 350 312 351 
<< m2 >>
rect 311 350 312 351 
<< m1 >>
rect 312 350 313 351 
<< m2 >>
rect 312 350 313 351 
<< m1 >>
rect 313 350 314 351 
<< m2 >>
rect 313 350 314 351 
<< m1 >>
rect 314 350 315 351 
<< m2 >>
rect 314 350 315 351 
<< m1 >>
rect 315 350 316 351 
<< m2 >>
rect 315 350 316 351 
<< m1 >>
rect 316 350 317 351 
<< m2 >>
rect 316 350 317 351 
<< m1 >>
rect 317 350 318 351 
<< m2 >>
rect 317 350 318 351 
<< m1 >>
rect 318 350 319 351 
<< m2 >>
rect 318 350 319 351 
<< m1 >>
rect 319 350 320 351 
<< m2 >>
rect 319 350 320 351 
<< m1 >>
rect 320 350 321 351 
<< m2 >>
rect 320 350 321 351 
<< m1 >>
rect 321 350 322 351 
<< m2 >>
rect 321 350 322 351 
<< m1 >>
rect 322 350 323 351 
<< m2 >>
rect 322 350 323 351 
<< m1 >>
rect 323 350 324 351 
<< m2 >>
rect 323 350 324 351 
<< m1 >>
rect 324 350 325 351 
<< m2 >>
rect 324 350 325 351 
<< m1 >>
rect 325 350 326 351 
<< m2 >>
rect 325 350 326 351 
<< m2 >>
rect 326 350 327 351 
<< m1 >>
rect 331 350 332 351 
<< m2 >>
rect 332 350 333 351 
<< m1 >>
rect 334 350 335 351 
<< m1 >>
rect 340 350 341 351 
<< m1 >>
rect 343 350 344 351 
<< m1 >>
rect 10 351 11 352 
<< m1 >>
rect 24 351 25 352 
<< m1 >>
rect 28 351 29 352 
<< m1 >>
rect 46 351 47 352 
<< m1 >>
rect 54 351 55 352 
<< m1 >>
rect 331 351 332 352 
<< m2 >>
rect 332 351 333 352 
<< m1 >>
rect 334 351 335 352 
<< m1 >>
rect 340 351 341 352 
<< m1 >>
rect 343 351 344 352 
<< m1 >>
rect 10 352 11 353 
<< m1 >>
rect 24 352 25 353 
<< m2 >>
rect 24 352 25 353 
<< m2c >>
rect 24 352 25 353 
<< m1 >>
rect 24 352 25 353 
<< m2 >>
rect 24 352 25 353 
<< m1 >>
rect 28 352 29 353 
<< m1 >>
rect 46 352 47 353 
<< m1 >>
rect 47 352 48 353 
<< m1 >>
rect 48 352 49 353 
<< m1 >>
rect 49 352 50 353 
<< m1 >>
rect 50 352 51 353 
<< m1 >>
rect 51 352 52 353 
<< m1 >>
rect 52 352 53 353 
<< m2 >>
rect 52 352 53 353 
<< m2c >>
rect 52 352 53 353 
<< m1 >>
rect 52 352 53 353 
<< m2 >>
rect 52 352 53 353 
<< m2 >>
rect 53 352 54 353 
<< m1 >>
rect 54 352 55 353 
<< m2 >>
rect 54 352 55 353 
<< m1 >>
rect 55 352 56 353 
<< m2 >>
rect 55 352 56 353 
<< m1 >>
rect 56 352 57 353 
<< m2 >>
rect 56 352 57 353 
<< m1 >>
rect 57 352 58 353 
<< m2 >>
rect 57 352 58 353 
<< m1 >>
rect 58 352 59 353 
<< m2 >>
rect 58 352 59 353 
<< m1 >>
rect 59 352 60 353 
<< m2 >>
rect 59 352 60 353 
<< m1 >>
rect 60 352 61 353 
<< m2 >>
rect 60 352 61 353 
<< m1 >>
rect 61 352 62 353 
<< m2 >>
rect 61 352 62 353 
<< m1 >>
rect 62 352 63 353 
<< m2 >>
rect 62 352 63 353 
<< m1 >>
rect 63 352 64 353 
<< m2 >>
rect 63 352 64 353 
<< m1 >>
rect 64 352 65 353 
<< m2 >>
rect 64 352 65 353 
<< m1 >>
rect 65 352 66 353 
<< m2 >>
rect 65 352 66 353 
<< m1 >>
rect 66 352 67 353 
<< m2 >>
rect 66 352 67 353 
<< m1 >>
rect 67 352 68 353 
<< m2 >>
rect 67 352 68 353 
<< m1 >>
rect 68 352 69 353 
<< m2 >>
rect 68 352 69 353 
<< m1 >>
rect 69 352 70 353 
<< m2 >>
rect 69 352 70 353 
<< m1 >>
rect 70 352 71 353 
<< m2 >>
rect 70 352 71 353 
<< m1 >>
rect 71 352 72 353 
<< m2 >>
rect 71 352 72 353 
<< m1 >>
rect 72 352 73 353 
<< m2 >>
rect 72 352 73 353 
<< m1 >>
rect 73 352 74 353 
<< m2 >>
rect 73 352 74 353 
<< m1 >>
rect 74 352 75 353 
<< m2 >>
rect 74 352 75 353 
<< m1 >>
rect 75 352 76 353 
<< m2 >>
rect 75 352 76 353 
<< m1 >>
rect 76 352 77 353 
<< m2 >>
rect 76 352 77 353 
<< m1 >>
rect 77 352 78 353 
<< m2 >>
rect 77 352 78 353 
<< m1 >>
rect 78 352 79 353 
<< m2 >>
rect 78 352 79 353 
<< m1 >>
rect 79 352 80 353 
<< m2 >>
rect 79 352 80 353 
<< m1 >>
rect 80 352 81 353 
<< m2 >>
rect 80 352 81 353 
<< m1 >>
rect 81 352 82 353 
<< m2 >>
rect 81 352 82 353 
<< m1 >>
rect 82 352 83 353 
<< m2 >>
rect 82 352 83 353 
<< m1 >>
rect 83 352 84 353 
<< m2 >>
rect 83 352 84 353 
<< m1 >>
rect 84 352 85 353 
<< m2 >>
rect 84 352 85 353 
<< m1 >>
rect 85 352 86 353 
<< m2 >>
rect 85 352 86 353 
<< m1 >>
rect 86 352 87 353 
<< m2 >>
rect 86 352 87 353 
<< m1 >>
rect 87 352 88 353 
<< m2 >>
rect 87 352 88 353 
<< m1 >>
rect 88 352 89 353 
<< m2 >>
rect 88 352 89 353 
<< m1 >>
rect 89 352 90 353 
<< m2 >>
rect 89 352 90 353 
<< m1 >>
rect 90 352 91 353 
<< m2 >>
rect 90 352 91 353 
<< m1 >>
rect 91 352 92 353 
<< m2 >>
rect 91 352 92 353 
<< m1 >>
rect 92 352 93 353 
<< m2 >>
rect 92 352 93 353 
<< m1 >>
rect 93 352 94 353 
<< m2 >>
rect 93 352 94 353 
<< m1 >>
rect 94 352 95 353 
<< m2 >>
rect 94 352 95 353 
<< m1 >>
rect 95 352 96 353 
<< m2 >>
rect 95 352 96 353 
<< m1 >>
rect 96 352 97 353 
<< m2 >>
rect 96 352 97 353 
<< m1 >>
rect 97 352 98 353 
<< m2 >>
rect 97 352 98 353 
<< m1 >>
rect 98 352 99 353 
<< m2 >>
rect 98 352 99 353 
<< m1 >>
rect 99 352 100 353 
<< m2 >>
rect 99 352 100 353 
<< m1 >>
rect 100 352 101 353 
<< m2 >>
rect 100 352 101 353 
<< m1 >>
rect 101 352 102 353 
<< m2 >>
rect 101 352 102 353 
<< m1 >>
rect 102 352 103 353 
<< m2 >>
rect 102 352 103 353 
<< m1 >>
rect 103 352 104 353 
<< m2 >>
rect 103 352 104 353 
<< m1 >>
rect 104 352 105 353 
<< m2 >>
rect 104 352 105 353 
<< m1 >>
rect 105 352 106 353 
<< m2 >>
rect 105 352 106 353 
<< m1 >>
rect 106 352 107 353 
<< m2 >>
rect 106 352 107 353 
<< m1 >>
rect 107 352 108 353 
<< m2 >>
rect 107 352 108 353 
<< m1 >>
rect 108 352 109 353 
<< m2 >>
rect 108 352 109 353 
<< m1 >>
rect 109 352 110 353 
<< m2 >>
rect 109 352 110 353 
<< m1 >>
rect 110 352 111 353 
<< m2 >>
rect 110 352 111 353 
<< m1 >>
rect 111 352 112 353 
<< m2 >>
rect 111 352 112 353 
<< m1 >>
rect 112 352 113 353 
<< m2 >>
rect 112 352 113 353 
<< m1 >>
rect 113 352 114 353 
<< m2 >>
rect 113 352 114 353 
<< m1 >>
rect 114 352 115 353 
<< m2 >>
rect 114 352 115 353 
<< m1 >>
rect 115 352 116 353 
<< m2 >>
rect 115 352 116 353 
<< m1 >>
rect 116 352 117 353 
<< m2 >>
rect 116 352 117 353 
<< m1 >>
rect 117 352 118 353 
<< m2 >>
rect 117 352 118 353 
<< m1 >>
rect 118 352 119 353 
<< m2 >>
rect 118 352 119 353 
<< m1 >>
rect 119 352 120 353 
<< m2 >>
rect 119 352 120 353 
<< m1 >>
rect 120 352 121 353 
<< m2 >>
rect 120 352 121 353 
<< m1 >>
rect 121 352 122 353 
<< m2 >>
rect 121 352 122 353 
<< m1 >>
rect 122 352 123 353 
<< m2 >>
rect 122 352 123 353 
<< m1 >>
rect 123 352 124 353 
<< m2 >>
rect 123 352 124 353 
<< m1 >>
rect 124 352 125 353 
<< m2 >>
rect 124 352 125 353 
<< m1 >>
rect 125 352 126 353 
<< m2 >>
rect 125 352 126 353 
<< m1 >>
rect 126 352 127 353 
<< m2 >>
rect 126 352 127 353 
<< m1 >>
rect 127 352 128 353 
<< m2 >>
rect 127 352 128 353 
<< m1 >>
rect 128 352 129 353 
<< m2 >>
rect 128 352 129 353 
<< m1 >>
rect 129 352 130 353 
<< m2 >>
rect 129 352 130 353 
<< m1 >>
rect 130 352 131 353 
<< m2 >>
rect 130 352 131 353 
<< m1 >>
rect 131 352 132 353 
<< m2 >>
rect 131 352 132 353 
<< m1 >>
rect 132 352 133 353 
<< m2 >>
rect 132 352 133 353 
<< m1 >>
rect 133 352 134 353 
<< m2 >>
rect 133 352 134 353 
<< m1 >>
rect 134 352 135 353 
<< m2 >>
rect 134 352 135 353 
<< m1 >>
rect 135 352 136 353 
<< m2 >>
rect 135 352 136 353 
<< m1 >>
rect 136 352 137 353 
<< m2 >>
rect 136 352 137 353 
<< m1 >>
rect 137 352 138 353 
<< m2 >>
rect 137 352 138 353 
<< m1 >>
rect 138 352 139 353 
<< m2 >>
rect 138 352 139 353 
<< m1 >>
rect 139 352 140 353 
<< m2 >>
rect 139 352 140 353 
<< m1 >>
rect 140 352 141 353 
<< m2 >>
rect 140 352 141 353 
<< m1 >>
rect 141 352 142 353 
<< m2 >>
rect 141 352 142 353 
<< m1 >>
rect 142 352 143 353 
<< m2 >>
rect 142 352 143 353 
<< m1 >>
rect 143 352 144 353 
<< m2 >>
rect 143 352 144 353 
<< m1 >>
rect 144 352 145 353 
<< m2 >>
rect 144 352 145 353 
<< m1 >>
rect 145 352 146 353 
<< m2 >>
rect 145 352 146 353 
<< m1 >>
rect 146 352 147 353 
<< m2 >>
rect 146 352 147 353 
<< m1 >>
rect 147 352 148 353 
<< m2 >>
rect 147 352 148 353 
<< m1 >>
rect 148 352 149 353 
<< m2 >>
rect 148 352 149 353 
<< m1 >>
rect 149 352 150 353 
<< m2 >>
rect 149 352 150 353 
<< m1 >>
rect 150 352 151 353 
<< m2 >>
rect 150 352 151 353 
<< m1 >>
rect 151 352 152 353 
<< m2 >>
rect 151 352 152 353 
<< m1 >>
rect 152 352 153 353 
<< m2 >>
rect 152 352 153 353 
<< m1 >>
rect 153 352 154 353 
<< m2 >>
rect 153 352 154 353 
<< m1 >>
rect 154 352 155 353 
<< m2 >>
rect 154 352 155 353 
<< m1 >>
rect 155 352 156 353 
<< m2 >>
rect 155 352 156 353 
<< m1 >>
rect 156 352 157 353 
<< m2 >>
rect 156 352 157 353 
<< m1 >>
rect 157 352 158 353 
<< m2 >>
rect 157 352 158 353 
<< m1 >>
rect 158 352 159 353 
<< m2 >>
rect 158 352 159 353 
<< m1 >>
rect 159 352 160 353 
<< m2 >>
rect 159 352 160 353 
<< m1 >>
rect 160 352 161 353 
<< m2 >>
rect 160 352 161 353 
<< m1 >>
rect 161 352 162 353 
<< m2 >>
rect 161 352 162 353 
<< m1 >>
rect 162 352 163 353 
<< m2 >>
rect 162 352 163 353 
<< m1 >>
rect 163 352 164 353 
<< m2 >>
rect 163 352 164 353 
<< m1 >>
rect 164 352 165 353 
<< m2 >>
rect 164 352 165 353 
<< m1 >>
rect 165 352 166 353 
<< m2 >>
rect 165 352 166 353 
<< m1 >>
rect 166 352 167 353 
<< m2 >>
rect 166 352 167 353 
<< m1 >>
rect 167 352 168 353 
<< m2 >>
rect 167 352 168 353 
<< m1 >>
rect 168 352 169 353 
<< m2 >>
rect 168 352 169 353 
<< m1 >>
rect 169 352 170 353 
<< m2 >>
rect 169 352 170 353 
<< m1 >>
rect 170 352 171 353 
<< m2 >>
rect 170 352 171 353 
<< m1 >>
rect 171 352 172 353 
<< m2 >>
rect 171 352 172 353 
<< m1 >>
rect 172 352 173 353 
<< m2 >>
rect 172 352 173 353 
<< m1 >>
rect 173 352 174 353 
<< m2 >>
rect 173 352 174 353 
<< m1 >>
rect 174 352 175 353 
<< m2 >>
rect 174 352 175 353 
<< m1 >>
rect 175 352 176 353 
<< m2 >>
rect 175 352 176 353 
<< m1 >>
rect 176 352 177 353 
<< m2 >>
rect 176 352 177 353 
<< m1 >>
rect 177 352 178 353 
<< m2 >>
rect 177 352 178 353 
<< m1 >>
rect 178 352 179 353 
<< m2 >>
rect 178 352 179 353 
<< m1 >>
rect 179 352 180 353 
<< m2 >>
rect 179 352 180 353 
<< m1 >>
rect 180 352 181 353 
<< m2 >>
rect 180 352 181 353 
<< m1 >>
rect 181 352 182 353 
<< m2 >>
rect 181 352 182 353 
<< m1 >>
rect 182 352 183 353 
<< m2 >>
rect 182 352 183 353 
<< m1 >>
rect 183 352 184 353 
<< m2 >>
rect 183 352 184 353 
<< m1 >>
rect 184 352 185 353 
<< m2 >>
rect 184 352 185 353 
<< m1 >>
rect 185 352 186 353 
<< m2 >>
rect 185 352 186 353 
<< m1 >>
rect 186 352 187 353 
<< m2 >>
rect 186 352 187 353 
<< m1 >>
rect 187 352 188 353 
<< m2 >>
rect 187 352 188 353 
<< m1 >>
rect 188 352 189 353 
<< m2 >>
rect 188 352 189 353 
<< m1 >>
rect 189 352 190 353 
<< m2 >>
rect 189 352 190 353 
<< m1 >>
rect 190 352 191 353 
<< m2 >>
rect 190 352 191 353 
<< m1 >>
rect 191 352 192 353 
<< m2 >>
rect 191 352 192 353 
<< m1 >>
rect 192 352 193 353 
<< m2 >>
rect 192 352 193 353 
<< m1 >>
rect 193 352 194 353 
<< m2 >>
rect 193 352 194 353 
<< m1 >>
rect 194 352 195 353 
<< m2 >>
rect 194 352 195 353 
<< m1 >>
rect 195 352 196 353 
<< m2 >>
rect 195 352 196 353 
<< m1 >>
rect 196 352 197 353 
<< m2 >>
rect 196 352 197 353 
<< m1 >>
rect 197 352 198 353 
<< m2 >>
rect 197 352 198 353 
<< m1 >>
rect 198 352 199 353 
<< m2 >>
rect 198 352 199 353 
<< m1 >>
rect 199 352 200 353 
<< m2 >>
rect 199 352 200 353 
<< m1 >>
rect 200 352 201 353 
<< m2 >>
rect 200 352 201 353 
<< m1 >>
rect 201 352 202 353 
<< m2 >>
rect 201 352 202 353 
<< m1 >>
rect 202 352 203 353 
<< m2 >>
rect 202 352 203 353 
<< m1 >>
rect 203 352 204 353 
<< m2 >>
rect 203 352 204 353 
<< m1 >>
rect 204 352 205 353 
<< m2 >>
rect 204 352 205 353 
<< m1 >>
rect 205 352 206 353 
<< m2 >>
rect 205 352 206 353 
<< m1 >>
rect 206 352 207 353 
<< m2 >>
rect 206 352 207 353 
<< m1 >>
rect 207 352 208 353 
<< m2 >>
rect 207 352 208 353 
<< m1 >>
rect 208 352 209 353 
<< m2 >>
rect 208 352 209 353 
<< m1 >>
rect 209 352 210 353 
<< m2 >>
rect 209 352 210 353 
<< m1 >>
rect 210 352 211 353 
<< m2 >>
rect 210 352 211 353 
<< m1 >>
rect 211 352 212 353 
<< m2 >>
rect 211 352 212 353 
<< m1 >>
rect 212 352 213 353 
<< m2 >>
rect 212 352 213 353 
<< m1 >>
rect 213 352 214 353 
<< m2 >>
rect 213 352 214 353 
<< m1 >>
rect 214 352 215 353 
<< m2 >>
rect 214 352 215 353 
<< m1 >>
rect 215 352 216 353 
<< m2 >>
rect 215 352 216 353 
<< m1 >>
rect 216 352 217 353 
<< m2 >>
rect 216 352 217 353 
<< m1 >>
rect 217 352 218 353 
<< m2 >>
rect 217 352 218 353 
<< m1 >>
rect 218 352 219 353 
<< m2 >>
rect 218 352 219 353 
<< m1 >>
rect 219 352 220 353 
<< m2 >>
rect 219 352 220 353 
<< m1 >>
rect 220 352 221 353 
<< m2 >>
rect 220 352 221 353 
<< m1 >>
rect 221 352 222 353 
<< m2 >>
rect 221 352 222 353 
<< m1 >>
rect 222 352 223 353 
<< m2 >>
rect 222 352 223 353 
<< m1 >>
rect 223 352 224 353 
<< m2 >>
rect 223 352 224 353 
<< m1 >>
rect 224 352 225 353 
<< m2 >>
rect 224 352 225 353 
<< m1 >>
rect 225 352 226 353 
<< m2 >>
rect 225 352 226 353 
<< m1 >>
rect 226 352 227 353 
<< m2 >>
rect 226 352 227 353 
<< m1 >>
rect 227 352 228 353 
<< m2 >>
rect 227 352 228 353 
<< m1 >>
rect 228 352 229 353 
<< m2 >>
rect 228 352 229 353 
<< m1 >>
rect 229 352 230 353 
<< m2 >>
rect 229 352 230 353 
<< m1 >>
rect 230 352 231 353 
<< m2 >>
rect 230 352 231 353 
<< m1 >>
rect 231 352 232 353 
<< m2 >>
rect 231 352 232 353 
<< m1 >>
rect 232 352 233 353 
<< m2 >>
rect 232 352 233 353 
<< m1 >>
rect 233 352 234 353 
<< m2 >>
rect 233 352 234 353 
<< m1 >>
rect 234 352 235 353 
<< m2 >>
rect 234 352 235 353 
<< m1 >>
rect 235 352 236 353 
<< m2 >>
rect 235 352 236 353 
<< m1 >>
rect 236 352 237 353 
<< m2 >>
rect 236 352 237 353 
<< m1 >>
rect 237 352 238 353 
<< m2 >>
rect 237 352 238 353 
<< m1 >>
rect 238 352 239 353 
<< m2 >>
rect 238 352 239 353 
<< m1 >>
rect 239 352 240 353 
<< m2 >>
rect 239 352 240 353 
<< m1 >>
rect 240 352 241 353 
<< m2 >>
rect 240 352 241 353 
<< m1 >>
rect 241 352 242 353 
<< m2 >>
rect 241 352 242 353 
<< m1 >>
rect 242 352 243 353 
<< m2 >>
rect 242 352 243 353 
<< m1 >>
rect 243 352 244 353 
<< m2 >>
rect 243 352 244 353 
<< m1 >>
rect 244 352 245 353 
<< m2 >>
rect 244 352 245 353 
<< m1 >>
rect 245 352 246 353 
<< m2 >>
rect 245 352 246 353 
<< m1 >>
rect 246 352 247 353 
<< m2 >>
rect 246 352 247 353 
<< m1 >>
rect 247 352 248 353 
<< m2 >>
rect 247 352 248 353 
<< m1 >>
rect 248 352 249 353 
<< m2 >>
rect 248 352 249 353 
<< m1 >>
rect 249 352 250 353 
<< m2 >>
rect 249 352 250 353 
<< m1 >>
rect 250 352 251 353 
<< m2 >>
rect 250 352 251 353 
<< m1 >>
rect 251 352 252 353 
<< m2 >>
rect 251 352 252 353 
<< m1 >>
rect 252 352 253 353 
<< m2 >>
rect 252 352 253 353 
<< m1 >>
rect 253 352 254 353 
<< m2 >>
rect 253 352 254 353 
<< m1 >>
rect 254 352 255 353 
<< m2 >>
rect 254 352 255 353 
<< m1 >>
rect 255 352 256 353 
<< m2 >>
rect 255 352 256 353 
<< m1 >>
rect 256 352 257 353 
<< m2 >>
rect 256 352 257 353 
<< m1 >>
rect 257 352 258 353 
<< m2 >>
rect 257 352 258 353 
<< m1 >>
rect 258 352 259 353 
<< m2 >>
rect 258 352 259 353 
<< m1 >>
rect 259 352 260 353 
<< m2 >>
rect 259 352 260 353 
<< m1 >>
rect 260 352 261 353 
<< m2 >>
rect 260 352 261 353 
<< m1 >>
rect 261 352 262 353 
<< m2 >>
rect 261 352 262 353 
<< m1 >>
rect 262 352 263 353 
<< m2 >>
rect 262 352 263 353 
<< m1 >>
rect 263 352 264 353 
<< m2 >>
rect 263 352 264 353 
<< m1 >>
rect 264 352 265 353 
<< m2 >>
rect 264 352 265 353 
<< m1 >>
rect 265 352 266 353 
<< m2 >>
rect 265 352 266 353 
<< m1 >>
rect 266 352 267 353 
<< m2 >>
rect 266 352 267 353 
<< m1 >>
rect 267 352 268 353 
<< m2 >>
rect 267 352 268 353 
<< m1 >>
rect 268 352 269 353 
<< m2 >>
rect 268 352 269 353 
<< m1 >>
rect 269 352 270 353 
<< m2 >>
rect 269 352 270 353 
<< m1 >>
rect 270 352 271 353 
<< m2 >>
rect 270 352 271 353 
<< m1 >>
rect 271 352 272 353 
<< m2 >>
rect 271 352 272 353 
<< m1 >>
rect 272 352 273 353 
<< m2 >>
rect 272 352 273 353 
<< m1 >>
rect 273 352 274 353 
<< m2 >>
rect 273 352 274 353 
<< m1 >>
rect 274 352 275 353 
<< m2 >>
rect 274 352 275 353 
<< m1 >>
rect 275 352 276 353 
<< m2 >>
rect 275 352 276 353 
<< m1 >>
rect 276 352 277 353 
<< m2 >>
rect 276 352 277 353 
<< m1 >>
rect 277 352 278 353 
<< m2 >>
rect 277 352 278 353 
<< m1 >>
rect 278 352 279 353 
<< m2 >>
rect 278 352 279 353 
<< m1 >>
rect 279 352 280 353 
<< m2 >>
rect 279 352 280 353 
<< m1 >>
rect 280 352 281 353 
<< m2 >>
rect 280 352 281 353 
<< m1 >>
rect 281 352 282 353 
<< m2 >>
rect 281 352 282 353 
<< m1 >>
rect 282 352 283 353 
<< m2 >>
rect 282 352 283 353 
<< m1 >>
rect 283 352 284 353 
<< m2 >>
rect 283 352 284 353 
<< m1 >>
rect 284 352 285 353 
<< m2 >>
rect 284 352 285 353 
<< m1 >>
rect 285 352 286 353 
<< m2 >>
rect 285 352 286 353 
<< m1 >>
rect 286 352 287 353 
<< m2 >>
rect 286 352 287 353 
<< m1 >>
rect 287 352 288 353 
<< m2 >>
rect 287 352 288 353 
<< m1 >>
rect 288 352 289 353 
<< m2 >>
rect 288 352 289 353 
<< m1 >>
rect 289 352 290 353 
<< m2 >>
rect 289 352 290 353 
<< m1 >>
rect 290 352 291 353 
<< m2 >>
rect 290 352 291 353 
<< m1 >>
rect 291 352 292 353 
<< m2 >>
rect 291 352 292 353 
<< m1 >>
rect 292 352 293 353 
<< m2 >>
rect 292 352 293 353 
<< m1 >>
rect 293 352 294 353 
<< m2 >>
rect 293 352 294 353 
<< m1 >>
rect 294 352 295 353 
<< m2 >>
rect 294 352 295 353 
<< m1 >>
rect 295 352 296 353 
<< m2 >>
rect 295 352 296 353 
<< m1 >>
rect 296 352 297 353 
<< m2 >>
rect 296 352 297 353 
<< m1 >>
rect 297 352 298 353 
<< m2 >>
rect 297 352 298 353 
<< m1 >>
rect 298 352 299 353 
<< m2 >>
rect 298 352 299 353 
<< m1 >>
rect 299 352 300 353 
<< m2 >>
rect 299 352 300 353 
<< m1 >>
rect 300 352 301 353 
<< m2 >>
rect 300 352 301 353 
<< m1 >>
rect 301 352 302 353 
<< m2 >>
rect 301 352 302 353 
<< m1 >>
rect 302 352 303 353 
<< m2 >>
rect 302 352 303 353 
<< m1 >>
rect 303 352 304 353 
<< m2 >>
rect 303 352 304 353 
<< m1 >>
rect 304 352 305 353 
<< m2 >>
rect 304 352 305 353 
<< m1 >>
rect 305 352 306 353 
<< m2 >>
rect 305 352 306 353 
<< m1 >>
rect 306 352 307 353 
<< m2 >>
rect 306 352 307 353 
<< m1 >>
rect 307 352 308 353 
<< m2 >>
rect 307 352 308 353 
<< m1 >>
rect 308 352 309 353 
<< m2 >>
rect 308 352 309 353 
<< m1 >>
rect 309 352 310 353 
<< m2 >>
rect 309 352 310 353 
<< m1 >>
rect 310 352 311 353 
<< m2 >>
rect 310 352 311 353 
<< m1 >>
rect 311 352 312 353 
<< m2 >>
rect 311 352 312 353 
<< m1 >>
rect 312 352 313 353 
<< m2 >>
rect 312 352 313 353 
<< m1 >>
rect 313 352 314 353 
<< m2 >>
rect 313 352 314 353 
<< m1 >>
rect 314 352 315 353 
<< m2 >>
rect 314 352 315 353 
<< m1 >>
rect 315 352 316 353 
<< m2 >>
rect 315 352 316 353 
<< m1 >>
rect 316 352 317 353 
<< m2 >>
rect 316 352 317 353 
<< m1 >>
rect 317 352 318 353 
<< m2 >>
rect 317 352 318 353 
<< m1 >>
rect 318 352 319 353 
<< m2 >>
rect 318 352 319 353 
<< m1 >>
rect 319 352 320 353 
<< m2 >>
rect 319 352 320 353 
<< m1 >>
rect 320 352 321 353 
<< m2 >>
rect 320 352 321 353 
<< m1 >>
rect 321 352 322 353 
<< m2 >>
rect 321 352 322 353 
<< m1 >>
rect 322 352 323 353 
<< m2 >>
rect 322 352 323 353 
<< m1 >>
rect 323 352 324 353 
<< m2 >>
rect 323 352 324 353 
<< m1 >>
rect 324 352 325 353 
<< m2 >>
rect 324 352 325 353 
<< m1 >>
rect 325 352 326 353 
<< m2 >>
rect 325 352 326 353 
<< m1 >>
rect 326 352 327 353 
<< m2 >>
rect 326 352 327 353 
<< m1 >>
rect 327 352 328 353 
<< m2 >>
rect 327 352 328 353 
<< m1 >>
rect 328 352 329 353 
<< m2 >>
rect 328 352 329 353 
<< m1 >>
rect 329 352 330 353 
<< m2 >>
rect 329 352 330 353 
<< m1 >>
rect 330 352 331 353 
<< m2 >>
rect 330 352 331 353 
<< m1 >>
rect 331 352 332 353 
<< m2 >>
rect 331 352 332 353 
<< m2 >>
rect 332 352 333 353 
<< m1 >>
rect 334 352 335 353 
<< m2 >>
rect 334 352 335 353 
<< m2c >>
rect 334 352 335 353 
<< m1 >>
rect 334 352 335 353 
<< m2 >>
rect 334 352 335 353 
<< m1 >>
rect 340 352 341 353 
<< m1 >>
rect 343 352 344 353 
<< m1 >>
rect 10 353 11 354 
<< m2 >>
rect 24 353 25 354 
<< m1 >>
rect 28 353 29 354 
<< m2 >>
rect 334 353 335 354 
<< m1 >>
rect 340 353 341 354 
<< m1 >>
rect 343 353 344 354 
<< m1 >>
rect 10 354 11 355 
<< m1 >>
rect 11 354 12 355 
<< m1 >>
rect 12 354 13 355 
<< m1 >>
rect 13 354 14 355 
<< m1 >>
rect 14 354 15 355 
<< m1 >>
rect 15 354 16 355 
<< m1 >>
rect 16 354 17 355 
<< m1 >>
rect 17 354 18 355 
<< m1 >>
rect 18 354 19 355 
<< m1 >>
rect 19 354 20 355 
<< m1 >>
rect 20 354 21 355 
<< m1 >>
rect 21 354 22 355 
<< m1 >>
rect 22 354 23 355 
<< m1 >>
rect 23 354 24 355 
<< m1 >>
rect 24 354 25 355 
<< m2 >>
rect 24 354 25 355 
<< m1 >>
rect 25 354 26 355 
<< m1 >>
rect 26 354 27 355 
<< m2 >>
rect 26 354 27 355 
<< m2c >>
rect 26 354 27 355 
<< m1 >>
rect 26 354 27 355 
<< m2 >>
rect 26 354 27 355 
<< m2 >>
rect 27 354 28 355 
<< m1 >>
rect 28 354 29 355 
<< m2 >>
rect 28 354 29 355 
<< m1 >>
rect 29 354 30 355 
<< m2 >>
rect 29 354 30 355 
<< m1 >>
rect 30 354 31 355 
<< m2 >>
rect 30 354 31 355 
<< m1 >>
rect 31 354 32 355 
<< m2 >>
rect 31 354 32 355 
<< m1 >>
rect 32 354 33 355 
<< m2 >>
rect 32 354 33 355 
<< m1 >>
rect 33 354 34 355 
<< m2 >>
rect 33 354 34 355 
<< m1 >>
rect 34 354 35 355 
<< m2 >>
rect 34 354 35 355 
<< m1 >>
rect 35 354 36 355 
<< m2 >>
rect 35 354 36 355 
<< m1 >>
rect 36 354 37 355 
<< m2 >>
rect 36 354 37 355 
<< m1 >>
rect 37 354 38 355 
<< m2 >>
rect 37 354 38 355 
<< m1 >>
rect 38 354 39 355 
<< m2 >>
rect 38 354 39 355 
<< m1 >>
rect 39 354 40 355 
<< m2 >>
rect 39 354 40 355 
<< m1 >>
rect 40 354 41 355 
<< m2 >>
rect 40 354 41 355 
<< m1 >>
rect 41 354 42 355 
<< m2 >>
rect 41 354 42 355 
<< m1 >>
rect 42 354 43 355 
<< m2 >>
rect 42 354 43 355 
<< m1 >>
rect 43 354 44 355 
<< m2 >>
rect 43 354 44 355 
<< m1 >>
rect 44 354 45 355 
<< m2 >>
rect 44 354 45 355 
<< m1 >>
rect 45 354 46 355 
<< m2 >>
rect 45 354 46 355 
<< m1 >>
rect 46 354 47 355 
<< m2 >>
rect 46 354 47 355 
<< m1 >>
rect 47 354 48 355 
<< m2 >>
rect 47 354 48 355 
<< m1 >>
rect 48 354 49 355 
<< m2 >>
rect 48 354 49 355 
<< m1 >>
rect 49 354 50 355 
<< m2 >>
rect 49 354 50 355 
<< m1 >>
rect 50 354 51 355 
<< m2 >>
rect 50 354 51 355 
<< m1 >>
rect 51 354 52 355 
<< m2 >>
rect 51 354 52 355 
<< m1 >>
rect 52 354 53 355 
<< m2 >>
rect 52 354 53 355 
<< m1 >>
rect 53 354 54 355 
<< m2 >>
rect 53 354 54 355 
<< m1 >>
rect 54 354 55 355 
<< m2 >>
rect 54 354 55 355 
<< m1 >>
rect 55 354 56 355 
<< m2 >>
rect 55 354 56 355 
<< m1 >>
rect 56 354 57 355 
<< m2 >>
rect 56 354 57 355 
<< m1 >>
rect 57 354 58 355 
<< m2 >>
rect 57 354 58 355 
<< m1 >>
rect 58 354 59 355 
<< m2 >>
rect 58 354 59 355 
<< m1 >>
rect 59 354 60 355 
<< m2 >>
rect 59 354 60 355 
<< m1 >>
rect 60 354 61 355 
<< m2 >>
rect 60 354 61 355 
<< m1 >>
rect 61 354 62 355 
<< m2 >>
rect 61 354 62 355 
<< m1 >>
rect 62 354 63 355 
<< m2 >>
rect 62 354 63 355 
<< m1 >>
rect 63 354 64 355 
<< m2 >>
rect 63 354 64 355 
<< m1 >>
rect 64 354 65 355 
<< m2 >>
rect 64 354 65 355 
<< m1 >>
rect 65 354 66 355 
<< m2 >>
rect 65 354 66 355 
<< m1 >>
rect 66 354 67 355 
<< m2 >>
rect 66 354 67 355 
<< m1 >>
rect 67 354 68 355 
<< m2 >>
rect 67 354 68 355 
<< m1 >>
rect 68 354 69 355 
<< m2 >>
rect 68 354 69 355 
<< m1 >>
rect 69 354 70 355 
<< m2 >>
rect 69 354 70 355 
<< m1 >>
rect 70 354 71 355 
<< m2 >>
rect 70 354 71 355 
<< m1 >>
rect 71 354 72 355 
<< m2 >>
rect 71 354 72 355 
<< m1 >>
rect 72 354 73 355 
<< m2 >>
rect 72 354 73 355 
<< m1 >>
rect 73 354 74 355 
<< m2 >>
rect 73 354 74 355 
<< m1 >>
rect 74 354 75 355 
<< m2 >>
rect 74 354 75 355 
<< m1 >>
rect 75 354 76 355 
<< m2 >>
rect 75 354 76 355 
<< m1 >>
rect 76 354 77 355 
<< m2 >>
rect 76 354 77 355 
<< m1 >>
rect 77 354 78 355 
<< m2 >>
rect 77 354 78 355 
<< m1 >>
rect 78 354 79 355 
<< m2 >>
rect 78 354 79 355 
<< m1 >>
rect 79 354 80 355 
<< m2 >>
rect 79 354 80 355 
<< m1 >>
rect 80 354 81 355 
<< m2 >>
rect 80 354 81 355 
<< m1 >>
rect 81 354 82 355 
<< m2 >>
rect 81 354 82 355 
<< m1 >>
rect 82 354 83 355 
<< m2 >>
rect 82 354 83 355 
<< m1 >>
rect 83 354 84 355 
<< m2 >>
rect 83 354 84 355 
<< m1 >>
rect 84 354 85 355 
<< m2 >>
rect 84 354 85 355 
<< m1 >>
rect 85 354 86 355 
<< m2 >>
rect 85 354 86 355 
<< m1 >>
rect 86 354 87 355 
<< m2 >>
rect 86 354 87 355 
<< m1 >>
rect 87 354 88 355 
<< m2 >>
rect 87 354 88 355 
<< m1 >>
rect 88 354 89 355 
<< m2 >>
rect 88 354 89 355 
<< m1 >>
rect 89 354 90 355 
<< m2 >>
rect 89 354 90 355 
<< m1 >>
rect 90 354 91 355 
<< m2 >>
rect 90 354 91 355 
<< m1 >>
rect 91 354 92 355 
<< m2 >>
rect 91 354 92 355 
<< m1 >>
rect 92 354 93 355 
<< m2 >>
rect 92 354 93 355 
<< m1 >>
rect 93 354 94 355 
<< m2 >>
rect 93 354 94 355 
<< m1 >>
rect 94 354 95 355 
<< m2 >>
rect 94 354 95 355 
<< m1 >>
rect 95 354 96 355 
<< m2 >>
rect 95 354 96 355 
<< m1 >>
rect 96 354 97 355 
<< m2 >>
rect 96 354 97 355 
<< m1 >>
rect 97 354 98 355 
<< m2 >>
rect 97 354 98 355 
<< m1 >>
rect 98 354 99 355 
<< m2 >>
rect 98 354 99 355 
<< m1 >>
rect 99 354 100 355 
<< m2 >>
rect 99 354 100 355 
<< m1 >>
rect 100 354 101 355 
<< m2 >>
rect 100 354 101 355 
<< m1 >>
rect 101 354 102 355 
<< m2 >>
rect 101 354 102 355 
<< m1 >>
rect 102 354 103 355 
<< m2 >>
rect 102 354 103 355 
<< m1 >>
rect 103 354 104 355 
<< m2 >>
rect 103 354 104 355 
<< m1 >>
rect 104 354 105 355 
<< m2 >>
rect 104 354 105 355 
<< m1 >>
rect 105 354 106 355 
<< m2 >>
rect 105 354 106 355 
<< m1 >>
rect 106 354 107 355 
<< m2 >>
rect 106 354 107 355 
<< m1 >>
rect 107 354 108 355 
<< m2 >>
rect 107 354 108 355 
<< m1 >>
rect 108 354 109 355 
<< m2 >>
rect 108 354 109 355 
<< m1 >>
rect 109 354 110 355 
<< m2 >>
rect 109 354 110 355 
<< m1 >>
rect 110 354 111 355 
<< m2 >>
rect 110 354 111 355 
<< m1 >>
rect 111 354 112 355 
<< m2 >>
rect 111 354 112 355 
<< m1 >>
rect 112 354 113 355 
<< m2 >>
rect 112 354 113 355 
<< m1 >>
rect 113 354 114 355 
<< m2 >>
rect 113 354 114 355 
<< m1 >>
rect 114 354 115 355 
<< m2 >>
rect 114 354 115 355 
<< m1 >>
rect 115 354 116 355 
<< m2 >>
rect 115 354 116 355 
<< m1 >>
rect 116 354 117 355 
<< m2 >>
rect 116 354 117 355 
<< m1 >>
rect 117 354 118 355 
<< m2 >>
rect 117 354 118 355 
<< m1 >>
rect 118 354 119 355 
<< m2 >>
rect 118 354 119 355 
<< m1 >>
rect 119 354 120 355 
<< m2 >>
rect 119 354 120 355 
<< m1 >>
rect 120 354 121 355 
<< m2 >>
rect 120 354 121 355 
<< m1 >>
rect 121 354 122 355 
<< m2 >>
rect 121 354 122 355 
<< m1 >>
rect 122 354 123 355 
<< m2 >>
rect 122 354 123 355 
<< m1 >>
rect 123 354 124 355 
<< m2 >>
rect 123 354 124 355 
<< m1 >>
rect 124 354 125 355 
<< m2 >>
rect 124 354 125 355 
<< m1 >>
rect 125 354 126 355 
<< m2 >>
rect 125 354 126 355 
<< m1 >>
rect 126 354 127 355 
<< m2 >>
rect 126 354 127 355 
<< m1 >>
rect 127 354 128 355 
<< m2 >>
rect 127 354 128 355 
<< m1 >>
rect 128 354 129 355 
<< m2 >>
rect 128 354 129 355 
<< m1 >>
rect 129 354 130 355 
<< m2 >>
rect 129 354 130 355 
<< m1 >>
rect 130 354 131 355 
<< m2 >>
rect 130 354 131 355 
<< m1 >>
rect 131 354 132 355 
<< m2 >>
rect 131 354 132 355 
<< m1 >>
rect 132 354 133 355 
<< m2 >>
rect 132 354 133 355 
<< m1 >>
rect 133 354 134 355 
<< m2 >>
rect 133 354 134 355 
<< m1 >>
rect 134 354 135 355 
<< m2 >>
rect 134 354 135 355 
<< m1 >>
rect 135 354 136 355 
<< m2 >>
rect 135 354 136 355 
<< m1 >>
rect 136 354 137 355 
<< m2 >>
rect 136 354 137 355 
<< m1 >>
rect 137 354 138 355 
<< m2 >>
rect 137 354 138 355 
<< m1 >>
rect 138 354 139 355 
<< m2 >>
rect 138 354 139 355 
<< m1 >>
rect 139 354 140 355 
<< m2 >>
rect 139 354 140 355 
<< m1 >>
rect 140 354 141 355 
<< m2 >>
rect 140 354 141 355 
<< m1 >>
rect 141 354 142 355 
<< m2 >>
rect 141 354 142 355 
<< m1 >>
rect 142 354 143 355 
<< m2 >>
rect 142 354 143 355 
<< m1 >>
rect 143 354 144 355 
<< m2 >>
rect 143 354 144 355 
<< m1 >>
rect 144 354 145 355 
<< m2 >>
rect 144 354 145 355 
<< m1 >>
rect 145 354 146 355 
<< m2 >>
rect 145 354 146 355 
<< m1 >>
rect 146 354 147 355 
<< m2 >>
rect 146 354 147 355 
<< m1 >>
rect 147 354 148 355 
<< m2 >>
rect 147 354 148 355 
<< m1 >>
rect 148 354 149 355 
<< m2 >>
rect 148 354 149 355 
<< m1 >>
rect 149 354 150 355 
<< m2 >>
rect 149 354 150 355 
<< m1 >>
rect 150 354 151 355 
<< m2 >>
rect 150 354 151 355 
<< m1 >>
rect 151 354 152 355 
<< m2 >>
rect 151 354 152 355 
<< m1 >>
rect 152 354 153 355 
<< m2 >>
rect 152 354 153 355 
<< m1 >>
rect 153 354 154 355 
<< m2 >>
rect 153 354 154 355 
<< m1 >>
rect 154 354 155 355 
<< m2 >>
rect 154 354 155 355 
<< m1 >>
rect 155 354 156 355 
<< m2 >>
rect 155 354 156 355 
<< m1 >>
rect 156 354 157 355 
<< m2 >>
rect 156 354 157 355 
<< m1 >>
rect 157 354 158 355 
<< m2 >>
rect 157 354 158 355 
<< m1 >>
rect 158 354 159 355 
<< m2 >>
rect 158 354 159 355 
<< m1 >>
rect 159 354 160 355 
<< m2 >>
rect 159 354 160 355 
<< m1 >>
rect 160 354 161 355 
<< m2 >>
rect 160 354 161 355 
<< m1 >>
rect 161 354 162 355 
<< m2 >>
rect 161 354 162 355 
<< m1 >>
rect 162 354 163 355 
<< m2 >>
rect 162 354 163 355 
<< m1 >>
rect 163 354 164 355 
<< m2 >>
rect 163 354 164 355 
<< m1 >>
rect 164 354 165 355 
<< m2 >>
rect 164 354 165 355 
<< m1 >>
rect 165 354 166 355 
<< m2 >>
rect 165 354 166 355 
<< m1 >>
rect 166 354 167 355 
<< m2 >>
rect 166 354 167 355 
<< m1 >>
rect 167 354 168 355 
<< m2 >>
rect 167 354 168 355 
<< m1 >>
rect 168 354 169 355 
<< m2 >>
rect 168 354 169 355 
<< m1 >>
rect 169 354 170 355 
<< m2 >>
rect 169 354 170 355 
<< m1 >>
rect 170 354 171 355 
<< m2 >>
rect 170 354 171 355 
<< m1 >>
rect 171 354 172 355 
<< m2 >>
rect 171 354 172 355 
<< m1 >>
rect 172 354 173 355 
<< m2 >>
rect 172 354 173 355 
<< m1 >>
rect 173 354 174 355 
<< m2 >>
rect 173 354 174 355 
<< m1 >>
rect 174 354 175 355 
<< m2 >>
rect 174 354 175 355 
<< m1 >>
rect 175 354 176 355 
<< m2 >>
rect 175 354 176 355 
<< m1 >>
rect 176 354 177 355 
<< m2 >>
rect 176 354 177 355 
<< m1 >>
rect 177 354 178 355 
<< m2 >>
rect 177 354 178 355 
<< m1 >>
rect 178 354 179 355 
<< m2 >>
rect 178 354 179 355 
<< m1 >>
rect 179 354 180 355 
<< m2 >>
rect 179 354 180 355 
<< m1 >>
rect 180 354 181 355 
<< m2 >>
rect 180 354 181 355 
<< m1 >>
rect 181 354 182 355 
<< m2 >>
rect 181 354 182 355 
<< m1 >>
rect 182 354 183 355 
<< m2 >>
rect 182 354 183 355 
<< m1 >>
rect 183 354 184 355 
<< m2 >>
rect 183 354 184 355 
<< m1 >>
rect 184 354 185 355 
<< m2 >>
rect 184 354 185 355 
<< m1 >>
rect 185 354 186 355 
<< m2 >>
rect 185 354 186 355 
<< m1 >>
rect 186 354 187 355 
<< m2 >>
rect 186 354 187 355 
<< m1 >>
rect 187 354 188 355 
<< m2 >>
rect 187 354 188 355 
<< m1 >>
rect 188 354 189 355 
<< m2 >>
rect 188 354 189 355 
<< m1 >>
rect 189 354 190 355 
<< m2 >>
rect 189 354 190 355 
<< m1 >>
rect 190 354 191 355 
<< m2 >>
rect 190 354 191 355 
<< m1 >>
rect 191 354 192 355 
<< m2 >>
rect 191 354 192 355 
<< m1 >>
rect 192 354 193 355 
<< m2 >>
rect 192 354 193 355 
<< m1 >>
rect 193 354 194 355 
<< m2 >>
rect 193 354 194 355 
<< m1 >>
rect 194 354 195 355 
<< m2 >>
rect 194 354 195 355 
<< m1 >>
rect 195 354 196 355 
<< m2 >>
rect 195 354 196 355 
<< m1 >>
rect 196 354 197 355 
<< m2 >>
rect 196 354 197 355 
<< m1 >>
rect 197 354 198 355 
<< m2 >>
rect 197 354 198 355 
<< m1 >>
rect 198 354 199 355 
<< m2 >>
rect 198 354 199 355 
<< m1 >>
rect 199 354 200 355 
<< m2 >>
rect 199 354 200 355 
<< m1 >>
rect 200 354 201 355 
<< m2 >>
rect 200 354 201 355 
<< m1 >>
rect 201 354 202 355 
<< m2 >>
rect 201 354 202 355 
<< m1 >>
rect 202 354 203 355 
<< m2 >>
rect 202 354 203 355 
<< m1 >>
rect 203 354 204 355 
<< m2 >>
rect 203 354 204 355 
<< m1 >>
rect 204 354 205 355 
<< m2 >>
rect 204 354 205 355 
<< m1 >>
rect 205 354 206 355 
<< m2 >>
rect 205 354 206 355 
<< m1 >>
rect 206 354 207 355 
<< m2 >>
rect 206 354 207 355 
<< m1 >>
rect 207 354 208 355 
<< m2 >>
rect 207 354 208 355 
<< m1 >>
rect 208 354 209 355 
<< m2 >>
rect 208 354 209 355 
<< m1 >>
rect 209 354 210 355 
<< m2 >>
rect 209 354 210 355 
<< m1 >>
rect 210 354 211 355 
<< m2 >>
rect 210 354 211 355 
<< m1 >>
rect 211 354 212 355 
<< m2 >>
rect 211 354 212 355 
<< m1 >>
rect 212 354 213 355 
<< m2 >>
rect 212 354 213 355 
<< m1 >>
rect 213 354 214 355 
<< m2 >>
rect 213 354 214 355 
<< m1 >>
rect 214 354 215 355 
<< m2 >>
rect 214 354 215 355 
<< m1 >>
rect 215 354 216 355 
<< m2 >>
rect 215 354 216 355 
<< m1 >>
rect 216 354 217 355 
<< m2 >>
rect 216 354 217 355 
<< m1 >>
rect 217 354 218 355 
<< m2 >>
rect 217 354 218 355 
<< m1 >>
rect 218 354 219 355 
<< m2 >>
rect 218 354 219 355 
<< m1 >>
rect 219 354 220 355 
<< m2 >>
rect 219 354 220 355 
<< m1 >>
rect 220 354 221 355 
<< m2 >>
rect 220 354 221 355 
<< m1 >>
rect 221 354 222 355 
<< m2 >>
rect 221 354 222 355 
<< m1 >>
rect 222 354 223 355 
<< m2 >>
rect 222 354 223 355 
<< m1 >>
rect 223 354 224 355 
<< m2 >>
rect 223 354 224 355 
<< m1 >>
rect 224 354 225 355 
<< m2 >>
rect 224 354 225 355 
<< m1 >>
rect 225 354 226 355 
<< m2 >>
rect 225 354 226 355 
<< m1 >>
rect 226 354 227 355 
<< m2 >>
rect 226 354 227 355 
<< m1 >>
rect 227 354 228 355 
<< m2 >>
rect 227 354 228 355 
<< m1 >>
rect 228 354 229 355 
<< m2 >>
rect 228 354 229 355 
<< m1 >>
rect 229 354 230 355 
<< m2 >>
rect 229 354 230 355 
<< m1 >>
rect 230 354 231 355 
<< m2 >>
rect 230 354 231 355 
<< m1 >>
rect 231 354 232 355 
<< m2 >>
rect 231 354 232 355 
<< m1 >>
rect 232 354 233 355 
<< m2 >>
rect 232 354 233 355 
<< m1 >>
rect 233 354 234 355 
<< m2 >>
rect 233 354 234 355 
<< m1 >>
rect 234 354 235 355 
<< m2 >>
rect 234 354 235 355 
<< m1 >>
rect 235 354 236 355 
<< m2 >>
rect 235 354 236 355 
<< m1 >>
rect 236 354 237 355 
<< m2 >>
rect 236 354 237 355 
<< m1 >>
rect 237 354 238 355 
<< m2 >>
rect 237 354 238 355 
<< m1 >>
rect 238 354 239 355 
<< m2 >>
rect 238 354 239 355 
<< m1 >>
rect 239 354 240 355 
<< m2 >>
rect 239 354 240 355 
<< m1 >>
rect 240 354 241 355 
<< m2 >>
rect 240 354 241 355 
<< m1 >>
rect 241 354 242 355 
<< m2 >>
rect 241 354 242 355 
<< m1 >>
rect 242 354 243 355 
<< m2 >>
rect 242 354 243 355 
<< m1 >>
rect 243 354 244 355 
<< m2 >>
rect 243 354 244 355 
<< m1 >>
rect 244 354 245 355 
<< m2 >>
rect 244 354 245 355 
<< m1 >>
rect 245 354 246 355 
<< m2 >>
rect 245 354 246 355 
<< m1 >>
rect 246 354 247 355 
<< m2 >>
rect 246 354 247 355 
<< m1 >>
rect 247 354 248 355 
<< m2 >>
rect 247 354 248 355 
<< m1 >>
rect 248 354 249 355 
<< m2 >>
rect 248 354 249 355 
<< m1 >>
rect 249 354 250 355 
<< m2 >>
rect 249 354 250 355 
<< m1 >>
rect 250 354 251 355 
<< m2 >>
rect 250 354 251 355 
<< m1 >>
rect 251 354 252 355 
<< m2 >>
rect 251 354 252 355 
<< m1 >>
rect 252 354 253 355 
<< m2 >>
rect 252 354 253 355 
<< m1 >>
rect 253 354 254 355 
<< m2 >>
rect 253 354 254 355 
<< m1 >>
rect 254 354 255 355 
<< m2 >>
rect 254 354 255 355 
<< m1 >>
rect 255 354 256 355 
<< m2 >>
rect 255 354 256 355 
<< m1 >>
rect 256 354 257 355 
<< m2 >>
rect 256 354 257 355 
<< m1 >>
rect 257 354 258 355 
<< m2 >>
rect 257 354 258 355 
<< m1 >>
rect 258 354 259 355 
<< m2 >>
rect 258 354 259 355 
<< m1 >>
rect 259 354 260 355 
<< m2 >>
rect 259 354 260 355 
<< m1 >>
rect 260 354 261 355 
<< m2 >>
rect 260 354 261 355 
<< m1 >>
rect 261 354 262 355 
<< m2 >>
rect 261 354 262 355 
<< m1 >>
rect 262 354 263 355 
<< m2 >>
rect 262 354 263 355 
<< m1 >>
rect 263 354 264 355 
<< m2 >>
rect 263 354 264 355 
<< m1 >>
rect 264 354 265 355 
<< m2 >>
rect 264 354 265 355 
<< m1 >>
rect 265 354 266 355 
<< m2 >>
rect 265 354 266 355 
<< m1 >>
rect 266 354 267 355 
<< m2 >>
rect 266 354 267 355 
<< m1 >>
rect 267 354 268 355 
<< m2 >>
rect 267 354 268 355 
<< m1 >>
rect 268 354 269 355 
<< m2 >>
rect 268 354 269 355 
<< m1 >>
rect 269 354 270 355 
<< m2 >>
rect 269 354 270 355 
<< m1 >>
rect 270 354 271 355 
<< m2 >>
rect 270 354 271 355 
<< m1 >>
rect 271 354 272 355 
<< m2 >>
rect 271 354 272 355 
<< m1 >>
rect 272 354 273 355 
<< m2 >>
rect 272 354 273 355 
<< m1 >>
rect 273 354 274 355 
<< m2 >>
rect 273 354 274 355 
<< m1 >>
rect 274 354 275 355 
<< m2 >>
rect 274 354 275 355 
<< m1 >>
rect 275 354 276 355 
<< m2 >>
rect 275 354 276 355 
<< m1 >>
rect 276 354 277 355 
<< m2 >>
rect 276 354 277 355 
<< m1 >>
rect 277 354 278 355 
<< m2 >>
rect 277 354 278 355 
<< m1 >>
rect 278 354 279 355 
<< m2 >>
rect 278 354 279 355 
<< m1 >>
rect 279 354 280 355 
<< m2 >>
rect 279 354 280 355 
<< m1 >>
rect 280 354 281 355 
<< m2 >>
rect 280 354 281 355 
<< m1 >>
rect 281 354 282 355 
<< m2 >>
rect 281 354 282 355 
<< m1 >>
rect 282 354 283 355 
<< m2 >>
rect 282 354 283 355 
<< m1 >>
rect 283 354 284 355 
<< m2 >>
rect 283 354 284 355 
<< m1 >>
rect 284 354 285 355 
<< m2 >>
rect 284 354 285 355 
<< m1 >>
rect 285 354 286 355 
<< m2 >>
rect 285 354 286 355 
<< m1 >>
rect 286 354 287 355 
<< m2 >>
rect 286 354 287 355 
<< m1 >>
rect 287 354 288 355 
<< m2 >>
rect 287 354 288 355 
<< m1 >>
rect 288 354 289 355 
<< m2 >>
rect 288 354 289 355 
<< m1 >>
rect 289 354 290 355 
<< m2 >>
rect 289 354 290 355 
<< m1 >>
rect 290 354 291 355 
<< m2 >>
rect 290 354 291 355 
<< m1 >>
rect 291 354 292 355 
<< m2 >>
rect 291 354 292 355 
<< m1 >>
rect 292 354 293 355 
<< m2 >>
rect 292 354 293 355 
<< m1 >>
rect 293 354 294 355 
<< m2 >>
rect 293 354 294 355 
<< m1 >>
rect 294 354 295 355 
<< m2 >>
rect 294 354 295 355 
<< m1 >>
rect 295 354 296 355 
<< m2 >>
rect 295 354 296 355 
<< m1 >>
rect 296 354 297 355 
<< m2 >>
rect 296 354 297 355 
<< m1 >>
rect 297 354 298 355 
<< m2 >>
rect 297 354 298 355 
<< m1 >>
rect 298 354 299 355 
<< m2 >>
rect 298 354 299 355 
<< m1 >>
rect 299 354 300 355 
<< m2 >>
rect 299 354 300 355 
<< m1 >>
rect 300 354 301 355 
<< m2 >>
rect 300 354 301 355 
<< m1 >>
rect 301 354 302 355 
<< m2 >>
rect 301 354 302 355 
<< m1 >>
rect 302 354 303 355 
<< m2 >>
rect 302 354 303 355 
<< m1 >>
rect 303 354 304 355 
<< m2 >>
rect 303 354 304 355 
<< m1 >>
rect 304 354 305 355 
<< m2 >>
rect 304 354 305 355 
<< m1 >>
rect 305 354 306 355 
<< m2 >>
rect 305 354 306 355 
<< m1 >>
rect 306 354 307 355 
<< m2 >>
rect 306 354 307 355 
<< m1 >>
rect 307 354 308 355 
<< m2 >>
rect 307 354 308 355 
<< m1 >>
rect 308 354 309 355 
<< m2 >>
rect 308 354 309 355 
<< m1 >>
rect 309 354 310 355 
<< m2 >>
rect 309 354 310 355 
<< m1 >>
rect 310 354 311 355 
<< m2 >>
rect 310 354 311 355 
<< m1 >>
rect 311 354 312 355 
<< m2 >>
rect 311 354 312 355 
<< m1 >>
rect 312 354 313 355 
<< m2 >>
rect 312 354 313 355 
<< m1 >>
rect 313 354 314 355 
<< m2 >>
rect 313 354 314 355 
<< m1 >>
rect 314 354 315 355 
<< m2 >>
rect 314 354 315 355 
<< m1 >>
rect 315 354 316 355 
<< m2 >>
rect 315 354 316 355 
<< m1 >>
rect 316 354 317 355 
<< m2 >>
rect 316 354 317 355 
<< m1 >>
rect 317 354 318 355 
<< m2 >>
rect 317 354 318 355 
<< m1 >>
rect 318 354 319 355 
<< m2 >>
rect 318 354 319 355 
<< m1 >>
rect 319 354 320 355 
<< m2 >>
rect 319 354 320 355 
<< m1 >>
rect 320 354 321 355 
<< m2 >>
rect 320 354 321 355 
<< m1 >>
rect 321 354 322 355 
<< m2 >>
rect 321 354 322 355 
<< m1 >>
rect 322 354 323 355 
<< m2 >>
rect 322 354 323 355 
<< m1 >>
rect 323 354 324 355 
<< m2 >>
rect 323 354 324 355 
<< m1 >>
rect 324 354 325 355 
<< m2 >>
rect 324 354 325 355 
<< m1 >>
rect 325 354 326 355 
<< m2 >>
rect 325 354 326 355 
<< m1 >>
rect 326 354 327 355 
<< m2 >>
rect 326 354 327 355 
<< m1 >>
rect 327 354 328 355 
<< m2 >>
rect 327 354 328 355 
<< m1 >>
rect 328 354 329 355 
<< m2 >>
rect 328 354 329 355 
<< m1 >>
rect 329 354 330 355 
<< m2 >>
rect 329 354 330 355 
<< m1 >>
rect 330 354 331 355 
<< m2 >>
rect 330 354 331 355 
<< m1 >>
rect 331 354 332 355 
<< m2 >>
rect 331 354 332 355 
<< m1 >>
rect 332 354 333 355 
<< m2 >>
rect 332 354 333 355 
<< m1 >>
rect 333 354 334 355 
<< m2 >>
rect 333 354 334 355 
<< m1 >>
rect 334 354 335 355 
<< m2 >>
rect 334 354 335 355 
<< m1 >>
rect 335 354 336 355 
<< m1 >>
rect 336 354 337 355 
<< m1 >>
rect 337 354 338 355 
<< m1 >>
rect 338 354 339 355 
<< m1 >>
rect 339 354 340 355 
<< m1 >>
rect 340 354 341 355 
<< m1 >>
rect 343 354 344 355 
<< m2 >>
rect 24 355 25 356 
<< m1 >>
rect 343 355 344 356 
<< m1 >>
rect 24 356 25 357 
<< m2 >>
rect 24 356 25 357 
<< m2c >>
rect 24 356 25 357 
<< m1 >>
rect 24 356 25 357 
<< m2 >>
rect 24 356 25 357 
<< m1 >>
rect 25 356 26 357 
<< m1 >>
rect 26 356 27 357 
<< m1 >>
rect 27 356 28 357 
<< m1 >>
rect 28 356 29 357 
<< m1 >>
rect 29 356 30 357 
<< m1 >>
rect 30 356 31 357 
<< m1 >>
rect 31 356 32 357 
<< m1 >>
rect 32 356 33 357 
<< m1 >>
rect 33 356 34 357 
<< m1 >>
rect 34 356 35 357 
<< m1 >>
rect 35 356 36 357 
<< m1 >>
rect 36 356 37 357 
<< m1 >>
rect 37 356 38 357 
<< m1 >>
rect 38 356 39 357 
<< m1 >>
rect 39 356 40 357 
<< m1 >>
rect 40 356 41 357 
<< m1 >>
rect 41 356 42 357 
<< m1 >>
rect 42 356 43 357 
<< m1 >>
rect 43 356 44 357 
<< m1 >>
rect 44 356 45 357 
<< m1 >>
rect 45 356 46 357 
<< m1 >>
rect 46 356 47 357 
<< m1 >>
rect 47 356 48 357 
<< m1 >>
rect 48 356 49 357 
<< m1 >>
rect 49 356 50 357 
<< m1 >>
rect 50 356 51 357 
<< m1 >>
rect 51 356 52 357 
<< m1 >>
rect 52 356 53 357 
<< m1 >>
rect 53 356 54 357 
<< m1 >>
rect 54 356 55 357 
<< m1 >>
rect 55 356 56 357 
<< m1 >>
rect 56 356 57 357 
<< m1 >>
rect 57 356 58 357 
<< m1 >>
rect 58 356 59 357 
<< m1 >>
rect 59 356 60 357 
<< m1 >>
rect 60 356 61 357 
<< m1 >>
rect 61 356 62 357 
<< m1 >>
rect 62 356 63 357 
<< m1 >>
rect 63 356 64 357 
<< m1 >>
rect 64 356 65 357 
<< m1 >>
rect 65 356 66 357 
<< m1 >>
rect 66 356 67 357 
<< m1 >>
rect 67 356 68 357 
<< m1 >>
rect 68 356 69 357 
<< m1 >>
rect 69 356 70 357 
<< m1 >>
rect 70 356 71 357 
<< m1 >>
rect 71 356 72 357 
<< m1 >>
rect 72 356 73 357 
<< m1 >>
rect 73 356 74 357 
<< m1 >>
rect 74 356 75 357 
<< m1 >>
rect 75 356 76 357 
<< m1 >>
rect 76 356 77 357 
<< m1 >>
rect 77 356 78 357 
<< m1 >>
rect 78 356 79 357 
<< m1 >>
rect 79 356 80 357 
<< m1 >>
rect 80 356 81 357 
<< m1 >>
rect 81 356 82 357 
<< m1 >>
rect 82 356 83 357 
<< m1 >>
rect 83 356 84 357 
<< m1 >>
rect 84 356 85 357 
<< m1 >>
rect 85 356 86 357 
<< m1 >>
rect 86 356 87 357 
<< m1 >>
rect 87 356 88 357 
<< m1 >>
rect 88 356 89 357 
<< m1 >>
rect 89 356 90 357 
<< m1 >>
rect 90 356 91 357 
<< m1 >>
rect 91 356 92 357 
<< m1 >>
rect 92 356 93 357 
<< m1 >>
rect 93 356 94 357 
<< m1 >>
rect 94 356 95 357 
<< m1 >>
rect 95 356 96 357 
<< m1 >>
rect 96 356 97 357 
<< m1 >>
rect 97 356 98 357 
<< m1 >>
rect 98 356 99 357 
<< m1 >>
rect 99 356 100 357 
<< m1 >>
rect 100 356 101 357 
<< m1 >>
rect 101 356 102 357 
<< m1 >>
rect 102 356 103 357 
<< m1 >>
rect 103 356 104 357 
<< m1 >>
rect 104 356 105 357 
<< m1 >>
rect 105 356 106 357 
<< m1 >>
rect 106 356 107 357 
<< m1 >>
rect 107 356 108 357 
<< m1 >>
rect 108 356 109 357 
<< m1 >>
rect 109 356 110 357 
<< m1 >>
rect 110 356 111 357 
<< m1 >>
rect 111 356 112 357 
<< m1 >>
rect 112 356 113 357 
<< m1 >>
rect 113 356 114 357 
<< m1 >>
rect 114 356 115 357 
<< m1 >>
rect 115 356 116 357 
<< m1 >>
rect 116 356 117 357 
<< m1 >>
rect 117 356 118 357 
<< m1 >>
rect 118 356 119 357 
<< m1 >>
rect 119 356 120 357 
<< m1 >>
rect 120 356 121 357 
<< m1 >>
rect 121 356 122 357 
<< m1 >>
rect 122 356 123 357 
<< m1 >>
rect 123 356 124 357 
<< m1 >>
rect 124 356 125 357 
<< m1 >>
rect 125 356 126 357 
<< m1 >>
rect 126 356 127 357 
<< m1 >>
rect 127 356 128 357 
<< m1 >>
rect 128 356 129 357 
<< m1 >>
rect 129 356 130 357 
<< m1 >>
rect 130 356 131 357 
<< m1 >>
rect 131 356 132 357 
<< m1 >>
rect 132 356 133 357 
<< m1 >>
rect 133 356 134 357 
<< m1 >>
rect 134 356 135 357 
<< m1 >>
rect 135 356 136 357 
<< m1 >>
rect 136 356 137 357 
<< m1 >>
rect 137 356 138 357 
<< m1 >>
rect 138 356 139 357 
<< m1 >>
rect 139 356 140 357 
<< m1 >>
rect 140 356 141 357 
<< m1 >>
rect 141 356 142 357 
<< m1 >>
rect 142 356 143 357 
<< m1 >>
rect 143 356 144 357 
<< m1 >>
rect 144 356 145 357 
<< m1 >>
rect 145 356 146 357 
<< m1 >>
rect 146 356 147 357 
<< m1 >>
rect 147 356 148 357 
<< m1 >>
rect 148 356 149 357 
<< m1 >>
rect 149 356 150 357 
<< m1 >>
rect 150 356 151 357 
<< m1 >>
rect 151 356 152 357 
<< m1 >>
rect 152 356 153 357 
<< m1 >>
rect 153 356 154 357 
<< m1 >>
rect 154 356 155 357 
<< m1 >>
rect 155 356 156 357 
<< m1 >>
rect 156 356 157 357 
<< m1 >>
rect 157 356 158 357 
<< m1 >>
rect 158 356 159 357 
<< m1 >>
rect 159 356 160 357 
<< m1 >>
rect 160 356 161 357 
<< m1 >>
rect 161 356 162 357 
<< m1 >>
rect 162 356 163 357 
<< m1 >>
rect 163 356 164 357 
<< m1 >>
rect 164 356 165 357 
<< m1 >>
rect 165 356 166 357 
<< m1 >>
rect 166 356 167 357 
<< m1 >>
rect 167 356 168 357 
<< m1 >>
rect 168 356 169 357 
<< m1 >>
rect 169 356 170 357 
<< m1 >>
rect 170 356 171 357 
<< m1 >>
rect 171 356 172 357 
<< m1 >>
rect 172 356 173 357 
<< m1 >>
rect 173 356 174 357 
<< m1 >>
rect 174 356 175 357 
<< m1 >>
rect 175 356 176 357 
<< m1 >>
rect 176 356 177 357 
<< m1 >>
rect 177 356 178 357 
<< m1 >>
rect 178 356 179 357 
<< m1 >>
rect 179 356 180 357 
<< m1 >>
rect 180 356 181 357 
<< m1 >>
rect 181 356 182 357 
<< m1 >>
rect 182 356 183 357 
<< m1 >>
rect 183 356 184 357 
<< m1 >>
rect 184 356 185 357 
<< m1 >>
rect 185 356 186 357 
<< m1 >>
rect 186 356 187 357 
<< m1 >>
rect 187 356 188 357 
<< m1 >>
rect 188 356 189 357 
<< m1 >>
rect 189 356 190 357 
<< m1 >>
rect 190 356 191 357 
<< m1 >>
rect 191 356 192 357 
<< m1 >>
rect 192 356 193 357 
<< m1 >>
rect 193 356 194 357 
<< m1 >>
rect 194 356 195 357 
<< m1 >>
rect 195 356 196 357 
<< m1 >>
rect 196 356 197 357 
<< m1 >>
rect 197 356 198 357 
<< m1 >>
rect 198 356 199 357 
<< m1 >>
rect 199 356 200 357 
<< m1 >>
rect 200 356 201 357 
<< m1 >>
rect 201 356 202 357 
<< m1 >>
rect 202 356 203 357 
<< m1 >>
rect 203 356 204 357 
<< m1 >>
rect 204 356 205 357 
<< m1 >>
rect 205 356 206 357 
<< m1 >>
rect 206 356 207 357 
<< m1 >>
rect 207 356 208 357 
<< m1 >>
rect 208 356 209 357 
<< m1 >>
rect 209 356 210 357 
<< m1 >>
rect 210 356 211 357 
<< m1 >>
rect 211 356 212 357 
<< m1 >>
rect 212 356 213 357 
<< m1 >>
rect 213 356 214 357 
<< m1 >>
rect 214 356 215 357 
<< m1 >>
rect 215 356 216 357 
<< m1 >>
rect 216 356 217 357 
<< m1 >>
rect 217 356 218 357 
<< m1 >>
rect 218 356 219 357 
<< m1 >>
rect 219 356 220 357 
<< m1 >>
rect 220 356 221 357 
<< m1 >>
rect 221 356 222 357 
<< m1 >>
rect 222 356 223 357 
<< m1 >>
rect 223 356 224 357 
<< m1 >>
rect 224 356 225 357 
<< m1 >>
rect 225 356 226 357 
<< m1 >>
rect 226 356 227 357 
<< m1 >>
rect 227 356 228 357 
<< m1 >>
rect 228 356 229 357 
<< m1 >>
rect 229 356 230 357 
<< m1 >>
rect 230 356 231 357 
<< m1 >>
rect 231 356 232 357 
<< m1 >>
rect 232 356 233 357 
<< m1 >>
rect 233 356 234 357 
<< m1 >>
rect 234 356 235 357 
<< m1 >>
rect 235 356 236 357 
<< m1 >>
rect 236 356 237 357 
<< m1 >>
rect 237 356 238 357 
<< m1 >>
rect 238 356 239 357 
<< m1 >>
rect 239 356 240 357 
<< m1 >>
rect 240 356 241 357 
<< m1 >>
rect 241 356 242 357 
<< m1 >>
rect 242 356 243 357 
<< m1 >>
rect 243 356 244 357 
<< m1 >>
rect 244 356 245 357 
<< m1 >>
rect 245 356 246 357 
<< m1 >>
rect 246 356 247 357 
<< m1 >>
rect 247 356 248 357 
<< m1 >>
rect 248 356 249 357 
<< m1 >>
rect 249 356 250 357 
<< m1 >>
rect 250 356 251 357 
<< m1 >>
rect 251 356 252 357 
<< m1 >>
rect 252 356 253 357 
<< m1 >>
rect 253 356 254 357 
<< m1 >>
rect 254 356 255 357 
<< m1 >>
rect 255 356 256 357 
<< m1 >>
rect 256 356 257 357 
<< m1 >>
rect 257 356 258 357 
<< m1 >>
rect 258 356 259 357 
<< m1 >>
rect 259 356 260 357 
<< m1 >>
rect 260 356 261 357 
<< m1 >>
rect 261 356 262 357 
<< m1 >>
rect 262 356 263 357 
<< m1 >>
rect 263 356 264 357 
<< m1 >>
rect 264 356 265 357 
<< m1 >>
rect 265 356 266 357 
<< m1 >>
rect 266 356 267 357 
<< m1 >>
rect 267 356 268 357 
<< m1 >>
rect 268 356 269 357 
<< m1 >>
rect 269 356 270 357 
<< m1 >>
rect 270 356 271 357 
<< m1 >>
rect 271 356 272 357 
<< m1 >>
rect 272 356 273 357 
<< m1 >>
rect 273 356 274 357 
<< m1 >>
rect 274 356 275 357 
<< m1 >>
rect 275 356 276 357 
<< m1 >>
rect 276 356 277 357 
<< m1 >>
rect 277 356 278 357 
<< m1 >>
rect 278 356 279 357 
<< m1 >>
rect 279 356 280 357 
<< m1 >>
rect 280 356 281 357 
<< m1 >>
rect 281 356 282 357 
<< m1 >>
rect 282 356 283 357 
<< m1 >>
rect 283 356 284 357 
<< m1 >>
rect 284 356 285 357 
<< m1 >>
rect 285 356 286 357 
<< m1 >>
rect 286 356 287 357 
<< m1 >>
rect 287 356 288 357 
<< m1 >>
rect 288 356 289 357 
<< m1 >>
rect 289 356 290 357 
<< m1 >>
rect 290 356 291 357 
<< m1 >>
rect 291 356 292 357 
<< m1 >>
rect 292 356 293 357 
<< m1 >>
rect 293 356 294 357 
<< m1 >>
rect 294 356 295 357 
<< m1 >>
rect 295 356 296 357 
<< m1 >>
rect 296 356 297 357 
<< m1 >>
rect 297 356 298 357 
<< m1 >>
rect 298 356 299 357 
<< m1 >>
rect 299 356 300 357 
<< m1 >>
rect 300 356 301 357 
<< m1 >>
rect 301 356 302 357 
<< m1 >>
rect 302 356 303 357 
<< m1 >>
rect 303 356 304 357 
<< m1 >>
rect 304 356 305 357 
<< m1 >>
rect 305 356 306 357 
<< m1 >>
rect 306 356 307 357 
<< m1 >>
rect 307 356 308 357 
<< m1 >>
rect 308 356 309 357 
<< m1 >>
rect 309 356 310 357 
<< m1 >>
rect 310 356 311 357 
<< m1 >>
rect 311 356 312 357 
<< m1 >>
rect 312 356 313 357 
<< m1 >>
rect 313 356 314 357 
<< m1 >>
rect 314 356 315 357 
<< m1 >>
rect 315 356 316 357 
<< m1 >>
rect 316 356 317 357 
<< m1 >>
rect 317 356 318 357 
<< m1 >>
rect 318 356 319 357 
<< m1 >>
rect 319 356 320 357 
<< m1 >>
rect 320 356 321 357 
<< m1 >>
rect 321 356 322 357 
<< m1 >>
rect 322 356 323 357 
<< m1 >>
rect 323 356 324 357 
<< m1 >>
rect 324 356 325 357 
<< m1 >>
rect 325 356 326 357 
<< m1 >>
rect 326 356 327 357 
<< m1 >>
rect 327 356 328 357 
<< m1 >>
rect 328 356 329 357 
<< m1 >>
rect 329 356 330 357 
<< m1 >>
rect 330 356 331 357 
<< m1 >>
rect 331 356 332 357 
<< m1 >>
rect 332 356 333 357 
<< m1 >>
rect 333 356 334 357 
<< m1 >>
rect 334 356 335 357 
<< m1 >>
rect 335 356 336 357 
<< m1 >>
rect 336 356 337 357 
<< m1 >>
rect 337 356 338 357 
<< m1 >>
rect 338 356 339 357 
<< m1 >>
rect 339 356 340 357 
<< m1 >>
rect 340 356 341 357 
<< m1 >>
rect 341 356 342 357 
<< m1 >>
rect 342 356 343 357 
<< m1 >>
rect 343 356 344 357 
<< labels >>
rlabel pdiffusion 283 174 284 175  0 t = 1
rlabel pdiffusion 286 174 287 175  0 t = 2
rlabel pdiffusion 283 179 284 180  0 t = 3
rlabel pdiffusion 286 179 287 180  0 t = 4
rlabel pdiffusion 282 174 288 180 0 cell no = 1
<< m1 >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< m2 >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< m2c >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< labels >>
rlabel pdiffusion 157 210 158 211  0 t = 1
rlabel pdiffusion 160 210 161 211  0 t = 2
rlabel pdiffusion 157 215 158 216  0 t = 3
rlabel pdiffusion 160 215 161 216  0 t = 4
rlabel pdiffusion 156 210 162 216 0 cell no = 2
<< m1 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2c >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< labels >>
rlabel pdiffusion 265 174 266 175  0 t = 1
rlabel pdiffusion 268 174 269 175  0 t = 2
rlabel pdiffusion 265 179 266 180  0 t = 3
rlabel pdiffusion 268 179 269 180  0 t = 4
rlabel pdiffusion 264 174 270 180 0 cell no = 3
<< m1 >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< m2 >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< m2c >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< labels >>
rlabel pdiffusion 175 48 176 49  0 t = 1
rlabel pdiffusion 178 48 179 49  0 t = 2
rlabel pdiffusion 175 53 176 54  0 t = 3
rlabel pdiffusion 178 53 179 54  0 t = 4
rlabel pdiffusion 174 48 180 54 0 cell no = 4
<< m1 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2c >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< labels >>
rlabel pdiffusion 283 318 284 319  0 t = 1
rlabel pdiffusion 286 318 287 319  0 t = 2
rlabel pdiffusion 283 323 284 324  0 t = 3
rlabel pdiffusion 286 323 287 324  0 t = 4
rlabel pdiffusion 282 318 288 324 0 cell no = 5
<< m1 >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< m2 >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< m2c >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< labels >>
rlabel pdiffusion 301 210 302 211  0 t = 1
rlabel pdiffusion 304 210 305 211  0 t = 2
rlabel pdiffusion 301 215 302 216  0 t = 3
rlabel pdiffusion 304 215 305 216  0 t = 4
rlabel pdiffusion 300 210 306 216 0 cell no = 6
<< m1 >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< m2 >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< m2c >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< labels >>
rlabel pdiffusion 301 228 302 229  0 t = 1
rlabel pdiffusion 304 228 305 229  0 t = 2
rlabel pdiffusion 301 233 302 234  0 t = 3
rlabel pdiffusion 304 233 305 234  0 t = 4
rlabel pdiffusion 300 228 306 234 0 cell no = 7
<< m1 >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< m2 >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< m2c >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< labels >>
rlabel pdiffusion 229 12 230 13  0 t = 1
rlabel pdiffusion 232 12 233 13  0 t = 2
rlabel pdiffusion 229 17 230 18  0 t = 3
rlabel pdiffusion 232 17 233 18  0 t = 4
rlabel pdiffusion 228 12 234 18 0 cell no = 8
<< m1 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2c >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< labels >>
rlabel pdiffusion 283 336 284 337  0 t = 1
rlabel pdiffusion 286 336 287 337  0 t = 2
rlabel pdiffusion 283 341 284 342  0 t = 3
rlabel pdiffusion 286 341 287 342  0 t = 4
rlabel pdiffusion 282 336 288 342 0 cell no = 9
<< m1 >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< m2 >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< m2c >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< labels >>
rlabel pdiffusion 103 192 104 193  0 t = 1
rlabel pdiffusion 106 192 107 193  0 t = 2
rlabel pdiffusion 103 197 104 198  0 t = 3
rlabel pdiffusion 106 197 107 198  0 t = 4
rlabel pdiffusion 102 192 108 198 0 cell no = 10
<< m1 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2c >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< labels >>
rlabel pdiffusion 49 318 50 319  0 t = 1
rlabel pdiffusion 52 318 53 319  0 t = 2
rlabel pdiffusion 49 323 50 324  0 t = 3
rlabel pdiffusion 52 323 53 324  0 t = 4
rlabel pdiffusion 48 318 54 324 0 cell no = 11
<< m1 >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< m2 >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< m2c >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 12
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 121 300 122 301  0 t = 1
rlabel pdiffusion 124 300 125 301  0 t = 2
rlabel pdiffusion 121 305 122 306  0 t = 3
rlabel pdiffusion 124 305 125 306  0 t = 4
rlabel pdiffusion 120 300 126 306 0 cell no = 13
<< m1 >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< m2 >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< m2c >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< labels >>
rlabel pdiffusion 211 84 212 85  0 t = 1
rlabel pdiffusion 214 84 215 85  0 t = 2
rlabel pdiffusion 211 89 212 90  0 t = 3
rlabel pdiffusion 214 89 215 90  0 t = 4
rlabel pdiffusion 210 84 216 90 0 cell no = 14
<< m1 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2c >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< labels >>
rlabel pdiffusion 283 210 284 211  0 t = 1
rlabel pdiffusion 286 210 287 211  0 t = 2
rlabel pdiffusion 283 215 284 216  0 t = 3
rlabel pdiffusion 286 215 287 216  0 t = 4
rlabel pdiffusion 282 210 288 216 0 cell no = 15
<< m1 >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< m2 >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< m2c >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< labels >>
rlabel pdiffusion 247 138 248 139  0 t = 1
rlabel pdiffusion 250 138 251 139  0 t = 2
rlabel pdiffusion 247 143 248 144  0 t = 3
rlabel pdiffusion 250 143 251 144  0 t = 4
rlabel pdiffusion 246 138 252 144 0 cell no = 16
<< m1 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2c >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< labels >>
rlabel pdiffusion 67 264 68 265  0 t = 1
rlabel pdiffusion 70 264 71 265  0 t = 2
rlabel pdiffusion 67 269 68 270  0 t = 3
rlabel pdiffusion 70 269 71 270  0 t = 4
rlabel pdiffusion 66 264 72 270 0 cell no = 17
<< m1 >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< m2 >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< m2c >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< labels >>
rlabel pdiffusion 247 174 248 175  0 t = 1
rlabel pdiffusion 250 174 251 175  0 t = 2
rlabel pdiffusion 247 179 248 180  0 t = 3
rlabel pdiffusion 250 179 251 180  0 t = 4
rlabel pdiffusion 246 174 252 180 0 cell no = 18
<< m1 >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< m2 >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< m2c >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< labels >>
rlabel pdiffusion 337 102 338 103  0 t = 1
rlabel pdiffusion 340 102 341 103  0 t = 2
rlabel pdiffusion 337 107 338 108  0 t = 3
rlabel pdiffusion 340 107 341 108  0 t = 4
rlabel pdiffusion 336 102 342 108 0 cell no = 19
<< m1 >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< m2 >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< m2c >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< labels >>
rlabel pdiffusion 175 174 176 175  0 t = 1
rlabel pdiffusion 178 174 179 175  0 t = 2
rlabel pdiffusion 175 179 176 180  0 t = 3
rlabel pdiffusion 178 179 179 180  0 t = 4
rlabel pdiffusion 174 174 180 180 0 cell no = 20
<< m1 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2c >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< labels >>
rlabel pdiffusion 229 318 230 319  0 t = 1
rlabel pdiffusion 232 318 233 319  0 t = 2
rlabel pdiffusion 229 323 230 324  0 t = 3
rlabel pdiffusion 232 323 233 324  0 t = 4
rlabel pdiffusion 228 318 234 324 0 cell no = 21
<< m1 >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< m2 >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< m2c >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< labels >>
rlabel pdiffusion 121 318 122 319  0 t = 1
rlabel pdiffusion 124 318 125 319  0 t = 2
rlabel pdiffusion 121 323 122 324  0 t = 3
rlabel pdiffusion 124 323 125 324  0 t = 4
rlabel pdiffusion 120 318 126 324 0 cell no = 22
<< m1 >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< m2 >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< m2c >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< labels >>
rlabel pdiffusion 337 84 338 85  0 t = 1
rlabel pdiffusion 340 84 341 85  0 t = 2
rlabel pdiffusion 337 89 338 90  0 t = 3
rlabel pdiffusion 340 89 341 90  0 t = 4
rlabel pdiffusion 336 84 342 90 0 cell no = 23
<< m1 >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< m2 >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< m2c >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< labels >>
rlabel pdiffusion 193 174 194 175  0 t = 1
rlabel pdiffusion 196 174 197 175  0 t = 2
rlabel pdiffusion 193 179 194 180  0 t = 3
rlabel pdiffusion 196 179 197 180  0 t = 4
rlabel pdiffusion 192 174 198 180 0 cell no = 24
<< m1 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2c >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< labels >>
rlabel pdiffusion 67 210 68 211  0 t = 1
rlabel pdiffusion 70 210 71 211  0 t = 2
rlabel pdiffusion 67 215 68 216  0 t = 3
rlabel pdiffusion 70 215 71 216  0 t = 4
rlabel pdiffusion 66 210 72 216 0 cell no = 25
<< m1 >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< m2 >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< m2c >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< labels >>
rlabel pdiffusion 121 228 122 229  0 t = 1
rlabel pdiffusion 124 228 125 229  0 t = 2
rlabel pdiffusion 121 233 122 234  0 t = 3
rlabel pdiffusion 124 233 125 234  0 t = 4
rlabel pdiffusion 120 228 126 234 0 cell no = 26
<< m1 >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< m2 >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< m2c >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< labels >>
rlabel pdiffusion 67 156 68 157  0 t = 1
rlabel pdiffusion 70 156 71 157  0 t = 2
rlabel pdiffusion 67 161 68 162  0 t = 3
rlabel pdiffusion 70 161 71 162  0 t = 4
rlabel pdiffusion 66 156 72 162 0 cell no = 27
<< m1 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2c >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< labels >>
rlabel pdiffusion 247 300 248 301  0 t = 1
rlabel pdiffusion 250 300 251 301  0 t = 2
rlabel pdiffusion 247 305 248 306  0 t = 3
rlabel pdiffusion 250 305 251 306  0 t = 4
rlabel pdiffusion 246 300 252 306 0 cell no = 28
<< m1 >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< m2 >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< m2c >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< labels >>
rlabel pdiffusion 139 102 140 103  0 t = 1
rlabel pdiffusion 142 102 143 103  0 t = 2
rlabel pdiffusion 139 107 140 108  0 t = 3
rlabel pdiffusion 142 107 143 108  0 t = 4
rlabel pdiffusion 138 102 144 108 0 cell no = 29
<< m1 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2c >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< labels >>
rlabel pdiffusion 229 156 230 157  0 t = 1
rlabel pdiffusion 232 156 233 157  0 t = 2
rlabel pdiffusion 229 161 230 162  0 t = 3
rlabel pdiffusion 232 161 233 162  0 t = 4
rlabel pdiffusion 228 156 234 162 0 cell no = 30
<< m1 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2c >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< labels >>
rlabel pdiffusion 49 300 50 301  0 t = 1
rlabel pdiffusion 52 300 53 301  0 t = 2
rlabel pdiffusion 49 305 50 306  0 t = 3
rlabel pdiffusion 52 305 53 306  0 t = 4
rlabel pdiffusion 48 300 54 306 0 cell no = 31
<< m1 >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< m2 >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< m2c >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< labels >>
rlabel pdiffusion 319 174 320 175  0 t = 1
rlabel pdiffusion 322 174 323 175  0 t = 2
rlabel pdiffusion 319 179 320 180  0 t = 3
rlabel pdiffusion 322 179 323 180  0 t = 4
rlabel pdiffusion 318 174 324 180 0 cell no = 32
<< m1 >>
rect 319 174 320 175 
rect 322 174 323 175 
rect 319 179 320 180 
rect 322 179 323 180 
<< m2 >>
rect 319 174 320 175 
rect 322 174 323 175 
rect 319 179 320 180 
rect 322 179 323 180 
<< m2c >>
rect 319 174 320 175 
rect 322 174 323 175 
rect 319 179 320 180 
rect 322 179 323 180 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 33
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 283 12 284 13  0 t = 1
rlabel pdiffusion 286 12 287 13  0 t = 2
rlabel pdiffusion 283 17 284 18  0 t = 3
rlabel pdiffusion 286 17 287 18  0 t = 4
rlabel pdiffusion 282 12 288 18 0 cell no = 34
<< m1 >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< m2 >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< m2c >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< labels >>
rlabel pdiffusion 283 138 284 139  0 t = 1
rlabel pdiffusion 286 138 287 139  0 t = 2
rlabel pdiffusion 283 143 284 144  0 t = 3
rlabel pdiffusion 286 143 287 144  0 t = 4
rlabel pdiffusion 282 138 288 144 0 cell no = 35
<< m1 >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< m2 >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< m2c >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< labels >>
rlabel pdiffusion 193 300 194 301  0 t = 1
rlabel pdiffusion 196 300 197 301  0 t = 2
rlabel pdiffusion 193 305 194 306  0 t = 3
rlabel pdiffusion 196 305 197 306  0 t = 4
rlabel pdiffusion 192 300 198 306 0 cell no = 36
<< m1 >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< m2 >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< m2c >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< labels >>
rlabel pdiffusion 319 120 320 121  0 t = 1
rlabel pdiffusion 322 120 323 121  0 t = 2
rlabel pdiffusion 319 125 320 126  0 t = 3
rlabel pdiffusion 322 125 323 126  0 t = 4
rlabel pdiffusion 318 120 324 126 0 cell no = 37
<< m1 >>
rect 319 120 320 121 
rect 322 120 323 121 
rect 319 125 320 126 
rect 322 125 323 126 
<< m2 >>
rect 319 120 320 121 
rect 322 120 323 121 
rect 319 125 320 126 
rect 322 125 323 126 
<< m2c >>
rect 319 120 320 121 
rect 322 120 323 121 
rect 319 125 320 126 
rect 322 125 323 126 
<< labels >>
rlabel pdiffusion 175 228 176 229  0 t = 1
rlabel pdiffusion 178 228 179 229  0 t = 2
rlabel pdiffusion 175 233 176 234  0 t = 3
rlabel pdiffusion 178 233 179 234  0 t = 4
rlabel pdiffusion 174 228 180 234 0 cell no = 38
<< m1 >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< m2 >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< m2c >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 39
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 211 12 212 13  0 t = 1
rlabel pdiffusion 214 12 215 13  0 t = 2
rlabel pdiffusion 211 17 212 18  0 t = 3
rlabel pdiffusion 214 17 215 18  0 t = 4
rlabel pdiffusion 210 12 216 18 0 cell no = 40
<< m1 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2c >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< labels >>
rlabel pdiffusion 319 138 320 139  0 t = 1
rlabel pdiffusion 322 138 323 139  0 t = 2
rlabel pdiffusion 319 143 320 144  0 t = 3
rlabel pdiffusion 322 143 323 144  0 t = 4
rlabel pdiffusion 318 138 324 144 0 cell no = 41
<< m1 >>
rect 319 138 320 139 
rect 322 138 323 139 
rect 319 143 320 144 
rect 322 143 323 144 
<< m2 >>
rect 319 138 320 139 
rect 322 138 323 139 
rect 319 143 320 144 
rect 322 143 323 144 
<< m2c >>
rect 319 138 320 139 
rect 322 138 323 139 
rect 319 143 320 144 
rect 322 143 323 144 
<< labels >>
rlabel pdiffusion 31 156 32 157  0 t = 1
rlabel pdiffusion 34 156 35 157  0 t = 2
rlabel pdiffusion 31 161 32 162  0 t = 3
rlabel pdiffusion 34 161 35 162  0 t = 4
rlabel pdiffusion 30 156 36 162 0 cell no = 42
<< m1 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2c >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< labels >>
rlabel pdiffusion 337 264 338 265  0 t = 1
rlabel pdiffusion 340 264 341 265  0 t = 2
rlabel pdiffusion 337 269 338 270  0 t = 3
rlabel pdiffusion 340 269 341 270  0 t = 4
rlabel pdiffusion 336 264 342 270 0 cell no = 43
<< m1 >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< m2 >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< m2c >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< labels >>
rlabel pdiffusion 193 102 194 103  0 t = 1
rlabel pdiffusion 196 102 197 103  0 t = 2
rlabel pdiffusion 193 107 194 108  0 t = 3
rlabel pdiffusion 196 107 197 108  0 t = 4
rlabel pdiffusion 192 102 198 108 0 cell no = 44
<< m1 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2c >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< labels >>
rlabel pdiffusion 301 264 302 265  0 t = 1
rlabel pdiffusion 304 264 305 265  0 t = 2
rlabel pdiffusion 301 269 302 270  0 t = 3
rlabel pdiffusion 304 269 305 270  0 t = 4
rlabel pdiffusion 300 264 306 270 0 cell no = 45
<< m1 >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< m2 >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< m2c >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< labels >>
rlabel pdiffusion 211 120 212 121  0 t = 1
rlabel pdiffusion 214 120 215 121  0 t = 2
rlabel pdiffusion 211 125 212 126  0 t = 3
rlabel pdiffusion 214 125 215 126  0 t = 4
rlabel pdiffusion 210 120 216 126 0 cell no = 46
<< m1 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2c >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< labels >>
rlabel pdiffusion 319 66 320 67  0 t = 1
rlabel pdiffusion 322 66 323 67  0 t = 2
rlabel pdiffusion 319 71 320 72  0 t = 3
rlabel pdiffusion 322 71 323 72  0 t = 4
rlabel pdiffusion 318 66 324 72 0 cell no = 47
<< m1 >>
rect 319 66 320 67 
rect 322 66 323 67 
rect 319 71 320 72 
rect 322 71 323 72 
<< m2 >>
rect 319 66 320 67 
rect 322 66 323 67 
rect 319 71 320 72 
rect 322 71 323 72 
<< m2c >>
rect 319 66 320 67 
rect 322 66 323 67 
rect 319 71 320 72 
rect 322 71 323 72 
<< labels >>
rlabel pdiffusion 31 30 32 31  0 t = 1
rlabel pdiffusion 34 30 35 31  0 t = 2
rlabel pdiffusion 31 35 32 36  0 t = 3
rlabel pdiffusion 34 35 35 36  0 t = 4
rlabel pdiffusion 30 30 36 36 0 cell no = 48
<< m1 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2c >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< labels >>
rlabel pdiffusion 67 282 68 283  0 t = 1
rlabel pdiffusion 70 282 71 283  0 t = 2
rlabel pdiffusion 67 287 68 288  0 t = 3
rlabel pdiffusion 70 287 71 288  0 t = 4
rlabel pdiffusion 66 282 72 288 0 cell no = 49
<< m1 >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< m2 >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< m2c >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< labels >>
rlabel pdiffusion 139 282 140 283  0 t = 1
rlabel pdiffusion 142 282 143 283  0 t = 2
rlabel pdiffusion 139 287 140 288  0 t = 3
rlabel pdiffusion 142 287 143 288  0 t = 4
rlabel pdiffusion 138 282 144 288 0 cell no = 50
<< m1 >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< m2 >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< m2c >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< labels >>
rlabel pdiffusion 103 120 104 121  0 t = 1
rlabel pdiffusion 106 120 107 121  0 t = 2
rlabel pdiffusion 103 125 104 126  0 t = 3
rlabel pdiffusion 106 125 107 126  0 t = 4
rlabel pdiffusion 102 120 108 126 0 cell no = 51
<< m1 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2c >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< labels >>
rlabel pdiffusion 31 300 32 301  0 t = 1
rlabel pdiffusion 34 300 35 301  0 t = 2
rlabel pdiffusion 31 305 32 306  0 t = 3
rlabel pdiffusion 34 305 35 306  0 t = 4
rlabel pdiffusion 30 300 36 306 0 cell no = 52
<< m1 >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< m2 >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< m2c >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< labels >>
rlabel pdiffusion 247 192 248 193  0 t = 1
rlabel pdiffusion 250 192 251 193  0 t = 2
rlabel pdiffusion 247 197 248 198  0 t = 3
rlabel pdiffusion 250 197 251 198  0 t = 4
rlabel pdiffusion 246 192 252 198 0 cell no = 53
<< m1 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2c >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< labels >>
rlabel pdiffusion 247 120 248 121  0 t = 1
rlabel pdiffusion 250 120 251 121  0 t = 2
rlabel pdiffusion 247 125 248 126  0 t = 3
rlabel pdiffusion 250 125 251 126  0 t = 4
rlabel pdiffusion 246 120 252 126 0 cell no = 54
<< m1 >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< m2 >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< m2c >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< labels >>
rlabel pdiffusion 13 264 14 265  0 t = 1
rlabel pdiffusion 16 264 17 265  0 t = 2
rlabel pdiffusion 13 269 14 270  0 t = 3
rlabel pdiffusion 16 269 17 270  0 t = 4
rlabel pdiffusion 12 264 18 270 0 cell no = 55
<< m1 >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< m2 >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< m2c >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< labels >>
rlabel pdiffusion 319 12 320 13  0 t = 1
rlabel pdiffusion 322 12 323 13  0 t = 2
rlabel pdiffusion 319 17 320 18  0 t = 3
rlabel pdiffusion 322 17 323 18  0 t = 4
rlabel pdiffusion 318 12 324 18 0 cell no = 56
<< m1 >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< m2 >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< m2c >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< labels >>
rlabel pdiffusion 13 156 14 157  0 t = 1
rlabel pdiffusion 16 156 17 157  0 t = 2
rlabel pdiffusion 13 161 14 162  0 t = 3
rlabel pdiffusion 16 161 17 162  0 t = 4
rlabel pdiffusion 12 156 18 162 0 cell no = 57
<< m1 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2c >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< labels >>
rlabel pdiffusion 175 30 176 31  0 t = 1
rlabel pdiffusion 178 30 179 31  0 t = 2
rlabel pdiffusion 175 35 176 36  0 t = 3
rlabel pdiffusion 178 35 179 36  0 t = 4
rlabel pdiffusion 174 30 180 36 0 cell no = 58
<< m1 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2c >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< labels >>
rlabel pdiffusion 247 30 248 31  0 t = 1
rlabel pdiffusion 250 30 251 31  0 t = 2
rlabel pdiffusion 247 35 248 36  0 t = 3
rlabel pdiffusion 250 35 251 36  0 t = 4
rlabel pdiffusion 246 30 252 36 0 cell no = 59
<< m1 >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< m2 >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< m2c >>
rect 247 30 248 31 
rect 250 30 251 31 
rect 247 35 248 36 
rect 250 35 251 36 
<< labels >>
rlabel pdiffusion 265 246 266 247  0 t = 1
rlabel pdiffusion 268 246 269 247  0 t = 2
rlabel pdiffusion 265 251 266 252  0 t = 3
rlabel pdiffusion 268 251 269 252  0 t = 4
rlabel pdiffusion 264 246 270 252 0 cell no = 60
<< m1 >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< m2 >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< m2c >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< labels >>
rlabel pdiffusion 211 102 212 103  0 t = 1
rlabel pdiffusion 214 102 215 103  0 t = 2
rlabel pdiffusion 211 107 212 108  0 t = 3
rlabel pdiffusion 214 107 215 108  0 t = 4
rlabel pdiffusion 210 102 216 108 0 cell no = 61
<< m1 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2c >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< labels >>
rlabel pdiffusion 67 138 68 139  0 t = 1
rlabel pdiffusion 70 138 71 139  0 t = 2
rlabel pdiffusion 67 143 68 144  0 t = 3
rlabel pdiffusion 70 143 71 144  0 t = 4
rlabel pdiffusion 66 138 72 144 0 cell no = 62
<< m1 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2c >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 63
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 64
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 211 282 212 283  0 t = 1
rlabel pdiffusion 214 282 215 283  0 t = 2
rlabel pdiffusion 211 287 212 288  0 t = 3
rlabel pdiffusion 214 287 215 288  0 t = 4
rlabel pdiffusion 210 282 216 288 0 cell no = 65
<< m1 >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< m2 >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< m2c >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< labels >>
rlabel pdiffusion 121 264 122 265  0 t = 1
rlabel pdiffusion 124 264 125 265  0 t = 2
rlabel pdiffusion 121 269 122 270  0 t = 3
rlabel pdiffusion 124 269 125 270  0 t = 4
rlabel pdiffusion 120 264 126 270 0 cell no = 66
<< m1 >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< m2 >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< m2c >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 67
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 211 210 212 211  0 t = 1
rlabel pdiffusion 214 210 215 211  0 t = 2
rlabel pdiffusion 211 215 212 216  0 t = 3
rlabel pdiffusion 214 215 215 216  0 t = 4
rlabel pdiffusion 210 210 216 216 0 cell no = 68
<< m1 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2c >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< labels >>
rlabel pdiffusion 229 282 230 283  0 t = 1
rlabel pdiffusion 232 282 233 283  0 t = 2
rlabel pdiffusion 229 287 230 288  0 t = 3
rlabel pdiffusion 232 287 233 288  0 t = 4
rlabel pdiffusion 228 282 234 288 0 cell no = 69
<< m1 >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< m2 >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< m2c >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< labels >>
rlabel pdiffusion 13 246 14 247  0 t = 1
rlabel pdiffusion 16 246 17 247  0 t = 2
rlabel pdiffusion 13 251 14 252  0 t = 3
rlabel pdiffusion 16 251 17 252  0 t = 4
rlabel pdiffusion 12 246 18 252 0 cell no = 70
<< m1 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2c >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< labels >>
rlabel pdiffusion 301 246 302 247  0 t = 1
rlabel pdiffusion 304 246 305 247  0 t = 2
rlabel pdiffusion 301 251 302 252  0 t = 3
rlabel pdiffusion 304 251 305 252  0 t = 4
rlabel pdiffusion 300 246 306 252 0 cell no = 71
<< m1 >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< m2 >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< m2c >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< labels >>
rlabel pdiffusion 193 30 194 31  0 t = 1
rlabel pdiffusion 196 30 197 31  0 t = 2
rlabel pdiffusion 193 35 194 36  0 t = 3
rlabel pdiffusion 196 35 197 36  0 t = 4
rlabel pdiffusion 192 30 198 36 0 cell no = 72
<< m1 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2c >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< labels >>
rlabel pdiffusion 283 66 284 67  0 t = 1
rlabel pdiffusion 286 66 287 67  0 t = 2
rlabel pdiffusion 283 71 284 72  0 t = 3
rlabel pdiffusion 286 71 287 72  0 t = 4
rlabel pdiffusion 282 66 288 72 0 cell no = 73
<< m1 >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< m2 >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< m2c >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< labels >>
rlabel pdiffusion 121 246 122 247  0 t = 1
rlabel pdiffusion 124 246 125 247  0 t = 2
rlabel pdiffusion 121 251 122 252  0 t = 3
rlabel pdiffusion 124 251 125 252  0 t = 4
rlabel pdiffusion 120 246 126 252 0 cell no = 74
<< m1 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2c >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< labels >>
rlabel pdiffusion 229 138 230 139  0 t = 1
rlabel pdiffusion 232 138 233 139  0 t = 2
rlabel pdiffusion 229 143 230 144  0 t = 3
rlabel pdiffusion 232 143 233 144  0 t = 4
rlabel pdiffusion 228 138 234 144 0 cell no = 75
<< m1 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2c >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 76
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 139 138 140 139  0 t = 1
rlabel pdiffusion 142 138 143 139  0 t = 2
rlabel pdiffusion 139 143 140 144  0 t = 3
rlabel pdiffusion 142 143 143 144  0 t = 4
rlabel pdiffusion 138 138 144 144 0 cell no = 77
<< m1 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2c >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< labels >>
rlabel pdiffusion 265 48 266 49  0 t = 1
rlabel pdiffusion 268 48 269 49  0 t = 2
rlabel pdiffusion 265 53 266 54  0 t = 3
rlabel pdiffusion 268 53 269 54  0 t = 4
rlabel pdiffusion 264 48 270 54 0 cell no = 78
<< m1 >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< m2 >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< m2c >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< labels >>
rlabel pdiffusion 67 228 68 229  0 t = 1
rlabel pdiffusion 70 228 71 229  0 t = 2
rlabel pdiffusion 67 233 68 234  0 t = 3
rlabel pdiffusion 70 233 71 234  0 t = 4
rlabel pdiffusion 66 228 72 234 0 cell no = 79
<< m1 >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< m2 >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< m2c >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< labels >>
rlabel pdiffusion 301 66 302 67  0 t = 1
rlabel pdiffusion 304 66 305 67  0 t = 2
rlabel pdiffusion 301 71 302 72  0 t = 3
rlabel pdiffusion 304 71 305 72  0 t = 4
rlabel pdiffusion 300 66 306 72 0 cell no = 80
<< m1 >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< m2 >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< m2c >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< labels >>
rlabel pdiffusion 49 282 50 283  0 t = 1
rlabel pdiffusion 52 282 53 283  0 t = 2
rlabel pdiffusion 49 287 50 288  0 t = 3
rlabel pdiffusion 52 287 53 288  0 t = 4
rlabel pdiffusion 48 282 54 288 0 cell no = 81
<< m1 >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< m2 >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< m2c >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< labels >>
rlabel pdiffusion 301 300 302 301  0 t = 1
rlabel pdiffusion 304 300 305 301  0 t = 2
rlabel pdiffusion 301 305 302 306  0 t = 3
rlabel pdiffusion 304 305 305 306  0 t = 4
rlabel pdiffusion 300 300 306 306 0 cell no = 82
<< m1 >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< m2 >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< m2c >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< labels >>
rlabel pdiffusion 157 48 158 49  0 t = 1
rlabel pdiffusion 160 48 161 49  0 t = 2
rlabel pdiffusion 157 53 158 54  0 t = 3
rlabel pdiffusion 160 53 161 54  0 t = 4
rlabel pdiffusion 156 48 162 54 0 cell no = 83
<< m1 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2c >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< labels >>
rlabel pdiffusion 121 210 122 211  0 t = 1
rlabel pdiffusion 124 210 125 211  0 t = 2
rlabel pdiffusion 121 215 122 216  0 t = 3
rlabel pdiffusion 124 215 125 216  0 t = 4
rlabel pdiffusion 120 210 126 216 0 cell no = 84
<< m1 >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< m2 >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< m2c >>
rect 121 210 122 211 
rect 124 210 125 211 
rect 121 215 122 216 
rect 124 215 125 216 
<< labels >>
rlabel pdiffusion 157 282 158 283  0 t = 1
rlabel pdiffusion 160 282 161 283  0 t = 2
rlabel pdiffusion 157 287 158 288  0 t = 3
rlabel pdiffusion 160 287 161 288  0 t = 4
rlabel pdiffusion 156 282 162 288 0 cell no = 85
<< m1 >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< m2 >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< m2c >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 86
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 319 30 320 31  0 t = 1
rlabel pdiffusion 322 30 323 31  0 t = 2
rlabel pdiffusion 319 35 320 36  0 t = 3
rlabel pdiffusion 322 35 323 36  0 t = 4
rlabel pdiffusion 318 30 324 36 0 cell no = 87
<< m1 >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< m2 >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< m2c >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< labels >>
rlabel pdiffusion 229 84 230 85  0 t = 1
rlabel pdiffusion 232 84 233 85  0 t = 2
rlabel pdiffusion 229 89 230 90  0 t = 3
rlabel pdiffusion 232 89 233 90  0 t = 4
rlabel pdiffusion 228 84 234 90 0 cell no = 88
<< m1 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2c >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< labels >>
rlabel pdiffusion 319 228 320 229  0 t = 1
rlabel pdiffusion 322 228 323 229  0 t = 2
rlabel pdiffusion 319 233 320 234  0 t = 3
rlabel pdiffusion 322 233 323 234  0 t = 4
rlabel pdiffusion 318 228 324 234 0 cell no = 89
<< m1 >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< m2 >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< m2c >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< labels >>
rlabel pdiffusion 103 156 104 157  0 t = 1
rlabel pdiffusion 106 156 107 157  0 t = 2
rlabel pdiffusion 103 161 104 162  0 t = 3
rlabel pdiffusion 106 161 107 162  0 t = 4
rlabel pdiffusion 102 156 108 162 0 cell no = 90
<< m1 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2c >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< labels >>
rlabel pdiffusion 139 174 140 175  0 t = 1
rlabel pdiffusion 142 174 143 175  0 t = 2
rlabel pdiffusion 139 179 140 180  0 t = 3
rlabel pdiffusion 142 179 143 180  0 t = 4
rlabel pdiffusion 138 174 144 180 0 cell no = 91
<< m1 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2c >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< labels >>
rlabel pdiffusion 301 318 302 319  0 t = 1
rlabel pdiffusion 304 318 305 319  0 t = 2
rlabel pdiffusion 301 323 302 324  0 t = 3
rlabel pdiffusion 304 323 305 324  0 t = 4
rlabel pdiffusion 300 318 306 324 0 cell no = 92
<< m1 >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< m2 >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< m2c >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< labels >>
rlabel pdiffusion 337 318 338 319  0 t = 1
rlabel pdiffusion 340 318 341 319  0 t = 2
rlabel pdiffusion 337 323 338 324  0 t = 3
rlabel pdiffusion 340 323 341 324  0 t = 4
rlabel pdiffusion 336 318 342 324 0 cell no = 93
<< m1 >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< m2 >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< m2c >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< labels >>
rlabel pdiffusion 13 282 14 283  0 t = 1
rlabel pdiffusion 16 282 17 283  0 t = 2
rlabel pdiffusion 13 287 14 288  0 t = 3
rlabel pdiffusion 16 287 17 288  0 t = 4
rlabel pdiffusion 12 282 18 288 0 cell no = 94
<< m1 >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< m2 >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< m2c >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< labels >>
rlabel pdiffusion 85 336 86 337  0 t = 1
rlabel pdiffusion 88 336 89 337  0 t = 2
rlabel pdiffusion 85 341 86 342  0 t = 3
rlabel pdiffusion 88 341 89 342  0 t = 4
rlabel pdiffusion 84 336 90 342 0 cell no = 95
<< m1 >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< m2 >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< m2c >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< labels >>
rlabel pdiffusion 139 246 140 247  0 t = 1
rlabel pdiffusion 142 246 143 247  0 t = 2
rlabel pdiffusion 139 251 140 252  0 t = 3
rlabel pdiffusion 142 251 143 252  0 t = 4
rlabel pdiffusion 138 246 144 252 0 cell no = 96
<< m1 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2c >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< labels >>
rlabel pdiffusion 283 228 284 229  0 t = 1
rlabel pdiffusion 286 228 287 229  0 t = 2
rlabel pdiffusion 283 233 284 234  0 t = 3
rlabel pdiffusion 286 233 287 234  0 t = 4
rlabel pdiffusion 282 228 288 234 0 cell no = 97
<< m1 >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< m2 >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< m2c >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< labels >>
rlabel pdiffusion 193 318 194 319  0 t = 1
rlabel pdiffusion 196 318 197 319  0 t = 2
rlabel pdiffusion 193 323 194 324  0 t = 3
rlabel pdiffusion 196 323 197 324  0 t = 4
rlabel pdiffusion 192 318 198 324 0 cell no = 98
<< m1 >>
rect 193 318 194 319 
rect 196 318 197 319 
rect 193 323 194 324 
rect 196 323 197 324 
<< m2 >>
rect 193 318 194 319 
rect 196 318 197 319 
rect 193 323 194 324 
rect 196 323 197 324 
<< m2c >>
rect 193 318 194 319 
rect 196 318 197 319 
rect 193 323 194 324 
rect 196 323 197 324 
<< labels >>
rlabel pdiffusion 157 264 158 265  0 t = 1
rlabel pdiffusion 160 264 161 265  0 t = 2
rlabel pdiffusion 157 269 158 270  0 t = 3
rlabel pdiffusion 160 269 161 270  0 t = 4
rlabel pdiffusion 156 264 162 270 0 cell no = 99
<< m1 >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< m2 >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< m2c >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< labels >>
rlabel pdiffusion 337 210 338 211  0 t = 1
rlabel pdiffusion 340 210 341 211  0 t = 2
rlabel pdiffusion 337 215 338 216  0 t = 3
rlabel pdiffusion 340 215 341 216  0 t = 4
rlabel pdiffusion 336 210 342 216 0 cell no = 100
<< m1 >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< m2 >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< m2c >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< labels >>
rlabel pdiffusion 67 246 68 247  0 t = 1
rlabel pdiffusion 70 246 71 247  0 t = 2
rlabel pdiffusion 67 251 68 252  0 t = 3
rlabel pdiffusion 70 251 71 252  0 t = 4
rlabel pdiffusion 66 246 72 252 0 cell no = 101
<< m1 >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< m2 >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< m2c >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< labels >>
rlabel pdiffusion 31 282 32 283  0 t = 1
rlabel pdiffusion 34 282 35 283  0 t = 2
rlabel pdiffusion 31 287 32 288  0 t = 3
rlabel pdiffusion 34 287 35 288  0 t = 4
rlabel pdiffusion 30 282 36 288 0 cell no = 102
<< m1 >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< m2 >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< m2c >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< labels >>
rlabel pdiffusion 157 246 158 247  0 t = 1
rlabel pdiffusion 160 246 161 247  0 t = 2
rlabel pdiffusion 157 251 158 252  0 t = 3
rlabel pdiffusion 160 251 161 252  0 t = 4
rlabel pdiffusion 156 246 162 252 0 cell no = 103
<< m1 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2c >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< labels >>
rlabel pdiffusion 31 246 32 247  0 t = 1
rlabel pdiffusion 34 246 35 247  0 t = 2
rlabel pdiffusion 31 251 32 252  0 t = 3
rlabel pdiffusion 34 251 35 252  0 t = 4
rlabel pdiffusion 30 246 36 252 0 cell no = 104
<< m1 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2c >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< labels >>
rlabel pdiffusion 121 138 122 139  0 t = 1
rlabel pdiffusion 124 138 125 139  0 t = 2
rlabel pdiffusion 121 143 122 144  0 t = 3
rlabel pdiffusion 124 143 125 144  0 t = 4
rlabel pdiffusion 120 138 126 144 0 cell no = 105
<< m1 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2c >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< labels >>
rlabel pdiffusion 193 210 194 211  0 t = 1
rlabel pdiffusion 196 210 197 211  0 t = 2
rlabel pdiffusion 193 215 194 216  0 t = 3
rlabel pdiffusion 196 215 197 216  0 t = 4
rlabel pdiffusion 192 210 198 216 0 cell no = 106
<< m1 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2c >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< labels >>
rlabel pdiffusion 337 300 338 301  0 t = 1
rlabel pdiffusion 340 300 341 301  0 t = 2
rlabel pdiffusion 337 305 338 306  0 t = 3
rlabel pdiffusion 340 305 341 306  0 t = 4
rlabel pdiffusion 336 300 342 306 0 cell no = 107
<< m1 >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< m2 >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< m2c >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< labels >>
rlabel pdiffusion 157 84 158 85  0 t = 1
rlabel pdiffusion 160 84 161 85  0 t = 2
rlabel pdiffusion 157 89 158 90  0 t = 3
rlabel pdiffusion 160 89 161 90  0 t = 4
rlabel pdiffusion 156 84 162 90 0 cell no = 108
<< m1 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2c >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< labels >>
rlabel pdiffusion 103 282 104 283  0 t = 1
rlabel pdiffusion 106 282 107 283  0 t = 2
rlabel pdiffusion 103 287 104 288  0 t = 3
rlabel pdiffusion 106 287 107 288  0 t = 4
rlabel pdiffusion 102 282 108 288 0 cell no = 109
<< m1 >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< m2 >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< m2c >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< labels >>
rlabel pdiffusion 103 300 104 301  0 t = 1
rlabel pdiffusion 106 300 107 301  0 t = 2
rlabel pdiffusion 103 305 104 306  0 t = 3
rlabel pdiffusion 106 305 107 306  0 t = 4
rlabel pdiffusion 102 300 108 306 0 cell no = 110
<< m1 >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< m2 >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< m2c >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< labels >>
rlabel pdiffusion 67 192 68 193  0 t = 1
rlabel pdiffusion 70 192 71 193  0 t = 2
rlabel pdiffusion 67 197 68 198  0 t = 3
rlabel pdiffusion 70 197 71 198  0 t = 4
rlabel pdiffusion 66 192 72 198 0 cell no = 111
<< m1 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2c >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< labels >>
rlabel pdiffusion 247 12 248 13  0 t = 1
rlabel pdiffusion 250 12 251 13  0 t = 2
rlabel pdiffusion 247 17 248 18  0 t = 3
rlabel pdiffusion 250 17 251 18  0 t = 4
rlabel pdiffusion 246 12 252 18 0 cell no = 112
<< m1 >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< m2 >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< m2c >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< labels >>
rlabel pdiffusion 85 282 86 283  0 t = 1
rlabel pdiffusion 88 282 89 283  0 t = 2
rlabel pdiffusion 85 287 86 288  0 t = 3
rlabel pdiffusion 88 287 89 288  0 t = 4
rlabel pdiffusion 84 282 90 288 0 cell no = 113
<< m1 >>
rect 85 282 86 283 
rect 88 282 89 283 
rect 85 287 86 288 
rect 88 287 89 288 
<< m2 >>
rect 85 282 86 283 
rect 88 282 89 283 
rect 85 287 86 288 
rect 88 287 89 288 
<< m2c >>
rect 85 282 86 283 
rect 88 282 89 283 
rect 85 287 86 288 
rect 88 287 89 288 
<< labels >>
rlabel pdiffusion 85 120 86 121  0 t = 1
rlabel pdiffusion 88 120 89 121  0 t = 2
rlabel pdiffusion 85 125 86 126  0 t = 3
rlabel pdiffusion 88 125 89 126  0 t = 4
rlabel pdiffusion 84 120 90 126 0 cell no = 114
<< m1 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2c >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< labels >>
rlabel pdiffusion 247 282 248 283  0 t = 1
rlabel pdiffusion 250 282 251 283  0 t = 2
rlabel pdiffusion 247 287 248 288  0 t = 3
rlabel pdiffusion 250 287 251 288  0 t = 4
rlabel pdiffusion 246 282 252 288 0 cell no = 115
<< m1 >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< m2 >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< m2c >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< labels >>
rlabel pdiffusion 247 264 248 265  0 t = 1
rlabel pdiffusion 250 264 251 265  0 t = 2
rlabel pdiffusion 247 269 248 270  0 t = 3
rlabel pdiffusion 250 269 251 270  0 t = 4
rlabel pdiffusion 246 264 252 270 0 cell no = 116
<< m1 >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< m2 >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< m2c >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< labels >>
rlabel pdiffusion 319 282 320 283  0 t = 1
rlabel pdiffusion 322 282 323 283  0 t = 2
rlabel pdiffusion 319 287 320 288  0 t = 3
rlabel pdiffusion 322 287 323 288  0 t = 4
rlabel pdiffusion 318 282 324 288 0 cell no = 117
<< m1 >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< m2 >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< m2c >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< labels >>
rlabel pdiffusion 175 12 176 13  0 t = 1
rlabel pdiffusion 178 12 179 13  0 t = 2
rlabel pdiffusion 175 17 176 18  0 t = 3
rlabel pdiffusion 178 17 179 18  0 t = 4
rlabel pdiffusion 174 12 180 18 0 cell no = 118
<< m1 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2c >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< labels >>
rlabel pdiffusion 337 282 338 283  0 t = 1
rlabel pdiffusion 340 282 341 283  0 t = 2
rlabel pdiffusion 337 287 338 288  0 t = 3
rlabel pdiffusion 340 287 341 288  0 t = 4
rlabel pdiffusion 336 282 342 288 0 cell no = 119
<< m1 >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< m2 >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< m2c >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< labels >>
rlabel pdiffusion 229 264 230 265  0 t = 1
rlabel pdiffusion 232 264 233 265  0 t = 2
rlabel pdiffusion 229 269 230 270  0 t = 3
rlabel pdiffusion 232 269 233 270  0 t = 4
rlabel pdiffusion 228 264 234 270 0 cell no = 120
<< m1 >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< m2 >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< m2c >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< labels >>
rlabel pdiffusion 229 120 230 121  0 t = 1
rlabel pdiffusion 232 120 233 121  0 t = 2
rlabel pdiffusion 229 125 230 126  0 t = 3
rlabel pdiffusion 232 125 233 126  0 t = 4
rlabel pdiffusion 228 120 234 126 0 cell no = 121
<< m1 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2c >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< labels >>
rlabel pdiffusion 139 66 140 67  0 t = 1
rlabel pdiffusion 142 66 143 67  0 t = 2
rlabel pdiffusion 139 71 140 72  0 t = 3
rlabel pdiffusion 142 71 143 72  0 t = 4
rlabel pdiffusion 138 66 144 72 0 cell no = 122
<< m1 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2c >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< labels >>
rlabel pdiffusion 229 102 230 103  0 t = 1
rlabel pdiffusion 232 102 233 103  0 t = 2
rlabel pdiffusion 229 107 230 108  0 t = 3
rlabel pdiffusion 232 107 233 108  0 t = 4
rlabel pdiffusion 228 102 234 108 0 cell no = 123
<< m1 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2c >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< labels >>
rlabel pdiffusion 49 138 50 139  0 t = 1
rlabel pdiffusion 52 138 53 139  0 t = 2
rlabel pdiffusion 49 143 50 144  0 t = 3
rlabel pdiffusion 52 143 53 144  0 t = 4
rlabel pdiffusion 48 138 54 144 0 cell no = 124
<< m1 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2c >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< labels >>
rlabel pdiffusion 337 228 338 229  0 t = 1
rlabel pdiffusion 340 228 341 229  0 t = 2
rlabel pdiffusion 337 233 338 234  0 t = 3
rlabel pdiffusion 340 233 341 234  0 t = 4
rlabel pdiffusion 336 228 342 234 0 cell no = 125
<< m1 >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< m2 >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< m2c >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< labels >>
rlabel pdiffusion 193 84 194 85  0 t = 1
rlabel pdiffusion 196 84 197 85  0 t = 2
rlabel pdiffusion 193 89 194 90  0 t = 3
rlabel pdiffusion 196 89 197 90  0 t = 4
rlabel pdiffusion 192 84 198 90 0 cell no = 126
<< m1 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2c >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< labels >>
rlabel pdiffusion 265 318 266 319  0 t = 1
rlabel pdiffusion 268 318 269 319  0 t = 2
rlabel pdiffusion 265 323 266 324  0 t = 3
rlabel pdiffusion 268 323 269 324  0 t = 4
rlabel pdiffusion 264 318 270 324 0 cell no = 127
<< m1 >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< m2 >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< m2c >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< labels >>
rlabel pdiffusion 85 300 86 301  0 t = 1
rlabel pdiffusion 88 300 89 301  0 t = 2
rlabel pdiffusion 85 305 86 306  0 t = 3
rlabel pdiffusion 88 305 89 306  0 t = 4
rlabel pdiffusion 84 300 90 306 0 cell no = 128
<< m1 >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< m2 >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< m2c >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< labels >>
rlabel pdiffusion 157 30 158 31  0 t = 1
rlabel pdiffusion 160 30 161 31  0 t = 2
rlabel pdiffusion 157 35 158 36  0 t = 3
rlabel pdiffusion 160 35 161 36  0 t = 4
rlabel pdiffusion 156 30 162 36 0 cell no = 129
<< m1 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2c >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< labels >>
rlabel pdiffusion 265 120 266 121  0 t = 1
rlabel pdiffusion 268 120 269 121  0 t = 2
rlabel pdiffusion 265 125 266 126  0 t = 3
rlabel pdiffusion 268 125 269 126  0 t = 4
rlabel pdiffusion 264 120 270 126 0 cell no = 130
<< m1 >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< m2 >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< m2c >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< labels >>
rlabel pdiffusion 283 120 284 121  0 t = 1
rlabel pdiffusion 286 120 287 121  0 t = 2
rlabel pdiffusion 283 125 284 126  0 t = 3
rlabel pdiffusion 286 125 287 126  0 t = 4
rlabel pdiffusion 282 120 288 126 0 cell no = 131
<< m1 >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< m2 >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< m2c >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 132
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 211 156 212 157  0 t = 1
rlabel pdiffusion 214 156 215 157  0 t = 2
rlabel pdiffusion 211 161 212 162  0 t = 3
rlabel pdiffusion 214 161 215 162  0 t = 4
rlabel pdiffusion 210 156 216 162 0 cell no = 133
<< m1 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2c >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< labels >>
rlabel pdiffusion 211 30 212 31  0 t = 1
rlabel pdiffusion 214 30 215 31  0 t = 2
rlabel pdiffusion 211 35 212 36  0 t = 3
rlabel pdiffusion 214 35 215 36  0 t = 4
rlabel pdiffusion 210 30 216 36 0 cell no = 134
<< m1 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2c >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 135
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 157 66 158 67  0 t = 1
rlabel pdiffusion 160 66 161 67  0 t = 2
rlabel pdiffusion 157 71 158 72  0 t = 3
rlabel pdiffusion 160 71 161 72  0 t = 4
rlabel pdiffusion 156 66 162 72 0 cell no = 136
<< m1 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2c >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< labels >>
rlabel pdiffusion 31 318 32 319  0 t = 1
rlabel pdiffusion 34 318 35 319  0 t = 2
rlabel pdiffusion 31 323 32 324  0 t = 3
rlabel pdiffusion 34 323 35 324  0 t = 4
rlabel pdiffusion 30 318 36 324 0 cell no = 137
<< m1 >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< m2 >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< m2c >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 138
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 265 12 266 13  0 t = 1
rlabel pdiffusion 268 12 269 13  0 t = 2
rlabel pdiffusion 265 17 266 18  0 t = 3
rlabel pdiffusion 268 17 269 18  0 t = 4
rlabel pdiffusion 264 12 270 18 0 cell no = 139
<< m1 >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< m2 >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< m2c >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< labels >>
rlabel pdiffusion 85 174 86 175  0 t = 1
rlabel pdiffusion 88 174 89 175  0 t = 2
rlabel pdiffusion 85 179 86 180  0 t = 3
rlabel pdiffusion 88 179 89 180  0 t = 4
rlabel pdiffusion 84 174 90 180 0 cell no = 140
<< m1 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2c >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< labels >>
rlabel pdiffusion 13 318 14 319  0 t = 1
rlabel pdiffusion 16 318 17 319  0 t = 2
rlabel pdiffusion 13 323 14 324  0 t = 3
rlabel pdiffusion 16 323 17 324  0 t = 4
rlabel pdiffusion 12 318 18 324 0 cell no = 141
<< m1 >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< m2 >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< m2c >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< labels >>
rlabel pdiffusion 247 66 248 67  0 t = 1
rlabel pdiffusion 250 66 251 67  0 t = 2
rlabel pdiffusion 247 71 248 72  0 t = 3
rlabel pdiffusion 250 71 251 72  0 t = 4
rlabel pdiffusion 246 66 252 72 0 cell no = 142
<< m1 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2c >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< labels >>
rlabel pdiffusion 175 336 176 337  0 t = 1
rlabel pdiffusion 178 336 179 337  0 t = 2
rlabel pdiffusion 175 341 176 342  0 t = 3
rlabel pdiffusion 178 341 179 342  0 t = 4
rlabel pdiffusion 174 336 180 342 0 cell no = 143
<< m1 >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< m2 >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< m2c >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< labels >>
rlabel pdiffusion 193 156 194 157  0 t = 1
rlabel pdiffusion 196 156 197 157  0 t = 2
rlabel pdiffusion 193 161 194 162  0 t = 3
rlabel pdiffusion 196 161 197 162  0 t = 4
rlabel pdiffusion 192 156 198 162 0 cell no = 144
<< m1 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2c >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< labels >>
rlabel pdiffusion 229 66 230 67  0 t = 1
rlabel pdiffusion 232 66 233 67  0 t = 2
rlabel pdiffusion 229 71 230 72  0 t = 3
rlabel pdiffusion 232 71 233 72  0 t = 4
rlabel pdiffusion 228 66 234 72 0 cell no = 145
<< m1 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2c >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< labels >>
rlabel pdiffusion 49 210 50 211  0 t = 1
rlabel pdiffusion 52 210 53 211  0 t = 2
rlabel pdiffusion 49 215 50 216  0 t = 3
rlabel pdiffusion 52 215 53 216  0 t = 4
rlabel pdiffusion 48 210 54 216 0 cell no = 146
<< m1 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2c >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< labels >>
rlabel pdiffusion 337 66 338 67  0 t = 1
rlabel pdiffusion 340 66 341 67  0 t = 2
rlabel pdiffusion 337 71 338 72  0 t = 3
rlabel pdiffusion 340 71 341 72  0 t = 4
rlabel pdiffusion 336 66 342 72 0 cell no = 147
<< m1 >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< m2 >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< m2c >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< labels >>
rlabel pdiffusion 265 66 266 67  0 t = 1
rlabel pdiffusion 268 66 269 67  0 t = 2
rlabel pdiffusion 265 71 266 72  0 t = 3
rlabel pdiffusion 268 71 269 72  0 t = 4
rlabel pdiffusion 264 66 270 72 0 cell no = 148
<< m1 >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< m2 >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< m2c >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< labels >>
rlabel pdiffusion 283 192 284 193  0 t = 1
rlabel pdiffusion 286 192 287 193  0 t = 2
rlabel pdiffusion 283 197 284 198  0 t = 3
rlabel pdiffusion 286 197 287 198  0 t = 4
rlabel pdiffusion 282 192 288 198 0 cell no = 149
<< m1 >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< m2 >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< m2c >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< labels >>
rlabel pdiffusion 175 66 176 67  0 t = 1
rlabel pdiffusion 178 66 179 67  0 t = 2
rlabel pdiffusion 175 71 176 72  0 t = 3
rlabel pdiffusion 178 71 179 72  0 t = 4
rlabel pdiffusion 174 66 180 72 0 cell no = 150
<< m1 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2c >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< labels >>
rlabel pdiffusion 301 84 302 85  0 t = 1
rlabel pdiffusion 304 84 305 85  0 t = 2
rlabel pdiffusion 301 89 302 90  0 t = 3
rlabel pdiffusion 304 89 305 90  0 t = 4
rlabel pdiffusion 300 84 306 90 0 cell no = 151
<< m1 >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< m2 >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< m2c >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 152
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 265 102 266 103  0 t = 1
rlabel pdiffusion 268 102 269 103  0 t = 2
rlabel pdiffusion 265 107 266 108  0 t = 3
rlabel pdiffusion 268 107 269 108  0 t = 4
rlabel pdiffusion 264 102 270 108 0 cell no = 153
<< m1 >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< m2 >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< m2c >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< labels >>
rlabel pdiffusion 175 300 176 301  0 t = 1
rlabel pdiffusion 178 300 179 301  0 t = 2
rlabel pdiffusion 175 305 176 306  0 t = 3
rlabel pdiffusion 178 305 179 306  0 t = 4
rlabel pdiffusion 174 300 180 306 0 cell no = 154
<< m1 >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< m2 >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< m2c >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 155
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 31 138 32 139  0 t = 1
rlabel pdiffusion 34 138 35 139  0 t = 2
rlabel pdiffusion 31 143 32 144  0 t = 3
rlabel pdiffusion 34 143 35 144  0 t = 4
rlabel pdiffusion 30 138 36 144 0 cell no = 156
<< m1 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2c >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< labels >>
rlabel pdiffusion 157 102 158 103  0 t = 1
rlabel pdiffusion 160 102 161 103  0 t = 2
rlabel pdiffusion 157 107 158 108  0 t = 3
rlabel pdiffusion 160 107 161 108  0 t = 4
rlabel pdiffusion 156 102 162 108 0 cell no = 157
<< m1 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2c >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< labels >>
rlabel pdiffusion 49 120 50 121  0 t = 1
rlabel pdiffusion 52 120 53 121  0 t = 2
rlabel pdiffusion 49 125 50 126  0 t = 3
rlabel pdiffusion 52 125 53 126  0 t = 4
rlabel pdiffusion 48 120 54 126 0 cell no = 158
<< m1 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2c >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< labels >>
rlabel pdiffusion 139 192 140 193  0 t = 1
rlabel pdiffusion 142 192 143 193  0 t = 2
rlabel pdiffusion 139 197 140 198  0 t = 3
rlabel pdiffusion 142 197 143 198  0 t = 4
rlabel pdiffusion 138 192 144 198 0 cell no = 159
<< m1 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2c >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< labels >>
rlabel pdiffusion 211 138 212 139  0 t = 1
rlabel pdiffusion 214 138 215 139  0 t = 2
rlabel pdiffusion 211 143 212 144  0 t = 3
rlabel pdiffusion 214 143 215 144  0 t = 4
rlabel pdiffusion 210 138 216 144 0 cell no = 160
<< m1 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2c >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< labels >>
rlabel pdiffusion 13 210 14 211  0 t = 1
rlabel pdiffusion 16 210 17 211  0 t = 2
rlabel pdiffusion 13 215 14 216  0 t = 3
rlabel pdiffusion 16 215 17 216  0 t = 4
rlabel pdiffusion 12 210 18 216 0 cell no = 161
<< m1 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2c >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< labels >>
rlabel pdiffusion 337 174 338 175  0 t = 1
rlabel pdiffusion 340 174 341 175  0 t = 2
rlabel pdiffusion 337 179 338 180  0 t = 3
rlabel pdiffusion 340 179 341 180  0 t = 4
rlabel pdiffusion 336 174 342 180 0 cell no = 162
<< m1 >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< m2 >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< m2c >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< labels >>
rlabel pdiffusion 211 318 212 319  0 t = 1
rlabel pdiffusion 214 318 215 319  0 t = 2
rlabel pdiffusion 211 323 212 324  0 t = 3
rlabel pdiffusion 214 323 215 324  0 t = 4
rlabel pdiffusion 210 318 216 324 0 cell no = 163
<< m1 >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< m2 >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< m2c >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< labels >>
rlabel pdiffusion 211 192 212 193  0 t = 1
rlabel pdiffusion 214 192 215 193  0 t = 2
rlabel pdiffusion 211 197 212 198  0 t = 3
rlabel pdiffusion 214 197 215 198  0 t = 4
rlabel pdiffusion 210 192 216 198 0 cell no = 164
<< m1 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2c >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< labels >>
rlabel pdiffusion 31 336 32 337  0 t = 1
rlabel pdiffusion 34 336 35 337  0 t = 2
rlabel pdiffusion 31 341 32 342  0 t = 3
rlabel pdiffusion 34 341 35 342  0 t = 4
rlabel pdiffusion 30 336 36 342 0 cell no = 165
<< m1 >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< m2 >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< m2c >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< labels >>
rlabel pdiffusion 319 246 320 247  0 t = 1
rlabel pdiffusion 322 246 323 247  0 t = 2
rlabel pdiffusion 319 251 320 252  0 t = 3
rlabel pdiffusion 322 251 323 252  0 t = 4
rlabel pdiffusion 318 246 324 252 0 cell no = 166
<< m1 >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< m2 >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< m2c >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< labels >>
rlabel pdiffusion 139 228 140 229  0 t = 1
rlabel pdiffusion 142 228 143 229  0 t = 2
rlabel pdiffusion 139 233 140 234  0 t = 3
rlabel pdiffusion 142 233 143 234  0 t = 4
rlabel pdiffusion 138 228 144 234 0 cell no = 167
<< m1 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2c >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< labels >>
rlabel pdiffusion 103 264 104 265  0 t = 1
rlabel pdiffusion 106 264 107 265  0 t = 2
rlabel pdiffusion 103 269 104 270  0 t = 3
rlabel pdiffusion 106 269 107 270  0 t = 4
rlabel pdiffusion 102 264 108 270 0 cell no = 168
<< m1 >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< m2 >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< m2c >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< labels >>
rlabel pdiffusion 139 336 140 337  0 t = 1
rlabel pdiffusion 142 336 143 337  0 t = 2
rlabel pdiffusion 139 341 140 342  0 t = 3
rlabel pdiffusion 142 341 143 342  0 t = 4
rlabel pdiffusion 138 336 144 342 0 cell no = 169
<< m1 >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< m2 >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< m2c >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 170
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 13 138 14 139  0 t = 1
rlabel pdiffusion 16 138 17 139  0 t = 2
rlabel pdiffusion 13 143 14 144  0 t = 3
rlabel pdiffusion 16 143 17 144  0 t = 4
rlabel pdiffusion 12 138 18 144 0 cell no = 171
<< m1 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2c >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< labels >>
rlabel pdiffusion 67 318 68 319  0 t = 1
rlabel pdiffusion 70 318 71 319  0 t = 2
rlabel pdiffusion 67 323 68 324  0 t = 3
rlabel pdiffusion 70 323 71 324  0 t = 4
rlabel pdiffusion 66 318 72 324 0 cell no = 172
<< m1 >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< m2 >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< m2c >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< labels >>
rlabel pdiffusion 175 210 176 211  0 t = 1
rlabel pdiffusion 178 210 179 211  0 t = 2
rlabel pdiffusion 175 215 176 216  0 t = 3
rlabel pdiffusion 178 215 179 216  0 t = 4
rlabel pdiffusion 174 210 180 216 0 cell no = 173
<< m1 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2c >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< labels >>
rlabel pdiffusion 229 30 230 31  0 t = 1
rlabel pdiffusion 232 30 233 31  0 t = 2
rlabel pdiffusion 229 35 230 36  0 t = 3
rlabel pdiffusion 232 35 233 36  0 t = 4
rlabel pdiffusion 228 30 234 36 0 cell no = 174
<< m1 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2c >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< labels >>
rlabel pdiffusion 283 282 284 283  0 t = 1
rlabel pdiffusion 286 282 287 283  0 t = 2
rlabel pdiffusion 283 287 284 288  0 t = 3
rlabel pdiffusion 286 287 287 288  0 t = 4
rlabel pdiffusion 282 282 288 288 0 cell no = 175
<< m1 >>
rect 283 282 284 283 
rect 286 282 287 283 
rect 283 287 284 288 
rect 286 287 287 288 
<< m2 >>
rect 283 282 284 283 
rect 286 282 287 283 
rect 283 287 284 288 
rect 286 287 287 288 
<< m2c >>
rect 283 282 284 283 
rect 286 282 287 283 
rect 283 287 284 288 
rect 286 287 287 288 
<< labels >>
rlabel pdiffusion 301 12 302 13  0 t = 1
rlabel pdiffusion 304 12 305 13  0 t = 2
rlabel pdiffusion 301 17 302 18  0 t = 3
rlabel pdiffusion 304 17 305 18  0 t = 4
rlabel pdiffusion 300 12 306 18 0 cell no = 176
<< m1 >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< m2 >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< m2c >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< labels >>
rlabel pdiffusion 103 174 104 175  0 t = 1
rlabel pdiffusion 106 174 107 175  0 t = 2
rlabel pdiffusion 103 179 104 180  0 t = 3
rlabel pdiffusion 106 179 107 180  0 t = 4
rlabel pdiffusion 102 174 108 180 0 cell no = 177
<< m1 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2c >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 178
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 31 264 32 265  0 t = 1
rlabel pdiffusion 34 264 35 265  0 t = 2
rlabel pdiffusion 31 269 32 270  0 t = 3
rlabel pdiffusion 34 269 35 270  0 t = 4
rlabel pdiffusion 30 264 36 270 0 cell no = 179
<< m1 >>
rect 31 264 32 265 
rect 34 264 35 265 
rect 31 269 32 270 
rect 34 269 35 270 
<< m2 >>
rect 31 264 32 265 
rect 34 264 35 265 
rect 31 269 32 270 
rect 34 269 35 270 
<< m2c >>
rect 31 264 32 265 
rect 34 264 35 265 
rect 31 269 32 270 
rect 34 269 35 270 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 180
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 49 246 50 247  0 t = 1
rlabel pdiffusion 52 246 53 247  0 t = 2
rlabel pdiffusion 49 251 50 252  0 t = 3
rlabel pdiffusion 52 251 53 252  0 t = 4
rlabel pdiffusion 48 246 54 252 0 cell no = 181
<< m1 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2c >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< labels >>
rlabel pdiffusion 229 210 230 211  0 t = 1
rlabel pdiffusion 232 210 233 211  0 t = 2
rlabel pdiffusion 229 215 230 216  0 t = 3
rlabel pdiffusion 232 215 233 216  0 t = 4
rlabel pdiffusion 228 210 234 216 0 cell no = 182
<< m1 >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< m2 >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< m2c >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< labels >>
rlabel pdiffusion 85 156 86 157  0 t = 1
rlabel pdiffusion 88 156 89 157  0 t = 2
rlabel pdiffusion 85 161 86 162  0 t = 3
rlabel pdiffusion 88 161 89 162  0 t = 4
rlabel pdiffusion 84 156 90 162 0 cell no = 183
<< m1 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2c >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< labels >>
rlabel pdiffusion 85 210 86 211  0 t = 1
rlabel pdiffusion 88 210 89 211  0 t = 2
rlabel pdiffusion 85 215 86 216  0 t = 3
rlabel pdiffusion 88 215 89 216  0 t = 4
rlabel pdiffusion 84 210 90 216 0 cell no = 184
<< m1 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2c >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 185
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 139 156 140 157  0 t = 1
rlabel pdiffusion 142 156 143 157  0 t = 2
rlabel pdiffusion 139 161 140 162  0 t = 3
rlabel pdiffusion 142 161 143 162  0 t = 4
rlabel pdiffusion 138 156 144 162 0 cell no = 186
<< m1 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2c >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< labels >>
rlabel pdiffusion 175 282 176 283  0 t = 1
rlabel pdiffusion 178 282 179 283  0 t = 2
rlabel pdiffusion 175 287 176 288  0 t = 3
rlabel pdiffusion 178 287 179 288  0 t = 4
rlabel pdiffusion 174 282 180 288 0 cell no = 187
<< m1 >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< m2 >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< m2c >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 188
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 189
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 139 12 140 13  0 t = 1
rlabel pdiffusion 142 12 143 13  0 t = 2
rlabel pdiffusion 139 17 140 18  0 t = 3
rlabel pdiffusion 142 17 143 18  0 t = 4
rlabel pdiffusion 138 12 144 18 0 cell no = 190
<< m1 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2c >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< labels >>
rlabel pdiffusion 121 336 122 337  0 t = 1
rlabel pdiffusion 124 336 125 337  0 t = 2
rlabel pdiffusion 121 341 122 342  0 t = 3
rlabel pdiffusion 124 341 125 342  0 t = 4
rlabel pdiffusion 120 336 126 342 0 cell no = 191
<< m1 >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< m2 >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< m2c >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< labels >>
rlabel pdiffusion 337 138 338 139  0 t = 1
rlabel pdiffusion 340 138 341 139  0 t = 2
rlabel pdiffusion 337 143 338 144  0 t = 3
rlabel pdiffusion 340 143 341 144  0 t = 4
rlabel pdiffusion 336 138 342 144 0 cell no = 192
<< m1 >>
rect 337 138 338 139 
rect 340 138 341 139 
rect 337 143 338 144 
rect 340 143 341 144 
<< m2 >>
rect 337 138 338 139 
rect 340 138 341 139 
rect 337 143 338 144 
rect 340 143 341 144 
<< m2c >>
rect 337 138 338 139 
rect 340 138 341 139 
rect 337 143 338 144 
rect 340 143 341 144 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 193
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 193 228 194 229  0 t = 1
rlabel pdiffusion 196 228 197 229  0 t = 2
rlabel pdiffusion 193 233 194 234  0 t = 3
rlabel pdiffusion 196 233 197 234  0 t = 4
rlabel pdiffusion 192 228 198 234 0 cell no = 194
<< m1 >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< m2 >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< m2c >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< labels >>
rlabel pdiffusion 247 102 248 103  0 t = 1
rlabel pdiffusion 250 102 251 103  0 t = 2
rlabel pdiffusion 247 107 248 108  0 t = 3
rlabel pdiffusion 250 107 251 108  0 t = 4
rlabel pdiffusion 246 102 252 108 0 cell no = 195
<< m1 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2c >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< labels >>
rlabel pdiffusion 157 12 158 13  0 t = 1
rlabel pdiffusion 160 12 161 13  0 t = 2
rlabel pdiffusion 157 17 158 18  0 t = 3
rlabel pdiffusion 160 17 161 18  0 t = 4
rlabel pdiffusion 156 12 162 18 0 cell no = 196
<< m1 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2c >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< labels >>
rlabel pdiffusion 67 120 68 121  0 t = 1
rlabel pdiffusion 70 120 71 121  0 t = 2
rlabel pdiffusion 67 125 68 126  0 t = 3
rlabel pdiffusion 70 125 71 126  0 t = 4
rlabel pdiffusion 66 120 72 126 0 cell no = 197
<< m1 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2c >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< labels >>
rlabel pdiffusion 13 336 14 337  0 t = 1
rlabel pdiffusion 16 336 17 337  0 t = 2
rlabel pdiffusion 13 341 14 342  0 t = 3
rlabel pdiffusion 16 341 17 342  0 t = 4
rlabel pdiffusion 12 336 18 342 0 cell no = 198
<< m1 >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< m2 >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< m2c >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< labels >>
rlabel pdiffusion 247 210 248 211  0 t = 1
rlabel pdiffusion 250 210 251 211  0 t = 2
rlabel pdiffusion 247 215 248 216  0 t = 3
rlabel pdiffusion 250 215 251 216  0 t = 4
rlabel pdiffusion 246 210 252 216 0 cell no = 199
<< m1 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2c >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< labels >>
rlabel pdiffusion 157 138 158 139  0 t = 1
rlabel pdiffusion 160 138 161 139  0 t = 2
rlabel pdiffusion 157 143 158 144  0 t = 3
rlabel pdiffusion 160 143 161 144  0 t = 4
rlabel pdiffusion 156 138 162 144 0 cell no = 200
<< m1 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2c >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< labels >>
rlabel pdiffusion 265 336 266 337  0 t = 1
rlabel pdiffusion 268 336 269 337  0 t = 2
rlabel pdiffusion 265 341 266 342  0 t = 3
rlabel pdiffusion 268 341 269 342  0 t = 4
rlabel pdiffusion 264 336 270 342 0 cell no = 201
<< m1 >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< m2 >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< m2c >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< labels >>
rlabel pdiffusion 337 192 338 193  0 t = 1
rlabel pdiffusion 340 192 341 193  0 t = 2
rlabel pdiffusion 337 197 338 198  0 t = 3
rlabel pdiffusion 340 197 341 198  0 t = 4
rlabel pdiffusion 336 192 342 198 0 cell no = 202
<< m1 >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< m2 >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< m2c >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< labels >>
rlabel pdiffusion 157 120 158 121  0 t = 1
rlabel pdiffusion 160 120 161 121  0 t = 2
rlabel pdiffusion 157 125 158 126  0 t = 3
rlabel pdiffusion 160 125 161 126  0 t = 4
rlabel pdiffusion 156 120 162 126 0 cell no = 203
<< m1 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2c >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< labels >>
rlabel pdiffusion 265 84 266 85  0 t = 1
rlabel pdiffusion 268 84 269 85  0 t = 2
rlabel pdiffusion 265 89 266 90  0 t = 3
rlabel pdiffusion 268 89 269 90  0 t = 4
rlabel pdiffusion 264 84 270 90 0 cell no = 204
<< m1 >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< m2 >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< m2c >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< labels >>
rlabel pdiffusion 301 192 302 193  0 t = 1
rlabel pdiffusion 304 192 305 193  0 t = 2
rlabel pdiffusion 301 197 302 198  0 t = 3
rlabel pdiffusion 304 197 305 198  0 t = 4
rlabel pdiffusion 300 192 306 198 0 cell no = 205
<< m1 >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< m2 >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< m2c >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< labels >>
rlabel pdiffusion 175 84 176 85  0 t = 1
rlabel pdiffusion 178 84 179 85  0 t = 2
rlabel pdiffusion 175 89 176 90  0 t = 3
rlabel pdiffusion 178 89 179 90  0 t = 4
rlabel pdiffusion 174 84 180 90 0 cell no = 206
<< m1 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2c >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< labels >>
rlabel pdiffusion 301 120 302 121  0 t = 1
rlabel pdiffusion 304 120 305 121  0 t = 2
rlabel pdiffusion 301 125 302 126  0 t = 3
rlabel pdiffusion 304 125 305 126  0 t = 4
rlabel pdiffusion 300 120 306 126 0 cell no = 207
<< m1 >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< m2 >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< m2c >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< labels >>
rlabel pdiffusion 31 174 32 175  0 t = 1
rlabel pdiffusion 34 174 35 175  0 t = 2
rlabel pdiffusion 31 179 32 180  0 t = 3
rlabel pdiffusion 34 179 35 180  0 t = 4
rlabel pdiffusion 30 174 36 180 0 cell no = 208
<< m1 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2c >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< labels >>
rlabel pdiffusion 247 246 248 247  0 t = 1
rlabel pdiffusion 250 246 251 247  0 t = 2
rlabel pdiffusion 247 251 248 252  0 t = 3
rlabel pdiffusion 250 251 251 252  0 t = 4
rlabel pdiffusion 246 246 252 252 0 cell no = 209
<< m1 >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< m2 >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< m2c >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< labels >>
rlabel pdiffusion 175 138 176 139  0 t = 1
rlabel pdiffusion 178 138 179 139  0 t = 2
rlabel pdiffusion 175 143 176 144  0 t = 3
rlabel pdiffusion 178 143 179 144  0 t = 4
rlabel pdiffusion 174 138 180 144 0 cell no = 210
<< m1 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2c >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< labels >>
rlabel pdiffusion 121 174 122 175  0 t = 1
rlabel pdiffusion 124 174 125 175  0 t = 2
rlabel pdiffusion 121 179 122 180  0 t = 3
rlabel pdiffusion 124 179 125 180  0 t = 4
rlabel pdiffusion 120 174 126 180 0 cell no = 211
<< m1 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2c >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< labels >>
rlabel pdiffusion 13 300 14 301  0 t = 1
rlabel pdiffusion 16 300 17 301  0 t = 2
rlabel pdiffusion 13 305 14 306  0 t = 3
rlabel pdiffusion 16 305 17 306  0 t = 4
rlabel pdiffusion 12 300 18 306 0 cell no = 212
<< m1 >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< m2 >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< m2c >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< labels >>
rlabel pdiffusion 319 156 320 157  0 t = 1
rlabel pdiffusion 322 156 323 157  0 t = 2
rlabel pdiffusion 319 161 320 162  0 t = 3
rlabel pdiffusion 322 161 323 162  0 t = 4
rlabel pdiffusion 318 156 324 162 0 cell no = 213
<< m1 >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< m2 >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< m2c >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< labels >>
rlabel pdiffusion 121 102 122 103  0 t = 1
rlabel pdiffusion 124 102 125 103  0 t = 2
rlabel pdiffusion 121 107 122 108  0 t = 3
rlabel pdiffusion 124 107 125 108  0 t = 4
rlabel pdiffusion 120 102 126 108 0 cell no = 214
<< m1 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2c >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< labels >>
rlabel pdiffusion 49 264 50 265  0 t = 1
rlabel pdiffusion 52 264 53 265  0 t = 2
rlabel pdiffusion 49 269 50 270  0 t = 3
rlabel pdiffusion 52 269 53 270  0 t = 4
rlabel pdiffusion 48 264 54 270 0 cell no = 215
<< m1 >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< m2 >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< m2c >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< labels >>
rlabel pdiffusion 157 318 158 319  0 t = 1
rlabel pdiffusion 160 318 161 319  0 t = 2
rlabel pdiffusion 157 323 158 324  0 t = 3
rlabel pdiffusion 160 323 161 324  0 t = 4
rlabel pdiffusion 156 318 162 324 0 cell no = 216
<< m1 >>
rect 157 318 158 319 
rect 160 318 161 319 
rect 157 323 158 324 
rect 160 323 161 324 
<< m2 >>
rect 157 318 158 319 
rect 160 318 161 319 
rect 157 323 158 324 
rect 160 323 161 324 
<< m2c >>
rect 157 318 158 319 
rect 160 318 161 319 
rect 157 323 158 324 
rect 160 323 161 324 
<< labels >>
rlabel pdiffusion 193 66 194 67  0 t = 1
rlabel pdiffusion 196 66 197 67  0 t = 2
rlabel pdiffusion 193 71 194 72  0 t = 3
rlabel pdiffusion 196 71 197 72  0 t = 4
rlabel pdiffusion 192 66 198 72 0 cell no = 217
<< m1 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2c >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< labels >>
rlabel pdiffusion 139 210 140 211  0 t = 1
rlabel pdiffusion 142 210 143 211  0 t = 2
rlabel pdiffusion 139 215 140 216  0 t = 3
rlabel pdiffusion 142 215 143 216  0 t = 4
rlabel pdiffusion 138 210 144 216 0 cell no = 218
<< m1 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2c >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< labels >>
rlabel pdiffusion 67 336 68 337  0 t = 1
rlabel pdiffusion 70 336 71 337  0 t = 2
rlabel pdiffusion 67 341 68 342  0 t = 3
rlabel pdiffusion 70 341 71 342  0 t = 4
rlabel pdiffusion 66 336 72 342 0 cell no = 219
<< m1 >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< m2 >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< m2c >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< labels >>
rlabel pdiffusion 193 138 194 139  0 t = 1
rlabel pdiffusion 196 138 197 139  0 t = 2
rlabel pdiffusion 193 143 194 144  0 t = 3
rlabel pdiffusion 196 143 197 144  0 t = 4
rlabel pdiffusion 192 138 198 144 0 cell no = 220
<< m1 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2c >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< labels >>
rlabel pdiffusion 283 102 284 103  0 t = 1
rlabel pdiffusion 286 102 287 103  0 t = 2
rlabel pdiffusion 283 107 284 108  0 t = 3
rlabel pdiffusion 286 107 287 108  0 t = 4
rlabel pdiffusion 282 102 288 108 0 cell no = 221
<< m1 >>
rect 283 102 284 103 
rect 286 102 287 103 
rect 283 107 284 108 
rect 286 107 287 108 
<< m2 >>
rect 283 102 284 103 
rect 286 102 287 103 
rect 283 107 284 108 
rect 286 107 287 108 
<< m2c >>
rect 283 102 284 103 
rect 286 102 287 103 
rect 283 107 284 108 
rect 286 107 287 108 
<< labels >>
rlabel pdiffusion 283 48 284 49  0 t = 1
rlabel pdiffusion 286 48 287 49  0 t = 2
rlabel pdiffusion 283 53 284 54  0 t = 3
rlabel pdiffusion 286 53 287 54  0 t = 4
rlabel pdiffusion 282 48 288 54 0 cell no = 222
<< m1 >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< m2 >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< m2c >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< labels >>
rlabel pdiffusion 337 30 338 31  0 t = 1
rlabel pdiffusion 340 30 341 31  0 t = 2
rlabel pdiffusion 337 35 338 36  0 t = 3
rlabel pdiffusion 340 35 341 36  0 t = 4
rlabel pdiffusion 336 30 342 36 0 cell no = 223
<< m1 >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< m2 >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< m2c >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< labels >>
rlabel pdiffusion 247 48 248 49  0 t = 1
rlabel pdiffusion 250 48 251 49  0 t = 2
rlabel pdiffusion 247 53 248 54  0 t = 3
rlabel pdiffusion 250 53 251 54  0 t = 4
rlabel pdiffusion 246 48 252 54 0 cell no = 224
<< m1 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2c >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< labels >>
rlabel pdiffusion 85 246 86 247  0 t = 1
rlabel pdiffusion 88 246 89 247  0 t = 2
rlabel pdiffusion 85 251 86 252  0 t = 3
rlabel pdiffusion 88 251 89 252  0 t = 4
rlabel pdiffusion 84 246 90 252 0 cell no = 225
<< m1 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2c >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< labels >>
rlabel pdiffusion 193 48 194 49  0 t = 1
rlabel pdiffusion 196 48 197 49  0 t = 2
rlabel pdiffusion 193 53 194 54  0 t = 3
rlabel pdiffusion 196 53 197 54  0 t = 4
rlabel pdiffusion 192 48 198 54 0 cell no = 226
<< m1 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2c >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< labels >>
rlabel pdiffusion 67 30 68 31  0 t = 1
rlabel pdiffusion 70 30 71 31  0 t = 2
rlabel pdiffusion 67 35 68 36  0 t = 3
rlabel pdiffusion 70 35 71 36  0 t = 4
rlabel pdiffusion 66 30 72 36 0 cell no = 227
<< m1 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2c >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< labels >>
rlabel pdiffusion 157 300 158 301  0 t = 1
rlabel pdiffusion 160 300 161 301  0 t = 2
rlabel pdiffusion 157 305 158 306  0 t = 3
rlabel pdiffusion 160 305 161 306  0 t = 4
rlabel pdiffusion 156 300 162 306 0 cell no = 228
<< m1 >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< m2 >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< m2c >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< labels >>
rlabel pdiffusion 49 228 50 229  0 t = 1
rlabel pdiffusion 52 228 53 229  0 t = 2
rlabel pdiffusion 49 233 50 234  0 t = 3
rlabel pdiffusion 52 233 53 234  0 t = 4
rlabel pdiffusion 48 228 54 234 0 cell no = 229
<< m1 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2c >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< labels >>
rlabel pdiffusion 85 192 86 193  0 t = 1
rlabel pdiffusion 88 192 89 193  0 t = 2
rlabel pdiffusion 85 197 86 198  0 t = 3
rlabel pdiffusion 88 197 89 198  0 t = 4
rlabel pdiffusion 84 192 90 198 0 cell no = 230
<< m1 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2c >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< labels >>
rlabel pdiffusion 103 246 104 247  0 t = 1
rlabel pdiffusion 106 246 107 247  0 t = 2
rlabel pdiffusion 103 251 104 252  0 t = 3
rlabel pdiffusion 106 251 107 252  0 t = 4
rlabel pdiffusion 102 246 108 252 0 cell no = 231
<< m1 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2c >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< labels >>
rlabel pdiffusion 121 282 122 283  0 t = 1
rlabel pdiffusion 124 282 125 283  0 t = 2
rlabel pdiffusion 121 287 122 288  0 t = 3
rlabel pdiffusion 124 287 125 288  0 t = 4
rlabel pdiffusion 120 282 126 288 0 cell no = 232
<< m1 >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< m2 >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< m2c >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< labels >>
rlabel pdiffusion 85 12 86 13  0 t = 1
rlabel pdiffusion 88 12 89 13  0 t = 2
rlabel pdiffusion 85 17 86 18  0 t = 3
rlabel pdiffusion 88 17 89 18  0 t = 4
rlabel pdiffusion 84 12 90 18 0 cell no = 233
<< m1 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2c >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< labels >>
rlabel pdiffusion 175 156 176 157  0 t = 1
rlabel pdiffusion 178 156 179 157  0 t = 2
rlabel pdiffusion 175 161 176 162  0 t = 3
rlabel pdiffusion 178 161 179 162  0 t = 4
rlabel pdiffusion 174 156 180 162 0 cell no = 234
<< m1 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2c >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 235
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 301 174 302 175  0 t = 1
rlabel pdiffusion 304 174 305 175  0 t = 2
rlabel pdiffusion 301 179 302 180  0 t = 3
rlabel pdiffusion 304 179 305 180  0 t = 4
rlabel pdiffusion 300 174 306 180 0 cell no = 236
<< m1 >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< m2 >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< m2c >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< labels >>
rlabel pdiffusion 49 192 50 193  0 t = 1
rlabel pdiffusion 52 192 53 193  0 t = 2
rlabel pdiffusion 49 197 50 198  0 t = 3
rlabel pdiffusion 52 197 53 198  0 t = 4
rlabel pdiffusion 48 192 54 198 0 cell no = 237
<< m1 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2c >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< labels >>
rlabel pdiffusion 337 156 338 157  0 t = 1
rlabel pdiffusion 340 156 341 157  0 t = 2
rlabel pdiffusion 337 161 338 162  0 t = 3
rlabel pdiffusion 340 161 341 162  0 t = 4
rlabel pdiffusion 336 156 342 162 0 cell no = 238
<< m1 >>
rect 337 156 338 157 
rect 340 156 341 157 
rect 337 161 338 162 
rect 340 161 341 162 
<< m2 >>
rect 337 156 338 157 
rect 340 156 341 157 
rect 337 161 338 162 
rect 340 161 341 162 
<< m2c >>
rect 337 156 338 157 
rect 340 156 341 157 
rect 337 161 338 162 
rect 340 161 341 162 
<< labels >>
rlabel pdiffusion 301 102 302 103  0 t = 1
rlabel pdiffusion 304 102 305 103  0 t = 2
rlabel pdiffusion 301 107 302 108  0 t = 3
rlabel pdiffusion 304 107 305 108  0 t = 4
rlabel pdiffusion 300 102 306 108 0 cell no = 239
<< m1 >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< m2 >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< m2c >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< labels >>
rlabel pdiffusion 247 84 248 85  0 t = 1
rlabel pdiffusion 250 84 251 85  0 t = 2
rlabel pdiffusion 247 89 248 90  0 t = 3
rlabel pdiffusion 250 89 251 90  0 t = 4
rlabel pdiffusion 246 84 252 90 0 cell no = 240
<< m1 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2c >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< labels >>
rlabel pdiffusion 193 246 194 247  0 t = 1
rlabel pdiffusion 196 246 197 247  0 t = 2
rlabel pdiffusion 193 251 194 252  0 t = 3
rlabel pdiffusion 196 251 197 252  0 t = 4
rlabel pdiffusion 192 246 198 252 0 cell no = 241
<< m1 >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< m2 >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< m2c >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< labels >>
rlabel pdiffusion 31 228 32 229  0 t = 1
rlabel pdiffusion 34 228 35 229  0 t = 2
rlabel pdiffusion 31 233 32 234  0 t = 3
rlabel pdiffusion 34 233 35 234  0 t = 4
rlabel pdiffusion 30 228 36 234 0 cell no = 242
<< m1 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2c >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< labels >>
rlabel pdiffusion 175 192 176 193  0 t = 1
rlabel pdiffusion 178 192 179 193  0 t = 2
rlabel pdiffusion 175 197 176 198  0 t = 3
rlabel pdiffusion 178 197 179 198  0 t = 4
rlabel pdiffusion 174 192 180 198 0 cell no = 243
<< m1 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2c >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< labels >>
rlabel pdiffusion 139 30 140 31  0 t = 1
rlabel pdiffusion 142 30 143 31  0 t = 2
rlabel pdiffusion 139 35 140 36  0 t = 3
rlabel pdiffusion 142 35 143 36  0 t = 4
rlabel pdiffusion 138 30 144 36 0 cell no = 244
<< m1 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2c >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< labels >>
rlabel pdiffusion 319 300 320 301  0 t = 1
rlabel pdiffusion 322 300 323 301  0 t = 2
rlabel pdiffusion 319 305 320 306  0 t = 3
rlabel pdiffusion 322 305 323 306  0 t = 4
rlabel pdiffusion 318 300 324 306 0 cell no = 245
<< m1 >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< m2 >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< m2c >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< labels >>
rlabel pdiffusion 193 120 194 121  0 t = 1
rlabel pdiffusion 196 120 197 121  0 t = 2
rlabel pdiffusion 193 125 194 126  0 t = 3
rlabel pdiffusion 196 125 197 126  0 t = 4
rlabel pdiffusion 192 120 198 126 0 cell no = 246
<< m1 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2c >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< labels >>
rlabel pdiffusion 85 138 86 139  0 t = 1
rlabel pdiffusion 88 138 89 139  0 t = 2
rlabel pdiffusion 85 143 86 144  0 t = 3
rlabel pdiffusion 88 143 89 144  0 t = 4
rlabel pdiffusion 84 138 90 144 0 cell no = 247
<< m1 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2 >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< m2c >>
rect 85 138 86 139 
rect 88 138 89 139 
rect 85 143 86 144 
rect 88 143 89 144 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 248
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 31 210 32 211  0 t = 1
rlabel pdiffusion 34 210 35 211  0 t = 2
rlabel pdiffusion 31 215 32 216  0 t = 3
rlabel pdiffusion 34 215 35 216  0 t = 4
rlabel pdiffusion 30 210 36 216 0 cell no = 249
<< m1 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2c >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< labels >>
rlabel pdiffusion 157 174 158 175  0 t = 1
rlabel pdiffusion 160 174 161 175  0 t = 2
rlabel pdiffusion 157 179 158 180  0 t = 3
rlabel pdiffusion 160 179 161 180  0 t = 4
rlabel pdiffusion 156 174 162 180 0 cell no = 250
<< m1 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2c >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< labels >>
rlabel pdiffusion 319 102 320 103  0 t = 1
rlabel pdiffusion 322 102 323 103  0 t = 2
rlabel pdiffusion 319 107 320 108  0 t = 3
rlabel pdiffusion 322 107 323 108  0 t = 4
rlabel pdiffusion 318 102 324 108 0 cell no = 251
<< m1 >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< m2 >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< m2c >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< labels >>
rlabel pdiffusion 229 246 230 247  0 t = 1
rlabel pdiffusion 232 246 233 247  0 t = 2
rlabel pdiffusion 229 251 230 252  0 t = 3
rlabel pdiffusion 232 251 233 252  0 t = 4
rlabel pdiffusion 228 246 234 252 0 cell no = 252
<< m1 >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< m2 >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< m2c >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< labels >>
rlabel pdiffusion 283 30 284 31  0 t = 1
rlabel pdiffusion 286 30 287 31  0 t = 2
rlabel pdiffusion 283 35 284 36  0 t = 3
rlabel pdiffusion 286 35 287 36  0 t = 4
rlabel pdiffusion 282 30 288 36 0 cell no = 253
<< m1 >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< m2 >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< m2c >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< labels >>
rlabel pdiffusion 13 228 14 229  0 t = 1
rlabel pdiffusion 16 228 17 229  0 t = 2
rlabel pdiffusion 13 233 14 234  0 t = 3
rlabel pdiffusion 16 233 17 234  0 t = 4
rlabel pdiffusion 12 228 18 234 0 cell no = 254
<< m1 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2c >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< labels >>
rlabel pdiffusion 337 336 338 337  0 t = 1
rlabel pdiffusion 340 336 341 337  0 t = 2
rlabel pdiffusion 337 341 338 342  0 t = 3
rlabel pdiffusion 340 341 341 342  0 t = 4
rlabel pdiffusion 336 336 342 342 0 cell no = 255
<< m1 >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< m2 >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< m2c >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< labels >>
rlabel pdiffusion 193 192 194 193  0 t = 1
rlabel pdiffusion 196 192 197 193  0 t = 2
rlabel pdiffusion 193 197 194 198  0 t = 3
rlabel pdiffusion 196 197 197 198  0 t = 4
rlabel pdiffusion 192 192 198 198 0 cell no = 256
<< m1 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2c >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< labels >>
rlabel pdiffusion 265 138 266 139  0 t = 1
rlabel pdiffusion 268 138 269 139  0 t = 2
rlabel pdiffusion 265 143 266 144  0 t = 3
rlabel pdiffusion 268 143 269 144  0 t = 4
rlabel pdiffusion 264 138 270 144 0 cell no = 257
<< m1 >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< m2 >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< m2c >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< labels >>
rlabel pdiffusion 139 264 140 265  0 t = 1
rlabel pdiffusion 142 264 143 265  0 t = 2
rlabel pdiffusion 139 269 140 270  0 t = 3
rlabel pdiffusion 142 269 143 270  0 t = 4
rlabel pdiffusion 138 264 144 270 0 cell no = 258
<< m1 >>
rect 139 264 140 265 
rect 142 264 143 265 
rect 139 269 140 270 
rect 142 269 143 270 
<< m2 >>
rect 139 264 140 265 
rect 142 264 143 265 
rect 139 269 140 270 
rect 142 269 143 270 
<< m2c >>
rect 139 264 140 265 
rect 142 264 143 265 
rect 139 269 140 270 
rect 142 269 143 270 
<< labels >>
rlabel pdiffusion 337 12 338 13  0 t = 1
rlabel pdiffusion 340 12 341 13  0 t = 2
rlabel pdiffusion 337 17 338 18  0 t = 3
rlabel pdiffusion 340 17 341 18  0 t = 4
rlabel pdiffusion 336 12 342 18 0 cell no = 259
<< m1 >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< m2 >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< m2c >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< labels >>
rlabel pdiffusion 229 300 230 301  0 t = 1
rlabel pdiffusion 232 300 233 301  0 t = 2
rlabel pdiffusion 229 305 230 306  0 t = 3
rlabel pdiffusion 232 305 233 306  0 t = 4
rlabel pdiffusion 228 300 234 306 0 cell no = 260
<< m1 >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< m2 >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< m2c >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< labels >>
rlabel pdiffusion 49 336 50 337  0 t = 1
rlabel pdiffusion 52 336 53 337  0 t = 2
rlabel pdiffusion 49 341 50 342  0 t = 3
rlabel pdiffusion 52 341 53 342  0 t = 4
rlabel pdiffusion 48 336 54 342 0 cell no = 261
<< m1 >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< m2 >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< m2c >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 262
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 157 192 158 193  0 t = 1
rlabel pdiffusion 160 192 161 193  0 t = 2
rlabel pdiffusion 157 197 158 198  0 t = 3
rlabel pdiffusion 160 197 161 198  0 t = 4
rlabel pdiffusion 156 192 162 198 0 cell no = 263
<< m1 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2c >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< labels >>
rlabel pdiffusion 265 156 266 157  0 t = 1
rlabel pdiffusion 268 156 269 157  0 t = 2
rlabel pdiffusion 265 161 266 162  0 t = 3
rlabel pdiffusion 268 161 269 162  0 t = 4
rlabel pdiffusion 264 156 270 162 0 cell no = 264
<< m1 >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< m2 >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< m2c >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< labels >>
rlabel pdiffusion 319 84 320 85  0 t = 1
rlabel pdiffusion 322 84 323 85  0 t = 2
rlabel pdiffusion 319 89 320 90  0 t = 3
rlabel pdiffusion 322 89 323 90  0 t = 4
rlabel pdiffusion 318 84 324 90 0 cell no = 265
<< m1 >>
rect 319 84 320 85 
rect 322 84 323 85 
rect 319 89 320 90 
rect 322 89 323 90 
<< m2 >>
rect 319 84 320 85 
rect 322 84 323 85 
rect 319 89 320 90 
rect 322 89 323 90 
<< m2c >>
rect 319 84 320 85 
rect 322 84 323 85 
rect 319 89 320 90 
rect 322 89 323 90 
<< labels >>
rlabel pdiffusion 283 264 284 265  0 t = 1
rlabel pdiffusion 286 264 287 265  0 t = 2
rlabel pdiffusion 283 269 284 270  0 t = 3
rlabel pdiffusion 286 269 287 270  0 t = 4
rlabel pdiffusion 282 264 288 270 0 cell no = 266
<< m1 >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< m2 >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< m2c >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< labels >>
rlabel pdiffusion 301 48 302 49  0 t = 1
rlabel pdiffusion 304 48 305 49  0 t = 2
rlabel pdiffusion 301 53 302 54  0 t = 3
rlabel pdiffusion 304 53 305 54  0 t = 4
rlabel pdiffusion 300 48 306 54 0 cell no = 267
<< m1 >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< m2 >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< m2c >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< labels >>
rlabel pdiffusion 13 192 14 193  0 t = 1
rlabel pdiffusion 16 192 17 193  0 t = 2
rlabel pdiffusion 13 197 14 198  0 t = 3
rlabel pdiffusion 16 197 17 198  0 t = 4
rlabel pdiffusion 12 192 18 198 0 cell no = 268
<< m1 >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< m2 >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< m2c >>
rect 13 192 14 193 
rect 16 192 17 193 
rect 13 197 14 198 
rect 16 197 17 198 
<< labels >>
rlabel pdiffusion 139 120 140 121  0 t = 1
rlabel pdiffusion 142 120 143 121  0 t = 2
rlabel pdiffusion 139 125 140 126  0 t = 3
rlabel pdiffusion 142 125 143 126  0 t = 4
rlabel pdiffusion 138 120 144 126 0 cell no = 269
<< m1 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2c >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< labels >>
rlabel pdiffusion 103 228 104 229  0 t = 1
rlabel pdiffusion 106 228 107 229  0 t = 2
rlabel pdiffusion 103 233 104 234  0 t = 3
rlabel pdiffusion 106 233 107 234  0 t = 4
rlabel pdiffusion 102 228 108 234 0 cell no = 270
<< m1 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2c >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< labels >>
rlabel pdiffusion 157 336 158 337  0 t = 1
rlabel pdiffusion 160 336 161 337  0 t = 2
rlabel pdiffusion 157 341 158 342  0 t = 3
rlabel pdiffusion 160 341 161 342  0 t = 4
rlabel pdiffusion 156 336 162 342 0 cell no = 271
<< m1 >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< m2 >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< m2c >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 272
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 103 30 104 31  0 t = 1
rlabel pdiffusion 106 30 107 31  0 t = 2
rlabel pdiffusion 103 35 104 36  0 t = 3
rlabel pdiffusion 106 35 107 36  0 t = 4
rlabel pdiffusion 102 30 108 36 0 cell no = 273
<< m1 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2c >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< labels >>
rlabel pdiffusion 175 120 176 121  0 t = 1
rlabel pdiffusion 178 120 179 121  0 t = 2
rlabel pdiffusion 175 125 176 126  0 t = 3
rlabel pdiffusion 178 125 179 126  0 t = 4
rlabel pdiffusion 174 120 180 126 0 cell no = 274
<< m1 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2c >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< labels >>
rlabel pdiffusion 175 102 176 103  0 t = 1
rlabel pdiffusion 178 102 179 103  0 t = 2
rlabel pdiffusion 175 107 176 108  0 t = 3
rlabel pdiffusion 178 107 179 108  0 t = 4
rlabel pdiffusion 174 102 180 108 0 cell no = 275
<< m1 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2c >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< labels >>
rlabel pdiffusion 157 228 158 229  0 t = 1
rlabel pdiffusion 160 228 161 229  0 t = 2
rlabel pdiffusion 157 233 158 234  0 t = 3
rlabel pdiffusion 160 233 161 234  0 t = 4
rlabel pdiffusion 156 228 162 234 0 cell no = 276
<< m1 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2c >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< labels >>
rlabel pdiffusion 103 210 104 211  0 t = 1
rlabel pdiffusion 106 210 107 211  0 t = 2
rlabel pdiffusion 103 215 104 216  0 t = 3
rlabel pdiffusion 106 215 107 216  0 t = 4
rlabel pdiffusion 102 210 108 216 0 cell no = 277
<< m1 >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< m2 >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< m2c >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< labels >>
rlabel pdiffusion 301 30 302 31  0 t = 1
rlabel pdiffusion 304 30 305 31  0 t = 2
rlabel pdiffusion 301 35 302 36  0 t = 3
rlabel pdiffusion 304 35 305 36  0 t = 4
rlabel pdiffusion 300 30 306 36 0 cell no = 278
<< m1 >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< m2 >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< m2c >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< labels >>
rlabel pdiffusion 247 156 248 157  0 t = 1
rlabel pdiffusion 250 156 251 157  0 t = 2
rlabel pdiffusion 247 161 248 162  0 t = 3
rlabel pdiffusion 250 161 251 162  0 t = 4
rlabel pdiffusion 246 156 252 162 0 cell no = 279
<< m1 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2c >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 280
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 265 282 266 283  0 t = 1
rlabel pdiffusion 268 282 269 283  0 t = 2
rlabel pdiffusion 265 287 266 288  0 t = 3
rlabel pdiffusion 268 287 269 288  0 t = 4
rlabel pdiffusion 264 282 270 288 0 cell no = 281
<< m1 >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< m2 >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< m2c >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< labels >>
rlabel pdiffusion 301 156 302 157  0 t = 1
rlabel pdiffusion 304 156 305 157  0 t = 2
rlabel pdiffusion 301 161 302 162  0 t = 3
rlabel pdiffusion 304 161 305 162  0 t = 4
rlabel pdiffusion 300 156 306 162 0 cell no = 282
<< m1 >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< m2 >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< m2c >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 283
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 284
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 319 264 320 265  0 t = 1
rlabel pdiffusion 322 264 323 265  0 t = 2
rlabel pdiffusion 319 269 320 270  0 t = 3
rlabel pdiffusion 322 269 323 270  0 t = 4
rlabel pdiffusion 318 264 324 270 0 cell no = 285
<< m1 >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< m2 >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< m2c >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< labels >>
rlabel pdiffusion 139 84 140 85  0 t = 1
rlabel pdiffusion 142 84 143 85  0 t = 2
rlabel pdiffusion 139 89 140 90  0 t = 3
rlabel pdiffusion 142 89 143 90  0 t = 4
rlabel pdiffusion 138 84 144 90 0 cell no = 286
<< m1 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2c >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< labels >>
rlabel pdiffusion 31 12 32 13  0 t = 1
rlabel pdiffusion 34 12 35 13  0 t = 2
rlabel pdiffusion 31 17 32 18  0 t = 3
rlabel pdiffusion 34 17 35 18  0 t = 4
rlabel pdiffusion 30 12 36 18 0 cell no = 287
<< m1 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2c >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< labels >>
rlabel pdiffusion 211 246 212 247  0 t = 1
rlabel pdiffusion 214 246 215 247  0 t = 2
rlabel pdiffusion 211 251 212 252  0 t = 3
rlabel pdiffusion 214 251 215 252  0 t = 4
rlabel pdiffusion 210 246 216 252 0 cell no = 288
<< m1 >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< m2 >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< m2c >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 289
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 337 246 338 247  0 t = 1
rlabel pdiffusion 340 246 341 247  0 t = 2
rlabel pdiffusion 337 251 338 252  0 t = 3
rlabel pdiffusion 340 251 341 252  0 t = 4
rlabel pdiffusion 336 246 342 252 0 cell no = 290
<< m1 >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< m2 >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< m2c >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< labels >>
rlabel pdiffusion 85 264 86 265  0 t = 1
rlabel pdiffusion 88 264 89 265  0 t = 2
rlabel pdiffusion 85 269 86 270  0 t = 3
rlabel pdiffusion 88 269 89 270  0 t = 4
rlabel pdiffusion 84 264 90 270 0 cell no = 291
<< m1 >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< m2 >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< m2c >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 292
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 121 156 122 157  0 t = 1
rlabel pdiffusion 124 156 125 157  0 t = 2
rlabel pdiffusion 121 161 122 162  0 t = 3
rlabel pdiffusion 124 161 125 162  0 t = 4
rlabel pdiffusion 120 156 126 162 0 cell no = 293
<< m1 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2c >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< labels >>
rlabel pdiffusion 283 300 284 301  0 t = 1
rlabel pdiffusion 286 300 287 301  0 t = 2
rlabel pdiffusion 283 305 284 306  0 t = 3
rlabel pdiffusion 286 305 287 306  0 t = 4
rlabel pdiffusion 282 300 288 306 0 cell no = 294
<< m1 >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< m2 >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< m2c >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< labels >>
rlabel pdiffusion 283 156 284 157  0 t = 1
rlabel pdiffusion 286 156 287 157  0 t = 2
rlabel pdiffusion 283 161 284 162  0 t = 3
rlabel pdiffusion 286 161 287 162  0 t = 4
rlabel pdiffusion 282 156 288 162 0 cell no = 295
<< m1 >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< m2 >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< m2c >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 296
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 103 318 104 319  0 t = 1
rlabel pdiffusion 106 318 107 319  0 t = 2
rlabel pdiffusion 103 323 104 324  0 t = 3
rlabel pdiffusion 106 323 107 324  0 t = 4
rlabel pdiffusion 102 318 108 324 0 cell no = 297
<< m1 >>
rect 103 318 104 319 
rect 106 318 107 319 
rect 103 323 104 324 
rect 106 323 107 324 
<< m2 >>
rect 103 318 104 319 
rect 106 318 107 319 
rect 103 323 104 324 
rect 106 323 107 324 
<< m2c >>
rect 103 318 104 319 
rect 106 318 107 319 
rect 103 323 104 324 
rect 106 323 107 324 
<< labels >>
rlabel pdiffusion 211 48 212 49  0 t = 1
rlabel pdiffusion 214 48 215 49  0 t = 2
rlabel pdiffusion 211 53 212 54  0 t = 3
rlabel pdiffusion 214 53 215 54  0 t = 4
rlabel pdiffusion 210 48 216 54 0 cell no = 298
<< m1 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2c >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< labels >>
rlabel pdiffusion 85 228 86 229  0 t = 1
rlabel pdiffusion 88 228 89 229  0 t = 2
rlabel pdiffusion 85 233 86 234  0 t = 3
rlabel pdiffusion 88 233 89 234  0 t = 4
rlabel pdiffusion 84 228 90 234 0 cell no = 299
<< m1 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2c >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< labels >>
rlabel pdiffusion 31 192 32 193  0 t = 1
rlabel pdiffusion 34 192 35 193  0 t = 2
rlabel pdiffusion 31 197 32 198  0 t = 3
rlabel pdiffusion 34 197 35 198  0 t = 4
rlabel pdiffusion 30 192 36 198 0 cell no = 300
<< m1 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2c >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< labels >>
rlabel pdiffusion 193 12 194 13  0 t = 1
rlabel pdiffusion 196 12 197 13  0 t = 2
rlabel pdiffusion 193 17 194 18  0 t = 3
rlabel pdiffusion 196 17 197 18  0 t = 4
rlabel pdiffusion 192 12 198 18 0 cell no = 301
<< m1 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2c >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< labels >>
rlabel pdiffusion 139 300 140 301  0 t = 1
rlabel pdiffusion 142 300 143 301  0 t = 2
rlabel pdiffusion 139 305 140 306  0 t = 3
rlabel pdiffusion 142 305 143 306  0 t = 4
rlabel pdiffusion 138 300 144 306 0 cell no = 302
<< m1 >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< m2 >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< m2c >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< labels >>
rlabel pdiffusion 121 84 122 85  0 t = 1
rlabel pdiffusion 124 84 125 85  0 t = 2
rlabel pdiffusion 121 89 122 90  0 t = 3
rlabel pdiffusion 124 89 125 90  0 t = 4
rlabel pdiffusion 120 84 126 90 0 cell no = 303
<< m1 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2c >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< labels >>
rlabel pdiffusion 103 336 104 337  0 t = 1
rlabel pdiffusion 106 336 107 337  0 t = 2
rlabel pdiffusion 103 341 104 342  0 t = 3
rlabel pdiffusion 106 341 107 342  0 t = 4
rlabel pdiffusion 102 336 108 342 0 cell no = 304
<< m1 >>
rect 103 336 104 337 
rect 106 336 107 337 
rect 103 341 104 342 
rect 106 341 107 342 
<< m2 >>
rect 103 336 104 337 
rect 106 336 107 337 
rect 103 341 104 342 
rect 106 341 107 342 
<< m2c >>
rect 103 336 104 337 
rect 106 336 107 337 
rect 103 341 104 342 
rect 106 341 107 342 
<< labels >>
rlabel pdiffusion 247 318 248 319  0 t = 1
rlabel pdiffusion 250 318 251 319  0 t = 2
rlabel pdiffusion 247 323 248 324  0 t = 3
rlabel pdiffusion 250 323 251 324  0 t = 4
rlabel pdiffusion 246 318 252 324 0 cell no = 305
<< m1 >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< m2 >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< m2c >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< labels >>
rlabel pdiffusion 229 336 230 337  0 t = 1
rlabel pdiffusion 232 336 233 337  0 t = 2
rlabel pdiffusion 229 341 230 342  0 t = 3
rlabel pdiffusion 232 341 233 342  0 t = 4
rlabel pdiffusion 228 336 234 342 0 cell no = 306
<< m1 >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< m2 >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< m2c >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< labels >>
rlabel pdiffusion 211 300 212 301  0 t = 1
rlabel pdiffusion 214 300 215 301  0 t = 2
rlabel pdiffusion 211 305 212 306  0 t = 3
rlabel pdiffusion 214 305 215 306  0 t = 4
rlabel pdiffusion 210 300 216 306 0 cell no = 307
<< m1 >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< m2 >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< m2c >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< labels >>
rlabel pdiffusion 175 246 176 247  0 t = 1
rlabel pdiffusion 178 246 179 247  0 t = 2
rlabel pdiffusion 175 251 176 252  0 t = 3
rlabel pdiffusion 178 251 179 252  0 t = 4
rlabel pdiffusion 174 246 180 252 0 cell no = 308
<< m1 >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< m2 >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< m2c >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< labels >>
rlabel pdiffusion 265 30 266 31  0 t = 1
rlabel pdiffusion 268 30 269 31  0 t = 2
rlabel pdiffusion 265 35 266 36  0 t = 3
rlabel pdiffusion 268 35 269 36  0 t = 4
rlabel pdiffusion 264 30 270 36 0 cell no = 309
<< m1 >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< m2 >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< m2c >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< labels >>
rlabel pdiffusion 103 84 104 85  0 t = 1
rlabel pdiffusion 106 84 107 85  0 t = 2
rlabel pdiffusion 103 89 104 90  0 t = 3
rlabel pdiffusion 106 89 107 90  0 t = 4
rlabel pdiffusion 102 84 108 90 0 cell no = 310
<< m1 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2c >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< labels >>
rlabel pdiffusion 319 336 320 337  0 t = 1
rlabel pdiffusion 322 336 323 337  0 t = 2
rlabel pdiffusion 319 341 320 342  0 t = 3
rlabel pdiffusion 322 341 323 342  0 t = 4
rlabel pdiffusion 318 336 324 342 0 cell no = 311
<< m1 >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< m2 >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< m2c >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< labels >>
rlabel pdiffusion 211 228 212 229  0 t = 1
rlabel pdiffusion 214 228 215 229  0 t = 2
rlabel pdiffusion 211 233 212 234  0 t = 3
rlabel pdiffusion 214 233 215 234  0 t = 4
rlabel pdiffusion 210 228 216 234 0 cell no = 312
<< m1 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2c >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< labels >>
rlabel pdiffusion 283 246 284 247  0 t = 1
rlabel pdiffusion 286 246 287 247  0 t = 2
rlabel pdiffusion 283 251 284 252  0 t = 3
rlabel pdiffusion 286 251 287 252  0 t = 4
rlabel pdiffusion 282 246 288 252 0 cell no = 313
<< m1 >>
rect 283 246 284 247 
rect 286 246 287 247 
rect 283 251 284 252 
rect 286 251 287 252 
<< m2 >>
rect 283 246 284 247 
rect 286 246 287 247 
rect 283 251 284 252 
rect 286 251 287 252 
<< m2c >>
rect 283 246 284 247 
rect 286 246 287 247 
rect 283 251 284 252 
rect 286 251 287 252 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 314
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 315
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 211 174 212 175  0 t = 1
rlabel pdiffusion 214 174 215 175  0 t = 2
rlabel pdiffusion 211 179 212 180  0 t = 3
rlabel pdiffusion 214 179 215 180  0 t = 4
rlabel pdiffusion 210 174 216 180 0 cell no = 316
<< m1 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2c >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< labels >>
rlabel pdiffusion 337 120 338 121  0 t = 1
rlabel pdiffusion 340 120 341 121  0 t = 2
rlabel pdiffusion 337 125 338 126  0 t = 3
rlabel pdiffusion 340 125 341 126  0 t = 4
rlabel pdiffusion 336 120 342 126 0 cell no = 317
<< m1 >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< m2 >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< m2c >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< labels >>
rlabel pdiffusion 265 210 266 211  0 t = 1
rlabel pdiffusion 268 210 269 211  0 t = 2
rlabel pdiffusion 265 215 266 216  0 t = 3
rlabel pdiffusion 268 215 269 216  0 t = 4
rlabel pdiffusion 264 210 270 216 0 cell no = 318
<< m1 >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< m2 >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< m2c >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< labels >>
rlabel pdiffusion 283 84 284 85  0 t = 1
rlabel pdiffusion 286 84 287 85  0 t = 2
rlabel pdiffusion 283 89 284 90  0 t = 3
rlabel pdiffusion 286 89 287 90  0 t = 4
rlabel pdiffusion 282 84 288 90 0 cell no = 319
<< m1 >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< m2 >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< m2c >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< labels >>
rlabel pdiffusion 67 174 68 175  0 t = 1
rlabel pdiffusion 70 174 71 175  0 t = 2
rlabel pdiffusion 67 179 68 180  0 t = 3
rlabel pdiffusion 70 179 71 180  0 t = 4
rlabel pdiffusion 66 174 72 180 0 cell no = 320
<< m1 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2c >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< labels >>
rlabel pdiffusion 265 264 266 265  0 t = 1
rlabel pdiffusion 268 264 269 265  0 t = 2
rlabel pdiffusion 265 269 266 270  0 t = 3
rlabel pdiffusion 268 269 269 270  0 t = 4
rlabel pdiffusion 264 264 270 270 0 cell no = 321
<< m1 >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< m2 >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< m2c >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< labels >>
rlabel pdiffusion 49 156 50 157  0 t = 1
rlabel pdiffusion 52 156 53 157  0 t = 2
rlabel pdiffusion 49 161 50 162  0 t = 3
rlabel pdiffusion 52 161 53 162  0 t = 4
rlabel pdiffusion 48 156 54 162 0 cell no = 322
<< m1 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2c >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< labels >>
rlabel pdiffusion 175 318 176 319  0 t = 1
rlabel pdiffusion 178 318 179 319  0 t = 2
rlabel pdiffusion 175 323 176 324  0 t = 3
rlabel pdiffusion 178 323 179 324  0 t = 4
rlabel pdiffusion 174 318 180 324 0 cell no = 323
<< m1 >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< m2 >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< m2c >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< labels >>
rlabel pdiffusion 319 210 320 211  0 t = 1
rlabel pdiffusion 322 210 323 211  0 t = 2
rlabel pdiffusion 319 215 320 216  0 t = 3
rlabel pdiffusion 322 215 323 216  0 t = 4
rlabel pdiffusion 318 210 324 216 0 cell no = 324
<< m1 >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< m2 >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< m2c >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< labels >>
rlabel pdiffusion 121 192 122 193  0 t = 1
rlabel pdiffusion 124 192 125 193  0 t = 2
rlabel pdiffusion 121 197 122 198  0 t = 3
rlabel pdiffusion 124 197 125 198  0 t = 4
rlabel pdiffusion 120 192 126 198 0 cell no = 325
<< m1 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2c >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< labels >>
rlabel pdiffusion 67 300 68 301  0 t = 1
rlabel pdiffusion 70 300 71 301  0 t = 2
rlabel pdiffusion 67 305 68 306  0 t = 3
rlabel pdiffusion 70 305 71 306  0 t = 4
rlabel pdiffusion 66 300 72 306 0 cell no = 326
<< m1 >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< m2 >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< m2c >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< labels >>
rlabel pdiffusion 265 228 266 229  0 t = 1
rlabel pdiffusion 268 228 269 229  0 t = 2
rlabel pdiffusion 265 233 266 234  0 t = 3
rlabel pdiffusion 268 233 269 234  0 t = 4
rlabel pdiffusion 264 228 270 234 0 cell no = 327
<< m1 >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< m2 >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< m2c >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< labels >>
rlabel pdiffusion 13 120 14 121  0 t = 1
rlabel pdiffusion 16 120 17 121  0 t = 2
rlabel pdiffusion 13 125 14 126  0 t = 3
rlabel pdiffusion 16 125 17 126  0 t = 4
rlabel pdiffusion 12 120 18 126 0 cell no = 328
<< m1 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2c >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< labels >>
rlabel pdiffusion 211 66 212 67  0 t = 1
rlabel pdiffusion 214 66 215 67  0 t = 2
rlabel pdiffusion 211 71 212 72  0 t = 3
rlabel pdiffusion 214 71 215 72  0 t = 4
rlabel pdiffusion 210 66 216 72 0 cell no = 329
<< m1 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2c >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 330
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 193 282 194 283  0 t = 1
rlabel pdiffusion 196 282 197 283  0 t = 2
rlabel pdiffusion 193 287 194 288  0 t = 3
rlabel pdiffusion 196 287 197 288  0 t = 4
rlabel pdiffusion 192 282 198 288 0 cell no = 331
<< m1 >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< m2 >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< m2c >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< labels >>
rlabel pdiffusion 139 48 140 49  0 t = 1
rlabel pdiffusion 142 48 143 49  0 t = 2
rlabel pdiffusion 139 53 140 54  0 t = 3
rlabel pdiffusion 142 53 143 54  0 t = 4
rlabel pdiffusion 138 48 144 54 0 cell no = 332
<< m1 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2c >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< labels >>
rlabel pdiffusion 229 228 230 229  0 t = 1
rlabel pdiffusion 232 228 233 229  0 t = 2
rlabel pdiffusion 229 233 230 234  0 t = 3
rlabel pdiffusion 232 233 233 234  0 t = 4
rlabel pdiffusion 228 228 234 234 0 cell no = 333
<< m1 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2c >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< labels >>
rlabel pdiffusion 103 138 104 139  0 t = 1
rlabel pdiffusion 106 138 107 139  0 t = 2
rlabel pdiffusion 103 143 104 144  0 t = 3
rlabel pdiffusion 106 143 107 144  0 t = 4
rlabel pdiffusion 102 138 108 144 0 cell no = 334
<< m1 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2c >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< labels >>
rlabel pdiffusion 265 192 266 193  0 t = 1
rlabel pdiffusion 268 192 269 193  0 t = 2
rlabel pdiffusion 265 197 266 198  0 t = 3
rlabel pdiffusion 268 197 269 198  0 t = 4
rlabel pdiffusion 264 192 270 198 0 cell no = 335
<< m1 >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< m2 >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< m2c >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< labels >>
rlabel pdiffusion 301 138 302 139  0 t = 1
rlabel pdiffusion 304 138 305 139  0 t = 2
rlabel pdiffusion 301 143 302 144  0 t = 3
rlabel pdiffusion 304 143 305 144  0 t = 4
rlabel pdiffusion 300 138 306 144 0 cell no = 336
<< m1 >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< m2 >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< m2c >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< labels >>
rlabel pdiffusion 229 174 230 175  0 t = 1
rlabel pdiffusion 232 174 233 175  0 t = 2
rlabel pdiffusion 229 179 230 180  0 t = 3
rlabel pdiffusion 232 179 233 180  0 t = 4
rlabel pdiffusion 228 174 234 180 0 cell no = 337
<< m1 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2c >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< labels >>
rlabel pdiffusion 193 336 194 337  0 t = 1
rlabel pdiffusion 196 336 197 337  0 t = 2
rlabel pdiffusion 193 341 194 342  0 t = 3
rlabel pdiffusion 196 341 197 342  0 t = 4
rlabel pdiffusion 192 336 198 342 0 cell no = 338
<< m1 >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< m2 >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< m2c >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< labels >>
rlabel pdiffusion 175 264 176 265  0 t = 1
rlabel pdiffusion 178 264 179 265  0 t = 2
rlabel pdiffusion 175 269 176 270  0 t = 3
rlabel pdiffusion 178 269 179 270  0 t = 4
rlabel pdiffusion 174 264 180 270 0 cell no = 339
<< m1 >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< m2 >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< m2c >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< labels >>
rlabel pdiffusion 247 336 248 337  0 t = 1
rlabel pdiffusion 250 336 251 337  0 t = 2
rlabel pdiffusion 247 341 248 342  0 t = 3
rlabel pdiffusion 250 341 251 342  0 t = 4
rlabel pdiffusion 246 336 252 342 0 cell no = 340
<< m1 >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< m2 >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< m2c >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< labels >>
rlabel pdiffusion 211 336 212 337  0 t = 1
rlabel pdiffusion 214 336 215 337  0 t = 2
rlabel pdiffusion 211 341 212 342  0 t = 3
rlabel pdiffusion 214 341 215 342  0 t = 4
rlabel pdiffusion 210 336 216 342 0 cell no = 341
<< m1 >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< m2 >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< m2c >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< labels >>
rlabel pdiffusion 85 318 86 319  0 t = 1
rlabel pdiffusion 88 318 89 319  0 t = 2
rlabel pdiffusion 85 323 86 324  0 t = 3
rlabel pdiffusion 88 323 89 324  0 t = 4
rlabel pdiffusion 84 318 90 324 0 cell no = 342
<< m1 >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< m2 >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< m2c >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< labels >>
rlabel pdiffusion 265 300 266 301  0 t = 1
rlabel pdiffusion 268 300 269 301  0 t = 2
rlabel pdiffusion 265 305 266 306  0 t = 3
rlabel pdiffusion 268 305 269 306  0 t = 4
rlabel pdiffusion 264 300 270 306 0 cell no = 343
<< m1 >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< m2 >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< m2c >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< labels >>
rlabel pdiffusion 319 318 320 319  0 t = 1
rlabel pdiffusion 322 318 323 319  0 t = 2
rlabel pdiffusion 319 323 320 324  0 t = 3
rlabel pdiffusion 322 323 323 324  0 t = 4
rlabel pdiffusion 318 318 324 324 0 cell no = 344
<< m1 >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< m2 >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< m2c >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< labels >>
rlabel pdiffusion 139 318 140 319  0 t = 1
rlabel pdiffusion 142 318 143 319  0 t = 2
rlabel pdiffusion 139 323 140 324  0 t = 3
rlabel pdiffusion 142 323 143 324  0 t = 4
rlabel pdiffusion 138 318 144 324 0 cell no = 345
<< m1 >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< m2 >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< m2c >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< labels >>
rlabel pdiffusion 157 156 158 157  0 t = 1
rlabel pdiffusion 160 156 161 157  0 t = 2
rlabel pdiffusion 157 161 158 162  0 t = 3
rlabel pdiffusion 160 161 161 162  0 t = 4
rlabel pdiffusion 156 156 162 162 0 cell no = 346
<< m1 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2c >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< labels >>
rlabel pdiffusion 13 174 14 175  0 t = 1
rlabel pdiffusion 16 174 17 175  0 t = 2
rlabel pdiffusion 13 179 14 180  0 t = 3
rlabel pdiffusion 16 179 17 180  0 t = 4
rlabel pdiffusion 12 174 18 180 0 cell no = 347
<< m1 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2c >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< labels >>
rlabel pdiffusion 211 264 212 265  0 t = 1
rlabel pdiffusion 214 264 215 265  0 t = 2
rlabel pdiffusion 211 269 212 270  0 t = 3
rlabel pdiffusion 214 269 215 270  0 t = 4
rlabel pdiffusion 210 264 216 270 0 cell no = 348
<< m1 >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< m2 >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< m2c >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< labels >>
rlabel pdiffusion 301 336 302 337  0 t = 1
rlabel pdiffusion 304 336 305 337  0 t = 2
rlabel pdiffusion 301 341 302 342  0 t = 3
rlabel pdiffusion 304 341 305 342  0 t = 4
rlabel pdiffusion 300 336 306 342 0 cell no = 349
<< m1 >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< m2 >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< m2c >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< labels >>
rlabel pdiffusion 193 264 194 265  0 t = 1
rlabel pdiffusion 196 264 197 265  0 t = 2
rlabel pdiffusion 193 269 194 270  0 t = 3
rlabel pdiffusion 196 269 197 270  0 t = 4
rlabel pdiffusion 192 264 198 270 0 cell no = 350
<< m1 >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< m2 >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< m2c >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< labels >>
rlabel pdiffusion 229 192 230 193  0 t = 1
rlabel pdiffusion 232 192 233 193  0 t = 2
rlabel pdiffusion 229 197 230 198  0 t = 3
rlabel pdiffusion 232 197 233 198  0 t = 4
rlabel pdiffusion 228 192 234 198 0 cell no = 351
<< m1 >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< m2 >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< m2c >>
rect 229 192 230 193 
rect 232 192 233 193 
rect 229 197 230 198 
rect 232 197 233 198 
<< labels >>
rlabel pdiffusion 247 228 248 229  0 t = 1
rlabel pdiffusion 250 228 251 229  0 t = 2
rlabel pdiffusion 247 233 248 234  0 t = 3
rlabel pdiffusion 250 233 251 234  0 t = 4
rlabel pdiffusion 246 228 252 234 0 cell no = 352
<< m1 >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< m2 >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< m2c >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< labels >>
rlabel pdiffusion 301 282 302 283  0 t = 1
rlabel pdiffusion 304 282 305 283  0 t = 2
rlabel pdiffusion 301 287 302 288  0 t = 3
rlabel pdiffusion 304 287 305 288  0 t = 4
rlabel pdiffusion 300 282 306 288 0 cell no = 353
<< m1 >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< m2 >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< m2c >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< labels >>
rlabel pdiffusion 319 192 320 193  0 t = 1
rlabel pdiffusion 322 192 323 193  0 t = 2
rlabel pdiffusion 319 197 320 198  0 t = 3
rlabel pdiffusion 322 197 323 198  0 t = 4
rlabel pdiffusion 318 192 324 198 0 cell no = 354
<< m1 >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< m2 >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< m2c >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< labels >>
rlabel pdiffusion 49 174 50 175  0 t = 1
rlabel pdiffusion 52 174 53 175  0 t = 2
rlabel pdiffusion 49 179 50 180  0 t = 3
rlabel pdiffusion 52 179 53 180  0 t = 4
rlabel pdiffusion 48 174 54 180 0 cell no = 355
<< m1 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2c >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 356
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 337 48 338 49  0 t = 1
rlabel pdiffusion 340 48 341 49  0 t = 2
rlabel pdiffusion 337 53 338 54  0 t = 3
rlabel pdiffusion 340 53 341 54  0 t = 4
rlabel pdiffusion 336 48 342 54 0 cell no = 357
<< m1 >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< m2 >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< m2c >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< labels >>
rlabel pdiffusion 319 48 320 49  0 t = 1
rlabel pdiffusion 322 48 323 49  0 t = 2
rlabel pdiffusion 319 53 320 54  0 t = 3
rlabel pdiffusion 322 53 323 54  0 t = 4
rlabel pdiffusion 318 48 324 54 0 cell no = 358
<< m1 >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< m2 >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< m2c >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 359
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 229 48 230 49  0 t = 1
rlabel pdiffusion 232 48 233 49  0 t = 2
rlabel pdiffusion 229 53 230 54  0 t = 3
rlabel pdiffusion 232 53 233 54  0 t = 4
rlabel pdiffusion 228 48 234 54 0 cell no = 360
<< m1 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2c >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< end >> 
