magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 30 7 31 8 
<< m1 >>
rect 31 7 32 8 
<< m1 >>
rect 32 7 33 8 
<< m1 >>
rect 33 7 34 8 
<< m1 >>
rect 34 7 35 8 
<< m1 >>
rect 35 7 36 8 
<< m1 >>
rect 36 7 37 8 
<< m1 >>
rect 37 7 38 8 
<< m1 >>
rect 38 7 39 8 
<< m1 >>
rect 39 7 40 8 
<< m1 >>
rect 40 7 41 8 
<< m1 >>
rect 41 7 42 8 
<< m1 >>
rect 42 7 43 8 
<< m2 >>
rect 42 7 43 8 
<< m2c >>
rect 42 7 43 8 
<< m1 >>
rect 42 7 43 8 
<< m2 >>
rect 42 7 43 8 
<< m2 >>
rect 43 7 44 8 
<< m1 >>
rect 44 7 45 8 
<< m2 >>
rect 44 7 45 8 
<< m1 >>
rect 45 7 46 8 
<< m2 >>
rect 45 7 46 8 
<< m1 >>
rect 46 7 47 8 
<< m2 >>
rect 46 7 47 8 
<< m1 >>
rect 47 7 48 8 
<< m2 >>
rect 47 7 48 8 
<< m1 >>
rect 48 7 49 8 
<< m2 >>
rect 48 7 49 8 
<< m1 >>
rect 49 7 50 8 
<< m2 >>
rect 49 7 50 8 
<< m1 >>
rect 50 7 51 8 
<< m2 >>
rect 50 7 51 8 
<< m1 >>
rect 51 7 52 8 
<< m2 >>
rect 51 7 52 8 
<< m1 >>
rect 52 7 53 8 
<< m2 >>
rect 52 7 53 8 
<< m1 >>
rect 53 7 54 8 
<< m2 >>
rect 53 7 54 8 
<< m1 >>
rect 54 7 55 8 
<< m2 >>
rect 54 7 55 8 
<< m1 >>
rect 55 7 56 8 
<< m2 >>
rect 55 7 56 8 
<< m1 >>
rect 56 7 57 8 
<< m2 >>
rect 56 7 57 8 
<< m1 >>
rect 57 7 58 8 
<< m2 >>
rect 57 7 58 8 
<< m1 >>
rect 58 7 59 8 
<< m2 >>
rect 58 7 59 8 
<< m1 >>
rect 59 7 60 8 
<< m2 >>
rect 59 7 60 8 
<< m1 >>
rect 60 7 61 8 
<< m2 >>
rect 60 7 61 8 
<< m1 >>
rect 61 7 62 8 
<< m2 >>
rect 61 7 62 8 
<< m1 >>
rect 62 7 63 8 
<< m2 >>
rect 62 7 63 8 
<< m1 >>
rect 63 7 64 8 
<< m2 >>
rect 63 7 64 8 
<< m1 >>
rect 64 7 65 8 
<< m2 >>
rect 64 7 65 8 
<< m1 >>
rect 65 7 66 8 
<< m2 >>
rect 65 7 66 8 
<< m1 >>
rect 66 7 67 8 
<< m2 >>
rect 66 7 67 8 
<< m1 >>
rect 67 7 68 8 
<< m2 >>
rect 67 7 68 8 
<< m1 >>
rect 68 7 69 8 
<< m2 >>
rect 68 7 69 8 
<< m1 >>
rect 69 7 70 8 
<< m2 >>
rect 69 7 70 8 
<< m1 >>
rect 70 7 71 8 
<< m2 >>
rect 70 7 71 8 
<< m1 >>
rect 71 7 72 8 
<< m2 >>
rect 71 7 72 8 
<< m1 >>
rect 72 7 73 8 
<< m2 >>
rect 72 7 73 8 
<< m1 >>
rect 73 7 74 8 
<< m2 >>
rect 73 7 74 8 
<< m1 >>
rect 74 7 75 8 
<< m2 >>
rect 74 7 75 8 
<< m1 >>
rect 75 7 76 8 
<< m2 >>
rect 75 7 76 8 
<< m1 >>
rect 76 7 77 8 
<< m2 >>
rect 76 7 77 8 
<< m1 >>
rect 77 7 78 8 
<< m2 >>
rect 77 7 78 8 
<< m1 >>
rect 78 7 79 8 
<< m2 >>
rect 78 7 79 8 
<< m1 >>
rect 79 7 80 8 
<< m2 >>
rect 79 7 80 8 
<< m1 >>
rect 80 7 81 8 
<< m2 >>
rect 80 7 81 8 
<< m1 >>
rect 81 7 82 8 
<< m2 >>
rect 81 7 82 8 
<< m1 >>
rect 82 7 83 8 
<< m2 >>
rect 82 7 83 8 
<< m2 >>
rect 83 7 84 8 
<< m1 >>
rect 84 7 85 8 
<< m2 >>
rect 84 7 85 8 
<< m2c >>
rect 84 7 85 8 
<< m1 >>
rect 84 7 85 8 
<< m2 >>
rect 84 7 85 8 
<< m1 >>
rect 85 7 86 8 
<< m1 >>
rect 86 7 87 8 
<< m1 >>
rect 87 7 88 8 
<< m1 >>
rect 88 7 89 8 
<< m1 >>
rect 89 7 90 8 
<< m1 >>
rect 90 7 91 8 
<< m1 >>
rect 91 7 92 8 
<< m1 >>
rect 92 7 93 8 
<< m1 >>
rect 93 7 94 8 
<< m1 >>
rect 94 7 95 8 
<< m1 >>
rect 95 7 96 8 
<< m1 >>
rect 96 7 97 8 
<< m1 >>
rect 97 7 98 8 
<< m1 >>
rect 98 7 99 8 
<< m1 >>
rect 99 7 100 8 
<< m1 >>
rect 100 7 101 8 
<< m1 >>
rect 101 7 102 8 
<< m1 >>
rect 102 7 103 8 
<< m1 >>
rect 103 7 104 8 
<< m1 >>
rect 104 7 105 8 
<< m1 >>
rect 105 7 106 8 
<< m1 >>
rect 106 7 107 8 
<< m1 >>
rect 107 7 108 8 
<< m1 >>
rect 108 7 109 8 
<< m1 >>
rect 109 7 110 8 
<< m1 >>
rect 110 7 111 8 
<< m1 >>
rect 111 7 112 8 
<< m1 >>
rect 112 7 113 8 
<< m1 >>
rect 113 7 114 8 
<< m1 >>
rect 114 7 115 8 
<< m1 >>
rect 115 7 116 8 
<< m1 >>
rect 116 7 117 8 
<< m1 >>
rect 117 7 118 8 
<< m1 >>
rect 118 7 119 8 
<< m1 >>
rect 119 7 120 8 
<< m1 >>
rect 120 7 121 8 
<< m1 >>
rect 121 7 122 8 
<< m1 >>
rect 122 7 123 8 
<< m1 >>
rect 123 7 124 8 
<< m1 >>
rect 124 7 125 8 
<< m1 >>
rect 125 7 126 8 
<< m1 >>
rect 126 7 127 8 
<< m1 >>
rect 127 7 128 8 
<< m2 >>
rect 16 8 17 9 
<< m2 >>
rect 17 8 18 9 
<< m2 >>
rect 18 8 19 9 
<< m2 >>
rect 19 8 20 9 
<< m2 >>
rect 20 8 21 9 
<< m2 >>
rect 21 8 22 9 
<< m2 >>
rect 22 8 23 9 
<< m2 >>
rect 23 8 24 9 
<< m2 >>
rect 24 8 25 9 
<< m2 >>
rect 25 8 26 9 
<< m2 >>
rect 26 8 27 9 
<< m2 >>
rect 27 8 28 9 
<< m2 >>
rect 28 8 29 9 
<< m2 >>
rect 29 8 30 9 
<< m1 >>
rect 30 8 31 9 
<< m2 >>
rect 30 8 31 9 
<< m2c >>
rect 30 8 31 9 
<< m1 >>
rect 30 8 31 9 
<< m2 >>
rect 30 8 31 9 
<< m1 >>
rect 44 8 45 9 
<< m1 >>
rect 82 8 83 9 
<< m1 >>
rect 127 8 128 9 
<< m1 >>
rect 13 9 14 10 
<< m1 >>
rect 14 9 15 10 
<< m1 >>
rect 15 9 16 10 
<< m1 >>
rect 16 9 17 10 
<< m2 >>
rect 16 9 17 10 
<< m1 >>
rect 17 9 18 10 
<< m1 >>
rect 18 9 19 10 
<< m1 >>
rect 19 9 20 10 
<< m1 >>
rect 20 9 21 10 
<< m1 >>
rect 21 9 22 10 
<< m1 >>
rect 22 9 23 10 
<< m1 >>
rect 23 9 24 10 
<< m1 >>
rect 24 9 25 10 
<< m1 >>
rect 25 9 26 10 
<< m1 >>
rect 26 9 27 10 
<< m1 >>
rect 27 9 28 10 
<< m1 >>
rect 28 9 29 10 
<< m1 >>
rect 44 9 45 10 
<< m1 >>
rect 82 9 83 10 
<< m1 >>
rect 85 9 86 10 
<< m1 >>
rect 86 9 87 10 
<< m1 >>
rect 87 9 88 10 
<< m1 >>
rect 88 9 89 10 
<< m1 >>
rect 89 9 90 10 
<< m1 >>
rect 90 9 91 10 
<< m1 >>
rect 91 9 92 10 
<< m1 >>
rect 103 9 104 10 
<< m1 >>
rect 104 9 105 10 
<< m1 >>
rect 105 9 106 10 
<< m1 >>
rect 106 9 107 10 
<< m1 >>
rect 107 9 108 10 
<< m1 >>
rect 108 9 109 10 
<< m1 >>
rect 109 9 110 10 
<< m1 >>
rect 127 9 128 10 
<< m1 >>
rect 13 10 14 11 
<< m2 >>
rect 16 10 17 11 
<< m1 >>
rect 28 10 29 11 
<< m1 >>
rect 34 10 35 11 
<< m1 >>
rect 35 10 36 11 
<< m1 >>
rect 36 10 37 11 
<< m1 >>
rect 37 10 38 11 
<< m1 >>
rect 44 10 45 11 
<< m1 >>
rect 46 10 47 11 
<< m1 >>
rect 47 10 48 11 
<< m1 >>
rect 48 10 49 11 
<< m1 >>
rect 49 10 50 11 
<< m1 >>
rect 70 10 71 11 
<< m1 >>
rect 71 10 72 11 
<< m1 >>
rect 72 10 73 11 
<< m1 >>
rect 73 10 74 11 
<< m1 >>
rect 82 10 83 11 
<< m1 >>
rect 85 10 86 11 
<< m1 >>
rect 91 10 92 11 
<< m1 >>
rect 103 10 104 11 
<< m1 >>
rect 109 10 110 11 
<< m1 >>
rect 127 10 128 11 
<< m1 >>
rect 13 11 14 12 
<< m1 >>
rect 16 11 17 12 
<< m2 >>
rect 16 11 17 12 
<< m2c >>
rect 16 11 17 12 
<< m1 >>
rect 16 11 17 12 
<< m2 >>
rect 16 11 17 12 
<< m1 >>
rect 28 11 29 12 
<< m1 >>
rect 34 11 35 12 
<< m1 >>
rect 37 11 38 12 
<< m1 >>
rect 44 11 45 12 
<< m1 >>
rect 46 11 47 12 
<< m1 >>
rect 49 11 50 12 
<< m1 >>
rect 70 11 71 12 
<< m1 >>
rect 73 11 74 12 
<< m1 >>
rect 82 11 83 12 
<< m1 >>
rect 85 11 86 12 
<< m1 >>
rect 91 11 92 12 
<< m1 >>
rect 103 11 104 12 
<< m1 >>
rect 109 11 110 12 
<< m1 >>
rect 127 11 128 12 
<< pdiffusion >>
rect 12 12 13 13 
<< m1 >>
rect 13 12 14 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< m1 >>
rect 16 12 17 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< m1 >>
rect 28 12 29 13 
<< pdiffusion >>
rect 30 12 31 13 
<< pdiffusion >>
rect 31 12 32 13 
<< pdiffusion >>
rect 32 12 33 13 
<< pdiffusion >>
rect 33 12 34 13 
<< m1 >>
rect 34 12 35 13 
<< pdiffusion >>
rect 34 12 35 13 
<< pdiffusion >>
rect 35 12 36 13 
<< m1 >>
rect 37 12 38 13 
<< m1 >>
rect 44 12 45 13 
<< m1 >>
rect 46 12 47 13 
<< pdiffusion >>
rect 48 12 49 13 
<< m1 >>
rect 49 12 50 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< pdiffusion >>
rect 51 12 52 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< pdiffusion >>
rect 66 12 67 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< m1 >>
rect 70 12 71 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< m1 >>
rect 73 12 74 13 
<< m1 >>
rect 82 12 83 13 
<< pdiffusion >>
rect 84 12 85 13 
<< m1 >>
rect 85 12 86 13 
<< pdiffusion >>
rect 85 12 86 13 
<< pdiffusion >>
rect 86 12 87 13 
<< pdiffusion >>
rect 87 12 88 13 
<< pdiffusion >>
rect 88 12 89 13 
<< pdiffusion >>
rect 89 12 90 13 
<< m1 >>
rect 91 12 92 13 
<< pdiffusion >>
rect 102 12 103 13 
<< m1 >>
rect 103 12 104 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< m1 >>
rect 109 12 110 13 
<< pdiffusion >>
rect 120 12 121 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< m1 >>
rect 127 12 128 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< m1 >>
rect 28 13 29 14 
<< pdiffusion >>
rect 30 13 31 14 
<< pdiffusion >>
rect 31 13 32 14 
<< pdiffusion >>
rect 32 13 33 14 
<< pdiffusion >>
rect 33 13 34 14 
<< pdiffusion >>
rect 34 13 35 14 
<< pdiffusion >>
rect 35 13 36 14 
<< m1 >>
rect 37 13 38 14 
<< m1 >>
rect 44 13 45 14 
<< m1 >>
rect 46 13 47 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< m1 >>
rect 73 13 74 14 
<< m1 >>
rect 82 13 83 14 
<< pdiffusion >>
rect 84 13 85 14 
<< pdiffusion >>
rect 85 13 86 14 
<< pdiffusion >>
rect 86 13 87 14 
<< pdiffusion >>
rect 87 13 88 14 
<< pdiffusion >>
rect 88 13 89 14 
<< pdiffusion >>
rect 89 13 90 14 
<< m1 >>
rect 91 13 92 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< m1 >>
rect 109 13 110 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< m1 >>
rect 127 13 128 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< m1 >>
rect 28 14 29 15 
<< pdiffusion >>
rect 30 14 31 15 
<< pdiffusion >>
rect 31 14 32 15 
<< pdiffusion >>
rect 32 14 33 15 
<< pdiffusion >>
rect 33 14 34 15 
<< pdiffusion >>
rect 34 14 35 15 
<< pdiffusion >>
rect 35 14 36 15 
<< m1 >>
rect 37 14 38 15 
<< m1 >>
rect 44 14 45 15 
<< m1 >>
rect 46 14 47 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< m1 >>
rect 73 14 74 15 
<< m1 >>
rect 82 14 83 15 
<< pdiffusion >>
rect 84 14 85 15 
<< pdiffusion >>
rect 85 14 86 15 
<< pdiffusion >>
rect 86 14 87 15 
<< pdiffusion >>
rect 87 14 88 15 
<< pdiffusion >>
rect 88 14 89 15 
<< pdiffusion >>
rect 89 14 90 15 
<< m1 >>
rect 91 14 92 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< m1 >>
rect 109 14 110 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< m1 >>
rect 127 14 128 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< m1 >>
rect 28 15 29 16 
<< pdiffusion >>
rect 30 15 31 16 
<< pdiffusion >>
rect 31 15 32 16 
<< pdiffusion >>
rect 32 15 33 16 
<< pdiffusion >>
rect 33 15 34 16 
<< pdiffusion >>
rect 34 15 35 16 
<< pdiffusion >>
rect 35 15 36 16 
<< m1 >>
rect 37 15 38 16 
<< m1 >>
rect 44 15 45 16 
<< m1 >>
rect 46 15 47 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< m1 >>
rect 73 15 74 16 
<< m1 >>
rect 82 15 83 16 
<< pdiffusion >>
rect 84 15 85 16 
<< pdiffusion >>
rect 85 15 86 16 
<< pdiffusion >>
rect 86 15 87 16 
<< pdiffusion >>
rect 87 15 88 16 
<< pdiffusion >>
rect 88 15 89 16 
<< pdiffusion >>
rect 89 15 90 16 
<< m1 >>
rect 91 15 92 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< m1 >>
rect 109 15 110 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< m1 >>
rect 127 15 128 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< m1 >>
rect 28 16 29 17 
<< pdiffusion >>
rect 30 16 31 17 
<< pdiffusion >>
rect 31 16 32 17 
<< pdiffusion >>
rect 32 16 33 17 
<< pdiffusion >>
rect 33 16 34 17 
<< pdiffusion >>
rect 34 16 35 17 
<< pdiffusion >>
rect 35 16 36 17 
<< m1 >>
rect 37 16 38 17 
<< m1 >>
rect 44 16 45 17 
<< m1 >>
rect 46 16 47 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< m1 >>
rect 73 16 74 17 
<< m1 >>
rect 82 16 83 17 
<< pdiffusion >>
rect 84 16 85 17 
<< pdiffusion >>
rect 85 16 86 17 
<< pdiffusion >>
rect 86 16 87 17 
<< pdiffusion >>
rect 87 16 88 17 
<< pdiffusion >>
rect 88 16 89 17 
<< pdiffusion >>
rect 89 16 90 17 
<< m1 >>
rect 91 16 92 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< m1 >>
rect 109 16 110 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< m1 >>
rect 127 16 128 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< m1 >>
rect 28 17 29 18 
<< pdiffusion >>
rect 30 17 31 18 
<< pdiffusion >>
rect 31 17 32 18 
<< pdiffusion >>
rect 32 17 33 18 
<< pdiffusion >>
rect 33 17 34 18 
<< m1 >>
rect 34 17 35 18 
<< pdiffusion >>
rect 34 17 35 18 
<< pdiffusion >>
rect 35 17 36 18 
<< m1 >>
rect 37 17 38 18 
<< m2 >>
rect 37 17 38 18 
<< m2c >>
rect 37 17 38 18 
<< m1 >>
rect 37 17 38 18 
<< m2 >>
rect 37 17 38 18 
<< m1 >>
rect 44 17 45 18 
<< m1 >>
rect 46 17 47 18 
<< pdiffusion >>
rect 48 17 49 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< m1 >>
rect 52 17 53 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< pdiffusion >>
rect 66 17 67 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< m1 >>
rect 73 17 74 18 
<< m1 >>
rect 82 17 83 18 
<< pdiffusion >>
rect 84 17 85 18 
<< m1 >>
rect 85 17 86 18 
<< pdiffusion >>
rect 85 17 86 18 
<< pdiffusion >>
rect 86 17 87 18 
<< pdiffusion >>
rect 87 17 88 18 
<< pdiffusion >>
rect 88 17 89 18 
<< pdiffusion >>
rect 89 17 90 18 
<< m1 >>
rect 91 17 92 18 
<< pdiffusion >>
rect 102 17 103 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< m1 >>
rect 109 17 110 18 
<< pdiffusion >>
rect 120 17 121 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< m1 >>
rect 124 17 125 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< m1 >>
rect 127 17 128 18 
<< m1 >>
rect 28 18 29 19 
<< m1 >>
rect 34 18 35 19 
<< m2 >>
rect 37 18 38 19 
<< m1 >>
rect 44 18 45 19 
<< m1 >>
rect 46 18 47 19 
<< m1 >>
rect 52 18 53 19 
<< m1 >>
rect 73 18 74 19 
<< m1 >>
rect 82 18 83 19 
<< m1 >>
rect 85 18 86 19 
<< m1 >>
rect 91 18 92 19 
<< m1 >>
rect 109 18 110 19 
<< m1 >>
rect 124 18 125 19 
<< m1 >>
rect 127 18 128 19 
<< m1 >>
rect 28 19 29 20 
<< m1 >>
rect 34 19 35 20 
<< m1 >>
rect 35 19 36 20 
<< m1 >>
rect 36 19 37 20 
<< m1 >>
rect 37 19 38 20 
<< m2 >>
rect 37 19 38 20 
<< m1 >>
rect 38 19 39 20 
<< m1 >>
rect 39 19 40 20 
<< m1 >>
rect 40 19 41 20 
<< m1 >>
rect 41 19 42 20 
<< m1 >>
rect 42 19 43 20 
<< m1 >>
rect 43 19 44 20 
<< m1 >>
rect 44 19 45 20 
<< m1 >>
rect 46 19 47 20 
<< m1 >>
rect 52 19 53 20 
<< m1 >>
rect 71 19 72 20 
<< m2 >>
rect 71 19 72 20 
<< m2c >>
rect 71 19 72 20 
<< m1 >>
rect 71 19 72 20 
<< m2 >>
rect 71 19 72 20 
<< m2 >>
rect 72 19 73 20 
<< m1 >>
rect 73 19 74 20 
<< m2 >>
rect 73 19 74 20 
<< m2 >>
rect 74 19 75 20 
<< m1 >>
rect 75 19 76 20 
<< m2 >>
rect 75 19 76 20 
<< m2c >>
rect 75 19 76 20 
<< m1 >>
rect 75 19 76 20 
<< m2 >>
rect 75 19 76 20 
<< m1 >>
rect 76 19 77 20 
<< m1 >>
rect 77 19 78 20 
<< m1 >>
rect 78 19 79 20 
<< m1 >>
rect 79 19 80 20 
<< m1 >>
rect 80 19 81 20 
<< m2 >>
rect 80 19 81 20 
<< m2c >>
rect 80 19 81 20 
<< m1 >>
rect 80 19 81 20 
<< m2 >>
rect 80 19 81 20 
<< m2 >>
rect 81 19 82 20 
<< m1 >>
rect 82 19 83 20 
<< m2 >>
rect 82 19 83 20 
<< m2 >>
rect 83 19 84 20 
<< m1 >>
rect 84 19 85 20 
<< m2 >>
rect 84 19 85 20 
<< m2c >>
rect 84 19 85 20 
<< m1 >>
rect 84 19 85 20 
<< m2 >>
rect 84 19 85 20 
<< m1 >>
rect 85 19 86 20 
<< m1 >>
rect 91 19 92 20 
<< m1 >>
rect 109 19 110 20 
<< m1 >>
rect 124 19 125 20 
<< m1 >>
rect 127 19 128 20 
<< m1 >>
rect 28 20 29 21 
<< m2 >>
rect 37 20 38 21 
<< m1 >>
rect 46 20 47 21 
<< m1 >>
rect 52 20 53 21 
<< m1 >>
rect 71 20 72 21 
<< m1 >>
rect 73 20 74 21 
<< m1 >>
rect 82 20 83 21 
<< m1 >>
rect 91 20 92 21 
<< m1 >>
rect 109 20 110 21 
<< m1 >>
rect 124 20 125 21 
<< m1 >>
rect 127 20 128 21 
<< m1 >>
rect 28 21 29 22 
<< m1 >>
rect 32 21 33 22 
<< m1 >>
rect 33 21 34 22 
<< m1 >>
rect 34 21 35 22 
<< m1 >>
rect 35 21 36 22 
<< m1 >>
rect 36 21 37 22 
<< m1 >>
rect 37 21 38 22 
<< m2 >>
rect 37 21 38 22 
<< m1 >>
rect 38 21 39 22 
<< m1 >>
rect 39 21 40 22 
<< m1 >>
rect 40 21 41 22 
<< m1 >>
rect 41 21 42 22 
<< m1 >>
rect 42 21 43 22 
<< m1 >>
rect 43 21 44 22 
<< m1 >>
rect 44 21 45 22 
<< m2 >>
rect 44 21 45 22 
<< m2c >>
rect 44 21 45 22 
<< m1 >>
rect 44 21 45 22 
<< m2 >>
rect 44 21 45 22 
<< m2 >>
rect 45 21 46 22 
<< m1 >>
rect 46 21 47 22 
<< m2 >>
rect 46 21 47 22 
<< m2 >>
rect 47 21 48 22 
<< m1 >>
rect 48 21 49 22 
<< m2 >>
rect 48 21 49 22 
<< m2c >>
rect 48 21 49 22 
<< m1 >>
rect 48 21 49 22 
<< m2 >>
rect 48 21 49 22 
<< m1 >>
rect 52 21 53 22 
<< m1 >>
rect 71 21 72 22 
<< m1 >>
rect 73 21 74 22 
<< m1 >>
rect 82 21 83 22 
<< m1 >>
rect 91 21 92 22 
<< m1 >>
rect 109 21 110 22 
<< m1 >>
rect 124 21 125 22 
<< m1 >>
rect 127 21 128 22 
<< m1 >>
rect 28 22 29 23 
<< m1 >>
rect 32 22 33 23 
<< m2 >>
rect 37 22 38 23 
<< m1 >>
rect 46 22 47 23 
<< m1 >>
rect 48 22 49 23 
<< m1 >>
rect 49 22 50 23 
<< m1 >>
rect 50 22 51 23 
<< m1 >>
rect 51 22 52 23 
<< m1 >>
rect 52 22 53 23 
<< m1 >>
rect 64 22 65 23 
<< m1 >>
rect 65 22 66 23 
<< m1 >>
rect 66 22 67 23 
<< m1 >>
rect 67 22 68 23 
<< m1 >>
rect 68 22 69 23 
<< m1 >>
rect 69 22 70 23 
<< m1 >>
rect 70 22 71 23 
<< m1 >>
rect 71 22 72 23 
<< m1 >>
rect 73 22 74 23 
<< m1 >>
rect 82 22 83 23 
<< m1 >>
rect 91 22 92 23 
<< m1 >>
rect 109 22 110 23 
<< m1 >>
rect 110 22 111 23 
<< m1 >>
rect 111 22 112 23 
<< m1 >>
rect 112 22 113 23 
<< m1 >>
rect 113 22 114 23 
<< m1 >>
rect 114 22 115 23 
<< m1 >>
rect 115 22 116 23 
<< m1 >>
rect 116 22 117 23 
<< m1 >>
rect 117 22 118 23 
<< m1 >>
rect 118 22 119 23 
<< m1 >>
rect 119 22 120 23 
<< m1 >>
rect 120 22 121 23 
<< m1 >>
rect 121 22 122 23 
<< m1 >>
rect 122 22 123 23 
<< m1 >>
rect 123 22 124 23 
<< m1 >>
rect 124 22 125 23 
<< m1 >>
rect 127 22 128 23 
<< m2 >>
rect 27 23 28 24 
<< m1 >>
rect 28 23 29 24 
<< m2 >>
rect 28 23 29 24 
<< m2 >>
rect 29 23 30 24 
<< m1 >>
rect 30 23 31 24 
<< m2 >>
rect 30 23 31 24 
<< m2c >>
rect 30 23 31 24 
<< m1 >>
rect 30 23 31 24 
<< m2 >>
rect 30 23 31 24 
<< m1 >>
rect 31 23 32 24 
<< m1 >>
rect 32 23 33 24 
<< m1 >>
rect 37 23 38 24 
<< m2 >>
rect 37 23 38 24 
<< m2c >>
rect 37 23 38 24 
<< m1 >>
rect 37 23 38 24 
<< m2 >>
rect 37 23 38 24 
<< m1 >>
rect 46 23 47 24 
<< m2 >>
rect 46 23 47 24 
<< m2c >>
rect 46 23 47 24 
<< m1 >>
rect 46 23 47 24 
<< m2 >>
rect 46 23 47 24 
<< m1 >>
rect 64 23 65 24 
<< m2 >>
rect 64 23 65 24 
<< m2c >>
rect 64 23 65 24 
<< m1 >>
rect 64 23 65 24 
<< m2 >>
rect 64 23 65 24 
<< m1 >>
rect 73 23 74 24 
<< m1 >>
rect 75 23 76 24 
<< m1 >>
rect 76 23 77 24 
<< m1 >>
rect 77 23 78 24 
<< m1 >>
rect 78 23 79 24 
<< m1 >>
rect 79 23 80 24 
<< m1 >>
rect 80 23 81 24 
<< m2 >>
rect 80 23 81 24 
<< m2c >>
rect 80 23 81 24 
<< m1 >>
rect 80 23 81 24 
<< m2 >>
rect 80 23 81 24 
<< m2 >>
rect 81 23 82 24 
<< m1 >>
rect 82 23 83 24 
<< m2 >>
rect 82 23 83 24 
<< m2 >>
rect 83 23 84 24 
<< m1 >>
rect 84 23 85 24 
<< m2 >>
rect 84 23 85 24 
<< m2c >>
rect 84 23 85 24 
<< m1 >>
rect 84 23 85 24 
<< m2 >>
rect 84 23 85 24 
<< m1 >>
rect 85 23 86 24 
<< m1 >>
rect 86 23 87 24 
<< m1 >>
rect 87 23 88 24 
<< m1 >>
rect 88 23 89 24 
<< m1 >>
rect 89 23 90 24 
<< m2 >>
rect 89 23 90 24 
<< m2c >>
rect 89 23 90 24 
<< m1 >>
rect 89 23 90 24 
<< m2 >>
rect 89 23 90 24 
<< m2 >>
rect 90 23 91 24 
<< m1 >>
rect 91 23 92 24 
<< m2 >>
rect 91 23 92 24 
<< m2 >>
rect 92 23 93 24 
<< m2 >>
rect 93 23 94 24 
<< m2 >>
rect 94 23 95 24 
<< m2 >>
rect 95 23 96 24 
<< m2 >>
rect 96 23 97 24 
<< m2 >>
rect 97 23 98 24 
<< m2 >>
rect 98 23 99 24 
<< m2 >>
rect 99 23 100 24 
<< m2 >>
rect 100 23 101 24 
<< m2 >>
rect 101 23 102 24 
<< m2 >>
rect 102 23 103 24 
<< m2 >>
rect 103 23 104 24 
<< m2 >>
rect 104 23 105 24 
<< m2 >>
rect 105 23 106 24 
<< m2 >>
rect 106 23 107 24 
<< m2 >>
rect 107 23 108 24 
<< m2 >>
rect 108 23 109 24 
<< m2 >>
rect 109 23 110 24 
<< m2 >>
rect 110 23 111 24 
<< m2 >>
rect 111 23 112 24 
<< m2 >>
rect 112 23 113 24 
<< m2 >>
rect 113 23 114 24 
<< m2 >>
rect 114 23 115 24 
<< m2 >>
rect 115 23 116 24 
<< m2 >>
rect 116 23 117 24 
<< m2 >>
rect 117 23 118 24 
<< m2 >>
rect 118 23 119 24 
<< m2 >>
rect 119 23 120 24 
<< m2 >>
rect 120 23 121 24 
<< m2 >>
rect 121 23 122 24 
<< m2 >>
rect 122 23 123 24 
<< m2 >>
rect 123 23 124 24 
<< m2 >>
rect 124 23 125 24 
<< m2 >>
rect 125 23 126 24 
<< m2 >>
rect 126 23 127 24 
<< m1 >>
rect 127 23 128 24 
<< m2 >>
rect 127 23 128 24 
<< m2 >>
rect 27 24 28 25 
<< m1 >>
rect 28 24 29 25 
<< m2 >>
rect 37 24 38 25 
<< m2 >>
rect 46 24 47 25 
<< m2 >>
rect 64 24 65 25 
<< m2 >>
rect 66 24 67 25 
<< m2 >>
rect 67 24 68 25 
<< m2 >>
rect 68 24 69 25 
<< m2 >>
rect 69 24 70 25 
<< m2 >>
rect 70 24 71 25 
<< m2 >>
rect 71 24 72 25 
<< m1 >>
rect 72 24 73 25 
<< m2 >>
rect 72 24 73 25 
<< m2c >>
rect 72 24 73 25 
<< m1 >>
rect 72 24 73 25 
<< m2 >>
rect 72 24 73 25 
<< m1 >>
rect 73 24 74 25 
<< m1 >>
rect 75 24 76 25 
<< m1 >>
rect 82 24 83 25 
<< m1 >>
rect 91 24 92 25 
<< m1 >>
rect 92 24 93 25 
<< m1 >>
rect 93 24 94 25 
<< m1 >>
rect 94 24 95 25 
<< m1 >>
rect 95 24 96 25 
<< m1 >>
rect 96 24 97 25 
<< m1 >>
rect 97 24 98 25 
<< m1 >>
rect 98 24 99 25 
<< m1 >>
rect 99 24 100 25 
<< m1 >>
rect 100 24 101 25 
<< m1 >>
rect 101 24 102 25 
<< m1 >>
rect 102 24 103 25 
<< m1 >>
rect 103 24 104 25 
<< m1 >>
rect 104 24 105 25 
<< m1 >>
rect 105 24 106 25 
<< m1 >>
rect 106 24 107 25 
<< m1 >>
rect 107 24 108 25 
<< m1 >>
rect 108 24 109 25 
<< m1 >>
rect 109 24 110 25 
<< m1 >>
rect 110 24 111 25 
<< m1 >>
rect 111 24 112 25 
<< m1 >>
rect 112 24 113 25 
<< m1 >>
rect 113 24 114 25 
<< m1 >>
rect 114 24 115 25 
<< m1 >>
rect 115 24 116 25 
<< m1 >>
rect 116 24 117 25 
<< m1 >>
rect 127 24 128 25 
<< m2 >>
rect 127 24 128 25 
<< m2 >>
rect 27 25 28 26 
<< m1 >>
rect 28 25 29 26 
<< m1 >>
rect 29 25 30 26 
<< m1 >>
rect 30 25 31 26 
<< m1 >>
rect 31 25 32 26 
<< m1 >>
rect 32 25 33 26 
<< m1 >>
rect 33 25 34 26 
<< m1 >>
rect 34 25 35 26 
<< m1 >>
rect 35 25 36 26 
<< m1 >>
rect 36 25 37 26 
<< m1 >>
rect 37 25 38 26 
<< m2 >>
rect 37 25 38 26 
<< m1 >>
rect 38 25 39 26 
<< m1 >>
rect 39 25 40 26 
<< m1 >>
rect 40 25 41 26 
<< m1 >>
rect 41 25 42 26 
<< m1 >>
rect 42 25 43 26 
<< m1 >>
rect 43 25 44 26 
<< m1 >>
rect 44 25 45 26 
<< m1 >>
rect 45 25 46 26 
<< m1 >>
rect 46 25 47 26 
<< m2 >>
rect 46 25 47 26 
<< m1 >>
rect 47 25 48 26 
<< m1 >>
rect 48 25 49 26 
<< m1 >>
rect 49 25 50 26 
<< m1 >>
rect 50 25 51 26 
<< m1 >>
rect 51 25 52 26 
<< m1 >>
rect 52 25 53 26 
<< m1 >>
rect 53 25 54 26 
<< m1 >>
rect 54 25 55 26 
<< m1 >>
rect 55 25 56 26 
<< m1 >>
rect 56 25 57 26 
<< m1 >>
rect 57 25 58 26 
<< m1 >>
rect 58 25 59 26 
<< m1 >>
rect 59 25 60 26 
<< m1 >>
rect 60 25 61 26 
<< m1 >>
rect 61 25 62 26 
<< m1 >>
rect 62 25 63 26 
<< m1 >>
rect 63 25 64 26 
<< m1 >>
rect 64 25 65 26 
<< m2 >>
rect 64 25 65 26 
<< m1 >>
rect 65 25 66 26 
<< m1 >>
rect 66 25 67 26 
<< m2 >>
rect 66 25 67 26 
<< m1 >>
rect 67 25 68 26 
<< m1 >>
rect 68 25 69 26 
<< m1 >>
rect 69 25 70 26 
<< m1 >>
rect 70 25 71 26 
<< m1 >>
rect 75 25 76 26 
<< m1 >>
rect 82 25 83 26 
<< m2 >>
rect 82 25 83 26 
<< m2 >>
rect 83 25 84 26 
<< m1 >>
rect 84 25 85 26 
<< m2 >>
rect 84 25 85 26 
<< m2c >>
rect 84 25 85 26 
<< m1 >>
rect 84 25 85 26 
<< m2 >>
rect 84 25 85 26 
<< m1 >>
rect 85 25 86 26 
<< m1 >>
rect 86 25 87 26 
<< m1 >>
rect 87 25 88 26 
<< m1 >>
rect 88 25 89 26 
<< m1 >>
rect 89 25 90 26 
<< m1 >>
rect 116 25 117 26 
<< m1 >>
rect 127 25 128 26 
<< m2 >>
rect 127 25 128 26 
<< m2 >>
rect 27 26 28 27 
<< m2 >>
rect 37 26 38 27 
<< m2 >>
rect 46 26 47 27 
<< m2 >>
rect 64 26 65 27 
<< m2 >>
rect 66 26 67 27 
<< m1 >>
rect 70 26 71 27 
<< m1 >>
rect 75 26 76 27 
<< m1 >>
rect 82 26 83 27 
<< m2 >>
rect 82 26 83 27 
<< m1 >>
rect 89 26 90 27 
<< m1 >>
rect 116 26 117 27 
<< m1 >>
rect 127 26 128 27 
<< m2 >>
rect 127 26 128 27 
<< m1 >>
rect 27 27 28 28 
<< m2 >>
rect 27 27 28 28 
<< m2c >>
rect 27 27 28 28 
<< m1 >>
rect 27 27 28 28 
<< m2 >>
rect 27 27 28 28 
<< m1 >>
rect 37 27 38 28 
<< m2 >>
rect 37 27 38 28 
<< m2c >>
rect 37 27 38 28 
<< m1 >>
rect 37 27 38 28 
<< m2 >>
rect 37 27 38 28 
<< m1 >>
rect 46 27 47 28 
<< m2 >>
rect 46 27 47 28 
<< m2c >>
rect 46 27 47 28 
<< m1 >>
rect 46 27 47 28 
<< m2 >>
rect 46 27 47 28 
<< m1 >>
rect 52 27 53 28 
<< m1 >>
rect 53 27 54 28 
<< m1 >>
rect 54 27 55 28 
<< m1 >>
rect 55 27 56 28 
<< m1 >>
rect 56 27 57 28 
<< m2 >>
rect 56 27 57 28 
<< m2c >>
rect 56 27 57 28 
<< m1 >>
rect 56 27 57 28 
<< m2 >>
rect 56 27 57 28 
<< m2 >>
rect 57 27 58 28 
<< m1 >>
rect 58 27 59 28 
<< m2 >>
rect 58 27 59 28 
<< m1 >>
rect 59 27 60 28 
<< m2 >>
rect 59 27 60 28 
<< m1 >>
rect 60 27 61 28 
<< m2 >>
rect 60 27 61 28 
<< m1 >>
rect 61 27 62 28 
<< m2 >>
rect 61 27 62 28 
<< m1 >>
rect 62 27 63 28 
<< m2 >>
rect 62 27 63 28 
<< m1 >>
rect 63 27 64 28 
<< m2 >>
rect 63 27 64 28 
<< m1 >>
rect 64 27 65 28 
<< m2 >>
rect 64 27 65 28 
<< m1 >>
rect 65 27 66 28 
<< m1 >>
rect 66 27 67 28 
<< m2 >>
rect 66 27 67 28 
<< m2c >>
rect 66 27 67 28 
<< m1 >>
rect 66 27 67 28 
<< m2 >>
rect 66 27 67 28 
<< m1 >>
rect 70 27 71 28 
<< m1 >>
rect 75 27 76 28 
<< m1 >>
rect 82 27 83 28 
<< m2 >>
rect 82 27 83 28 
<< m1 >>
rect 89 27 90 28 
<< m1 >>
rect 116 27 117 28 
<< m1 >>
rect 127 27 128 28 
<< m2 >>
rect 127 27 128 28 
<< m1 >>
rect 16 28 17 29 
<< m1 >>
rect 17 28 18 29 
<< m1 >>
rect 18 28 19 29 
<< m1 >>
rect 19 28 20 29 
<< m1 >>
rect 20 28 21 29 
<< m1 >>
rect 21 28 22 29 
<< m1 >>
rect 27 28 28 29 
<< m1 >>
rect 37 28 38 29 
<< m1 >>
rect 46 28 47 29 
<< m1 >>
rect 52 28 53 29 
<< m1 >>
rect 58 28 59 29 
<< m1 >>
rect 70 28 71 29 
<< m1 >>
rect 75 28 76 29 
<< m1 >>
rect 82 28 83 29 
<< m2 >>
rect 82 28 83 29 
<< m1 >>
rect 83 28 84 29 
<< m1 >>
rect 84 28 85 29 
<< m1 >>
rect 85 28 86 29 
<< m1 >>
rect 89 28 90 29 
<< m1 >>
rect 90 28 91 29 
<< m1 >>
rect 91 28 92 29 
<< m1 >>
rect 92 28 93 29 
<< m1 >>
rect 93 28 94 29 
<< m1 >>
rect 94 28 95 29 
<< m1 >>
rect 95 28 96 29 
<< m1 >>
rect 96 28 97 29 
<< m1 >>
rect 97 28 98 29 
<< m1 >>
rect 98 28 99 29 
<< m1 >>
rect 99 28 100 29 
<< m1 >>
rect 100 28 101 29 
<< m1 >>
rect 101 28 102 29 
<< m1 >>
rect 102 28 103 29 
<< m1 >>
rect 103 28 104 29 
<< m1 >>
rect 104 28 105 29 
<< m1 >>
rect 105 28 106 29 
<< m1 >>
rect 106 28 107 29 
<< m1 >>
rect 107 28 108 29 
<< m1 >>
rect 108 28 109 29 
<< m1 >>
rect 109 28 110 29 
<< m1 >>
rect 110 28 111 29 
<< m1 >>
rect 111 28 112 29 
<< m1 >>
rect 112 28 113 29 
<< m1 >>
rect 113 28 114 29 
<< m1 >>
rect 114 28 115 29 
<< m1 >>
rect 116 28 117 29 
<< m1 >>
rect 127 28 128 29 
<< m2 >>
rect 127 28 128 29 
<< m1 >>
rect 16 29 17 30 
<< m1 >>
rect 21 29 22 30 
<< m1 >>
rect 27 29 28 30 
<< m1 >>
rect 37 29 38 30 
<< m1 >>
rect 46 29 47 30 
<< m1 >>
rect 52 29 53 30 
<< m1 >>
rect 58 29 59 30 
<< m1 >>
rect 70 29 71 30 
<< m1 >>
rect 75 29 76 30 
<< m2 >>
rect 82 29 83 30 
<< m1 >>
rect 85 29 86 30 
<< m1 >>
rect 114 29 115 30 
<< m1 >>
rect 116 29 117 30 
<< m1 >>
rect 127 29 128 30 
<< m2 >>
rect 127 29 128 30 
<< pdiffusion >>
rect 12 30 13 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< pdiffusion >>
rect 15 30 16 31 
<< m1 >>
rect 16 30 17 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< m1 >>
rect 21 30 22 31 
<< m1 >>
rect 27 30 28 31 
<< m1 >>
rect 37 30 38 31 
<< m1 >>
rect 46 30 47 31 
<< pdiffusion >>
rect 48 30 49 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< m1 >>
rect 52 30 53 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 58 30 59 31 
<< pdiffusion >>
rect 66 30 67 31 
<< pdiffusion >>
rect 67 30 68 31 
<< pdiffusion >>
rect 68 30 69 31 
<< pdiffusion >>
rect 69 30 70 31 
<< m1 >>
rect 70 30 71 31 
<< pdiffusion >>
rect 70 30 71 31 
<< pdiffusion >>
rect 71 30 72 31 
<< m1 >>
rect 75 30 76 31 
<< m1 >>
rect 82 30 83 31 
<< m2 >>
rect 82 30 83 31 
<< m2c >>
rect 82 30 83 31 
<< m1 >>
rect 82 30 83 31 
<< m2 >>
rect 82 30 83 31 
<< pdiffusion >>
rect 84 30 85 31 
<< m1 >>
rect 85 30 86 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< m1 >>
rect 114 30 115 31 
<< m1 >>
rect 116 30 117 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< m1 >>
rect 127 30 128 31 
<< m2 >>
rect 127 30 128 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< m1 >>
rect 21 31 22 32 
<< m1 >>
rect 27 31 28 32 
<< m1 >>
rect 37 31 38 32 
<< m1 >>
rect 46 31 47 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 58 31 59 32 
<< pdiffusion >>
rect 66 31 67 32 
<< pdiffusion >>
rect 67 31 68 32 
<< pdiffusion >>
rect 68 31 69 32 
<< pdiffusion >>
rect 69 31 70 32 
<< pdiffusion >>
rect 70 31 71 32 
<< pdiffusion >>
rect 71 31 72 32 
<< m1 >>
rect 75 31 76 32 
<< m1 >>
rect 82 31 83 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< m1 >>
rect 114 31 115 32 
<< m1 >>
rect 116 31 117 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< m1 >>
rect 127 31 128 32 
<< m2 >>
rect 127 31 128 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< m1 >>
rect 21 32 22 33 
<< m1 >>
rect 27 32 28 33 
<< m1 >>
rect 37 32 38 33 
<< m1 >>
rect 46 32 47 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 58 32 59 33 
<< pdiffusion >>
rect 66 32 67 33 
<< pdiffusion >>
rect 67 32 68 33 
<< pdiffusion >>
rect 68 32 69 33 
<< pdiffusion >>
rect 69 32 70 33 
<< pdiffusion >>
rect 70 32 71 33 
<< pdiffusion >>
rect 71 32 72 33 
<< m1 >>
rect 75 32 76 33 
<< m1 >>
rect 82 32 83 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< m1 >>
rect 114 32 115 33 
<< m1 >>
rect 116 32 117 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< m1 >>
rect 127 32 128 33 
<< m2 >>
rect 127 32 128 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< m1 >>
rect 21 33 22 34 
<< m1 >>
rect 27 33 28 34 
<< m1 >>
rect 37 33 38 34 
<< m1 >>
rect 46 33 47 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 58 33 59 34 
<< pdiffusion >>
rect 66 33 67 34 
<< pdiffusion >>
rect 67 33 68 34 
<< pdiffusion >>
rect 68 33 69 34 
<< pdiffusion >>
rect 69 33 70 34 
<< pdiffusion >>
rect 70 33 71 34 
<< pdiffusion >>
rect 71 33 72 34 
<< m1 >>
rect 75 33 76 34 
<< m1 >>
rect 82 33 83 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< m1 >>
rect 114 33 115 34 
<< m1 >>
rect 116 33 117 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< m1 >>
rect 127 33 128 34 
<< m2 >>
rect 127 33 128 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< m1 >>
rect 21 34 22 35 
<< m1 >>
rect 27 34 28 35 
<< m1 >>
rect 37 34 38 35 
<< m1 >>
rect 46 34 47 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 58 34 59 35 
<< pdiffusion >>
rect 66 34 67 35 
<< pdiffusion >>
rect 67 34 68 35 
<< pdiffusion >>
rect 68 34 69 35 
<< pdiffusion >>
rect 69 34 70 35 
<< pdiffusion >>
rect 70 34 71 35 
<< pdiffusion >>
rect 71 34 72 35 
<< m1 >>
rect 75 34 76 35 
<< m1 >>
rect 82 34 83 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< m1 >>
rect 114 34 115 35 
<< m1 >>
rect 116 34 117 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< m1 >>
rect 127 34 128 35 
<< m2 >>
rect 127 34 128 35 
<< pdiffusion >>
rect 12 35 13 36 
<< m1 >>
rect 13 35 14 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< m1 >>
rect 16 35 17 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< m1 >>
rect 21 35 22 36 
<< m1 >>
rect 27 35 28 36 
<< m1 >>
rect 37 35 38 36 
<< m1 >>
rect 46 35 47 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< m1 >>
rect 52 35 53 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 58 35 59 36 
<< pdiffusion >>
rect 66 35 67 36 
<< m1 >>
rect 67 35 68 36 
<< pdiffusion >>
rect 67 35 68 36 
<< pdiffusion >>
rect 68 35 69 36 
<< m1 >>
rect 69 35 70 36 
<< m2 >>
rect 69 35 70 36 
<< m2c >>
rect 69 35 70 36 
<< m1 >>
rect 69 35 70 36 
<< m2 >>
rect 69 35 70 36 
<< pdiffusion >>
rect 69 35 70 36 
<< m1 >>
rect 70 35 71 36 
<< pdiffusion >>
rect 70 35 71 36 
<< pdiffusion >>
rect 71 35 72 36 
<< m1 >>
rect 75 35 76 36 
<< m1 >>
rect 82 35 83 36 
<< pdiffusion >>
rect 84 35 85 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< m1 >>
rect 88 35 89 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< m1 >>
rect 114 35 115 36 
<< m1 >>
rect 116 35 117 36 
<< pdiffusion >>
rect 120 35 121 36 
<< m1 >>
rect 121 35 122 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< m1 >>
rect 124 35 125 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< m1 >>
rect 127 35 128 36 
<< m2 >>
rect 127 35 128 36 
<< m1 >>
rect 13 36 14 37 
<< m1 >>
rect 16 36 17 37 
<< m1 >>
rect 21 36 22 37 
<< m1 >>
rect 27 36 28 37 
<< m1 >>
rect 37 36 38 37 
<< m1 >>
rect 46 36 47 37 
<< m1 >>
rect 52 36 53 37 
<< m1 >>
rect 58 36 59 37 
<< m1 >>
rect 67 36 68 37 
<< m1 >>
rect 70 36 71 37 
<< m2 >>
rect 70 36 71 37 
<< m1 >>
rect 73 36 74 37 
<< m2 >>
rect 73 36 74 37 
<< m2c >>
rect 73 36 74 37 
<< m1 >>
rect 73 36 74 37 
<< m2 >>
rect 73 36 74 37 
<< m1 >>
rect 74 36 75 37 
<< m1 >>
rect 75 36 76 37 
<< m1 >>
rect 82 36 83 37 
<< m2 >>
rect 82 36 83 37 
<< m2c >>
rect 82 36 83 37 
<< m1 >>
rect 82 36 83 37 
<< m2 >>
rect 82 36 83 37 
<< m1 >>
rect 88 36 89 37 
<< m1 >>
rect 114 36 115 37 
<< m1 >>
rect 116 36 117 37 
<< m1 >>
rect 121 36 122 37 
<< m1 >>
rect 124 36 125 37 
<< m1 >>
rect 127 36 128 37 
<< m2 >>
rect 127 36 128 37 
<< m1 >>
rect 13 37 14 38 
<< m1 >>
rect 16 37 17 38 
<< m1 >>
rect 21 37 22 38 
<< m1 >>
rect 27 37 28 38 
<< m1 >>
rect 37 37 38 38 
<< m1 >>
rect 46 37 47 38 
<< m1 >>
rect 52 37 53 38 
<< m1 >>
rect 58 37 59 38 
<< m1 >>
rect 67 37 68 38 
<< m2 >>
rect 70 37 71 38 
<< m2 >>
rect 71 37 72 38 
<< m2 >>
rect 72 37 73 38 
<< m2 >>
rect 73 37 74 38 
<< m2 >>
rect 82 37 83 38 
<< m1 >>
rect 88 37 89 38 
<< m1 >>
rect 114 37 115 38 
<< m1 >>
rect 116 37 117 38 
<< m1 >>
rect 121 37 122 38 
<< m1 >>
rect 124 37 125 38 
<< m1 >>
rect 125 37 126 38 
<< m2 >>
rect 125 37 126 38 
<< m2c >>
rect 125 37 126 38 
<< m1 >>
rect 125 37 126 38 
<< m2 >>
rect 125 37 126 38 
<< m2 >>
rect 126 37 127 38 
<< m1 >>
rect 127 37 128 38 
<< m2 >>
rect 127 37 128 38 
<< m1 >>
rect 13 38 14 39 
<< m1 >>
rect 14 38 15 39 
<< m2 >>
rect 14 38 15 39 
<< m2c >>
rect 14 38 15 39 
<< m1 >>
rect 14 38 15 39 
<< m2 >>
rect 14 38 15 39 
<< m2 >>
rect 15 38 16 39 
<< m1 >>
rect 16 38 17 39 
<< m2 >>
rect 16 38 17 39 
<< m1 >>
rect 21 38 22 39 
<< m1 >>
rect 27 38 28 39 
<< m1 >>
rect 37 38 38 39 
<< m1 >>
rect 46 38 47 39 
<< m1 >>
rect 52 38 53 39 
<< m1 >>
rect 58 38 59 39 
<< m1 >>
rect 67 38 68 39 
<< m1 >>
rect 68 38 69 39 
<< m1 >>
rect 69 38 70 39 
<< m1 >>
rect 70 38 71 39 
<< m1 >>
rect 71 38 72 39 
<< m1 >>
rect 72 38 73 39 
<< m1 >>
rect 73 38 74 39 
<< m1 >>
rect 74 38 75 39 
<< m1 >>
rect 75 38 76 39 
<< m1 >>
rect 76 38 77 39 
<< m1 >>
rect 77 38 78 39 
<< m1 >>
rect 78 38 79 39 
<< m1 >>
rect 79 38 80 39 
<< m1 >>
rect 80 38 81 39 
<< m1 >>
rect 81 38 82 39 
<< m1 >>
rect 82 38 83 39 
<< m2 >>
rect 82 38 83 39 
<< m1 >>
rect 83 38 84 39 
<< m1 >>
rect 84 38 85 39 
<< m2 >>
rect 84 38 85 39 
<< m2c >>
rect 84 38 85 39 
<< m1 >>
rect 84 38 85 39 
<< m2 >>
rect 84 38 85 39 
<< m1 >>
rect 88 38 89 39 
<< m1 >>
rect 114 38 115 39 
<< m2 >>
rect 114 38 115 39 
<< m2c >>
rect 114 38 115 39 
<< m1 >>
rect 114 38 115 39 
<< m2 >>
rect 114 38 115 39 
<< m2 >>
rect 115 38 116 39 
<< m1 >>
rect 116 38 117 39 
<< m2 >>
rect 116 38 117 39 
<< m2 >>
rect 117 38 118 39 
<< m1 >>
rect 118 38 119 39 
<< m2 >>
rect 118 38 119 39 
<< m2c >>
rect 118 38 119 39 
<< m1 >>
rect 118 38 119 39 
<< m2 >>
rect 118 38 119 39 
<< m1 >>
rect 119 38 120 39 
<< m1 >>
rect 121 38 122 39 
<< m1 >>
rect 127 38 128 39 
<< m1 >>
rect 16 39 17 40 
<< m2 >>
rect 16 39 17 40 
<< m1 >>
rect 21 39 22 40 
<< m2 >>
rect 21 39 22 40 
<< m2c >>
rect 21 39 22 40 
<< m1 >>
rect 21 39 22 40 
<< m2 >>
rect 21 39 22 40 
<< m1 >>
rect 27 39 28 40 
<< m1 >>
rect 37 39 38 40 
<< m1 >>
rect 44 39 45 40 
<< m2 >>
rect 44 39 45 40 
<< m2c >>
rect 44 39 45 40 
<< m1 >>
rect 44 39 45 40 
<< m2 >>
rect 44 39 45 40 
<< m2 >>
rect 45 39 46 40 
<< m1 >>
rect 46 39 47 40 
<< m2 >>
rect 46 39 47 40 
<< m2 >>
rect 47 39 48 40 
<< m1 >>
rect 48 39 49 40 
<< m2 >>
rect 48 39 49 40 
<< m2c >>
rect 48 39 49 40 
<< m1 >>
rect 48 39 49 40 
<< m2 >>
rect 48 39 49 40 
<< m1 >>
rect 52 39 53 40 
<< m1 >>
rect 58 39 59 40 
<< m2 >>
rect 82 39 83 40 
<< m2 >>
rect 84 39 85 40 
<< m1 >>
rect 88 39 89 40 
<< m1 >>
rect 116 39 117 40 
<< m1 >>
rect 119 39 120 40 
<< m1 >>
rect 121 39 122 40 
<< m1 >>
rect 127 39 128 40 
<< m1 >>
rect 10 40 11 41 
<< m1 >>
rect 11 40 12 41 
<< m1 >>
rect 12 40 13 41 
<< m1 >>
rect 13 40 14 41 
<< m1 >>
rect 14 40 15 41 
<< m1 >>
rect 15 40 16 41 
<< m1 >>
rect 16 40 17 41 
<< m2 >>
rect 16 40 17 41 
<< m2 >>
rect 21 40 22 41 
<< m1 >>
rect 27 40 28 41 
<< m1 >>
rect 37 40 38 41 
<< m1 >>
rect 44 40 45 41 
<< m1 >>
rect 46 40 47 41 
<< m1 >>
rect 48 40 49 41 
<< m1 >>
rect 49 40 50 41 
<< m1 >>
rect 50 40 51 41 
<< m2 >>
rect 50 40 51 41 
<< m2c >>
rect 50 40 51 41 
<< m1 >>
rect 50 40 51 41 
<< m2 >>
rect 50 40 51 41 
<< m2 >>
rect 51 40 52 41 
<< m1 >>
rect 52 40 53 41 
<< m2 >>
rect 52 40 53 41 
<< m2 >>
rect 53 40 54 41 
<< m1 >>
rect 54 40 55 41 
<< m2 >>
rect 54 40 55 41 
<< m2c >>
rect 54 40 55 41 
<< m1 >>
rect 54 40 55 41 
<< m2 >>
rect 54 40 55 41 
<< m1 >>
rect 55 40 56 41 
<< m1 >>
rect 56 40 57 41 
<< m2 >>
rect 56 40 57 41 
<< m2c >>
rect 56 40 57 41 
<< m1 >>
rect 56 40 57 41 
<< m2 >>
rect 56 40 57 41 
<< m2 >>
rect 57 40 58 41 
<< m1 >>
rect 58 40 59 41 
<< m2 >>
rect 58 40 59 41 
<< m2 >>
rect 59 40 60 41 
<< m1 >>
rect 60 40 61 41 
<< m2 >>
rect 60 40 61 41 
<< m1 >>
rect 61 40 62 41 
<< m2 >>
rect 61 40 62 41 
<< m1 >>
rect 62 40 63 41 
<< m2 >>
rect 62 40 63 41 
<< m1 >>
rect 63 40 64 41 
<< m2 >>
rect 63 40 64 41 
<< m1 >>
rect 64 40 65 41 
<< m2 >>
rect 64 40 65 41 
<< m1 >>
rect 65 40 66 41 
<< m2 >>
rect 65 40 66 41 
<< m1 >>
rect 66 40 67 41 
<< m2 >>
rect 66 40 67 41 
<< m1 >>
rect 67 40 68 41 
<< m2 >>
rect 67 40 68 41 
<< m1 >>
rect 68 40 69 41 
<< m2 >>
rect 68 40 69 41 
<< m1 >>
rect 69 40 70 41 
<< m2 >>
rect 69 40 70 41 
<< m1 >>
rect 70 40 71 41 
<< m2 >>
rect 70 40 71 41 
<< m1 >>
rect 71 40 72 41 
<< m2 >>
rect 71 40 72 41 
<< m1 >>
rect 72 40 73 41 
<< m2 >>
rect 72 40 73 41 
<< m1 >>
rect 73 40 74 41 
<< m2 >>
rect 73 40 74 41 
<< m1 >>
rect 74 40 75 41 
<< m2 >>
rect 74 40 75 41 
<< m1 >>
rect 75 40 76 41 
<< m2 >>
rect 75 40 76 41 
<< m1 >>
rect 76 40 77 41 
<< m2 >>
rect 76 40 77 41 
<< m1 >>
rect 77 40 78 41 
<< m2 >>
rect 77 40 78 41 
<< m1 >>
rect 78 40 79 41 
<< m2 >>
rect 78 40 79 41 
<< m1 >>
rect 79 40 80 41 
<< m2 >>
rect 79 40 80 41 
<< m1 >>
rect 80 40 81 41 
<< m2 >>
rect 80 40 81 41 
<< m1 >>
rect 81 40 82 41 
<< m2 >>
rect 81 40 82 41 
<< m1 >>
rect 82 40 83 41 
<< m2 >>
rect 82 40 83 41 
<< m1 >>
rect 83 40 84 41 
<< m1 >>
rect 84 40 85 41 
<< m2 >>
rect 84 40 85 41 
<< m1 >>
rect 85 40 86 41 
<< m2 >>
rect 85 40 86 41 
<< m1 >>
rect 86 40 87 41 
<< m2 >>
rect 86 40 87 41 
<< m1 >>
rect 87 40 88 41 
<< m2 >>
rect 87 40 88 41 
<< m1 >>
rect 88 40 89 41 
<< m2 >>
rect 88 40 89 41 
<< m2 >>
rect 89 40 90 41 
<< m1 >>
rect 90 40 91 41 
<< m2 >>
rect 90 40 91 41 
<< m2c >>
rect 90 40 91 41 
<< m1 >>
rect 90 40 91 41 
<< m2 >>
rect 90 40 91 41 
<< m1 >>
rect 91 40 92 41 
<< m1 >>
rect 92 40 93 41 
<< m1 >>
rect 93 40 94 41 
<< m1 >>
rect 94 40 95 41 
<< m1 >>
rect 95 40 96 41 
<< m1 >>
rect 96 40 97 41 
<< m1 >>
rect 97 40 98 41 
<< m1 >>
rect 98 40 99 41 
<< m1 >>
rect 99 40 100 41 
<< m1 >>
rect 100 40 101 41 
<< m1 >>
rect 101 40 102 41 
<< m1 >>
rect 102 40 103 41 
<< m1 >>
rect 103 40 104 41 
<< m1 >>
rect 104 40 105 41 
<< m1 >>
rect 105 40 106 41 
<< m1 >>
rect 106 40 107 41 
<< m1 >>
rect 107 40 108 41 
<< m1 >>
rect 108 40 109 41 
<< m1 >>
rect 109 40 110 41 
<< m1 >>
rect 110 40 111 41 
<< m1 >>
rect 111 40 112 41 
<< m1 >>
rect 112 40 113 41 
<< m1 >>
rect 113 40 114 41 
<< m1 >>
rect 114 40 115 41 
<< m2 >>
rect 114 40 115 41 
<< m2c >>
rect 114 40 115 41 
<< m1 >>
rect 114 40 115 41 
<< m2 >>
rect 114 40 115 41 
<< m1 >>
rect 116 40 117 41 
<< m2 >>
rect 116 40 117 41 
<< m2c >>
rect 116 40 117 41 
<< m1 >>
rect 116 40 117 41 
<< m2 >>
rect 116 40 117 41 
<< m1 >>
rect 119 40 120 41 
<< m2 >>
rect 119 40 120 41 
<< m2c >>
rect 119 40 120 41 
<< m1 >>
rect 119 40 120 41 
<< m2 >>
rect 119 40 120 41 
<< m2 >>
rect 120 40 121 41 
<< m1 >>
rect 121 40 122 41 
<< m2 >>
rect 121 40 122 41 
<< m2 >>
rect 122 40 123 41 
<< m1 >>
rect 127 40 128 41 
<< m1 >>
rect 10 41 11 42 
<< m2 >>
rect 16 41 17 42 
<< m1 >>
rect 19 41 20 42 
<< m2 >>
rect 19 41 20 42 
<< m2c >>
rect 19 41 20 42 
<< m1 >>
rect 19 41 20 42 
<< m2 >>
rect 19 41 20 42 
<< m1 >>
rect 20 41 21 42 
<< m1 >>
rect 21 41 22 42 
<< m2 >>
rect 21 41 22 42 
<< m1 >>
rect 22 41 23 42 
<< m1 >>
rect 23 41 24 42 
<< m1 >>
rect 24 41 25 42 
<< m1 >>
rect 25 41 26 42 
<< m1 >>
rect 26 41 27 42 
<< m1 >>
rect 27 41 28 42 
<< m1 >>
rect 37 41 38 42 
<< m2 >>
rect 37 41 38 42 
<< m2c >>
rect 37 41 38 42 
<< m1 >>
rect 37 41 38 42 
<< m2 >>
rect 37 41 38 42 
<< m1 >>
rect 44 41 45 42 
<< m2 >>
rect 44 41 45 42 
<< m2c >>
rect 44 41 45 42 
<< m1 >>
rect 44 41 45 42 
<< m2 >>
rect 44 41 45 42 
<< m1 >>
rect 46 41 47 42 
<< m2 >>
rect 46 41 47 42 
<< m2c >>
rect 46 41 47 42 
<< m1 >>
rect 46 41 47 42 
<< m2 >>
rect 46 41 47 42 
<< m1 >>
rect 52 41 53 42 
<< m1 >>
rect 58 41 59 42 
<< m1 >>
rect 60 41 61 42 
<< m2 >>
rect 114 41 115 42 
<< m2 >>
rect 116 41 117 42 
<< m1 >>
rect 121 41 122 42 
<< m2 >>
rect 122 41 123 42 
<< m1 >>
rect 125 41 126 42 
<< m2 >>
rect 125 41 126 42 
<< m2c >>
rect 125 41 126 42 
<< m1 >>
rect 125 41 126 42 
<< m2 >>
rect 125 41 126 42 
<< m1 >>
rect 126 41 127 42 
<< m1 >>
rect 127 41 128 42 
<< m1 >>
rect 10 42 11 43 
<< m1 >>
rect 16 42 17 43 
<< m2 >>
rect 16 42 17 43 
<< m2c >>
rect 16 42 17 43 
<< m1 >>
rect 16 42 17 43 
<< m2 >>
rect 16 42 17 43 
<< m2 >>
rect 19 42 20 43 
<< m2 >>
rect 21 42 22 43 
<< m2 >>
rect 37 42 38 43 
<< m2 >>
rect 44 42 45 43 
<< m2 >>
rect 46 42 47 43 
<< m1 >>
rect 52 42 53 43 
<< m1 >>
rect 58 42 59 43 
<< m1 >>
rect 60 42 61 43 
<< m1 >>
rect 82 42 83 43 
<< m1 >>
rect 83 42 84 43 
<< m1 >>
rect 84 42 85 43 
<< m1 >>
rect 85 42 86 43 
<< m1 >>
rect 86 42 87 43 
<< m1 >>
rect 87 42 88 43 
<< m1 >>
rect 88 42 89 43 
<< m1 >>
rect 89 42 90 43 
<< m2 >>
rect 89 42 90 43 
<< m2c >>
rect 89 42 90 43 
<< m1 >>
rect 89 42 90 43 
<< m2 >>
rect 89 42 90 43 
<< m2 >>
rect 90 42 91 43 
<< m2 >>
rect 91 42 92 43 
<< m2 >>
rect 92 42 93 43 
<< m2 >>
rect 93 42 94 43 
<< m2 >>
rect 94 42 95 43 
<< m2 >>
rect 95 42 96 43 
<< m2 >>
rect 96 42 97 43 
<< m2 >>
rect 97 42 98 43 
<< m2 >>
rect 98 42 99 43 
<< m2 >>
rect 99 42 100 43 
<< m2 >>
rect 100 42 101 43 
<< m2 >>
rect 101 42 102 43 
<< m2 >>
rect 102 42 103 43 
<< m2 >>
rect 103 42 104 43 
<< m2 >>
rect 104 42 105 43 
<< m2 >>
rect 105 42 106 43 
<< m2 >>
rect 106 42 107 43 
<< m2 >>
rect 107 42 108 43 
<< m2 >>
rect 108 42 109 43 
<< m2 >>
rect 109 42 110 43 
<< m2 >>
rect 110 42 111 43 
<< m1 >>
rect 111 42 112 43 
<< m2 >>
rect 111 42 112 43 
<< m2c >>
rect 111 42 112 43 
<< m1 >>
rect 111 42 112 43 
<< m2 >>
rect 111 42 112 43 
<< m1 >>
rect 112 42 113 43 
<< m1 >>
rect 113 42 114 43 
<< m1 >>
rect 114 42 115 43 
<< m2 >>
rect 114 42 115 43 
<< m1 >>
rect 115 42 116 43 
<< m1 >>
rect 116 42 117 43 
<< m2 >>
rect 116 42 117 43 
<< m1 >>
rect 117 42 118 43 
<< m1 >>
rect 118 42 119 43 
<< m1 >>
rect 119 42 120 43 
<< m1 >>
rect 120 42 121 43 
<< m1 >>
rect 121 42 122 43 
<< m2 >>
rect 122 42 123 43 
<< m2 >>
rect 125 42 126 43 
<< m1 >>
rect 10 43 11 44 
<< m1 >>
rect 16 43 17 44 
<< m1 >>
rect 19 43 20 44 
<< m2 >>
rect 19 43 20 44 
<< m1 >>
rect 20 43 21 44 
<< m1 >>
rect 21 43 22 44 
<< m2 >>
rect 21 43 22 44 
<< m1 >>
rect 22 43 23 44 
<< m1 >>
rect 23 43 24 44 
<< m1 >>
rect 24 43 25 44 
<< m1 >>
rect 25 43 26 44 
<< m1 >>
rect 26 43 27 44 
<< m1 >>
rect 27 43 28 44 
<< m1 >>
rect 28 43 29 44 
<< m1 >>
rect 29 43 30 44 
<< m1 >>
rect 30 43 31 44 
<< m1 >>
rect 31 43 32 44 
<< m1 >>
rect 32 43 33 44 
<< m1 >>
rect 33 43 34 44 
<< m1 >>
rect 34 43 35 44 
<< m1 >>
rect 35 43 36 44 
<< m1 >>
rect 36 43 37 44 
<< m1 >>
rect 37 43 38 44 
<< m2 >>
rect 37 43 38 44 
<< m1 >>
rect 38 43 39 44 
<< m1 >>
rect 39 43 40 44 
<< m1 >>
rect 40 43 41 44 
<< m1 >>
rect 41 43 42 44 
<< m1 >>
rect 42 43 43 44 
<< m1 >>
rect 43 43 44 44 
<< m1 >>
rect 44 43 45 44 
<< m2 >>
rect 44 43 45 44 
<< m1 >>
rect 45 43 46 44 
<< m1 >>
rect 46 43 47 44 
<< m2 >>
rect 46 43 47 44 
<< m1 >>
rect 47 43 48 44 
<< m1 >>
rect 48 43 49 44 
<< m1 >>
rect 49 43 50 44 
<< m1 >>
rect 50 43 51 44 
<< m1 >>
rect 51 43 52 44 
<< m1 >>
rect 52 43 53 44 
<< m1 >>
rect 56 43 57 44 
<< m2 >>
rect 56 43 57 44 
<< m2c >>
rect 56 43 57 44 
<< m1 >>
rect 56 43 57 44 
<< m2 >>
rect 56 43 57 44 
<< m2 >>
rect 57 43 58 44 
<< m1 >>
rect 58 43 59 44 
<< m2 >>
rect 58 43 59 44 
<< m2 >>
rect 59 43 60 44 
<< m1 >>
rect 60 43 61 44 
<< m2 >>
rect 60 43 61 44 
<< m2 >>
rect 61 43 62 44 
<< m1 >>
rect 62 43 63 44 
<< m2 >>
rect 62 43 63 44 
<< m2c >>
rect 62 43 63 44 
<< m1 >>
rect 62 43 63 44 
<< m2 >>
rect 62 43 63 44 
<< m1 >>
rect 63 43 64 44 
<< m1 >>
rect 64 43 65 44 
<< m1 >>
rect 65 43 66 44 
<< m1 >>
rect 66 43 67 44 
<< m2 >>
rect 66 43 67 44 
<< m1 >>
rect 67 43 68 44 
<< m2 >>
rect 67 43 68 44 
<< m1 >>
rect 68 43 69 44 
<< m2 >>
rect 68 43 69 44 
<< m1 >>
rect 69 43 70 44 
<< m2 >>
rect 69 43 70 44 
<< m1 >>
rect 70 43 71 44 
<< m2 >>
rect 70 43 71 44 
<< m1 >>
rect 71 43 72 44 
<< m2 >>
rect 71 43 72 44 
<< m1 >>
rect 72 43 73 44 
<< m2 >>
rect 72 43 73 44 
<< m1 >>
rect 73 43 74 44 
<< m2 >>
rect 73 43 74 44 
<< m1 >>
rect 74 43 75 44 
<< m2 >>
rect 74 43 75 44 
<< m1 >>
rect 75 43 76 44 
<< m2 >>
rect 75 43 76 44 
<< m1 >>
rect 76 43 77 44 
<< m2 >>
rect 76 43 77 44 
<< m1 >>
rect 77 43 78 44 
<< m2 >>
rect 77 43 78 44 
<< m1 >>
rect 78 43 79 44 
<< m2 >>
rect 78 43 79 44 
<< m1 >>
rect 79 43 80 44 
<< m1 >>
rect 80 43 81 44 
<< m2 >>
rect 80 43 81 44 
<< m2c >>
rect 80 43 81 44 
<< m1 >>
rect 80 43 81 44 
<< m2 >>
rect 80 43 81 44 
<< m2 >>
rect 81 43 82 44 
<< m1 >>
rect 82 43 83 44 
<< m2 >>
rect 82 43 83 44 
<< m2 >>
rect 83 43 84 44 
<< m2 >>
rect 84 43 85 44 
<< m2 >>
rect 85 43 86 44 
<< m2 >>
rect 86 43 87 44 
<< m2 >>
rect 87 43 88 44 
<< m1 >>
rect 91 43 92 44 
<< m1 >>
rect 92 43 93 44 
<< m1 >>
rect 93 43 94 44 
<< m1 >>
rect 94 43 95 44 
<< m1 >>
rect 95 43 96 44 
<< m1 >>
rect 96 43 97 44 
<< m1 >>
rect 97 43 98 44 
<< m1 >>
rect 98 43 99 44 
<< m1 >>
rect 99 43 100 44 
<< m1 >>
rect 100 43 101 44 
<< m1 >>
rect 101 43 102 44 
<< m1 >>
rect 102 43 103 44 
<< m1 >>
rect 103 43 104 44 
<< m1 >>
rect 104 43 105 44 
<< m1 >>
rect 105 43 106 44 
<< m1 >>
rect 106 43 107 44 
<< m1 >>
rect 107 43 108 44 
<< m1 >>
rect 108 43 109 44 
<< m1 >>
rect 109 43 110 44 
<< m2 >>
rect 114 43 115 44 
<< m2 >>
rect 116 43 117 44 
<< m2 >>
rect 122 43 123 44 
<< m1 >>
rect 123 43 124 44 
<< m2 >>
rect 123 43 124 44 
<< m2c >>
rect 123 43 124 44 
<< m1 >>
rect 123 43 124 44 
<< m2 >>
rect 123 43 124 44 
<< m1 >>
rect 124 43 125 44 
<< m1 >>
rect 125 43 126 44 
<< m2 >>
rect 125 43 126 44 
<< m1 >>
rect 126 43 127 44 
<< m1 >>
rect 127 43 128 44 
<< m1 >>
rect 10 44 11 45 
<< m1 >>
rect 16 44 17 45 
<< m1 >>
rect 19 44 20 45 
<< m2 >>
rect 19 44 20 45 
<< m2 >>
rect 21 44 22 45 
<< m2 >>
rect 37 44 38 45 
<< m2 >>
rect 44 44 45 45 
<< m2 >>
rect 46 44 47 45 
<< m1 >>
rect 56 44 57 45 
<< m1 >>
rect 58 44 59 45 
<< m1 >>
rect 60 44 61 45 
<< m2 >>
rect 66 44 67 45 
<< m2 >>
rect 78 44 79 45 
<< m1 >>
rect 82 44 83 45 
<< m1 >>
rect 87 44 88 45 
<< m2 >>
rect 87 44 88 45 
<< m2c >>
rect 87 44 88 45 
<< m1 >>
rect 87 44 88 45 
<< m2 >>
rect 87 44 88 45 
<< m1 >>
rect 91 44 92 45 
<< m1 >>
rect 109 44 110 45 
<< m1 >>
rect 114 44 115 45 
<< m2 >>
rect 114 44 115 45 
<< m2c >>
rect 114 44 115 45 
<< m1 >>
rect 114 44 115 45 
<< m2 >>
rect 114 44 115 45 
<< m1 >>
rect 116 44 117 45 
<< m2 >>
rect 116 44 117 45 
<< m2c >>
rect 116 44 117 45 
<< m1 >>
rect 116 44 117 45 
<< m2 >>
rect 116 44 117 45 
<< m2 >>
rect 125 44 126 45 
<< m1 >>
rect 127 44 128 45 
<< m1 >>
rect 10 45 11 46 
<< m1 >>
rect 16 45 17 46 
<< m1 >>
rect 19 45 20 46 
<< m2 >>
rect 19 45 20 46 
<< m1 >>
rect 21 45 22 46 
<< m2 >>
rect 21 45 22 46 
<< m2c >>
rect 21 45 22 46 
<< m1 >>
rect 21 45 22 46 
<< m2 >>
rect 21 45 22 46 
<< m1 >>
rect 34 45 35 46 
<< m1 >>
rect 35 45 36 46 
<< m1 >>
rect 36 45 37 46 
<< m1 >>
rect 37 45 38 46 
<< m2 >>
rect 37 45 38 46 
<< m2c >>
rect 37 45 38 46 
<< m1 >>
rect 37 45 38 46 
<< m2 >>
rect 37 45 38 46 
<< m1 >>
rect 44 45 45 46 
<< m2 >>
rect 44 45 45 46 
<< m2c >>
rect 44 45 45 46 
<< m1 >>
rect 44 45 45 46 
<< m2 >>
rect 44 45 45 46 
<< m1 >>
rect 46 45 47 46 
<< m2 >>
rect 46 45 47 46 
<< m2c >>
rect 46 45 47 46 
<< m1 >>
rect 46 45 47 46 
<< m2 >>
rect 46 45 47 46 
<< m1 >>
rect 49 45 50 46 
<< m1 >>
rect 50 45 51 46 
<< m1 >>
rect 51 45 52 46 
<< m1 >>
rect 52 45 53 46 
<< m1 >>
rect 53 45 54 46 
<< m1 >>
rect 54 45 55 46 
<< m2 >>
rect 54 45 55 46 
<< m2c >>
rect 54 45 55 46 
<< m1 >>
rect 54 45 55 46 
<< m2 >>
rect 54 45 55 46 
<< m2 >>
rect 55 45 56 46 
<< m1 >>
rect 56 45 57 46 
<< m2 >>
rect 56 45 57 46 
<< m2 >>
rect 57 45 58 46 
<< m1 >>
rect 58 45 59 46 
<< m2 >>
rect 58 45 59 46 
<< m2 >>
rect 59 45 60 46 
<< m1 >>
rect 60 45 61 46 
<< m2 >>
rect 60 45 61 46 
<< m2 >>
rect 61 45 62 46 
<< m1 >>
rect 62 45 63 46 
<< m2 >>
rect 62 45 63 46 
<< m2c >>
rect 62 45 63 46 
<< m1 >>
rect 62 45 63 46 
<< m2 >>
rect 62 45 63 46 
<< m1 >>
rect 63 45 64 46 
<< m1 >>
rect 64 45 65 46 
<< m1 >>
rect 65 45 66 46 
<< m1 >>
rect 66 45 67 46 
<< m2 >>
rect 66 45 67 46 
<< m2c >>
rect 66 45 67 46 
<< m1 >>
rect 66 45 67 46 
<< m2 >>
rect 66 45 67 46 
<< m1 >>
rect 78 45 79 46 
<< m2 >>
rect 78 45 79 46 
<< m2c >>
rect 78 45 79 46 
<< m1 >>
rect 78 45 79 46 
<< m2 >>
rect 78 45 79 46 
<< m1 >>
rect 82 45 83 46 
<< m1 >>
rect 87 45 88 46 
<< m1 >>
rect 91 45 92 46 
<< m1 >>
rect 109 45 110 46 
<< m1 >>
rect 114 45 115 46 
<< m1 >>
rect 116 45 117 46 
<< m1 >>
rect 121 45 122 46 
<< m1 >>
rect 122 45 123 46 
<< m1 >>
rect 123 45 124 46 
<< m1 >>
rect 124 45 125 46 
<< m1 >>
rect 125 45 126 46 
<< m2 >>
rect 125 45 126 46 
<< m2c >>
rect 125 45 126 46 
<< m1 >>
rect 125 45 126 46 
<< m2 >>
rect 125 45 126 46 
<< m1 >>
rect 127 45 128 46 
<< m1 >>
rect 10 46 11 47 
<< m1 >>
rect 16 46 17 47 
<< m1 >>
rect 19 46 20 47 
<< m2 >>
rect 19 46 20 47 
<< m1 >>
rect 21 46 22 47 
<< m1 >>
rect 28 46 29 47 
<< m1 >>
rect 29 46 30 47 
<< m1 >>
rect 30 46 31 47 
<< m1 >>
rect 31 46 32 47 
<< m1 >>
rect 34 46 35 47 
<< m1 >>
rect 44 46 45 47 
<< m1 >>
rect 46 46 47 47 
<< m1 >>
rect 49 46 50 47 
<< m1 >>
rect 56 46 57 47 
<< m1 >>
rect 58 46 59 47 
<< m1 >>
rect 60 46 61 47 
<< m1 >>
rect 78 46 79 47 
<< m1 >>
rect 79 46 80 47 
<< m1 >>
rect 80 46 81 47 
<< m2 >>
rect 80 46 81 47 
<< m2c >>
rect 80 46 81 47 
<< m1 >>
rect 80 46 81 47 
<< m2 >>
rect 80 46 81 47 
<< m2 >>
rect 81 46 82 47 
<< m1 >>
rect 82 46 83 47 
<< m2 >>
rect 82 46 83 47 
<< m2 >>
rect 83 46 84 47 
<< m1 >>
rect 84 46 85 47 
<< m2 >>
rect 84 46 85 47 
<< m2c >>
rect 84 46 85 47 
<< m1 >>
rect 84 46 85 47 
<< m2 >>
rect 84 46 85 47 
<< m1 >>
rect 85 46 86 47 
<< m1 >>
rect 87 46 88 47 
<< m1 >>
rect 88 46 89 47 
<< m1 >>
rect 91 46 92 47 
<< m1 >>
rect 109 46 110 47 
<< m1 >>
rect 112 46 113 47 
<< m2 >>
rect 112 46 113 47 
<< m2c >>
rect 112 46 113 47 
<< m1 >>
rect 112 46 113 47 
<< m2 >>
rect 112 46 113 47 
<< m2 >>
rect 113 46 114 47 
<< m1 >>
rect 114 46 115 47 
<< m2 >>
rect 114 46 115 47 
<< m2 >>
rect 115 46 116 47 
<< m1 >>
rect 116 46 117 47 
<< m2 >>
rect 116 46 117 47 
<< m2c >>
rect 116 46 117 47 
<< m1 >>
rect 116 46 117 47 
<< m2 >>
rect 116 46 117 47 
<< m1 >>
rect 121 46 122 47 
<< m1 >>
rect 127 46 128 47 
<< m1 >>
rect 10 47 11 48 
<< m1 >>
rect 16 47 17 48 
<< m1 >>
rect 19 47 20 48 
<< m2 >>
rect 19 47 20 48 
<< m1 >>
rect 21 47 22 48 
<< m1 >>
rect 28 47 29 48 
<< m1 >>
rect 31 47 32 48 
<< m1 >>
rect 34 47 35 48 
<< m1 >>
rect 44 47 45 48 
<< m1 >>
rect 46 47 47 48 
<< m1 >>
rect 49 47 50 48 
<< m1 >>
rect 56 47 57 48 
<< m1 >>
rect 58 47 59 48 
<< m1 >>
rect 60 47 61 48 
<< m1 >>
rect 82 47 83 48 
<< m1 >>
rect 85 47 86 48 
<< m1 >>
rect 88 47 89 48 
<< m1 >>
rect 91 47 92 48 
<< m1 >>
rect 109 47 110 48 
<< m1 >>
rect 112 47 113 48 
<< m1 >>
rect 114 47 115 48 
<< m1 >>
rect 121 47 122 48 
<< m1 >>
rect 127 47 128 48 
<< m1 >>
rect 10 48 11 49 
<< pdiffusion >>
rect 12 48 13 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< m1 >>
rect 16 48 17 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< m1 >>
rect 19 48 20 49 
<< m2 >>
rect 19 48 20 49 
<< m1 >>
rect 21 48 22 49 
<< m1 >>
rect 28 48 29 49 
<< pdiffusion >>
rect 30 48 31 49 
<< m1 >>
rect 31 48 32 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< m1 >>
rect 34 48 35 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< m1 >>
rect 44 48 45 49 
<< m1 >>
rect 46 48 47 49 
<< pdiffusion >>
rect 48 48 49 49 
<< m1 >>
rect 49 48 50 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 56 48 57 49 
<< m1 >>
rect 58 48 59 49 
<< m1 >>
rect 60 48 61 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< m1 >>
rect 82 48 83 49 
<< pdiffusion >>
rect 84 48 85 49 
<< m1 >>
rect 85 48 86 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< m1 >>
rect 88 48 89 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< pdiffusion >>
rect 102 48 103 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< m1 >>
rect 109 48 110 49 
<< m1 >>
rect 112 48 113 49 
<< m1 >>
rect 114 48 115 49 
<< pdiffusion >>
rect 120 48 121 49 
<< m1 >>
rect 121 48 122 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< m1 >>
rect 127 48 128 49 
<< m1 >>
rect 10 49 11 50 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< m1 >>
rect 19 49 20 50 
<< m2 >>
rect 19 49 20 50 
<< m1 >>
rect 21 49 22 50 
<< m1 >>
rect 28 49 29 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< m1 >>
rect 44 49 45 50 
<< m1 >>
rect 46 49 47 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 56 49 57 50 
<< m1 >>
rect 58 49 59 50 
<< m1 >>
rect 60 49 61 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< m1 >>
rect 82 49 83 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< m1 >>
rect 109 49 110 50 
<< m1 >>
rect 112 49 113 50 
<< m1 >>
rect 114 49 115 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< m1 >>
rect 127 49 128 50 
<< m1 >>
rect 10 50 11 51 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< m1 >>
rect 19 50 20 51 
<< m2 >>
rect 19 50 20 51 
<< m1 >>
rect 21 50 22 51 
<< m1 >>
rect 28 50 29 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< m1 >>
rect 44 50 45 51 
<< m1 >>
rect 46 50 47 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 56 50 57 51 
<< m1 >>
rect 58 50 59 51 
<< m1 >>
rect 60 50 61 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< m1 >>
rect 82 50 83 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< m1 >>
rect 109 50 110 51 
<< m1 >>
rect 112 50 113 51 
<< m1 >>
rect 114 50 115 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< m1 >>
rect 127 50 128 51 
<< m1 >>
rect 10 51 11 52 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< m1 >>
rect 19 51 20 52 
<< m2 >>
rect 19 51 20 52 
<< m1 >>
rect 21 51 22 52 
<< m1 >>
rect 28 51 29 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< m1 >>
rect 44 51 45 52 
<< m1 >>
rect 46 51 47 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 56 51 57 52 
<< m1 >>
rect 58 51 59 52 
<< m1 >>
rect 60 51 61 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< m1 >>
rect 82 51 83 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< m1 >>
rect 109 51 110 52 
<< m1 >>
rect 112 51 113 52 
<< m1 >>
rect 114 51 115 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< m1 >>
rect 127 51 128 52 
<< m1 >>
rect 10 52 11 53 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< m1 >>
rect 19 52 20 53 
<< m2 >>
rect 19 52 20 53 
<< m1 >>
rect 21 52 22 53 
<< m1 >>
rect 28 52 29 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< m1 >>
rect 44 52 45 53 
<< m1 >>
rect 46 52 47 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 56 52 57 53 
<< m1 >>
rect 58 52 59 53 
<< m1 >>
rect 60 52 61 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< m1 >>
rect 82 52 83 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< m1 >>
rect 109 52 110 53 
<< m1 >>
rect 112 52 113 53 
<< m1 >>
rect 114 52 115 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< m1 >>
rect 127 52 128 53 
<< m1 >>
rect 10 53 11 54 
<< pdiffusion >>
rect 12 53 13 54 
<< m1 >>
rect 13 53 14 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< m1 >>
rect 19 53 20 54 
<< m2 >>
rect 19 53 20 54 
<< m1 >>
rect 21 53 22 54 
<< m1 >>
rect 28 53 29 54 
<< pdiffusion >>
rect 30 53 31 54 
<< m1 >>
rect 31 53 32 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< m1 >>
rect 34 53 35 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< m1 >>
rect 44 53 45 54 
<< m1 >>
rect 46 53 47 54 
<< pdiffusion >>
rect 48 53 49 54 
<< m1 >>
rect 49 53 50 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 56 53 57 54 
<< m1 >>
rect 58 53 59 54 
<< m1 >>
rect 60 53 61 54 
<< pdiffusion >>
rect 66 53 67 54 
<< m1 >>
rect 67 53 68 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< m1 >>
rect 82 53 83 54 
<< pdiffusion >>
rect 84 53 85 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< m1 >>
rect 88 53 89 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< pdiffusion >>
rect 102 53 103 54 
<< m1 >>
rect 103 53 104 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< m1 >>
rect 106 53 107 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< m1 >>
rect 109 53 110 54 
<< m1 >>
rect 112 53 113 54 
<< m1 >>
rect 114 53 115 54 
<< pdiffusion >>
rect 120 53 121 54 
<< m1 >>
rect 121 53 122 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< m1 >>
rect 124 53 125 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< m1 >>
rect 127 53 128 54 
<< m1 >>
rect 10 54 11 55 
<< m1 >>
rect 13 54 14 55 
<< m1 >>
rect 19 54 20 55 
<< m2 >>
rect 19 54 20 55 
<< m1 >>
rect 21 54 22 55 
<< m1 >>
rect 28 54 29 55 
<< m1 >>
rect 31 54 32 55 
<< m1 >>
rect 34 54 35 55 
<< m1 >>
rect 44 54 45 55 
<< m1 >>
rect 46 54 47 55 
<< m1 >>
rect 49 54 50 55 
<< m1 >>
rect 56 54 57 55 
<< m1 >>
rect 58 54 59 55 
<< m1 >>
rect 60 54 61 55 
<< m1 >>
rect 67 54 68 55 
<< m1 >>
rect 82 54 83 55 
<< m1 >>
rect 88 54 89 55 
<< m1 >>
rect 91 54 92 55 
<< m1 >>
rect 103 54 104 55 
<< m1 >>
rect 106 54 107 55 
<< m1 >>
rect 109 54 110 55 
<< m2 >>
rect 109 54 110 55 
<< m2c >>
rect 109 54 110 55 
<< m1 >>
rect 109 54 110 55 
<< m2 >>
rect 109 54 110 55 
<< m1 >>
rect 112 54 113 55 
<< m2 >>
rect 112 54 113 55 
<< m2c >>
rect 112 54 113 55 
<< m1 >>
rect 112 54 113 55 
<< m2 >>
rect 112 54 113 55 
<< m1 >>
rect 114 54 115 55 
<< m2 >>
rect 114 54 115 55 
<< m2c >>
rect 114 54 115 55 
<< m1 >>
rect 114 54 115 55 
<< m2 >>
rect 114 54 115 55 
<< m1 >>
rect 121 54 122 55 
<< m1 >>
rect 124 54 125 55 
<< m1 >>
rect 127 54 128 55 
<< m1 >>
rect 10 55 11 56 
<< m1 >>
rect 13 55 14 56 
<< m1 >>
rect 19 55 20 56 
<< m2 >>
rect 19 55 20 56 
<< m1 >>
rect 21 55 22 56 
<< m1 >>
rect 28 55 29 56 
<< m1 >>
rect 31 55 32 56 
<< m1 >>
rect 34 55 35 56 
<< m1 >>
rect 44 55 45 56 
<< m1 >>
rect 46 55 47 56 
<< m1 >>
rect 49 55 50 56 
<< m1 >>
rect 56 55 57 56 
<< m1 >>
rect 58 55 59 56 
<< m1 >>
rect 60 55 61 56 
<< m1 >>
rect 67 55 68 56 
<< m1 >>
rect 82 55 83 56 
<< m1 >>
rect 88 55 89 56 
<< m1 >>
rect 89 55 90 56 
<< m1 >>
rect 90 55 91 56 
<< m1 >>
rect 91 55 92 56 
<< m1 >>
rect 103 55 104 56 
<< m1 >>
rect 106 55 107 56 
<< m2 >>
rect 109 55 110 56 
<< m2 >>
rect 112 55 113 56 
<< m2 >>
rect 114 55 115 56 
<< m1 >>
rect 121 55 122 56 
<< m1 >>
rect 122 55 123 56 
<< m2 >>
rect 122 55 123 56 
<< m2c >>
rect 122 55 123 56 
<< m1 >>
rect 122 55 123 56 
<< m2 >>
rect 122 55 123 56 
<< m2 >>
rect 123 55 124 56 
<< m1 >>
rect 124 55 125 56 
<< m1 >>
rect 127 55 128 56 
<< m1 >>
rect 10 56 11 57 
<< m1 >>
rect 13 56 14 57 
<< m1 >>
rect 14 56 15 57 
<< m1 >>
rect 15 56 16 57 
<< m1 >>
rect 16 56 17 57 
<< m1 >>
rect 17 56 18 57 
<< m1 >>
rect 18 56 19 57 
<< m1 >>
rect 19 56 20 57 
<< m2 >>
rect 19 56 20 57 
<< m1 >>
rect 21 56 22 57 
<< m1 >>
rect 28 56 29 57 
<< m1 >>
rect 31 56 32 57 
<< m1 >>
rect 34 56 35 57 
<< m1 >>
rect 44 56 45 57 
<< m1 >>
rect 46 56 47 57 
<< m2 >>
rect 46 56 47 57 
<< m2c >>
rect 46 56 47 57 
<< m1 >>
rect 46 56 47 57 
<< m2 >>
rect 46 56 47 57 
<< m1 >>
rect 49 56 50 57 
<< m1 >>
rect 50 56 51 57 
<< m1 >>
rect 51 56 52 57 
<< m1 >>
rect 52 56 53 57 
<< m1 >>
rect 53 56 54 57 
<< m1 >>
rect 54 56 55 57 
<< m2 >>
rect 54 56 55 57 
<< m2c >>
rect 54 56 55 57 
<< m1 >>
rect 54 56 55 57 
<< m2 >>
rect 54 56 55 57 
<< m1 >>
rect 56 56 57 57 
<< m2 >>
rect 56 56 57 57 
<< m2c >>
rect 56 56 57 57 
<< m1 >>
rect 56 56 57 57 
<< m2 >>
rect 56 56 57 57 
<< m1 >>
rect 58 56 59 57 
<< m2 >>
rect 58 56 59 57 
<< m2c >>
rect 58 56 59 57 
<< m1 >>
rect 58 56 59 57 
<< m2 >>
rect 58 56 59 57 
<< m1 >>
rect 60 56 61 57 
<< m2 >>
rect 60 56 61 57 
<< m2c >>
rect 60 56 61 57 
<< m1 >>
rect 60 56 61 57 
<< m2 >>
rect 60 56 61 57 
<< m1 >>
rect 67 56 68 57 
<< m1 >>
rect 68 56 69 57 
<< m1 >>
rect 69 56 70 57 
<< m1 >>
rect 70 56 71 57 
<< m1 >>
rect 71 56 72 57 
<< m1 >>
rect 72 56 73 57 
<< m1 >>
rect 73 56 74 57 
<< m1 >>
rect 74 56 75 57 
<< m1 >>
rect 75 56 76 57 
<< m1 >>
rect 76 56 77 57 
<< m1 >>
rect 77 56 78 57 
<< m1 >>
rect 78 56 79 57 
<< m1 >>
rect 79 56 80 57 
<< m1 >>
rect 80 56 81 57 
<< m1 >>
rect 81 56 82 57 
<< m1 >>
rect 82 56 83 57 
<< m1 >>
rect 103 56 104 57 
<< m1 >>
rect 106 56 107 57 
<< m1 >>
rect 107 56 108 57 
<< m1 >>
rect 108 56 109 57 
<< m1 >>
rect 109 56 110 57 
<< m2 >>
rect 109 56 110 57 
<< m1 >>
rect 110 56 111 57 
<< m1 >>
rect 111 56 112 57 
<< m1 >>
rect 112 56 113 57 
<< m2 >>
rect 112 56 113 57 
<< m1 >>
rect 113 56 114 57 
<< m1 >>
rect 114 56 115 57 
<< m2 >>
rect 114 56 115 57 
<< m1 >>
rect 115 56 116 57 
<< m1 >>
rect 116 56 117 57 
<< m1 >>
rect 117 56 118 57 
<< m1 >>
rect 118 56 119 57 
<< m2 >>
rect 118 56 119 57 
<< m2c >>
rect 118 56 119 57 
<< m1 >>
rect 118 56 119 57 
<< m2 >>
rect 118 56 119 57 
<< m2 >>
rect 123 56 124 57 
<< m1 >>
rect 124 56 125 57 
<< m2 >>
rect 124 56 125 57 
<< m2 >>
rect 125 56 126 57 
<< m1 >>
rect 126 56 127 57 
<< m2 >>
rect 126 56 127 57 
<< m2c >>
rect 126 56 127 57 
<< m1 >>
rect 126 56 127 57 
<< m2 >>
rect 126 56 127 57 
<< m1 >>
rect 127 56 128 57 
<< m1 >>
rect 10 57 11 58 
<< m2 >>
rect 19 57 20 58 
<< m1 >>
rect 21 57 22 58 
<< m1 >>
rect 28 57 29 58 
<< m1 >>
rect 31 57 32 58 
<< m1 >>
rect 34 57 35 58 
<< m1 >>
rect 44 57 45 58 
<< m2 >>
rect 46 57 47 58 
<< m2 >>
rect 54 57 55 58 
<< m2 >>
rect 56 57 57 58 
<< m2 >>
rect 58 57 59 58 
<< m2 >>
rect 60 57 61 58 
<< m1 >>
rect 103 57 104 58 
<< m2 >>
rect 109 57 110 58 
<< m2 >>
rect 112 57 113 58 
<< m2 >>
rect 114 57 115 58 
<< m2 >>
rect 118 57 119 58 
<< m1 >>
rect 124 57 125 58 
<< m1 >>
rect 10 58 11 59 
<< m1 >>
rect 19 58 20 59 
<< m2 >>
rect 19 58 20 59 
<< m2c >>
rect 19 58 20 59 
<< m1 >>
rect 19 58 20 59 
<< m2 >>
rect 19 58 20 59 
<< m1 >>
rect 21 58 22 59 
<< m1 >>
rect 28 58 29 59 
<< m1 >>
rect 31 58 32 59 
<< m1 >>
rect 34 58 35 59 
<< m1 >>
rect 44 58 45 59 
<< m1 >>
rect 46 58 47 59 
<< m2 >>
rect 46 58 47 59 
<< m1 >>
rect 47 58 48 59 
<< m1 >>
rect 48 58 49 59 
<< m1 >>
rect 49 58 50 59 
<< m1 >>
rect 50 58 51 59 
<< m1 >>
rect 51 58 52 59 
<< m1 >>
rect 52 58 53 59 
<< m1 >>
rect 53 58 54 59 
<< m1 >>
rect 54 58 55 59 
<< m2 >>
rect 54 58 55 59 
<< m1 >>
rect 55 58 56 59 
<< m1 >>
rect 56 58 57 59 
<< m2 >>
rect 56 58 57 59 
<< m1 >>
rect 57 58 58 59 
<< m1 >>
rect 58 58 59 59 
<< m2 >>
rect 58 58 59 59 
<< m1 >>
rect 59 58 60 59 
<< m1 >>
rect 60 58 61 59 
<< m2 >>
rect 60 58 61 59 
<< m1 >>
rect 61 58 62 59 
<< m1 >>
rect 62 58 63 59 
<< m2 >>
rect 62 58 63 59 
<< m2c >>
rect 62 58 63 59 
<< m1 >>
rect 62 58 63 59 
<< m2 >>
rect 62 58 63 59 
<< m2 >>
rect 63 58 64 59 
<< m1 >>
rect 64 58 65 59 
<< m2 >>
rect 64 58 65 59 
<< m1 >>
rect 65 58 66 59 
<< m2 >>
rect 65 58 66 59 
<< m1 >>
rect 66 58 67 59 
<< m2 >>
rect 66 58 67 59 
<< m1 >>
rect 67 58 68 59 
<< m2 >>
rect 67 58 68 59 
<< m1 >>
rect 68 58 69 59 
<< m2 >>
rect 68 58 69 59 
<< m1 >>
rect 69 58 70 59 
<< m2 >>
rect 69 58 70 59 
<< m1 >>
rect 70 58 71 59 
<< m2 >>
rect 70 58 71 59 
<< m1 >>
rect 71 58 72 59 
<< m2 >>
rect 71 58 72 59 
<< m1 >>
rect 72 58 73 59 
<< m2 >>
rect 72 58 73 59 
<< m1 >>
rect 73 58 74 59 
<< m2 >>
rect 73 58 74 59 
<< m1 >>
rect 74 58 75 59 
<< m2 >>
rect 74 58 75 59 
<< m1 >>
rect 75 58 76 59 
<< m2 >>
rect 75 58 76 59 
<< m1 >>
rect 76 58 77 59 
<< m2 >>
rect 76 58 77 59 
<< m1 >>
rect 77 58 78 59 
<< m2 >>
rect 77 58 78 59 
<< m1 >>
rect 78 58 79 59 
<< m2 >>
rect 78 58 79 59 
<< m1 >>
rect 79 58 80 59 
<< m2 >>
rect 79 58 80 59 
<< m1 >>
rect 80 58 81 59 
<< m2 >>
rect 80 58 81 59 
<< m1 >>
rect 81 58 82 59 
<< m2 >>
rect 81 58 82 59 
<< m1 >>
rect 82 58 83 59 
<< m2 >>
rect 82 58 83 59 
<< m1 >>
rect 83 58 84 59 
<< m2 >>
rect 83 58 84 59 
<< m1 >>
rect 84 58 85 59 
<< m2 >>
rect 84 58 85 59 
<< m1 >>
rect 85 58 86 59 
<< m2 >>
rect 85 58 86 59 
<< m1 >>
rect 86 58 87 59 
<< m2 >>
rect 86 58 87 59 
<< m1 >>
rect 87 58 88 59 
<< m2 >>
rect 87 58 88 59 
<< m1 >>
rect 88 58 89 59 
<< m2 >>
rect 88 58 89 59 
<< m1 >>
rect 89 58 90 59 
<< m2 >>
rect 89 58 90 59 
<< m1 >>
rect 90 58 91 59 
<< m2 >>
rect 90 58 91 59 
<< m1 >>
rect 91 58 92 59 
<< m2 >>
rect 91 58 92 59 
<< m1 >>
rect 92 58 93 59 
<< m2 >>
rect 92 58 93 59 
<< m1 >>
rect 93 58 94 59 
<< m2 >>
rect 93 58 94 59 
<< m1 >>
rect 94 58 95 59 
<< m2 >>
rect 94 58 95 59 
<< m1 >>
rect 95 58 96 59 
<< m2 >>
rect 95 58 96 59 
<< m1 >>
rect 96 58 97 59 
<< m2 >>
rect 96 58 97 59 
<< m1 >>
rect 97 58 98 59 
<< m2 >>
rect 97 58 98 59 
<< m1 >>
rect 98 58 99 59 
<< m2 >>
rect 98 58 99 59 
<< m1 >>
rect 99 58 100 59 
<< m2 >>
rect 99 58 100 59 
<< m1 >>
rect 100 58 101 59 
<< m2 >>
rect 100 58 101 59 
<< m1 >>
rect 101 58 102 59 
<< m2 >>
rect 101 58 102 59 
<< m1 >>
rect 102 58 103 59 
<< m2 >>
rect 102 58 103 59 
<< m1 >>
rect 103 58 104 59 
<< m2 >>
rect 103 58 104 59 
<< m2 >>
rect 104 58 105 59 
<< m1 >>
rect 105 58 106 59 
<< m2 >>
rect 105 58 106 59 
<< m2c >>
rect 105 58 106 59 
<< m1 >>
rect 105 58 106 59 
<< m2 >>
rect 105 58 106 59 
<< m1 >>
rect 106 58 107 59 
<< m1 >>
rect 107 58 108 59 
<< m1 >>
rect 108 58 109 59 
<< m1 >>
rect 109 58 110 59 
<< m2 >>
rect 109 58 110 59 
<< m1 >>
rect 110 58 111 59 
<< m1 >>
rect 111 58 112 59 
<< m1 >>
rect 112 58 113 59 
<< m2 >>
rect 112 58 113 59 
<< m1 >>
rect 113 58 114 59 
<< m1 >>
rect 114 58 115 59 
<< m2 >>
rect 114 58 115 59 
<< m1 >>
rect 115 58 116 59 
<< m1 >>
rect 116 58 117 59 
<< m1 >>
rect 117 58 118 59 
<< m1 >>
rect 118 58 119 59 
<< m2 >>
rect 118 58 119 59 
<< m1 >>
rect 119 58 120 59 
<< m1 >>
rect 120 58 121 59 
<< m1 >>
rect 121 58 122 59 
<< m1 >>
rect 122 58 123 59 
<< m1 >>
rect 123 58 124 59 
<< m1 >>
rect 124 58 125 59 
<< m1 >>
rect 10 59 11 60 
<< m1 >>
rect 19 59 20 60 
<< m1 >>
rect 21 59 22 60 
<< m1 >>
rect 28 59 29 60 
<< m1 >>
rect 31 59 32 60 
<< m1 >>
rect 34 59 35 60 
<< m1 >>
rect 35 59 36 60 
<< m1 >>
rect 36 59 37 60 
<< m1 >>
rect 37 59 38 60 
<< m1 >>
rect 38 59 39 60 
<< m2 >>
rect 38 59 39 60 
<< m2c >>
rect 38 59 39 60 
<< m1 >>
rect 38 59 39 60 
<< m2 >>
rect 38 59 39 60 
<< m1 >>
rect 44 59 45 60 
<< m2 >>
rect 44 59 45 60 
<< m2c >>
rect 44 59 45 60 
<< m1 >>
rect 44 59 45 60 
<< m2 >>
rect 44 59 45 60 
<< m1 >>
rect 46 59 47 60 
<< m2 >>
rect 46 59 47 60 
<< m2 >>
rect 54 59 55 60 
<< m2 >>
rect 56 59 57 60 
<< m2 >>
rect 58 59 59 60 
<< m2 >>
rect 60 59 61 60 
<< m1 >>
rect 64 59 65 60 
<< m2 >>
rect 109 59 110 60 
<< m2 >>
rect 112 59 113 60 
<< m2 >>
rect 114 59 115 60 
<< m2 >>
rect 118 59 119 60 
<< m1 >>
rect 10 60 11 61 
<< m1 >>
rect 19 60 20 61 
<< m1 >>
rect 21 60 22 61 
<< m1 >>
rect 28 60 29 61 
<< m1 >>
rect 31 60 32 61 
<< m2 >>
rect 38 60 39 61 
<< m2 >>
rect 40 60 41 61 
<< m2 >>
rect 41 60 42 61 
<< m2 >>
rect 42 60 43 61 
<< m2 >>
rect 43 60 44 61 
<< m2 >>
rect 44 60 45 61 
<< m1 >>
rect 46 60 47 61 
<< m2 >>
rect 46 60 47 61 
<< m1 >>
rect 54 60 55 61 
<< m2 >>
rect 54 60 55 61 
<< m2c >>
rect 54 60 55 61 
<< m1 >>
rect 54 60 55 61 
<< m2 >>
rect 54 60 55 61 
<< m1 >>
rect 56 60 57 61 
<< m2 >>
rect 56 60 57 61 
<< m2c >>
rect 56 60 57 61 
<< m1 >>
rect 56 60 57 61 
<< m2 >>
rect 56 60 57 61 
<< m1 >>
rect 58 60 59 61 
<< m2 >>
rect 58 60 59 61 
<< m2c >>
rect 58 60 59 61 
<< m1 >>
rect 58 60 59 61 
<< m2 >>
rect 58 60 59 61 
<< m1 >>
rect 60 60 61 61 
<< m2 >>
rect 60 60 61 61 
<< m2c >>
rect 60 60 61 61 
<< m1 >>
rect 60 60 61 61 
<< m2 >>
rect 60 60 61 61 
<< m1 >>
rect 61 60 62 61 
<< m1 >>
rect 62 60 63 61 
<< m2 >>
rect 62 60 63 61 
<< m2c >>
rect 62 60 63 61 
<< m1 >>
rect 62 60 63 61 
<< m2 >>
rect 62 60 63 61 
<< m2 >>
rect 63 60 64 61 
<< m1 >>
rect 64 60 65 61 
<< m2 >>
rect 64 60 65 61 
<< m2 >>
rect 65 60 66 61 
<< m1 >>
rect 66 60 67 61 
<< m2 >>
rect 66 60 67 61 
<< m2c >>
rect 66 60 67 61 
<< m1 >>
rect 66 60 67 61 
<< m2 >>
rect 66 60 67 61 
<< m1 >>
rect 67 60 68 61 
<< m1 >>
rect 68 60 69 61 
<< m1 >>
rect 69 60 70 61 
<< m1 >>
rect 70 60 71 61 
<< m1 >>
rect 109 60 110 61 
<< m2 >>
rect 109 60 110 61 
<< m2c >>
rect 109 60 110 61 
<< m1 >>
rect 109 60 110 61 
<< m2 >>
rect 109 60 110 61 
<< m1 >>
rect 112 60 113 61 
<< m2 >>
rect 112 60 113 61 
<< m2c >>
rect 112 60 113 61 
<< m1 >>
rect 112 60 113 61 
<< m2 >>
rect 112 60 113 61 
<< m1 >>
rect 114 60 115 61 
<< m2 >>
rect 114 60 115 61 
<< m2c >>
rect 114 60 115 61 
<< m1 >>
rect 114 60 115 61 
<< m2 >>
rect 114 60 115 61 
<< m1 >>
rect 118 60 119 61 
<< m2 >>
rect 118 60 119 61 
<< m2c >>
rect 118 60 119 61 
<< m1 >>
rect 118 60 119 61 
<< m2 >>
rect 118 60 119 61 
<< m1 >>
rect 10 61 11 62 
<< m1 >>
rect 19 61 20 62 
<< m1 >>
rect 21 61 22 62 
<< m1 >>
rect 28 61 29 62 
<< m1 >>
rect 31 61 32 62 
<< m1 >>
rect 32 61 33 62 
<< m1 >>
rect 33 61 34 62 
<< m1 >>
rect 34 61 35 62 
<< m1 >>
rect 35 61 36 62 
<< m1 >>
rect 36 61 37 62 
<< m1 >>
rect 37 61 38 62 
<< m1 >>
rect 38 61 39 62 
<< m2 >>
rect 38 61 39 62 
<< m1 >>
rect 39 61 40 62 
<< m1 >>
rect 40 61 41 62 
<< m2 >>
rect 40 61 41 62 
<< m1 >>
rect 41 61 42 62 
<< m1 >>
rect 42 61 43 62 
<< m1 >>
rect 43 61 44 62 
<< m1 >>
rect 44 61 45 62 
<< m1 >>
rect 46 61 47 62 
<< m2 >>
rect 46 61 47 62 
<< m1 >>
rect 54 61 55 62 
<< m1 >>
rect 56 61 57 62 
<< m1 >>
rect 58 61 59 62 
<< m1 >>
rect 64 61 65 62 
<< m1 >>
rect 70 61 71 62 
<< m1 >>
rect 100 61 101 62 
<< m1 >>
rect 101 61 102 62 
<< m2 >>
rect 101 61 102 62 
<< m2c >>
rect 101 61 102 62 
<< m1 >>
rect 101 61 102 62 
<< m2 >>
rect 101 61 102 62 
<< m2 >>
rect 102 61 103 62 
<< m2 >>
rect 103 61 104 62 
<< m2 >>
rect 104 61 105 62 
<< m2 >>
rect 105 61 106 62 
<< m1 >>
rect 109 61 110 62 
<< m1 >>
rect 112 61 113 62 
<< m1 >>
rect 114 61 115 62 
<< m1 >>
rect 118 61 119 62 
<< m1 >>
rect 10 62 11 63 
<< m1 >>
rect 19 62 20 63 
<< m1 >>
rect 21 62 22 63 
<< m1 >>
rect 28 62 29 63 
<< m2 >>
rect 38 62 39 63 
<< m2 >>
rect 40 62 41 63 
<< m1 >>
rect 44 62 45 63 
<< m1 >>
rect 46 62 47 63 
<< m2 >>
rect 46 62 47 63 
<< m1 >>
rect 54 62 55 63 
<< m1 >>
rect 56 62 57 63 
<< m2 >>
rect 56 62 57 63 
<< m2c >>
rect 56 62 57 63 
<< m1 >>
rect 56 62 57 63 
<< m2 >>
rect 56 62 57 63 
<< m2 >>
rect 57 62 58 63 
<< m1 >>
rect 58 62 59 63 
<< m2 >>
rect 58 62 59 63 
<< m2 >>
rect 59 62 60 63 
<< m1 >>
rect 60 62 61 63 
<< m2 >>
rect 60 62 61 63 
<< m2c >>
rect 60 62 61 63 
<< m1 >>
rect 60 62 61 63 
<< m2 >>
rect 60 62 61 63 
<< m1 >>
rect 61 62 62 63 
<< m1 >>
rect 62 62 63 63 
<< m2 >>
rect 62 62 63 63 
<< m2c >>
rect 62 62 63 63 
<< m1 >>
rect 62 62 63 63 
<< m2 >>
rect 62 62 63 63 
<< m2 >>
rect 63 62 64 63 
<< m1 >>
rect 64 62 65 63 
<< m1 >>
rect 70 62 71 63 
<< m1 >>
rect 100 62 101 63 
<< m1 >>
rect 103 62 104 63 
<< m1 >>
rect 104 62 105 63 
<< m1 >>
rect 105 62 106 63 
<< m2 >>
rect 105 62 106 63 
<< m1 >>
rect 106 62 107 63 
<< m1 >>
rect 107 62 108 63 
<< m2 >>
rect 107 62 108 63 
<< m2c >>
rect 107 62 108 63 
<< m1 >>
rect 107 62 108 63 
<< m2 >>
rect 107 62 108 63 
<< m2 >>
rect 108 62 109 63 
<< m1 >>
rect 109 62 110 63 
<< m2 >>
rect 109 62 110 63 
<< m2 >>
rect 110 62 111 63 
<< m1 >>
rect 111 62 112 63 
<< m2 >>
rect 111 62 112 63 
<< m2c >>
rect 111 62 112 63 
<< m1 >>
rect 111 62 112 63 
<< m2 >>
rect 111 62 112 63 
<< m1 >>
rect 112 62 113 63 
<< m1 >>
rect 114 62 115 63 
<< m1 >>
rect 118 62 119 63 
<< m1 >>
rect 10 63 11 64 
<< m1 >>
rect 13 63 14 64 
<< m1 >>
rect 14 63 15 64 
<< m1 >>
rect 15 63 16 64 
<< m1 >>
rect 16 63 17 64 
<< m1 >>
rect 17 63 18 64 
<< m2 >>
rect 17 63 18 64 
<< m2c >>
rect 17 63 18 64 
<< m1 >>
rect 17 63 18 64 
<< m2 >>
rect 17 63 18 64 
<< m2 >>
rect 18 63 19 64 
<< m1 >>
rect 19 63 20 64 
<< m2 >>
rect 19 63 20 64 
<< m2 >>
rect 20 63 21 64 
<< m1 >>
rect 21 63 22 64 
<< m2 >>
rect 21 63 22 64 
<< m2 >>
rect 22 63 23 64 
<< m1 >>
rect 23 63 24 64 
<< m2 >>
rect 23 63 24 64 
<< m2c >>
rect 23 63 24 64 
<< m1 >>
rect 23 63 24 64 
<< m2 >>
rect 23 63 24 64 
<< m1 >>
rect 24 63 25 64 
<< m1 >>
rect 25 63 26 64 
<< m1 >>
rect 26 63 27 64 
<< m2 >>
rect 26 63 27 64 
<< m2c >>
rect 26 63 27 64 
<< m1 >>
rect 26 63 27 64 
<< m2 >>
rect 26 63 27 64 
<< m2 >>
rect 27 63 28 64 
<< m1 >>
rect 28 63 29 64 
<< m1 >>
rect 34 63 35 64 
<< m1 >>
rect 35 63 36 64 
<< m1 >>
rect 36 63 37 64 
<< m1 >>
rect 37 63 38 64 
<< m1 >>
rect 38 63 39 64 
<< m2 >>
rect 38 63 39 64 
<< m1 >>
rect 39 63 40 64 
<< m1 >>
rect 40 63 41 64 
<< m2 >>
rect 40 63 41 64 
<< m1 >>
rect 41 63 42 64 
<< m1 >>
rect 42 63 43 64 
<< m2 >>
rect 42 63 43 64 
<< m2c >>
rect 42 63 43 64 
<< m1 >>
rect 42 63 43 64 
<< m2 >>
rect 42 63 43 64 
<< m2 >>
rect 43 63 44 64 
<< m1 >>
rect 44 63 45 64 
<< m2 >>
rect 44 63 45 64 
<< m2 >>
rect 45 63 46 64 
<< m1 >>
rect 46 63 47 64 
<< m2 >>
rect 46 63 47 64 
<< m1 >>
rect 49 63 50 64 
<< m1 >>
rect 50 63 51 64 
<< m1 >>
rect 51 63 52 64 
<< m1 >>
rect 52 63 53 64 
<< m2 >>
rect 52 63 53 64 
<< m2c >>
rect 52 63 53 64 
<< m1 >>
rect 52 63 53 64 
<< m2 >>
rect 52 63 53 64 
<< m2 >>
rect 53 63 54 64 
<< m1 >>
rect 54 63 55 64 
<< m2 >>
rect 54 63 55 64 
<< m1 >>
rect 58 63 59 64 
<< m2 >>
rect 63 63 64 64 
<< m1 >>
rect 64 63 65 64 
<< m1 >>
rect 70 63 71 64 
<< m1 >>
rect 100 63 101 64 
<< m1 >>
rect 103 63 104 64 
<< m2 >>
rect 105 63 106 64 
<< m1 >>
rect 109 63 110 64 
<< m1 >>
rect 114 63 115 64 
<< m1 >>
rect 118 63 119 64 
<< m1 >>
rect 10 64 11 65 
<< m1 >>
rect 13 64 14 65 
<< m1 >>
rect 19 64 20 65 
<< m1 >>
rect 21 64 22 65 
<< m2 >>
rect 27 64 28 65 
<< m1 >>
rect 28 64 29 65 
<< m1 >>
rect 34 64 35 65 
<< m2 >>
rect 38 64 39 65 
<< m2 >>
rect 40 64 41 65 
<< m1 >>
rect 44 64 45 65 
<< m1 >>
rect 46 64 47 65 
<< m1 >>
rect 49 64 50 65 
<< m1 >>
rect 54 64 55 65 
<< m2 >>
rect 54 64 55 65 
<< m1 >>
rect 55 64 56 65 
<< m2 >>
rect 55 64 56 65 
<< m1 >>
rect 56 64 57 65 
<< m2 >>
rect 56 64 57 65 
<< m2 >>
rect 57 64 58 65 
<< m1 >>
rect 58 64 59 65 
<< m2 >>
rect 58 64 59 65 
<< m2 >>
rect 59 64 60 65 
<< m2 >>
rect 63 64 64 65 
<< m1 >>
rect 64 64 65 65 
<< m1 >>
rect 70 64 71 65 
<< m1 >>
rect 100 64 101 65 
<< m1 >>
rect 103 64 104 65 
<< m1 >>
rect 105 64 106 65 
<< m2 >>
rect 105 64 106 65 
<< m2c >>
rect 105 64 106 65 
<< m1 >>
rect 105 64 106 65 
<< m2 >>
rect 105 64 106 65 
<< m1 >>
rect 106 64 107 65 
<< m1 >>
rect 109 64 110 65 
<< m1 >>
rect 114 64 115 65 
<< m1 >>
rect 118 64 119 65 
<< m1 >>
rect 10 65 11 66 
<< m1 >>
rect 13 65 14 66 
<< m1 >>
rect 19 65 20 66 
<< m1 >>
rect 21 65 22 66 
<< m2 >>
rect 27 65 28 66 
<< m1 >>
rect 28 65 29 66 
<< m1 >>
rect 34 65 35 66 
<< m1 >>
rect 38 65 39 66 
<< m2 >>
rect 38 65 39 66 
<< m1 >>
rect 39 65 40 66 
<< m1 >>
rect 40 65 41 66 
<< m2 >>
rect 40 65 41 66 
<< m2c >>
rect 40 65 41 66 
<< m1 >>
rect 40 65 41 66 
<< m2 >>
rect 40 65 41 66 
<< m1 >>
rect 44 65 45 66 
<< m1 >>
rect 46 65 47 66 
<< m1 >>
rect 49 65 50 66 
<< m1 >>
rect 56 65 57 66 
<< m1 >>
rect 58 65 59 66 
<< m2 >>
rect 59 65 60 66 
<< m2 >>
rect 63 65 64 66 
<< m1 >>
rect 64 65 65 66 
<< m1 >>
rect 70 65 71 66 
<< m1 >>
rect 100 65 101 66 
<< m1 >>
rect 103 65 104 66 
<< m1 >>
rect 106 65 107 66 
<< m1 >>
rect 109 65 110 66 
<< m1 >>
rect 114 65 115 66 
<< m1 >>
rect 118 65 119 66 
<< m1 >>
rect 10 66 11 67 
<< pdiffusion >>
rect 12 66 13 67 
<< m1 >>
rect 13 66 14 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< m1 >>
rect 19 66 20 67 
<< m1 >>
rect 21 66 22 67 
<< m2 >>
rect 27 66 28 67 
<< m1 >>
rect 28 66 29 67 
<< pdiffusion >>
rect 30 66 31 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< m1 >>
rect 34 66 35 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< m1 >>
rect 38 66 39 67 
<< m2 >>
rect 38 66 39 67 
<< m1 >>
rect 44 66 45 67 
<< m1 >>
rect 46 66 47 67 
<< pdiffusion >>
rect 48 66 49 67 
<< m1 >>
rect 49 66 50 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 56 66 57 67 
<< m1 >>
rect 58 66 59 67 
<< m2 >>
rect 59 66 60 67 
<< m2 >>
rect 63 66 64 67 
<< m1 >>
rect 64 66 65 67 
<< pdiffusion >>
rect 66 66 67 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< m1 >>
rect 70 66 71 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< pdiffusion >>
rect 84 66 85 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< m1 >>
rect 100 66 101 67 
<< pdiffusion >>
rect 102 66 103 67 
<< m1 >>
rect 103 66 104 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< m1 >>
rect 106 66 107 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< m1 >>
rect 109 66 110 67 
<< m1 >>
rect 114 66 115 67 
<< m1 >>
rect 118 66 119 67 
<< pdiffusion >>
rect 120 66 121 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< m1 >>
rect 10 67 11 68 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< m1 >>
rect 19 67 20 68 
<< m1 >>
rect 21 67 22 68 
<< m2 >>
rect 27 67 28 68 
<< m1 >>
rect 28 67 29 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< m1 >>
rect 38 67 39 68 
<< m2 >>
rect 38 67 39 68 
<< m1 >>
rect 44 67 45 68 
<< m1 >>
rect 46 67 47 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 56 67 57 68 
<< m1 >>
rect 58 67 59 68 
<< m2 >>
rect 59 67 60 68 
<< m2 >>
rect 63 67 64 68 
<< m1 >>
rect 64 67 65 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< m1 >>
rect 100 67 101 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< m1 >>
rect 109 67 110 68 
<< m1 >>
rect 114 67 115 68 
<< m1 >>
rect 118 67 119 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< m1 >>
rect 10 68 11 69 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< m1 >>
rect 19 68 20 69 
<< m1 >>
rect 21 68 22 69 
<< m2 >>
rect 27 68 28 69 
<< m1 >>
rect 28 68 29 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< m1 >>
rect 38 68 39 69 
<< m2 >>
rect 38 68 39 69 
<< m1 >>
rect 44 68 45 69 
<< m1 >>
rect 46 68 47 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 56 68 57 69 
<< m1 >>
rect 58 68 59 69 
<< m2 >>
rect 59 68 60 69 
<< m2 >>
rect 63 68 64 69 
<< m1 >>
rect 64 68 65 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< m1 >>
rect 100 68 101 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< m1 >>
rect 109 68 110 69 
<< m1 >>
rect 114 68 115 69 
<< m1 >>
rect 118 68 119 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< m1 >>
rect 10 69 11 70 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< m1 >>
rect 19 69 20 70 
<< m1 >>
rect 21 69 22 70 
<< m2 >>
rect 27 69 28 70 
<< m1 >>
rect 28 69 29 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< m1 >>
rect 38 69 39 70 
<< m2 >>
rect 38 69 39 70 
<< m1 >>
rect 44 69 45 70 
<< m1 >>
rect 46 69 47 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 56 69 57 70 
<< m1 >>
rect 58 69 59 70 
<< m2 >>
rect 59 69 60 70 
<< m2 >>
rect 63 69 64 70 
<< m1 >>
rect 64 69 65 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< m1 >>
rect 100 69 101 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< m1 >>
rect 109 69 110 70 
<< m1 >>
rect 114 69 115 70 
<< m1 >>
rect 118 69 119 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< m1 >>
rect 10 70 11 71 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< m1 >>
rect 19 70 20 71 
<< m1 >>
rect 21 70 22 71 
<< m2 >>
rect 27 70 28 71 
<< m1 >>
rect 28 70 29 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< m1 >>
rect 38 70 39 71 
<< m2 >>
rect 38 70 39 71 
<< m1 >>
rect 44 70 45 71 
<< m1 >>
rect 46 70 47 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 56 70 57 71 
<< m1 >>
rect 58 70 59 71 
<< m2 >>
rect 59 70 60 71 
<< m2 >>
rect 63 70 64 71 
<< m1 >>
rect 64 70 65 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< m1 >>
rect 100 70 101 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< m1 >>
rect 109 70 110 71 
<< m1 >>
rect 114 70 115 71 
<< m1 >>
rect 118 70 119 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< m1 >>
rect 10 71 11 72 
<< pdiffusion >>
rect 12 71 13 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< m1 >>
rect 16 71 17 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< m1 >>
rect 19 71 20 72 
<< m1 >>
rect 21 71 22 72 
<< m2 >>
rect 27 71 28 72 
<< m1 >>
rect 28 71 29 72 
<< pdiffusion >>
rect 30 71 31 72 
<< m1 >>
rect 31 71 32 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< m1 >>
rect 34 71 35 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< m1 >>
rect 38 71 39 72 
<< m2 >>
rect 38 71 39 72 
<< m1 >>
rect 44 71 45 72 
<< m1 >>
rect 46 71 47 72 
<< pdiffusion >>
rect 48 71 49 72 
<< m1 >>
rect 49 71 50 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< m1 >>
rect 52 71 53 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 56 71 57 72 
<< m1 >>
rect 58 71 59 72 
<< m2 >>
rect 59 71 60 72 
<< m2 >>
rect 63 71 64 72 
<< m1 >>
rect 64 71 65 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< m1 >>
rect 88 71 89 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< m1 >>
rect 100 71 101 72 
<< pdiffusion >>
rect 102 71 103 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< m1 >>
rect 109 71 110 72 
<< m1 >>
rect 114 71 115 72 
<< m2 >>
rect 114 71 115 72 
<< m2c >>
rect 114 71 115 72 
<< m1 >>
rect 114 71 115 72 
<< m2 >>
rect 114 71 115 72 
<< m1 >>
rect 118 71 119 72 
<< pdiffusion >>
rect 120 71 121 72 
<< m1 >>
rect 121 71 122 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< m1 >>
rect 10 72 11 73 
<< m1 >>
rect 16 72 17 73 
<< m1 >>
rect 19 72 20 73 
<< m1 >>
rect 21 72 22 73 
<< m2 >>
rect 27 72 28 73 
<< m1 >>
rect 28 72 29 73 
<< m1 >>
rect 31 72 32 73 
<< m1 >>
rect 34 72 35 73 
<< m1 >>
rect 38 72 39 73 
<< m2 >>
rect 38 72 39 73 
<< m1 >>
rect 44 72 45 73 
<< m1 >>
rect 46 72 47 73 
<< m1 >>
rect 49 72 50 73 
<< m1 >>
rect 52 72 53 73 
<< m1 >>
rect 56 72 57 73 
<< m1 >>
rect 58 72 59 73 
<< m2 >>
rect 59 72 60 73 
<< m2 >>
rect 63 72 64 73 
<< m1 >>
rect 64 72 65 73 
<< m1 >>
rect 88 72 89 73 
<< m1 >>
rect 100 72 101 73 
<< m1 >>
rect 109 72 110 73 
<< m2 >>
rect 114 72 115 73 
<< m1 >>
rect 118 72 119 73 
<< m1 >>
rect 121 72 122 73 
<< m1 >>
rect 10 73 11 74 
<< m1 >>
rect 16 73 17 74 
<< m1 >>
rect 17 73 18 74 
<< m1 >>
rect 18 73 19 74 
<< m1 >>
rect 19 73 20 74 
<< m1 >>
rect 21 73 22 74 
<< m2 >>
rect 27 73 28 74 
<< m1 >>
rect 28 73 29 74 
<< m1 >>
rect 29 73 30 74 
<< m1 >>
rect 30 73 31 74 
<< m1 >>
rect 31 73 32 74 
<< m1 >>
rect 34 73 35 74 
<< m1 >>
rect 38 73 39 74 
<< m2 >>
rect 38 73 39 74 
<< m2 >>
rect 39 73 40 74 
<< m1 >>
rect 40 73 41 74 
<< m2 >>
rect 40 73 41 74 
<< m2c >>
rect 40 73 41 74 
<< m1 >>
rect 40 73 41 74 
<< m2 >>
rect 40 73 41 74 
<< m1 >>
rect 41 73 42 74 
<< m1 >>
rect 42 73 43 74 
<< m2 >>
rect 42 73 43 74 
<< m2c >>
rect 42 73 43 74 
<< m1 >>
rect 42 73 43 74 
<< m2 >>
rect 42 73 43 74 
<< m2 >>
rect 43 73 44 74 
<< m1 >>
rect 44 73 45 74 
<< m2 >>
rect 44 73 45 74 
<< m2 >>
rect 45 73 46 74 
<< m1 >>
rect 46 73 47 74 
<< m2 >>
rect 46 73 47 74 
<< m2 >>
rect 47 73 48 74 
<< m1 >>
rect 48 73 49 74 
<< m2 >>
rect 48 73 49 74 
<< m2c >>
rect 48 73 49 74 
<< m1 >>
rect 48 73 49 74 
<< m2 >>
rect 48 73 49 74 
<< m1 >>
rect 49 73 50 74 
<< m1 >>
rect 52 73 53 74 
<< m1 >>
rect 56 73 57 74 
<< m1 >>
rect 58 73 59 74 
<< m2 >>
rect 59 73 60 74 
<< m1 >>
rect 60 73 61 74 
<< m2 >>
rect 60 73 61 74 
<< m2c >>
rect 60 73 61 74 
<< m1 >>
rect 60 73 61 74 
<< m2 >>
rect 60 73 61 74 
<< m1 >>
rect 61 73 62 74 
<< m1 >>
rect 62 73 63 74 
<< m2 >>
rect 63 73 64 74 
<< m1 >>
rect 64 73 65 74 
<< m2 >>
rect 64 73 65 74 
<< m2 >>
rect 65 73 66 74 
<< m1 >>
rect 66 73 67 74 
<< m2 >>
rect 66 73 67 74 
<< m2c >>
rect 66 73 67 74 
<< m1 >>
rect 66 73 67 74 
<< m2 >>
rect 66 73 67 74 
<< m1 >>
rect 88 73 89 74 
<< m1 >>
rect 89 73 90 74 
<< m1 >>
rect 90 73 91 74 
<< m1 >>
rect 91 73 92 74 
<< m1 >>
rect 92 73 93 74 
<< m1 >>
rect 93 73 94 74 
<< m1 >>
rect 94 73 95 74 
<< m1 >>
rect 95 73 96 74 
<< m1 >>
rect 96 73 97 74 
<< m1 >>
rect 97 73 98 74 
<< m1 >>
rect 98 73 99 74 
<< m1 >>
rect 99 73 100 74 
<< m1 >>
rect 100 73 101 74 
<< m1 >>
rect 107 73 108 74 
<< m2 >>
rect 107 73 108 74 
<< m2c >>
rect 107 73 108 74 
<< m1 >>
rect 107 73 108 74 
<< m2 >>
rect 107 73 108 74 
<< m2 >>
rect 108 73 109 74 
<< m1 >>
rect 109 73 110 74 
<< m2 >>
rect 109 73 110 74 
<< m2 >>
rect 110 73 111 74 
<< m1 >>
rect 111 73 112 74 
<< m2 >>
rect 111 73 112 74 
<< m2c >>
rect 111 73 112 74 
<< m1 >>
rect 111 73 112 74 
<< m2 >>
rect 111 73 112 74 
<< m1 >>
rect 112 73 113 74 
<< m1 >>
rect 113 73 114 74 
<< m1 >>
rect 114 73 115 74 
<< m2 >>
rect 114 73 115 74 
<< m1 >>
rect 115 73 116 74 
<< m1 >>
rect 116 73 117 74 
<< m2 >>
rect 116 73 117 74 
<< m2c >>
rect 116 73 117 74 
<< m1 >>
rect 116 73 117 74 
<< m2 >>
rect 116 73 117 74 
<< m2 >>
rect 117 73 118 74 
<< m1 >>
rect 118 73 119 74 
<< m2 >>
rect 118 73 119 74 
<< m2 >>
rect 119 73 120 74 
<< m1 >>
rect 120 73 121 74 
<< m2 >>
rect 120 73 121 74 
<< m2c >>
rect 120 73 121 74 
<< m1 >>
rect 120 73 121 74 
<< m2 >>
rect 120 73 121 74 
<< m1 >>
rect 121 73 122 74 
<< m1 >>
rect 10 74 11 75 
<< m1 >>
rect 21 74 22 75 
<< m2 >>
rect 27 74 28 75 
<< m1 >>
rect 34 74 35 75 
<< m1 >>
rect 38 74 39 75 
<< m1 >>
rect 44 74 45 75 
<< m1 >>
rect 46 74 47 75 
<< m1 >>
rect 52 74 53 75 
<< m1 >>
rect 56 74 57 75 
<< m1 >>
rect 58 74 59 75 
<< m1 >>
rect 62 74 63 75 
<< m1 >>
rect 64 74 65 75 
<< m1 >>
rect 66 74 67 75 
<< m1 >>
rect 107 74 108 75 
<< m1 >>
rect 109 74 110 75 
<< m2 >>
rect 114 74 115 75 
<< m1 >>
rect 118 74 119 75 
<< m1 >>
rect 10 75 11 76 
<< m1 >>
rect 21 75 22 76 
<< m2 >>
rect 27 75 28 76 
<< m1 >>
rect 34 75 35 76 
<< m1 >>
rect 38 75 39 76 
<< m1 >>
rect 44 75 45 76 
<< m1 >>
rect 46 75 47 76 
<< m1 >>
rect 52 75 53 76 
<< m1 >>
rect 56 75 57 76 
<< m2 >>
rect 56 75 57 76 
<< m2c >>
rect 56 75 57 76 
<< m1 >>
rect 56 75 57 76 
<< m2 >>
rect 56 75 57 76 
<< m2 >>
rect 57 75 58 76 
<< m1 >>
rect 58 75 59 76 
<< m2 >>
rect 58 75 59 76 
<< m2 >>
rect 59 75 60 76 
<< m1 >>
rect 60 75 61 76 
<< m2 >>
rect 60 75 61 76 
<< m2c >>
rect 60 75 61 76 
<< m1 >>
rect 60 75 61 76 
<< m2 >>
rect 60 75 61 76 
<< m1 >>
rect 62 75 63 76 
<< m1 >>
rect 64 75 65 76 
<< m1 >>
rect 66 75 67 76 
<< m1 >>
rect 107 75 108 76 
<< m1 >>
rect 109 75 110 76 
<< m1 >>
rect 114 75 115 76 
<< m2 >>
rect 114 75 115 76 
<< m2c >>
rect 114 75 115 76 
<< m1 >>
rect 114 75 115 76 
<< m2 >>
rect 114 75 115 76 
<< m1 >>
rect 118 75 119 76 
<< m1 >>
rect 10 76 11 77 
<< m1 >>
rect 21 76 22 77 
<< m2 >>
rect 27 76 28 77 
<< m1 >>
rect 28 76 29 77 
<< m1 >>
rect 29 76 30 77 
<< m1 >>
rect 30 76 31 77 
<< m1 >>
rect 31 76 32 77 
<< m1 >>
rect 32 76 33 77 
<< m1 >>
rect 33 76 34 77 
<< m1 >>
rect 34 76 35 77 
<< m1 >>
rect 38 76 39 77 
<< m1 >>
rect 44 76 45 77 
<< m1 >>
rect 46 76 47 77 
<< m1 >>
rect 52 76 53 77 
<< m1 >>
rect 58 76 59 77 
<< m1 >>
rect 60 76 61 77 
<< m1 >>
rect 62 76 63 77 
<< m1 >>
rect 64 76 65 77 
<< m1 >>
rect 66 76 67 77 
<< m1 >>
rect 67 76 68 77 
<< m1 >>
rect 68 76 69 77 
<< m1 >>
rect 69 76 70 77 
<< m1 >>
rect 70 76 71 77 
<< m1 >>
rect 71 76 72 77 
<< m1 >>
rect 72 76 73 77 
<< m1 >>
rect 73 76 74 77 
<< m1 >>
rect 100 76 101 77 
<< m1 >>
rect 101 76 102 77 
<< m1 >>
rect 102 76 103 77 
<< m1 >>
rect 103 76 104 77 
<< m1 >>
rect 104 76 105 77 
<< m1 >>
rect 105 76 106 77 
<< m1 >>
rect 106 76 107 77 
<< m1 >>
rect 107 76 108 77 
<< m1 >>
rect 109 76 110 77 
<< m1 >>
rect 114 76 115 77 
<< m1 >>
rect 118 76 119 77 
<< m1 >>
rect 10 77 11 78 
<< m1 >>
rect 21 77 22 78 
<< m2 >>
rect 27 77 28 78 
<< m1 >>
rect 28 77 29 78 
<< m1 >>
rect 38 77 39 78 
<< m2 >>
rect 38 77 39 78 
<< m2c >>
rect 38 77 39 78 
<< m1 >>
rect 38 77 39 78 
<< m2 >>
rect 38 77 39 78 
<< m1 >>
rect 42 77 43 78 
<< m2 >>
rect 42 77 43 78 
<< m2c >>
rect 42 77 43 78 
<< m1 >>
rect 42 77 43 78 
<< m2 >>
rect 42 77 43 78 
<< m2 >>
rect 43 77 44 78 
<< m1 >>
rect 44 77 45 78 
<< m2 >>
rect 44 77 45 78 
<< m2 >>
rect 45 77 46 78 
<< m1 >>
rect 46 77 47 78 
<< m2 >>
rect 46 77 47 78 
<< m2 >>
rect 47 77 48 78 
<< m1 >>
rect 48 77 49 78 
<< m2 >>
rect 48 77 49 78 
<< m2c >>
rect 48 77 49 78 
<< m1 >>
rect 48 77 49 78 
<< m2 >>
rect 48 77 49 78 
<< m1 >>
rect 49 77 50 78 
<< m1 >>
rect 50 77 51 78 
<< m2 >>
rect 50 77 51 78 
<< m2c >>
rect 50 77 51 78 
<< m1 >>
rect 50 77 51 78 
<< m2 >>
rect 50 77 51 78 
<< m2 >>
rect 51 77 52 78 
<< m1 >>
rect 52 77 53 78 
<< m2 >>
rect 52 77 53 78 
<< m1 >>
rect 53 77 54 78 
<< m1 >>
rect 54 77 55 78 
<< m1 >>
rect 55 77 56 78 
<< m1 >>
rect 56 77 57 78 
<< m2 >>
rect 56 77 57 78 
<< m2c >>
rect 56 77 57 78 
<< m1 >>
rect 56 77 57 78 
<< m2 >>
rect 56 77 57 78 
<< m1 >>
rect 58 77 59 78 
<< m2 >>
rect 58 77 59 78 
<< m2c >>
rect 58 77 59 78 
<< m1 >>
rect 58 77 59 78 
<< m2 >>
rect 58 77 59 78 
<< m1 >>
rect 60 77 61 78 
<< m2 >>
rect 60 77 61 78 
<< m2c >>
rect 60 77 61 78 
<< m1 >>
rect 60 77 61 78 
<< m2 >>
rect 60 77 61 78 
<< m1 >>
rect 62 77 63 78 
<< m2 >>
rect 62 77 63 78 
<< m2c >>
rect 62 77 63 78 
<< m1 >>
rect 62 77 63 78 
<< m2 >>
rect 62 77 63 78 
<< m2 >>
rect 63 77 64 78 
<< m1 >>
rect 64 77 65 78 
<< m2 >>
rect 64 77 65 78 
<< m2 >>
rect 65 77 66 78 
<< m2 >>
rect 66 77 67 78 
<< m2 >>
rect 67 77 68 78 
<< m2 >>
rect 68 77 69 78 
<< m2 >>
rect 69 77 70 78 
<< m2 >>
rect 70 77 71 78 
<< m2 >>
rect 71 77 72 78 
<< m2 >>
rect 72 77 73 78 
<< m1 >>
rect 73 77 74 78 
<< m2 >>
rect 73 77 74 78 
<< m1 >>
rect 100 77 101 78 
<< m1 >>
rect 109 77 110 78 
<< m1 >>
rect 114 77 115 78 
<< m1 >>
rect 118 77 119 78 
<< m1 >>
rect 10 78 11 79 
<< m1 >>
rect 21 78 22 79 
<< m2 >>
rect 27 78 28 79 
<< m1 >>
rect 28 78 29 79 
<< m2 >>
rect 28 78 29 79 
<< m2 >>
rect 29 78 30 79 
<< m1 >>
rect 30 78 31 79 
<< m2 >>
rect 30 78 31 79 
<< m2c >>
rect 30 78 31 79 
<< m1 >>
rect 30 78 31 79 
<< m2 >>
rect 30 78 31 79 
<< m2 >>
rect 38 78 39 79 
<< m1 >>
rect 42 78 43 79 
<< m1 >>
rect 44 78 45 79 
<< m1 >>
rect 46 78 47 79 
<< m2 >>
rect 52 78 53 79 
<< m2 >>
rect 56 78 57 79 
<< m2 >>
rect 58 78 59 79 
<< m2 >>
rect 60 78 61 79 
<< m1 >>
rect 64 78 65 79 
<< m1 >>
rect 73 78 74 79 
<< m2 >>
rect 73 78 74 79 
<< m1 >>
rect 100 78 101 79 
<< m1 >>
rect 109 78 110 79 
<< m1 >>
rect 114 78 115 79 
<< m1 >>
rect 118 78 119 79 
<< m1 >>
rect 10 79 11 80 
<< m1 >>
rect 21 79 22 80 
<< m1 >>
rect 28 79 29 80 
<< m1 >>
rect 30 79 31 80 
<< m1 >>
rect 31 79 32 80 
<< m1 >>
rect 32 79 33 80 
<< m1 >>
rect 33 79 34 80 
<< m1 >>
rect 34 79 35 80 
<< m1 >>
rect 35 79 36 80 
<< m1 >>
rect 36 79 37 80 
<< m1 >>
rect 37 79 38 80 
<< m1 >>
rect 38 79 39 80 
<< m2 >>
rect 38 79 39 80 
<< m1 >>
rect 39 79 40 80 
<< m1 >>
rect 40 79 41 80 
<< m2 >>
rect 40 79 41 80 
<< m2c >>
rect 40 79 41 80 
<< m1 >>
rect 40 79 41 80 
<< m2 >>
rect 40 79 41 80 
<< m2 >>
rect 41 79 42 80 
<< m1 >>
rect 42 79 43 80 
<< m1 >>
rect 44 79 45 80 
<< m2 >>
rect 44 79 45 80 
<< m2c >>
rect 44 79 45 80 
<< m1 >>
rect 44 79 45 80 
<< m2 >>
rect 44 79 45 80 
<< m2 >>
rect 45 79 46 80 
<< m1 >>
rect 46 79 47 80 
<< m2 >>
rect 46 79 47 80 
<< m2 >>
rect 47 79 48 80 
<< m1 >>
rect 48 79 49 80 
<< m2 >>
rect 48 79 49 80 
<< m2c >>
rect 48 79 49 80 
<< m1 >>
rect 48 79 49 80 
<< m2 >>
rect 48 79 49 80 
<< m1 >>
rect 49 79 50 80 
<< m1 >>
rect 50 79 51 80 
<< m1 >>
rect 51 79 52 80 
<< m1 >>
rect 52 79 53 80 
<< m2 >>
rect 52 79 53 80 
<< m1 >>
rect 53 79 54 80 
<< m1 >>
rect 54 79 55 80 
<< m1 >>
rect 55 79 56 80 
<< m1 >>
rect 56 79 57 80 
<< m2 >>
rect 56 79 57 80 
<< m1 >>
rect 57 79 58 80 
<< m1 >>
rect 58 79 59 80 
<< m2 >>
rect 58 79 59 80 
<< m1 >>
rect 59 79 60 80 
<< m1 >>
rect 60 79 61 80 
<< m2 >>
rect 60 79 61 80 
<< m1 >>
rect 61 79 62 80 
<< m1 >>
rect 62 79 63 80 
<< m2 >>
rect 62 79 63 80 
<< m2c >>
rect 62 79 63 80 
<< m1 >>
rect 62 79 63 80 
<< m2 >>
rect 62 79 63 80 
<< m2 >>
rect 63 79 64 80 
<< m1 >>
rect 64 79 65 80 
<< m2 >>
rect 64 79 65 80 
<< m2 >>
rect 65 79 66 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m2c >>
rect 66 79 67 80 
<< m1 >>
rect 66 79 67 80 
<< m2 >>
rect 66 79 67 80 
<< m1 >>
rect 67 79 68 80 
<< m1 >>
rect 68 79 69 80 
<< m1 >>
rect 69 79 70 80 
<< m1 >>
rect 70 79 71 80 
<< m1 >>
rect 73 79 74 80 
<< m2 >>
rect 73 79 74 80 
<< m1 >>
rect 100 79 101 80 
<< m2 >>
rect 100 79 101 80 
<< m2 >>
rect 101 79 102 80 
<< m1 >>
rect 102 79 103 80 
<< m2 >>
rect 102 79 103 80 
<< m2c >>
rect 102 79 103 80 
<< m1 >>
rect 102 79 103 80 
<< m2 >>
rect 102 79 103 80 
<< m1 >>
rect 103 79 104 80 
<< m1 >>
rect 104 79 105 80 
<< m1 >>
rect 105 79 106 80 
<< m1 >>
rect 106 79 107 80 
<< m1 >>
rect 109 79 110 80 
<< m1 >>
rect 114 79 115 80 
<< m1 >>
rect 118 79 119 80 
<< m1 >>
rect 10 80 11 81 
<< m1 >>
rect 21 80 22 81 
<< m2 >>
rect 21 80 22 81 
<< m2c >>
rect 21 80 22 81 
<< m1 >>
rect 21 80 22 81 
<< m2 >>
rect 21 80 22 81 
<< m1 >>
rect 28 80 29 81 
<< m2 >>
rect 38 80 39 81 
<< m2 >>
rect 41 80 42 81 
<< m1 >>
rect 42 80 43 81 
<< m1 >>
rect 46 80 47 81 
<< m2 >>
rect 52 80 53 81 
<< m2 >>
rect 56 80 57 81 
<< m2 >>
rect 58 80 59 81 
<< m2 >>
rect 60 80 61 81 
<< m1 >>
rect 64 80 65 81 
<< m1 >>
rect 70 80 71 81 
<< m1 >>
rect 73 80 74 81 
<< m2 >>
rect 73 80 74 81 
<< m1 >>
rect 100 80 101 81 
<< m2 >>
rect 100 80 101 81 
<< m1 >>
rect 106 80 107 81 
<< m1 >>
rect 109 80 110 81 
<< m1 >>
rect 114 80 115 81 
<< m1 >>
rect 118 80 119 81 
<< m1 >>
rect 10 81 11 82 
<< m2 >>
rect 21 81 22 82 
<< m1 >>
rect 28 81 29 82 
<< m1 >>
rect 34 81 35 82 
<< m1 >>
rect 35 81 36 82 
<< m1 >>
rect 36 81 37 82 
<< m1 >>
rect 37 81 38 82 
<< m1 >>
rect 38 81 39 82 
<< m2 >>
rect 38 81 39 82 
<< m2c >>
rect 38 81 39 82 
<< m1 >>
rect 38 81 39 82 
<< m2 >>
rect 38 81 39 82 
<< m2 >>
rect 41 81 42 82 
<< m1 >>
rect 42 81 43 82 
<< m2 >>
rect 42 81 43 82 
<< m2 >>
rect 43 81 44 82 
<< m1 >>
rect 44 81 45 82 
<< m2 >>
rect 44 81 45 82 
<< m2c >>
rect 44 81 45 82 
<< m1 >>
rect 44 81 45 82 
<< m2 >>
rect 44 81 45 82 
<< m1 >>
rect 46 81 47 82 
<< m1 >>
rect 52 81 53 82 
<< m2 >>
rect 52 81 53 82 
<< m2c >>
rect 52 81 53 82 
<< m1 >>
rect 52 81 53 82 
<< m2 >>
rect 52 81 53 82 
<< m1 >>
rect 56 81 57 82 
<< m2 >>
rect 56 81 57 82 
<< m2c >>
rect 56 81 57 82 
<< m1 >>
rect 56 81 57 82 
<< m2 >>
rect 56 81 57 82 
<< m1 >>
rect 58 81 59 82 
<< m2 >>
rect 58 81 59 82 
<< m2c >>
rect 58 81 59 82 
<< m1 >>
rect 58 81 59 82 
<< m2 >>
rect 58 81 59 82 
<< m1 >>
rect 60 81 61 82 
<< m2 >>
rect 60 81 61 82 
<< m2c >>
rect 60 81 61 82 
<< m1 >>
rect 60 81 61 82 
<< m2 >>
rect 60 81 61 82 
<< m1 >>
rect 64 81 65 82 
<< m1 >>
rect 70 81 71 82 
<< m1 >>
rect 73 81 74 82 
<< m2 >>
rect 73 81 74 82 
<< m1 >>
rect 100 81 101 82 
<< m2 >>
rect 100 81 101 82 
<< m1 >>
rect 106 81 107 82 
<< m1 >>
rect 109 81 110 82 
<< m1 >>
rect 114 81 115 82 
<< m1 >>
rect 118 81 119 82 
<< m1 >>
rect 10 82 11 83 
<< m1 >>
rect 16 82 17 83 
<< m1 >>
rect 17 82 18 83 
<< m1 >>
rect 18 82 19 83 
<< m1 >>
rect 19 82 20 83 
<< m1 >>
rect 20 82 21 83 
<< m1 >>
rect 21 82 22 83 
<< m2 >>
rect 21 82 22 83 
<< m1 >>
rect 22 82 23 83 
<< m1 >>
rect 23 82 24 83 
<< m1 >>
rect 24 82 25 83 
<< m1 >>
rect 25 82 26 83 
<< m1 >>
rect 26 82 27 83 
<< m2 >>
rect 26 82 27 83 
<< m2c >>
rect 26 82 27 83 
<< m1 >>
rect 26 82 27 83 
<< m2 >>
rect 26 82 27 83 
<< m2 >>
rect 27 82 28 83 
<< m1 >>
rect 28 82 29 83 
<< m1 >>
rect 34 82 35 83 
<< m1 >>
rect 42 82 43 83 
<< m1 >>
rect 44 82 45 83 
<< m1 >>
rect 46 82 47 83 
<< m1 >>
rect 52 82 53 83 
<< m1 >>
rect 56 82 57 83 
<< m1 >>
rect 58 82 59 83 
<< m1 >>
rect 60 82 61 83 
<< m1 >>
rect 64 82 65 83 
<< m1 >>
rect 70 82 71 83 
<< m1 >>
rect 73 82 74 83 
<< m2 >>
rect 73 82 74 83 
<< m1 >>
rect 100 82 101 83 
<< m2 >>
rect 100 82 101 83 
<< m1 >>
rect 106 82 107 83 
<< m1 >>
rect 109 82 110 83 
<< m1 >>
rect 114 82 115 83 
<< m1 >>
rect 118 82 119 83 
<< m1 >>
rect 119 82 120 83 
<< m1 >>
rect 120 82 121 83 
<< m1 >>
rect 121 82 122 83 
<< m1 >>
rect 10 83 11 84 
<< m1 >>
rect 16 83 17 84 
<< m2 >>
rect 21 83 22 84 
<< m2 >>
rect 27 83 28 84 
<< m1 >>
rect 28 83 29 84 
<< m1 >>
rect 34 83 35 84 
<< m1 >>
rect 42 83 43 84 
<< m1 >>
rect 44 83 45 84 
<< m1 >>
rect 46 83 47 84 
<< m1 >>
rect 52 83 53 84 
<< m1 >>
rect 56 83 57 84 
<< m1 >>
rect 58 83 59 84 
<< m1 >>
rect 60 83 61 84 
<< m1 >>
rect 64 83 65 84 
<< m1 >>
rect 70 83 71 84 
<< m1 >>
rect 73 83 74 84 
<< m2 >>
rect 73 83 74 84 
<< m1 >>
rect 100 83 101 84 
<< m2 >>
rect 100 83 101 84 
<< m1 >>
rect 106 83 107 84 
<< m1 >>
rect 109 83 110 84 
<< m1 >>
rect 114 83 115 84 
<< m1 >>
rect 121 83 122 84 
<< m1 >>
rect 10 84 11 85 
<< pdiffusion >>
rect 12 84 13 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< m1 >>
rect 16 84 17 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< m1 >>
rect 21 84 22 85 
<< m2 >>
rect 21 84 22 85 
<< m2c >>
rect 21 84 22 85 
<< m1 >>
rect 21 84 22 85 
<< m2 >>
rect 21 84 22 85 
<< m2 >>
rect 27 84 28 85 
<< m1 >>
rect 28 84 29 85 
<< pdiffusion >>
rect 30 84 31 85 
<< pdiffusion >>
rect 31 84 32 85 
<< pdiffusion >>
rect 32 84 33 85 
<< pdiffusion >>
rect 33 84 34 85 
<< m1 >>
rect 34 84 35 85 
<< pdiffusion >>
rect 34 84 35 85 
<< pdiffusion >>
rect 35 84 36 85 
<< m1 >>
rect 42 84 43 85 
<< m1 >>
rect 44 84 45 85 
<< m1 >>
rect 46 84 47 85 
<< pdiffusion >>
rect 48 84 49 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< m1 >>
rect 52 84 53 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< m1 >>
rect 56 84 57 85 
<< m1 >>
rect 58 84 59 85 
<< m1 >>
rect 60 84 61 85 
<< m1 >>
rect 64 84 65 85 
<< pdiffusion >>
rect 66 84 67 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< m1 >>
rect 70 84 71 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< m1 >>
rect 73 84 74 85 
<< m2 >>
rect 73 84 74 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 100 84 101 85 
<< m2 >>
rect 100 84 101 85 
<< pdiffusion >>
rect 102 84 103 85 
<< pdiffusion >>
rect 103 84 104 85 
<< pdiffusion >>
rect 104 84 105 85 
<< pdiffusion >>
rect 105 84 106 85 
<< m1 >>
rect 106 84 107 85 
<< pdiffusion >>
rect 106 84 107 85 
<< pdiffusion >>
rect 107 84 108 85 
<< m1 >>
rect 109 84 110 85 
<< m1 >>
rect 114 84 115 85 
<< pdiffusion >>
rect 120 84 121 85 
<< m1 >>
rect 121 84 122 85 
<< pdiffusion >>
rect 121 84 122 85 
<< pdiffusion >>
rect 122 84 123 85 
<< pdiffusion >>
rect 123 84 124 85 
<< pdiffusion >>
rect 124 84 125 85 
<< pdiffusion >>
rect 125 84 126 85 
<< m1 >>
rect 10 85 11 86 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< m1 >>
rect 21 85 22 86 
<< m2 >>
rect 27 85 28 86 
<< m1 >>
rect 28 85 29 86 
<< pdiffusion >>
rect 30 85 31 86 
<< pdiffusion >>
rect 31 85 32 86 
<< pdiffusion >>
rect 32 85 33 86 
<< pdiffusion >>
rect 33 85 34 86 
<< pdiffusion >>
rect 34 85 35 86 
<< pdiffusion >>
rect 35 85 36 86 
<< m1 >>
rect 42 85 43 86 
<< m1 >>
rect 44 85 45 86 
<< m1 >>
rect 46 85 47 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< m1 >>
rect 56 85 57 86 
<< m1 >>
rect 58 85 59 86 
<< m1 >>
rect 60 85 61 86 
<< m1 >>
rect 64 85 65 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< m1 >>
rect 73 85 74 86 
<< m2 >>
rect 73 85 74 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 100 85 101 86 
<< m2 >>
rect 100 85 101 86 
<< pdiffusion >>
rect 102 85 103 86 
<< pdiffusion >>
rect 103 85 104 86 
<< pdiffusion >>
rect 104 85 105 86 
<< pdiffusion >>
rect 105 85 106 86 
<< pdiffusion >>
rect 106 85 107 86 
<< pdiffusion >>
rect 107 85 108 86 
<< m1 >>
rect 109 85 110 86 
<< m1 >>
rect 114 85 115 86 
<< pdiffusion >>
rect 120 85 121 86 
<< pdiffusion >>
rect 121 85 122 86 
<< pdiffusion >>
rect 122 85 123 86 
<< pdiffusion >>
rect 123 85 124 86 
<< pdiffusion >>
rect 124 85 125 86 
<< pdiffusion >>
rect 125 85 126 86 
<< m1 >>
rect 10 86 11 87 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< m1 >>
rect 21 86 22 87 
<< m2 >>
rect 27 86 28 87 
<< m1 >>
rect 28 86 29 87 
<< pdiffusion >>
rect 30 86 31 87 
<< pdiffusion >>
rect 31 86 32 87 
<< pdiffusion >>
rect 32 86 33 87 
<< pdiffusion >>
rect 33 86 34 87 
<< pdiffusion >>
rect 34 86 35 87 
<< pdiffusion >>
rect 35 86 36 87 
<< m1 >>
rect 42 86 43 87 
<< m1 >>
rect 44 86 45 87 
<< m1 >>
rect 46 86 47 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< m1 >>
rect 56 86 57 87 
<< m1 >>
rect 58 86 59 87 
<< m1 >>
rect 60 86 61 87 
<< m1 >>
rect 64 86 65 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< m1 >>
rect 73 86 74 87 
<< m2 >>
rect 73 86 74 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 100 86 101 87 
<< m2 >>
rect 100 86 101 87 
<< pdiffusion >>
rect 102 86 103 87 
<< pdiffusion >>
rect 103 86 104 87 
<< pdiffusion >>
rect 104 86 105 87 
<< pdiffusion >>
rect 105 86 106 87 
<< pdiffusion >>
rect 106 86 107 87 
<< pdiffusion >>
rect 107 86 108 87 
<< m1 >>
rect 109 86 110 87 
<< m1 >>
rect 114 86 115 87 
<< pdiffusion >>
rect 120 86 121 87 
<< pdiffusion >>
rect 121 86 122 87 
<< pdiffusion >>
rect 122 86 123 87 
<< pdiffusion >>
rect 123 86 124 87 
<< pdiffusion >>
rect 124 86 125 87 
<< pdiffusion >>
rect 125 86 126 87 
<< m1 >>
rect 10 87 11 88 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< m1 >>
rect 21 87 22 88 
<< m2 >>
rect 27 87 28 88 
<< m1 >>
rect 28 87 29 88 
<< pdiffusion >>
rect 30 87 31 88 
<< pdiffusion >>
rect 31 87 32 88 
<< pdiffusion >>
rect 32 87 33 88 
<< pdiffusion >>
rect 33 87 34 88 
<< pdiffusion >>
rect 34 87 35 88 
<< pdiffusion >>
rect 35 87 36 88 
<< m1 >>
rect 42 87 43 88 
<< m1 >>
rect 44 87 45 88 
<< m1 >>
rect 46 87 47 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< m1 >>
rect 56 87 57 88 
<< m1 >>
rect 58 87 59 88 
<< m1 >>
rect 60 87 61 88 
<< m1 >>
rect 64 87 65 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< m1 >>
rect 73 87 74 88 
<< m2 >>
rect 73 87 74 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 100 87 101 88 
<< m2 >>
rect 100 87 101 88 
<< pdiffusion >>
rect 102 87 103 88 
<< pdiffusion >>
rect 103 87 104 88 
<< pdiffusion >>
rect 104 87 105 88 
<< pdiffusion >>
rect 105 87 106 88 
<< pdiffusion >>
rect 106 87 107 88 
<< pdiffusion >>
rect 107 87 108 88 
<< m1 >>
rect 109 87 110 88 
<< m1 >>
rect 114 87 115 88 
<< pdiffusion >>
rect 120 87 121 88 
<< pdiffusion >>
rect 121 87 122 88 
<< pdiffusion >>
rect 122 87 123 88 
<< pdiffusion >>
rect 123 87 124 88 
<< pdiffusion >>
rect 124 87 125 88 
<< pdiffusion >>
rect 125 87 126 88 
<< m1 >>
rect 10 88 11 89 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< m1 >>
rect 21 88 22 89 
<< m2 >>
rect 27 88 28 89 
<< m1 >>
rect 28 88 29 89 
<< pdiffusion >>
rect 30 88 31 89 
<< pdiffusion >>
rect 31 88 32 89 
<< pdiffusion >>
rect 32 88 33 89 
<< pdiffusion >>
rect 33 88 34 89 
<< pdiffusion >>
rect 34 88 35 89 
<< pdiffusion >>
rect 35 88 36 89 
<< m1 >>
rect 42 88 43 89 
<< m1 >>
rect 44 88 45 89 
<< m1 >>
rect 46 88 47 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< m1 >>
rect 56 88 57 89 
<< m1 >>
rect 58 88 59 89 
<< m1 >>
rect 60 88 61 89 
<< m1 >>
rect 64 88 65 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< m1 >>
rect 73 88 74 89 
<< m2 >>
rect 73 88 74 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 100 88 101 89 
<< m2 >>
rect 100 88 101 89 
<< pdiffusion >>
rect 102 88 103 89 
<< pdiffusion >>
rect 103 88 104 89 
<< pdiffusion >>
rect 104 88 105 89 
<< pdiffusion >>
rect 105 88 106 89 
<< pdiffusion >>
rect 106 88 107 89 
<< pdiffusion >>
rect 107 88 108 89 
<< m1 >>
rect 109 88 110 89 
<< m1 >>
rect 114 88 115 89 
<< pdiffusion >>
rect 120 88 121 89 
<< pdiffusion >>
rect 121 88 122 89 
<< pdiffusion >>
rect 122 88 123 89 
<< pdiffusion >>
rect 123 88 124 89 
<< pdiffusion >>
rect 124 88 125 89 
<< pdiffusion >>
rect 125 88 126 89 
<< m1 >>
rect 10 89 11 90 
<< pdiffusion >>
rect 12 89 13 90 
<< m1 >>
rect 13 89 14 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< m1 >>
rect 21 89 22 90 
<< m2 >>
rect 27 89 28 90 
<< m1 >>
rect 28 89 29 90 
<< pdiffusion >>
rect 30 89 31 90 
<< m1 >>
rect 31 89 32 90 
<< pdiffusion >>
rect 31 89 32 90 
<< pdiffusion >>
rect 32 89 33 90 
<< pdiffusion >>
rect 33 89 34 90 
<< pdiffusion >>
rect 34 89 35 90 
<< pdiffusion >>
rect 35 89 36 90 
<< m1 >>
rect 42 89 43 90 
<< m1 >>
rect 44 89 45 90 
<< m1 >>
rect 46 89 47 90 
<< pdiffusion >>
rect 48 89 49 90 
<< m1 >>
rect 49 89 50 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< m1 >>
rect 56 89 57 90 
<< m1 >>
rect 58 89 59 90 
<< m1 >>
rect 60 89 61 90 
<< m1 >>
rect 64 89 65 90 
<< pdiffusion >>
rect 66 89 67 90 
<< m1 >>
rect 67 89 68 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< m1 >>
rect 73 89 74 90 
<< m2 >>
rect 73 89 74 90 
<< pdiffusion >>
rect 84 89 85 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< m1 >>
rect 88 89 89 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 100 89 101 90 
<< m2 >>
rect 100 89 101 90 
<< pdiffusion >>
rect 102 89 103 90 
<< pdiffusion >>
rect 103 89 104 90 
<< pdiffusion >>
rect 104 89 105 90 
<< pdiffusion >>
rect 105 89 106 90 
<< m1 >>
rect 106 89 107 90 
<< pdiffusion >>
rect 106 89 107 90 
<< pdiffusion >>
rect 107 89 108 90 
<< m1 >>
rect 109 89 110 90 
<< m1 >>
rect 114 89 115 90 
<< pdiffusion >>
rect 120 89 121 90 
<< m1 >>
rect 121 89 122 90 
<< pdiffusion >>
rect 121 89 122 90 
<< pdiffusion >>
rect 122 89 123 90 
<< pdiffusion >>
rect 123 89 124 90 
<< pdiffusion >>
rect 124 89 125 90 
<< pdiffusion >>
rect 125 89 126 90 
<< m1 >>
rect 10 90 11 91 
<< m1 >>
rect 13 90 14 91 
<< m1 >>
rect 21 90 22 91 
<< m2 >>
rect 27 90 28 91 
<< m1 >>
rect 28 90 29 91 
<< m1 >>
rect 31 90 32 91 
<< m1 >>
rect 42 90 43 91 
<< m2 >>
rect 42 90 43 91 
<< m2c >>
rect 42 90 43 91 
<< m1 >>
rect 42 90 43 91 
<< m2 >>
rect 42 90 43 91 
<< m1 >>
rect 44 90 45 91 
<< m2 >>
rect 44 90 45 91 
<< m2c >>
rect 44 90 45 91 
<< m1 >>
rect 44 90 45 91 
<< m2 >>
rect 44 90 45 91 
<< m1 >>
rect 46 90 47 91 
<< m1 >>
rect 49 90 50 91 
<< m1 >>
rect 56 90 57 91 
<< m2 >>
rect 56 90 57 91 
<< m2c >>
rect 56 90 57 91 
<< m1 >>
rect 56 90 57 91 
<< m2 >>
rect 56 90 57 91 
<< m1 >>
rect 58 90 59 91 
<< m2 >>
rect 58 90 59 91 
<< m2c >>
rect 58 90 59 91 
<< m1 >>
rect 58 90 59 91 
<< m2 >>
rect 58 90 59 91 
<< m1 >>
rect 60 90 61 91 
<< m2 >>
rect 60 90 61 91 
<< m2c >>
rect 60 90 61 91 
<< m1 >>
rect 60 90 61 91 
<< m2 >>
rect 60 90 61 91 
<< m1 >>
rect 64 90 65 91 
<< m1 >>
rect 67 90 68 91 
<< m1 >>
rect 73 90 74 91 
<< m2 >>
rect 73 90 74 91 
<< m1 >>
rect 88 90 89 91 
<< m1 >>
rect 100 90 101 91 
<< m2 >>
rect 100 90 101 91 
<< m1 >>
rect 106 90 107 91 
<< m1 >>
rect 109 90 110 91 
<< m1 >>
rect 114 90 115 91 
<< m1 >>
rect 121 90 122 91 
<< m1 >>
rect 10 91 11 92 
<< m1 >>
rect 13 91 14 92 
<< m1 >>
rect 21 91 22 92 
<< m2 >>
rect 27 91 28 92 
<< m1 >>
rect 28 91 29 92 
<< m1 >>
rect 31 91 32 92 
<< m2 >>
rect 42 91 43 92 
<< m2 >>
rect 44 91 45 92 
<< m1 >>
rect 46 91 47 92 
<< m1 >>
rect 49 91 50 92 
<< m2 >>
rect 56 91 57 92 
<< m2 >>
rect 58 91 59 92 
<< m2 >>
rect 60 91 61 92 
<< m1 >>
rect 64 91 65 92 
<< m1 >>
rect 67 91 68 92 
<< m1 >>
rect 73 91 74 92 
<< m2 >>
rect 73 91 74 92 
<< m1 >>
rect 74 91 75 92 
<< m1 >>
rect 75 91 76 92 
<< m1 >>
rect 76 91 77 92 
<< m1 >>
rect 77 91 78 92 
<< m1 >>
rect 78 91 79 92 
<< m1 >>
rect 79 91 80 92 
<< m1 >>
rect 80 91 81 92 
<< m1 >>
rect 81 91 82 92 
<< m1 >>
rect 82 91 83 92 
<< m1 >>
rect 83 91 84 92 
<< m1 >>
rect 88 91 89 92 
<< m2 >>
rect 89 91 90 92 
<< m1 >>
rect 90 91 91 92 
<< m2 >>
rect 90 91 91 92 
<< m2c >>
rect 90 91 91 92 
<< m1 >>
rect 90 91 91 92 
<< m2 >>
rect 90 91 91 92 
<< m1 >>
rect 91 91 92 92 
<< m1 >>
rect 92 91 93 92 
<< m1 >>
rect 93 91 94 92 
<< m1 >>
rect 94 91 95 92 
<< m1 >>
rect 95 91 96 92 
<< m1 >>
rect 96 91 97 92 
<< m1 >>
rect 97 91 98 92 
<< m1 >>
rect 98 91 99 92 
<< m1 >>
rect 99 91 100 92 
<< m1 >>
rect 100 91 101 92 
<< m2 >>
rect 100 91 101 92 
<< m1 >>
rect 106 91 107 92 
<< m1 >>
rect 107 91 108 92 
<< m2 >>
rect 107 91 108 92 
<< m2c >>
rect 107 91 108 92 
<< m1 >>
rect 107 91 108 92 
<< m2 >>
rect 107 91 108 92 
<< m2 >>
rect 108 91 109 92 
<< m1 >>
rect 109 91 110 92 
<< m2 >>
rect 109 91 110 92 
<< m1 >>
rect 114 91 115 92 
<< m1 >>
rect 118 91 119 92 
<< m1 >>
rect 119 91 120 92 
<< m1 >>
rect 120 91 121 92 
<< m1 >>
rect 121 91 122 92 
<< m1 >>
rect 10 92 11 93 
<< m1 >>
rect 13 92 14 93 
<< m1 >>
rect 14 92 15 93 
<< m1 >>
rect 15 92 16 93 
<< m1 >>
rect 16 92 17 93 
<< m1 >>
rect 17 92 18 93 
<< m1 >>
rect 18 92 19 93 
<< m1 >>
rect 19 92 20 93 
<< m1 >>
rect 20 92 21 93 
<< m1 >>
rect 21 92 22 93 
<< m2 >>
rect 27 92 28 93 
<< m1 >>
rect 28 92 29 93 
<< m1 >>
rect 31 92 32 93 
<< m1 >>
rect 32 92 33 93 
<< m1 >>
rect 33 92 34 93 
<< m1 >>
rect 34 92 35 93 
<< m1 >>
rect 35 92 36 93 
<< m1 >>
rect 36 92 37 93 
<< m1 >>
rect 37 92 38 93 
<< m1 >>
rect 38 92 39 93 
<< m1 >>
rect 39 92 40 93 
<< m1 >>
rect 40 92 41 93 
<< m1 >>
rect 41 92 42 93 
<< m1 >>
rect 42 92 43 93 
<< m2 >>
rect 42 92 43 93 
<< m1 >>
rect 43 92 44 93 
<< m1 >>
rect 44 92 45 93 
<< m2 >>
rect 44 92 45 93 
<< m1 >>
rect 45 92 46 93 
<< m1 >>
rect 46 92 47 93 
<< m1 >>
rect 49 92 50 93 
<< m1 >>
rect 50 92 51 93 
<< m1 >>
rect 51 92 52 93 
<< m1 >>
rect 52 92 53 93 
<< m1 >>
rect 53 92 54 93 
<< m1 >>
rect 54 92 55 93 
<< m1 >>
rect 55 92 56 93 
<< m1 >>
rect 56 92 57 93 
<< m2 >>
rect 56 92 57 93 
<< m1 >>
rect 57 92 58 93 
<< m1 >>
rect 58 92 59 93 
<< m2 >>
rect 58 92 59 93 
<< m1 >>
rect 59 92 60 93 
<< m1 >>
rect 60 92 61 93 
<< m2 >>
rect 60 92 61 93 
<< m1 >>
rect 61 92 62 93 
<< m1 >>
rect 62 92 63 93 
<< m1 >>
rect 63 92 64 93 
<< m1 >>
rect 64 92 65 93 
<< m1 >>
rect 67 92 68 93 
<< m2 >>
rect 72 92 73 93 
<< m2 >>
rect 73 92 74 93 
<< m1 >>
rect 83 92 84 93 
<< m2 >>
rect 83 92 84 93 
<< m2c >>
rect 83 92 84 93 
<< m1 >>
rect 83 92 84 93 
<< m2 >>
rect 83 92 84 93 
<< m1 >>
rect 86 92 87 93 
<< m2 >>
rect 86 92 87 93 
<< m2c >>
rect 86 92 87 93 
<< m1 >>
rect 86 92 87 93 
<< m2 >>
rect 86 92 87 93 
<< m2 >>
rect 87 92 88 93 
<< m1 >>
rect 88 92 89 93 
<< m2 >>
rect 88 92 89 93 
<< m2 >>
rect 89 92 90 93 
<< m2 >>
rect 100 92 101 93 
<< m1 >>
rect 109 92 110 93 
<< m2 >>
rect 109 92 110 93 
<< m1 >>
rect 114 92 115 93 
<< m1 >>
rect 118 92 119 93 
<< m1 >>
rect 10 93 11 94 
<< m2 >>
rect 27 93 28 94 
<< m1 >>
rect 28 93 29 94 
<< m2 >>
rect 42 93 43 94 
<< m2 >>
rect 44 93 45 94 
<< m2 >>
rect 56 93 57 94 
<< m2 >>
rect 58 93 59 94 
<< m2 >>
rect 60 93 61 94 
<< m1 >>
rect 67 93 68 94 
<< m1 >>
rect 72 93 73 94 
<< m2 >>
rect 72 93 73 94 
<< m2c >>
rect 72 93 73 94 
<< m1 >>
rect 72 93 73 94 
<< m2 >>
rect 72 93 73 94 
<< m2 >>
rect 83 93 84 94 
<< m1 >>
rect 86 93 87 94 
<< m1 >>
rect 88 93 89 94 
<< m1 >>
rect 100 93 101 94 
<< m2 >>
rect 100 93 101 94 
<< m2c >>
rect 100 93 101 94 
<< m1 >>
rect 100 93 101 94 
<< m2 >>
rect 100 93 101 94 
<< m1 >>
rect 109 93 110 94 
<< m2 >>
rect 109 93 110 94 
<< m1 >>
rect 114 93 115 94 
<< m1 >>
rect 118 93 119 94 
<< m1 >>
rect 10 94 11 95 
<< m2 >>
rect 27 94 28 95 
<< m1 >>
rect 28 94 29 95 
<< m2 >>
rect 28 94 29 95 
<< m2 >>
rect 29 94 30 95 
<< m1 >>
rect 30 94 31 95 
<< m2 >>
rect 30 94 31 95 
<< m2c >>
rect 30 94 31 95 
<< m1 >>
rect 30 94 31 95 
<< m2 >>
rect 30 94 31 95 
<< m1 >>
rect 31 94 32 95 
<< m1 >>
rect 32 94 33 95 
<< m1 >>
rect 33 94 34 95 
<< m1 >>
rect 34 94 35 95 
<< m1 >>
rect 35 94 36 95 
<< m1 >>
rect 36 94 37 95 
<< m1 >>
rect 37 94 38 95 
<< m1 >>
rect 38 94 39 95 
<< m1 >>
rect 39 94 40 95 
<< m1 >>
rect 40 94 41 95 
<< m1 >>
rect 41 94 42 95 
<< m1 >>
rect 42 94 43 95 
<< m2 >>
rect 42 94 43 95 
<< m1 >>
rect 43 94 44 95 
<< m1 >>
rect 44 94 45 95 
<< m2 >>
rect 44 94 45 95 
<< m1 >>
rect 45 94 46 95 
<< m1 >>
rect 46 94 47 95 
<< m1 >>
rect 47 94 48 95 
<< m1 >>
rect 48 94 49 95 
<< m1 >>
rect 49 94 50 95 
<< m1 >>
rect 50 94 51 95 
<< m1 >>
rect 51 94 52 95 
<< m1 >>
rect 52 94 53 95 
<< m1 >>
rect 53 94 54 95 
<< m1 >>
rect 54 94 55 95 
<< m1 >>
rect 55 94 56 95 
<< m1 >>
rect 56 94 57 95 
<< m2 >>
rect 56 94 57 95 
<< m1 >>
rect 57 94 58 95 
<< m1 >>
rect 58 94 59 95 
<< m2 >>
rect 58 94 59 95 
<< m1 >>
rect 59 94 60 95 
<< m1 >>
rect 60 94 61 95 
<< m2 >>
rect 60 94 61 95 
<< m1 >>
rect 61 94 62 95 
<< m1 >>
rect 62 94 63 95 
<< m1 >>
rect 63 94 64 95 
<< m1 >>
rect 64 94 65 95 
<< m1 >>
rect 65 94 66 95 
<< m1 >>
rect 66 94 67 95 
<< m1 >>
rect 67 94 68 95 
<< m1 >>
rect 72 94 73 95 
<< m2 >>
rect 83 94 84 95 
<< m1 >>
rect 84 94 85 95 
<< m2 >>
rect 84 94 85 95 
<< m1 >>
rect 85 94 86 95 
<< m2 >>
rect 85 94 86 95 
<< m1 >>
rect 86 94 87 95 
<< m2 >>
rect 86 94 87 95 
<< m2 >>
rect 87 94 88 95 
<< m1 >>
rect 88 94 89 95 
<< m2 >>
rect 88 94 89 95 
<< m2 >>
rect 89 94 90 95 
<< m1 >>
rect 90 94 91 95 
<< m2 >>
rect 90 94 91 95 
<< m2c >>
rect 90 94 91 95 
<< m1 >>
rect 90 94 91 95 
<< m2 >>
rect 90 94 91 95 
<< m1 >>
rect 100 94 101 95 
<< m1 >>
rect 109 94 110 95 
<< m2 >>
rect 109 94 110 95 
<< m1 >>
rect 114 94 115 95 
<< m1 >>
rect 118 94 119 95 
<< m1 >>
rect 10 95 11 96 
<< m1 >>
rect 28 95 29 96 
<< m2 >>
rect 42 95 43 96 
<< m2 >>
rect 44 95 45 96 
<< m2 >>
rect 56 95 57 96 
<< m2 >>
rect 58 95 59 96 
<< m2 >>
rect 60 95 61 96 
<< m2 >>
rect 62 95 63 96 
<< m2 >>
rect 63 95 64 96 
<< m2 >>
rect 64 95 65 96 
<< m2 >>
rect 65 95 66 96 
<< m2 >>
rect 66 95 67 96 
<< m2 >>
rect 67 95 68 96 
<< m2 >>
rect 68 95 69 96 
<< m2 >>
rect 69 95 70 96 
<< m1 >>
rect 70 95 71 96 
<< m2 >>
rect 70 95 71 96 
<< m2c >>
rect 70 95 71 96 
<< m1 >>
rect 70 95 71 96 
<< m2 >>
rect 70 95 71 96 
<< m1 >>
rect 71 95 72 96 
<< m1 >>
rect 72 95 73 96 
<< m1 >>
rect 84 95 85 96 
<< m1 >>
rect 88 95 89 96 
<< m1 >>
rect 90 95 91 96 
<< m1 >>
rect 91 95 92 96 
<< m1 >>
rect 92 95 93 96 
<< m1 >>
rect 93 95 94 96 
<< m1 >>
rect 94 95 95 96 
<< m1 >>
rect 95 95 96 96 
<< m1 >>
rect 96 95 97 96 
<< m1 >>
rect 97 95 98 96 
<< m1 >>
rect 98 95 99 96 
<< m2 >>
rect 98 95 99 96 
<< m2c >>
rect 98 95 99 96 
<< m1 >>
rect 98 95 99 96 
<< m2 >>
rect 98 95 99 96 
<< m2 >>
rect 99 95 100 96 
<< m1 >>
rect 100 95 101 96 
<< m2 >>
rect 100 95 101 96 
<< m2 >>
rect 101 95 102 96 
<< m1 >>
rect 102 95 103 96 
<< m2 >>
rect 102 95 103 96 
<< m2c >>
rect 102 95 103 96 
<< m1 >>
rect 102 95 103 96 
<< m2 >>
rect 102 95 103 96 
<< m1 >>
rect 103 95 104 96 
<< m1 >>
rect 109 95 110 96 
<< m2 >>
rect 109 95 110 96 
<< m1 >>
rect 114 95 115 96 
<< m1 >>
rect 118 95 119 96 
<< m1 >>
rect 10 96 11 97 
<< m1 >>
rect 11 96 12 97 
<< m1 >>
rect 12 96 13 97 
<< m1 >>
rect 13 96 14 97 
<< m1 >>
rect 14 96 15 97 
<< m1 >>
rect 15 96 16 97 
<< m1 >>
rect 16 96 17 97 
<< m1 >>
rect 17 96 18 97 
<< m1 >>
rect 18 96 19 97 
<< m1 >>
rect 19 96 20 97 
<< m1 >>
rect 20 96 21 97 
<< m1 >>
rect 21 96 22 97 
<< m1 >>
rect 22 96 23 97 
<< m1 >>
rect 23 96 24 97 
<< m1 >>
rect 24 96 25 97 
<< m1 >>
rect 25 96 26 97 
<< m1 >>
rect 26 96 27 97 
<< m2 >>
rect 26 96 27 97 
<< m2c >>
rect 26 96 27 97 
<< m1 >>
rect 26 96 27 97 
<< m2 >>
rect 26 96 27 97 
<< m2 >>
rect 27 96 28 97 
<< m1 >>
rect 28 96 29 97 
<< m2 >>
rect 28 96 29 97 
<< m2 >>
rect 29 96 30 97 
<< m1 >>
rect 30 96 31 97 
<< m2 >>
rect 30 96 31 97 
<< m2c >>
rect 30 96 31 97 
<< m1 >>
rect 30 96 31 97 
<< m2 >>
rect 30 96 31 97 
<< m1 >>
rect 31 96 32 97 
<< m1 >>
rect 32 96 33 97 
<< m1 >>
rect 42 96 43 97 
<< m2 >>
rect 42 96 43 97 
<< m2c >>
rect 42 96 43 97 
<< m1 >>
rect 42 96 43 97 
<< m2 >>
rect 42 96 43 97 
<< m1 >>
rect 44 96 45 97 
<< m2 >>
rect 44 96 45 97 
<< m2c >>
rect 44 96 45 97 
<< m1 >>
rect 44 96 45 97 
<< m2 >>
rect 44 96 45 97 
<< m1 >>
rect 56 96 57 97 
<< m2 >>
rect 56 96 57 97 
<< m2c >>
rect 56 96 57 97 
<< m1 >>
rect 56 96 57 97 
<< m2 >>
rect 56 96 57 97 
<< m1 >>
rect 58 96 59 97 
<< m2 >>
rect 58 96 59 97 
<< m2c >>
rect 58 96 59 97 
<< m1 >>
rect 58 96 59 97 
<< m2 >>
rect 58 96 59 97 
<< m1 >>
rect 59 96 60 97 
<< m1 >>
rect 60 96 61 97 
<< m2 >>
rect 60 96 61 97 
<< m1 >>
rect 61 96 62 97 
<< m1 >>
rect 62 96 63 97 
<< m2 >>
rect 62 96 63 97 
<< m1 >>
rect 63 96 64 97 
<< m1 >>
rect 64 96 65 97 
<< m1 >>
rect 65 96 66 97 
<< m1 >>
rect 66 96 67 97 
<< m1 >>
rect 67 96 68 97 
<< m1 >>
rect 68 96 69 97 
<< m1 >>
rect 84 96 85 97 
<< m1 >>
rect 88 96 89 97 
<< m1 >>
rect 100 96 101 97 
<< m1 >>
rect 103 96 104 97 
<< m1 >>
rect 109 96 110 97 
<< m2 >>
rect 109 96 110 97 
<< m1 >>
rect 114 96 115 97 
<< m1 >>
rect 118 96 119 97 
<< m1 >>
rect 28 97 29 98 
<< m1 >>
rect 32 97 33 98 
<< m1 >>
rect 42 97 43 98 
<< m1 >>
rect 44 97 45 98 
<< m1 >>
rect 56 97 57 98 
<< m2 >>
rect 60 97 61 98 
<< m2 >>
rect 62 97 63 98 
<< m1 >>
rect 68 97 69 98 
<< m2 >>
rect 68 97 69 98 
<< m2c >>
rect 68 97 69 98 
<< m1 >>
rect 68 97 69 98 
<< m2 >>
rect 68 97 69 98 
<< m1 >>
rect 84 97 85 98 
<< m1 >>
rect 88 97 89 98 
<< m1 >>
rect 100 97 101 98 
<< m1 >>
rect 103 97 104 98 
<< m1 >>
rect 109 97 110 98 
<< m2 >>
rect 109 97 110 98 
<< m1 >>
rect 114 97 115 98 
<< m1 >>
rect 118 97 119 98 
<< m1 >>
rect 28 98 29 99 
<< m1 >>
rect 32 98 33 99 
<< m1 >>
rect 33 98 34 99 
<< m1 >>
rect 34 98 35 99 
<< m1 >>
rect 35 98 36 99 
<< m1 >>
rect 36 98 37 99 
<< m1 >>
rect 37 98 38 99 
<< m1 >>
rect 38 98 39 99 
<< m1 >>
rect 39 98 40 99 
<< m1 >>
rect 40 98 41 99 
<< m2 >>
rect 40 98 41 99 
<< m2c >>
rect 40 98 41 99 
<< m1 >>
rect 40 98 41 99 
<< m2 >>
rect 40 98 41 99 
<< m2 >>
rect 41 98 42 99 
<< m1 >>
rect 42 98 43 99 
<< m1 >>
rect 44 98 45 99 
<< m1 >>
rect 56 98 57 99 
<< m1 >>
rect 60 98 61 99 
<< m2 >>
rect 60 98 61 99 
<< m2c >>
rect 60 98 61 99 
<< m1 >>
rect 60 98 61 99 
<< m2 >>
rect 60 98 61 99 
<< m1 >>
rect 62 98 63 99 
<< m2 >>
rect 62 98 63 99 
<< m2c >>
rect 62 98 63 99 
<< m1 >>
rect 62 98 63 99 
<< m2 >>
rect 62 98 63 99 
<< m2 >>
rect 68 98 69 99 
<< m2 >>
rect 69 98 70 99 
<< m2 >>
rect 70 98 71 99 
<< m2 >>
rect 82 98 83 99 
<< m2 >>
rect 83 98 84 99 
<< m1 >>
rect 84 98 85 99 
<< m2 >>
rect 84 98 85 99 
<< m2c >>
rect 84 98 85 99 
<< m1 >>
rect 84 98 85 99 
<< m2 >>
rect 84 98 85 99 
<< m1 >>
rect 88 98 89 99 
<< m1 >>
rect 100 98 101 99 
<< m1 >>
rect 103 98 104 99 
<< m1 >>
rect 109 98 110 99 
<< m2 >>
rect 109 98 110 99 
<< m1 >>
rect 114 98 115 99 
<< m1 >>
rect 118 98 119 99 
<< m1 >>
rect 28 99 29 100 
<< m2 >>
rect 41 99 42 100 
<< m1 >>
rect 42 99 43 100 
<< m1 >>
rect 44 99 45 100 
<< m1 >>
rect 49 99 50 100 
<< m1 >>
rect 50 99 51 100 
<< m1 >>
rect 51 99 52 100 
<< m1 >>
rect 52 99 53 100 
<< m1 >>
rect 53 99 54 100 
<< m1 >>
rect 54 99 55 100 
<< m2 >>
rect 54 99 55 100 
<< m2c >>
rect 54 99 55 100 
<< m1 >>
rect 54 99 55 100 
<< m2 >>
rect 54 99 55 100 
<< m2 >>
rect 55 99 56 100 
<< m1 >>
rect 56 99 57 100 
<< m1 >>
rect 60 99 61 100 
<< m1 >>
rect 62 99 63 100 
<< m1 >>
rect 67 99 68 100 
<< m1 >>
rect 68 99 69 100 
<< m1 >>
rect 69 99 70 100 
<< m1 >>
rect 70 99 71 100 
<< m2 >>
rect 70 99 71 100 
<< m1 >>
rect 71 99 72 100 
<< m1 >>
rect 72 99 73 100 
<< m1 >>
rect 73 99 74 100 
<< m1 >>
rect 74 99 75 100 
<< m1 >>
rect 75 99 76 100 
<< m1 >>
rect 76 99 77 100 
<< m1 >>
rect 77 99 78 100 
<< m1 >>
rect 78 99 79 100 
<< m1 >>
rect 79 99 80 100 
<< m1 >>
rect 80 99 81 100 
<< m1 >>
rect 81 99 82 100 
<< m1 >>
rect 82 99 83 100 
<< m2 >>
rect 82 99 83 100 
<< m1 >>
rect 88 99 89 100 
<< m1 >>
rect 100 99 101 100 
<< m1 >>
rect 103 99 104 100 
<< m1 >>
rect 109 99 110 100 
<< m2 >>
rect 109 99 110 100 
<< m1 >>
rect 114 99 115 100 
<< m1 >>
rect 118 99 119 100 
<< m1 >>
rect 28 100 29 101 
<< m2 >>
rect 41 100 42 101 
<< m1 >>
rect 42 100 43 101 
<< m1 >>
rect 44 100 45 101 
<< m1 >>
rect 49 100 50 101 
<< m2 >>
rect 55 100 56 101 
<< m1 >>
rect 56 100 57 101 
<< m1 >>
rect 60 100 61 101 
<< m1 >>
rect 62 100 63 101 
<< m1 >>
rect 67 100 68 101 
<< m2 >>
rect 70 100 71 101 
<< m1 >>
rect 82 100 83 101 
<< m2 >>
rect 82 100 83 101 
<< m1 >>
rect 88 100 89 101 
<< m1 >>
rect 100 100 101 101 
<< m1 >>
rect 103 100 104 101 
<< m1 >>
rect 109 100 110 101 
<< m2 >>
rect 109 100 110 101 
<< m1 >>
rect 114 100 115 101 
<< m1 >>
rect 118 100 119 101 
<< m1 >>
rect 28 101 29 102 
<< m2 >>
rect 41 101 42 102 
<< m1 >>
rect 42 101 43 102 
<< m1 >>
rect 44 101 45 102 
<< m1 >>
rect 49 101 50 102 
<< m2 >>
rect 55 101 56 102 
<< m1 >>
rect 56 101 57 102 
<< m1 >>
rect 60 101 61 102 
<< m1 >>
rect 62 101 63 102 
<< m1 >>
rect 67 101 68 102 
<< m1 >>
rect 70 101 71 102 
<< m2 >>
rect 70 101 71 102 
<< m2c >>
rect 70 101 71 102 
<< m1 >>
rect 70 101 71 102 
<< m2 >>
rect 70 101 71 102 
<< m1 >>
rect 80 101 81 102 
<< m2 >>
rect 80 101 81 102 
<< m2c >>
rect 80 101 81 102 
<< m1 >>
rect 80 101 81 102 
<< m2 >>
rect 80 101 81 102 
<< m2 >>
rect 81 101 82 102 
<< m1 >>
rect 82 101 83 102 
<< m2 >>
rect 82 101 83 102 
<< m1 >>
rect 88 101 89 102 
<< m1 >>
rect 100 101 101 102 
<< m1 >>
rect 103 101 104 102 
<< m1 >>
rect 109 101 110 102 
<< m2 >>
rect 109 101 110 102 
<< m1 >>
rect 114 101 115 102 
<< m1 >>
rect 118 101 119 102 
<< pdiffusion >>
rect 12 102 13 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< m1 >>
rect 28 102 29 103 
<< pdiffusion >>
rect 30 102 31 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< pdiffusion >>
rect 33 102 34 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< m2 >>
rect 41 102 42 103 
<< m1 >>
rect 42 102 43 103 
<< m1 >>
rect 44 102 45 103 
<< pdiffusion >>
rect 48 102 49 103 
<< m1 >>
rect 49 102 50 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m2 >>
rect 55 102 56 103 
<< m1 >>
rect 56 102 57 103 
<< m1 >>
rect 60 102 61 103 
<< m1 >>
rect 62 102 63 103 
<< pdiffusion >>
rect 66 102 67 103 
<< m1 >>
rect 67 102 68 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< m1 >>
rect 70 102 71 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< m1 >>
rect 80 102 81 103 
<< m1 >>
rect 82 102 83 103 
<< pdiffusion >>
rect 84 102 85 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< m1 >>
rect 88 102 89 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< m1 >>
rect 100 102 101 103 
<< pdiffusion >>
rect 102 102 103 103 
<< m1 >>
rect 103 102 104 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< m1 >>
rect 109 102 110 103 
<< m2 >>
rect 109 102 110 103 
<< m1 >>
rect 114 102 115 103 
<< m1 >>
rect 118 102 119 103 
<< pdiffusion >>
rect 120 102 121 103 
<< pdiffusion >>
rect 121 102 122 103 
<< pdiffusion >>
rect 122 102 123 103 
<< pdiffusion >>
rect 123 102 124 103 
<< pdiffusion >>
rect 124 102 125 103 
<< pdiffusion >>
rect 125 102 126 103 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< m1 >>
rect 28 103 29 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< m2 >>
rect 41 103 42 104 
<< m1 >>
rect 42 103 43 104 
<< m1 >>
rect 44 103 45 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m2 >>
rect 55 103 56 104 
<< m1 >>
rect 56 103 57 104 
<< m1 >>
rect 60 103 61 104 
<< m1 >>
rect 62 103 63 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< m1 >>
rect 80 103 81 104 
<< m1 >>
rect 82 103 83 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< m1 >>
rect 100 103 101 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< m1 >>
rect 109 103 110 104 
<< m2 >>
rect 109 103 110 104 
<< m1 >>
rect 114 103 115 104 
<< m1 >>
rect 118 103 119 104 
<< pdiffusion >>
rect 120 103 121 104 
<< pdiffusion >>
rect 121 103 122 104 
<< pdiffusion >>
rect 122 103 123 104 
<< pdiffusion >>
rect 123 103 124 104 
<< pdiffusion >>
rect 124 103 125 104 
<< pdiffusion >>
rect 125 103 126 104 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< m1 >>
rect 28 104 29 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< m2 >>
rect 41 104 42 105 
<< m1 >>
rect 42 104 43 105 
<< m1 >>
rect 44 104 45 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m2 >>
rect 55 104 56 105 
<< m1 >>
rect 56 104 57 105 
<< m1 >>
rect 60 104 61 105 
<< m1 >>
rect 62 104 63 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< m1 >>
rect 80 104 81 105 
<< m1 >>
rect 82 104 83 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< m1 >>
rect 100 104 101 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< m1 >>
rect 109 104 110 105 
<< m2 >>
rect 109 104 110 105 
<< m1 >>
rect 114 104 115 105 
<< m1 >>
rect 118 104 119 105 
<< pdiffusion >>
rect 120 104 121 105 
<< pdiffusion >>
rect 121 104 122 105 
<< pdiffusion >>
rect 122 104 123 105 
<< pdiffusion >>
rect 123 104 124 105 
<< pdiffusion >>
rect 124 104 125 105 
<< pdiffusion >>
rect 125 104 126 105 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< m1 >>
rect 28 105 29 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< m2 >>
rect 41 105 42 106 
<< m1 >>
rect 42 105 43 106 
<< m1 >>
rect 44 105 45 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m2 >>
rect 55 105 56 106 
<< m1 >>
rect 56 105 57 106 
<< m1 >>
rect 60 105 61 106 
<< m1 >>
rect 62 105 63 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< m1 >>
rect 80 105 81 106 
<< m1 >>
rect 82 105 83 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< m1 >>
rect 100 105 101 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< m1 >>
rect 109 105 110 106 
<< m2 >>
rect 109 105 110 106 
<< m1 >>
rect 114 105 115 106 
<< m1 >>
rect 118 105 119 106 
<< pdiffusion >>
rect 120 105 121 106 
<< pdiffusion >>
rect 121 105 122 106 
<< pdiffusion >>
rect 122 105 123 106 
<< pdiffusion >>
rect 123 105 124 106 
<< pdiffusion >>
rect 124 105 125 106 
<< pdiffusion >>
rect 125 105 126 106 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< m1 >>
rect 28 106 29 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< m2 >>
rect 41 106 42 107 
<< m1 >>
rect 42 106 43 107 
<< m1 >>
rect 44 106 45 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m2 >>
rect 55 106 56 107 
<< m1 >>
rect 56 106 57 107 
<< m1 >>
rect 60 106 61 107 
<< m1 >>
rect 62 106 63 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< m1 >>
rect 80 106 81 107 
<< m1 >>
rect 82 106 83 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< m1 >>
rect 100 106 101 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< m1 >>
rect 109 106 110 107 
<< m2 >>
rect 109 106 110 107 
<< m1 >>
rect 114 106 115 107 
<< m1 >>
rect 118 106 119 107 
<< pdiffusion >>
rect 120 106 121 107 
<< pdiffusion >>
rect 121 106 122 107 
<< pdiffusion >>
rect 122 106 123 107 
<< pdiffusion >>
rect 123 106 124 107 
<< pdiffusion >>
rect 124 106 125 107 
<< pdiffusion >>
rect 125 106 126 107 
<< pdiffusion >>
rect 12 107 13 108 
<< m1 >>
rect 13 107 14 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< m1 >>
rect 28 107 29 108 
<< pdiffusion >>
rect 30 107 31 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< m1 >>
rect 34 107 35 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< m2 >>
rect 41 107 42 108 
<< m1 >>
rect 42 107 43 108 
<< m1 >>
rect 44 107 45 108 
<< pdiffusion >>
rect 48 107 49 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m2 >>
rect 55 107 56 108 
<< m1 >>
rect 56 107 57 108 
<< m1 >>
rect 60 107 61 108 
<< m1 >>
rect 62 107 63 108 
<< pdiffusion >>
rect 66 107 67 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< m1 >>
rect 80 107 81 108 
<< m1 >>
rect 82 107 83 108 
<< pdiffusion >>
rect 84 107 85 108 
<< m1 >>
rect 85 107 86 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< m1 >>
rect 100 107 101 108 
<< pdiffusion >>
rect 102 107 103 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< m1 >>
rect 106 107 107 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< m1 >>
rect 109 107 110 108 
<< m2 >>
rect 109 107 110 108 
<< m1 >>
rect 114 107 115 108 
<< m1 >>
rect 118 107 119 108 
<< pdiffusion >>
rect 120 107 121 108 
<< pdiffusion >>
rect 121 107 122 108 
<< pdiffusion >>
rect 122 107 123 108 
<< pdiffusion >>
rect 123 107 124 108 
<< m1 >>
rect 124 107 125 108 
<< pdiffusion >>
rect 124 107 125 108 
<< pdiffusion >>
rect 125 107 126 108 
<< m1 >>
rect 13 108 14 109 
<< m1 >>
rect 28 108 29 109 
<< m1 >>
rect 34 108 35 109 
<< m2 >>
rect 41 108 42 109 
<< m1 >>
rect 42 108 43 109 
<< m1 >>
rect 44 108 45 109 
<< m2 >>
rect 55 108 56 109 
<< m1 >>
rect 56 108 57 109 
<< m1 >>
rect 60 108 61 109 
<< m1 >>
rect 62 108 63 109 
<< m1 >>
rect 80 108 81 109 
<< m1 >>
rect 82 108 83 109 
<< m1 >>
rect 85 108 86 109 
<< m1 >>
rect 100 108 101 109 
<< m1 >>
rect 106 108 107 109 
<< m1 >>
rect 109 108 110 109 
<< m2 >>
rect 109 108 110 109 
<< m1 >>
rect 114 108 115 109 
<< m1 >>
rect 118 108 119 109 
<< m2 >>
rect 118 108 119 109 
<< m2c >>
rect 118 108 119 109 
<< m1 >>
rect 118 108 119 109 
<< m2 >>
rect 118 108 119 109 
<< m1 >>
rect 124 108 125 109 
<< m1 >>
rect 13 109 14 110 
<< m1 >>
rect 28 109 29 110 
<< m1 >>
rect 34 109 35 110 
<< m2 >>
rect 41 109 42 110 
<< m1 >>
rect 42 109 43 110 
<< m1 >>
rect 44 109 45 110 
<< m2 >>
rect 55 109 56 110 
<< m1 >>
rect 56 109 57 110 
<< m1 >>
rect 60 109 61 110 
<< m1 >>
rect 62 109 63 110 
<< m1 >>
rect 80 109 81 110 
<< m1 >>
rect 82 109 83 110 
<< m1 >>
rect 85 109 86 110 
<< m1 >>
rect 100 109 101 110 
<< m1 >>
rect 106 109 107 110 
<< m1 >>
rect 107 109 108 110 
<< m1 >>
rect 108 109 109 110 
<< m1 >>
rect 109 109 110 110 
<< m2 >>
rect 109 109 110 110 
<< m1 >>
rect 114 109 115 110 
<< m2 >>
rect 118 109 119 110 
<< m1 >>
rect 124 109 125 110 
<< m1 >>
rect 13 110 14 111 
<< m1 >>
rect 28 110 29 111 
<< m1 >>
rect 34 110 35 111 
<< m2 >>
rect 41 110 42 111 
<< m1 >>
rect 42 110 43 111 
<< m1 >>
rect 44 110 45 111 
<< m2 >>
rect 55 110 56 111 
<< m1 >>
rect 56 110 57 111 
<< m1 >>
rect 60 110 61 111 
<< m1 >>
rect 62 110 63 111 
<< m1 >>
rect 70 110 71 111 
<< m1 >>
rect 71 110 72 111 
<< m1 >>
rect 72 110 73 111 
<< m1 >>
rect 73 110 74 111 
<< m1 >>
rect 74 110 75 111 
<< m1 >>
rect 75 110 76 111 
<< m1 >>
rect 76 110 77 111 
<< m1 >>
rect 77 110 78 111 
<< m1 >>
rect 78 110 79 111 
<< m1 >>
rect 79 110 80 111 
<< m1 >>
rect 80 110 81 111 
<< m1 >>
rect 82 110 83 111 
<< m1 >>
rect 85 110 86 111 
<< m1 >>
rect 86 110 87 111 
<< m1 >>
rect 87 110 88 111 
<< m1 >>
rect 88 110 89 111 
<< m1 >>
rect 89 110 90 111 
<< m1 >>
rect 90 110 91 111 
<< m1 >>
rect 91 110 92 111 
<< m1 >>
rect 92 110 93 111 
<< m1 >>
rect 93 110 94 111 
<< m1 >>
rect 94 110 95 111 
<< m1 >>
rect 95 110 96 111 
<< m1 >>
rect 96 110 97 111 
<< m1 >>
rect 97 110 98 111 
<< m1 >>
rect 98 110 99 111 
<< m1 >>
rect 99 110 100 111 
<< m1 >>
rect 100 110 101 111 
<< m2 >>
rect 109 110 110 111 
<< m1 >>
rect 114 110 115 111 
<< m1 >>
rect 115 110 116 111 
<< m1 >>
rect 116 110 117 111 
<< m1 >>
rect 117 110 118 111 
<< m1 >>
rect 118 110 119 111 
<< m2 >>
rect 118 110 119 111 
<< m1 >>
rect 119 110 120 111 
<< m1 >>
rect 120 110 121 111 
<< m2 >>
rect 120 110 121 111 
<< m2c >>
rect 120 110 121 111 
<< m1 >>
rect 120 110 121 111 
<< m2 >>
rect 120 110 121 111 
<< m1 >>
rect 124 110 125 111 
<< m1 >>
rect 13 111 14 112 
<< m1 >>
rect 28 111 29 112 
<< m1 >>
rect 34 111 35 112 
<< m2 >>
rect 41 111 42 112 
<< m1 >>
rect 42 111 43 112 
<< m1 >>
rect 44 111 45 112 
<< m2 >>
rect 55 111 56 112 
<< m1 >>
rect 56 111 57 112 
<< m1 >>
rect 60 111 61 112 
<< m1 >>
rect 62 111 63 112 
<< m1 >>
rect 70 111 71 112 
<< m1 >>
rect 82 111 83 112 
<< m2 >>
rect 109 111 110 112 
<< m2 >>
rect 118 111 119 112 
<< m2 >>
rect 120 111 121 112 
<< m1 >>
rect 124 111 125 112 
<< m1 >>
rect 13 112 14 113 
<< m1 >>
rect 14 112 15 113 
<< m1 >>
rect 15 112 16 113 
<< m1 >>
rect 16 112 17 113 
<< m1 >>
rect 17 112 18 113 
<< m1 >>
rect 18 112 19 113 
<< m1 >>
rect 19 112 20 113 
<< m1 >>
rect 20 112 21 113 
<< m1 >>
rect 21 112 22 113 
<< m1 >>
rect 22 112 23 113 
<< m1 >>
rect 23 112 24 113 
<< m1 >>
rect 24 112 25 113 
<< m1 >>
rect 25 112 26 113 
<< m1 >>
rect 26 112 27 113 
<< m2 >>
rect 26 112 27 113 
<< m2c >>
rect 26 112 27 113 
<< m1 >>
rect 26 112 27 113 
<< m2 >>
rect 26 112 27 113 
<< m2 >>
rect 27 112 28 113 
<< m1 >>
rect 28 112 29 113 
<< m2 >>
rect 28 112 29 113 
<< m2 >>
rect 29 112 30 113 
<< m1 >>
rect 30 112 31 113 
<< m2 >>
rect 30 112 31 113 
<< m2c >>
rect 30 112 31 113 
<< m1 >>
rect 30 112 31 113 
<< m2 >>
rect 30 112 31 113 
<< m1 >>
rect 31 112 32 113 
<< m1 >>
rect 32 112 33 113 
<< m1 >>
rect 33 112 34 113 
<< m1 >>
rect 34 112 35 113 
<< m2 >>
rect 41 112 42 113 
<< m1 >>
rect 42 112 43 113 
<< m1 >>
rect 44 112 45 113 
<< m2 >>
rect 55 112 56 113 
<< m1 >>
rect 56 112 57 113 
<< m1 >>
rect 60 112 61 113 
<< m1 >>
rect 62 112 63 113 
<< m1 >>
rect 70 112 71 113 
<< m1 >>
rect 82 112 83 113 
<< m1 >>
rect 83 112 84 113 
<< m1 >>
rect 84 112 85 113 
<< m1 >>
rect 85 112 86 113 
<< m1 >>
rect 86 112 87 113 
<< m1 >>
rect 87 112 88 113 
<< m1 >>
rect 88 112 89 113 
<< m1 >>
rect 89 112 90 113 
<< m1 >>
rect 90 112 91 113 
<< m1 >>
rect 91 112 92 113 
<< m1 >>
rect 92 112 93 113 
<< m1 >>
rect 93 112 94 113 
<< m1 >>
rect 94 112 95 113 
<< m1 >>
rect 95 112 96 113 
<< m1 >>
rect 96 112 97 113 
<< m1 >>
rect 97 112 98 113 
<< m1 >>
rect 98 112 99 113 
<< m1 >>
rect 99 112 100 113 
<< m1 >>
rect 100 112 101 113 
<< m1 >>
rect 101 112 102 113 
<< m1 >>
rect 102 112 103 113 
<< m1 >>
rect 103 112 104 113 
<< m1 >>
rect 104 112 105 113 
<< m1 >>
rect 105 112 106 113 
<< m1 >>
rect 106 112 107 113 
<< m1 >>
rect 107 112 108 113 
<< m1 >>
rect 108 112 109 113 
<< m1 >>
rect 109 112 110 113 
<< m2 >>
rect 109 112 110 113 
<< m1 >>
rect 110 112 111 113 
<< m1 >>
rect 111 112 112 113 
<< m1 >>
rect 112 112 113 113 
<< m1 >>
rect 113 112 114 113 
<< m1 >>
rect 114 112 115 113 
<< m1 >>
rect 115 112 116 113 
<< m1 >>
rect 116 112 117 113 
<< m1 >>
rect 117 112 118 113 
<< m1 >>
rect 118 112 119 113 
<< m2 >>
rect 118 112 119 113 
<< m1 >>
rect 119 112 120 113 
<< m1 >>
rect 120 112 121 113 
<< m2 >>
rect 120 112 121 113 
<< m1 >>
rect 121 112 122 113 
<< m1 >>
rect 122 112 123 113 
<< m1 >>
rect 123 112 124 113 
<< m1 >>
rect 124 112 125 113 
<< m1 >>
rect 28 113 29 114 
<< m2 >>
rect 41 113 42 114 
<< m1 >>
rect 42 113 43 114 
<< m1 >>
rect 44 113 45 114 
<< m2 >>
rect 55 113 56 114 
<< m1 >>
rect 56 113 57 114 
<< m2 >>
rect 57 113 58 114 
<< m1 >>
rect 58 113 59 114 
<< m2 >>
rect 58 113 59 114 
<< m2c >>
rect 58 113 59 114 
<< m1 >>
rect 58 113 59 114 
<< m2 >>
rect 58 113 59 114 
<< m1 >>
rect 59 113 60 114 
<< m1 >>
rect 60 113 61 114 
<< m2 >>
rect 60 113 61 114 
<< m2 >>
rect 61 113 62 114 
<< m1 >>
rect 62 113 63 114 
<< m2 >>
rect 62 113 63 114 
<< m2c >>
rect 62 113 63 114 
<< m1 >>
rect 62 113 63 114 
<< m2 >>
rect 62 113 63 114 
<< m1 >>
rect 70 113 71 114 
<< m2 >>
rect 109 113 110 114 
<< m2 >>
rect 118 113 119 114 
<< m2 >>
rect 120 113 121 114 
<< m2 >>
rect 121 113 122 114 
<< m2 >>
rect 122 113 123 114 
<< m2 >>
rect 123 113 124 114 
<< m2 >>
rect 124 113 125 114 
<< m1 >>
rect 28 114 29 115 
<< m2 >>
rect 41 114 42 115 
<< m1 >>
rect 42 114 43 115 
<< m1 >>
rect 44 114 45 115 
<< m2 >>
rect 55 114 56 115 
<< m1 >>
rect 56 114 57 115 
<< m2 >>
rect 57 114 58 115 
<< m2 >>
rect 60 114 61 115 
<< m1 >>
rect 70 114 71 115 
<< m2 >>
rect 109 114 110 115 
<< m2 >>
rect 118 114 119 115 
<< m1 >>
rect 124 114 125 115 
<< m2 >>
rect 124 114 125 115 
<< m2c >>
rect 124 114 125 115 
<< m1 >>
rect 124 114 125 115 
<< m2 >>
rect 124 114 125 115 
<< m1 >>
rect 28 115 29 116 
<< m2 >>
rect 41 115 42 116 
<< m1 >>
rect 42 115 43 116 
<< m1 >>
rect 44 115 45 116 
<< m2 >>
rect 55 115 56 116 
<< m1 >>
rect 56 115 57 116 
<< m1 >>
rect 57 115 58 116 
<< m2 >>
rect 57 115 58 116 
<< m1 >>
rect 58 115 59 116 
<< m1 >>
rect 59 115 60 116 
<< m1 >>
rect 60 115 61 116 
<< m2 >>
rect 60 115 61 116 
<< m1 >>
rect 61 115 62 116 
<< m1 >>
rect 62 115 63 116 
<< m1 >>
rect 63 115 64 116 
<< m1 >>
rect 64 115 65 116 
<< m1 >>
rect 65 115 66 116 
<< m1 >>
rect 66 115 67 116 
<< m1 >>
rect 67 115 68 116 
<< m1 >>
rect 68 115 69 116 
<< m2 >>
rect 68 115 69 116 
<< m2c >>
rect 68 115 69 116 
<< m1 >>
rect 68 115 69 116 
<< m2 >>
rect 68 115 69 116 
<< m2 >>
rect 69 115 70 116 
<< m1 >>
rect 70 115 71 116 
<< m2 >>
rect 70 115 71 116 
<< m2 >>
rect 71 115 72 116 
<< m1 >>
rect 72 115 73 116 
<< m2 >>
rect 72 115 73 116 
<< m2c >>
rect 72 115 73 116 
<< m1 >>
rect 72 115 73 116 
<< m2 >>
rect 72 115 73 116 
<< m1 >>
rect 73 115 74 116 
<< m1 >>
rect 74 115 75 116 
<< m1 >>
rect 75 115 76 116 
<< m1 >>
rect 76 115 77 116 
<< m1 >>
rect 77 115 78 116 
<< m1 >>
rect 78 115 79 116 
<< m1 >>
rect 79 115 80 116 
<< m1 >>
rect 80 115 81 116 
<< m1 >>
rect 81 115 82 116 
<< m1 >>
rect 82 115 83 116 
<< m1 >>
rect 83 115 84 116 
<< m1 >>
rect 84 115 85 116 
<< m1 >>
rect 85 115 86 116 
<< m1 >>
rect 86 115 87 116 
<< m1 >>
rect 87 115 88 116 
<< m1 >>
rect 88 115 89 116 
<< m1 >>
rect 89 115 90 116 
<< m1 >>
rect 90 115 91 116 
<< m1 >>
rect 91 115 92 116 
<< m1 >>
rect 92 115 93 116 
<< m1 >>
rect 93 115 94 116 
<< m1 >>
rect 94 115 95 116 
<< m1 >>
rect 95 115 96 116 
<< m1 >>
rect 96 115 97 116 
<< m1 >>
rect 97 115 98 116 
<< m1 >>
rect 98 115 99 116 
<< m1 >>
rect 99 115 100 116 
<< m1 >>
rect 100 115 101 116 
<< m1 >>
rect 101 115 102 116 
<< m1 >>
rect 102 115 103 116 
<< m1 >>
rect 103 115 104 116 
<< m1 >>
rect 104 115 105 116 
<< m1 >>
rect 105 115 106 116 
<< m1 >>
rect 106 115 107 116 
<< m1 >>
rect 107 115 108 116 
<< m1 >>
rect 108 115 109 116 
<< m1 >>
rect 109 115 110 116 
<< m2 >>
rect 109 115 110 116 
<< m1 >>
rect 110 115 111 116 
<< m1 >>
rect 111 115 112 116 
<< m1 >>
rect 112 115 113 116 
<< m1 >>
rect 113 115 114 116 
<< m1 >>
rect 114 115 115 116 
<< m1 >>
rect 115 115 116 116 
<< m1 >>
rect 116 115 117 116 
<< m1 >>
rect 117 115 118 116 
<< m1 >>
rect 118 115 119 116 
<< m2 >>
rect 118 115 119 116 
<< m1 >>
rect 119 115 120 116 
<< m1 >>
rect 120 115 121 116 
<< m1 >>
rect 121 115 122 116 
<< m1 >>
rect 124 115 125 116 
<< m1 >>
rect 28 116 29 117 
<< m2 >>
rect 41 116 42 117 
<< m1 >>
rect 42 116 43 117 
<< m1 >>
rect 44 116 45 117 
<< m2 >>
rect 55 116 56 117 
<< m2 >>
rect 57 116 58 117 
<< m2 >>
rect 60 116 61 117 
<< m1 >>
rect 70 116 71 117 
<< m2 >>
rect 109 116 110 117 
<< m2 >>
rect 118 116 119 117 
<< m1 >>
rect 121 116 122 117 
<< m1 >>
rect 124 116 125 117 
<< m1 >>
rect 28 117 29 118 
<< m2 >>
rect 41 117 42 118 
<< m1 >>
rect 42 117 43 118 
<< m1 >>
rect 44 117 45 118 
<< m1 >>
rect 55 117 56 118 
<< m2 >>
rect 55 117 56 118 
<< m2c >>
rect 55 117 56 118 
<< m1 >>
rect 55 117 56 118 
<< m2 >>
rect 55 117 56 118 
<< m1 >>
rect 56 117 57 118 
<< m1 >>
rect 57 117 58 118 
<< m2 >>
rect 57 117 58 118 
<< m1 >>
rect 58 117 59 118 
<< m1 >>
rect 59 117 60 118 
<< m1 >>
rect 60 117 61 118 
<< m2 >>
rect 60 117 61 118 
<< m1 >>
rect 61 117 62 118 
<< m1 >>
rect 62 117 63 118 
<< m1 >>
rect 63 117 64 118 
<< m1 >>
rect 64 117 65 118 
<< m1 >>
rect 65 117 66 118 
<< m1 >>
rect 66 117 67 118 
<< m1 >>
rect 67 117 68 118 
<< m1 >>
rect 70 117 71 118 
<< m1 >>
rect 106 117 107 118 
<< m1 >>
rect 107 117 108 118 
<< m1 >>
rect 108 117 109 118 
<< m1 >>
rect 109 117 110 118 
<< m2 >>
rect 109 117 110 118 
<< m2c >>
rect 109 117 110 118 
<< m1 >>
rect 109 117 110 118 
<< m2 >>
rect 109 117 110 118 
<< m1 >>
rect 118 117 119 118 
<< m2 >>
rect 118 117 119 118 
<< m2c >>
rect 118 117 119 118 
<< m1 >>
rect 118 117 119 118 
<< m2 >>
rect 118 117 119 118 
<< m1 >>
rect 121 117 122 118 
<< m1 >>
rect 124 117 125 118 
<< m1 >>
rect 28 118 29 119 
<< m2 >>
rect 41 118 42 119 
<< m1 >>
rect 42 118 43 119 
<< m1 >>
rect 44 118 45 119 
<< m2 >>
rect 57 118 58 119 
<< m2 >>
rect 59 118 60 119 
<< m2 >>
rect 60 118 61 119 
<< m1 >>
rect 67 118 68 119 
<< m1 >>
rect 70 118 71 119 
<< m1 >>
rect 106 118 107 119 
<< m1 >>
rect 118 118 119 119 
<< m1 >>
rect 121 118 122 119 
<< m1 >>
rect 124 118 125 119 
<< m1 >>
rect 28 119 29 120 
<< m2 >>
rect 41 119 42 120 
<< m1 >>
rect 42 119 43 120 
<< m1 >>
rect 44 119 45 120 
<< m1 >>
rect 45 119 46 120 
<< m1 >>
rect 46 119 47 120 
<< m1 >>
rect 47 119 48 120 
<< m1 >>
rect 48 119 49 120 
<< m1 >>
rect 49 119 50 120 
<< m1 >>
rect 50 119 51 120 
<< m1 >>
rect 51 119 52 120 
<< m1 >>
rect 52 119 53 120 
<< m1 >>
rect 53 119 54 120 
<< m1 >>
rect 54 119 55 120 
<< m1 >>
rect 55 119 56 120 
<< m1 >>
rect 56 119 57 120 
<< m1 >>
rect 57 119 58 120 
<< m2 >>
rect 57 119 58 120 
<< m2c >>
rect 57 119 58 120 
<< m1 >>
rect 57 119 58 120 
<< m2 >>
rect 57 119 58 120 
<< m1 >>
rect 59 119 60 120 
<< m2 >>
rect 59 119 60 120 
<< m2c >>
rect 59 119 60 120 
<< m1 >>
rect 59 119 60 120 
<< m2 >>
rect 59 119 60 120 
<< m1 >>
rect 67 119 68 120 
<< m1 >>
rect 70 119 71 120 
<< m1 >>
rect 106 119 107 120 
<< m1 >>
rect 118 119 119 120 
<< m1 >>
rect 121 119 122 120 
<< m1 >>
rect 124 119 125 120 
<< pdiffusion >>
rect 12 120 13 121 
<< pdiffusion >>
rect 13 120 14 121 
<< pdiffusion >>
rect 14 120 15 121 
<< pdiffusion >>
rect 15 120 16 121 
<< pdiffusion >>
rect 16 120 17 121 
<< pdiffusion >>
rect 17 120 18 121 
<< m1 >>
rect 28 120 29 121 
<< pdiffusion >>
rect 30 120 31 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< m2 >>
rect 41 120 42 121 
<< m1 >>
rect 42 120 43 121 
<< m1 >>
rect 59 120 60 121 
<< pdiffusion >>
rect 66 120 67 121 
<< m1 >>
rect 67 120 68 121 
<< pdiffusion >>
rect 67 120 68 121 
<< pdiffusion >>
rect 68 120 69 121 
<< pdiffusion >>
rect 69 120 70 121 
<< m1 >>
rect 70 120 71 121 
<< pdiffusion >>
rect 70 120 71 121 
<< pdiffusion >>
rect 71 120 72 121 
<< pdiffusion >>
rect 102 120 103 121 
<< pdiffusion >>
rect 103 120 104 121 
<< pdiffusion >>
rect 104 120 105 121 
<< pdiffusion >>
rect 105 120 106 121 
<< m1 >>
rect 106 120 107 121 
<< pdiffusion >>
rect 106 120 107 121 
<< pdiffusion >>
rect 107 120 108 121 
<< m1 >>
rect 118 120 119 121 
<< pdiffusion >>
rect 120 120 121 121 
<< m1 >>
rect 121 120 122 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< m1 >>
rect 124 120 125 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< pdiffusion >>
rect 12 121 13 122 
<< pdiffusion >>
rect 13 121 14 122 
<< pdiffusion >>
rect 14 121 15 122 
<< pdiffusion >>
rect 15 121 16 122 
<< pdiffusion >>
rect 16 121 17 122 
<< pdiffusion >>
rect 17 121 18 122 
<< m1 >>
rect 28 121 29 122 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< m2 >>
rect 41 121 42 122 
<< m1 >>
rect 42 121 43 122 
<< m2 >>
rect 42 121 43 122 
<< m2 >>
rect 43 121 44 122 
<< m1 >>
rect 44 121 45 122 
<< m2 >>
rect 44 121 45 122 
<< m2c >>
rect 44 121 45 122 
<< m1 >>
rect 44 121 45 122 
<< m2 >>
rect 44 121 45 122 
<< m1 >>
rect 45 121 46 122 
<< m1 >>
rect 46 121 47 122 
<< m1 >>
rect 47 121 48 122 
<< m1 >>
rect 48 121 49 122 
<< m1 >>
rect 49 121 50 122 
<< m1 >>
rect 50 121 51 122 
<< m1 >>
rect 51 121 52 122 
<< m1 >>
rect 52 121 53 122 
<< m1 >>
rect 53 121 54 122 
<< m1 >>
rect 54 121 55 122 
<< m1 >>
rect 55 121 56 122 
<< m1 >>
rect 56 121 57 122 
<< m1 >>
rect 57 121 58 122 
<< m1 >>
rect 58 121 59 122 
<< m1 >>
rect 59 121 60 122 
<< pdiffusion >>
rect 66 121 67 122 
<< pdiffusion >>
rect 67 121 68 122 
<< pdiffusion >>
rect 68 121 69 122 
<< pdiffusion >>
rect 69 121 70 122 
<< pdiffusion >>
rect 70 121 71 122 
<< pdiffusion >>
rect 71 121 72 122 
<< pdiffusion >>
rect 102 121 103 122 
<< pdiffusion >>
rect 103 121 104 122 
<< pdiffusion >>
rect 104 121 105 122 
<< pdiffusion >>
rect 105 121 106 122 
<< pdiffusion >>
rect 106 121 107 122 
<< pdiffusion >>
rect 107 121 108 122 
<< m1 >>
rect 118 121 119 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< pdiffusion >>
rect 12 122 13 123 
<< pdiffusion >>
rect 13 122 14 123 
<< pdiffusion >>
rect 14 122 15 123 
<< pdiffusion >>
rect 15 122 16 123 
<< pdiffusion >>
rect 16 122 17 123 
<< pdiffusion >>
rect 17 122 18 123 
<< m1 >>
rect 28 122 29 123 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< m1 >>
rect 42 122 43 123 
<< pdiffusion >>
rect 66 122 67 123 
<< pdiffusion >>
rect 67 122 68 123 
<< pdiffusion >>
rect 68 122 69 123 
<< pdiffusion >>
rect 69 122 70 123 
<< pdiffusion >>
rect 70 122 71 123 
<< pdiffusion >>
rect 71 122 72 123 
<< pdiffusion >>
rect 102 122 103 123 
<< pdiffusion >>
rect 103 122 104 123 
<< pdiffusion >>
rect 104 122 105 123 
<< pdiffusion >>
rect 105 122 106 123 
<< pdiffusion >>
rect 106 122 107 123 
<< pdiffusion >>
rect 107 122 108 123 
<< m1 >>
rect 118 122 119 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< pdiffusion >>
rect 12 123 13 124 
<< pdiffusion >>
rect 13 123 14 124 
<< pdiffusion >>
rect 14 123 15 124 
<< pdiffusion >>
rect 15 123 16 124 
<< pdiffusion >>
rect 16 123 17 124 
<< pdiffusion >>
rect 17 123 18 124 
<< m1 >>
rect 28 123 29 124 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< m1 >>
rect 42 123 43 124 
<< pdiffusion >>
rect 66 123 67 124 
<< pdiffusion >>
rect 67 123 68 124 
<< pdiffusion >>
rect 68 123 69 124 
<< pdiffusion >>
rect 69 123 70 124 
<< pdiffusion >>
rect 70 123 71 124 
<< pdiffusion >>
rect 71 123 72 124 
<< pdiffusion >>
rect 102 123 103 124 
<< pdiffusion >>
rect 103 123 104 124 
<< pdiffusion >>
rect 104 123 105 124 
<< pdiffusion >>
rect 105 123 106 124 
<< pdiffusion >>
rect 106 123 107 124 
<< pdiffusion >>
rect 107 123 108 124 
<< m1 >>
rect 118 123 119 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< pdiffusion >>
rect 12 124 13 125 
<< pdiffusion >>
rect 13 124 14 125 
<< pdiffusion >>
rect 14 124 15 125 
<< pdiffusion >>
rect 15 124 16 125 
<< pdiffusion >>
rect 16 124 17 125 
<< pdiffusion >>
rect 17 124 18 125 
<< m1 >>
rect 28 124 29 125 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< m1 >>
rect 42 124 43 125 
<< pdiffusion >>
rect 66 124 67 125 
<< pdiffusion >>
rect 67 124 68 125 
<< pdiffusion >>
rect 68 124 69 125 
<< pdiffusion >>
rect 69 124 70 125 
<< pdiffusion >>
rect 70 124 71 125 
<< pdiffusion >>
rect 71 124 72 125 
<< pdiffusion >>
rect 102 124 103 125 
<< pdiffusion >>
rect 103 124 104 125 
<< pdiffusion >>
rect 104 124 105 125 
<< pdiffusion >>
rect 105 124 106 125 
<< pdiffusion >>
rect 106 124 107 125 
<< pdiffusion >>
rect 107 124 108 125 
<< m1 >>
rect 118 124 119 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< pdiffusion >>
rect 12 125 13 126 
<< m1 >>
rect 13 125 14 126 
<< pdiffusion >>
rect 13 125 14 126 
<< pdiffusion >>
rect 14 125 15 126 
<< pdiffusion >>
rect 15 125 16 126 
<< pdiffusion >>
rect 16 125 17 126 
<< pdiffusion >>
rect 17 125 18 126 
<< m1 >>
rect 28 125 29 126 
<< pdiffusion >>
rect 30 125 31 126 
<< m1 >>
rect 31 125 32 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< m1 >>
rect 42 125 43 126 
<< pdiffusion >>
rect 66 125 67 126 
<< pdiffusion >>
rect 67 125 68 126 
<< pdiffusion >>
rect 68 125 69 126 
<< pdiffusion >>
rect 69 125 70 126 
<< pdiffusion >>
rect 70 125 71 126 
<< pdiffusion >>
rect 71 125 72 126 
<< pdiffusion >>
rect 102 125 103 126 
<< pdiffusion >>
rect 103 125 104 126 
<< pdiffusion >>
rect 104 125 105 126 
<< pdiffusion >>
rect 105 125 106 126 
<< pdiffusion >>
rect 106 125 107 126 
<< pdiffusion >>
rect 107 125 108 126 
<< m1 >>
rect 118 125 119 126 
<< pdiffusion >>
rect 120 125 121 126 
<< m1 >>
rect 121 125 122 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< m1 >>
rect 13 126 14 127 
<< m1 >>
rect 28 126 29 127 
<< m1 >>
rect 31 126 32 127 
<< m1 >>
rect 42 126 43 127 
<< m1 >>
rect 118 126 119 127 
<< m1 >>
rect 121 126 122 127 
<< m1 >>
rect 13 127 14 128 
<< m1 >>
rect 28 127 29 128 
<< m1 >>
rect 31 127 32 128 
<< m1 >>
rect 42 127 43 128 
<< m1 >>
rect 118 127 119 128 
<< m1 >>
rect 119 127 120 128 
<< m1 >>
rect 120 127 121 128 
<< m1 >>
rect 121 127 122 128 
<< m1 >>
rect 13 128 14 129 
<< m1 >>
rect 14 128 15 129 
<< m1 >>
rect 15 128 16 129 
<< m1 >>
rect 16 128 17 129 
<< m1 >>
rect 17 128 18 129 
<< m1 >>
rect 18 128 19 129 
<< m1 >>
rect 19 128 20 129 
<< m1 >>
rect 20 128 21 129 
<< m1 >>
rect 21 128 22 129 
<< m1 >>
rect 22 128 23 129 
<< m1 >>
rect 23 128 24 129 
<< m1 >>
rect 24 128 25 129 
<< m1 >>
rect 25 128 26 129 
<< m1 >>
rect 26 128 27 129 
<< m1 >>
rect 27 128 28 129 
<< m1 >>
rect 28 128 29 129 
<< m1 >>
rect 31 128 32 129 
<< m1 >>
rect 32 128 33 129 
<< m1 >>
rect 33 128 34 129 
<< m1 >>
rect 34 128 35 129 
<< m1 >>
rect 35 128 36 129 
<< m1 >>
rect 36 128 37 129 
<< m1 >>
rect 37 128 38 129 
<< m1 >>
rect 38 128 39 129 
<< m1 >>
rect 39 128 40 129 
<< m1 >>
rect 40 128 41 129 
<< m1 >>
rect 41 128 42 129 
<< m1 >>
rect 42 128 43 129 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 1
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 103 84 104 85  0 t = 1
rlabel pdiffusion 106 84 107 85  0 t = 2
rlabel pdiffusion 103 89 104 90  0 t = 3
rlabel pdiffusion 106 89 107 90  0 t = 4
rlabel pdiffusion 102 84 108 90 0 cell no = 2
<< m1 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2c >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 3
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 4
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 5
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 85 12 86 13  0 t = 1
rlabel pdiffusion 88 12 89 13  0 t = 2
rlabel pdiffusion 85 17 86 18  0 t = 3
rlabel pdiffusion 88 17 89 18  0 t = 4
rlabel pdiffusion 84 12 90 18 0 cell no = 6
<< m1 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2 >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< m2c >>
rect 85 12 86 13 
rect 88 12 89 13 
rect 85 17 86 18 
rect 88 17 89 18 
<< labels >>
rlabel pdiffusion 121 84 122 85  0 t = 1
rlabel pdiffusion 124 84 125 85  0 t = 2
rlabel pdiffusion 121 89 122 90  0 t = 3
rlabel pdiffusion 124 89 125 90  0 t = 4
rlabel pdiffusion 120 84 126 90 0 cell no = 7
<< m1 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2c >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 8
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 9
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 10
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 11
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 12
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 13
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 14
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 15
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 16
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 17
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 67 30 68 31  0 t = 1
rlabel pdiffusion 70 30 71 31  0 t = 2
rlabel pdiffusion 67 35 68 36  0 t = 3
rlabel pdiffusion 70 35 71 36  0 t = 4
rlabel pdiffusion 66 30 72 36 0 cell no = 18
<< m1 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2c >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 19
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 20
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 21
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 13 120 14 121  0 t = 1
rlabel pdiffusion 16 120 17 121  0 t = 2
rlabel pdiffusion 13 125 14 126  0 t = 3
rlabel pdiffusion 16 125 17 126  0 t = 4
rlabel pdiffusion 12 120 18 126 0 cell no = 22
<< m1 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2c >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 23
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 24
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 25
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 26
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 27
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 121 102 122 103  0 t = 1
rlabel pdiffusion 124 102 125 103  0 t = 2
rlabel pdiffusion 121 107 122 108  0 t = 3
rlabel pdiffusion 124 107 125 108  0 t = 4
rlabel pdiffusion 120 102 126 108 0 cell no = 28
<< m1 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2 >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< m2c >>
rect 121 102 122 103 
rect 124 102 125 103 
rect 121 107 122 108 
rect 124 107 125 108 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 29
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 31 84 32 85  0 t = 1
rlabel pdiffusion 34 84 35 85  0 t = 2
rlabel pdiffusion 31 89 32 90  0 t = 3
rlabel pdiffusion 34 89 35 90  0 t = 4
rlabel pdiffusion 30 84 36 90 0 cell no = 30
<< m1 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2c >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 31
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 32
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 33
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 34
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 67 120 68 121  0 t = 1
rlabel pdiffusion 70 120 71 121  0 t = 2
rlabel pdiffusion 67 125 68 126  0 t = 3
rlabel pdiffusion 70 125 71 126  0 t = 4
rlabel pdiffusion 66 120 72 126 0 cell no = 35
<< m1 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2c >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 36
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 37
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 38
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 103 120 104 121  0 t = 1
rlabel pdiffusion 106 120 107 121  0 t = 2
rlabel pdiffusion 103 125 104 126  0 t = 3
rlabel pdiffusion 106 125 107 126  0 t = 4
rlabel pdiffusion 102 120 108 126 0 cell no = 39
<< m1 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2c >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 40
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 41
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 31 12 32 13  0 t = 1
rlabel pdiffusion 34 12 35 13  0 t = 2
rlabel pdiffusion 31 17 32 18  0 t = 3
rlabel pdiffusion 34 17 35 18  0 t = 4
rlabel pdiffusion 30 12 36 18 0 cell no = 42
<< m1 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2c >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 43
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 44
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 45
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< end >> 
