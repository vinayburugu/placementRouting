magic
tech scmos
timestamp 11111111111
<< m1 >>
rect 142 10 143 11 
<< m1 >>
rect 143 10 144 11 
<< m1 >>
rect 144 10 145 11 
<< m1 >>
rect 145 10 146 11 
<< m1 >>
rect 280 10 281 11 
<< m1 >>
rect 281 10 282 11 
<< m1 >>
rect 282 10 283 11 
<< m1 >>
rect 283 10 284 11 
<< m1 >>
rect 289 10 290 11 
<< m1 >>
rect 290 10 291 11 
<< m1 >>
rect 291 10 292 11 
<< m1 >>
rect 292 10 293 11 
<< m1 >>
rect 293 10 294 11 
<< m1 >>
rect 294 10 295 11 
<< m1 >>
rect 295 10 296 11 
<< m1 >>
rect 296 10 297 11 
<< m1 >>
rect 297 10 298 11 
<< m1 >>
rect 298 10 299 11 
<< m1 >>
rect 299 10 300 11 
<< m1 >>
rect 300 10 301 11 
<< m1 >>
rect 301 10 302 11 
<< m1 >>
rect 505 10 506 11 
<< m1 >>
rect 506 10 507 11 
<< m1 >>
rect 507 10 508 11 
<< m1 >>
rect 508 10 509 11 
<< m1 >>
rect 509 10 510 11 
<< m1 >>
rect 510 10 511 11 
<< m1 >>
rect 511 10 512 11 
<< m1 >>
rect 512 10 513 11 
<< m1 >>
rect 513 10 514 11 
<< m1 >>
rect 514 10 515 11 
<< m1 >>
rect 515 10 516 11 
<< m1 >>
rect 516 10 517 11 
<< m1 >>
rect 517 10 518 11 
<< m1 >>
rect 142 11 143 12 
<< m1 >>
rect 145 11 146 12 
<< m1 >>
rect 280 11 281 12 
<< m1 >>
rect 283 11 284 12 
<< m1 >>
rect 289 11 290 12 
<< m1 >>
rect 301 11 302 12 
<< m1 >>
rect 505 11 506 12 
<< m1 >>
rect 517 11 518 12 
<< pdiffusion >>
rect 12 12 13 13 
<< pdiffusion >>
rect 13 12 14 13 
<< pdiffusion >>
rect 14 12 15 13 
<< pdiffusion >>
rect 15 12 16 13 
<< pdiffusion >>
rect 16 12 17 13 
<< pdiffusion >>
rect 17 12 18 13 
<< pdiffusion >>
rect 30 12 31 13 
<< pdiffusion >>
rect 31 12 32 13 
<< pdiffusion >>
rect 32 12 33 13 
<< pdiffusion >>
rect 33 12 34 13 
<< pdiffusion >>
rect 34 12 35 13 
<< pdiffusion >>
rect 35 12 36 13 
<< pdiffusion >>
rect 48 12 49 13 
<< pdiffusion >>
rect 49 12 50 13 
<< pdiffusion >>
rect 50 12 51 13 
<< pdiffusion >>
rect 51 12 52 13 
<< pdiffusion >>
rect 52 12 53 13 
<< pdiffusion >>
rect 53 12 54 13 
<< pdiffusion >>
rect 66 12 67 13 
<< pdiffusion >>
rect 67 12 68 13 
<< pdiffusion >>
rect 68 12 69 13 
<< pdiffusion >>
rect 69 12 70 13 
<< pdiffusion >>
rect 70 12 71 13 
<< pdiffusion >>
rect 71 12 72 13 
<< pdiffusion >>
rect 102 12 103 13 
<< pdiffusion >>
rect 103 12 104 13 
<< pdiffusion >>
rect 104 12 105 13 
<< pdiffusion >>
rect 105 12 106 13 
<< pdiffusion >>
rect 106 12 107 13 
<< pdiffusion >>
rect 107 12 108 13 
<< pdiffusion >>
rect 120 12 121 13 
<< pdiffusion >>
rect 121 12 122 13 
<< pdiffusion >>
rect 122 12 123 13 
<< pdiffusion >>
rect 123 12 124 13 
<< pdiffusion >>
rect 124 12 125 13 
<< pdiffusion >>
rect 125 12 126 13 
<< pdiffusion >>
rect 138 12 139 13 
<< pdiffusion >>
rect 139 12 140 13 
<< pdiffusion >>
rect 140 12 141 13 
<< pdiffusion >>
rect 141 12 142 13 
<< m1 >>
rect 142 12 143 13 
<< pdiffusion >>
rect 142 12 143 13 
<< pdiffusion >>
rect 143 12 144 13 
<< m1 >>
rect 145 12 146 13 
<< pdiffusion >>
rect 156 12 157 13 
<< pdiffusion >>
rect 157 12 158 13 
<< pdiffusion >>
rect 158 12 159 13 
<< pdiffusion >>
rect 159 12 160 13 
<< pdiffusion >>
rect 160 12 161 13 
<< pdiffusion >>
rect 161 12 162 13 
<< pdiffusion >>
rect 174 12 175 13 
<< pdiffusion >>
rect 175 12 176 13 
<< pdiffusion >>
rect 176 12 177 13 
<< pdiffusion >>
rect 177 12 178 13 
<< pdiffusion >>
rect 178 12 179 13 
<< pdiffusion >>
rect 179 12 180 13 
<< pdiffusion >>
rect 192 12 193 13 
<< pdiffusion >>
rect 193 12 194 13 
<< pdiffusion >>
rect 194 12 195 13 
<< pdiffusion >>
rect 195 12 196 13 
<< pdiffusion >>
rect 196 12 197 13 
<< pdiffusion >>
rect 197 12 198 13 
<< pdiffusion >>
rect 210 12 211 13 
<< pdiffusion >>
rect 211 12 212 13 
<< pdiffusion >>
rect 212 12 213 13 
<< pdiffusion >>
rect 213 12 214 13 
<< pdiffusion >>
rect 214 12 215 13 
<< pdiffusion >>
rect 215 12 216 13 
<< pdiffusion >>
rect 228 12 229 13 
<< pdiffusion >>
rect 229 12 230 13 
<< pdiffusion >>
rect 230 12 231 13 
<< pdiffusion >>
rect 231 12 232 13 
<< pdiffusion >>
rect 232 12 233 13 
<< pdiffusion >>
rect 233 12 234 13 
<< pdiffusion >>
rect 246 12 247 13 
<< pdiffusion >>
rect 247 12 248 13 
<< pdiffusion >>
rect 248 12 249 13 
<< pdiffusion >>
rect 249 12 250 13 
<< pdiffusion >>
rect 250 12 251 13 
<< pdiffusion >>
rect 251 12 252 13 
<< pdiffusion >>
rect 264 12 265 13 
<< pdiffusion >>
rect 265 12 266 13 
<< pdiffusion >>
rect 266 12 267 13 
<< pdiffusion >>
rect 267 12 268 13 
<< pdiffusion >>
rect 268 12 269 13 
<< pdiffusion >>
rect 269 12 270 13 
<< m1 >>
rect 280 12 281 13 
<< pdiffusion >>
rect 282 12 283 13 
<< m1 >>
rect 283 12 284 13 
<< pdiffusion >>
rect 283 12 284 13 
<< pdiffusion >>
rect 284 12 285 13 
<< pdiffusion >>
rect 285 12 286 13 
<< pdiffusion >>
rect 286 12 287 13 
<< pdiffusion >>
rect 287 12 288 13 
<< m1 >>
rect 289 12 290 13 
<< pdiffusion >>
rect 300 12 301 13 
<< m1 >>
rect 301 12 302 13 
<< pdiffusion >>
rect 301 12 302 13 
<< pdiffusion >>
rect 302 12 303 13 
<< pdiffusion >>
rect 303 12 304 13 
<< pdiffusion >>
rect 304 12 305 13 
<< pdiffusion >>
rect 305 12 306 13 
<< pdiffusion >>
rect 318 12 319 13 
<< pdiffusion >>
rect 319 12 320 13 
<< pdiffusion >>
rect 320 12 321 13 
<< pdiffusion >>
rect 321 12 322 13 
<< pdiffusion >>
rect 322 12 323 13 
<< pdiffusion >>
rect 323 12 324 13 
<< pdiffusion >>
rect 336 12 337 13 
<< pdiffusion >>
rect 337 12 338 13 
<< pdiffusion >>
rect 338 12 339 13 
<< pdiffusion >>
rect 339 12 340 13 
<< pdiffusion >>
rect 340 12 341 13 
<< pdiffusion >>
rect 341 12 342 13 
<< pdiffusion >>
rect 354 12 355 13 
<< pdiffusion >>
rect 355 12 356 13 
<< pdiffusion >>
rect 356 12 357 13 
<< pdiffusion >>
rect 357 12 358 13 
<< pdiffusion >>
rect 358 12 359 13 
<< pdiffusion >>
rect 359 12 360 13 
<< pdiffusion >>
rect 372 12 373 13 
<< pdiffusion >>
rect 373 12 374 13 
<< pdiffusion >>
rect 374 12 375 13 
<< pdiffusion >>
rect 375 12 376 13 
<< pdiffusion >>
rect 376 12 377 13 
<< pdiffusion >>
rect 377 12 378 13 
<< pdiffusion >>
rect 390 12 391 13 
<< pdiffusion >>
rect 391 12 392 13 
<< pdiffusion >>
rect 392 12 393 13 
<< pdiffusion >>
rect 393 12 394 13 
<< pdiffusion >>
rect 394 12 395 13 
<< pdiffusion >>
rect 395 12 396 13 
<< pdiffusion >>
rect 408 12 409 13 
<< pdiffusion >>
rect 409 12 410 13 
<< pdiffusion >>
rect 410 12 411 13 
<< pdiffusion >>
rect 411 12 412 13 
<< pdiffusion >>
rect 412 12 413 13 
<< pdiffusion >>
rect 413 12 414 13 
<< pdiffusion >>
rect 426 12 427 13 
<< pdiffusion >>
rect 427 12 428 13 
<< pdiffusion >>
rect 428 12 429 13 
<< pdiffusion >>
rect 429 12 430 13 
<< pdiffusion >>
rect 430 12 431 13 
<< pdiffusion >>
rect 431 12 432 13 
<< pdiffusion >>
rect 444 12 445 13 
<< pdiffusion >>
rect 445 12 446 13 
<< pdiffusion >>
rect 446 12 447 13 
<< pdiffusion >>
rect 447 12 448 13 
<< pdiffusion >>
rect 448 12 449 13 
<< pdiffusion >>
rect 449 12 450 13 
<< pdiffusion >>
rect 462 12 463 13 
<< pdiffusion >>
rect 463 12 464 13 
<< pdiffusion >>
rect 464 12 465 13 
<< pdiffusion >>
rect 465 12 466 13 
<< pdiffusion >>
rect 466 12 467 13 
<< pdiffusion >>
rect 467 12 468 13 
<< pdiffusion >>
rect 480 12 481 13 
<< pdiffusion >>
rect 481 12 482 13 
<< pdiffusion >>
rect 482 12 483 13 
<< pdiffusion >>
rect 483 12 484 13 
<< pdiffusion >>
rect 484 12 485 13 
<< pdiffusion >>
rect 485 12 486 13 
<< pdiffusion >>
rect 498 12 499 13 
<< pdiffusion >>
rect 499 12 500 13 
<< pdiffusion >>
rect 500 12 501 13 
<< pdiffusion >>
rect 501 12 502 13 
<< pdiffusion >>
rect 502 12 503 13 
<< pdiffusion >>
rect 503 12 504 13 
<< m1 >>
rect 505 12 506 13 
<< pdiffusion >>
rect 516 12 517 13 
<< m1 >>
rect 517 12 518 13 
<< pdiffusion >>
rect 517 12 518 13 
<< pdiffusion >>
rect 518 12 519 13 
<< pdiffusion >>
rect 519 12 520 13 
<< pdiffusion >>
rect 520 12 521 13 
<< pdiffusion >>
rect 521 12 522 13 
<< pdiffusion >>
rect 12 13 13 14 
<< pdiffusion >>
rect 13 13 14 14 
<< pdiffusion >>
rect 14 13 15 14 
<< pdiffusion >>
rect 15 13 16 14 
<< pdiffusion >>
rect 16 13 17 14 
<< pdiffusion >>
rect 17 13 18 14 
<< pdiffusion >>
rect 30 13 31 14 
<< pdiffusion >>
rect 31 13 32 14 
<< pdiffusion >>
rect 32 13 33 14 
<< pdiffusion >>
rect 33 13 34 14 
<< pdiffusion >>
rect 34 13 35 14 
<< pdiffusion >>
rect 35 13 36 14 
<< pdiffusion >>
rect 48 13 49 14 
<< pdiffusion >>
rect 49 13 50 14 
<< pdiffusion >>
rect 50 13 51 14 
<< pdiffusion >>
rect 51 13 52 14 
<< pdiffusion >>
rect 52 13 53 14 
<< pdiffusion >>
rect 53 13 54 14 
<< pdiffusion >>
rect 66 13 67 14 
<< pdiffusion >>
rect 67 13 68 14 
<< pdiffusion >>
rect 68 13 69 14 
<< pdiffusion >>
rect 69 13 70 14 
<< pdiffusion >>
rect 70 13 71 14 
<< pdiffusion >>
rect 71 13 72 14 
<< pdiffusion >>
rect 102 13 103 14 
<< pdiffusion >>
rect 103 13 104 14 
<< pdiffusion >>
rect 104 13 105 14 
<< pdiffusion >>
rect 105 13 106 14 
<< pdiffusion >>
rect 106 13 107 14 
<< pdiffusion >>
rect 107 13 108 14 
<< pdiffusion >>
rect 120 13 121 14 
<< pdiffusion >>
rect 121 13 122 14 
<< pdiffusion >>
rect 122 13 123 14 
<< pdiffusion >>
rect 123 13 124 14 
<< pdiffusion >>
rect 124 13 125 14 
<< pdiffusion >>
rect 125 13 126 14 
<< pdiffusion >>
rect 138 13 139 14 
<< pdiffusion >>
rect 139 13 140 14 
<< pdiffusion >>
rect 140 13 141 14 
<< pdiffusion >>
rect 141 13 142 14 
<< pdiffusion >>
rect 142 13 143 14 
<< pdiffusion >>
rect 143 13 144 14 
<< m1 >>
rect 145 13 146 14 
<< pdiffusion >>
rect 156 13 157 14 
<< pdiffusion >>
rect 157 13 158 14 
<< pdiffusion >>
rect 158 13 159 14 
<< pdiffusion >>
rect 159 13 160 14 
<< pdiffusion >>
rect 160 13 161 14 
<< pdiffusion >>
rect 161 13 162 14 
<< pdiffusion >>
rect 174 13 175 14 
<< pdiffusion >>
rect 175 13 176 14 
<< pdiffusion >>
rect 176 13 177 14 
<< pdiffusion >>
rect 177 13 178 14 
<< pdiffusion >>
rect 178 13 179 14 
<< pdiffusion >>
rect 179 13 180 14 
<< pdiffusion >>
rect 192 13 193 14 
<< pdiffusion >>
rect 193 13 194 14 
<< pdiffusion >>
rect 194 13 195 14 
<< pdiffusion >>
rect 195 13 196 14 
<< pdiffusion >>
rect 196 13 197 14 
<< pdiffusion >>
rect 197 13 198 14 
<< pdiffusion >>
rect 210 13 211 14 
<< pdiffusion >>
rect 211 13 212 14 
<< pdiffusion >>
rect 212 13 213 14 
<< pdiffusion >>
rect 213 13 214 14 
<< pdiffusion >>
rect 214 13 215 14 
<< pdiffusion >>
rect 215 13 216 14 
<< pdiffusion >>
rect 228 13 229 14 
<< pdiffusion >>
rect 229 13 230 14 
<< pdiffusion >>
rect 230 13 231 14 
<< pdiffusion >>
rect 231 13 232 14 
<< pdiffusion >>
rect 232 13 233 14 
<< pdiffusion >>
rect 233 13 234 14 
<< pdiffusion >>
rect 246 13 247 14 
<< pdiffusion >>
rect 247 13 248 14 
<< pdiffusion >>
rect 248 13 249 14 
<< pdiffusion >>
rect 249 13 250 14 
<< pdiffusion >>
rect 250 13 251 14 
<< pdiffusion >>
rect 251 13 252 14 
<< pdiffusion >>
rect 264 13 265 14 
<< pdiffusion >>
rect 265 13 266 14 
<< pdiffusion >>
rect 266 13 267 14 
<< pdiffusion >>
rect 267 13 268 14 
<< pdiffusion >>
rect 268 13 269 14 
<< pdiffusion >>
rect 269 13 270 14 
<< m1 >>
rect 280 13 281 14 
<< pdiffusion >>
rect 282 13 283 14 
<< pdiffusion >>
rect 283 13 284 14 
<< pdiffusion >>
rect 284 13 285 14 
<< pdiffusion >>
rect 285 13 286 14 
<< pdiffusion >>
rect 286 13 287 14 
<< pdiffusion >>
rect 287 13 288 14 
<< m1 >>
rect 289 13 290 14 
<< pdiffusion >>
rect 300 13 301 14 
<< pdiffusion >>
rect 301 13 302 14 
<< pdiffusion >>
rect 302 13 303 14 
<< pdiffusion >>
rect 303 13 304 14 
<< pdiffusion >>
rect 304 13 305 14 
<< pdiffusion >>
rect 305 13 306 14 
<< pdiffusion >>
rect 318 13 319 14 
<< pdiffusion >>
rect 319 13 320 14 
<< pdiffusion >>
rect 320 13 321 14 
<< pdiffusion >>
rect 321 13 322 14 
<< pdiffusion >>
rect 322 13 323 14 
<< pdiffusion >>
rect 323 13 324 14 
<< pdiffusion >>
rect 336 13 337 14 
<< pdiffusion >>
rect 337 13 338 14 
<< pdiffusion >>
rect 338 13 339 14 
<< pdiffusion >>
rect 339 13 340 14 
<< pdiffusion >>
rect 340 13 341 14 
<< pdiffusion >>
rect 341 13 342 14 
<< pdiffusion >>
rect 354 13 355 14 
<< pdiffusion >>
rect 355 13 356 14 
<< pdiffusion >>
rect 356 13 357 14 
<< pdiffusion >>
rect 357 13 358 14 
<< pdiffusion >>
rect 358 13 359 14 
<< pdiffusion >>
rect 359 13 360 14 
<< pdiffusion >>
rect 372 13 373 14 
<< pdiffusion >>
rect 373 13 374 14 
<< pdiffusion >>
rect 374 13 375 14 
<< pdiffusion >>
rect 375 13 376 14 
<< pdiffusion >>
rect 376 13 377 14 
<< pdiffusion >>
rect 377 13 378 14 
<< pdiffusion >>
rect 390 13 391 14 
<< pdiffusion >>
rect 391 13 392 14 
<< pdiffusion >>
rect 392 13 393 14 
<< pdiffusion >>
rect 393 13 394 14 
<< pdiffusion >>
rect 394 13 395 14 
<< pdiffusion >>
rect 395 13 396 14 
<< pdiffusion >>
rect 408 13 409 14 
<< pdiffusion >>
rect 409 13 410 14 
<< pdiffusion >>
rect 410 13 411 14 
<< pdiffusion >>
rect 411 13 412 14 
<< pdiffusion >>
rect 412 13 413 14 
<< pdiffusion >>
rect 413 13 414 14 
<< pdiffusion >>
rect 426 13 427 14 
<< pdiffusion >>
rect 427 13 428 14 
<< pdiffusion >>
rect 428 13 429 14 
<< pdiffusion >>
rect 429 13 430 14 
<< pdiffusion >>
rect 430 13 431 14 
<< pdiffusion >>
rect 431 13 432 14 
<< pdiffusion >>
rect 444 13 445 14 
<< pdiffusion >>
rect 445 13 446 14 
<< pdiffusion >>
rect 446 13 447 14 
<< pdiffusion >>
rect 447 13 448 14 
<< pdiffusion >>
rect 448 13 449 14 
<< pdiffusion >>
rect 449 13 450 14 
<< pdiffusion >>
rect 462 13 463 14 
<< pdiffusion >>
rect 463 13 464 14 
<< pdiffusion >>
rect 464 13 465 14 
<< pdiffusion >>
rect 465 13 466 14 
<< pdiffusion >>
rect 466 13 467 14 
<< pdiffusion >>
rect 467 13 468 14 
<< pdiffusion >>
rect 480 13 481 14 
<< pdiffusion >>
rect 481 13 482 14 
<< pdiffusion >>
rect 482 13 483 14 
<< pdiffusion >>
rect 483 13 484 14 
<< pdiffusion >>
rect 484 13 485 14 
<< pdiffusion >>
rect 485 13 486 14 
<< pdiffusion >>
rect 498 13 499 14 
<< pdiffusion >>
rect 499 13 500 14 
<< pdiffusion >>
rect 500 13 501 14 
<< pdiffusion >>
rect 501 13 502 14 
<< pdiffusion >>
rect 502 13 503 14 
<< pdiffusion >>
rect 503 13 504 14 
<< m1 >>
rect 505 13 506 14 
<< pdiffusion >>
rect 516 13 517 14 
<< pdiffusion >>
rect 517 13 518 14 
<< pdiffusion >>
rect 518 13 519 14 
<< pdiffusion >>
rect 519 13 520 14 
<< pdiffusion >>
rect 520 13 521 14 
<< pdiffusion >>
rect 521 13 522 14 
<< pdiffusion >>
rect 12 14 13 15 
<< pdiffusion >>
rect 13 14 14 15 
<< pdiffusion >>
rect 14 14 15 15 
<< pdiffusion >>
rect 15 14 16 15 
<< pdiffusion >>
rect 16 14 17 15 
<< pdiffusion >>
rect 17 14 18 15 
<< pdiffusion >>
rect 30 14 31 15 
<< pdiffusion >>
rect 31 14 32 15 
<< pdiffusion >>
rect 32 14 33 15 
<< pdiffusion >>
rect 33 14 34 15 
<< pdiffusion >>
rect 34 14 35 15 
<< pdiffusion >>
rect 35 14 36 15 
<< pdiffusion >>
rect 48 14 49 15 
<< pdiffusion >>
rect 49 14 50 15 
<< pdiffusion >>
rect 50 14 51 15 
<< pdiffusion >>
rect 51 14 52 15 
<< pdiffusion >>
rect 52 14 53 15 
<< pdiffusion >>
rect 53 14 54 15 
<< pdiffusion >>
rect 66 14 67 15 
<< pdiffusion >>
rect 67 14 68 15 
<< pdiffusion >>
rect 68 14 69 15 
<< pdiffusion >>
rect 69 14 70 15 
<< pdiffusion >>
rect 70 14 71 15 
<< pdiffusion >>
rect 71 14 72 15 
<< pdiffusion >>
rect 102 14 103 15 
<< pdiffusion >>
rect 103 14 104 15 
<< pdiffusion >>
rect 104 14 105 15 
<< pdiffusion >>
rect 105 14 106 15 
<< pdiffusion >>
rect 106 14 107 15 
<< pdiffusion >>
rect 107 14 108 15 
<< pdiffusion >>
rect 120 14 121 15 
<< pdiffusion >>
rect 121 14 122 15 
<< pdiffusion >>
rect 122 14 123 15 
<< pdiffusion >>
rect 123 14 124 15 
<< pdiffusion >>
rect 124 14 125 15 
<< pdiffusion >>
rect 125 14 126 15 
<< pdiffusion >>
rect 138 14 139 15 
<< pdiffusion >>
rect 139 14 140 15 
<< pdiffusion >>
rect 140 14 141 15 
<< pdiffusion >>
rect 141 14 142 15 
<< pdiffusion >>
rect 142 14 143 15 
<< pdiffusion >>
rect 143 14 144 15 
<< m1 >>
rect 145 14 146 15 
<< pdiffusion >>
rect 156 14 157 15 
<< pdiffusion >>
rect 157 14 158 15 
<< pdiffusion >>
rect 158 14 159 15 
<< pdiffusion >>
rect 159 14 160 15 
<< pdiffusion >>
rect 160 14 161 15 
<< pdiffusion >>
rect 161 14 162 15 
<< pdiffusion >>
rect 174 14 175 15 
<< pdiffusion >>
rect 175 14 176 15 
<< pdiffusion >>
rect 176 14 177 15 
<< pdiffusion >>
rect 177 14 178 15 
<< pdiffusion >>
rect 178 14 179 15 
<< pdiffusion >>
rect 179 14 180 15 
<< pdiffusion >>
rect 192 14 193 15 
<< pdiffusion >>
rect 193 14 194 15 
<< pdiffusion >>
rect 194 14 195 15 
<< pdiffusion >>
rect 195 14 196 15 
<< pdiffusion >>
rect 196 14 197 15 
<< pdiffusion >>
rect 197 14 198 15 
<< pdiffusion >>
rect 210 14 211 15 
<< pdiffusion >>
rect 211 14 212 15 
<< pdiffusion >>
rect 212 14 213 15 
<< pdiffusion >>
rect 213 14 214 15 
<< pdiffusion >>
rect 214 14 215 15 
<< pdiffusion >>
rect 215 14 216 15 
<< pdiffusion >>
rect 228 14 229 15 
<< pdiffusion >>
rect 229 14 230 15 
<< pdiffusion >>
rect 230 14 231 15 
<< pdiffusion >>
rect 231 14 232 15 
<< pdiffusion >>
rect 232 14 233 15 
<< pdiffusion >>
rect 233 14 234 15 
<< pdiffusion >>
rect 246 14 247 15 
<< pdiffusion >>
rect 247 14 248 15 
<< pdiffusion >>
rect 248 14 249 15 
<< pdiffusion >>
rect 249 14 250 15 
<< pdiffusion >>
rect 250 14 251 15 
<< pdiffusion >>
rect 251 14 252 15 
<< pdiffusion >>
rect 264 14 265 15 
<< pdiffusion >>
rect 265 14 266 15 
<< pdiffusion >>
rect 266 14 267 15 
<< pdiffusion >>
rect 267 14 268 15 
<< pdiffusion >>
rect 268 14 269 15 
<< pdiffusion >>
rect 269 14 270 15 
<< m1 >>
rect 280 14 281 15 
<< pdiffusion >>
rect 282 14 283 15 
<< pdiffusion >>
rect 283 14 284 15 
<< pdiffusion >>
rect 284 14 285 15 
<< pdiffusion >>
rect 285 14 286 15 
<< pdiffusion >>
rect 286 14 287 15 
<< pdiffusion >>
rect 287 14 288 15 
<< m1 >>
rect 289 14 290 15 
<< pdiffusion >>
rect 300 14 301 15 
<< pdiffusion >>
rect 301 14 302 15 
<< pdiffusion >>
rect 302 14 303 15 
<< pdiffusion >>
rect 303 14 304 15 
<< pdiffusion >>
rect 304 14 305 15 
<< pdiffusion >>
rect 305 14 306 15 
<< pdiffusion >>
rect 318 14 319 15 
<< pdiffusion >>
rect 319 14 320 15 
<< pdiffusion >>
rect 320 14 321 15 
<< pdiffusion >>
rect 321 14 322 15 
<< pdiffusion >>
rect 322 14 323 15 
<< pdiffusion >>
rect 323 14 324 15 
<< pdiffusion >>
rect 336 14 337 15 
<< pdiffusion >>
rect 337 14 338 15 
<< pdiffusion >>
rect 338 14 339 15 
<< pdiffusion >>
rect 339 14 340 15 
<< pdiffusion >>
rect 340 14 341 15 
<< pdiffusion >>
rect 341 14 342 15 
<< pdiffusion >>
rect 354 14 355 15 
<< pdiffusion >>
rect 355 14 356 15 
<< pdiffusion >>
rect 356 14 357 15 
<< pdiffusion >>
rect 357 14 358 15 
<< pdiffusion >>
rect 358 14 359 15 
<< pdiffusion >>
rect 359 14 360 15 
<< pdiffusion >>
rect 372 14 373 15 
<< pdiffusion >>
rect 373 14 374 15 
<< pdiffusion >>
rect 374 14 375 15 
<< pdiffusion >>
rect 375 14 376 15 
<< pdiffusion >>
rect 376 14 377 15 
<< pdiffusion >>
rect 377 14 378 15 
<< pdiffusion >>
rect 390 14 391 15 
<< pdiffusion >>
rect 391 14 392 15 
<< pdiffusion >>
rect 392 14 393 15 
<< pdiffusion >>
rect 393 14 394 15 
<< pdiffusion >>
rect 394 14 395 15 
<< pdiffusion >>
rect 395 14 396 15 
<< pdiffusion >>
rect 408 14 409 15 
<< pdiffusion >>
rect 409 14 410 15 
<< pdiffusion >>
rect 410 14 411 15 
<< pdiffusion >>
rect 411 14 412 15 
<< pdiffusion >>
rect 412 14 413 15 
<< pdiffusion >>
rect 413 14 414 15 
<< pdiffusion >>
rect 426 14 427 15 
<< pdiffusion >>
rect 427 14 428 15 
<< pdiffusion >>
rect 428 14 429 15 
<< pdiffusion >>
rect 429 14 430 15 
<< pdiffusion >>
rect 430 14 431 15 
<< pdiffusion >>
rect 431 14 432 15 
<< pdiffusion >>
rect 444 14 445 15 
<< pdiffusion >>
rect 445 14 446 15 
<< pdiffusion >>
rect 446 14 447 15 
<< pdiffusion >>
rect 447 14 448 15 
<< pdiffusion >>
rect 448 14 449 15 
<< pdiffusion >>
rect 449 14 450 15 
<< pdiffusion >>
rect 462 14 463 15 
<< pdiffusion >>
rect 463 14 464 15 
<< pdiffusion >>
rect 464 14 465 15 
<< pdiffusion >>
rect 465 14 466 15 
<< pdiffusion >>
rect 466 14 467 15 
<< pdiffusion >>
rect 467 14 468 15 
<< pdiffusion >>
rect 480 14 481 15 
<< pdiffusion >>
rect 481 14 482 15 
<< pdiffusion >>
rect 482 14 483 15 
<< pdiffusion >>
rect 483 14 484 15 
<< pdiffusion >>
rect 484 14 485 15 
<< pdiffusion >>
rect 485 14 486 15 
<< pdiffusion >>
rect 498 14 499 15 
<< pdiffusion >>
rect 499 14 500 15 
<< pdiffusion >>
rect 500 14 501 15 
<< pdiffusion >>
rect 501 14 502 15 
<< pdiffusion >>
rect 502 14 503 15 
<< pdiffusion >>
rect 503 14 504 15 
<< m1 >>
rect 505 14 506 15 
<< pdiffusion >>
rect 516 14 517 15 
<< pdiffusion >>
rect 517 14 518 15 
<< pdiffusion >>
rect 518 14 519 15 
<< pdiffusion >>
rect 519 14 520 15 
<< pdiffusion >>
rect 520 14 521 15 
<< pdiffusion >>
rect 521 14 522 15 
<< pdiffusion >>
rect 12 15 13 16 
<< pdiffusion >>
rect 13 15 14 16 
<< pdiffusion >>
rect 14 15 15 16 
<< pdiffusion >>
rect 15 15 16 16 
<< pdiffusion >>
rect 16 15 17 16 
<< pdiffusion >>
rect 17 15 18 16 
<< pdiffusion >>
rect 30 15 31 16 
<< pdiffusion >>
rect 31 15 32 16 
<< pdiffusion >>
rect 32 15 33 16 
<< pdiffusion >>
rect 33 15 34 16 
<< pdiffusion >>
rect 34 15 35 16 
<< pdiffusion >>
rect 35 15 36 16 
<< pdiffusion >>
rect 48 15 49 16 
<< pdiffusion >>
rect 49 15 50 16 
<< pdiffusion >>
rect 50 15 51 16 
<< pdiffusion >>
rect 51 15 52 16 
<< pdiffusion >>
rect 52 15 53 16 
<< pdiffusion >>
rect 53 15 54 16 
<< pdiffusion >>
rect 66 15 67 16 
<< pdiffusion >>
rect 67 15 68 16 
<< pdiffusion >>
rect 68 15 69 16 
<< pdiffusion >>
rect 69 15 70 16 
<< pdiffusion >>
rect 70 15 71 16 
<< pdiffusion >>
rect 71 15 72 16 
<< pdiffusion >>
rect 102 15 103 16 
<< pdiffusion >>
rect 103 15 104 16 
<< pdiffusion >>
rect 104 15 105 16 
<< pdiffusion >>
rect 105 15 106 16 
<< pdiffusion >>
rect 106 15 107 16 
<< pdiffusion >>
rect 107 15 108 16 
<< pdiffusion >>
rect 120 15 121 16 
<< pdiffusion >>
rect 121 15 122 16 
<< pdiffusion >>
rect 122 15 123 16 
<< pdiffusion >>
rect 123 15 124 16 
<< pdiffusion >>
rect 124 15 125 16 
<< pdiffusion >>
rect 125 15 126 16 
<< pdiffusion >>
rect 138 15 139 16 
<< pdiffusion >>
rect 139 15 140 16 
<< pdiffusion >>
rect 140 15 141 16 
<< pdiffusion >>
rect 141 15 142 16 
<< pdiffusion >>
rect 142 15 143 16 
<< pdiffusion >>
rect 143 15 144 16 
<< m1 >>
rect 145 15 146 16 
<< pdiffusion >>
rect 156 15 157 16 
<< pdiffusion >>
rect 157 15 158 16 
<< pdiffusion >>
rect 158 15 159 16 
<< pdiffusion >>
rect 159 15 160 16 
<< pdiffusion >>
rect 160 15 161 16 
<< pdiffusion >>
rect 161 15 162 16 
<< pdiffusion >>
rect 174 15 175 16 
<< pdiffusion >>
rect 175 15 176 16 
<< pdiffusion >>
rect 176 15 177 16 
<< pdiffusion >>
rect 177 15 178 16 
<< pdiffusion >>
rect 178 15 179 16 
<< pdiffusion >>
rect 179 15 180 16 
<< pdiffusion >>
rect 192 15 193 16 
<< pdiffusion >>
rect 193 15 194 16 
<< pdiffusion >>
rect 194 15 195 16 
<< pdiffusion >>
rect 195 15 196 16 
<< pdiffusion >>
rect 196 15 197 16 
<< pdiffusion >>
rect 197 15 198 16 
<< pdiffusion >>
rect 210 15 211 16 
<< pdiffusion >>
rect 211 15 212 16 
<< pdiffusion >>
rect 212 15 213 16 
<< pdiffusion >>
rect 213 15 214 16 
<< pdiffusion >>
rect 214 15 215 16 
<< pdiffusion >>
rect 215 15 216 16 
<< pdiffusion >>
rect 228 15 229 16 
<< pdiffusion >>
rect 229 15 230 16 
<< pdiffusion >>
rect 230 15 231 16 
<< pdiffusion >>
rect 231 15 232 16 
<< pdiffusion >>
rect 232 15 233 16 
<< pdiffusion >>
rect 233 15 234 16 
<< pdiffusion >>
rect 246 15 247 16 
<< pdiffusion >>
rect 247 15 248 16 
<< pdiffusion >>
rect 248 15 249 16 
<< pdiffusion >>
rect 249 15 250 16 
<< pdiffusion >>
rect 250 15 251 16 
<< pdiffusion >>
rect 251 15 252 16 
<< pdiffusion >>
rect 264 15 265 16 
<< pdiffusion >>
rect 265 15 266 16 
<< pdiffusion >>
rect 266 15 267 16 
<< pdiffusion >>
rect 267 15 268 16 
<< pdiffusion >>
rect 268 15 269 16 
<< pdiffusion >>
rect 269 15 270 16 
<< m1 >>
rect 280 15 281 16 
<< pdiffusion >>
rect 282 15 283 16 
<< pdiffusion >>
rect 283 15 284 16 
<< pdiffusion >>
rect 284 15 285 16 
<< pdiffusion >>
rect 285 15 286 16 
<< pdiffusion >>
rect 286 15 287 16 
<< pdiffusion >>
rect 287 15 288 16 
<< m1 >>
rect 289 15 290 16 
<< pdiffusion >>
rect 300 15 301 16 
<< pdiffusion >>
rect 301 15 302 16 
<< pdiffusion >>
rect 302 15 303 16 
<< pdiffusion >>
rect 303 15 304 16 
<< pdiffusion >>
rect 304 15 305 16 
<< pdiffusion >>
rect 305 15 306 16 
<< pdiffusion >>
rect 318 15 319 16 
<< pdiffusion >>
rect 319 15 320 16 
<< pdiffusion >>
rect 320 15 321 16 
<< pdiffusion >>
rect 321 15 322 16 
<< pdiffusion >>
rect 322 15 323 16 
<< pdiffusion >>
rect 323 15 324 16 
<< pdiffusion >>
rect 336 15 337 16 
<< pdiffusion >>
rect 337 15 338 16 
<< pdiffusion >>
rect 338 15 339 16 
<< pdiffusion >>
rect 339 15 340 16 
<< pdiffusion >>
rect 340 15 341 16 
<< pdiffusion >>
rect 341 15 342 16 
<< pdiffusion >>
rect 354 15 355 16 
<< pdiffusion >>
rect 355 15 356 16 
<< pdiffusion >>
rect 356 15 357 16 
<< pdiffusion >>
rect 357 15 358 16 
<< pdiffusion >>
rect 358 15 359 16 
<< pdiffusion >>
rect 359 15 360 16 
<< pdiffusion >>
rect 372 15 373 16 
<< pdiffusion >>
rect 373 15 374 16 
<< pdiffusion >>
rect 374 15 375 16 
<< pdiffusion >>
rect 375 15 376 16 
<< pdiffusion >>
rect 376 15 377 16 
<< pdiffusion >>
rect 377 15 378 16 
<< pdiffusion >>
rect 390 15 391 16 
<< pdiffusion >>
rect 391 15 392 16 
<< pdiffusion >>
rect 392 15 393 16 
<< pdiffusion >>
rect 393 15 394 16 
<< pdiffusion >>
rect 394 15 395 16 
<< pdiffusion >>
rect 395 15 396 16 
<< pdiffusion >>
rect 408 15 409 16 
<< pdiffusion >>
rect 409 15 410 16 
<< pdiffusion >>
rect 410 15 411 16 
<< pdiffusion >>
rect 411 15 412 16 
<< pdiffusion >>
rect 412 15 413 16 
<< pdiffusion >>
rect 413 15 414 16 
<< pdiffusion >>
rect 426 15 427 16 
<< pdiffusion >>
rect 427 15 428 16 
<< pdiffusion >>
rect 428 15 429 16 
<< pdiffusion >>
rect 429 15 430 16 
<< pdiffusion >>
rect 430 15 431 16 
<< pdiffusion >>
rect 431 15 432 16 
<< pdiffusion >>
rect 444 15 445 16 
<< pdiffusion >>
rect 445 15 446 16 
<< pdiffusion >>
rect 446 15 447 16 
<< pdiffusion >>
rect 447 15 448 16 
<< pdiffusion >>
rect 448 15 449 16 
<< pdiffusion >>
rect 449 15 450 16 
<< pdiffusion >>
rect 462 15 463 16 
<< pdiffusion >>
rect 463 15 464 16 
<< pdiffusion >>
rect 464 15 465 16 
<< pdiffusion >>
rect 465 15 466 16 
<< pdiffusion >>
rect 466 15 467 16 
<< pdiffusion >>
rect 467 15 468 16 
<< pdiffusion >>
rect 480 15 481 16 
<< pdiffusion >>
rect 481 15 482 16 
<< pdiffusion >>
rect 482 15 483 16 
<< pdiffusion >>
rect 483 15 484 16 
<< pdiffusion >>
rect 484 15 485 16 
<< pdiffusion >>
rect 485 15 486 16 
<< pdiffusion >>
rect 498 15 499 16 
<< pdiffusion >>
rect 499 15 500 16 
<< pdiffusion >>
rect 500 15 501 16 
<< pdiffusion >>
rect 501 15 502 16 
<< pdiffusion >>
rect 502 15 503 16 
<< pdiffusion >>
rect 503 15 504 16 
<< m1 >>
rect 505 15 506 16 
<< pdiffusion >>
rect 516 15 517 16 
<< pdiffusion >>
rect 517 15 518 16 
<< pdiffusion >>
rect 518 15 519 16 
<< pdiffusion >>
rect 519 15 520 16 
<< pdiffusion >>
rect 520 15 521 16 
<< pdiffusion >>
rect 521 15 522 16 
<< pdiffusion >>
rect 12 16 13 17 
<< pdiffusion >>
rect 13 16 14 17 
<< pdiffusion >>
rect 14 16 15 17 
<< pdiffusion >>
rect 15 16 16 17 
<< pdiffusion >>
rect 16 16 17 17 
<< pdiffusion >>
rect 17 16 18 17 
<< pdiffusion >>
rect 30 16 31 17 
<< pdiffusion >>
rect 31 16 32 17 
<< pdiffusion >>
rect 32 16 33 17 
<< pdiffusion >>
rect 33 16 34 17 
<< pdiffusion >>
rect 34 16 35 17 
<< pdiffusion >>
rect 35 16 36 17 
<< pdiffusion >>
rect 48 16 49 17 
<< pdiffusion >>
rect 49 16 50 17 
<< pdiffusion >>
rect 50 16 51 17 
<< pdiffusion >>
rect 51 16 52 17 
<< pdiffusion >>
rect 52 16 53 17 
<< pdiffusion >>
rect 53 16 54 17 
<< pdiffusion >>
rect 66 16 67 17 
<< pdiffusion >>
rect 67 16 68 17 
<< pdiffusion >>
rect 68 16 69 17 
<< pdiffusion >>
rect 69 16 70 17 
<< pdiffusion >>
rect 70 16 71 17 
<< pdiffusion >>
rect 71 16 72 17 
<< pdiffusion >>
rect 102 16 103 17 
<< pdiffusion >>
rect 103 16 104 17 
<< pdiffusion >>
rect 104 16 105 17 
<< pdiffusion >>
rect 105 16 106 17 
<< pdiffusion >>
rect 106 16 107 17 
<< pdiffusion >>
rect 107 16 108 17 
<< pdiffusion >>
rect 120 16 121 17 
<< pdiffusion >>
rect 121 16 122 17 
<< pdiffusion >>
rect 122 16 123 17 
<< pdiffusion >>
rect 123 16 124 17 
<< pdiffusion >>
rect 124 16 125 17 
<< pdiffusion >>
rect 125 16 126 17 
<< pdiffusion >>
rect 138 16 139 17 
<< pdiffusion >>
rect 139 16 140 17 
<< pdiffusion >>
rect 140 16 141 17 
<< pdiffusion >>
rect 141 16 142 17 
<< pdiffusion >>
rect 142 16 143 17 
<< pdiffusion >>
rect 143 16 144 17 
<< m1 >>
rect 145 16 146 17 
<< pdiffusion >>
rect 156 16 157 17 
<< pdiffusion >>
rect 157 16 158 17 
<< pdiffusion >>
rect 158 16 159 17 
<< pdiffusion >>
rect 159 16 160 17 
<< pdiffusion >>
rect 160 16 161 17 
<< pdiffusion >>
rect 161 16 162 17 
<< pdiffusion >>
rect 174 16 175 17 
<< pdiffusion >>
rect 175 16 176 17 
<< pdiffusion >>
rect 176 16 177 17 
<< pdiffusion >>
rect 177 16 178 17 
<< pdiffusion >>
rect 178 16 179 17 
<< pdiffusion >>
rect 179 16 180 17 
<< pdiffusion >>
rect 192 16 193 17 
<< pdiffusion >>
rect 193 16 194 17 
<< pdiffusion >>
rect 194 16 195 17 
<< pdiffusion >>
rect 195 16 196 17 
<< pdiffusion >>
rect 196 16 197 17 
<< pdiffusion >>
rect 197 16 198 17 
<< pdiffusion >>
rect 210 16 211 17 
<< pdiffusion >>
rect 211 16 212 17 
<< pdiffusion >>
rect 212 16 213 17 
<< pdiffusion >>
rect 213 16 214 17 
<< pdiffusion >>
rect 214 16 215 17 
<< pdiffusion >>
rect 215 16 216 17 
<< pdiffusion >>
rect 228 16 229 17 
<< pdiffusion >>
rect 229 16 230 17 
<< pdiffusion >>
rect 230 16 231 17 
<< pdiffusion >>
rect 231 16 232 17 
<< pdiffusion >>
rect 232 16 233 17 
<< pdiffusion >>
rect 233 16 234 17 
<< pdiffusion >>
rect 246 16 247 17 
<< pdiffusion >>
rect 247 16 248 17 
<< pdiffusion >>
rect 248 16 249 17 
<< pdiffusion >>
rect 249 16 250 17 
<< pdiffusion >>
rect 250 16 251 17 
<< pdiffusion >>
rect 251 16 252 17 
<< pdiffusion >>
rect 264 16 265 17 
<< pdiffusion >>
rect 265 16 266 17 
<< pdiffusion >>
rect 266 16 267 17 
<< pdiffusion >>
rect 267 16 268 17 
<< pdiffusion >>
rect 268 16 269 17 
<< pdiffusion >>
rect 269 16 270 17 
<< m1 >>
rect 280 16 281 17 
<< pdiffusion >>
rect 282 16 283 17 
<< pdiffusion >>
rect 283 16 284 17 
<< pdiffusion >>
rect 284 16 285 17 
<< pdiffusion >>
rect 285 16 286 17 
<< pdiffusion >>
rect 286 16 287 17 
<< pdiffusion >>
rect 287 16 288 17 
<< m1 >>
rect 289 16 290 17 
<< pdiffusion >>
rect 300 16 301 17 
<< pdiffusion >>
rect 301 16 302 17 
<< pdiffusion >>
rect 302 16 303 17 
<< pdiffusion >>
rect 303 16 304 17 
<< pdiffusion >>
rect 304 16 305 17 
<< pdiffusion >>
rect 305 16 306 17 
<< pdiffusion >>
rect 318 16 319 17 
<< pdiffusion >>
rect 319 16 320 17 
<< pdiffusion >>
rect 320 16 321 17 
<< pdiffusion >>
rect 321 16 322 17 
<< pdiffusion >>
rect 322 16 323 17 
<< pdiffusion >>
rect 323 16 324 17 
<< pdiffusion >>
rect 336 16 337 17 
<< pdiffusion >>
rect 337 16 338 17 
<< pdiffusion >>
rect 338 16 339 17 
<< pdiffusion >>
rect 339 16 340 17 
<< pdiffusion >>
rect 340 16 341 17 
<< pdiffusion >>
rect 341 16 342 17 
<< pdiffusion >>
rect 354 16 355 17 
<< pdiffusion >>
rect 355 16 356 17 
<< pdiffusion >>
rect 356 16 357 17 
<< pdiffusion >>
rect 357 16 358 17 
<< pdiffusion >>
rect 358 16 359 17 
<< pdiffusion >>
rect 359 16 360 17 
<< pdiffusion >>
rect 372 16 373 17 
<< pdiffusion >>
rect 373 16 374 17 
<< pdiffusion >>
rect 374 16 375 17 
<< pdiffusion >>
rect 375 16 376 17 
<< pdiffusion >>
rect 376 16 377 17 
<< pdiffusion >>
rect 377 16 378 17 
<< pdiffusion >>
rect 390 16 391 17 
<< pdiffusion >>
rect 391 16 392 17 
<< pdiffusion >>
rect 392 16 393 17 
<< pdiffusion >>
rect 393 16 394 17 
<< pdiffusion >>
rect 394 16 395 17 
<< pdiffusion >>
rect 395 16 396 17 
<< pdiffusion >>
rect 408 16 409 17 
<< pdiffusion >>
rect 409 16 410 17 
<< pdiffusion >>
rect 410 16 411 17 
<< pdiffusion >>
rect 411 16 412 17 
<< pdiffusion >>
rect 412 16 413 17 
<< pdiffusion >>
rect 413 16 414 17 
<< pdiffusion >>
rect 426 16 427 17 
<< pdiffusion >>
rect 427 16 428 17 
<< pdiffusion >>
rect 428 16 429 17 
<< pdiffusion >>
rect 429 16 430 17 
<< pdiffusion >>
rect 430 16 431 17 
<< pdiffusion >>
rect 431 16 432 17 
<< pdiffusion >>
rect 444 16 445 17 
<< pdiffusion >>
rect 445 16 446 17 
<< pdiffusion >>
rect 446 16 447 17 
<< pdiffusion >>
rect 447 16 448 17 
<< pdiffusion >>
rect 448 16 449 17 
<< pdiffusion >>
rect 449 16 450 17 
<< pdiffusion >>
rect 462 16 463 17 
<< pdiffusion >>
rect 463 16 464 17 
<< pdiffusion >>
rect 464 16 465 17 
<< pdiffusion >>
rect 465 16 466 17 
<< pdiffusion >>
rect 466 16 467 17 
<< pdiffusion >>
rect 467 16 468 17 
<< pdiffusion >>
rect 480 16 481 17 
<< pdiffusion >>
rect 481 16 482 17 
<< pdiffusion >>
rect 482 16 483 17 
<< pdiffusion >>
rect 483 16 484 17 
<< pdiffusion >>
rect 484 16 485 17 
<< pdiffusion >>
rect 485 16 486 17 
<< pdiffusion >>
rect 498 16 499 17 
<< pdiffusion >>
rect 499 16 500 17 
<< pdiffusion >>
rect 500 16 501 17 
<< pdiffusion >>
rect 501 16 502 17 
<< pdiffusion >>
rect 502 16 503 17 
<< pdiffusion >>
rect 503 16 504 17 
<< m1 >>
rect 505 16 506 17 
<< pdiffusion >>
rect 516 16 517 17 
<< pdiffusion >>
rect 517 16 518 17 
<< pdiffusion >>
rect 518 16 519 17 
<< pdiffusion >>
rect 519 16 520 17 
<< pdiffusion >>
rect 520 16 521 17 
<< pdiffusion >>
rect 521 16 522 17 
<< pdiffusion >>
rect 12 17 13 18 
<< pdiffusion >>
rect 13 17 14 18 
<< pdiffusion >>
rect 14 17 15 18 
<< pdiffusion >>
rect 15 17 16 18 
<< pdiffusion >>
rect 16 17 17 18 
<< pdiffusion >>
rect 17 17 18 18 
<< pdiffusion >>
rect 30 17 31 18 
<< pdiffusion >>
rect 31 17 32 18 
<< pdiffusion >>
rect 32 17 33 18 
<< pdiffusion >>
rect 33 17 34 18 
<< pdiffusion >>
rect 34 17 35 18 
<< pdiffusion >>
rect 35 17 36 18 
<< pdiffusion >>
rect 48 17 49 18 
<< pdiffusion >>
rect 49 17 50 18 
<< pdiffusion >>
rect 50 17 51 18 
<< pdiffusion >>
rect 51 17 52 18 
<< pdiffusion >>
rect 52 17 53 18 
<< pdiffusion >>
rect 53 17 54 18 
<< pdiffusion >>
rect 66 17 67 18 
<< pdiffusion >>
rect 67 17 68 18 
<< pdiffusion >>
rect 68 17 69 18 
<< pdiffusion >>
rect 69 17 70 18 
<< pdiffusion >>
rect 70 17 71 18 
<< pdiffusion >>
rect 71 17 72 18 
<< pdiffusion >>
rect 102 17 103 18 
<< pdiffusion >>
rect 103 17 104 18 
<< pdiffusion >>
rect 104 17 105 18 
<< pdiffusion >>
rect 105 17 106 18 
<< m1 >>
rect 106 17 107 18 
<< pdiffusion >>
rect 106 17 107 18 
<< pdiffusion >>
rect 107 17 108 18 
<< pdiffusion >>
rect 120 17 121 18 
<< pdiffusion >>
rect 121 17 122 18 
<< pdiffusion >>
rect 122 17 123 18 
<< pdiffusion >>
rect 123 17 124 18 
<< pdiffusion >>
rect 124 17 125 18 
<< pdiffusion >>
rect 125 17 126 18 
<< pdiffusion >>
rect 138 17 139 18 
<< pdiffusion >>
rect 139 17 140 18 
<< pdiffusion >>
rect 140 17 141 18 
<< pdiffusion >>
rect 141 17 142 18 
<< pdiffusion >>
rect 142 17 143 18 
<< pdiffusion >>
rect 143 17 144 18 
<< m1 >>
rect 145 17 146 18 
<< pdiffusion >>
rect 156 17 157 18 
<< pdiffusion >>
rect 157 17 158 18 
<< pdiffusion >>
rect 158 17 159 18 
<< pdiffusion >>
rect 159 17 160 18 
<< pdiffusion >>
rect 160 17 161 18 
<< pdiffusion >>
rect 161 17 162 18 
<< pdiffusion >>
rect 174 17 175 18 
<< pdiffusion >>
rect 175 17 176 18 
<< pdiffusion >>
rect 176 17 177 18 
<< pdiffusion >>
rect 177 17 178 18 
<< pdiffusion >>
rect 178 17 179 18 
<< pdiffusion >>
rect 179 17 180 18 
<< pdiffusion >>
rect 192 17 193 18 
<< pdiffusion >>
rect 193 17 194 18 
<< pdiffusion >>
rect 194 17 195 18 
<< pdiffusion >>
rect 195 17 196 18 
<< pdiffusion >>
rect 196 17 197 18 
<< pdiffusion >>
rect 197 17 198 18 
<< pdiffusion >>
rect 210 17 211 18 
<< pdiffusion >>
rect 211 17 212 18 
<< pdiffusion >>
rect 212 17 213 18 
<< pdiffusion >>
rect 213 17 214 18 
<< m1 >>
rect 214 17 215 18 
<< pdiffusion >>
rect 214 17 215 18 
<< pdiffusion >>
rect 215 17 216 18 
<< pdiffusion >>
rect 228 17 229 18 
<< m1 >>
rect 229 17 230 18 
<< pdiffusion >>
rect 229 17 230 18 
<< pdiffusion >>
rect 230 17 231 18 
<< pdiffusion >>
rect 231 17 232 18 
<< pdiffusion >>
rect 232 17 233 18 
<< pdiffusion >>
rect 233 17 234 18 
<< pdiffusion >>
rect 246 17 247 18 
<< pdiffusion >>
rect 247 17 248 18 
<< pdiffusion >>
rect 248 17 249 18 
<< pdiffusion >>
rect 249 17 250 18 
<< pdiffusion >>
rect 250 17 251 18 
<< pdiffusion >>
rect 251 17 252 18 
<< pdiffusion >>
rect 264 17 265 18 
<< m1 >>
rect 265 17 266 18 
<< pdiffusion >>
rect 265 17 266 18 
<< pdiffusion >>
rect 266 17 267 18 
<< pdiffusion >>
rect 267 17 268 18 
<< pdiffusion >>
rect 268 17 269 18 
<< pdiffusion >>
rect 269 17 270 18 
<< m1 >>
rect 280 17 281 18 
<< pdiffusion >>
rect 282 17 283 18 
<< pdiffusion >>
rect 283 17 284 18 
<< pdiffusion >>
rect 284 17 285 18 
<< pdiffusion >>
rect 285 17 286 18 
<< pdiffusion >>
rect 286 17 287 18 
<< pdiffusion >>
rect 287 17 288 18 
<< m1 >>
rect 289 17 290 18 
<< pdiffusion >>
rect 300 17 301 18 
<< pdiffusion >>
rect 301 17 302 18 
<< pdiffusion >>
rect 302 17 303 18 
<< pdiffusion >>
rect 303 17 304 18 
<< pdiffusion >>
rect 304 17 305 18 
<< pdiffusion >>
rect 305 17 306 18 
<< pdiffusion >>
rect 318 17 319 18 
<< pdiffusion >>
rect 319 17 320 18 
<< pdiffusion >>
rect 320 17 321 18 
<< pdiffusion >>
rect 321 17 322 18 
<< pdiffusion >>
rect 322 17 323 18 
<< pdiffusion >>
rect 323 17 324 18 
<< pdiffusion >>
rect 336 17 337 18 
<< pdiffusion >>
rect 337 17 338 18 
<< pdiffusion >>
rect 338 17 339 18 
<< pdiffusion >>
rect 339 17 340 18 
<< m1 >>
rect 340 17 341 18 
<< pdiffusion >>
rect 340 17 341 18 
<< pdiffusion >>
rect 341 17 342 18 
<< pdiffusion >>
rect 354 17 355 18 
<< pdiffusion >>
rect 355 17 356 18 
<< pdiffusion >>
rect 356 17 357 18 
<< pdiffusion >>
rect 357 17 358 18 
<< pdiffusion >>
rect 358 17 359 18 
<< pdiffusion >>
rect 359 17 360 18 
<< pdiffusion >>
rect 372 17 373 18 
<< pdiffusion >>
rect 373 17 374 18 
<< pdiffusion >>
rect 374 17 375 18 
<< pdiffusion >>
rect 375 17 376 18 
<< pdiffusion >>
rect 376 17 377 18 
<< pdiffusion >>
rect 377 17 378 18 
<< pdiffusion >>
rect 390 17 391 18 
<< m1 >>
rect 391 17 392 18 
<< pdiffusion >>
rect 391 17 392 18 
<< pdiffusion >>
rect 392 17 393 18 
<< pdiffusion >>
rect 393 17 394 18 
<< pdiffusion >>
rect 394 17 395 18 
<< pdiffusion >>
rect 395 17 396 18 
<< pdiffusion >>
rect 408 17 409 18 
<< m1 >>
rect 409 17 410 18 
<< pdiffusion >>
rect 409 17 410 18 
<< pdiffusion >>
rect 410 17 411 18 
<< pdiffusion >>
rect 411 17 412 18 
<< pdiffusion >>
rect 412 17 413 18 
<< pdiffusion >>
rect 413 17 414 18 
<< pdiffusion >>
rect 426 17 427 18 
<< pdiffusion >>
rect 427 17 428 18 
<< pdiffusion >>
rect 428 17 429 18 
<< pdiffusion >>
rect 429 17 430 18 
<< pdiffusion >>
rect 430 17 431 18 
<< pdiffusion >>
rect 431 17 432 18 
<< pdiffusion >>
rect 444 17 445 18 
<< pdiffusion >>
rect 445 17 446 18 
<< pdiffusion >>
rect 446 17 447 18 
<< pdiffusion >>
rect 447 17 448 18 
<< m1 >>
rect 448 17 449 18 
<< pdiffusion >>
rect 448 17 449 18 
<< pdiffusion >>
rect 449 17 450 18 
<< pdiffusion >>
rect 462 17 463 18 
<< pdiffusion >>
rect 463 17 464 18 
<< pdiffusion >>
rect 464 17 465 18 
<< pdiffusion >>
rect 465 17 466 18 
<< pdiffusion >>
rect 466 17 467 18 
<< pdiffusion >>
rect 467 17 468 18 
<< pdiffusion >>
rect 480 17 481 18 
<< pdiffusion >>
rect 481 17 482 18 
<< pdiffusion >>
rect 482 17 483 18 
<< pdiffusion >>
rect 483 17 484 18 
<< pdiffusion >>
rect 484 17 485 18 
<< pdiffusion >>
rect 485 17 486 18 
<< pdiffusion >>
rect 498 17 499 18 
<< pdiffusion >>
rect 499 17 500 18 
<< pdiffusion >>
rect 500 17 501 18 
<< pdiffusion >>
rect 501 17 502 18 
<< pdiffusion >>
rect 502 17 503 18 
<< pdiffusion >>
rect 503 17 504 18 
<< m1 >>
rect 505 17 506 18 
<< pdiffusion >>
rect 516 17 517 18 
<< pdiffusion >>
rect 517 17 518 18 
<< pdiffusion >>
rect 518 17 519 18 
<< pdiffusion >>
rect 519 17 520 18 
<< pdiffusion >>
rect 520 17 521 18 
<< pdiffusion >>
rect 521 17 522 18 
<< m1 >>
rect 106 18 107 19 
<< m1 >>
rect 145 18 146 19 
<< m1 >>
rect 214 18 215 19 
<< m1 >>
rect 229 18 230 19 
<< m1 >>
rect 265 18 266 19 
<< m1 >>
rect 280 18 281 19 
<< m1 >>
rect 289 18 290 19 
<< m1 >>
rect 340 18 341 19 
<< m1 >>
rect 391 18 392 19 
<< m1 >>
rect 409 18 410 19 
<< m1 >>
rect 448 18 449 19 
<< m1 >>
rect 505 18 506 19 
<< m1 >>
rect 106 19 107 20 
<< m1 >>
rect 145 19 146 20 
<< m1 >>
rect 214 19 215 20 
<< m1 >>
rect 229 19 230 20 
<< m1 >>
rect 265 19 266 20 
<< m1 >>
rect 280 19 281 20 
<< m1 >>
rect 289 19 290 20 
<< m1 >>
rect 340 19 341 20 
<< m1 >>
rect 388 19 389 20 
<< m1 >>
rect 389 19 390 20 
<< m1 >>
rect 390 19 391 20 
<< m1 >>
rect 391 19 392 20 
<< m1 >>
rect 409 19 410 20 
<< m1 >>
rect 448 19 449 20 
<< m1 >>
rect 505 19 506 20 
<< m1 >>
rect 106 20 107 21 
<< m1 >>
rect 145 20 146 21 
<< m1 >>
rect 214 20 215 21 
<< m1 >>
rect 229 20 230 21 
<< m2 >>
rect 229 20 230 21 
<< m2c >>
rect 229 20 230 21 
<< m1 >>
rect 229 20 230 21 
<< m2 >>
rect 229 20 230 21 
<< m1 >>
rect 265 20 266 21 
<< m1 >>
rect 280 20 281 21 
<< m1 >>
rect 289 20 290 21 
<< m1 >>
rect 340 20 341 21 
<< m1 >>
rect 388 20 389 21 
<< m1 >>
rect 409 20 410 21 
<< m1 >>
rect 448 20 449 21 
<< m1 >>
rect 505 20 506 21 
<< m1 >>
rect 106 21 107 22 
<< m1 >>
rect 145 21 146 22 
<< m1 >>
rect 214 21 215 22 
<< m2 >>
rect 229 21 230 22 
<< m1 >>
rect 265 21 266 22 
<< m1 >>
rect 280 21 281 22 
<< m1 >>
rect 289 21 290 22 
<< m1 >>
rect 340 21 341 22 
<< m1 >>
rect 388 21 389 22 
<< m1 >>
rect 409 21 410 22 
<< m1 >>
rect 448 21 449 22 
<< m1 >>
rect 505 21 506 22 
<< m1 >>
rect 106 22 107 23 
<< m1 >>
rect 107 22 108 23 
<< m1 >>
rect 108 22 109 23 
<< m1 >>
rect 109 22 110 23 
<< m1 >>
rect 110 22 111 23 
<< m1 >>
rect 111 22 112 23 
<< m1 >>
rect 112 22 113 23 
<< m1 >>
rect 113 22 114 23 
<< m1 >>
rect 114 22 115 23 
<< m1 >>
rect 115 22 116 23 
<< m1 >>
rect 116 22 117 23 
<< m1 >>
rect 117 22 118 23 
<< m1 >>
rect 118 22 119 23 
<< m1 >>
rect 119 22 120 23 
<< m1 >>
rect 120 22 121 23 
<< m1 >>
rect 121 22 122 23 
<< m1 >>
rect 122 22 123 23 
<< m1 >>
rect 123 22 124 23 
<< m1 >>
rect 124 22 125 23 
<< m1 >>
rect 145 22 146 23 
<< m1 >>
rect 214 22 215 23 
<< m1 >>
rect 228 22 229 23 
<< m1 >>
rect 229 22 230 23 
<< m2 >>
rect 229 22 230 23 
<< m1 >>
rect 230 22 231 23 
<< m1 >>
rect 231 22 232 23 
<< m1 >>
rect 232 22 233 23 
<< m1 >>
rect 233 22 234 23 
<< m1 >>
rect 234 22 235 23 
<< m1 >>
rect 235 22 236 23 
<< m1 >>
rect 236 22 237 23 
<< m1 >>
rect 237 22 238 23 
<< m1 >>
rect 238 22 239 23 
<< m1 >>
rect 239 22 240 23 
<< m1 >>
rect 240 22 241 23 
<< m1 >>
rect 241 22 242 23 
<< m1 >>
rect 242 22 243 23 
<< m1 >>
rect 243 22 244 23 
<< m1 >>
rect 244 22 245 23 
<< m1 >>
rect 245 22 246 23 
<< m1 >>
rect 246 22 247 23 
<< m1 >>
rect 247 22 248 23 
<< m1 >>
rect 248 22 249 23 
<< m1 >>
rect 249 22 250 23 
<< m1 >>
rect 250 22 251 23 
<< m1 >>
rect 251 22 252 23 
<< m1 >>
rect 252 22 253 23 
<< m1 >>
rect 253 22 254 23 
<< m1 >>
rect 254 22 255 23 
<< m1 >>
rect 255 22 256 23 
<< m1 >>
rect 256 22 257 23 
<< m1 >>
rect 257 22 258 23 
<< m1 >>
rect 258 22 259 23 
<< m1 >>
rect 259 22 260 23 
<< m1 >>
rect 260 22 261 23 
<< m1 >>
rect 261 22 262 23 
<< m1 >>
rect 262 22 263 23 
<< m1 >>
rect 263 22 264 23 
<< m1 >>
rect 264 22 265 23 
<< m1 >>
rect 265 22 266 23 
<< m1 >>
rect 278 22 279 23 
<< m2 >>
rect 278 22 279 23 
<< m2c >>
rect 278 22 279 23 
<< m1 >>
rect 278 22 279 23 
<< m2 >>
rect 278 22 279 23 
<< m2 >>
rect 279 22 280 23 
<< m1 >>
rect 280 22 281 23 
<< m2 >>
rect 280 22 281 23 
<< m2 >>
rect 281 22 282 23 
<< m1 >>
rect 282 22 283 23 
<< m2 >>
rect 282 22 283 23 
<< m2c >>
rect 282 22 283 23 
<< m1 >>
rect 282 22 283 23 
<< m2 >>
rect 282 22 283 23 
<< m1 >>
rect 283 22 284 23 
<< m1 >>
rect 284 22 285 23 
<< m1 >>
rect 285 22 286 23 
<< m1 >>
rect 286 22 287 23 
<< m1 >>
rect 287 22 288 23 
<< m2 >>
rect 287 22 288 23 
<< m2c >>
rect 287 22 288 23 
<< m1 >>
rect 287 22 288 23 
<< m2 >>
rect 287 22 288 23 
<< m2 >>
rect 288 22 289 23 
<< m1 >>
rect 289 22 290 23 
<< m2 >>
rect 289 22 290 23 
<< m2 >>
rect 290 22 291 23 
<< m1 >>
rect 291 22 292 23 
<< m2 >>
rect 291 22 292 23 
<< m2c >>
rect 291 22 292 23 
<< m1 >>
rect 291 22 292 23 
<< m2 >>
rect 291 22 292 23 
<< m1 >>
rect 292 22 293 23 
<< m1 >>
rect 293 22 294 23 
<< m1 >>
rect 294 22 295 23 
<< m1 >>
rect 295 22 296 23 
<< m1 >>
rect 296 22 297 23 
<< m1 >>
rect 297 22 298 23 
<< m1 >>
rect 298 22 299 23 
<< m1 >>
rect 299 22 300 23 
<< m1 >>
rect 300 22 301 23 
<< m1 >>
rect 301 22 302 23 
<< m1 >>
rect 302 22 303 23 
<< m1 >>
rect 303 22 304 23 
<< m1 >>
rect 304 22 305 23 
<< m1 >>
rect 305 22 306 23 
<< m1 >>
rect 306 22 307 23 
<< m1 >>
rect 307 22 308 23 
<< m1 >>
rect 308 22 309 23 
<< m1 >>
rect 309 22 310 23 
<< m1 >>
rect 310 22 311 23 
<< m1 >>
rect 311 22 312 23 
<< m1 >>
rect 312 22 313 23 
<< m1 >>
rect 313 22 314 23 
<< m1 >>
rect 314 22 315 23 
<< m1 >>
rect 315 22 316 23 
<< m1 >>
rect 316 22 317 23 
<< m1 >>
rect 317 22 318 23 
<< m1 >>
rect 318 22 319 23 
<< m1 >>
rect 319 22 320 23 
<< m1 >>
rect 320 22 321 23 
<< m1 >>
rect 321 22 322 23 
<< m1 >>
rect 322 22 323 23 
<< m1 >>
rect 323 22 324 23 
<< m1 >>
rect 324 22 325 23 
<< m1 >>
rect 325 22 326 23 
<< m1 >>
rect 326 22 327 23 
<< m1 >>
rect 327 22 328 23 
<< m1 >>
rect 328 22 329 23 
<< m1 >>
rect 329 22 330 23 
<< m1 >>
rect 330 22 331 23 
<< m1 >>
rect 331 22 332 23 
<< m1 >>
rect 332 22 333 23 
<< m2 >>
rect 332 22 333 23 
<< m2c >>
rect 332 22 333 23 
<< m1 >>
rect 332 22 333 23 
<< m2 >>
rect 332 22 333 23 
<< m2 >>
rect 333 22 334 23 
<< m1 >>
rect 334 22 335 23 
<< m2 >>
rect 334 22 335 23 
<< m1 >>
rect 335 22 336 23 
<< m2 >>
rect 335 22 336 23 
<< m1 >>
rect 336 22 337 23 
<< m2 >>
rect 336 22 337 23 
<< m1 >>
rect 337 22 338 23 
<< m2 >>
rect 337 22 338 23 
<< m1 >>
rect 338 22 339 23 
<< m2 >>
rect 338 22 339 23 
<< m1 >>
rect 339 22 340 23 
<< m2 >>
rect 339 22 340 23 
<< m1 >>
rect 340 22 341 23 
<< m2 >>
rect 340 22 341 23 
<< m2 >>
rect 341 22 342 23 
<< m1 >>
rect 342 22 343 23 
<< m2 >>
rect 342 22 343 23 
<< m2c >>
rect 342 22 343 23 
<< m1 >>
rect 342 22 343 23 
<< m2 >>
rect 342 22 343 23 
<< m1 >>
rect 343 22 344 23 
<< m1 >>
rect 344 22 345 23 
<< m1 >>
rect 345 22 346 23 
<< m1 >>
rect 346 22 347 23 
<< m1 >>
rect 347 22 348 23 
<< m1 >>
rect 348 22 349 23 
<< m1 >>
rect 349 22 350 23 
<< m1 >>
rect 350 22 351 23 
<< m1 >>
rect 351 22 352 23 
<< m1 >>
rect 352 22 353 23 
<< m1 >>
rect 353 22 354 23 
<< m1 >>
rect 354 22 355 23 
<< m1 >>
rect 355 22 356 23 
<< m1 >>
rect 356 22 357 23 
<< m1 >>
rect 357 22 358 23 
<< m1 >>
rect 358 22 359 23 
<< m1 >>
rect 359 22 360 23 
<< m1 >>
rect 360 22 361 23 
<< m1 >>
rect 361 22 362 23 
<< m1 >>
rect 362 22 363 23 
<< m1 >>
rect 363 22 364 23 
<< m1 >>
rect 364 22 365 23 
<< m1 >>
rect 365 22 366 23 
<< m1 >>
rect 366 22 367 23 
<< m1 >>
rect 367 22 368 23 
<< m1 >>
rect 368 22 369 23 
<< m1 >>
rect 369 22 370 23 
<< m1 >>
rect 370 22 371 23 
<< m1 >>
rect 371 22 372 23 
<< m1 >>
rect 372 22 373 23 
<< m1 >>
rect 373 22 374 23 
<< m1 >>
rect 374 22 375 23 
<< m1 >>
rect 375 22 376 23 
<< m1 >>
rect 376 22 377 23 
<< m1 >>
rect 377 22 378 23 
<< m1 >>
rect 378 22 379 23 
<< m1 >>
rect 379 22 380 23 
<< m1 >>
rect 380 22 381 23 
<< m1 >>
rect 381 22 382 23 
<< m1 >>
rect 382 22 383 23 
<< m1 >>
rect 383 22 384 23 
<< m1 >>
rect 384 22 385 23 
<< m1 >>
rect 385 22 386 23 
<< m1 >>
rect 386 22 387 23 
<< m2 >>
rect 386 22 387 23 
<< m2c >>
rect 386 22 387 23 
<< m1 >>
rect 386 22 387 23 
<< m2 >>
rect 386 22 387 23 
<< m2 >>
rect 387 22 388 23 
<< m1 >>
rect 388 22 389 23 
<< m2 >>
rect 388 22 389 23 
<< m2 >>
rect 389 22 390 23 
<< m1 >>
rect 390 22 391 23 
<< m2 >>
rect 390 22 391 23 
<< m2c >>
rect 390 22 391 23 
<< m1 >>
rect 390 22 391 23 
<< m2 >>
rect 390 22 391 23 
<< m1 >>
rect 391 22 392 23 
<< m1 >>
rect 392 22 393 23 
<< m1 >>
rect 393 22 394 23 
<< m1 >>
rect 394 22 395 23 
<< m1 >>
rect 395 22 396 23 
<< m1 >>
rect 396 22 397 23 
<< m1 >>
rect 397 22 398 23 
<< m1 >>
rect 398 22 399 23 
<< m1 >>
rect 399 22 400 23 
<< m1 >>
rect 400 22 401 23 
<< m1 >>
rect 401 22 402 23 
<< m1 >>
rect 402 22 403 23 
<< m1 >>
rect 403 22 404 23 
<< m1 >>
rect 404 22 405 23 
<< m1 >>
rect 405 22 406 23 
<< m1 >>
rect 406 22 407 23 
<< m1 >>
rect 407 22 408 23 
<< m1 >>
rect 408 22 409 23 
<< m1 >>
rect 409 22 410 23 
<< m1 >>
rect 448 22 449 23 
<< m1 >>
rect 505 22 506 23 
<< m1 >>
rect 124 23 125 24 
<< m1 >>
rect 145 23 146 24 
<< m1 >>
rect 214 23 215 24 
<< m1 >>
rect 228 23 229 24 
<< m2 >>
rect 229 23 230 24 
<< m1 >>
rect 278 23 279 24 
<< m1 >>
rect 280 23 281 24 
<< m1 >>
rect 289 23 290 24 
<< m1 >>
rect 334 23 335 24 
<< m1 >>
rect 388 23 389 24 
<< m1 >>
rect 448 23 449 24 
<< m1 >>
rect 487 23 488 24 
<< m1 >>
rect 488 23 489 24 
<< m1 >>
rect 489 23 490 24 
<< m1 >>
rect 490 23 491 24 
<< m1 >>
rect 491 23 492 24 
<< m1 >>
rect 492 23 493 24 
<< m1 >>
rect 493 23 494 24 
<< m1 >>
rect 494 23 495 24 
<< m1 >>
rect 495 23 496 24 
<< m1 >>
rect 496 23 497 24 
<< m1 >>
rect 497 23 498 24 
<< m1 >>
rect 498 23 499 24 
<< m1 >>
rect 499 23 500 24 
<< m1 >>
rect 500 23 501 24 
<< m1 >>
rect 501 23 502 24 
<< m1 >>
rect 502 23 503 24 
<< m1 >>
rect 503 23 504 24 
<< m1 >>
rect 504 23 505 24 
<< m1 >>
rect 505 23 506 24 
<< m1 >>
rect 124 24 125 25 
<< m1 >>
rect 145 24 146 25 
<< m1 >>
rect 214 24 215 25 
<< m1 >>
rect 228 24 229 25 
<< m2 >>
rect 229 24 230 25 
<< m1 >>
rect 230 24 231 25 
<< m2 >>
rect 230 24 231 25 
<< m2c >>
rect 230 24 231 25 
<< m1 >>
rect 230 24 231 25 
<< m2 >>
rect 230 24 231 25 
<< m1 >>
rect 231 24 232 25 
<< m1 >>
rect 232 24 233 25 
<< m1 >>
rect 233 24 234 25 
<< m1 >>
rect 234 24 235 25 
<< m1 >>
rect 235 24 236 25 
<< m1 >>
rect 278 24 279 25 
<< m1 >>
rect 280 24 281 25 
<< m1 >>
rect 289 24 290 25 
<< m1 >>
rect 334 24 335 25 
<< m1 >>
rect 388 24 389 25 
<< m1 >>
rect 448 24 449 25 
<< m1 >>
rect 487 24 488 25 
<< m1 >>
rect 124 25 125 26 
<< m1 >>
rect 127 25 128 26 
<< m1 >>
rect 128 25 129 26 
<< m1 >>
rect 129 25 130 26 
<< m1 >>
rect 130 25 131 26 
<< m1 >>
rect 131 25 132 26 
<< m1 >>
rect 132 25 133 26 
<< m1 >>
rect 133 25 134 26 
<< m1 >>
rect 134 25 135 26 
<< m1 >>
rect 135 25 136 26 
<< m1 >>
rect 136 25 137 26 
<< m1 >>
rect 137 25 138 26 
<< m1 >>
rect 138 25 139 26 
<< m1 >>
rect 139 25 140 26 
<< m1 >>
rect 140 25 141 26 
<< m1 >>
rect 141 25 142 26 
<< m1 >>
rect 142 25 143 26 
<< m1 >>
rect 145 25 146 26 
<< m1 >>
rect 214 25 215 26 
<< m1 >>
rect 228 25 229 26 
<< m1 >>
rect 235 25 236 26 
<< m1 >>
rect 278 25 279 26 
<< m1 >>
rect 280 25 281 26 
<< m1 >>
rect 289 25 290 26 
<< m1 >>
rect 334 25 335 26 
<< m1 >>
rect 388 25 389 26 
<< m1 >>
rect 448 25 449 26 
<< m1 >>
rect 487 25 488 26 
<< m1 >>
rect 505 25 506 26 
<< m1 >>
rect 506 25 507 26 
<< m1 >>
rect 507 25 508 26 
<< m1 >>
rect 508 25 509 26 
<< m1 >>
rect 509 25 510 26 
<< m1 >>
rect 510 25 511 26 
<< m1 >>
rect 511 25 512 26 
<< m1 >>
rect 512 25 513 26 
<< m1 >>
rect 513 25 514 26 
<< m1 >>
rect 514 25 515 26 
<< m1 >>
rect 515 25 516 26 
<< m1 >>
rect 516 25 517 26 
<< m1 >>
rect 517 25 518 26 
<< m1 >>
rect 518 25 519 26 
<< m1 >>
rect 519 25 520 26 
<< m1 >>
rect 520 25 521 26 
<< m1 >>
rect 124 26 125 27 
<< m1 >>
rect 127 26 128 27 
<< m1 >>
rect 142 26 143 27 
<< m1 >>
rect 145 26 146 27 
<< m1 >>
rect 214 26 215 27 
<< m2 >>
rect 225 26 226 27 
<< m2 >>
rect 226 26 227 27 
<< m2 >>
rect 227 26 228 27 
<< m1 >>
rect 228 26 229 27 
<< m2 >>
rect 228 26 229 27 
<< m2c >>
rect 228 26 229 27 
<< m1 >>
rect 228 26 229 27 
<< m2 >>
rect 228 26 229 27 
<< m1 >>
rect 235 26 236 27 
<< m1 >>
rect 278 26 279 27 
<< m1 >>
rect 280 26 281 27 
<< m1 >>
rect 289 26 290 27 
<< m1 >>
rect 334 26 335 27 
<< m1 >>
rect 388 26 389 27 
<< m1 >>
rect 448 26 449 27 
<< m1 >>
rect 487 26 488 27 
<< m1 >>
rect 505 26 506 27 
<< m1 >>
rect 520 26 521 27 
<< m1 >>
rect 124 27 125 28 
<< m1 >>
rect 127 27 128 28 
<< m1 >>
rect 142 27 143 28 
<< m1 >>
rect 145 27 146 28 
<< m1 >>
rect 193 27 194 28 
<< m1 >>
rect 194 27 195 28 
<< m1 >>
rect 195 27 196 28 
<< m1 >>
rect 196 27 197 28 
<< m1 >>
rect 197 27 198 28 
<< m1 >>
rect 198 27 199 28 
<< m1 >>
rect 199 27 200 28 
<< m1 >>
rect 200 27 201 28 
<< m1 >>
rect 201 27 202 28 
<< m1 >>
rect 202 27 203 28 
<< m1 >>
rect 203 27 204 28 
<< m1 >>
rect 204 27 205 28 
<< m1 >>
rect 205 27 206 28 
<< m1 >>
rect 206 27 207 28 
<< m1 >>
rect 207 27 208 28 
<< m1 >>
rect 208 27 209 28 
<< m1 >>
rect 214 27 215 28 
<< m1 >>
rect 215 27 216 28 
<< m1 >>
rect 216 27 217 28 
<< m1 >>
rect 217 27 218 28 
<< m1 >>
rect 218 27 219 28 
<< m1 >>
rect 219 27 220 28 
<< m1 >>
rect 220 27 221 28 
<< m1 >>
rect 221 27 222 28 
<< m1 >>
rect 222 27 223 28 
<< m1 >>
rect 223 27 224 28 
<< m1 >>
rect 224 27 225 28 
<< m1 >>
rect 225 27 226 28 
<< m2 >>
rect 225 27 226 28 
<< m1 >>
rect 226 27 227 28 
<< m1 >>
rect 235 27 236 28 
<< m1 >>
rect 278 27 279 28 
<< m1 >>
rect 280 27 281 28 
<< m1 >>
rect 289 27 290 28 
<< m1 >>
rect 334 27 335 28 
<< m1 >>
rect 388 27 389 28 
<< m1 >>
rect 448 27 449 28 
<< m1 >>
rect 487 27 488 28 
<< m1 >>
rect 505 27 506 28 
<< m1 >>
rect 520 27 521 28 
<< m1 >>
rect 64 28 65 29 
<< m1 >>
rect 65 28 66 29 
<< m1 >>
rect 66 28 67 29 
<< m1 >>
rect 67 28 68 29 
<< m1 >>
rect 106 28 107 29 
<< m1 >>
rect 107 28 108 29 
<< m1 >>
rect 108 28 109 29 
<< m1 >>
rect 109 28 110 29 
<< m1 >>
rect 110 28 111 29 
<< m1 >>
rect 111 28 112 29 
<< m1 >>
rect 124 28 125 29 
<< m1 >>
rect 127 28 128 29 
<< m1 >>
rect 142 28 143 29 
<< m1 >>
rect 145 28 146 29 
<< m1 >>
rect 193 28 194 29 
<< m1 >>
rect 208 28 209 29 
<< m2 >>
rect 225 28 226 29 
<< m1 >>
rect 226 28 227 29 
<< m1 >>
rect 235 28 236 29 
<< m1 >>
rect 278 28 279 29 
<< m1 >>
rect 280 28 281 29 
<< m1 >>
rect 286 28 287 29 
<< m1 >>
rect 287 28 288 29 
<< m1 >>
rect 288 28 289 29 
<< m1 >>
rect 289 28 290 29 
<< m1 >>
rect 334 28 335 29 
<< m1 >>
rect 388 28 389 29 
<< m1 >>
rect 406 28 407 29 
<< m1 >>
rect 407 28 408 29 
<< m1 >>
rect 408 28 409 29 
<< m1 >>
rect 409 28 410 29 
<< m1 >>
rect 430 28 431 29 
<< m1 >>
rect 431 28 432 29 
<< m1 >>
rect 432 28 433 29 
<< m1 >>
rect 433 28 434 29 
<< m1 >>
rect 448 28 449 29 
<< m1 >>
rect 487 28 488 29 
<< m1 >>
rect 505 28 506 29 
<< m1 >>
rect 520 28 521 29 
<< m1 >>
rect 64 29 65 30 
<< m1 >>
rect 67 29 68 30 
<< m1 >>
rect 106 29 107 30 
<< m1 >>
rect 111 29 112 30 
<< m1 >>
rect 124 29 125 30 
<< m1 >>
rect 127 29 128 30 
<< m1 >>
rect 142 29 143 30 
<< m1 >>
rect 145 29 146 30 
<< m1 >>
rect 193 29 194 30 
<< m1 >>
rect 208 29 209 30 
<< m2 >>
rect 225 29 226 30 
<< m1 >>
rect 226 29 227 30 
<< m1 >>
rect 235 29 236 30 
<< m1 >>
rect 278 29 279 30 
<< m1 >>
rect 280 29 281 30 
<< m1 >>
rect 286 29 287 30 
<< m1 >>
rect 334 29 335 30 
<< m1 >>
rect 388 29 389 30 
<< m1 >>
rect 406 29 407 30 
<< m1 >>
rect 409 29 410 30 
<< m1 >>
rect 430 29 431 30 
<< m1 >>
rect 433 29 434 30 
<< m1 >>
rect 448 29 449 30 
<< m1 >>
rect 487 29 488 30 
<< m1 >>
rect 505 29 506 30 
<< m1 >>
rect 520 29 521 30 
<< pdiffusion >>
rect 12 30 13 31 
<< pdiffusion >>
rect 13 30 14 31 
<< pdiffusion >>
rect 14 30 15 31 
<< pdiffusion >>
rect 15 30 16 31 
<< pdiffusion >>
rect 16 30 17 31 
<< pdiffusion >>
rect 17 30 18 31 
<< pdiffusion >>
rect 30 30 31 31 
<< pdiffusion >>
rect 31 30 32 31 
<< pdiffusion >>
rect 32 30 33 31 
<< pdiffusion >>
rect 33 30 34 31 
<< pdiffusion >>
rect 34 30 35 31 
<< pdiffusion >>
rect 35 30 36 31 
<< pdiffusion >>
rect 48 30 49 31 
<< pdiffusion >>
rect 49 30 50 31 
<< pdiffusion >>
rect 50 30 51 31 
<< pdiffusion >>
rect 51 30 52 31 
<< pdiffusion >>
rect 52 30 53 31 
<< pdiffusion >>
rect 53 30 54 31 
<< m1 >>
rect 64 30 65 31 
<< pdiffusion >>
rect 66 30 67 31 
<< m1 >>
rect 67 30 68 31 
<< pdiffusion >>
rect 67 30 68 31 
<< pdiffusion >>
rect 68 30 69 31 
<< pdiffusion >>
rect 69 30 70 31 
<< pdiffusion >>
rect 70 30 71 31 
<< pdiffusion >>
rect 71 30 72 31 
<< pdiffusion >>
rect 84 30 85 31 
<< pdiffusion >>
rect 85 30 86 31 
<< pdiffusion >>
rect 86 30 87 31 
<< pdiffusion >>
rect 87 30 88 31 
<< pdiffusion >>
rect 88 30 89 31 
<< pdiffusion >>
rect 89 30 90 31 
<< pdiffusion >>
rect 102 30 103 31 
<< pdiffusion >>
rect 103 30 104 31 
<< pdiffusion >>
rect 104 30 105 31 
<< pdiffusion >>
rect 105 30 106 31 
<< m1 >>
rect 106 30 107 31 
<< pdiffusion >>
rect 106 30 107 31 
<< pdiffusion >>
rect 107 30 108 31 
<< m1 >>
rect 111 30 112 31 
<< pdiffusion >>
rect 120 30 121 31 
<< pdiffusion >>
rect 121 30 122 31 
<< pdiffusion >>
rect 122 30 123 31 
<< pdiffusion >>
rect 123 30 124 31 
<< m1 >>
rect 124 30 125 31 
<< pdiffusion >>
rect 124 30 125 31 
<< pdiffusion >>
rect 125 30 126 31 
<< m1 >>
rect 127 30 128 31 
<< pdiffusion >>
rect 138 30 139 31 
<< pdiffusion >>
rect 139 30 140 31 
<< pdiffusion >>
rect 140 30 141 31 
<< pdiffusion >>
rect 141 30 142 31 
<< m1 >>
rect 142 30 143 31 
<< pdiffusion >>
rect 142 30 143 31 
<< pdiffusion >>
rect 143 30 144 31 
<< m1 >>
rect 145 30 146 31 
<< pdiffusion >>
rect 156 30 157 31 
<< pdiffusion >>
rect 157 30 158 31 
<< pdiffusion >>
rect 158 30 159 31 
<< pdiffusion >>
rect 159 30 160 31 
<< pdiffusion >>
rect 160 30 161 31 
<< pdiffusion >>
rect 161 30 162 31 
<< pdiffusion >>
rect 174 30 175 31 
<< pdiffusion >>
rect 175 30 176 31 
<< pdiffusion >>
rect 176 30 177 31 
<< pdiffusion >>
rect 177 30 178 31 
<< pdiffusion >>
rect 178 30 179 31 
<< pdiffusion >>
rect 179 30 180 31 
<< pdiffusion >>
rect 192 30 193 31 
<< m1 >>
rect 193 30 194 31 
<< pdiffusion >>
rect 193 30 194 31 
<< pdiffusion >>
rect 194 30 195 31 
<< pdiffusion >>
rect 195 30 196 31 
<< pdiffusion >>
rect 196 30 197 31 
<< pdiffusion >>
rect 197 30 198 31 
<< m1 >>
rect 208 30 209 31 
<< pdiffusion >>
rect 210 30 211 31 
<< pdiffusion >>
rect 211 30 212 31 
<< pdiffusion >>
rect 212 30 213 31 
<< pdiffusion >>
rect 213 30 214 31 
<< pdiffusion >>
rect 214 30 215 31 
<< pdiffusion >>
rect 215 30 216 31 
<< m2 >>
rect 225 30 226 31 
<< m1 >>
rect 226 30 227 31 
<< pdiffusion >>
rect 228 30 229 31 
<< pdiffusion >>
rect 229 30 230 31 
<< pdiffusion >>
rect 230 30 231 31 
<< pdiffusion >>
rect 231 30 232 31 
<< pdiffusion >>
rect 232 30 233 31 
<< pdiffusion >>
rect 233 30 234 31 
<< m1 >>
rect 235 30 236 31 
<< pdiffusion >>
rect 264 30 265 31 
<< pdiffusion >>
rect 265 30 266 31 
<< pdiffusion >>
rect 266 30 267 31 
<< pdiffusion >>
rect 267 30 268 31 
<< pdiffusion >>
rect 268 30 269 31 
<< pdiffusion >>
rect 269 30 270 31 
<< m1 >>
rect 278 30 279 31 
<< m1 >>
rect 280 30 281 31 
<< pdiffusion >>
rect 282 30 283 31 
<< pdiffusion >>
rect 283 30 284 31 
<< pdiffusion >>
rect 284 30 285 31 
<< pdiffusion >>
rect 285 30 286 31 
<< m1 >>
rect 286 30 287 31 
<< pdiffusion >>
rect 286 30 287 31 
<< pdiffusion >>
rect 287 30 288 31 
<< pdiffusion >>
rect 300 30 301 31 
<< pdiffusion >>
rect 301 30 302 31 
<< pdiffusion >>
rect 302 30 303 31 
<< pdiffusion >>
rect 303 30 304 31 
<< pdiffusion >>
rect 304 30 305 31 
<< pdiffusion >>
rect 305 30 306 31 
<< pdiffusion >>
rect 318 30 319 31 
<< pdiffusion >>
rect 319 30 320 31 
<< pdiffusion >>
rect 320 30 321 31 
<< pdiffusion >>
rect 321 30 322 31 
<< pdiffusion >>
rect 322 30 323 31 
<< pdiffusion >>
rect 323 30 324 31 
<< m1 >>
rect 334 30 335 31 
<< pdiffusion >>
rect 336 30 337 31 
<< pdiffusion >>
rect 337 30 338 31 
<< pdiffusion >>
rect 338 30 339 31 
<< pdiffusion >>
rect 339 30 340 31 
<< pdiffusion >>
rect 340 30 341 31 
<< pdiffusion >>
rect 341 30 342 31 
<< pdiffusion >>
rect 354 30 355 31 
<< pdiffusion >>
rect 355 30 356 31 
<< pdiffusion >>
rect 356 30 357 31 
<< pdiffusion >>
rect 357 30 358 31 
<< pdiffusion >>
rect 358 30 359 31 
<< pdiffusion >>
rect 359 30 360 31 
<< pdiffusion >>
rect 372 30 373 31 
<< pdiffusion >>
rect 373 30 374 31 
<< pdiffusion >>
rect 374 30 375 31 
<< pdiffusion >>
rect 375 30 376 31 
<< pdiffusion >>
rect 376 30 377 31 
<< pdiffusion >>
rect 377 30 378 31 
<< m1 >>
rect 388 30 389 31 
<< pdiffusion >>
rect 390 30 391 31 
<< pdiffusion >>
rect 391 30 392 31 
<< pdiffusion >>
rect 392 30 393 31 
<< pdiffusion >>
rect 393 30 394 31 
<< pdiffusion >>
rect 394 30 395 31 
<< pdiffusion >>
rect 395 30 396 31 
<< m1 >>
rect 406 30 407 31 
<< pdiffusion >>
rect 408 30 409 31 
<< m1 >>
rect 409 30 410 31 
<< pdiffusion >>
rect 409 30 410 31 
<< pdiffusion >>
rect 410 30 411 31 
<< pdiffusion >>
rect 411 30 412 31 
<< pdiffusion >>
rect 412 30 413 31 
<< pdiffusion >>
rect 413 30 414 31 
<< pdiffusion >>
rect 426 30 427 31 
<< pdiffusion >>
rect 427 30 428 31 
<< pdiffusion >>
rect 428 30 429 31 
<< pdiffusion >>
rect 429 30 430 31 
<< m1 >>
rect 430 30 431 31 
<< pdiffusion >>
rect 430 30 431 31 
<< pdiffusion >>
rect 431 30 432 31 
<< m1 >>
rect 433 30 434 31 
<< pdiffusion >>
rect 444 30 445 31 
<< pdiffusion >>
rect 445 30 446 31 
<< pdiffusion >>
rect 446 30 447 31 
<< pdiffusion >>
rect 447 30 448 31 
<< m1 >>
rect 448 30 449 31 
<< pdiffusion >>
rect 448 30 449 31 
<< pdiffusion >>
rect 449 30 450 31 
<< pdiffusion >>
rect 462 30 463 31 
<< pdiffusion >>
rect 463 30 464 31 
<< pdiffusion >>
rect 464 30 465 31 
<< pdiffusion >>
rect 465 30 466 31 
<< pdiffusion >>
rect 466 30 467 31 
<< pdiffusion >>
rect 467 30 468 31 
<< pdiffusion >>
rect 480 30 481 31 
<< pdiffusion >>
rect 481 30 482 31 
<< pdiffusion >>
rect 482 30 483 31 
<< pdiffusion >>
rect 483 30 484 31 
<< pdiffusion >>
rect 484 30 485 31 
<< pdiffusion >>
rect 485 30 486 31 
<< m1 >>
rect 487 30 488 31 
<< m1 >>
rect 505 30 506 31 
<< pdiffusion >>
rect 516 30 517 31 
<< pdiffusion >>
rect 517 30 518 31 
<< pdiffusion >>
rect 518 30 519 31 
<< pdiffusion >>
rect 519 30 520 31 
<< m1 >>
rect 520 30 521 31 
<< pdiffusion >>
rect 520 30 521 31 
<< pdiffusion >>
rect 521 30 522 31 
<< pdiffusion >>
rect 12 31 13 32 
<< pdiffusion >>
rect 13 31 14 32 
<< pdiffusion >>
rect 14 31 15 32 
<< pdiffusion >>
rect 15 31 16 32 
<< pdiffusion >>
rect 16 31 17 32 
<< pdiffusion >>
rect 17 31 18 32 
<< pdiffusion >>
rect 30 31 31 32 
<< pdiffusion >>
rect 31 31 32 32 
<< pdiffusion >>
rect 32 31 33 32 
<< pdiffusion >>
rect 33 31 34 32 
<< pdiffusion >>
rect 34 31 35 32 
<< pdiffusion >>
rect 35 31 36 32 
<< pdiffusion >>
rect 48 31 49 32 
<< pdiffusion >>
rect 49 31 50 32 
<< pdiffusion >>
rect 50 31 51 32 
<< pdiffusion >>
rect 51 31 52 32 
<< pdiffusion >>
rect 52 31 53 32 
<< pdiffusion >>
rect 53 31 54 32 
<< m1 >>
rect 64 31 65 32 
<< pdiffusion >>
rect 66 31 67 32 
<< pdiffusion >>
rect 67 31 68 32 
<< pdiffusion >>
rect 68 31 69 32 
<< pdiffusion >>
rect 69 31 70 32 
<< pdiffusion >>
rect 70 31 71 32 
<< pdiffusion >>
rect 71 31 72 32 
<< pdiffusion >>
rect 84 31 85 32 
<< pdiffusion >>
rect 85 31 86 32 
<< pdiffusion >>
rect 86 31 87 32 
<< pdiffusion >>
rect 87 31 88 32 
<< pdiffusion >>
rect 88 31 89 32 
<< pdiffusion >>
rect 89 31 90 32 
<< pdiffusion >>
rect 102 31 103 32 
<< pdiffusion >>
rect 103 31 104 32 
<< pdiffusion >>
rect 104 31 105 32 
<< pdiffusion >>
rect 105 31 106 32 
<< pdiffusion >>
rect 106 31 107 32 
<< pdiffusion >>
rect 107 31 108 32 
<< m1 >>
rect 111 31 112 32 
<< pdiffusion >>
rect 120 31 121 32 
<< pdiffusion >>
rect 121 31 122 32 
<< pdiffusion >>
rect 122 31 123 32 
<< pdiffusion >>
rect 123 31 124 32 
<< pdiffusion >>
rect 124 31 125 32 
<< pdiffusion >>
rect 125 31 126 32 
<< m1 >>
rect 127 31 128 32 
<< pdiffusion >>
rect 138 31 139 32 
<< pdiffusion >>
rect 139 31 140 32 
<< pdiffusion >>
rect 140 31 141 32 
<< pdiffusion >>
rect 141 31 142 32 
<< pdiffusion >>
rect 142 31 143 32 
<< pdiffusion >>
rect 143 31 144 32 
<< m1 >>
rect 145 31 146 32 
<< pdiffusion >>
rect 156 31 157 32 
<< pdiffusion >>
rect 157 31 158 32 
<< pdiffusion >>
rect 158 31 159 32 
<< pdiffusion >>
rect 159 31 160 32 
<< pdiffusion >>
rect 160 31 161 32 
<< pdiffusion >>
rect 161 31 162 32 
<< pdiffusion >>
rect 174 31 175 32 
<< pdiffusion >>
rect 175 31 176 32 
<< pdiffusion >>
rect 176 31 177 32 
<< pdiffusion >>
rect 177 31 178 32 
<< pdiffusion >>
rect 178 31 179 32 
<< pdiffusion >>
rect 179 31 180 32 
<< pdiffusion >>
rect 192 31 193 32 
<< pdiffusion >>
rect 193 31 194 32 
<< pdiffusion >>
rect 194 31 195 32 
<< pdiffusion >>
rect 195 31 196 32 
<< pdiffusion >>
rect 196 31 197 32 
<< pdiffusion >>
rect 197 31 198 32 
<< m1 >>
rect 208 31 209 32 
<< pdiffusion >>
rect 210 31 211 32 
<< pdiffusion >>
rect 211 31 212 32 
<< pdiffusion >>
rect 212 31 213 32 
<< pdiffusion >>
rect 213 31 214 32 
<< pdiffusion >>
rect 214 31 215 32 
<< pdiffusion >>
rect 215 31 216 32 
<< m2 >>
rect 225 31 226 32 
<< m1 >>
rect 226 31 227 32 
<< pdiffusion >>
rect 228 31 229 32 
<< pdiffusion >>
rect 229 31 230 32 
<< pdiffusion >>
rect 230 31 231 32 
<< pdiffusion >>
rect 231 31 232 32 
<< pdiffusion >>
rect 232 31 233 32 
<< pdiffusion >>
rect 233 31 234 32 
<< m1 >>
rect 235 31 236 32 
<< pdiffusion >>
rect 264 31 265 32 
<< pdiffusion >>
rect 265 31 266 32 
<< pdiffusion >>
rect 266 31 267 32 
<< pdiffusion >>
rect 267 31 268 32 
<< pdiffusion >>
rect 268 31 269 32 
<< pdiffusion >>
rect 269 31 270 32 
<< m1 >>
rect 278 31 279 32 
<< m1 >>
rect 280 31 281 32 
<< pdiffusion >>
rect 282 31 283 32 
<< pdiffusion >>
rect 283 31 284 32 
<< pdiffusion >>
rect 284 31 285 32 
<< pdiffusion >>
rect 285 31 286 32 
<< pdiffusion >>
rect 286 31 287 32 
<< pdiffusion >>
rect 287 31 288 32 
<< pdiffusion >>
rect 300 31 301 32 
<< pdiffusion >>
rect 301 31 302 32 
<< pdiffusion >>
rect 302 31 303 32 
<< pdiffusion >>
rect 303 31 304 32 
<< pdiffusion >>
rect 304 31 305 32 
<< pdiffusion >>
rect 305 31 306 32 
<< pdiffusion >>
rect 318 31 319 32 
<< pdiffusion >>
rect 319 31 320 32 
<< pdiffusion >>
rect 320 31 321 32 
<< pdiffusion >>
rect 321 31 322 32 
<< pdiffusion >>
rect 322 31 323 32 
<< pdiffusion >>
rect 323 31 324 32 
<< m1 >>
rect 334 31 335 32 
<< pdiffusion >>
rect 336 31 337 32 
<< pdiffusion >>
rect 337 31 338 32 
<< pdiffusion >>
rect 338 31 339 32 
<< pdiffusion >>
rect 339 31 340 32 
<< pdiffusion >>
rect 340 31 341 32 
<< pdiffusion >>
rect 341 31 342 32 
<< pdiffusion >>
rect 354 31 355 32 
<< pdiffusion >>
rect 355 31 356 32 
<< pdiffusion >>
rect 356 31 357 32 
<< pdiffusion >>
rect 357 31 358 32 
<< pdiffusion >>
rect 358 31 359 32 
<< pdiffusion >>
rect 359 31 360 32 
<< pdiffusion >>
rect 372 31 373 32 
<< pdiffusion >>
rect 373 31 374 32 
<< pdiffusion >>
rect 374 31 375 32 
<< pdiffusion >>
rect 375 31 376 32 
<< pdiffusion >>
rect 376 31 377 32 
<< pdiffusion >>
rect 377 31 378 32 
<< m1 >>
rect 388 31 389 32 
<< pdiffusion >>
rect 390 31 391 32 
<< pdiffusion >>
rect 391 31 392 32 
<< pdiffusion >>
rect 392 31 393 32 
<< pdiffusion >>
rect 393 31 394 32 
<< pdiffusion >>
rect 394 31 395 32 
<< pdiffusion >>
rect 395 31 396 32 
<< m1 >>
rect 406 31 407 32 
<< pdiffusion >>
rect 408 31 409 32 
<< pdiffusion >>
rect 409 31 410 32 
<< pdiffusion >>
rect 410 31 411 32 
<< pdiffusion >>
rect 411 31 412 32 
<< pdiffusion >>
rect 412 31 413 32 
<< pdiffusion >>
rect 413 31 414 32 
<< pdiffusion >>
rect 426 31 427 32 
<< pdiffusion >>
rect 427 31 428 32 
<< pdiffusion >>
rect 428 31 429 32 
<< pdiffusion >>
rect 429 31 430 32 
<< pdiffusion >>
rect 430 31 431 32 
<< pdiffusion >>
rect 431 31 432 32 
<< m1 >>
rect 433 31 434 32 
<< pdiffusion >>
rect 444 31 445 32 
<< pdiffusion >>
rect 445 31 446 32 
<< pdiffusion >>
rect 446 31 447 32 
<< pdiffusion >>
rect 447 31 448 32 
<< pdiffusion >>
rect 448 31 449 32 
<< pdiffusion >>
rect 449 31 450 32 
<< pdiffusion >>
rect 462 31 463 32 
<< pdiffusion >>
rect 463 31 464 32 
<< pdiffusion >>
rect 464 31 465 32 
<< pdiffusion >>
rect 465 31 466 32 
<< pdiffusion >>
rect 466 31 467 32 
<< pdiffusion >>
rect 467 31 468 32 
<< pdiffusion >>
rect 480 31 481 32 
<< pdiffusion >>
rect 481 31 482 32 
<< pdiffusion >>
rect 482 31 483 32 
<< pdiffusion >>
rect 483 31 484 32 
<< pdiffusion >>
rect 484 31 485 32 
<< pdiffusion >>
rect 485 31 486 32 
<< m1 >>
rect 487 31 488 32 
<< m1 >>
rect 505 31 506 32 
<< pdiffusion >>
rect 516 31 517 32 
<< pdiffusion >>
rect 517 31 518 32 
<< pdiffusion >>
rect 518 31 519 32 
<< pdiffusion >>
rect 519 31 520 32 
<< pdiffusion >>
rect 520 31 521 32 
<< pdiffusion >>
rect 521 31 522 32 
<< pdiffusion >>
rect 12 32 13 33 
<< pdiffusion >>
rect 13 32 14 33 
<< pdiffusion >>
rect 14 32 15 33 
<< pdiffusion >>
rect 15 32 16 33 
<< pdiffusion >>
rect 16 32 17 33 
<< pdiffusion >>
rect 17 32 18 33 
<< pdiffusion >>
rect 30 32 31 33 
<< pdiffusion >>
rect 31 32 32 33 
<< pdiffusion >>
rect 32 32 33 33 
<< pdiffusion >>
rect 33 32 34 33 
<< pdiffusion >>
rect 34 32 35 33 
<< pdiffusion >>
rect 35 32 36 33 
<< pdiffusion >>
rect 48 32 49 33 
<< pdiffusion >>
rect 49 32 50 33 
<< pdiffusion >>
rect 50 32 51 33 
<< pdiffusion >>
rect 51 32 52 33 
<< pdiffusion >>
rect 52 32 53 33 
<< pdiffusion >>
rect 53 32 54 33 
<< m1 >>
rect 64 32 65 33 
<< pdiffusion >>
rect 66 32 67 33 
<< pdiffusion >>
rect 67 32 68 33 
<< pdiffusion >>
rect 68 32 69 33 
<< pdiffusion >>
rect 69 32 70 33 
<< pdiffusion >>
rect 70 32 71 33 
<< pdiffusion >>
rect 71 32 72 33 
<< pdiffusion >>
rect 84 32 85 33 
<< pdiffusion >>
rect 85 32 86 33 
<< pdiffusion >>
rect 86 32 87 33 
<< pdiffusion >>
rect 87 32 88 33 
<< pdiffusion >>
rect 88 32 89 33 
<< pdiffusion >>
rect 89 32 90 33 
<< pdiffusion >>
rect 102 32 103 33 
<< pdiffusion >>
rect 103 32 104 33 
<< pdiffusion >>
rect 104 32 105 33 
<< pdiffusion >>
rect 105 32 106 33 
<< pdiffusion >>
rect 106 32 107 33 
<< pdiffusion >>
rect 107 32 108 33 
<< m1 >>
rect 111 32 112 33 
<< pdiffusion >>
rect 120 32 121 33 
<< pdiffusion >>
rect 121 32 122 33 
<< pdiffusion >>
rect 122 32 123 33 
<< pdiffusion >>
rect 123 32 124 33 
<< pdiffusion >>
rect 124 32 125 33 
<< pdiffusion >>
rect 125 32 126 33 
<< m1 >>
rect 127 32 128 33 
<< pdiffusion >>
rect 138 32 139 33 
<< pdiffusion >>
rect 139 32 140 33 
<< pdiffusion >>
rect 140 32 141 33 
<< pdiffusion >>
rect 141 32 142 33 
<< pdiffusion >>
rect 142 32 143 33 
<< pdiffusion >>
rect 143 32 144 33 
<< m1 >>
rect 145 32 146 33 
<< pdiffusion >>
rect 156 32 157 33 
<< pdiffusion >>
rect 157 32 158 33 
<< pdiffusion >>
rect 158 32 159 33 
<< pdiffusion >>
rect 159 32 160 33 
<< pdiffusion >>
rect 160 32 161 33 
<< pdiffusion >>
rect 161 32 162 33 
<< pdiffusion >>
rect 174 32 175 33 
<< pdiffusion >>
rect 175 32 176 33 
<< pdiffusion >>
rect 176 32 177 33 
<< pdiffusion >>
rect 177 32 178 33 
<< pdiffusion >>
rect 178 32 179 33 
<< pdiffusion >>
rect 179 32 180 33 
<< pdiffusion >>
rect 192 32 193 33 
<< pdiffusion >>
rect 193 32 194 33 
<< pdiffusion >>
rect 194 32 195 33 
<< pdiffusion >>
rect 195 32 196 33 
<< pdiffusion >>
rect 196 32 197 33 
<< pdiffusion >>
rect 197 32 198 33 
<< m1 >>
rect 208 32 209 33 
<< pdiffusion >>
rect 210 32 211 33 
<< pdiffusion >>
rect 211 32 212 33 
<< pdiffusion >>
rect 212 32 213 33 
<< pdiffusion >>
rect 213 32 214 33 
<< pdiffusion >>
rect 214 32 215 33 
<< pdiffusion >>
rect 215 32 216 33 
<< m2 >>
rect 225 32 226 33 
<< m1 >>
rect 226 32 227 33 
<< pdiffusion >>
rect 228 32 229 33 
<< pdiffusion >>
rect 229 32 230 33 
<< pdiffusion >>
rect 230 32 231 33 
<< pdiffusion >>
rect 231 32 232 33 
<< pdiffusion >>
rect 232 32 233 33 
<< pdiffusion >>
rect 233 32 234 33 
<< m1 >>
rect 235 32 236 33 
<< pdiffusion >>
rect 264 32 265 33 
<< pdiffusion >>
rect 265 32 266 33 
<< pdiffusion >>
rect 266 32 267 33 
<< pdiffusion >>
rect 267 32 268 33 
<< pdiffusion >>
rect 268 32 269 33 
<< pdiffusion >>
rect 269 32 270 33 
<< m1 >>
rect 278 32 279 33 
<< m1 >>
rect 280 32 281 33 
<< pdiffusion >>
rect 282 32 283 33 
<< pdiffusion >>
rect 283 32 284 33 
<< pdiffusion >>
rect 284 32 285 33 
<< pdiffusion >>
rect 285 32 286 33 
<< pdiffusion >>
rect 286 32 287 33 
<< pdiffusion >>
rect 287 32 288 33 
<< pdiffusion >>
rect 300 32 301 33 
<< pdiffusion >>
rect 301 32 302 33 
<< pdiffusion >>
rect 302 32 303 33 
<< pdiffusion >>
rect 303 32 304 33 
<< pdiffusion >>
rect 304 32 305 33 
<< pdiffusion >>
rect 305 32 306 33 
<< pdiffusion >>
rect 318 32 319 33 
<< pdiffusion >>
rect 319 32 320 33 
<< pdiffusion >>
rect 320 32 321 33 
<< pdiffusion >>
rect 321 32 322 33 
<< pdiffusion >>
rect 322 32 323 33 
<< pdiffusion >>
rect 323 32 324 33 
<< m1 >>
rect 334 32 335 33 
<< pdiffusion >>
rect 336 32 337 33 
<< pdiffusion >>
rect 337 32 338 33 
<< pdiffusion >>
rect 338 32 339 33 
<< pdiffusion >>
rect 339 32 340 33 
<< pdiffusion >>
rect 340 32 341 33 
<< pdiffusion >>
rect 341 32 342 33 
<< pdiffusion >>
rect 354 32 355 33 
<< pdiffusion >>
rect 355 32 356 33 
<< pdiffusion >>
rect 356 32 357 33 
<< pdiffusion >>
rect 357 32 358 33 
<< pdiffusion >>
rect 358 32 359 33 
<< pdiffusion >>
rect 359 32 360 33 
<< pdiffusion >>
rect 372 32 373 33 
<< pdiffusion >>
rect 373 32 374 33 
<< pdiffusion >>
rect 374 32 375 33 
<< pdiffusion >>
rect 375 32 376 33 
<< pdiffusion >>
rect 376 32 377 33 
<< pdiffusion >>
rect 377 32 378 33 
<< m1 >>
rect 388 32 389 33 
<< pdiffusion >>
rect 390 32 391 33 
<< pdiffusion >>
rect 391 32 392 33 
<< pdiffusion >>
rect 392 32 393 33 
<< pdiffusion >>
rect 393 32 394 33 
<< pdiffusion >>
rect 394 32 395 33 
<< pdiffusion >>
rect 395 32 396 33 
<< m1 >>
rect 406 32 407 33 
<< pdiffusion >>
rect 408 32 409 33 
<< pdiffusion >>
rect 409 32 410 33 
<< pdiffusion >>
rect 410 32 411 33 
<< pdiffusion >>
rect 411 32 412 33 
<< pdiffusion >>
rect 412 32 413 33 
<< pdiffusion >>
rect 413 32 414 33 
<< pdiffusion >>
rect 426 32 427 33 
<< pdiffusion >>
rect 427 32 428 33 
<< pdiffusion >>
rect 428 32 429 33 
<< pdiffusion >>
rect 429 32 430 33 
<< pdiffusion >>
rect 430 32 431 33 
<< pdiffusion >>
rect 431 32 432 33 
<< m1 >>
rect 433 32 434 33 
<< pdiffusion >>
rect 444 32 445 33 
<< pdiffusion >>
rect 445 32 446 33 
<< pdiffusion >>
rect 446 32 447 33 
<< pdiffusion >>
rect 447 32 448 33 
<< pdiffusion >>
rect 448 32 449 33 
<< pdiffusion >>
rect 449 32 450 33 
<< pdiffusion >>
rect 462 32 463 33 
<< pdiffusion >>
rect 463 32 464 33 
<< pdiffusion >>
rect 464 32 465 33 
<< pdiffusion >>
rect 465 32 466 33 
<< pdiffusion >>
rect 466 32 467 33 
<< pdiffusion >>
rect 467 32 468 33 
<< pdiffusion >>
rect 480 32 481 33 
<< pdiffusion >>
rect 481 32 482 33 
<< pdiffusion >>
rect 482 32 483 33 
<< pdiffusion >>
rect 483 32 484 33 
<< pdiffusion >>
rect 484 32 485 33 
<< pdiffusion >>
rect 485 32 486 33 
<< m1 >>
rect 487 32 488 33 
<< m1 >>
rect 505 32 506 33 
<< pdiffusion >>
rect 516 32 517 33 
<< pdiffusion >>
rect 517 32 518 33 
<< pdiffusion >>
rect 518 32 519 33 
<< pdiffusion >>
rect 519 32 520 33 
<< pdiffusion >>
rect 520 32 521 33 
<< pdiffusion >>
rect 521 32 522 33 
<< pdiffusion >>
rect 12 33 13 34 
<< pdiffusion >>
rect 13 33 14 34 
<< pdiffusion >>
rect 14 33 15 34 
<< pdiffusion >>
rect 15 33 16 34 
<< pdiffusion >>
rect 16 33 17 34 
<< pdiffusion >>
rect 17 33 18 34 
<< pdiffusion >>
rect 30 33 31 34 
<< pdiffusion >>
rect 31 33 32 34 
<< pdiffusion >>
rect 32 33 33 34 
<< pdiffusion >>
rect 33 33 34 34 
<< pdiffusion >>
rect 34 33 35 34 
<< pdiffusion >>
rect 35 33 36 34 
<< pdiffusion >>
rect 48 33 49 34 
<< pdiffusion >>
rect 49 33 50 34 
<< pdiffusion >>
rect 50 33 51 34 
<< pdiffusion >>
rect 51 33 52 34 
<< pdiffusion >>
rect 52 33 53 34 
<< pdiffusion >>
rect 53 33 54 34 
<< m1 >>
rect 64 33 65 34 
<< pdiffusion >>
rect 66 33 67 34 
<< pdiffusion >>
rect 67 33 68 34 
<< pdiffusion >>
rect 68 33 69 34 
<< pdiffusion >>
rect 69 33 70 34 
<< pdiffusion >>
rect 70 33 71 34 
<< pdiffusion >>
rect 71 33 72 34 
<< pdiffusion >>
rect 84 33 85 34 
<< pdiffusion >>
rect 85 33 86 34 
<< pdiffusion >>
rect 86 33 87 34 
<< pdiffusion >>
rect 87 33 88 34 
<< pdiffusion >>
rect 88 33 89 34 
<< pdiffusion >>
rect 89 33 90 34 
<< pdiffusion >>
rect 102 33 103 34 
<< pdiffusion >>
rect 103 33 104 34 
<< pdiffusion >>
rect 104 33 105 34 
<< pdiffusion >>
rect 105 33 106 34 
<< pdiffusion >>
rect 106 33 107 34 
<< pdiffusion >>
rect 107 33 108 34 
<< m1 >>
rect 111 33 112 34 
<< pdiffusion >>
rect 120 33 121 34 
<< pdiffusion >>
rect 121 33 122 34 
<< pdiffusion >>
rect 122 33 123 34 
<< pdiffusion >>
rect 123 33 124 34 
<< pdiffusion >>
rect 124 33 125 34 
<< pdiffusion >>
rect 125 33 126 34 
<< m1 >>
rect 127 33 128 34 
<< pdiffusion >>
rect 138 33 139 34 
<< pdiffusion >>
rect 139 33 140 34 
<< pdiffusion >>
rect 140 33 141 34 
<< pdiffusion >>
rect 141 33 142 34 
<< pdiffusion >>
rect 142 33 143 34 
<< pdiffusion >>
rect 143 33 144 34 
<< m1 >>
rect 145 33 146 34 
<< pdiffusion >>
rect 156 33 157 34 
<< pdiffusion >>
rect 157 33 158 34 
<< pdiffusion >>
rect 158 33 159 34 
<< pdiffusion >>
rect 159 33 160 34 
<< pdiffusion >>
rect 160 33 161 34 
<< pdiffusion >>
rect 161 33 162 34 
<< pdiffusion >>
rect 174 33 175 34 
<< pdiffusion >>
rect 175 33 176 34 
<< pdiffusion >>
rect 176 33 177 34 
<< pdiffusion >>
rect 177 33 178 34 
<< pdiffusion >>
rect 178 33 179 34 
<< pdiffusion >>
rect 179 33 180 34 
<< pdiffusion >>
rect 192 33 193 34 
<< pdiffusion >>
rect 193 33 194 34 
<< pdiffusion >>
rect 194 33 195 34 
<< pdiffusion >>
rect 195 33 196 34 
<< pdiffusion >>
rect 196 33 197 34 
<< pdiffusion >>
rect 197 33 198 34 
<< m1 >>
rect 208 33 209 34 
<< pdiffusion >>
rect 210 33 211 34 
<< pdiffusion >>
rect 211 33 212 34 
<< pdiffusion >>
rect 212 33 213 34 
<< pdiffusion >>
rect 213 33 214 34 
<< pdiffusion >>
rect 214 33 215 34 
<< pdiffusion >>
rect 215 33 216 34 
<< m2 >>
rect 225 33 226 34 
<< m1 >>
rect 226 33 227 34 
<< pdiffusion >>
rect 228 33 229 34 
<< pdiffusion >>
rect 229 33 230 34 
<< pdiffusion >>
rect 230 33 231 34 
<< pdiffusion >>
rect 231 33 232 34 
<< pdiffusion >>
rect 232 33 233 34 
<< pdiffusion >>
rect 233 33 234 34 
<< m1 >>
rect 235 33 236 34 
<< pdiffusion >>
rect 264 33 265 34 
<< pdiffusion >>
rect 265 33 266 34 
<< pdiffusion >>
rect 266 33 267 34 
<< pdiffusion >>
rect 267 33 268 34 
<< pdiffusion >>
rect 268 33 269 34 
<< pdiffusion >>
rect 269 33 270 34 
<< m1 >>
rect 278 33 279 34 
<< m1 >>
rect 280 33 281 34 
<< pdiffusion >>
rect 282 33 283 34 
<< pdiffusion >>
rect 283 33 284 34 
<< pdiffusion >>
rect 284 33 285 34 
<< pdiffusion >>
rect 285 33 286 34 
<< pdiffusion >>
rect 286 33 287 34 
<< pdiffusion >>
rect 287 33 288 34 
<< pdiffusion >>
rect 300 33 301 34 
<< pdiffusion >>
rect 301 33 302 34 
<< pdiffusion >>
rect 302 33 303 34 
<< pdiffusion >>
rect 303 33 304 34 
<< pdiffusion >>
rect 304 33 305 34 
<< pdiffusion >>
rect 305 33 306 34 
<< pdiffusion >>
rect 318 33 319 34 
<< pdiffusion >>
rect 319 33 320 34 
<< pdiffusion >>
rect 320 33 321 34 
<< pdiffusion >>
rect 321 33 322 34 
<< pdiffusion >>
rect 322 33 323 34 
<< pdiffusion >>
rect 323 33 324 34 
<< m1 >>
rect 334 33 335 34 
<< pdiffusion >>
rect 336 33 337 34 
<< pdiffusion >>
rect 337 33 338 34 
<< pdiffusion >>
rect 338 33 339 34 
<< pdiffusion >>
rect 339 33 340 34 
<< pdiffusion >>
rect 340 33 341 34 
<< pdiffusion >>
rect 341 33 342 34 
<< pdiffusion >>
rect 354 33 355 34 
<< pdiffusion >>
rect 355 33 356 34 
<< pdiffusion >>
rect 356 33 357 34 
<< pdiffusion >>
rect 357 33 358 34 
<< pdiffusion >>
rect 358 33 359 34 
<< pdiffusion >>
rect 359 33 360 34 
<< pdiffusion >>
rect 372 33 373 34 
<< pdiffusion >>
rect 373 33 374 34 
<< pdiffusion >>
rect 374 33 375 34 
<< pdiffusion >>
rect 375 33 376 34 
<< pdiffusion >>
rect 376 33 377 34 
<< pdiffusion >>
rect 377 33 378 34 
<< m1 >>
rect 388 33 389 34 
<< pdiffusion >>
rect 390 33 391 34 
<< pdiffusion >>
rect 391 33 392 34 
<< pdiffusion >>
rect 392 33 393 34 
<< pdiffusion >>
rect 393 33 394 34 
<< pdiffusion >>
rect 394 33 395 34 
<< pdiffusion >>
rect 395 33 396 34 
<< m1 >>
rect 406 33 407 34 
<< pdiffusion >>
rect 408 33 409 34 
<< pdiffusion >>
rect 409 33 410 34 
<< pdiffusion >>
rect 410 33 411 34 
<< pdiffusion >>
rect 411 33 412 34 
<< pdiffusion >>
rect 412 33 413 34 
<< pdiffusion >>
rect 413 33 414 34 
<< pdiffusion >>
rect 426 33 427 34 
<< pdiffusion >>
rect 427 33 428 34 
<< pdiffusion >>
rect 428 33 429 34 
<< pdiffusion >>
rect 429 33 430 34 
<< pdiffusion >>
rect 430 33 431 34 
<< pdiffusion >>
rect 431 33 432 34 
<< m1 >>
rect 433 33 434 34 
<< pdiffusion >>
rect 444 33 445 34 
<< pdiffusion >>
rect 445 33 446 34 
<< pdiffusion >>
rect 446 33 447 34 
<< pdiffusion >>
rect 447 33 448 34 
<< pdiffusion >>
rect 448 33 449 34 
<< pdiffusion >>
rect 449 33 450 34 
<< pdiffusion >>
rect 462 33 463 34 
<< pdiffusion >>
rect 463 33 464 34 
<< pdiffusion >>
rect 464 33 465 34 
<< pdiffusion >>
rect 465 33 466 34 
<< pdiffusion >>
rect 466 33 467 34 
<< pdiffusion >>
rect 467 33 468 34 
<< pdiffusion >>
rect 480 33 481 34 
<< pdiffusion >>
rect 481 33 482 34 
<< pdiffusion >>
rect 482 33 483 34 
<< pdiffusion >>
rect 483 33 484 34 
<< pdiffusion >>
rect 484 33 485 34 
<< pdiffusion >>
rect 485 33 486 34 
<< m1 >>
rect 487 33 488 34 
<< m1 >>
rect 505 33 506 34 
<< pdiffusion >>
rect 516 33 517 34 
<< pdiffusion >>
rect 517 33 518 34 
<< pdiffusion >>
rect 518 33 519 34 
<< pdiffusion >>
rect 519 33 520 34 
<< pdiffusion >>
rect 520 33 521 34 
<< pdiffusion >>
rect 521 33 522 34 
<< pdiffusion >>
rect 12 34 13 35 
<< pdiffusion >>
rect 13 34 14 35 
<< pdiffusion >>
rect 14 34 15 35 
<< pdiffusion >>
rect 15 34 16 35 
<< pdiffusion >>
rect 16 34 17 35 
<< pdiffusion >>
rect 17 34 18 35 
<< pdiffusion >>
rect 30 34 31 35 
<< pdiffusion >>
rect 31 34 32 35 
<< pdiffusion >>
rect 32 34 33 35 
<< pdiffusion >>
rect 33 34 34 35 
<< pdiffusion >>
rect 34 34 35 35 
<< pdiffusion >>
rect 35 34 36 35 
<< pdiffusion >>
rect 48 34 49 35 
<< pdiffusion >>
rect 49 34 50 35 
<< pdiffusion >>
rect 50 34 51 35 
<< pdiffusion >>
rect 51 34 52 35 
<< pdiffusion >>
rect 52 34 53 35 
<< pdiffusion >>
rect 53 34 54 35 
<< m1 >>
rect 64 34 65 35 
<< pdiffusion >>
rect 66 34 67 35 
<< pdiffusion >>
rect 67 34 68 35 
<< pdiffusion >>
rect 68 34 69 35 
<< pdiffusion >>
rect 69 34 70 35 
<< pdiffusion >>
rect 70 34 71 35 
<< pdiffusion >>
rect 71 34 72 35 
<< pdiffusion >>
rect 84 34 85 35 
<< pdiffusion >>
rect 85 34 86 35 
<< pdiffusion >>
rect 86 34 87 35 
<< pdiffusion >>
rect 87 34 88 35 
<< pdiffusion >>
rect 88 34 89 35 
<< pdiffusion >>
rect 89 34 90 35 
<< pdiffusion >>
rect 102 34 103 35 
<< pdiffusion >>
rect 103 34 104 35 
<< pdiffusion >>
rect 104 34 105 35 
<< pdiffusion >>
rect 105 34 106 35 
<< pdiffusion >>
rect 106 34 107 35 
<< pdiffusion >>
rect 107 34 108 35 
<< m1 >>
rect 111 34 112 35 
<< pdiffusion >>
rect 120 34 121 35 
<< pdiffusion >>
rect 121 34 122 35 
<< pdiffusion >>
rect 122 34 123 35 
<< pdiffusion >>
rect 123 34 124 35 
<< pdiffusion >>
rect 124 34 125 35 
<< pdiffusion >>
rect 125 34 126 35 
<< m1 >>
rect 127 34 128 35 
<< pdiffusion >>
rect 138 34 139 35 
<< pdiffusion >>
rect 139 34 140 35 
<< pdiffusion >>
rect 140 34 141 35 
<< pdiffusion >>
rect 141 34 142 35 
<< pdiffusion >>
rect 142 34 143 35 
<< pdiffusion >>
rect 143 34 144 35 
<< m1 >>
rect 145 34 146 35 
<< pdiffusion >>
rect 156 34 157 35 
<< pdiffusion >>
rect 157 34 158 35 
<< pdiffusion >>
rect 158 34 159 35 
<< pdiffusion >>
rect 159 34 160 35 
<< pdiffusion >>
rect 160 34 161 35 
<< pdiffusion >>
rect 161 34 162 35 
<< pdiffusion >>
rect 174 34 175 35 
<< pdiffusion >>
rect 175 34 176 35 
<< pdiffusion >>
rect 176 34 177 35 
<< pdiffusion >>
rect 177 34 178 35 
<< pdiffusion >>
rect 178 34 179 35 
<< pdiffusion >>
rect 179 34 180 35 
<< pdiffusion >>
rect 192 34 193 35 
<< pdiffusion >>
rect 193 34 194 35 
<< pdiffusion >>
rect 194 34 195 35 
<< pdiffusion >>
rect 195 34 196 35 
<< pdiffusion >>
rect 196 34 197 35 
<< pdiffusion >>
rect 197 34 198 35 
<< m1 >>
rect 208 34 209 35 
<< pdiffusion >>
rect 210 34 211 35 
<< pdiffusion >>
rect 211 34 212 35 
<< pdiffusion >>
rect 212 34 213 35 
<< pdiffusion >>
rect 213 34 214 35 
<< pdiffusion >>
rect 214 34 215 35 
<< pdiffusion >>
rect 215 34 216 35 
<< m2 >>
rect 225 34 226 35 
<< m1 >>
rect 226 34 227 35 
<< pdiffusion >>
rect 228 34 229 35 
<< pdiffusion >>
rect 229 34 230 35 
<< pdiffusion >>
rect 230 34 231 35 
<< pdiffusion >>
rect 231 34 232 35 
<< pdiffusion >>
rect 232 34 233 35 
<< pdiffusion >>
rect 233 34 234 35 
<< m1 >>
rect 235 34 236 35 
<< pdiffusion >>
rect 264 34 265 35 
<< pdiffusion >>
rect 265 34 266 35 
<< pdiffusion >>
rect 266 34 267 35 
<< pdiffusion >>
rect 267 34 268 35 
<< pdiffusion >>
rect 268 34 269 35 
<< pdiffusion >>
rect 269 34 270 35 
<< m1 >>
rect 278 34 279 35 
<< m1 >>
rect 280 34 281 35 
<< pdiffusion >>
rect 282 34 283 35 
<< pdiffusion >>
rect 283 34 284 35 
<< pdiffusion >>
rect 284 34 285 35 
<< pdiffusion >>
rect 285 34 286 35 
<< pdiffusion >>
rect 286 34 287 35 
<< pdiffusion >>
rect 287 34 288 35 
<< pdiffusion >>
rect 300 34 301 35 
<< pdiffusion >>
rect 301 34 302 35 
<< pdiffusion >>
rect 302 34 303 35 
<< pdiffusion >>
rect 303 34 304 35 
<< pdiffusion >>
rect 304 34 305 35 
<< pdiffusion >>
rect 305 34 306 35 
<< pdiffusion >>
rect 318 34 319 35 
<< pdiffusion >>
rect 319 34 320 35 
<< pdiffusion >>
rect 320 34 321 35 
<< pdiffusion >>
rect 321 34 322 35 
<< pdiffusion >>
rect 322 34 323 35 
<< pdiffusion >>
rect 323 34 324 35 
<< m1 >>
rect 334 34 335 35 
<< pdiffusion >>
rect 336 34 337 35 
<< pdiffusion >>
rect 337 34 338 35 
<< pdiffusion >>
rect 338 34 339 35 
<< pdiffusion >>
rect 339 34 340 35 
<< pdiffusion >>
rect 340 34 341 35 
<< pdiffusion >>
rect 341 34 342 35 
<< pdiffusion >>
rect 354 34 355 35 
<< pdiffusion >>
rect 355 34 356 35 
<< pdiffusion >>
rect 356 34 357 35 
<< pdiffusion >>
rect 357 34 358 35 
<< pdiffusion >>
rect 358 34 359 35 
<< pdiffusion >>
rect 359 34 360 35 
<< pdiffusion >>
rect 372 34 373 35 
<< pdiffusion >>
rect 373 34 374 35 
<< pdiffusion >>
rect 374 34 375 35 
<< pdiffusion >>
rect 375 34 376 35 
<< pdiffusion >>
rect 376 34 377 35 
<< pdiffusion >>
rect 377 34 378 35 
<< m1 >>
rect 388 34 389 35 
<< pdiffusion >>
rect 390 34 391 35 
<< pdiffusion >>
rect 391 34 392 35 
<< pdiffusion >>
rect 392 34 393 35 
<< pdiffusion >>
rect 393 34 394 35 
<< pdiffusion >>
rect 394 34 395 35 
<< pdiffusion >>
rect 395 34 396 35 
<< m1 >>
rect 406 34 407 35 
<< pdiffusion >>
rect 408 34 409 35 
<< pdiffusion >>
rect 409 34 410 35 
<< pdiffusion >>
rect 410 34 411 35 
<< pdiffusion >>
rect 411 34 412 35 
<< pdiffusion >>
rect 412 34 413 35 
<< pdiffusion >>
rect 413 34 414 35 
<< pdiffusion >>
rect 426 34 427 35 
<< pdiffusion >>
rect 427 34 428 35 
<< pdiffusion >>
rect 428 34 429 35 
<< pdiffusion >>
rect 429 34 430 35 
<< pdiffusion >>
rect 430 34 431 35 
<< pdiffusion >>
rect 431 34 432 35 
<< m1 >>
rect 433 34 434 35 
<< pdiffusion >>
rect 444 34 445 35 
<< pdiffusion >>
rect 445 34 446 35 
<< pdiffusion >>
rect 446 34 447 35 
<< pdiffusion >>
rect 447 34 448 35 
<< pdiffusion >>
rect 448 34 449 35 
<< pdiffusion >>
rect 449 34 450 35 
<< pdiffusion >>
rect 462 34 463 35 
<< pdiffusion >>
rect 463 34 464 35 
<< pdiffusion >>
rect 464 34 465 35 
<< pdiffusion >>
rect 465 34 466 35 
<< pdiffusion >>
rect 466 34 467 35 
<< pdiffusion >>
rect 467 34 468 35 
<< pdiffusion >>
rect 480 34 481 35 
<< pdiffusion >>
rect 481 34 482 35 
<< pdiffusion >>
rect 482 34 483 35 
<< pdiffusion >>
rect 483 34 484 35 
<< pdiffusion >>
rect 484 34 485 35 
<< pdiffusion >>
rect 485 34 486 35 
<< m1 >>
rect 487 34 488 35 
<< m1 >>
rect 505 34 506 35 
<< pdiffusion >>
rect 516 34 517 35 
<< pdiffusion >>
rect 517 34 518 35 
<< pdiffusion >>
rect 518 34 519 35 
<< pdiffusion >>
rect 519 34 520 35 
<< pdiffusion >>
rect 520 34 521 35 
<< pdiffusion >>
rect 521 34 522 35 
<< pdiffusion >>
rect 12 35 13 36 
<< pdiffusion >>
rect 13 35 14 36 
<< pdiffusion >>
rect 14 35 15 36 
<< pdiffusion >>
rect 15 35 16 36 
<< pdiffusion >>
rect 16 35 17 36 
<< pdiffusion >>
rect 17 35 18 36 
<< pdiffusion >>
rect 30 35 31 36 
<< pdiffusion >>
rect 31 35 32 36 
<< pdiffusion >>
rect 32 35 33 36 
<< pdiffusion >>
rect 33 35 34 36 
<< pdiffusion >>
rect 34 35 35 36 
<< pdiffusion >>
rect 35 35 36 36 
<< pdiffusion >>
rect 48 35 49 36 
<< pdiffusion >>
rect 49 35 50 36 
<< pdiffusion >>
rect 50 35 51 36 
<< pdiffusion >>
rect 51 35 52 36 
<< pdiffusion >>
rect 52 35 53 36 
<< pdiffusion >>
rect 53 35 54 36 
<< m1 >>
rect 64 35 65 36 
<< pdiffusion >>
rect 66 35 67 36 
<< pdiffusion >>
rect 67 35 68 36 
<< pdiffusion >>
rect 68 35 69 36 
<< pdiffusion >>
rect 69 35 70 36 
<< pdiffusion >>
rect 70 35 71 36 
<< pdiffusion >>
rect 71 35 72 36 
<< pdiffusion >>
rect 84 35 85 36 
<< m1 >>
rect 85 35 86 36 
<< pdiffusion >>
rect 85 35 86 36 
<< pdiffusion >>
rect 86 35 87 36 
<< pdiffusion >>
rect 87 35 88 36 
<< pdiffusion >>
rect 88 35 89 36 
<< pdiffusion >>
rect 89 35 90 36 
<< pdiffusion >>
rect 102 35 103 36 
<< pdiffusion >>
rect 103 35 104 36 
<< pdiffusion >>
rect 104 35 105 36 
<< pdiffusion >>
rect 105 35 106 36 
<< m1 >>
rect 106 35 107 36 
<< pdiffusion >>
rect 106 35 107 36 
<< pdiffusion >>
rect 107 35 108 36 
<< m1 >>
rect 111 35 112 36 
<< pdiffusion >>
rect 120 35 121 36 
<< pdiffusion >>
rect 121 35 122 36 
<< pdiffusion >>
rect 122 35 123 36 
<< pdiffusion >>
rect 123 35 124 36 
<< pdiffusion >>
rect 124 35 125 36 
<< pdiffusion >>
rect 125 35 126 36 
<< m1 >>
rect 127 35 128 36 
<< pdiffusion >>
rect 138 35 139 36 
<< pdiffusion >>
rect 139 35 140 36 
<< pdiffusion >>
rect 140 35 141 36 
<< pdiffusion >>
rect 141 35 142 36 
<< pdiffusion >>
rect 142 35 143 36 
<< pdiffusion >>
rect 143 35 144 36 
<< m1 >>
rect 145 35 146 36 
<< pdiffusion >>
rect 156 35 157 36 
<< m1 >>
rect 157 35 158 36 
<< pdiffusion >>
rect 157 35 158 36 
<< pdiffusion >>
rect 158 35 159 36 
<< pdiffusion >>
rect 159 35 160 36 
<< m1 >>
rect 160 35 161 36 
<< pdiffusion >>
rect 160 35 161 36 
<< pdiffusion >>
rect 161 35 162 36 
<< pdiffusion >>
rect 174 35 175 36 
<< pdiffusion >>
rect 175 35 176 36 
<< pdiffusion >>
rect 176 35 177 36 
<< pdiffusion >>
rect 177 35 178 36 
<< pdiffusion >>
rect 178 35 179 36 
<< pdiffusion >>
rect 179 35 180 36 
<< pdiffusion >>
rect 192 35 193 36 
<< m1 >>
rect 193 35 194 36 
<< pdiffusion >>
rect 193 35 194 36 
<< pdiffusion >>
rect 194 35 195 36 
<< pdiffusion >>
rect 195 35 196 36 
<< pdiffusion >>
rect 196 35 197 36 
<< pdiffusion >>
rect 197 35 198 36 
<< m1 >>
rect 208 35 209 36 
<< pdiffusion >>
rect 210 35 211 36 
<< pdiffusion >>
rect 211 35 212 36 
<< pdiffusion >>
rect 212 35 213 36 
<< pdiffusion >>
rect 213 35 214 36 
<< m1 >>
rect 214 35 215 36 
<< pdiffusion >>
rect 214 35 215 36 
<< pdiffusion >>
rect 215 35 216 36 
<< m2 >>
rect 225 35 226 36 
<< m1 >>
rect 226 35 227 36 
<< pdiffusion >>
rect 228 35 229 36 
<< pdiffusion >>
rect 229 35 230 36 
<< pdiffusion >>
rect 230 35 231 36 
<< pdiffusion >>
rect 231 35 232 36 
<< pdiffusion >>
rect 232 35 233 36 
<< pdiffusion >>
rect 233 35 234 36 
<< m1 >>
rect 235 35 236 36 
<< pdiffusion >>
rect 264 35 265 36 
<< pdiffusion >>
rect 265 35 266 36 
<< pdiffusion >>
rect 266 35 267 36 
<< pdiffusion >>
rect 267 35 268 36 
<< pdiffusion >>
rect 268 35 269 36 
<< pdiffusion >>
rect 269 35 270 36 
<< m1 >>
rect 278 35 279 36 
<< m1 >>
rect 280 35 281 36 
<< pdiffusion >>
rect 282 35 283 36 
<< pdiffusion >>
rect 283 35 284 36 
<< pdiffusion >>
rect 284 35 285 36 
<< pdiffusion >>
rect 285 35 286 36 
<< pdiffusion >>
rect 286 35 287 36 
<< pdiffusion >>
rect 287 35 288 36 
<< pdiffusion >>
rect 300 35 301 36 
<< m1 >>
rect 301 35 302 36 
<< pdiffusion >>
rect 301 35 302 36 
<< pdiffusion >>
rect 302 35 303 36 
<< pdiffusion >>
rect 303 35 304 36 
<< pdiffusion >>
rect 304 35 305 36 
<< pdiffusion >>
rect 305 35 306 36 
<< pdiffusion >>
rect 318 35 319 36 
<< pdiffusion >>
rect 319 35 320 36 
<< pdiffusion >>
rect 320 35 321 36 
<< pdiffusion >>
rect 321 35 322 36 
<< pdiffusion >>
rect 322 35 323 36 
<< pdiffusion >>
rect 323 35 324 36 
<< m1 >>
rect 334 35 335 36 
<< pdiffusion >>
rect 336 35 337 36 
<< pdiffusion >>
rect 337 35 338 36 
<< pdiffusion >>
rect 338 35 339 36 
<< pdiffusion >>
rect 339 35 340 36 
<< m1 >>
rect 340 35 341 36 
<< pdiffusion >>
rect 340 35 341 36 
<< pdiffusion >>
rect 341 35 342 36 
<< pdiffusion >>
rect 354 35 355 36 
<< pdiffusion >>
rect 355 35 356 36 
<< pdiffusion >>
rect 356 35 357 36 
<< pdiffusion >>
rect 357 35 358 36 
<< pdiffusion >>
rect 358 35 359 36 
<< pdiffusion >>
rect 359 35 360 36 
<< pdiffusion >>
rect 372 35 373 36 
<< m1 >>
rect 373 35 374 36 
<< pdiffusion >>
rect 373 35 374 36 
<< pdiffusion >>
rect 374 35 375 36 
<< pdiffusion >>
rect 375 35 376 36 
<< pdiffusion >>
rect 376 35 377 36 
<< pdiffusion >>
rect 377 35 378 36 
<< m1 >>
rect 388 35 389 36 
<< pdiffusion >>
rect 390 35 391 36 
<< pdiffusion >>
rect 391 35 392 36 
<< pdiffusion >>
rect 392 35 393 36 
<< pdiffusion >>
rect 393 35 394 36 
<< pdiffusion >>
rect 394 35 395 36 
<< pdiffusion >>
rect 395 35 396 36 
<< m1 >>
rect 406 35 407 36 
<< pdiffusion >>
rect 408 35 409 36 
<< pdiffusion >>
rect 409 35 410 36 
<< pdiffusion >>
rect 410 35 411 36 
<< pdiffusion >>
rect 411 35 412 36 
<< pdiffusion >>
rect 412 35 413 36 
<< pdiffusion >>
rect 413 35 414 36 
<< pdiffusion >>
rect 426 35 427 36 
<< pdiffusion >>
rect 427 35 428 36 
<< pdiffusion >>
rect 428 35 429 36 
<< pdiffusion >>
rect 429 35 430 36 
<< pdiffusion >>
rect 430 35 431 36 
<< pdiffusion >>
rect 431 35 432 36 
<< m1 >>
rect 433 35 434 36 
<< pdiffusion >>
rect 444 35 445 36 
<< pdiffusion >>
rect 445 35 446 36 
<< pdiffusion >>
rect 446 35 447 36 
<< pdiffusion >>
rect 447 35 448 36 
<< pdiffusion >>
rect 448 35 449 36 
<< pdiffusion >>
rect 449 35 450 36 
<< pdiffusion >>
rect 462 35 463 36 
<< pdiffusion >>
rect 463 35 464 36 
<< pdiffusion >>
rect 464 35 465 36 
<< pdiffusion >>
rect 465 35 466 36 
<< m1 >>
rect 466 35 467 36 
<< pdiffusion >>
rect 466 35 467 36 
<< pdiffusion >>
rect 467 35 468 36 
<< pdiffusion >>
rect 480 35 481 36 
<< pdiffusion >>
rect 481 35 482 36 
<< pdiffusion >>
rect 482 35 483 36 
<< pdiffusion >>
rect 483 35 484 36 
<< m1 >>
rect 484 35 485 36 
<< pdiffusion >>
rect 484 35 485 36 
<< pdiffusion >>
rect 485 35 486 36 
<< m1 >>
rect 487 35 488 36 
<< m1 >>
rect 505 35 506 36 
<< pdiffusion >>
rect 516 35 517 36 
<< pdiffusion >>
rect 517 35 518 36 
<< pdiffusion >>
rect 518 35 519 36 
<< pdiffusion >>
rect 519 35 520 36 
<< pdiffusion >>
rect 520 35 521 36 
<< pdiffusion >>
rect 521 35 522 36 
<< m1 >>
rect 64 36 65 37 
<< m1 >>
rect 85 36 86 37 
<< m1 >>
rect 106 36 107 37 
<< m1 >>
rect 111 36 112 37 
<< m1 >>
rect 127 36 128 37 
<< m1 >>
rect 145 36 146 37 
<< m1 >>
rect 157 36 158 37 
<< m1 >>
rect 160 36 161 37 
<< m1 >>
rect 193 36 194 37 
<< m1 >>
rect 208 36 209 37 
<< m1 >>
rect 214 36 215 37 
<< m2 >>
rect 225 36 226 37 
<< m1 >>
rect 226 36 227 37 
<< m1 >>
rect 235 36 236 37 
<< m1 >>
rect 278 36 279 37 
<< m1 >>
rect 280 36 281 37 
<< m1 >>
rect 301 36 302 37 
<< m1 >>
rect 334 36 335 37 
<< m1 >>
rect 340 36 341 37 
<< m1 >>
rect 373 36 374 37 
<< m1 >>
rect 388 36 389 37 
<< m1 >>
rect 406 36 407 37 
<< m1 >>
rect 433 36 434 37 
<< m1 >>
rect 466 36 467 37 
<< m1 >>
rect 484 36 485 37 
<< m1 >>
rect 487 36 488 37 
<< m1 >>
rect 505 36 506 37 
<< m1 >>
rect 64 37 65 38 
<< m1 >>
rect 85 37 86 38 
<< m1 >>
rect 106 37 107 38 
<< m1 >>
rect 111 37 112 38 
<< m1 >>
rect 127 37 128 38 
<< m1 >>
rect 145 37 146 38 
<< m1 >>
rect 146 37 147 38 
<< m1 >>
rect 147 37 148 38 
<< m1 >>
rect 148 37 149 38 
<< m1 >>
rect 149 37 150 38 
<< m1 >>
rect 150 37 151 38 
<< m1 >>
rect 151 37 152 38 
<< m1 >>
rect 152 37 153 38 
<< m1 >>
rect 153 37 154 38 
<< m1 >>
rect 154 37 155 38 
<< m1 >>
rect 155 37 156 38 
<< m1 >>
rect 156 37 157 38 
<< m1 >>
rect 157 37 158 38 
<< m1 >>
rect 160 37 161 38 
<< m1 >>
rect 161 37 162 38 
<< m1 >>
rect 162 37 163 38 
<< m1 >>
rect 163 37 164 38 
<< m1 >>
rect 193 37 194 38 
<< m1 >>
rect 208 37 209 38 
<< m1 >>
rect 214 37 215 38 
<< m2 >>
rect 225 37 226 38 
<< m1 >>
rect 226 37 227 38 
<< m1 >>
rect 235 37 236 38 
<< m1 >>
rect 278 37 279 38 
<< m1 >>
rect 280 37 281 38 
<< m1 >>
rect 301 37 302 38 
<< m1 >>
rect 334 37 335 38 
<< m1 >>
rect 340 37 341 38 
<< m1 >>
rect 373 37 374 38 
<< m1 >>
rect 388 37 389 38 
<< m1 >>
rect 406 37 407 38 
<< m1 >>
rect 433 37 434 38 
<< m1 >>
rect 466 37 467 38 
<< m1 >>
rect 484 37 485 38 
<< m1 >>
rect 485 37 486 38 
<< m1 >>
rect 486 37 487 38 
<< m1 >>
rect 487 37 488 38 
<< m1 >>
rect 505 37 506 38 
<< m1 >>
rect 64 38 65 39 
<< m1 >>
rect 85 38 86 39 
<< m1 >>
rect 86 38 87 39 
<< m1 >>
rect 87 38 88 39 
<< m1 >>
rect 88 38 89 39 
<< m1 >>
rect 89 38 90 39 
<< m1 >>
rect 90 38 91 39 
<< m1 >>
rect 91 38 92 39 
<< m1 >>
rect 106 38 107 39 
<< m1 >>
rect 111 38 112 39 
<< m1 >>
rect 127 38 128 39 
<< m1 >>
rect 163 38 164 39 
<< m1 >>
rect 193 38 194 39 
<< m1 >>
rect 208 38 209 39 
<< m1 >>
rect 214 38 215 39 
<< m2 >>
rect 225 38 226 39 
<< m1 >>
rect 226 38 227 39 
<< m1 >>
rect 235 38 236 39 
<< m1 >>
rect 278 38 279 39 
<< m1 >>
rect 280 38 281 39 
<< m1 >>
rect 301 38 302 39 
<< m1 >>
rect 334 38 335 39 
<< m1 >>
rect 340 38 341 39 
<< m1 >>
rect 373 38 374 39 
<< m1 >>
rect 374 38 375 39 
<< m1 >>
rect 375 38 376 39 
<< m1 >>
rect 376 38 377 39 
<< m1 >>
rect 377 38 378 39 
<< m1 >>
rect 378 38 379 39 
<< m1 >>
rect 379 38 380 39 
<< m1 >>
rect 380 38 381 39 
<< m1 >>
rect 381 38 382 39 
<< m1 >>
rect 382 38 383 39 
<< m1 >>
rect 383 38 384 39 
<< m1 >>
rect 384 38 385 39 
<< m1 >>
rect 385 38 386 39 
<< m1 >>
rect 386 38 387 39 
<< m1 >>
rect 387 38 388 39 
<< m1 >>
rect 388 38 389 39 
<< m1 >>
rect 406 38 407 39 
<< m1 >>
rect 433 38 434 39 
<< m1 >>
rect 466 38 467 39 
<< m1 >>
rect 505 38 506 39 
<< m1 >>
rect 64 39 65 40 
<< m1 >>
rect 91 39 92 40 
<< m1 >>
rect 106 39 107 40 
<< m1 >>
rect 111 39 112 40 
<< m1 >>
rect 127 39 128 40 
<< m1 >>
rect 163 39 164 40 
<< m1 >>
rect 193 39 194 40 
<< m1 >>
rect 208 39 209 40 
<< m1 >>
rect 214 39 215 40 
<< m2 >>
rect 225 39 226 40 
<< m1 >>
rect 226 39 227 40 
<< m1 >>
rect 235 39 236 40 
<< m1 >>
rect 278 39 279 40 
<< m1 >>
rect 280 39 281 40 
<< m1 >>
rect 301 39 302 40 
<< m1 >>
rect 334 39 335 40 
<< m1 >>
rect 340 39 341 40 
<< m1 >>
rect 406 39 407 40 
<< m1 >>
rect 433 39 434 40 
<< m1 >>
rect 466 39 467 40 
<< m1 >>
rect 505 39 506 40 
<< m1 >>
rect 64 40 65 41 
<< m1 >>
rect 91 40 92 41 
<< m1 >>
rect 100 40 101 41 
<< m1 >>
rect 101 40 102 41 
<< m1 >>
rect 102 40 103 41 
<< m1 >>
rect 103 40 104 41 
<< m1 >>
rect 104 40 105 41 
<< m1 >>
rect 105 40 106 41 
<< m1 >>
rect 106 40 107 41 
<< m1 >>
rect 111 40 112 41 
<< m1 >>
rect 127 40 128 41 
<< m1 >>
rect 163 40 164 41 
<< m1 >>
rect 193 40 194 41 
<< m1 >>
rect 208 40 209 41 
<< m1 >>
rect 209 40 210 41 
<< m1 >>
rect 210 40 211 41 
<< m1 >>
rect 211 40 212 41 
<< m1 >>
rect 212 40 213 41 
<< m1 >>
rect 213 40 214 41 
<< m1 >>
rect 214 40 215 41 
<< m2 >>
rect 225 40 226 41 
<< m1 >>
rect 226 40 227 41 
<< m1 >>
rect 235 40 236 41 
<< m1 >>
rect 278 40 279 41 
<< m1 >>
rect 280 40 281 41 
<< m1 >>
rect 301 40 302 41 
<< m1 >>
rect 334 40 335 41 
<< m1 >>
rect 340 40 341 41 
<< m1 >>
rect 406 40 407 41 
<< m1 >>
rect 407 40 408 41 
<< m1 >>
rect 408 40 409 41 
<< m1 >>
rect 409 40 410 41 
<< m1 >>
rect 433 40 434 41 
<< m1 >>
rect 466 40 467 41 
<< m1 >>
rect 505 40 506 41 
<< m1 >>
rect 64 41 65 42 
<< m1 >>
rect 91 41 92 42 
<< m1 >>
rect 100 41 101 42 
<< m1 >>
rect 111 41 112 42 
<< m1 >>
rect 127 41 128 42 
<< m1 >>
rect 163 41 164 42 
<< m1 >>
rect 193 41 194 42 
<< m2 >>
rect 225 41 226 42 
<< m1 >>
rect 226 41 227 42 
<< m1 >>
rect 235 41 236 42 
<< m2 >>
rect 235 41 236 42 
<< m2c >>
rect 235 41 236 42 
<< m1 >>
rect 235 41 236 42 
<< m2 >>
rect 235 41 236 42 
<< m1 >>
rect 278 41 279 42 
<< m2 >>
rect 278 41 279 42 
<< m2c >>
rect 278 41 279 42 
<< m1 >>
rect 278 41 279 42 
<< m2 >>
rect 278 41 279 42 
<< m1 >>
rect 280 41 281 42 
<< m2 >>
rect 280 41 281 42 
<< m2c >>
rect 280 41 281 42 
<< m1 >>
rect 280 41 281 42 
<< m2 >>
rect 280 41 281 42 
<< m1 >>
rect 301 41 302 42 
<< m1 >>
rect 302 41 303 42 
<< m1 >>
rect 303 41 304 42 
<< m1 >>
rect 304 41 305 42 
<< m1 >>
rect 305 41 306 42 
<< m1 >>
rect 306 41 307 42 
<< m1 >>
rect 307 41 308 42 
<< m1 >>
rect 308 41 309 42 
<< m1 >>
rect 309 41 310 42 
<< m1 >>
rect 310 41 311 42 
<< m1 >>
rect 311 41 312 42 
<< m1 >>
rect 312 41 313 42 
<< m1 >>
rect 313 41 314 42 
<< m1 >>
rect 314 41 315 42 
<< m1 >>
rect 315 41 316 42 
<< m1 >>
rect 316 41 317 42 
<< m1 >>
rect 317 41 318 42 
<< m1 >>
rect 318 41 319 42 
<< m1 >>
rect 319 41 320 42 
<< m1 >>
rect 320 41 321 42 
<< m1 >>
rect 321 41 322 42 
<< m1 >>
rect 322 41 323 42 
<< m1 >>
rect 323 41 324 42 
<< m1 >>
rect 324 41 325 42 
<< m1 >>
rect 325 41 326 42 
<< m1 >>
rect 326 41 327 42 
<< m1 >>
rect 327 41 328 42 
<< m1 >>
rect 328 41 329 42 
<< m1 >>
rect 329 41 330 42 
<< m1 >>
rect 330 41 331 42 
<< m1 >>
rect 331 41 332 42 
<< m1 >>
rect 332 41 333 42 
<< m2 >>
rect 332 41 333 42 
<< m2c >>
rect 332 41 333 42 
<< m1 >>
rect 332 41 333 42 
<< m2 >>
rect 332 41 333 42 
<< m1 >>
rect 334 41 335 42 
<< m2 >>
rect 334 41 335 42 
<< m2c >>
rect 334 41 335 42 
<< m1 >>
rect 334 41 335 42 
<< m2 >>
rect 334 41 335 42 
<< m1 >>
rect 340 41 341 42 
<< m1 >>
rect 409 41 410 42 
<< m1 >>
rect 433 41 434 42 
<< m1 >>
rect 466 41 467 42 
<< m1 >>
rect 505 41 506 42 
<< m2 >>
rect 505 41 506 42 
<< m2c >>
rect 505 41 506 42 
<< m1 >>
rect 505 41 506 42 
<< m2 >>
rect 505 41 506 42 
<< m1 >>
rect 64 42 65 43 
<< m1 >>
rect 91 42 92 43 
<< m1 >>
rect 100 42 101 43 
<< m1 >>
rect 111 42 112 43 
<< m1 >>
rect 127 42 128 43 
<< m1 >>
rect 163 42 164 43 
<< m1 >>
rect 193 42 194 43 
<< m2 >>
rect 225 42 226 43 
<< m1 >>
rect 226 42 227 43 
<< m2 >>
rect 235 42 236 43 
<< m2 >>
rect 246 42 247 43 
<< m2 >>
rect 247 42 248 43 
<< m2 >>
rect 248 42 249 43 
<< m2 >>
rect 249 42 250 43 
<< m2 >>
rect 250 42 251 43 
<< m2 >>
rect 251 42 252 43 
<< m2 >>
rect 252 42 253 43 
<< m2 >>
rect 253 42 254 43 
<< m2 >>
rect 254 42 255 43 
<< m2 >>
rect 255 42 256 43 
<< m2 >>
rect 256 42 257 43 
<< m2 >>
rect 257 42 258 43 
<< m2 >>
rect 258 42 259 43 
<< m2 >>
rect 259 42 260 43 
<< m2 >>
rect 260 42 261 43 
<< m2 >>
rect 261 42 262 43 
<< m2 >>
rect 262 42 263 43 
<< m2 >>
rect 263 42 264 43 
<< m2 >>
rect 264 42 265 43 
<< m2 >>
rect 265 42 266 43 
<< m2 >>
rect 266 42 267 43 
<< m2 >>
rect 267 42 268 43 
<< m2 >>
rect 268 42 269 43 
<< m2 >>
rect 269 42 270 43 
<< m2 >>
rect 270 42 271 43 
<< m2 >>
rect 271 42 272 43 
<< m2 >>
rect 272 42 273 43 
<< m2 >>
rect 273 42 274 43 
<< m2 >>
rect 274 42 275 43 
<< m2 >>
rect 275 42 276 43 
<< m2 >>
rect 276 42 277 43 
<< m2 >>
rect 277 42 278 43 
<< m2 >>
rect 278 42 279 43 
<< m2 >>
rect 280 42 281 43 
<< m2 >>
rect 332 42 333 43 
<< m2 >>
rect 334 42 335 43 
<< m1 >>
rect 340 42 341 43 
<< m1 >>
rect 409 42 410 43 
<< m1 >>
rect 433 42 434 43 
<< m1 >>
rect 466 42 467 43 
<< m2 >>
rect 505 42 506 43 
<< m1 >>
rect 19 43 20 44 
<< m1 >>
rect 20 43 21 44 
<< m1 >>
rect 21 43 22 44 
<< m1 >>
rect 22 43 23 44 
<< m1 >>
rect 23 43 24 44 
<< m1 >>
rect 24 43 25 44 
<< m1 >>
rect 25 43 26 44 
<< m1 >>
rect 26 43 27 44 
<< m1 >>
rect 27 43 28 44 
<< m1 >>
rect 28 43 29 44 
<< m1 >>
rect 29 43 30 44 
<< m1 >>
rect 30 43 31 44 
<< m1 >>
rect 31 43 32 44 
<< m1 >>
rect 32 43 33 44 
<< m1 >>
rect 33 43 34 44 
<< m1 >>
rect 34 43 35 44 
<< m1 >>
rect 52 43 53 44 
<< m1 >>
rect 53 43 54 44 
<< m1 >>
rect 54 43 55 44 
<< m1 >>
rect 55 43 56 44 
<< m1 >>
rect 56 43 57 44 
<< m1 >>
rect 57 43 58 44 
<< m1 >>
rect 58 43 59 44 
<< m1 >>
rect 59 43 60 44 
<< m1 >>
rect 60 43 61 44 
<< m1 >>
rect 61 43 62 44 
<< m1 >>
rect 62 43 63 44 
<< m2 >>
rect 62 43 63 44 
<< m2c >>
rect 62 43 63 44 
<< m1 >>
rect 62 43 63 44 
<< m2 >>
rect 62 43 63 44 
<< m2 >>
rect 63 43 64 44 
<< m1 >>
rect 64 43 65 44 
<< m2 >>
rect 64 43 65 44 
<< m2 >>
rect 65 43 66 44 
<< m1 >>
rect 66 43 67 44 
<< m2 >>
rect 66 43 67 44 
<< m2c >>
rect 66 43 67 44 
<< m1 >>
rect 66 43 67 44 
<< m2 >>
rect 66 43 67 44 
<< m1 >>
rect 67 43 68 44 
<< m1 >>
rect 68 43 69 44 
<< m1 >>
rect 69 43 70 44 
<< m1 >>
rect 70 43 71 44 
<< m1 >>
rect 91 43 92 44 
<< m1 >>
rect 100 43 101 44 
<< m1 >>
rect 111 43 112 44 
<< m1 >>
rect 127 43 128 44 
<< m1 >>
rect 163 43 164 44 
<< m1 >>
rect 165 43 166 44 
<< m1 >>
rect 166 43 167 44 
<< m1 >>
rect 167 43 168 44 
<< m1 >>
rect 168 43 169 44 
<< m1 >>
rect 169 43 170 44 
<< m1 >>
rect 170 43 171 44 
<< m1 >>
rect 171 43 172 44 
<< m1 >>
rect 172 43 173 44 
<< m1 >>
rect 173 43 174 44 
<< m1 >>
rect 174 43 175 44 
<< m1 >>
rect 175 43 176 44 
<< m1 >>
rect 176 43 177 44 
<< m1 >>
rect 177 43 178 44 
<< m1 >>
rect 178 43 179 44 
<< m1 >>
rect 179 43 180 44 
<< m1 >>
rect 180 43 181 44 
<< m1 >>
rect 181 43 182 44 
<< m1 >>
rect 182 43 183 44 
<< m1 >>
rect 183 43 184 44 
<< m1 >>
rect 184 43 185 44 
<< m1 >>
rect 185 43 186 44 
<< m1 >>
rect 186 43 187 44 
<< m1 >>
rect 187 43 188 44 
<< m1 >>
rect 188 43 189 44 
<< m1 >>
rect 189 43 190 44 
<< m1 >>
rect 190 43 191 44 
<< m1 >>
rect 191 43 192 44 
<< m1 >>
rect 192 43 193 44 
<< m1 >>
rect 193 43 194 44 
<< m2 >>
rect 225 43 226 44 
<< m1 >>
rect 226 43 227 44 
<< m1 >>
rect 235 43 236 44 
<< m2 >>
rect 235 43 236 44 
<< m1 >>
rect 236 43 237 44 
<< m1 >>
rect 237 43 238 44 
<< m1 >>
rect 238 43 239 44 
<< m1 >>
rect 239 43 240 44 
<< m1 >>
rect 240 43 241 44 
<< m1 >>
rect 241 43 242 44 
<< m1 >>
rect 242 43 243 44 
<< m1 >>
rect 243 43 244 44 
<< m1 >>
rect 244 43 245 44 
<< m1 >>
rect 245 43 246 44 
<< m1 >>
rect 246 43 247 44 
<< m2 >>
rect 246 43 247 44 
<< m1 >>
rect 247 43 248 44 
<< m1 >>
rect 248 43 249 44 
<< m1 >>
rect 249 43 250 44 
<< m1 >>
rect 250 43 251 44 
<< m1 >>
rect 251 43 252 44 
<< m1 >>
rect 252 43 253 44 
<< m1 >>
rect 253 43 254 44 
<< m1 >>
rect 254 43 255 44 
<< m1 >>
rect 255 43 256 44 
<< m1 >>
rect 256 43 257 44 
<< m1 >>
rect 257 43 258 44 
<< m1 >>
rect 258 43 259 44 
<< m1 >>
rect 259 43 260 44 
<< m1 >>
rect 260 43 261 44 
<< m1 >>
rect 261 43 262 44 
<< m1 >>
rect 262 43 263 44 
<< m1 >>
rect 263 43 264 44 
<< m1 >>
rect 264 43 265 44 
<< m1 >>
rect 265 43 266 44 
<< m1 >>
rect 266 43 267 44 
<< m1 >>
rect 267 43 268 44 
<< m1 >>
rect 268 43 269 44 
<< m1 >>
rect 269 43 270 44 
<< m1 >>
rect 270 43 271 44 
<< m1 >>
rect 271 43 272 44 
<< m1 >>
rect 272 43 273 44 
<< m1 >>
rect 273 43 274 44 
<< m1 >>
rect 274 43 275 44 
<< m1 >>
rect 275 43 276 44 
<< m1 >>
rect 276 43 277 44 
<< m1 >>
rect 277 43 278 44 
<< m1 >>
rect 278 43 279 44 
<< m1 >>
rect 279 43 280 44 
<< m1 >>
rect 280 43 281 44 
<< m2 >>
rect 280 43 281 44 
<< m1 >>
rect 281 43 282 44 
<< m1 >>
rect 282 43 283 44 
<< m1 >>
rect 283 43 284 44 
<< m1 >>
rect 284 43 285 44 
<< m1 >>
rect 285 43 286 44 
<< m1 >>
rect 286 43 287 44 
<< m1 >>
rect 287 43 288 44 
<< m1 >>
rect 288 43 289 44 
<< m1 >>
rect 289 43 290 44 
<< m1 >>
rect 290 43 291 44 
<< m1 >>
rect 291 43 292 44 
<< m1 >>
rect 292 43 293 44 
<< m1 >>
rect 293 43 294 44 
<< m1 >>
rect 294 43 295 44 
<< m1 >>
rect 295 43 296 44 
<< m1 >>
rect 296 43 297 44 
<< m1 >>
rect 297 43 298 44 
<< m1 >>
rect 298 43 299 44 
<< m1 >>
rect 299 43 300 44 
<< m1 >>
rect 300 43 301 44 
<< m1 >>
rect 301 43 302 44 
<< m1 >>
rect 302 43 303 44 
<< m1 >>
rect 303 43 304 44 
<< m1 >>
rect 304 43 305 44 
<< m1 >>
rect 305 43 306 44 
<< m1 >>
rect 306 43 307 44 
<< m1 >>
rect 307 43 308 44 
<< m1 >>
rect 308 43 309 44 
<< m1 >>
rect 309 43 310 44 
<< m1 >>
rect 310 43 311 44 
<< m1 >>
rect 311 43 312 44 
<< m1 >>
rect 312 43 313 44 
<< m1 >>
rect 313 43 314 44 
<< m1 >>
rect 314 43 315 44 
<< m1 >>
rect 315 43 316 44 
<< m1 >>
rect 316 43 317 44 
<< m1 >>
rect 317 43 318 44 
<< m1 >>
rect 318 43 319 44 
<< m1 >>
rect 319 43 320 44 
<< m1 >>
rect 320 43 321 44 
<< m1 >>
rect 321 43 322 44 
<< m1 >>
rect 322 43 323 44 
<< m1 >>
rect 323 43 324 44 
<< m1 >>
rect 324 43 325 44 
<< m1 >>
rect 325 43 326 44 
<< m1 >>
rect 326 43 327 44 
<< m1 >>
rect 327 43 328 44 
<< m1 >>
rect 328 43 329 44 
<< m1 >>
rect 329 43 330 44 
<< m1 >>
rect 330 43 331 44 
<< m1 >>
rect 331 43 332 44 
<< m1 >>
rect 332 43 333 44 
<< m2 >>
rect 332 43 333 44 
<< m1 >>
rect 333 43 334 44 
<< m1 >>
rect 334 43 335 44 
<< m2 >>
rect 334 43 335 44 
<< m1 >>
rect 335 43 336 44 
<< m1 >>
rect 336 43 337 44 
<< m1 >>
rect 337 43 338 44 
<< m1 >>
rect 338 43 339 44 
<< m1 >>
rect 339 43 340 44 
<< m1 >>
rect 340 43 341 44 
<< m1 >>
rect 409 43 410 44 
<< m1 >>
rect 433 43 434 44 
<< m1 >>
rect 466 43 467 44 
<< m1 >>
rect 487 43 488 44 
<< m1 >>
rect 488 43 489 44 
<< m1 >>
rect 489 43 490 44 
<< m1 >>
rect 490 43 491 44 
<< m1 >>
rect 491 43 492 44 
<< m1 >>
rect 492 43 493 44 
<< m1 >>
rect 493 43 494 44 
<< m1 >>
rect 494 43 495 44 
<< m1 >>
rect 495 43 496 44 
<< m1 >>
rect 496 43 497 44 
<< m1 >>
rect 497 43 498 44 
<< m1 >>
rect 498 43 499 44 
<< m1 >>
rect 499 43 500 44 
<< m1 >>
rect 500 43 501 44 
<< m1 >>
rect 501 43 502 44 
<< m1 >>
rect 502 43 503 44 
<< m1 >>
rect 503 43 504 44 
<< m1 >>
rect 504 43 505 44 
<< m1 >>
rect 505 43 506 44 
<< m2 >>
rect 505 43 506 44 
<< m1 >>
rect 506 43 507 44 
<< m1 >>
rect 507 43 508 44 
<< m1 >>
rect 508 43 509 44 
<< m1 >>
rect 509 43 510 44 
<< m1 >>
rect 510 43 511 44 
<< m1 >>
rect 511 43 512 44 
<< m1 >>
rect 512 43 513 44 
<< m1 >>
rect 513 43 514 44 
<< m1 >>
rect 514 43 515 44 
<< m1 >>
rect 515 43 516 44 
<< m1 >>
rect 516 43 517 44 
<< m1 >>
rect 517 43 518 44 
<< m1 >>
rect 518 43 519 44 
<< m1 >>
rect 519 43 520 44 
<< m1 >>
rect 520 43 521 44 
<< m1 >>
rect 19 44 20 45 
<< m1 >>
rect 34 44 35 45 
<< m1 >>
rect 52 44 53 45 
<< m1 >>
rect 64 44 65 45 
<< m1 >>
rect 70 44 71 45 
<< m1 >>
rect 91 44 92 45 
<< m1 >>
rect 100 44 101 45 
<< m1 >>
rect 111 44 112 45 
<< m1 >>
rect 127 44 128 45 
<< m1 >>
rect 163 44 164 45 
<< m1 >>
rect 165 44 166 45 
<< m2 >>
rect 225 44 226 45 
<< m1 >>
rect 226 44 227 45 
<< m1 >>
rect 235 44 236 45 
<< m2 >>
rect 235 44 236 45 
<< m2 >>
rect 246 44 247 45 
<< m2 >>
rect 280 44 281 45 
<< m2 >>
rect 332 44 333 45 
<< m2 >>
rect 334 44 335 45 
<< m1 >>
rect 409 44 410 45 
<< m1 >>
rect 433 44 434 45 
<< m1 >>
rect 466 44 467 45 
<< m1 >>
rect 487 44 488 45 
<< m2 >>
rect 505 44 506 45 
<< m1 >>
rect 520 44 521 45 
<< m1 >>
rect 19 45 20 46 
<< m1 >>
rect 34 45 35 46 
<< m1 >>
rect 52 45 53 46 
<< m1 >>
rect 64 45 65 46 
<< m1 >>
rect 70 45 71 46 
<< m1 >>
rect 91 45 92 46 
<< m1 >>
rect 100 45 101 46 
<< m1 >>
rect 103 45 104 46 
<< m1 >>
rect 104 45 105 46 
<< m1 >>
rect 105 45 106 46 
<< m1 >>
rect 106 45 107 46 
<< m1 >>
rect 107 45 108 46 
<< m1 >>
rect 108 45 109 46 
<< m1 >>
rect 109 45 110 46 
<< m1 >>
rect 111 45 112 46 
<< m1 >>
rect 127 45 128 46 
<< m1 >>
rect 163 45 164 46 
<< m1 >>
rect 165 45 166 46 
<< m2 >>
rect 225 45 226 46 
<< m1 >>
rect 226 45 227 46 
<< m1 >>
rect 235 45 236 46 
<< m2 >>
rect 235 45 236 46 
<< m2 >>
rect 236 45 237 46 
<< m1 >>
rect 237 45 238 46 
<< m2 >>
rect 237 45 238 46 
<< m2c >>
rect 237 45 238 46 
<< m1 >>
rect 237 45 238 46 
<< m2 >>
rect 237 45 238 46 
<< m1 >>
rect 244 45 245 46 
<< m1 >>
rect 245 45 246 46 
<< m1 >>
rect 246 45 247 46 
<< m2 >>
rect 246 45 247 46 
<< m2c >>
rect 246 45 247 46 
<< m1 >>
rect 246 45 247 46 
<< m2 >>
rect 246 45 247 46 
<< m1 >>
rect 280 45 281 46 
<< m2 >>
rect 280 45 281 46 
<< m2c >>
rect 280 45 281 46 
<< m1 >>
rect 280 45 281 46 
<< m2 >>
rect 280 45 281 46 
<< m1 >>
rect 283 45 284 46 
<< m1 >>
rect 284 45 285 46 
<< m1 >>
rect 285 45 286 46 
<< m1 >>
rect 286 45 287 46 
<< m1 >>
rect 287 45 288 46 
<< m1 >>
rect 288 45 289 46 
<< m1 >>
rect 289 45 290 46 
<< m1 >>
rect 332 45 333 46 
<< m2 >>
rect 332 45 333 46 
<< m2c >>
rect 332 45 333 46 
<< m1 >>
rect 332 45 333 46 
<< m2 >>
rect 332 45 333 46 
<< m1 >>
rect 334 45 335 46 
<< m2 >>
rect 334 45 335 46 
<< m2c >>
rect 334 45 335 46 
<< m1 >>
rect 334 45 335 46 
<< m2 >>
rect 334 45 335 46 
<< m1 >>
rect 409 45 410 46 
<< m1 >>
rect 433 45 434 46 
<< m1 >>
rect 466 45 467 46 
<< m1 >>
rect 487 45 488 46 
<< m1 >>
rect 505 45 506 46 
<< m2 >>
rect 505 45 506 46 
<< m2c >>
rect 505 45 506 46 
<< m1 >>
rect 505 45 506 46 
<< m2 >>
rect 505 45 506 46 
<< m1 >>
rect 520 45 521 46 
<< m1 >>
rect 19 46 20 47 
<< m1 >>
rect 34 46 35 47 
<< m1 >>
rect 52 46 53 47 
<< m1 >>
rect 64 46 65 47 
<< m1 >>
rect 70 46 71 47 
<< m1 >>
rect 91 46 92 47 
<< m1 >>
rect 100 46 101 47 
<< m1 >>
rect 103 46 104 47 
<< m1 >>
rect 109 46 110 47 
<< m1 >>
rect 111 46 112 47 
<< m1 >>
rect 124 46 125 47 
<< m1 >>
rect 125 46 126 47 
<< m1 >>
rect 126 46 127 47 
<< m1 >>
rect 127 46 128 47 
<< m1 >>
rect 163 46 164 47 
<< m1 >>
rect 165 46 166 47 
<< m1 >>
rect 178 46 179 47 
<< m1 >>
rect 179 46 180 47 
<< m1 >>
rect 180 46 181 47 
<< m1 >>
rect 181 46 182 47 
<< m1 >>
rect 182 46 183 47 
<< m1 >>
rect 183 46 184 47 
<< m1 >>
rect 184 46 185 47 
<< m1 >>
rect 185 46 186 47 
<< m1 >>
rect 186 46 187 47 
<< m1 >>
rect 187 46 188 47 
<< m1 >>
rect 188 46 189 47 
<< m1 >>
rect 189 46 190 47 
<< m1 >>
rect 190 46 191 47 
<< m2 >>
rect 225 46 226 47 
<< m1 >>
rect 226 46 227 47 
<< m1 >>
rect 235 46 236 47 
<< m1 >>
rect 237 46 238 47 
<< m1 >>
rect 244 46 245 47 
<< m1 >>
rect 250 46 251 47 
<< m1 >>
rect 251 46 252 47 
<< m1 >>
rect 252 46 253 47 
<< m1 >>
rect 253 46 254 47 
<< m1 >>
rect 280 46 281 47 
<< m1 >>
rect 283 46 284 47 
<< m1 >>
rect 289 46 290 47 
<< m1 >>
rect 332 46 333 47 
<< m1 >>
rect 334 46 335 47 
<< m1 >>
rect 388 46 389 47 
<< m1 >>
rect 389 46 390 47 
<< m1 >>
rect 390 46 391 47 
<< m1 >>
rect 391 46 392 47 
<< m1 >>
rect 409 46 410 47 
<< m1 >>
rect 433 46 434 47 
<< m1 >>
rect 466 46 467 47 
<< m1 >>
rect 487 46 488 47 
<< m1 >>
rect 505 46 506 47 
<< m1 >>
rect 520 46 521 47 
<< m1 >>
rect 19 47 20 48 
<< m1 >>
rect 34 47 35 48 
<< m1 >>
rect 52 47 53 48 
<< m1 >>
rect 64 47 65 48 
<< m1 >>
rect 70 47 71 48 
<< m1 >>
rect 91 47 92 48 
<< m1 >>
rect 100 47 101 48 
<< m1 >>
rect 103 47 104 48 
<< m1 >>
rect 109 47 110 48 
<< m1 >>
rect 111 47 112 48 
<< m1 >>
rect 124 47 125 48 
<< m1 >>
rect 163 47 164 48 
<< m1 >>
rect 165 47 166 48 
<< m1 >>
rect 178 47 179 48 
<< m1 >>
rect 190 47 191 48 
<< m2 >>
rect 225 47 226 48 
<< m1 >>
rect 226 47 227 48 
<< m1 >>
rect 235 47 236 48 
<< m1 >>
rect 237 47 238 48 
<< m1 >>
rect 244 47 245 48 
<< m1 >>
rect 250 47 251 48 
<< m1 >>
rect 253 47 254 48 
<< m1 >>
rect 280 47 281 48 
<< m1 >>
rect 283 47 284 48 
<< m1 >>
rect 289 47 290 48 
<< m1 >>
rect 332 47 333 48 
<< m1 >>
rect 334 47 335 48 
<< m1 >>
rect 388 47 389 48 
<< m1 >>
rect 391 47 392 48 
<< m1 >>
rect 409 47 410 48 
<< m1 >>
rect 433 47 434 48 
<< m1 >>
rect 466 47 467 48 
<< m1 >>
rect 487 47 488 48 
<< m1 >>
rect 505 47 506 48 
<< m1 >>
rect 520 47 521 48 
<< pdiffusion >>
rect 12 48 13 49 
<< pdiffusion >>
rect 13 48 14 49 
<< pdiffusion >>
rect 14 48 15 49 
<< pdiffusion >>
rect 15 48 16 49 
<< pdiffusion >>
rect 16 48 17 49 
<< pdiffusion >>
rect 17 48 18 49 
<< m1 >>
rect 19 48 20 49 
<< pdiffusion >>
rect 30 48 31 49 
<< pdiffusion >>
rect 31 48 32 49 
<< pdiffusion >>
rect 32 48 33 49 
<< pdiffusion >>
rect 33 48 34 49 
<< m1 >>
rect 34 48 35 49 
<< pdiffusion >>
rect 34 48 35 49 
<< pdiffusion >>
rect 35 48 36 49 
<< pdiffusion >>
rect 48 48 49 49 
<< pdiffusion >>
rect 49 48 50 49 
<< pdiffusion >>
rect 50 48 51 49 
<< pdiffusion >>
rect 51 48 52 49 
<< m1 >>
rect 52 48 53 49 
<< pdiffusion >>
rect 52 48 53 49 
<< pdiffusion >>
rect 53 48 54 49 
<< m1 >>
rect 64 48 65 49 
<< pdiffusion >>
rect 66 48 67 49 
<< pdiffusion >>
rect 67 48 68 49 
<< pdiffusion >>
rect 68 48 69 49 
<< pdiffusion >>
rect 69 48 70 49 
<< m1 >>
rect 70 48 71 49 
<< pdiffusion >>
rect 70 48 71 49 
<< pdiffusion >>
rect 71 48 72 49 
<< pdiffusion >>
rect 84 48 85 49 
<< pdiffusion >>
rect 85 48 86 49 
<< pdiffusion >>
rect 86 48 87 49 
<< pdiffusion >>
rect 87 48 88 49 
<< pdiffusion >>
rect 88 48 89 49 
<< pdiffusion >>
rect 89 48 90 49 
<< m1 >>
rect 91 48 92 49 
<< m1 >>
rect 100 48 101 49 
<< pdiffusion >>
rect 102 48 103 49 
<< m1 >>
rect 103 48 104 49 
<< pdiffusion >>
rect 103 48 104 49 
<< pdiffusion >>
rect 104 48 105 49 
<< pdiffusion >>
rect 105 48 106 49 
<< pdiffusion >>
rect 106 48 107 49 
<< pdiffusion >>
rect 107 48 108 49 
<< m1 >>
rect 109 48 110 49 
<< m1 >>
rect 111 48 112 49 
<< pdiffusion >>
rect 120 48 121 49 
<< pdiffusion >>
rect 121 48 122 49 
<< pdiffusion >>
rect 122 48 123 49 
<< pdiffusion >>
rect 123 48 124 49 
<< m1 >>
rect 124 48 125 49 
<< pdiffusion >>
rect 124 48 125 49 
<< pdiffusion >>
rect 125 48 126 49 
<< pdiffusion >>
rect 138 48 139 49 
<< pdiffusion >>
rect 139 48 140 49 
<< pdiffusion >>
rect 140 48 141 49 
<< pdiffusion >>
rect 141 48 142 49 
<< pdiffusion >>
rect 142 48 143 49 
<< pdiffusion >>
rect 143 48 144 49 
<< pdiffusion >>
rect 156 48 157 49 
<< pdiffusion >>
rect 157 48 158 49 
<< pdiffusion >>
rect 158 48 159 49 
<< pdiffusion >>
rect 159 48 160 49 
<< pdiffusion >>
rect 160 48 161 49 
<< pdiffusion >>
rect 161 48 162 49 
<< m1 >>
rect 163 48 164 49 
<< m1 >>
rect 165 48 166 49 
<< pdiffusion >>
rect 174 48 175 49 
<< pdiffusion >>
rect 175 48 176 49 
<< pdiffusion >>
rect 176 48 177 49 
<< pdiffusion >>
rect 177 48 178 49 
<< m1 >>
rect 178 48 179 49 
<< pdiffusion >>
rect 178 48 179 49 
<< pdiffusion >>
rect 179 48 180 49 
<< m1 >>
rect 190 48 191 49 
<< pdiffusion >>
rect 192 48 193 49 
<< pdiffusion >>
rect 193 48 194 49 
<< pdiffusion >>
rect 194 48 195 49 
<< pdiffusion >>
rect 195 48 196 49 
<< pdiffusion >>
rect 196 48 197 49 
<< pdiffusion >>
rect 197 48 198 49 
<< pdiffusion >>
rect 210 48 211 49 
<< pdiffusion >>
rect 211 48 212 49 
<< pdiffusion >>
rect 212 48 213 49 
<< pdiffusion >>
rect 213 48 214 49 
<< pdiffusion >>
rect 214 48 215 49 
<< pdiffusion >>
rect 215 48 216 49 
<< m2 >>
rect 225 48 226 49 
<< m1 >>
rect 226 48 227 49 
<< pdiffusion >>
rect 228 48 229 49 
<< pdiffusion >>
rect 229 48 230 49 
<< pdiffusion >>
rect 230 48 231 49 
<< pdiffusion >>
rect 231 48 232 49 
<< pdiffusion >>
rect 232 48 233 49 
<< pdiffusion >>
rect 233 48 234 49 
<< m1 >>
rect 235 48 236 49 
<< m1 >>
rect 237 48 238 49 
<< m1 >>
rect 244 48 245 49 
<< pdiffusion >>
rect 246 48 247 49 
<< pdiffusion >>
rect 247 48 248 49 
<< pdiffusion >>
rect 248 48 249 49 
<< pdiffusion >>
rect 249 48 250 49 
<< m1 >>
rect 250 48 251 49 
<< pdiffusion >>
rect 250 48 251 49 
<< pdiffusion >>
rect 251 48 252 49 
<< m1 >>
rect 253 48 254 49 
<< pdiffusion >>
rect 264 48 265 49 
<< pdiffusion >>
rect 265 48 266 49 
<< pdiffusion >>
rect 266 48 267 49 
<< pdiffusion >>
rect 267 48 268 49 
<< pdiffusion >>
rect 268 48 269 49 
<< pdiffusion >>
rect 269 48 270 49 
<< m1 >>
rect 280 48 281 49 
<< pdiffusion >>
rect 282 48 283 49 
<< m1 >>
rect 283 48 284 49 
<< pdiffusion >>
rect 283 48 284 49 
<< pdiffusion >>
rect 284 48 285 49 
<< pdiffusion >>
rect 285 48 286 49 
<< pdiffusion >>
rect 286 48 287 49 
<< pdiffusion >>
rect 287 48 288 49 
<< m1 >>
rect 289 48 290 49 
<< pdiffusion >>
rect 300 48 301 49 
<< pdiffusion >>
rect 301 48 302 49 
<< pdiffusion >>
rect 302 48 303 49 
<< pdiffusion >>
rect 303 48 304 49 
<< pdiffusion >>
rect 304 48 305 49 
<< pdiffusion >>
rect 305 48 306 49 
<< pdiffusion >>
rect 318 48 319 49 
<< pdiffusion >>
rect 319 48 320 49 
<< pdiffusion >>
rect 320 48 321 49 
<< pdiffusion >>
rect 321 48 322 49 
<< pdiffusion >>
rect 322 48 323 49 
<< pdiffusion >>
rect 323 48 324 49 
<< m1 >>
rect 332 48 333 49 
<< m1 >>
rect 334 48 335 49 
<< pdiffusion >>
rect 336 48 337 49 
<< pdiffusion >>
rect 337 48 338 49 
<< pdiffusion >>
rect 338 48 339 49 
<< pdiffusion >>
rect 339 48 340 49 
<< pdiffusion >>
rect 340 48 341 49 
<< pdiffusion >>
rect 341 48 342 49 
<< pdiffusion >>
rect 354 48 355 49 
<< pdiffusion >>
rect 355 48 356 49 
<< pdiffusion >>
rect 356 48 357 49 
<< pdiffusion >>
rect 357 48 358 49 
<< pdiffusion >>
rect 358 48 359 49 
<< pdiffusion >>
rect 359 48 360 49 
<< pdiffusion >>
rect 372 48 373 49 
<< pdiffusion >>
rect 373 48 374 49 
<< pdiffusion >>
rect 374 48 375 49 
<< pdiffusion >>
rect 375 48 376 49 
<< pdiffusion >>
rect 376 48 377 49 
<< pdiffusion >>
rect 377 48 378 49 
<< m1 >>
rect 388 48 389 49 
<< pdiffusion >>
rect 390 48 391 49 
<< m1 >>
rect 391 48 392 49 
<< pdiffusion >>
rect 391 48 392 49 
<< pdiffusion >>
rect 392 48 393 49 
<< pdiffusion >>
rect 393 48 394 49 
<< pdiffusion >>
rect 394 48 395 49 
<< pdiffusion >>
rect 395 48 396 49 
<< pdiffusion >>
rect 408 48 409 49 
<< m1 >>
rect 409 48 410 49 
<< pdiffusion >>
rect 409 48 410 49 
<< pdiffusion >>
rect 410 48 411 49 
<< pdiffusion >>
rect 411 48 412 49 
<< pdiffusion >>
rect 412 48 413 49 
<< pdiffusion >>
rect 413 48 414 49 
<< pdiffusion >>
rect 426 48 427 49 
<< pdiffusion >>
rect 427 48 428 49 
<< pdiffusion >>
rect 428 48 429 49 
<< pdiffusion >>
rect 429 48 430 49 
<< pdiffusion >>
rect 430 48 431 49 
<< pdiffusion >>
rect 431 48 432 49 
<< m1 >>
rect 433 48 434 49 
<< pdiffusion >>
rect 444 48 445 49 
<< pdiffusion >>
rect 445 48 446 49 
<< pdiffusion >>
rect 446 48 447 49 
<< pdiffusion >>
rect 447 48 448 49 
<< pdiffusion >>
rect 448 48 449 49 
<< pdiffusion >>
rect 449 48 450 49 
<< pdiffusion >>
rect 462 48 463 49 
<< pdiffusion >>
rect 463 48 464 49 
<< pdiffusion >>
rect 464 48 465 49 
<< pdiffusion >>
rect 465 48 466 49 
<< m1 >>
rect 466 48 467 49 
<< pdiffusion >>
rect 466 48 467 49 
<< pdiffusion >>
rect 467 48 468 49 
<< pdiffusion >>
rect 480 48 481 49 
<< pdiffusion >>
rect 481 48 482 49 
<< pdiffusion >>
rect 482 48 483 49 
<< pdiffusion >>
rect 483 48 484 49 
<< pdiffusion >>
rect 484 48 485 49 
<< pdiffusion >>
rect 485 48 486 49 
<< m1 >>
rect 487 48 488 49 
<< pdiffusion >>
rect 498 48 499 49 
<< pdiffusion >>
rect 499 48 500 49 
<< pdiffusion >>
rect 500 48 501 49 
<< pdiffusion >>
rect 501 48 502 49 
<< pdiffusion >>
rect 502 48 503 49 
<< pdiffusion >>
rect 503 48 504 49 
<< m1 >>
rect 505 48 506 49 
<< pdiffusion >>
rect 516 48 517 49 
<< pdiffusion >>
rect 517 48 518 49 
<< pdiffusion >>
rect 518 48 519 49 
<< pdiffusion >>
rect 519 48 520 49 
<< m1 >>
rect 520 48 521 49 
<< pdiffusion >>
rect 520 48 521 49 
<< pdiffusion >>
rect 521 48 522 49 
<< pdiffusion >>
rect 12 49 13 50 
<< pdiffusion >>
rect 13 49 14 50 
<< pdiffusion >>
rect 14 49 15 50 
<< pdiffusion >>
rect 15 49 16 50 
<< pdiffusion >>
rect 16 49 17 50 
<< pdiffusion >>
rect 17 49 18 50 
<< m1 >>
rect 19 49 20 50 
<< pdiffusion >>
rect 30 49 31 50 
<< pdiffusion >>
rect 31 49 32 50 
<< pdiffusion >>
rect 32 49 33 50 
<< pdiffusion >>
rect 33 49 34 50 
<< pdiffusion >>
rect 34 49 35 50 
<< pdiffusion >>
rect 35 49 36 50 
<< pdiffusion >>
rect 48 49 49 50 
<< pdiffusion >>
rect 49 49 50 50 
<< pdiffusion >>
rect 50 49 51 50 
<< pdiffusion >>
rect 51 49 52 50 
<< pdiffusion >>
rect 52 49 53 50 
<< pdiffusion >>
rect 53 49 54 50 
<< m1 >>
rect 64 49 65 50 
<< pdiffusion >>
rect 66 49 67 50 
<< pdiffusion >>
rect 67 49 68 50 
<< pdiffusion >>
rect 68 49 69 50 
<< pdiffusion >>
rect 69 49 70 50 
<< pdiffusion >>
rect 70 49 71 50 
<< pdiffusion >>
rect 71 49 72 50 
<< pdiffusion >>
rect 84 49 85 50 
<< pdiffusion >>
rect 85 49 86 50 
<< pdiffusion >>
rect 86 49 87 50 
<< pdiffusion >>
rect 87 49 88 50 
<< pdiffusion >>
rect 88 49 89 50 
<< pdiffusion >>
rect 89 49 90 50 
<< m1 >>
rect 91 49 92 50 
<< m1 >>
rect 100 49 101 50 
<< pdiffusion >>
rect 102 49 103 50 
<< pdiffusion >>
rect 103 49 104 50 
<< pdiffusion >>
rect 104 49 105 50 
<< pdiffusion >>
rect 105 49 106 50 
<< pdiffusion >>
rect 106 49 107 50 
<< pdiffusion >>
rect 107 49 108 50 
<< m1 >>
rect 109 49 110 50 
<< m1 >>
rect 111 49 112 50 
<< pdiffusion >>
rect 120 49 121 50 
<< pdiffusion >>
rect 121 49 122 50 
<< pdiffusion >>
rect 122 49 123 50 
<< pdiffusion >>
rect 123 49 124 50 
<< pdiffusion >>
rect 124 49 125 50 
<< pdiffusion >>
rect 125 49 126 50 
<< pdiffusion >>
rect 138 49 139 50 
<< pdiffusion >>
rect 139 49 140 50 
<< pdiffusion >>
rect 140 49 141 50 
<< pdiffusion >>
rect 141 49 142 50 
<< pdiffusion >>
rect 142 49 143 50 
<< pdiffusion >>
rect 143 49 144 50 
<< pdiffusion >>
rect 156 49 157 50 
<< pdiffusion >>
rect 157 49 158 50 
<< pdiffusion >>
rect 158 49 159 50 
<< pdiffusion >>
rect 159 49 160 50 
<< pdiffusion >>
rect 160 49 161 50 
<< pdiffusion >>
rect 161 49 162 50 
<< m1 >>
rect 163 49 164 50 
<< m1 >>
rect 165 49 166 50 
<< pdiffusion >>
rect 174 49 175 50 
<< pdiffusion >>
rect 175 49 176 50 
<< pdiffusion >>
rect 176 49 177 50 
<< pdiffusion >>
rect 177 49 178 50 
<< pdiffusion >>
rect 178 49 179 50 
<< pdiffusion >>
rect 179 49 180 50 
<< m1 >>
rect 190 49 191 50 
<< pdiffusion >>
rect 192 49 193 50 
<< pdiffusion >>
rect 193 49 194 50 
<< pdiffusion >>
rect 194 49 195 50 
<< pdiffusion >>
rect 195 49 196 50 
<< pdiffusion >>
rect 196 49 197 50 
<< pdiffusion >>
rect 197 49 198 50 
<< pdiffusion >>
rect 210 49 211 50 
<< pdiffusion >>
rect 211 49 212 50 
<< pdiffusion >>
rect 212 49 213 50 
<< pdiffusion >>
rect 213 49 214 50 
<< pdiffusion >>
rect 214 49 215 50 
<< pdiffusion >>
rect 215 49 216 50 
<< m2 >>
rect 225 49 226 50 
<< m1 >>
rect 226 49 227 50 
<< pdiffusion >>
rect 228 49 229 50 
<< pdiffusion >>
rect 229 49 230 50 
<< pdiffusion >>
rect 230 49 231 50 
<< pdiffusion >>
rect 231 49 232 50 
<< pdiffusion >>
rect 232 49 233 50 
<< pdiffusion >>
rect 233 49 234 50 
<< m1 >>
rect 235 49 236 50 
<< m1 >>
rect 237 49 238 50 
<< m1 >>
rect 244 49 245 50 
<< pdiffusion >>
rect 246 49 247 50 
<< pdiffusion >>
rect 247 49 248 50 
<< pdiffusion >>
rect 248 49 249 50 
<< pdiffusion >>
rect 249 49 250 50 
<< pdiffusion >>
rect 250 49 251 50 
<< pdiffusion >>
rect 251 49 252 50 
<< m1 >>
rect 253 49 254 50 
<< pdiffusion >>
rect 264 49 265 50 
<< pdiffusion >>
rect 265 49 266 50 
<< pdiffusion >>
rect 266 49 267 50 
<< pdiffusion >>
rect 267 49 268 50 
<< pdiffusion >>
rect 268 49 269 50 
<< pdiffusion >>
rect 269 49 270 50 
<< m1 >>
rect 280 49 281 50 
<< pdiffusion >>
rect 282 49 283 50 
<< pdiffusion >>
rect 283 49 284 50 
<< pdiffusion >>
rect 284 49 285 50 
<< pdiffusion >>
rect 285 49 286 50 
<< pdiffusion >>
rect 286 49 287 50 
<< pdiffusion >>
rect 287 49 288 50 
<< m1 >>
rect 289 49 290 50 
<< pdiffusion >>
rect 300 49 301 50 
<< pdiffusion >>
rect 301 49 302 50 
<< pdiffusion >>
rect 302 49 303 50 
<< pdiffusion >>
rect 303 49 304 50 
<< pdiffusion >>
rect 304 49 305 50 
<< pdiffusion >>
rect 305 49 306 50 
<< pdiffusion >>
rect 318 49 319 50 
<< pdiffusion >>
rect 319 49 320 50 
<< pdiffusion >>
rect 320 49 321 50 
<< pdiffusion >>
rect 321 49 322 50 
<< pdiffusion >>
rect 322 49 323 50 
<< pdiffusion >>
rect 323 49 324 50 
<< m1 >>
rect 332 49 333 50 
<< m1 >>
rect 334 49 335 50 
<< pdiffusion >>
rect 336 49 337 50 
<< pdiffusion >>
rect 337 49 338 50 
<< pdiffusion >>
rect 338 49 339 50 
<< pdiffusion >>
rect 339 49 340 50 
<< pdiffusion >>
rect 340 49 341 50 
<< pdiffusion >>
rect 341 49 342 50 
<< pdiffusion >>
rect 354 49 355 50 
<< pdiffusion >>
rect 355 49 356 50 
<< pdiffusion >>
rect 356 49 357 50 
<< pdiffusion >>
rect 357 49 358 50 
<< pdiffusion >>
rect 358 49 359 50 
<< pdiffusion >>
rect 359 49 360 50 
<< pdiffusion >>
rect 372 49 373 50 
<< pdiffusion >>
rect 373 49 374 50 
<< pdiffusion >>
rect 374 49 375 50 
<< pdiffusion >>
rect 375 49 376 50 
<< pdiffusion >>
rect 376 49 377 50 
<< pdiffusion >>
rect 377 49 378 50 
<< m1 >>
rect 388 49 389 50 
<< pdiffusion >>
rect 390 49 391 50 
<< pdiffusion >>
rect 391 49 392 50 
<< pdiffusion >>
rect 392 49 393 50 
<< pdiffusion >>
rect 393 49 394 50 
<< pdiffusion >>
rect 394 49 395 50 
<< pdiffusion >>
rect 395 49 396 50 
<< pdiffusion >>
rect 408 49 409 50 
<< pdiffusion >>
rect 409 49 410 50 
<< pdiffusion >>
rect 410 49 411 50 
<< pdiffusion >>
rect 411 49 412 50 
<< pdiffusion >>
rect 412 49 413 50 
<< pdiffusion >>
rect 413 49 414 50 
<< pdiffusion >>
rect 426 49 427 50 
<< pdiffusion >>
rect 427 49 428 50 
<< pdiffusion >>
rect 428 49 429 50 
<< pdiffusion >>
rect 429 49 430 50 
<< pdiffusion >>
rect 430 49 431 50 
<< pdiffusion >>
rect 431 49 432 50 
<< m1 >>
rect 433 49 434 50 
<< pdiffusion >>
rect 444 49 445 50 
<< pdiffusion >>
rect 445 49 446 50 
<< pdiffusion >>
rect 446 49 447 50 
<< pdiffusion >>
rect 447 49 448 50 
<< pdiffusion >>
rect 448 49 449 50 
<< pdiffusion >>
rect 449 49 450 50 
<< pdiffusion >>
rect 462 49 463 50 
<< pdiffusion >>
rect 463 49 464 50 
<< pdiffusion >>
rect 464 49 465 50 
<< pdiffusion >>
rect 465 49 466 50 
<< pdiffusion >>
rect 466 49 467 50 
<< pdiffusion >>
rect 467 49 468 50 
<< pdiffusion >>
rect 480 49 481 50 
<< pdiffusion >>
rect 481 49 482 50 
<< pdiffusion >>
rect 482 49 483 50 
<< pdiffusion >>
rect 483 49 484 50 
<< pdiffusion >>
rect 484 49 485 50 
<< pdiffusion >>
rect 485 49 486 50 
<< m1 >>
rect 487 49 488 50 
<< pdiffusion >>
rect 498 49 499 50 
<< pdiffusion >>
rect 499 49 500 50 
<< pdiffusion >>
rect 500 49 501 50 
<< pdiffusion >>
rect 501 49 502 50 
<< pdiffusion >>
rect 502 49 503 50 
<< pdiffusion >>
rect 503 49 504 50 
<< m1 >>
rect 505 49 506 50 
<< pdiffusion >>
rect 516 49 517 50 
<< pdiffusion >>
rect 517 49 518 50 
<< pdiffusion >>
rect 518 49 519 50 
<< pdiffusion >>
rect 519 49 520 50 
<< pdiffusion >>
rect 520 49 521 50 
<< pdiffusion >>
rect 521 49 522 50 
<< pdiffusion >>
rect 12 50 13 51 
<< pdiffusion >>
rect 13 50 14 51 
<< pdiffusion >>
rect 14 50 15 51 
<< pdiffusion >>
rect 15 50 16 51 
<< pdiffusion >>
rect 16 50 17 51 
<< pdiffusion >>
rect 17 50 18 51 
<< m1 >>
rect 19 50 20 51 
<< pdiffusion >>
rect 30 50 31 51 
<< pdiffusion >>
rect 31 50 32 51 
<< pdiffusion >>
rect 32 50 33 51 
<< pdiffusion >>
rect 33 50 34 51 
<< pdiffusion >>
rect 34 50 35 51 
<< pdiffusion >>
rect 35 50 36 51 
<< pdiffusion >>
rect 48 50 49 51 
<< pdiffusion >>
rect 49 50 50 51 
<< pdiffusion >>
rect 50 50 51 51 
<< pdiffusion >>
rect 51 50 52 51 
<< pdiffusion >>
rect 52 50 53 51 
<< pdiffusion >>
rect 53 50 54 51 
<< m1 >>
rect 64 50 65 51 
<< pdiffusion >>
rect 66 50 67 51 
<< pdiffusion >>
rect 67 50 68 51 
<< pdiffusion >>
rect 68 50 69 51 
<< pdiffusion >>
rect 69 50 70 51 
<< pdiffusion >>
rect 70 50 71 51 
<< pdiffusion >>
rect 71 50 72 51 
<< pdiffusion >>
rect 84 50 85 51 
<< pdiffusion >>
rect 85 50 86 51 
<< pdiffusion >>
rect 86 50 87 51 
<< pdiffusion >>
rect 87 50 88 51 
<< pdiffusion >>
rect 88 50 89 51 
<< pdiffusion >>
rect 89 50 90 51 
<< m1 >>
rect 91 50 92 51 
<< m1 >>
rect 100 50 101 51 
<< pdiffusion >>
rect 102 50 103 51 
<< pdiffusion >>
rect 103 50 104 51 
<< pdiffusion >>
rect 104 50 105 51 
<< pdiffusion >>
rect 105 50 106 51 
<< pdiffusion >>
rect 106 50 107 51 
<< pdiffusion >>
rect 107 50 108 51 
<< m1 >>
rect 109 50 110 51 
<< m1 >>
rect 111 50 112 51 
<< pdiffusion >>
rect 120 50 121 51 
<< pdiffusion >>
rect 121 50 122 51 
<< pdiffusion >>
rect 122 50 123 51 
<< pdiffusion >>
rect 123 50 124 51 
<< pdiffusion >>
rect 124 50 125 51 
<< pdiffusion >>
rect 125 50 126 51 
<< pdiffusion >>
rect 138 50 139 51 
<< pdiffusion >>
rect 139 50 140 51 
<< pdiffusion >>
rect 140 50 141 51 
<< pdiffusion >>
rect 141 50 142 51 
<< pdiffusion >>
rect 142 50 143 51 
<< pdiffusion >>
rect 143 50 144 51 
<< pdiffusion >>
rect 156 50 157 51 
<< pdiffusion >>
rect 157 50 158 51 
<< pdiffusion >>
rect 158 50 159 51 
<< pdiffusion >>
rect 159 50 160 51 
<< pdiffusion >>
rect 160 50 161 51 
<< pdiffusion >>
rect 161 50 162 51 
<< m1 >>
rect 163 50 164 51 
<< m1 >>
rect 165 50 166 51 
<< pdiffusion >>
rect 174 50 175 51 
<< pdiffusion >>
rect 175 50 176 51 
<< pdiffusion >>
rect 176 50 177 51 
<< pdiffusion >>
rect 177 50 178 51 
<< pdiffusion >>
rect 178 50 179 51 
<< pdiffusion >>
rect 179 50 180 51 
<< m1 >>
rect 190 50 191 51 
<< pdiffusion >>
rect 192 50 193 51 
<< pdiffusion >>
rect 193 50 194 51 
<< pdiffusion >>
rect 194 50 195 51 
<< pdiffusion >>
rect 195 50 196 51 
<< pdiffusion >>
rect 196 50 197 51 
<< pdiffusion >>
rect 197 50 198 51 
<< pdiffusion >>
rect 210 50 211 51 
<< pdiffusion >>
rect 211 50 212 51 
<< pdiffusion >>
rect 212 50 213 51 
<< pdiffusion >>
rect 213 50 214 51 
<< pdiffusion >>
rect 214 50 215 51 
<< pdiffusion >>
rect 215 50 216 51 
<< m2 >>
rect 225 50 226 51 
<< m1 >>
rect 226 50 227 51 
<< pdiffusion >>
rect 228 50 229 51 
<< pdiffusion >>
rect 229 50 230 51 
<< pdiffusion >>
rect 230 50 231 51 
<< pdiffusion >>
rect 231 50 232 51 
<< pdiffusion >>
rect 232 50 233 51 
<< pdiffusion >>
rect 233 50 234 51 
<< m1 >>
rect 235 50 236 51 
<< m1 >>
rect 237 50 238 51 
<< m1 >>
rect 244 50 245 51 
<< pdiffusion >>
rect 246 50 247 51 
<< pdiffusion >>
rect 247 50 248 51 
<< pdiffusion >>
rect 248 50 249 51 
<< pdiffusion >>
rect 249 50 250 51 
<< pdiffusion >>
rect 250 50 251 51 
<< pdiffusion >>
rect 251 50 252 51 
<< m1 >>
rect 253 50 254 51 
<< pdiffusion >>
rect 264 50 265 51 
<< pdiffusion >>
rect 265 50 266 51 
<< pdiffusion >>
rect 266 50 267 51 
<< pdiffusion >>
rect 267 50 268 51 
<< pdiffusion >>
rect 268 50 269 51 
<< pdiffusion >>
rect 269 50 270 51 
<< m1 >>
rect 280 50 281 51 
<< pdiffusion >>
rect 282 50 283 51 
<< pdiffusion >>
rect 283 50 284 51 
<< pdiffusion >>
rect 284 50 285 51 
<< pdiffusion >>
rect 285 50 286 51 
<< pdiffusion >>
rect 286 50 287 51 
<< pdiffusion >>
rect 287 50 288 51 
<< m1 >>
rect 289 50 290 51 
<< pdiffusion >>
rect 300 50 301 51 
<< pdiffusion >>
rect 301 50 302 51 
<< pdiffusion >>
rect 302 50 303 51 
<< pdiffusion >>
rect 303 50 304 51 
<< pdiffusion >>
rect 304 50 305 51 
<< pdiffusion >>
rect 305 50 306 51 
<< pdiffusion >>
rect 318 50 319 51 
<< pdiffusion >>
rect 319 50 320 51 
<< pdiffusion >>
rect 320 50 321 51 
<< pdiffusion >>
rect 321 50 322 51 
<< pdiffusion >>
rect 322 50 323 51 
<< pdiffusion >>
rect 323 50 324 51 
<< m1 >>
rect 332 50 333 51 
<< m1 >>
rect 334 50 335 51 
<< pdiffusion >>
rect 336 50 337 51 
<< pdiffusion >>
rect 337 50 338 51 
<< pdiffusion >>
rect 338 50 339 51 
<< pdiffusion >>
rect 339 50 340 51 
<< pdiffusion >>
rect 340 50 341 51 
<< pdiffusion >>
rect 341 50 342 51 
<< pdiffusion >>
rect 354 50 355 51 
<< pdiffusion >>
rect 355 50 356 51 
<< pdiffusion >>
rect 356 50 357 51 
<< pdiffusion >>
rect 357 50 358 51 
<< pdiffusion >>
rect 358 50 359 51 
<< pdiffusion >>
rect 359 50 360 51 
<< pdiffusion >>
rect 372 50 373 51 
<< pdiffusion >>
rect 373 50 374 51 
<< pdiffusion >>
rect 374 50 375 51 
<< pdiffusion >>
rect 375 50 376 51 
<< pdiffusion >>
rect 376 50 377 51 
<< pdiffusion >>
rect 377 50 378 51 
<< m1 >>
rect 388 50 389 51 
<< pdiffusion >>
rect 390 50 391 51 
<< pdiffusion >>
rect 391 50 392 51 
<< pdiffusion >>
rect 392 50 393 51 
<< pdiffusion >>
rect 393 50 394 51 
<< pdiffusion >>
rect 394 50 395 51 
<< pdiffusion >>
rect 395 50 396 51 
<< pdiffusion >>
rect 408 50 409 51 
<< pdiffusion >>
rect 409 50 410 51 
<< pdiffusion >>
rect 410 50 411 51 
<< pdiffusion >>
rect 411 50 412 51 
<< pdiffusion >>
rect 412 50 413 51 
<< pdiffusion >>
rect 413 50 414 51 
<< pdiffusion >>
rect 426 50 427 51 
<< pdiffusion >>
rect 427 50 428 51 
<< pdiffusion >>
rect 428 50 429 51 
<< pdiffusion >>
rect 429 50 430 51 
<< pdiffusion >>
rect 430 50 431 51 
<< pdiffusion >>
rect 431 50 432 51 
<< m1 >>
rect 433 50 434 51 
<< pdiffusion >>
rect 444 50 445 51 
<< pdiffusion >>
rect 445 50 446 51 
<< pdiffusion >>
rect 446 50 447 51 
<< pdiffusion >>
rect 447 50 448 51 
<< pdiffusion >>
rect 448 50 449 51 
<< pdiffusion >>
rect 449 50 450 51 
<< pdiffusion >>
rect 462 50 463 51 
<< pdiffusion >>
rect 463 50 464 51 
<< pdiffusion >>
rect 464 50 465 51 
<< pdiffusion >>
rect 465 50 466 51 
<< pdiffusion >>
rect 466 50 467 51 
<< pdiffusion >>
rect 467 50 468 51 
<< pdiffusion >>
rect 480 50 481 51 
<< pdiffusion >>
rect 481 50 482 51 
<< pdiffusion >>
rect 482 50 483 51 
<< pdiffusion >>
rect 483 50 484 51 
<< pdiffusion >>
rect 484 50 485 51 
<< pdiffusion >>
rect 485 50 486 51 
<< m1 >>
rect 487 50 488 51 
<< pdiffusion >>
rect 498 50 499 51 
<< pdiffusion >>
rect 499 50 500 51 
<< pdiffusion >>
rect 500 50 501 51 
<< pdiffusion >>
rect 501 50 502 51 
<< pdiffusion >>
rect 502 50 503 51 
<< pdiffusion >>
rect 503 50 504 51 
<< m1 >>
rect 505 50 506 51 
<< pdiffusion >>
rect 516 50 517 51 
<< pdiffusion >>
rect 517 50 518 51 
<< pdiffusion >>
rect 518 50 519 51 
<< pdiffusion >>
rect 519 50 520 51 
<< pdiffusion >>
rect 520 50 521 51 
<< pdiffusion >>
rect 521 50 522 51 
<< pdiffusion >>
rect 12 51 13 52 
<< pdiffusion >>
rect 13 51 14 52 
<< pdiffusion >>
rect 14 51 15 52 
<< pdiffusion >>
rect 15 51 16 52 
<< pdiffusion >>
rect 16 51 17 52 
<< pdiffusion >>
rect 17 51 18 52 
<< m1 >>
rect 19 51 20 52 
<< pdiffusion >>
rect 30 51 31 52 
<< pdiffusion >>
rect 31 51 32 52 
<< pdiffusion >>
rect 32 51 33 52 
<< pdiffusion >>
rect 33 51 34 52 
<< pdiffusion >>
rect 34 51 35 52 
<< pdiffusion >>
rect 35 51 36 52 
<< pdiffusion >>
rect 48 51 49 52 
<< pdiffusion >>
rect 49 51 50 52 
<< pdiffusion >>
rect 50 51 51 52 
<< pdiffusion >>
rect 51 51 52 52 
<< pdiffusion >>
rect 52 51 53 52 
<< pdiffusion >>
rect 53 51 54 52 
<< m1 >>
rect 64 51 65 52 
<< pdiffusion >>
rect 66 51 67 52 
<< pdiffusion >>
rect 67 51 68 52 
<< pdiffusion >>
rect 68 51 69 52 
<< pdiffusion >>
rect 69 51 70 52 
<< pdiffusion >>
rect 70 51 71 52 
<< pdiffusion >>
rect 71 51 72 52 
<< pdiffusion >>
rect 84 51 85 52 
<< pdiffusion >>
rect 85 51 86 52 
<< pdiffusion >>
rect 86 51 87 52 
<< pdiffusion >>
rect 87 51 88 52 
<< pdiffusion >>
rect 88 51 89 52 
<< pdiffusion >>
rect 89 51 90 52 
<< m1 >>
rect 91 51 92 52 
<< m1 >>
rect 100 51 101 52 
<< pdiffusion >>
rect 102 51 103 52 
<< pdiffusion >>
rect 103 51 104 52 
<< pdiffusion >>
rect 104 51 105 52 
<< pdiffusion >>
rect 105 51 106 52 
<< pdiffusion >>
rect 106 51 107 52 
<< pdiffusion >>
rect 107 51 108 52 
<< m1 >>
rect 109 51 110 52 
<< m1 >>
rect 111 51 112 52 
<< pdiffusion >>
rect 120 51 121 52 
<< pdiffusion >>
rect 121 51 122 52 
<< pdiffusion >>
rect 122 51 123 52 
<< pdiffusion >>
rect 123 51 124 52 
<< pdiffusion >>
rect 124 51 125 52 
<< pdiffusion >>
rect 125 51 126 52 
<< pdiffusion >>
rect 138 51 139 52 
<< pdiffusion >>
rect 139 51 140 52 
<< pdiffusion >>
rect 140 51 141 52 
<< pdiffusion >>
rect 141 51 142 52 
<< pdiffusion >>
rect 142 51 143 52 
<< pdiffusion >>
rect 143 51 144 52 
<< pdiffusion >>
rect 156 51 157 52 
<< pdiffusion >>
rect 157 51 158 52 
<< pdiffusion >>
rect 158 51 159 52 
<< pdiffusion >>
rect 159 51 160 52 
<< pdiffusion >>
rect 160 51 161 52 
<< pdiffusion >>
rect 161 51 162 52 
<< m1 >>
rect 163 51 164 52 
<< m1 >>
rect 165 51 166 52 
<< pdiffusion >>
rect 174 51 175 52 
<< pdiffusion >>
rect 175 51 176 52 
<< pdiffusion >>
rect 176 51 177 52 
<< pdiffusion >>
rect 177 51 178 52 
<< pdiffusion >>
rect 178 51 179 52 
<< pdiffusion >>
rect 179 51 180 52 
<< m1 >>
rect 190 51 191 52 
<< pdiffusion >>
rect 192 51 193 52 
<< pdiffusion >>
rect 193 51 194 52 
<< pdiffusion >>
rect 194 51 195 52 
<< pdiffusion >>
rect 195 51 196 52 
<< pdiffusion >>
rect 196 51 197 52 
<< pdiffusion >>
rect 197 51 198 52 
<< pdiffusion >>
rect 210 51 211 52 
<< pdiffusion >>
rect 211 51 212 52 
<< pdiffusion >>
rect 212 51 213 52 
<< pdiffusion >>
rect 213 51 214 52 
<< pdiffusion >>
rect 214 51 215 52 
<< pdiffusion >>
rect 215 51 216 52 
<< m2 >>
rect 225 51 226 52 
<< m1 >>
rect 226 51 227 52 
<< pdiffusion >>
rect 228 51 229 52 
<< pdiffusion >>
rect 229 51 230 52 
<< pdiffusion >>
rect 230 51 231 52 
<< pdiffusion >>
rect 231 51 232 52 
<< pdiffusion >>
rect 232 51 233 52 
<< pdiffusion >>
rect 233 51 234 52 
<< m1 >>
rect 235 51 236 52 
<< m1 >>
rect 237 51 238 52 
<< m1 >>
rect 244 51 245 52 
<< pdiffusion >>
rect 246 51 247 52 
<< pdiffusion >>
rect 247 51 248 52 
<< pdiffusion >>
rect 248 51 249 52 
<< pdiffusion >>
rect 249 51 250 52 
<< pdiffusion >>
rect 250 51 251 52 
<< pdiffusion >>
rect 251 51 252 52 
<< m1 >>
rect 253 51 254 52 
<< pdiffusion >>
rect 264 51 265 52 
<< pdiffusion >>
rect 265 51 266 52 
<< pdiffusion >>
rect 266 51 267 52 
<< pdiffusion >>
rect 267 51 268 52 
<< pdiffusion >>
rect 268 51 269 52 
<< pdiffusion >>
rect 269 51 270 52 
<< m1 >>
rect 280 51 281 52 
<< pdiffusion >>
rect 282 51 283 52 
<< pdiffusion >>
rect 283 51 284 52 
<< pdiffusion >>
rect 284 51 285 52 
<< pdiffusion >>
rect 285 51 286 52 
<< pdiffusion >>
rect 286 51 287 52 
<< pdiffusion >>
rect 287 51 288 52 
<< m1 >>
rect 289 51 290 52 
<< pdiffusion >>
rect 300 51 301 52 
<< pdiffusion >>
rect 301 51 302 52 
<< pdiffusion >>
rect 302 51 303 52 
<< pdiffusion >>
rect 303 51 304 52 
<< pdiffusion >>
rect 304 51 305 52 
<< pdiffusion >>
rect 305 51 306 52 
<< pdiffusion >>
rect 318 51 319 52 
<< pdiffusion >>
rect 319 51 320 52 
<< pdiffusion >>
rect 320 51 321 52 
<< pdiffusion >>
rect 321 51 322 52 
<< pdiffusion >>
rect 322 51 323 52 
<< pdiffusion >>
rect 323 51 324 52 
<< m1 >>
rect 332 51 333 52 
<< m1 >>
rect 334 51 335 52 
<< pdiffusion >>
rect 336 51 337 52 
<< pdiffusion >>
rect 337 51 338 52 
<< pdiffusion >>
rect 338 51 339 52 
<< pdiffusion >>
rect 339 51 340 52 
<< pdiffusion >>
rect 340 51 341 52 
<< pdiffusion >>
rect 341 51 342 52 
<< pdiffusion >>
rect 354 51 355 52 
<< pdiffusion >>
rect 355 51 356 52 
<< pdiffusion >>
rect 356 51 357 52 
<< pdiffusion >>
rect 357 51 358 52 
<< pdiffusion >>
rect 358 51 359 52 
<< pdiffusion >>
rect 359 51 360 52 
<< pdiffusion >>
rect 372 51 373 52 
<< pdiffusion >>
rect 373 51 374 52 
<< pdiffusion >>
rect 374 51 375 52 
<< pdiffusion >>
rect 375 51 376 52 
<< pdiffusion >>
rect 376 51 377 52 
<< pdiffusion >>
rect 377 51 378 52 
<< m1 >>
rect 388 51 389 52 
<< pdiffusion >>
rect 390 51 391 52 
<< pdiffusion >>
rect 391 51 392 52 
<< pdiffusion >>
rect 392 51 393 52 
<< pdiffusion >>
rect 393 51 394 52 
<< pdiffusion >>
rect 394 51 395 52 
<< pdiffusion >>
rect 395 51 396 52 
<< pdiffusion >>
rect 408 51 409 52 
<< pdiffusion >>
rect 409 51 410 52 
<< pdiffusion >>
rect 410 51 411 52 
<< pdiffusion >>
rect 411 51 412 52 
<< pdiffusion >>
rect 412 51 413 52 
<< pdiffusion >>
rect 413 51 414 52 
<< pdiffusion >>
rect 426 51 427 52 
<< pdiffusion >>
rect 427 51 428 52 
<< pdiffusion >>
rect 428 51 429 52 
<< pdiffusion >>
rect 429 51 430 52 
<< pdiffusion >>
rect 430 51 431 52 
<< pdiffusion >>
rect 431 51 432 52 
<< m1 >>
rect 433 51 434 52 
<< pdiffusion >>
rect 444 51 445 52 
<< pdiffusion >>
rect 445 51 446 52 
<< pdiffusion >>
rect 446 51 447 52 
<< pdiffusion >>
rect 447 51 448 52 
<< pdiffusion >>
rect 448 51 449 52 
<< pdiffusion >>
rect 449 51 450 52 
<< pdiffusion >>
rect 462 51 463 52 
<< pdiffusion >>
rect 463 51 464 52 
<< pdiffusion >>
rect 464 51 465 52 
<< pdiffusion >>
rect 465 51 466 52 
<< pdiffusion >>
rect 466 51 467 52 
<< pdiffusion >>
rect 467 51 468 52 
<< pdiffusion >>
rect 480 51 481 52 
<< pdiffusion >>
rect 481 51 482 52 
<< pdiffusion >>
rect 482 51 483 52 
<< pdiffusion >>
rect 483 51 484 52 
<< pdiffusion >>
rect 484 51 485 52 
<< pdiffusion >>
rect 485 51 486 52 
<< m1 >>
rect 487 51 488 52 
<< pdiffusion >>
rect 498 51 499 52 
<< pdiffusion >>
rect 499 51 500 52 
<< pdiffusion >>
rect 500 51 501 52 
<< pdiffusion >>
rect 501 51 502 52 
<< pdiffusion >>
rect 502 51 503 52 
<< pdiffusion >>
rect 503 51 504 52 
<< m1 >>
rect 505 51 506 52 
<< pdiffusion >>
rect 516 51 517 52 
<< pdiffusion >>
rect 517 51 518 52 
<< pdiffusion >>
rect 518 51 519 52 
<< pdiffusion >>
rect 519 51 520 52 
<< pdiffusion >>
rect 520 51 521 52 
<< pdiffusion >>
rect 521 51 522 52 
<< pdiffusion >>
rect 12 52 13 53 
<< pdiffusion >>
rect 13 52 14 53 
<< pdiffusion >>
rect 14 52 15 53 
<< pdiffusion >>
rect 15 52 16 53 
<< pdiffusion >>
rect 16 52 17 53 
<< pdiffusion >>
rect 17 52 18 53 
<< m1 >>
rect 19 52 20 53 
<< pdiffusion >>
rect 30 52 31 53 
<< pdiffusion >>
rect 31 52 32 53 
<< pdiffusion >>
rect 32 52 33 53 
<< pdiffusion >>
rect 33 52 34 53 
<< pdiffusion >>
rect 34 52 35 53 
<< pdiffusion >>
rect 35 52 36 53 
<< pdiffusion >>
rect 48 52 49 53 
<< pdiffusion >>
rect 49 52 50 53 
<< pdiffusion >>
rect 50 52 51 53 
<< pdiffusion >>
rect 51 52 52 53 
<< pdiffusion >>
rect 52 52 53 53 
<< pdiffusion >>
rect 53 52 54 53 
<< m1 >>
rect 64 52 65 53 
<< pdiffusion >>
rect 66 52 67 53 
<< pdiffusion >>
rect 67 52 68 53 
<< pdiffusion >>
rect 68 52 69 53 
<< pdiffusion >>
rect 69 52 70 53 
<< pdiffusion >>
rect 70 52 71 53 
<< pdiffusion >>
rect 71 52 72 53 
<< pdiffusion >>
rect 84 52 85 53 
<< pdiffusion >>
rect 85 52 86 53 
<< pdiffusion >>
rect 86 52 87 53 
<< pdiffusion >>
rect 87 52 88 53 
<< pdiffusion >>
rect 88 52 89 53 
<< pdiffusion >>
rect 89 52 90 53 
<< m1 >>
rect 91 52 92 53 
<< m1 >>
rect 100 52 101 53 
<< pdiffusion >>
rect 102 52 103 53 
<< pdiffusion >>
rect 103 52 104 53 
<< pdiffusion >>
rect 104 52 105 53 
<< pdiffusion >>
rect 105 52 106 53 
<< pdiffusion >>
rect 106 52 107 53 
<< pdiffusion >>
rect 107 52 108 53 
<< m1 >>
rect 109 52 110 53 
<< m1 >>
rect 111 52 112 53 
<< pdiffusion >>
rect 120 52 121 53 
<< pdiffusion >>
rect 121 52 122 53 
<< pdiffusion >>
rect 122 52 123 53 
<< pdiffusion >>
rect 123 52 124 53 
<< pdiffusion >>
rect 124 52 125 53 
<< pdiffusion >>
rect 125 52 126 53 
<< pdiffusion >>
rect 138 52 139 53 
<< pdiffusion >>
rect 139 52 140 53 
<< pdiffusion >>
rect 140 52 141 53 
<< pdiffusion >>
rect 141 52 142 53 
<< pdiffusion >>
rect 142 52 143 53 
<< pdiffusion >>
rect 143 52 144 53 
<< pdiffusion >>
rect 156 52 157 53 
<< pdiffusion >>
rect 157 52 158 53 
<< pdiffusion >>
rect 158 52 159 53 
<< pdiffusion >>
rect 159 52 160 53 
<< pdiffusion >>
rect 160 52 161 53 
<< pdiffusion >>
rect 161 52 162 53 
<< m1 >>
rect 163 52 164 53 
<< m1 >>
rect 165 52 166 53 
<< pdiffusion >>
rect 174 52 175 53 
<< pdiffusion >>
rect 175 52 176 53 
<< pdiffusion >>
rect 176 52 177 53 
<< pdiffusion >>
rect 177 52 178 53 
<< pdiffusion >>
rect 178 52 179 53 
<< pdiffusion >>
rect 179 52 180 53 
<< m1 >>
rect 190 52 191 53 
<< pdiffusion >>
rect 192 52 193 53 
<< pdiffusion >>
rect 193 52 194 53 
<< pdiffusion >>
rect 194 52 195 53 
<< pdiffusion >>
rect 195 52 196 53 
<< pdiffusion >>
rect 196 52 197 53 
<< pdiffusion >>
rect 197 52 198 53 
<< pdiffusion >>
rect 210 52 211 53 
<< pdiffusion >>
rect 211 52 212 53 
<< pdiffusion >>
rect 212 52 213 53 
<< pdiffusion >>
rect 213 52 214 53 
<< pdiffusion >>
rect 214 52 215 53 
<< pdiffusion >>
rect 215 52 216 53 
<< m2 >>
rect 225 52 226 53 
<< m1 >>
rect 226 52 227 53 
<< pdiffusion >>
rect 228 52 229 53 
<< pdiffusion >>
rect 229 52 230 53 
<< pdiffusion >>
rect 230 52 231 53 
<< pdiffusion >>
rect 231 52 232 53 
<< pdiffusion >>
rect 232 52 233 53 
<< pdiffusion >>
rect 233 52 234 53 
<< m1 >>
rect 235 52 236 53 
<< m1 >>
rect 237 52 238 53 
<< m1 >>
rect 244 52 245 53 
<< pdiffusion >>
rect 246 52 247 53 
<< pdiffusion >>
rect 247 52 248 53 
<< pdiffusion >>
rect 248 52 249 53 
<< pdiffusion >>
rect 249 52 250 53 
<< pdiffusion >>
rect 250 52 251 53 
<< pdiffusion >>
rect 251 52 252 53 
<< m1 >>
rect 253 52 254 53 
<< pdiffusion >>
rect 264 52 265 53 
<< pdiffusion >>
rect 265 52 266 53 
<< pdiffusion >>
rect 266 52 267 53 
<< pdiffusion >>
rect 267 52 268 53 
<< pdiffusion >>
rect 268 52 269 53 
<< pdiffusion >>
rect 269 52 270 53 
<< m1 >>
rect 280 52 281 53 
<< pdiffusion >>
rect 282 52 283 53 
<< pdiffusion >>
rect 283 52 284 53 
<< pdiffusion >>
rect 284 52 285 53 
<< pdiffusion >>
rect 285 52 286 53 
<< pdiffusion >>
rect 286 52 287 53 
<< pdiffusion >>
rect 287 52 288 53 
<< m1 >>
rect 289 52 290 53 
<< pdiffusion >>
rect 300 52 301 53 
<< pdiffusion >>
rect 301 52 302 53 
<< pdiffusion >>
rect 302 52 303 53 
<< pdiffusion >>
rect 303 52 304 53 
<< pdiffusion >>
rect 304 52 305 53 
<< pdiffusion >>
rect 305 52 306 53 
<< pdiffusion >>
rect 318 52 319 53 
<< pdiffusion >>
rect 319 52 320 53 
<< pdiffusion >>
rect 320 52 321 53 
<< pdiffusion >>
rect 321 52 322 53 
<< pdiffusion >>
rect 322 52 323 53 
<< pdiffusion >>
rect 323 52 324 53 
<< m1 >>
rect 332 52 333 53 
<< m1 >>
rect 334 52 335 53 
<< pdiffusion >>
rect 336 52 337 53 
<< pdiffusion >>
rect 337 52 338 53 
<< pdiffusion >>
rect 338 52 339 53 
<< pdiffusion >>
rect 339 52 340 53 
<< pdiffusion >>
rect 340 52 341 53 
<< pdiffusion >>
rect 341 52 342 53 
<< pdiffusion >>
rect 354 52 355 53 
<< pdiffusion >>
rect 355 52 356 53 
<< pdiffusion >>
rect 356 52 357 53 
<< pdiffusion >>
rect 357 52 358 53 
<< pdiffusion >>
rect 358 52 359 53 
<< pdiffusion >>
rect 359 52 360 53 
<< pdiffusion >>
rect 372 52 373 53 
<< pdiffusion >>
rect 373 52 374 53 
<< pdiffusion >>
rect 374 52 375 53 
<< pdiffusion >>
rect 375 52 376 53 
<< pdiffusion >>
rect 376 52 377 53 
<< pdiffusion >>
rect 377 52 378 53 
<< m1 >>
rect 388 52 389 53 
<< pdiffusion >>
rect 390 52 391 53 
<< pdiffusion >>
rect 391 52 392 53 
<< pdiffusion >>
rect 392 52 393 53 
<< pdiffusion >>
rect 393 52 394 53 
<< pdiffusion >>
rect 394 52 395 53 
<< pdiffusion >>
rect 395 52 396 53 
<< pdiffusion >>
rect 408 52 409 53 
<< pdiffusion >>
rect 409 52 410 53 
<< pdiffusion >>
rect 410 52 411 53 
<< pdiffusion >>
rect 411 52 412 53 
<< pdiffusion >>
rect 412 52 413 53 
<< pdiffusion >>
rect 413 52 414 53 
<< pdiffusion >>
rect 426 52 427 53 
<< pdiffusion >>
rect 427 52 428 53 
<< pdiffusion >>
rect 428 52 429 53 
<< pdiffusion >>
rect 429 52 430 53 
<< pdiffusion >>
rect 430 52 431 53 
<< pdiffusion >>
rect 431 52 432 53 
<< m1 >>
rect 433 52 434 53 
<< pdiffusion >>
rect 444 52 445 53 
<< pdiffusion >>
rect 445 52 446 53 
<< pdiffusion >>
rect 446 52 447 53 
<< pdiffusion >>
rect 447 52 448 53 
<< pdiffusion >>
rect 448 52 449 53 
<< pdiffusion >>
rect 449 52 450 53 
<< pdiffusion >>
rect 462 52 463 53 
<< pdiffusion >>
rect 463 52 464 53 
<< pdiffusion >>
rect 464 52 465 53 
<< pdiffusion >>
rect 465 52 466 53 
<< pdiffusion >>
rect 466 52 467 53 
<< pdiffusion >>
rect 467 52 468 53 
<< pdiffusion >>
rect 480 52 481 53 
<< pdiffusion >>
rect 481 52 482 53 
<< pdiffusion >>
rect 482 52 483 53 
<< pdiffusion >>
rect 483 52 484 53 
<< pdiffusion >>
rect 484 52 485 53 
<< pdiffusion >>
rect 485 52 486 53 
<< m1 >>
rect 487 52 488 53 
<< pdiffusion >>
rect 498 52 499 53 
<< pdiffusion >>
rect 499 52 500 53 
<< pdiffusion >>
rect 500 52 501 53 
<< pdiffusion >>
rect 501 52 502 53 
<< pdiffusion >>
rect 502 52 503 53 
<< pdiffusion >>
rect 503 52 504 53 
<< m1 >>
rect 505 52 506 53 
<< pdiffusion >>
rect 516 52 517 53 
<< pdiffusion >>
rect 517 52 518 53 
<< pdiffusion >>
rect 518 52 519 53 
<< pdiffusion >>
rect 519 52 520 53 
<< pdiffusion >>
rect 520 52 521 53 
<< pdiffusion >>
rect 521 52 522 53 
<< pdiffusion >>
rect 12 53 13 54 
<< pdiffusion >>
rect 13 53 14 54 
<< pdiffusion >>
rect 14 53 15 54 
<< pdiffusion >>
rect 15 53 16 54 
<< m1 >>
rect 16 53 17 54 
<< pdiffusion >>
rect 16 53 17 54 
<< pdiffusion >>
rect 17 53 18 54 
<< m1 >>
rect 19 53 20 54 
<< pdiffusion >>
rect 30 53 31 54 
<< pdiffusion >>
rect 31 53 32 54 
<< pdiffusion >>
rect 32 53 33 54 
<< pdiffusion >>
rect 33 53 34 54 
<< pdiffusion >>
rect 34 53 35 54 
<< pdiffusion >>
rect 35 53 36 54 
<< pdiffusion >>
rect 48 53 49 54 
<< pdiffusion >>
rect 49 53 50 54 
<< pdiffusion >>
rect 50 53 51 54 
<< pdiffusion >>
rect 51 53 52 54 
<< pdiffusion >>
rect 52 53 53 54 
<< pdiffusion >>
rect 53 53 54 54 
<< m1 >>
rect 64 53 65 54 
<< pdiffusion >>
rect 66 53 67 54 
<< pdiffusion >>
rect 67 53 68 54 
<< pdiffusion >>
rect 68 53 69 54 
<< pdiffusion >>
rect 69 53 70 54 
<< pdiffusion >>
rect 70 53 71 54 
<< pdiffusion >>
rect 71 53 72 54 
<< pdiffusion >>
rect 84 53 85 54 
<< m1 >>
rect 85 53 86 54 
<< pdiffusion >>
rect 85 53 86 54 
<< pdiffusion >>
rect 86 53 87 54 
<< pdiffusion >>
rect 87 53 88 54 
<< pdiffusion >>
rect 88 53 89 54 
<< pdiffusion >>
rect 89 53 90 54 
<< m1 >>
rect 91 53 92 54 
<< m1 >>
rect 100 53 101 54 
<< pdiffusion >>
rect 102 53 103 54 
<< pdiffusion >>
rect 103 53 104 54 
<< pdiffusion >>
rect 104 53 105 54 
<< pdiffusion >>
rect 105 53 106 54 
<< pdiffusion >>
rect 106 53 107 54 
<< pdiffusion >>
rect 107 53 108 54 
<< m1 >>
rect 109 53 110 54 
<< m1 >>
rect 111 53 112 54 
<< pdiffusion >>
rect 120 53 121 54 
<< pdiffusion >>
rect 121 53 122 54 
<< pdiffusion >>
rect 122 53 123 54 
<< pdiffusion >>
rect 123 53 124 54 
<< pdiffusion >>
rect 124 53 125 54 
<< pdiffusion >>
rect 125 53 126 54 
<< pdiffusion >>
rect 138 53 139 54 
<< pdiffusion >>
rect 139 53 140 54 
<< pdiffusion >>
rect 140 53 141 54 
<< pdiffusion >>
rect 141 53 142 54 
<< pdiffusion >>
rect 142 53 143 54 
<< pdiffusion >>
rect 143 53 144 54 
<< pdiffusion >>
rect 156 53 157 54 
<< pdiffusion >>
rect 157 53 158 54 
<< pdiffusion >>
rect 158 53 159 54 
<< pdiffusion >>
rect 159 53 160 54 
<< pdiffusion >>
rect 160 53 161 54 
<< pdiffusion >>
rect 161 53 162 54 
<< m1 >>
rect 163 53 164 54 
<< m1 >>
rect 165 53 166 54 
<< pdiffusion >>
rect 174 53 175 54 
<< pdiffusion >>
rect 175 53 176 54 
<< pdiffusion >>
rect 176 53 177 54 
<< pdiffusion >>
rect 177 53 178 54 
<< pdiffusion >>
rect 178 53 179 54 
<< pdiffusion >>
rect 179 53 180 54 
<< m1 >>
rect 190 53 191 54 
<< pdiffusion >>
rect 192 53 193 54 
<< pdiffusion >>
rect 193 53 194 54 
<< pdiffusion >>
rect 194 53 195 54 
<< pdiffusion >>
rect 195 53 196 54 
<< pdiffusion >>
rect 196 53 197 54 
<< pdiffusion >>
rect 197 53 198 54 
<< pdiffusion >>
rect 210 53 211 54 
<< pdiffusion >>
rect 211 53 212 54 
<< pdiffusion >>
rect 212 53 213 54 
<< pdiffusion >>
rect 213 53 214 54 
<< pdiffusion >>
rect 214 53 215 54 
<< pdiffusion >>
rect 215 53 216 54 
<< m2 >>
rect 225 53 226 54 
<< m1 >>
rect 226 53 227 54 
<< pdiffusion >>
rect 228 53 229 54 
<< m1 >>
rect 229 53 230 54 
<< pdiffusion >>
rect 229 53 230 54 
<< pdiffusion >>
rect 230 53 231 54 
<< pdiffusion >>
rect 231 53 232 54 
<< m1 >>
rect 232 53 233 54 
<< pdiffusion >>
rect 232 53 233 54 
<< pdiffusion >>
rect 233 53 234 54 
<< m1 >>
rect 235 53 236 54 
<< m1 >>
rect 237 53 238 54 
<< m1 >>
rect 244 53 245 54 
<< pdiffusion >>
rect 246 53 247 54 
<< pdiffusion >>
rect 247 53 248 54 
<< pdiffusion >>
rect 248 53 249 54 
<< pdiffusion >>
rect 249 53 250 54 
<< pdiffusion >>
rect 250 53 251 54 
<< pdiffusion >>
rect 251 53 252 54 
<< m1 >>
rect 253 53 254 54 
<< pdiffusion >>
rect 264 53 265 54 
<< m1 >>
rect 265 53 266 54 
<< pdiffusion >>
rect 265 53 266 54 
<< pdiffusion >>
rect 266 53 267 54 
<< pdiffusion >>
rect 267 53 268 54 
<< m1 >>
rect 268 53 269 54 
<< pdiffusion >>
rect 268 53 269 54 
<< pdiffusion >>
rect 269 53 270 54 
<< m1 >>
rect 280 53 281 54 
<< pdiffusion >>
rect 282 53 283 54 
<< pdiffusion >>
rect 283 53 284 54 
<< pdiffusion >>
rect 284 53 285 54 
<< pdiffusion >>
rect 285 53 286 54 
<< pdiffusion >>
rect 286 53 287 54 
<< pdiffusion >>
rect 287 53 288 54 
<< m1 >>
rect 289 53 290 54 
<< pdiffusion >>
rect 300 53 301 54 
<< pdiffusion >>
rect 301 53 302 54 
<< pdiffusion >>
rect 302 53 303 54 
<< pdiffusion >>
rect 303 53 304 54 
<< pdiffusion >>
rect 304 53 305 54 
<< pdiffusion >>
rect 305 53 306 54 
<< pdiffusion >>
rect 318 53 319 54 
<< pdiffusion >>
rect 319 53 320 54 
<< pdiffusion >>
rect 320 53 321 54 
<< pdiffusion >>
rect 321 53 322 54 
<< pdiffusion >>
rect 322 53 323 54 
<< pdiffusion >>
rect 323 53 324 54 
<< m1 >>
rect 332 53 333 54 
<< m1 >>
rect 334 53 335 54 
<< pdiffusion >>
rect 336 53 337 54 
<< pdiffusion >>
rect 337 53 338 54 
<< pdiffusion >>
rect 338 53 339 54 
<< pdiffusion >>
rect 339 53 340 54 
<< pdiffusion >>
rect 340 53 341 54 
<< pdiffusion >>
rect 341 53 342 54 
<< pdiffusion >>
rect 354 53 355 54 
<< pdiffusion >>
rect 355 53 356 54 
<< pdiffusion >>
rect 356 53 357 54 
<< pdiffusion >>
rect 357 53 358 54 
<< pdiffusion >>
rect 358 53 359 54 
<< pdiffusion >>
rect 359 53 360 54 
<< pdiffusion >>
rect 372 53 373 54 
<< pdiffusion >>
rect 373 53 374 54 
<< pdiffusion >>
rect 374 53 375 54 
<< pdiffusion >>
rect 375 53 376 54 
<< pdiffusion >>
rect 376 53 377 54 
<< pdiffusion >>
rect 377 53 378 54 
<< m1 >>
rect 388 53 389 54 
<< pdiffusion >>
rect 390 53 391 54 
<< pdiffusion >>
rect 391 53 392 54 
<< pdiffusion >>
rect 392 53 393 54 
<< pdiffusion >>
rect 393 53 394 54 
<< pdiffusion >>
rect 394 53 395 54 
<< pdiffusion >>
rect 395 53 396 54 
<< pdiffusion >>
rect 408 53 409 54 
<< pdiffusion >>
rect 409 53 410 54 
<< pdiffusion >>
rect 410 53 411 54 
<< pdiffusion >>
rect 411 53 412 54 
<< pdiffusion >>
rect 412 53 413 54 
<< pdiffusion >>
rect 413 53 414 54 
<< pdiffusion >>
rect 426 53 427 54 
<< pdiffusion >>
rect 427 53 428 54 
<< pdiffusion >>
rect 428 53 429 54 
<< pdiffusion >>
rect 429 53 430 54 
<< pdiffusion >>
rect 430 53 431 54 
<< pdiffusion >>
rect 431 53 432 54 
<< m1 >>
rect 433 53 434 54 
<< pdiffusion >>
rect 444 53 445 54 
<< pdiffusion >>
rect 445 53 446 54 
<< pdiffusion >>
rect 446 53 447 54 
<< pdiffusion >>
rect 447 53 448 54 
<< pdiffusion >>
rect 448 53 449 54 
<< pdiffusion >>
rect 449 53 450 54 
<< pdiffusion >>
rect 462 53 463 54 
<< pdiffusion >>
rect 463 53 464 54 
<< pdiffusion >>
rect 464 53 465 54 
<< pdiffusion >>
rect 465 53 466 54 
<< pdiffusion >>
rect 466 53 467 54 
<< pdiffusion >>
rect 467 53 468 54 
<< pdiffusion >>
rect 480 53 481 54 
<< pdiffusion >>
rect 481 53 482 54 
<< pdiffusion >>
rect 482 53 483 54 
<< pdiffusion >>
rect 483 53 484 54 
<< pdiffusion >>
rect 484 53 485 54 
<< pdiffusion >>
rect 485 53 486 54 
<< m1 >>
rect 487 53 488 54 
<< pdiffusion >>
rect 498 53 499 54 
<< m1 >>
rect 499 53 500 54 
<< pdiffusion >>
rect 499 53 500 54 
<< pdiffusion >>
rect 500 53 501 54 
<< pdiffusion >>
rect 501 53 502 54 
<< pdiffusion >>
rect 502 53 503 54 
<< pdiffusion >>
rect 503 53 504 54 
<< m1 >>
rect 505 53 506 54 
<< pdiffusion >>
rect 516 53 517 54 
<< pdiffusion >>
rect 517 53 518 54 
<< pdiffusion >>
rect 518 53 519 54 
<< pdiffusion >>
rect 519 53 520 54 
<< pdiffusion >>
rect 520 53 521 54 
<< pdiffusion >>
rect 521 53 522 54 
<< m1 >>
rect 16 54 17 55 
<< m1 >>
rect 19 54 20 55 
<< m1 >>
rect 64 54 65 55 
<< m1 >>
rect 85 54 86 55 
<< m1 >>
rect 91 54 92 55 
<< m1 >>
rect 100 54 101 55 
<< m1 >>
rect 109 54 110 55 
<< m1 >>
rect 111 54 112 55 
<< m1 >>
rect 163 54 164 55 
<< m1 >>
rect 165 54 166 55 
<< m1 >>
rect 190 54 191 55 
<< m2 >>
rect 225 54 226 55 
<< m1 >>
rect 226 54 227 55 
<< m1 >>
rect 229 54 230 55 
<< m1 >>
rect 232 54 233 55 
<< m1 >>
rect 235 54 236 55 
<< m1 >>
rect 237 54 238 55 
<< m1 >>
rect 244 54 245 55 
<< m1 >>
rect 253 54 254 55 
<< m1 >>
rect 265 54 266 55 
<< m1 >>
rect 268 54 269 55 
<< m1 >>
rect 280 54 281 55 
<< m1 >>
rect 289 54 290 55 
<< m1 >>
rect 332 54 333 55 
<< m1 >>
rect 334 54 335 55 
<< m1 >>
rect 388 54 389 55 
<< m1 >>
rect 433 54 434 55 
<< m1 >>
rect 487 54 488 55 
<< m1 >>
rect 499 54 500 55 
<< m1 >>
rect 505 54 506 55 
<< m1 >>
rect 16 55 17 56 
<< m1 >>
rect 17 55 18 56 
<< m1 >>
rect 18 55 19 56 
<< m1 >>
rect 19 55 20 56 
<< m1 >>
rect 64 55 65 56 
<< m1 >>
rect 85 55 86 56 
<< m1 >>
rect 91 55 92 56 
<< m1 >>
rect 100 55 101 56 
<< m1 >>
rect 109 55 110 56 
<< m1 >>
rect 111 55 112 56 
<< m1 >>
rect 163 55 164 56 
<< m1 >>
rect 165 55 166 56 
<< m1 >>
rect 190 55 191 56 
<< m2 >>
rect 225 55 226 56 
<< m1 >>
rect 226 55 227 56 
<< m1 >>
rect 229 55 230 56 
<< m1 >>
rect 232 55 233 56 
<< m1 >>
rect 233 55 234 56 
<< m1 >>
rect 234 55 235 56 
<< m1 >>
rect 235 55 236 56 
<< m1 >>
rect 237 55 238 56 
<< m1 >>
rect 244 55 245 56 
<< m1 >>
rect 253 55 254 56 
<< m1 >>
rect 265 55 266 56 
<< m1 >>
rect 268 55 269 56 
<< m1 >>
rect 280 55 281 56 
<< m1 >>
rect 289 55 290 56 
<< m1 >>
rect 332 55 333 56 
<< m1 >>
rect 334 55 335 56 
<< m1 >>
rect 388 55 389 56 
<< m1 >>
rect 433 55 434 56 
<< m1 >>
rect 487 55 488 56 
<< m1 >>
rect 499 55 500 56 
<< m1 >>
rect 505 55 506 56 
<< m1 >>
rect 64 56 65 57 
<< m1 >>
rect 85 56 86 57 
<< m1 >>
rect 91 56 92 57 
<< m1 >>
rect 100 56 101 57 
<< m1 >>
rect 109 56 110 57 
<< m1 >>
rect 111 56 112 57 
<< m1 >>
rect 163 56 164 57 
<< m1 >>
rect 165 56 166 57 
<< m1 >>
rect 190 56 191 57 
<< m2 >>
rect 225 56 226 57 
<< m1 >>
rect 226 56 227 57 
<< m1 >>
rect 229 56 230 57 
<< m1 >>
rect 237 56 238 57 
<< m1 >>
rect 244 56 245 57 
<< m1 >>
rect 253 56 254 57 
<< m1 >>
rect 265 56 266 57 
<< m1 >>
rect 268 56 269 57 
<< m1 >>
rect 280 56 281 57 
<< m1 >>
rect 289 56 290 57 
<< m1 >>
rect 332 56 333 57 
<< m1 >>
rect 334 56 335 57 
<< m1 >>
rect 388 56 389 57 
<< m1 >>
rect 433 56 434 57 
<< m1 >>
rect 487 56 488 57 
<< m1 >>
rect 499 56 500 57 
<< m1 >>
rect 500 56 501 57 
<< m1 >>
rect 501 56 502 57 
<< m1 >>
rect 502 56 503 57 
<< m1 >>
rect 503 56 504 57 
<< m1 >>
rect 504 56 505 57 
<< m1 >>
rect 505 56 506 57 
<< m1 >>
rect 64 57 65 58 
<< m1 >>
rect 85 57 86 58 
<< m1 >>
rect 91 57 92 58 
<< m1 >>
rect 100 57 101 58 
<< m1 >>
rect 109 57 110 58 
<< m1 >>
rect 111 57 112 58 
<< m1 >>
rect 158 57 159 58 
<< m1 >>
rect 159 57 160 58 
<< m1 >>
rect 160 57 161 58 
<< m1 >>
rect 161 57 162 58 
<< m2 >>
rect 161 57 162 58 
<< m2c >>
rect 161 57 162 58 
<< m1 >>
rect 161 57 162 58 
<< m2 >>
rect 161 57 162 58 
<< m2 >>
rect 162 57 163 58 
<< m1 >>
rect 163 57 164 58 
<< m2 >>
rect 163 57 164 58 
<< m2 >>
rect 164 57 165 58 
<< m1 >>
rect 165 57 166 58 
<< m2 >>
rect 165 57 166 58 
<< m2c >>
rect 165 57 166 58 
<< m1 >>
rect 165 57 166 58 
<< m2 >>
rect 165 57 166 58 
<< m1 >>
rect 190 57 191 58 
<< m2 >>
rect 225 57 226 58 
<< m1 >>
rect 226 57 227 58 
<< m1 >>
rect 229 57 230 58 
<< m1 >>
rect 237 57 238 58 
<< m2 >>
rect 237 57 238 58 
<< m2c >>
rect 237 57 238 58 
<< m1 >>
rect 237 57 238 58 
<< m2 >>
rect 237 57 238 58 
<< m1 >>
rect 244 57 245 58 
<< m2 >>
rect 244 57 245 58 
<< m2c >>
rect 244 57 245 58 
<< m1 >>
rect 244 57 245 58 
<< m2 >>
rect 244 57 245 58 
<< m1 >>
rect 248 57 249 58 
<< m1 >>
rect 249 57 250 58 
<< m1 >>
rect 250 57 251 58 
<< m1 >>
rect 251 57 252 58 
<< m2 >>
rect 251 57 252 58 
<< m2c >>
rect 251 57 252 58 
<< m1 >>
rect 251 57 252 58 
<< m2 >>
rect 251 57 252 58 
<< m2 >>
rect 252 57 253 58 
<< m1 >>
rect 253 57 254 58 
<< m2 >>
rect 253 57 254 58 
<< m2 >>
rect 254 57 255 58 
<< m1 >>
rect 255 57 256 58 
<< m2 >>
rect 255 57 256 58 
<< m2c >>
rect 255 57 256 58 
<< m1 >>
rect 255 57 256 58 
<< m2 >>
rect 255 57 256 58 
<< m1 >>
rect 256 57 257 58 
<< m1 >>
rect 257 57 258 58 
<< m1 >>
rect 258 57 259 58 
<< m1 >>
rect 259 57 260 58 
<< m1 >>
rect 260 57 261 58 
<< m1 >>
rect 261 57 262 58 
<< m1 >>
rect 262 57 263 58 
<< m1 >>
rect 263 57 264 58 
<< m1 >>
rect 264 57 265 58 
<< m1 >>
rect 265 57 266 58 
<< m1 >>
rect 268 57 269 58 
<< m2 >>
rect 269 57 270 58 
<< m1 >>
rect 270 57 271 58 
<< m2 >>
rect 270 57 271 58 
<< m2c >>
rect 270 57 271 58 
<< m1 >>
rect 270 57 271 58 
<< m2 >>
rect 270 57 271 58 
<< m1 >>
rect 271 57 272 58 
<< m1 >>
rect 272 57 273 58 
<< m1 >>
rect 273 57 274 58 
<< m1 >>
rect 274 57 275 58 
<< m1 >>
rect 275 57 276 58 
<< m1 >>
rect 276 57 277 58 
<< m1 >>
rect 277 57 278 58 
<< m1 >>
rect 278 57 279 58 
<< m2 >>
rect 278 57 279 58 
<< m2c >>
rect 278 57 279 58 
<< m1 >>
rect 278 57 279 58 
<< m2 >>
rect 278 57 279 58 
<< m2 >>
rect 279 57 280 58 
<< m1 >>
rect 280 57 281 58 
<< m2 >>
rect 280 57 281 58 
<< m2 >>
rect 281 57 282 58 
<< m1 >>
rect 282 57 283 58 
<< m2 >>
rect 282 57 283 58 
<< m2c >>
rect 282 57 283 58 
<< m1 >>
rect 282 57 283 58 
<< m2 >>
rect 282 57 283 58 
<< m1 >>
rect 289 57 290 58 
<< m1 >>
rect 330 57 331 58 
<< m2 >>
rect 330 57 331 58 
<< m2c >>
rect 330 57 331 58 
<< m1 >>
rect 330 57 331 58 
<< m2 >>
rect 330 57 331 58 
<< m2 >>
rect 331 57 332 58 
<< m1 >>
rect 332 57 333 58 
<< m2 >>
rect 332 57 333 58 
<< m2 >>
rect 333 57 334 58 
<< m1 >>
rect 334 57 335 58 
<< m2 >>
rect 334 57 335 58 
<< m2 >>
rect 335 57 336 58 
<< m1 >>
rect 336 57 337 58 
<< m2 >>
rect 336 57 337 58 
<< m2c >>
rect 336 57 337 58 
<< m1 >>
rect 336 57 337 58 
<< m2 >>
rect 336 57 337 58 
<< m1 >>
rect 388 57 389 58 
<< m1 >>
rect 433 57 434 58 
<< m1 >>
rect 487 57 488 58 
<< m1 >>
rect 64 58 65 59 
<< m1 >>
rect 85 58 86 59 
<< m1 >>
rect 91 58 92 59 
<< m1 >>
rect 100 58 101 59 
<< m1 >>
rect 109 58 110 59 
<< m1 >>
rect 111 58 112 59 
<< m1 >>
rect 112 58 113 59 
<< m1 >>
rect 113 58 114 59 
<< m1 >>
rect 114 58 115 59 
<< m1 >>
rect 115 58 116 59 
<< m1 >>
rect 116 58 117 59 
<< m1 >>
rect 117 58 118 59 
<< m1 >>
rect 118 58 119 59 
<< m1 >>
rect 119 58 120 59 
<< m1 >>
rect 120 58 121 59 
<< m1 >>
rect 121 58 122 59 
<< m1 >>
rect 122 58 123 59 
<< m1 >>
rect 123 58 124 59 
<< m1 >>
rect 124 58 125 59 
<< m1 >>
rect 158 58 159 59 
<< m1 >>
rect 163 58 164 59 
<< m1 >>
rect 190 58 191 59 
<< m2 >>
rect 225 58 226 59 
<< m1 >>
rect 226 58 227 59 
<< m1 >>
rect 229 58 230 59 
<< m2 >>
rect 237 58 238 59 
<< m2 >>
rect 244 58 245 59 
<< m1 >>
rect 248 58 249 59 
<< m1 >>
rect 253 58 254 59 
<< m2 >>
rect 264 58 265 59 
<< m2 >>
rect 265 58 266 59 
<< m2 >>
rect 266 58 267 59 
<< m2 >>
rect 267 58 268 59 
<< m1 >>
rect 268 58 269 59 
<< m2 >>
rect 268 58 269 59 
<< m2 >>
rect 269 58 270 59 
<< m1 >>
rect 280 58 281 59 
<< m1 >>
rect 282 58 283 59 
<< m1 >>
rect 283 58 284 59 
<< m1 >>
rect 284 58 285 59 
<< m1 >>
rect 285 58 286 59 
<< m1 >>
rect 286 58 287 59 
<< m1 >>
rect 287 58 288 59 
<< m2 >>
rect 287 58 288 59 
<< m2c >>
rect 287 58 288 59 
<< m1 >>
rect 287 58 288 59 
<< m2 >>
rect 287 58 288 59 
<< m2 >>
rect 288 58 289 59 
<< m1 >>
rect 289 58 290 59 
<< m2 >>
rect 289 58 290 59 
<< m2 >>
rect 290 58 291 59 
<< m1 >>
rect 291 58 292 59 
<< m2 >>
rect 291 58 292 59 
<< m2c >>
rect 291 58 292 59 
<< m1 >>
rect 291 58 292 59 
<< m2 >>
rect 291 58 292 59 
<< m1 >>
rect 292 58 293 59 
<< m1 >>
rect 293 58 294 59 
<< m1 >>
rect 294 58 295 59 
<< m1 >>
rect 295 58 296 59 
<< m1 >>
rect 296 58 297 59 
<< m1 >>
rect 297 58 298 59 
<< m1 >>
rect 298 58 299 59 
<< m1 >>
rect 299 58 300 59 
<< m1 >>
rect 300 58 301 59 
<< m1 >>
rect 301 58 302 59 
<< m1 >>
rect 302 58 303 59 
<< m1 >>
rect 303 58 304 59 
<< m1 >>
rect 304 58 305 59 
<< m1 >>
rect 305 58 306 59 
<< m1 >>
rect 306 58 307 59 
<< m1 >>
rect 307 58 308 59 
<< m1 >>
rect 308 58 309 59 
<< m1 >>
rect 309 58 310 59 
<< m1 >>
rect 310 58 311 59 
<< m1 >>
rect 311 58 312 59 
<< m1 >>
rect 312 58 313 59 
<< m1 >>
rect 313 58 314 59 
<< m1 >>
rect 314 58 315 59 
<< m1 >>
rect 315 58 316 59 
<< m1 >>
rect 316 58 317 59 
<< m1 >>
rect 317 58 318 59 
<< m1 >>
rect 318 58 319 59 
<< m1 >>
rect 319 58 320 59 
<< m1 >>
rect 320 58 321 59 
<< m1 >>
rect 321 58 322 59 
<< m1 >>
rect 322 58 323 59 
<< m1 >>
rect 323 58 324 59 
<< m1 >>
rect 324 58 325 59 
<< m1 >>
rect 325 58 326 59 
<< m1 >>
rect 326 58 327 59 
<< m1 >>
rect 327 58 328 59 
<< m1 >>
rect 328 58 329 59 
<< m1 >>
rect 329 58 330 59 
<< m1 >>
rect 330 58 331 59 
<< m1 >>
rect 332 58 333 59 
<< m1 >>
rect 334 58 335 59 
<< m1 >>
rect 336 58 337 59 
<< m2 >>
rect 371 58 372 59 
<< m2 >>
rect 372 58 373 59 
<< m2 >>
rect 373 58 374 59 
<< m2 >>
rect 374 58 375 59 
<< m2 >>
rect 375 58 376 59 
<< m2 >>
rect 376 58 377 59 
<< m2 >>
rect 377 58 378 59 
<< m1 >>
rect 378 58 379 59 
<< m2 >>
rect 378 58 379 59 
<< m2c >>
rect 378 58 379 59 
<< m1 >>
rect 378 58 379 59 
<< m2 >>
rect 378 58 379 59 
<< m1 >>
rect 379 58 380 59 
<< m1 >>
rect 380 58 381 59 
<< m1 >>
rect 381 58 382 59 
<< m1 >>
rect 382 58 383 59 
<< m1 >>
rect 383 58 384 59 
<< m1 >>
rect 384 58 385 59 
<< m1 >>
rect 385 58 386 59 
<< m1 >>
rect 386 58 387 59 
<< m1 >>
rect 387 58 388 59 
<< m1 >>
rect 388 58 389 59 
<< m1 >>
rect 433 58 434 59 
<< m1 >>
rect 487 58 488 59 
<< m1 >>
rect 64 59 65 60 
<< m1 >>
rect 85 59 86 60 
<< m1 >>
rect 91 59 92 60 
<< m2 >>
rect 91 59 92 60 
<< m2c >>
rect 91 59 92 60 
<< m1 >>
rect 91 59 92 60 
<< m2 >>
rect 91 59 92 60 
<< m1 >>
rect 100 59 101 60 
<< m2 >>
rect 100 59 101 60 
<< m2c >>
rect 100 59 101 60 
<< m1 >>
rect 100 59 101 60 
<< m2 >>
rect 100 59 101 60 
<< m1 >>
rect 109 59 110 60 
<< m2 >>
rect 109 59 110 60 
<< m2c >>
rect 109 59 110 60 
<< m1 >>
rect 109 59 110 60 
<< m2 >>
rect 109 59 110 60 
<< m1 >>
rect 124 59 125 60 
<< m2 >>
rect 124 59 125 60 
<< m2c >>
rect 124 59 125 60 
<< m1 >>
rect 124 59 125 60 
<< m2 >>
rect 124 59 125 60 
<< m1 >>
rect 145 59 146 60 
<< m2 >>
rect 145 59 146 60 
<< m2c >>
rect 145 59 146 60 
<< m1 >>
rect 145 59 146 60 
<< m2 >>
rect 145 59 146 60 
<< m1 >>
rect 146 59 147 60 
<< m1 >>
rect 147 59 148 60 
<< m1 >>
rect 148 59 149 60 
<< m1 >>
rect 149 59 150 60 
<< m1 >>
rect 150 59 151 60 
<< m1 >>
rect 151 59 152 60 
<< m1 >>
rect 152 59 153 60 
<< m1 >>
rect 153 59 154 60 
<< m1 >>
rect 154 59 155 60 
<< m1 >>
rect 155 59 156 60 
<< m1 >>
rect 156 59 157 60 
<< m1 >>
rect 157 59 158 60 
<< m1 >>
rect 158 59 159 60 
<< m1 >>
rect 163 59 164 60 
<< m2 >>
rect 163 59 164 60 
<< m2c >>
rect 163 59 164 60 
<< m1 >>
rect 163 59 164 60 
<< m2 >>
rect 163 59 164 60 
<< m1 >>
rect 190 59 191 60 
<< m1 >>
rect 191 59 192 60 
<< m1 >>
rect 192 59 193 60 
<< m1 >>
rect 193 59 194 60 
<< m1 >>
rect 194 59 195 60 
<< m1 >>
rect 195 59 196 60 
<< m1 >>
rect 196 59 197 60 
<< m1 >>
rect 197 59 198 60 
<< m1 >>
rect 198 59 199 60 
<< m1 >>
rect 199 59 200 60 
<< m1 >>
rect 200 59 201 60 
<< m1 >>
rect 201 59 202 60 
<< m2 >>
rect 201 59 202 60 
<< m2c >>
rect 201 59 202 60 
<< m1 >>
rect 201 59 202 60 
<< m2 >>
rect 201 59 202 60 
<< m2 >>
rect 225 59 226 60 
<< m1 >>
rect 226 59 227 60 
<< m1 >>
rect 227 59 228 60 
<< m2 >>
rect 227 59 228 60 
<< m2c >>
rect 227 59 228 60 
<< m1 >>
rect 227 59 228 60 
<< m2 >>
rect 227 59 228 60 
<< m2 >>
rect 228 59 229 60 
<< m1 >>
rect 229 59 230 60 
<< m2 >>
rect 229 59 230 60 
<< m2 >>
rect 230 59 231 60 
<< m1 >>
rect 235 59 236 60 
<< m2 >>
rect 235 59 236 60 
<< m2c >>
rect 235 59 236 60 
<< m1 >>
rect 235 59 236 60 
<< m2 >>
rect 235 59 236 60 
<< m1 >>
rect 236 59 237 60 
<< m1 >>
rect 237 59 238 60 
<< m2 >>
rect 237 59 238 60 
<< m1 >>
rect 238 59 239 60 
<< m1 >>
rect 239 59 240 60 
<< m1 >>
rect 240 59 241 60 
<< m1 >>
rect 241 59 242 60 
<< m1 >>
rect 242 59 243 60 
<< m1 >>
rect 243 59 244 60 
<< m1 >>
rect 244 59 245 60 
<< m2 >>
rect 244 59 245 60 
<< m1 >>
rect 245 59 246 60 
<< m1 >>
rect 246 59 247 60 
<< m1 >>
rect 247 59 248 60 
<< m1 >>
rect 248 59 249 60 
<< m1 >>
rect 253 59 254 60 
<< m2 >>
rect 253 59 254 60 
<< m2c >>
rect 253 59 254 60 
<< m1 >>
rect 253 59 254 60 
<< m2 >>
rect 253 59 254 60 
<< m1 >>
rect 255 59 256 60 
<< m2 >>
rect 255 59 256 60 
<< m2c >>
rect 255 59 256 60 
<< m1 >>
rect 255 59 256 60 
<< m2 >>
rect 255 59 256 60 
<< m1 >>
rect 256 59 257 60 
<< m1 >>
rect 257 59 258 60 
<< m1 >>
rect 258 59 259 60 
<< m1 >>
rect 259 59 260 60 
<< m1 >>
rect 260 59 261 60 
<< m1 >>
rect 261 59 262 60 
<< m1 >>
rect 262 59 263 60 
<< m1 >>
rect 263 59 264 60 
<< m1 >>
rect 264 59 265 60 
<< m2 >>
rect 264 59 265 60 
<< m1 >>
rect 265 59 266 60 
<< m1 >>
rect 266 59 267 60 
<< m1 >>
rect 267 59 268 60 
<< m1 >>
rect 268 59 269 60 
<< m1 >>
rect 280 59 281 60 
<< m2 >>
rect 280 59 281 60 
<< m2c >>
rect 280 59 281 60 
<< m1 >>
rect 280 59 281 60 
<< m2 >>
rect 280 59 281 60 
<< m1 >>
rect 289 59 290 60 
<< m1 >>
rect 332 59 333 60 
<< m2 >>
rect 332 59 333 60 
<< m2c >>
rect 332 59 333 60 
<< m1 >>
rect 332 59 333 60 
<< m2 >>
rect 332 59 333 60 
<< m2 >>
rect 333 59 334 60 
<< m1 >>
rect 334 59 335 60 
<< m2 >>
rect 334 59 335 60 
<< m2 >>
rect 335 59 336 60 
<< m1 >>
rect 336 59 337 60 
<< m1 >>
rect 337 59 338 60 
<< m1 >>
rect 338 59 339 60 
<< m1 >>
rect 339 59 340 60 
<< m1 >>
rect 340 59 341 60 
<< m1 >>
rect 341 59 342 60 
<< m1 >>
rect 342 59 343 60 
<< m1 >>
rect 343 59 344 60 
<< m1 >>
rect 344 59 345 60 
<< m1 >>
rect 345 59 346 60 
<< m1 >>
rect 346 59 347 60 
<< m1 >>
rect 347 59 348 60 
<< m1 >>
rect 348 59 349 60 
<< m1 >>
rect 349 59 350 60 
<< m1 >>
rect 350 59 351 60 
<< m1 >>
rect 351 59 352 60 
<< m1 >>
rect 352 59 353 60 
<< m1 >>
rect 353 59 354 60 
<< m1 >>
rect 354 59 355 60 
<< m1 >>
rect 355 59 356 60 
<< m1 >>
rect 356 59 357 60 
<< m1 >>
rect 357 59 358 60 
<< m1 >>
rect 358 59 359 60 
<< m1 >>
rect 359 59 360 60 
<< m1 >>
rect 360 59 361 60 
<< m1 >>
rect 361 59 362 60 
<< m1 >>
rect 362 59 363 60 
<< m1 >>
rect 363 59 364 60 
<< m1 >>
rect 364 59 365 60 
<< m1 >>
rect 365 59 366 60 
<< m1 >>
rect 366 59 367 60 
<< m1 >>
rect 367 59 368 60 
<< m1 >>
rect 368 59 369 60 
<< m1 >>
rect 369 59 370 60 
<< m1 >>
rect 370 59 371 60 
<< m1 >>
rect 371 59 372 60 
<< m2 >>
rect 371 59 372 60 
<< m1 >>
rect 372 59 373 60 
<< m1 >>
rect 373 59 374 60 
<< m1 >>
rect 374 59 375 60 
<< m1 >>
rect 375 59 376 60 
<< m1 >>
rect 376 59 377 60 
<< m1 >>
rect 433 59 434 60 
<< m1 >>
rect 487 59 488 60 
<< m1 >>
rect 64 60 65 61 
<< m1 >>
rect 85 60 86 61 
<< m2 >>
rect 91 60 92 61 
<< m2 >>
rect 92 60 93 61 
<< m2 >>
rect 100 60 101 61 
<< m2 >>
rect 109 60 110 61 
<< m2 >>
rect 110 60 111 61 
<< m2 >>
rect 111 60 112 61 
<< m2 >>
rect 112 60 113 61 
<< m2 >>
rect 113 60 114 61 
<< m2 >>
rect 114 60 115 61 
<< m2 >>
rect 115 60 116 61 
<< m2 >>
rect 116 60 117 61 
<< m2 >>
rect 117 60 118 61 
<< m2 >>
rect 118 60 119 61 
<< m2 >>
rect 119 60 120 61 
<< m2 >>
rect 120 60 121 61 
<< m2 >>
rect 121 60 122 61 
<< m2 >>
rect 122 60 123 61 
<< m2 >>
rect 124 60 125 61 
<< m2 >>
rect 145 60 146 61 
<< m2 >>
rect 163 60 164 61 
<< m2 >>
rect 164 60 165 61 
<< m2 >>
rect 165 60 166 61 
<< m2 >>
rect 166 60 167 61 
<< m2 >>
rect 167 60 168 61 
<< m2 >>
rect 168 60 169 61 
<< m2 >>
rect 169 60 170 61 
<< m2 >>
rect 170 60 171 61 
<< m2 >>
rect 171 60 172 61 
<< m2 >>
rect 172 60 173 61 
<< m2 >>
rect 173 60 174 61 
<< m2 >>
rect 174 60 175 61 
<< m2 >>
rect 175 60 176 61 
<< m2 >>
rect 176 60 177 61 
<< m2 >>
rect 177 60 178 61 
<< m2 >>
rect 178 60 179 61 
<< m2 >>
rect 179 60 180 61 
<< m2 >>
rect 180 60 181 61 
<< m2 >>
rect 181 60 182 61 
<< m2 >>
rect 182 60 183 61 
<< m2 >>
rect 183 60 184 61 
<< m2 >>
rect 184 60 185 61 
<< m2 >>
rect 185 60 186 61 
<< m2 >>
rect 186 60 187 61 
<< m2 >>
rect 187 60 188 61 
<< m2 >>
rect 188 60 189 61 
<< m2 >>
rect 189 60 190 61 
<< m2 >>
rect 190 60 191 61 
<< m2 >>
rect 191 60 192 61 
<< m2 >>
rect 192 60 193 61 
<< m2 >>
rect 193 60 194 61 
<< m2 >>
rect 194 60 195 61 
<< m2 >>
rect 201 60 202 61 
<< m2 >>
rect 208 60 209 61 
<< m2 >>
rect 209 60 210 61 
<< m2 >>
rect 210 60 211 61 
<< m2 >>
rect 211 60 212 61 
<< m2 >>
rect 212 60 213 61 
<< m2 >>
rect 213 60 214 61 
<< m2 >>
rect 214 60 215 61 
<< m2 >>
rect 215 60 216 61 
<< m2 >>
rect 216 60 217 61 
<< m2 >>
rect 217 60 218 61 
<< m2 >>
rect 218 60 219 61 
<< m2 >>
rect 219 60 220 61 
<< m2 >>
rect 220 60 221 61 
<< m2 >>
rect 221 60 222 61 
<< m2 >>
rect 222 60 223 61 
<< m2 >>
rect 223 60 224 61 
<< m2 >>
rect 224 60 225 61 
<< m2 >>
rect 225 60 226 61 
<< m1 >>
rect 229 60 230 61 
<< m2 >>
rect 230 60 231 61 
<< m2 >>
rect 235 60 236 61 
<< m2 >>
rect 237 60 238 61 
<< m2 >>
rect 244 60 245 61 
<< m2 >>
rect 246 60 247 61 
<< m2 >>
rect 247 60 248 61 
<< m2 >>
rect 248 60 249 61 
<< m2 >>
rect 249 60 250 61 
<< m2 >>
rect 250 60 251 61 
<< m2 >>
rect 251 60 252 61 
<< m2 >>
rect 252 60 253 61 
<< m2 >>
rect 253 60 254 61 
<< m2 >>
rect 255 60 256 61 
<< m2 >>
rect 264 60 265 61 
<< m2 >>
rect 280 60 281 61 
<< m1 >>
rect 289 60 290 61 
<< m1 >>
rect 334 60 335 61 
<< m2 >>
rect 335 60 336 61 
<< m2 >>
rect 371 60 372 61 
<< m1 >>
rect 376 60 377 61 
<< m1 >>
rect 433 60 434 61 
<< m1 >>
rect 487 60 488 61 
<< m1 >>
rect 64 61 65 62 
<< m1 >>
rect 85 61 86 62 
<< m1 >>
rect 86 61 87 62 
<< m1 >>
rect 88 61 89 62 
<< m1 >>
rect 89 61 90 62 
<< m1 >>
rect 90 61 91 62 
<< m1 >>
rect 91 61 92 62 
<< m1 >>
rect 92 61 93 62 
<< m2 >>
rect 92 61 93 62 
<< m1 >>
rect 93 61 94 62 
<< m1 >>
rect 94 61 95 62 
<< m1 >>
rect 95 61 96 62 
<< m1 >>
rect 96 61 97 62 
<< m1 >>
rect 97 61 98 62 
<< m1 >>
rect 98 61 99 62 
<< m1 >>
rect 99 61 100 62 
<< m1 >>
rect 100 61 101 62 
<< m2 >>
rect 100 61 101 62 
<< m1 >>
rect 101 61 102 62 
<< m1 >>
rect 102 61 103 62 
<< m1 >>
rect 103 61 104 62 
<< m1 >>
rect 104 61 105 62 
<< m1 >>
rect 105 61 106 62 
<< m1 >>
rect 106 61 107 62 
<< m1 >>
rect 107 61 108 62 
<< m1 >>
rect 108 61 109 62 
<< m1 >>
rect 109 61 110 62 
<< m1 >>
rect 110 61 111 62 
<< m1 >>
rect 111 61 112 62 
<< m1 >>
rect 112 61 113 62 
<< m1 >>
rect 113 61 114 62 
<< m1 >>
rect 114 61 115 62 
<< m1 >>
rect 115 61 116 62 
<< m1 >>
rect 116 61 117 62 
<< m1 >>
rect 117 61 118 62 
<< m1 >>
rect 118 61 119 62 
<< m1 >>
rect 119 61 120 62 
<< m1 >>
rect 120 61 121 62 
<< m1 >>
rect 121 61 122 62 
<< m1 >>
rect 122 61 123 62 
<< m2 >>
rect 122 61 123 62 
<< m1 >>
rect 123 61 124 62 
<< m1 >>
rect 124 61 125 62 
<< m2 >>
rect 124 61 125 62 
<< m1 >>
rect 125 61 126 62 
<< m1 >>
rect 126 61 127 62 
<< m1 >>
rect 127 61 128 62 
<< m1 >>
rect 128 61 129 62 
<< m1 >>
rect 129 61 130 62 
<< m1 >>
rect 130 61 131 62 
<< m1 >>
rect 131 61 132 62 
<< m1 >>
rect 132 61 133 62 
<< m1 >>
rect 133 61 134 62 
<< m1 >>
rect 134 61 135 62 
<< m1 >>
rect 135 61 136 62 
<< m1 >>
rect 136 61 137 62 
<< m1 >>
rect 137 61 138 62 
<< m1 >>
rect 138 61 139 62 
<< m1 >>
rect 139 61 140 62 
<< m1 >>
rect 140 61 141 62 
<< m1 >>
rect 141 61 142 62 
<< m1 >>
rect 142 61 143 62 
<< m1 >>
rect 143 61 144 62 
<< m1 >>
rect 144 61 145 62 
<< m1 >>
rect 145 61 146 62 
<< m2 >>
rect 145 61 146 62 
<< m1 >>
rect 146 61 147 62 
<< m1 >>
rect 147 61 148 62 
<< m1 >>
rect 148 61 149 62 
<< m1 >>
rect 149 61 150 62 
<< m1 >>
rect 150 61 151 62 
<< m1 >>
rect 151 61 152 62 
<< m1 >>
rect 152 61 153 62 
<< m1 >>
rect 153 61 154 62 
<< m1 >>
rect 154 61 155 62 
<< m1 >>
rect 155 61 156 62 
<< m1 >>
rect 156 61 157 62 
<< m1 >>
rect 157 61 158 62 
<< m1 >>
rect 158 61 159 62 
<< m1 >>
rect 159 61 160 62 
<< m1 >>
rect 160 61 161 62 
<< m1 >>
rect 161 61 162 62 
<< m1 >>
rect 162 61 163 62 
<< m1 >>
rect 163 61 164 62 
<< m1 >>
rect 164 61 165 62 
<< m1 >>
rect 165 61 166 62 
<< m1 >>
rect 166 61 167 62 
<< m1 >>
rect 167 61 168 62 
<< m1 >>
rect 168 61 169 62 
<< m1 >>
rect 169 61 170 62 
<< m1 >>
rect 170 61 171 62 
<< m1 >>
rect 171 61 172 62 
<< m1 >>
rect 172 61 173 62 
<< m1 >>
rect 173 61 174 62 
<< m1 >>
rect 174 61 175 62 
<< m1 >>
rect 175 61 176 62 
<< m1 >>
rect 176 61 177 62 
<< m1 >>
rect 177 61 178 62 
<< m1 >>
rect 178 61 179 62 
<< m1 >>
rect 179 61 180 62 
<< m1 >>
rect 180 61 181 62 
<< m1 >>
rect 181 61 182 62 
<< m1 >>
rect 182 61 183 62 
<< m1 >>
rect 183 61 184 62 
<< m1 >>
rect 184 61 185 62 
<< m1 >>
rect 185 61 186 62 
<< m1 >>
rect 186 61 187 62 
<< m1 >>
rect 187 61 188 62 
<< m1 >>
rect 188 61 189 62 
<< m1 >>
rect 189 61 190 62 
<< m1 >>
rect 190 61 191 62 
<< m1 >>
rect 191 61 192 62 
<< m1 >>
rect 192 61 193 62 
<< m1 >>
rect 193 61 194 62 
<< m1 >>
rect 194 61 195 62 
<< m2 >>
rect 194 61 195 62 
<< m1 >>
rect 195 61 196 62 
<< m1 >>
rect 196 61 197 62 
<< m1 >>
rect 197 61 198 62 
<< m1 >>
rect 198 61 199 62 
<< m1 >>
rect 199 61 200 62 
<< m1 >>
rect 200 61 201 62 
<< m1 >>
rect 201 61 202 62 
<< m2 >>
rect 201 61 202 62 
<< m1 >>
rect 202 61 203 62 
<< m1 >>
rect 203 61 204 62 
<< m1 >>
rect 204 61 205 62 
<< m1 >>
rect 205 61 206 62 
<< m1 >>
rect 206 61 207 62 
<< m1 >>
rect 207 61 208 62 
<< m1 >>
rect 208 61 209 62 
<< m2 >>
rect 208 61 209 62 
<< m1 >>
rect 209 61 210 62 
<< m1 >>
rect 210 61 211 62 
<< m1 >>
rect 211 61 212 62 
<< m1 >>
rect 212 61 213 62 
<< m1 >>
rect 213 61 214 62 
<< m1 >>
rect 214 61 215 62 
<< m1 >>
rect 215 61 216 62 
<< m1 >>
rect 216 61 217 62 
<< m1 >>
rect 217 61 218 62 
<< m1 >>
rect 218 61 219 62 
<< m1 >>
rect 219 61 220 62 
<< m1 >>
rect 220 61 221 62 
<< m1 >>
rect 221 61 222 62 
<< m1 >>
rect 222 61 223 62 
<< m1 >>
rect 223 61 224 62 
<< m1 >>
rect 224 61 225 62 
<< m1 >>
rect 225 61 226 62 
<< m1 >>
rect 226 61 227 62 
<< m1 >>
rect 227 61 228 62 
<< m1 >>
rect 228 61 229 62 
<< m1 >>
rect 229 61 230 62 
<< m2 >>
rect 230 61 231 62 
<< m1 >>
rect 231 61 232 62 
<< m2 >>
rect 231 61 232 62 
<< m2c >>
rect 231 61 232 62 
<< m1 >>
rect 231 61 232 62 
<< m2 >>
rect 231 61 232 62 
<< m1 >>
rect 232 61 233 62 
<< m1 >>
rect 233 61 234 62 
<< m1 >>
rect 234 61 235 62 
<< m1 >>
rect 235 61 236 62 
<< m2 >>
rect 235 61 236 62 
<< m1 >>
rect 236 61 237 62 
<< m1 >>
rect 237 61 238 62 
<< m2 >>
rect 237 61 238 62 
<< m1 >>
rect 238 61 239 62 
<< m1 >>
rect 239 61 240 62 
<< m1 >>
rect 240 61 241 62 
<< m1 >>
rect 241 61 242 62 
<< m1 >>
rect 242 61 243 62 
<< m1 >>
rect 243 61 244 62 
<< m1 >>
rect 244 61 245 62 
<< m2 >>
rect 244 61 245 62 
<< m1 >>
rect 245 61 246 62 
<< m1 >>
rect 246 61 247 62 
<< m2 >>
rect 246 61 247 62 
<< m1 >>
rect 247 61 248 62 
<< m1 >>
rect 248 61 249 62 
<< m1 >>
rect 249 61 250 62 
<< m1 >>
rect 250 61 251 62 
<< m1 >>
rect 251 61 252 62 
<< m1 >>
rect 252 61 253 62 
<< m1 >>
rect 253 61 254 62 
<< m1 >>
rect 254 61 255 62 
<< m1 >>
rect 255 61 256 62 
<< m2 >>
rect 255 61 256 62 
<< m1 >>
rect 256 61 257 62 
<< m1 >>
rect 257 61 258 62 
<< m1 >>
rect 258 61 259 62 
<< m1 >>
rect 259 61 260 62 
<< m1 >>
rect 260 61 261 62 
<< m1 >>
rect 261 61 262 62 
<< m1 >>
rect 262 61 263 62 
<< m1 >>
rect 263 61 264 62 
<< m1 >>
rect 264 61 265 62 
<< m2 >>
rect 264 61 265 62 
<< m1 >>
rect 265 61 266 62 
<< m1 >>
rect 266 61 267 62 
<< m1 >>
rect 267 61 268 62 
<< m1 >>
rect 268 61 269 62 
<< m1 >>
rect 269 61 270 62 
<< m1 >>
rect 270 61 271 62 
<< m1 >>
rect 271 61 272 62 
<< m1 >>
rect 272 61 273 62 
<< m1 >>
rect 273 61 274 62 
<< m1 >>
rect 274 61 275 62 
<< m1 >>
rect 275 61 276 62 
<< m1 >>
rect 276 61 277 62 
<< m1 >>
rect 277 61 278 62 
<< m1 >>
rect 278 61 279 62 
<< m1 >>
rect 279 61 280 62 
<< m1 >>
rect 280 61 281 62 
<< m2 >>
rect 280 61 281 62 
<< m1 >>
rect 281 61 282 62 
<< m1 >>
rect 282 61 283 62 
<< m1 >>
rect 283 61 284 62 
<< m1 >>
rect 284 61 285 62 
<< m1 >>
rect 285 61 286 62 
<< m1 >>
rect 286 61 287 62 
<< m1 >>
rect 287 61 288 62 
<< m2 >>
rect 287 61 288 62 
<< m2c >>
rect 287 61 288 62 
<< m1 >>
rect 287 61 288 62 
<< m2 >>
rect 287 61 288 62 
<< m2 >>
rect 288 61 289 62 
<< m1 >>
rect 289 61 290 62 
<< m2 >>
rect 289 61 290 62 
<< m2 >>
rect 290 61 291 62 
<< m1 >>
rect 291 61 292 62 
<< m2 >>
rect 291 61 292 62 
<< m2c >>
rect 291 61 292 62 
<< m1 >>
rect 291 61 292 62 
<< m2 >>
rect 291 61 292 62 
<< m1 >>
rect 292 61 293 62 
<< m1 >>
rect 293 61 294 62 
<< m1 >>
rect 294 61 295 62 
<< m1 >>
rect 295 61 296 62 
<< m1 >>
rect 296 61 297 62 
<< m1 >>
rect 297 61 298 62 
<< m1 >>
rect 298 61 299 62 
<< m1 >>
rect 299 61 300 62 
<< m1 >>
rect 300 61 301 62 
<< m1 >>
rect 301 61 302 62 
<< m1 >>
rect 302 61 303 62 
<< m1 >>
rect 303 61 304 62 
<< m1 >>
rect 304 61 305 62 
<< m1 >>
rect 305 61 306 62 
<< m1 >>
rect 306 61 307 62 
<< m1 >>
rect 307 61 308 62 
<< m1 >>
rect 308 61 309 62 
<< m1 >>
rect 309 61 310 62 
<< m1 >>
rect 310 61 311 62 
<< m1 >>
rect 311 61 312 62 
<< m1 >>
rect 312 61 313 62 
<< m1 >>
rect 313 61 314 62 
<< m1 >>
rect 314 61 315 62 
<< m1 >>
rect 315 61 316 62 
<< m1 >>
rect 316 61 317 62 
<< m1 >>
rect 317 61 318 62 
<< m1 >>
rect 318 61 319 62 
<< m1 >>
rect 319 61 320 62 
<< m1 >>
rect 320 61 321 62 
<< m1 >>
rect 321 61 322 62 
<< m1 >>
rect 322 61 323 62 
<< m1 >>
rect 323 61 324 62 
<< m1 >>
rect 324 61 325 62 
<< m1 >>
rect 325 61 326 62 
<< m1 >>
rect 326 61 327 62 
<< m1 >>
rect 327 61 328 62 
<< m1 >>
rect 328 61 329 62 
<< m1 >>
rect 329 61 330 62 
<< m1 >>
rect 330 61 331 62 
<< m1 >>
rect 331 61 332 62 
<< m1 >>
rect 332 61 333 62 
<< m1 >>
rect 334 61 335 62 
<< m2 >>
rect 335 61 336 62 
<< m1 >>
rect 336 61 337 62 
<< m2 >>
rect 336 61 337 62 
<< m2c >>
rect 336 61 337 62 
<< m1 >>
rect 336 61 337 62 
<< m2 >>
rect 336 61 337 62 
<< m1 >>
rect 337 61 338 62 
<< m1 >>
rect 338 61 339 62 
<< m1 >>
rect 339 61 340 62 
<< m1 >>
rect 340 61 341 62 
<< m1 >>
rect 341 61 342 62 
<< m1 >>
rect 342 61 343 62 
<< m1 >>
rect 343 61 344 62 
<< m1 >>
rect 344 61 345 62 
<< m1 >>
rect 345 61 346 62 
<< m1 >>
rect 346 61 347 62 
<< m1 >>
rect 347 61 348 62 
<< m1 >>
rect 348 61 349 62 
<< m1 >>
rect 349 61 350 62 
<< m1 >>
rect 350 61 351 62 
<< m1 >>
rect 351 61 352 62 
<< m1 >>
rect 352 61 353 62 
<< m1 >>
rect 353 61 354 62 
<< m1 >>
rect 354 61 355 62 
<< m1 >>
rect 355 61 356 62 
<< m1 >>
rect 356 61 357 62 
<< m1 >>
rect 357 61 358 62 
<< m1 >>
rect 358 61 359 62 
<< m1 >>
rect 359 61 360 62 
<< m1 >>
rect 360 61 361 62 
<< m1 >>
rect 361 61 362 62 
<< m1 >>
rect 362 61 363 62 
<< m1 >>
rect 363 61 364 62 
<< m1 >>
rect 364 61 365 62 
<< m1 >>
rect 365 61 366 62 
<< m1 >>
rect 366 61 367 62 
<< m1 >>
rect 367 61 368 62 
<< m1 >>
rect 368 61 369 62 
<< m1 >>
rect 369 61 370 62 
<< m1 >>
rect 370 61 371 62 
<< m2 >>
rect 371 61 372 62 
<< m1 >>
rect 376 61 377 62 
<< m1 >>
rect 433 61 434 62 
<< m1 >>
rect 487 61 488 62 
<< m1 >>
rect 64 62 65 63 
<< m1 >>
rect 86 62 87 63 
<< m1 >>
rect 88 62 89 63 
<< m2 >>
rect 92 62 93 63 
<< m2 >>
rect 100 62 101 63 
<< m2 >>
rect 122 62 123 63 
<< m2 >>
rect 124 62 125 63 
<< m2 >>
rect 145 62 146 63 
<< m2 >>
rect 194 62 195 63 
<< m2 >>
rect 201 62 202 63 
<< m2 >>
rect 208 62 209 63 
<< m2 >>
rect 235 62 236 63 
<< m2 >>
rect 237 62 238 63 
<< m2 >>
rect 244 62 245 63 
<< m2 >>
rect 246 62 247 63 
<< m2 >>
rect 255 62 256 63 
<< m2 >>
rect 264 62 265 63 
<< m2 >>
rect 280 62 281 63 
<< m1 >>
rect 289 62 290 63 
<< m1 >>
rect 332 62 333 63 
<< m1 >>
rect 334 62 335 63 
<< m1 >>
rect 370 62 371 63 
<< m2 >>
rect 371 62 372 63 
<< m1 >>
rect 376 62 377 63 
<< m1 >>
rect 433 62 434 63 
<< m1 >>
rect 487 62 488 63 
<< m1 >>
rect 13 63 14 64 
<< m1 >>
rect 14 63 15 64 
<< m1 >>
rect 15 63 16 64 
<< m1 >>
rect 16 63 17 64 
<< m1 >>
rect 17 63 18 64 
<< m1 >>
rect 18 63 19 64 
<< m1 >>
rect 19 63 20 64 
<< m1 >>
rect 20 63 21 64 
<< m1 >>
rect 21 63 22 64 
<< m1 >>
rect 22 63 23 64 
<< m1 >>
rect 23 63 24 64 
<< m1 >>
rect 24 63 25 64 
<< m1 >>
rect 25 63 26 64 
<< m1 >>
rect 26 63 27 64 
<< m1 >>
rect 27 63 28 64 
<< m1 >>
rect 28 63 29 64 
<< m1 >>
rect 64 63 65 64 
<< m1 >>
rect 86 63 87 64 
<< m2 >>
rect 86 63 87 64 
<< m2c >>
rect 86 63 87 64 
<< m1 >>
rect 86 63 87 64 
<< m2 >>
rect 86 63 87 64 
<< m2 >>
rect 87 63 88 64 
<< m1 >>
rect 88 63 89 64 
<< m2 >>
rect 88 63 89 64 
<< m2 >>
rect 89 63 90 64 
<< m2 >>
rect 92 63 93 64 
<< m2 >>
rect 100 63 101 64 
<< m1 >>
rect 122 63 123 64 
<< m2 >>
rect 122 63 123 64 
<< m2c >>
rect 122 63 123 64 
<< m1 >>
rect 122 63 123 64 
<< m2 >>
rect 122 63 123 64 
<< m1 >>
rect 123 63 124 64 
<< m1 >>
rect 124 63 125 64 
<< m2 >>
rect 124 63 125 64 
<< m1 >>
rect 125 63 126 64 
<< m2 >>
rect 125 63 126 64 
<< m1 >>
rect 126 63 127 64 
<< m2 >>
rect 126 63 127 64 
<< m1 >>
rect 127 63 128 64 
<< m2 >>
rect 127 63 128 64 
<< m1 >>
rect 128 63 129 64 
<< m2 >>
rect 128 63 129 64 
<< m1 >>
rect 129 63 130 64 
<< m2 >>
rect 129 63 130 64 
<< m2 >>
rect 130 63 131 64 
<< m1 >>
rect 131 63 132 64 
<< m2 >>
rect 131 63 132 64 
<< m2c >>
rect 131 63 132 64 
<< m1 >>
rect 131 63 132 64 
<< m2 >>
rect 131 63 132 64 
<< m1 >>
rect 145 63 146 64 
<< m2 >>
rect 145 63 146 64 
<< m2c >>
rect 145 63 146 64 
<< m1 >>
rect 145 63 146 64 
<< m2 >>
rect 145 63 146 64 
<< m1 >>
rect 194 63 195 64 
<< m2 >>
rect 194 63 195 64 
<< m2c >>
rect 194 63 195 64 
<< m1 >>
rect 194 63 195 64 
<< m2 >>
rect 194 63 195 64 
<< m1 >>
rect 195 63 196 64 
<< m1 >>
rect 196 63 197 64 
<< m1 >>
rect 197 63 198 64 
<< m1 >>
rect 198 63 199 64 
<< m1 >>
rect 199 63 200 64 
<< m1 >>
rect 200 63 201 64 
<< m1 >>
rect 201 63 202 64 
<< m2 >>
rect 201 63 202 64 
<< m1 >>
rect 202 63 203 64 
<< m1 >>
rect 203 63 204 64 
<< m1 >>
rect 204 63 205 64 
<< m1 >>
rect 205 63 206 64 
<< m1 >>
rect 206 63 207 64 
<< m1 >>
rect 207 63 208 64 
<< m1 >>
rect 208 63 209 64 
<< m2 >>
rect 208 63 209 64 
<< m1 >>
rect 209 63 210 64 
<< m1 >>
rect 210 63 211 64 
<< m1 >>
rect 211 63 212 64 
<< m1 >>
rect 229 63 230 64 
<< m1 >>
rect 230 63 231 64 
<< m1 >>
rect 231 63 232 64 
<< m1 >>
rect 232 63 233 64 
<< m1 >>
rect 233 63 234 64 
<< m1 >>
rect 234 63 235 64 
<< m1 >>
rect 235 63 236 64 
<< m2 >>
rect 235 63 236 64 
<< m1 >>
rect 236 63 237 64 
<< m1 >>
rect 237 63 238 64 
<< m2 >>
rect 237 63 238 64 
<< m1 >>
rect 238 63 239 64 
<< m1 >>
rect 239 63 240 64 
<< m1 >>
rect 240 63 241 64 
<< m1 >>
rect 241 63 242 64 
<< m1 >>
rect 242 63 243 64 
<< m1 >>
rect 243 63 244 64 
<< m1 >>
rect 244 63 245 64 
<< m2 >>
rect 244 63 245 64 
<< m1 >>
rect 245 63 246 64 
<< m1 >>
rect 246 63 247 64 
<< m2 >>
rect 246 63 247 64 
<< m2c >>
rect 246 63 247 64 
<< m1 >>
rect 246 63 247 64 
<< m2 >>
rect 246 63 247 64 
<< m1 >>
rect 255 63 256 64 
<< m2 >>
rect 255 63 256 64 
<< m2c >>
rect 255 63 256 64 
<< m1 >>
rect 255 63 256 64 
<< m2 >>
rect 255 63 256 64 
<< m1 >>
rect 262 63 263 64 
<< m1 >>
rect 263 63 264 64 
<< m1 >>
rect 264 63 265 64 
<< m2 >>
rect 264 63 265 64 
<< m2c >>
rect 264 63 265 64 
<< m1 >>
rect 264 63 265 64 
<< m2 >>
rect 264 63 265 64 
<< m1 >>
rect 280 63 281 64 
<< m2 >>
rect 280 63 281 64 
<< m2c >>
rect 280 63 281 64 
<< m1 >>
rect 280 63 281 64 
<< m2 >>
rect 280 63 281 64 
<< m1 >>
rect 289 63 290 64 
<< m1 >>
rect 332 63 333 64 
<< m1 >>
rect 334 63 335 64 
<< m1 >>
rect 366 63 367 64 
<< m1 >>
rect 367 63 368 64 
<< m1 >>
rect 368 63 369 64 
<< m2 >>
rect 368 63 369 64 
<< m2c >>
rect 368 63 369 64 
<< m1 >>
rect 368 63 369 64 
<< m2 >>
rect 368 63 369 64 
<< m2 >>
rect 369 63 370 64 
<< m1 >>
rect 370 63 371 64 
<< m2 >>
rect 370 63 371 64 
<< m2 >>
rect 371 63 372 64 
<< m1 >>
rect 376 63 377 64 
<< m1 >>
rect 433 63 434 64 
<< m1 >>
rect 487 63 488 64 
<< m1 >>
rect 13 64 14 65 
<< m1 >>
rect 28 64 29 65 
<< m1 >>
rect 64 64 65 65 
<< m1 >>
rect 88 64 89 65 
<< m2 >>
rect 89 64 90 65 
<< m1 >>
rect 90 64 91 65 
<< m2 >>
rect 90 64 91 65 
<< m2c >>
rect 90 64 91 65 
<< m1 >>
rect 90 64 91 65 
<< m2 >>
rect 90 64 91 65 
<< m1 >>
rect 91 64 92 65 
<< m1 >>
rect 92 64 93 65 
<< m2 >>
rect 92 64 93 65 
<< m1 >>
rect 93 64 94 65 
<< m1 >>
rect 94 64 95 65 
<< m1 >>
rect 95 64 96 65 
<< m1 >>
rect 96 64 97 65 
<< m1 >>
rect 97 64 98 65 
<< m1 >>
rect 98 64 99 65 
<< m1 >>
rect 99 64 100 65 
<< m1 >>
rect 100 64 101 65 
<< m2 >>
rect 100 64 101 65 
<< m1 >>
rect 129 64 130 65 
<< m1 >>
rect 131 64 132 65 
<< m1 >>
rect 145 64 146 65 
<< m2 >>
rect 196 64 197 65 
<< m2 >>
rect 197 64 198 65 
<< m2 >>
rect 198 64 199 65 
<< m2 >>
rect 199 64 200 65 
<< m2 >>
rect 201 64 202 65 
<< m2 >>
rect 208 64 209 65 
<< m1 >>
rect 211 64 212 65 
<< m1 >>
rect 229 64 230 65 
<< m2 >>
rect 235 64 236 65 
<< m2 >>
rect 237 64 238 65 
<< m2 >>
rect 244 64 245 65 
<< m1 >>
rect 255 64 256 65 
<< m1 >>
rect 262 64 263 65 
<< m1 >>
rect 280 64 281 65 
<< m1 >>
rect 289 64 290 65 
<< m1 >>
rect 332 64 333 65 
<< m1 >>
rect 334 64 335 65 
<< m1 >>
rect 366 64 367 65 
<< m1 >>
rect 370 64 371 65 
<< m1 >>
rect 376 64 377 65 
<< m1 >>
rect 412 64 413 65 
<< m1 >>
rect 413 64 414 65 
<< m1 >>
rect 414 64 415 65 
<< m1 >>
rect 415 64 416 65 
<< m1 >>
rect 433 64 434 65 
<< m1 >>
rect 484 64 485 65 
<< m1 >>
rect 485 64 486 65 
<< m2 >>
rect 485 64 486 65 
<< m2c >>
rect 485 64 486 65 
<< m1 >>
rect 485 64 486 65 
<< m2 >>
rect 485 64 486 65 
<< m2 >>
rect 486 64 487 65 
<< m1 >>
rect 487 64 488 65 
<< m2 >>
rect 487 64 488 65 
<< m1 >>
rect 13 65 14 66 
<< m1 >>
rect 28 65 29 66 
<< m1 >>
rect 64 65 65 66 
<< m1 >>
rect 88 65 89 66 
<< m2 >>
rect 92 65 93 66 
<< m1 >>
rect 100 65 101 66 
<< m2 >>
rect 100 65 101 66 
<< m1 >>
rect 129 65 130 66 
<< m1 >>
rect 131 65 132 66 
<< m1 >>
rect 145 65 146 66 
<< m1 >>
rect 196 65 197 66 
<< m2 >>
rect 196 65 197 66 
<< m2c >>
rect 196 65 197 66 
<< m1 >>
rect 196 65 197 66 
<< m2 >>
rect 196 65 197 66 
<< m1 >>
rect 199 65 200 66 
<< m2 >>
rect 199 65 200 66 
<< m2c >>
rect 199 65 200 66 
<< m1 >>
rect 199 65 200 66 
<< m2 >>
rect 199 65 200 66 
<< m1 >>
rect 201 65 202 66 
<< m2 >>
rect 201 65 202 66 
<< m2c >>
rect 201 65 202 66 
<< m1 >>
rect 201 65 202 66 
<< m2 >>
rect 201 65 202 66 
<< m1 >>
rect 208 65 209 66 
<< m2 >>
rect 208 65 209 66 
<< m2c >>
rect 208 65 209 66 
<< m1 >>
rect 208 65 209 66 
<< m2 >>
rect 208 65 209 66 
<< m1 >>
rect 211 65 212 66 
<< m1 >>
rect 229 65 230 66 
<< m1 >>
rect 235 65 236 66 
<< m2 >>
rect 235 65 236 66 
<< m2c >>
rect 235 65 236 66 
<< m1 >>
rect 235 65 236 66 
<< m2 >>
rect 235 65 236 66 
<< m1 >>
rect 237 65 238 66 
<< m2 >>
rect 237 65 238 66 
<< m2c >>
rect 237 65 238 66 
<< m1 >>
rect 237 65 238 66 
<< m2 >>
rect 237 65 238 66 
<< m1 >>
rect 244 65 245 66 
<< m2 >>
rect 244 65 245 66 
<< m2c >>
rect 244 65 245 66 
<< m1 >>
rect 244 65 245 66 
<< m2 >>
rect 244 65 245 66 
<< m1 >>
rect 253 65 254 66 
<< m2 >>
rect 253 65 254 66 
<< m2c >>
rect 253 65 254 66 
<< m1 >>
rect 253 65 254 66 
<< m2 >>
rect 253 65 254 66 
<< m2 >>
rect 254 65 255 66 
<< m1 >>
rect 255 65 256 66 
<< m2 >>
rect 255 65 256 66 
<< m2 >>
rect 256 65 257 66 
<< m1 >>
rect 257 65 258 66 
<< m2 >>
rect 257 65 258 66 
<< m2c >>
rect 257 65 258 66 
<< m1 >>
rect 257 65 258 66 
<< m2 >>
rect 257 65 258 66 
<< m1 >>
rect 258 65 259 66 
<< m1 >>
rect 259 65 260 66 
<< m1 >>
rect 260 65 261 66 
<< m1 >>
rect 261 65 262 66 
<< m1 >>
rect 262 65 263 66 
<< m1 >>
rect 280 65 281 66 
<< m1 >>
rect 289 65 290 66 
<< m1 >>
rect 332 65 333 66 
<< m1 >>
rect 334 65 335 66 
<< m1 >>
rect 366 65 367 66 
<< m1 >>
rect 370 65 371 66 
<< m1 >>
rect 376 65 377 66 
<< m1 >>
rect 412 65 413 66 
<< m1 >>
rect 415 65 416 66 
<< m1 >>
rect 433 65 434 66 
<< m1 >>
rect 484 65 485 66 
<< m1 >>
rect 487 65 488 66 
<< m2 >>
rect 487 65 488 66 
<< pdiffusion >>
rect 12 66 13 67 
<< m1 >>
rect 13 66 14 67 
<< pdiffusion >>
rect 13 66 14 67 
<< pdiffusion >>
rect 14 66 15 67 
<< pdiffusion >>
rect 15 66 16 67 
<< pdiffusion >>
rect 16 66 17 67 
<< pdiffusion >>
rect 17 66 18 67 
<< m1 >>
rect 28 66 29 67 
<< pdiffusion >>
rect 30 66 31 67 
<< pdiffusion >>
rect 31 66 32 67 
<< pdiffusion >>
rect 32 66 33 67 
<< pdiffusion >>
rect 33 66 34 67 
<< pdiffusion >>
rect 34 66 35 67 
<< pdiffusion >>
rect 35 66 36 67 
<< pdiffusion >>
rect 48 66 49 67 
<< pdiffusion >>
rect 49 66 50 67 
<< pdiffusion >>
rect 50 66 51 67 
<< pdiffusion >>
rect 51 66 52 67 
<< pdiffusion >>
rect 52 66 53 67 
<< pdiffusion >>
rect 53 66 54 67 
<< m1 >>
rect 64 66 65 67 
<< pdiffusion >>
rect 66 66 67 67 
<< pdiffusion >>
rect 67 66 68 67 
<< pdiffusion >>
rect 68 66 69 67 
<< pdiffusion >>
rect 69 66 70 67 
<< pdiffusion >>
rect 70 66 71 67 
<< pdiffusion >>
rect 71 66 72 67 
<< pdiffusion >>
rect 84 66 85 67 
<< pdiffusion >>
rect 85 66 86 67 
<< pdiffusion >>
rect 86 66 87 67 
<< pdiffusion >>
rect 87 66 88 67 
<< m1 >>
rect 88 66 89 67 
<< pdiffusion >>
rect 88 66 89 67 
<< pdiffusion >>
rect 89 66 90 67 
<< m1 >>
rect 92 66 93 67 
<< m2 >>
rect 92 66 93 67 
<< m2c >>
rect 92 66 93 67 
<< m1 >>
rect 92 66 93 67 
<< m2 >>
rect 92 66 93 67 
<< m1 >>
rect 100 66 101 67 
<< m2 >>
rect 100 66 101 67 
<< pdiffusion >>
rect 102 66 103 67 
<< pdiffusion >>
rect 103 66 104 67 
<< pdiffusion >>
rect 104 66 105 67 
<< pdiffusion >>
rect 105 66 106 67 
<< pdiffusion >>
rect 106 66 107 67 
<< pdiffusion >>
rect 107 66 108 67 
<< pdiffusion >>
rect 120 66 121 67 
<< pdiffusion >>
rect 121 66 122 67 
<< pdiffusion >>
rect 122 66 123 67 
<< pdiffusion >>
rect 123 66 124 67 
<< pdiffusion >>
rect 124 66 125 67 
<< pdiffusion >>
rect 125 66 126 67 
<< m1 >>
rect 129 66 130 67 
<< m1 >>
rect 131 66 132 67 
<< pdiffusion >>
rect 138 66 139 67 
<< pdiffusion >>
rect 139 66 140 67 
<< pdiffusion >>
rect 140 66 141 67 
<< pdiffusion >>
rect 141 66 142 67 
<< pdiffusion >>
rect 142 66 143 67 
<< pdiffusion >>
rect 143 66 144 67 
<< m1 >>
rect 145 66 146 67 
<< pdiffusion >>
rect 156 66 157 67 
<< pdiffusion >>
rect 157 66 158 67 
<< pdiffusion >>
rect 158 66 159 67 
<< pdiffusion >>
rect 159 66 160 67 
<< pdiffusion >>
rect 160 66 161 67 
<< pdiffusion >>
rect 161 66 162 67 
<< pdiffusion >>
rect 174 66 175 67 
<< pdiffusion >>
rect 175 66 176 67 
<< pdiffusion >>
rect 176 66 177 67 
<< pdiffusion >>
rect 177 66 178 67 
<< pdiffusion >>
rect 178 66 179 67 
<< pdiffusion >>
rect 179 66 180 67 
<< pdiffusion >>
rect 192 66 193 67 
<< pdiffusion >>
rect 193 66 194 67 
<< pdiffusion >>
rect 194 66 195 67 
<< pdiffusion >>
rect 195 66 196 67 
<< m1 >>
rect 196 66 197 67 
<< pdiffusion >>
rect 196 66 197 67 
<< pdiffusion >>
rect 197 66 198 67 
<< m1 >>
rect 199 66 200 67 
<< m1 >>
rect 201 66 202 67 
<< m1 >>
rect 208 66 209 67 
<< pdiffusion >>
rect 210 66 211 67 
<< m1 >>
rect 211 66 212 67 
<< pdiffusion >>
rect 211 66 212 67 
<< pdiffusion >>
rect 212 66 213 67 
<< pdiffusion >>
rect 213 66 214 67 
<< pdiffusion >>
rect 214 66 215 67 
<< pdiffusion >>
rect 215 66 216 67 
<< pdiffusion >>
rect 228 66 229 67 
<< m1 >>
rect 229 66 230 67 
<< pdiffusion >>
rect 229 66 230 67 
<< pdiffusion >>
rect 230 66 231 67 
<< pdiffusion >>
rect 231 66 232 67 
<< pdiffusion >>
rect 232 66 233 67 
<< pdiffusion >>
rect 233 66 234 67 
<< m1 >>
rect 235 66 236 67 
<< m1 >>
rect 237 66 238 67 
<< m1 >>
rect 244 66 245 67 
<< pdiffusion >>
rect 246 66 247 67 
<< pdiffusion >>
rect 247 66 248 67 
<< pdiffusion >>
rect 248 66 249 67 
<< pdiffusion >>
rect 249 66 250 67 
<< pdiffusion >>
rect 250 66 251 67 
<< pdiffusion >>
rect 251 66 252 67 
<< m1 >>
rect 253 66 254 67 
<< m1 >>
rect 255 66 256 67 
<< pdiffusion >>
rect 264 66 265 67 
<< pdiffusion >>
rect 265 66 266 67 
<< pdiffusion >>
rect 266 66 267 67 
<< pdiffusion >>
rect 267 66 268 67 
<< pdiffusion >>
rect 268 66 269 67 
<< pdiffusion >>
rect 269 66 270 67 
<< m1 >>
rect 280 66 281 67 
<< pdiffusion >>
rect 282 66 283 67 
<< pdiffusion >>
rect 283 66 284 67 
<< pdiffusion >>
rect 284 66 285 67 
<< pdiffusion >>
rect 285 66 286 67 
<< pdiffusion >>
rect 286 66 287 67 
<< pdiffusion >>
rect 287 66 288 67 
<< m1 >>
rect 289 66 290 67 
<< pdiffusion >>
rect 300 66 301 67 
<< pdiffusion >>
rect 301 66 302 67 
<< pdiffusion >>
rect 302 66 303 67 
<< pdiffusion >>
rect 303 66 304 67 
<< pdiffusion >>
rect 304 66 305 67 
<< pdiffusion >>
rect 305 66 306 67 
<< pdiffusion >>
rect 318 66 319 67 
<< pdiffusion >>
rect 319 66 320 67 
<< pdiffusion >>
rect 320 66 321 67 
<< pdiffusion >>
rect 321 66 322 67 
<< pdiffusion >>
rect 322 66 323 67 
<< pdiffusion >>
rect 323 66 324 67 
<< m1 >>
rect 332 66 333 67 
<< m1 >>
rect 334 66 335 67 
<< pdiffusion >>
rect 336 66 337 67 
<< pdiffusion >>
rect 337 66 338 67 
<< pdiffusion >>
rect 338 66 339 67 
<< pdiffusion >>
rect 339 66 340 67 
<< pdiffusion >>
rect 340 66 341 67 
<< pdiffusion >>
rect 341 66 342 67 
<< pdiffusion >>
rect 354 66 355 67 
<< pdiffusion >>
rect 355 66 356 67 
<< pdiffusion >>
rect 356 66 357 67 
<< pdiffusion >>
rect 357 66 358 67 
<< pdiffusion >>
rect 358 66 359 67 
<< pdiffusion >>
rect 359 66 360 67 
<< m1 >>
rect 366 66 367 67 
<< m1 >>
rect 370 66 371 67 
<< pdiffusion >>
rect 372 66 373 67 
<< pdiffusion >>
rect 373 66 374 67 
<< pdiffusion >>
rect 374 66 375 67 
<< pdiffusion >>
rect 375 66 376 67 
<< m1 >>
rect 376 66 377 67 
<< pdiffusion >>
rect 376 66 377 67 
<< pdiffusion >>
rect 377 66 378 67 
<< pdiffusion >>
rect 390 66 391 67 
<< pdiffusion >>
rect 391 66 392 67 
<< pdiffusion >>
rect 392 66 393 67 
<< pdiffusion >>
rect 393 66 394 67 
<< pdiffusion >>
rect 394 66 395 67 
<< pdiffusion >>
rect 395 66 396 67 
<< pdiffusion >>
rect 408 66 409 67 
<< pdiffusion >>
rect 409 66 410 67 
<< pdiffusion >>
rect 410 66 411 67 
<< pdiffusion >>
rect 411 66 412 67 
<< m1 >>
rect 412 66 413 67 
<< pdiffusion >>
rect 412 66 413 67 
<< pdiffusion >>
rect 413 66 414 67 
<< m1 >>
rect 415 66 416 67 
<< pdiffusion >>
rect 426 66 427 67 
<< pdiffusion >>
rect 427 66 428 67 
<< pdiffusion >>
rect 428 66 429 67 
<< pdiffusion >>
rect 429 66 430 67 
<< pdiffusion >>
rect 430 66 431 67 
<< pdiffusion >>
rect 431 66 432 67 
<< m1 >>
rect 433 66 434 67 
<< pdiffusion >>
rect 462 66 463 67 
<< pdiffusion >>
rect 463 66 464 67 
<< pdiffusion >>
rect 464 66 465 67 
<< pdiffusion >>
rect 465 66 466 67 
<< pdiffusion >>
rect 466 66 467 67 
<< pdiffusion >>
rect 467 66 468 67 
<< pdiffusion >>
rect 480 66 481 67 
<< pdiffusion >>
rect 481 66 482 67 
<< pdiffusion >>
rect 482 66 483 67 
<< pdiffusion >>
rect 483 66 484 67 
<< m1 >>
rect 484 66 485 67 
<< pdiffusion >>
rect 484 66 485 67 
<< pdiffusion >>
rect 485 66 486 67 
<< m1 >>
rect 487 66 488 67 
<< m2 >>
rect 487 66 488 67 
<< pdiffusion >>
rect 498 66 499 67 
<< pdiffusion >>
rect 499 66 500 67 
<< pdiffusion >>
rect 500 66 501 67 
<< pdiffusion >>
rect 501 66 502 67 
<< pdiffusion >>
rect 502 66 503 67 
<< pdiffusion >>
rect 503 66 504 67 
<< pdiffusion >>
rect 516 66 517 67 
<< pdiffusion >>
rect 517 66 518 67 
<< pdiffusion >>
rect 518 66 519 67 
<< pdiffusion >>
rect 519 66 520 67 
<< pdiffusion >>
rect 520 66 521 67 
<< pdiffusion >>
rect 521 66 522 67 
<< pdiffusion >>
rect 12 67 13 68 
<< pdiffusion >>
rect 13 67 14 68 
<< pdiffusion >>
rect 14 67 15 68 
<< pdiffusion >>
rect 15 67 16 68 
<< pdiffusion >>
rect 16 67 17 68 
<< pdiffusion >>
rect 17 67 18 68 
<< m1 >>
rect 28 67 29 68 
<< pdiffusion >>
rect 30 67 31 68 
<< pdiffusion >>
rect 31 67 32 68 
<< pdiffusion >>
rect 32 67 33 68 
<< pdiffusion >>
rect 33 67 34 68 
<< pdiffusion >>
rect 34 67 35 68 
<< pdiffusion >>
rect 35 67 36 68 
<< pdiffusion >>
rect 48 67 49 68 
<< pdiffusion >>
rect 49 67 50 68 
<< pdiffusion >>
rect 50 67 51 68 
<< pdiffusion >>
rect 51 67 52 68 
<< pdiffusion >>
rect 52 67 53 68 
<< pdiffusion >>
rect 53 67 54 68 
<< m1 >>
rect 64 67 65 68 
<< pdiffusion >>
rect 66 67 67 68 
<< pdiffusion >>
rect 67 67 68 68 
<< pdiffusion >>
rect 68 67 69 68 
<< pdiffusion >>
rect 69 67 70 68 
<< pdiffusion >>
rect 70 67 71 68 
<< pdiffusion >>
rect 71 67 72 68 
<< pdiffusion >>
rect 84 67 85 68 
<< pdiffusion >>
rect 85 67 86 68 
<< pdiffusion >>
rect 86 67 87 68 
<< pdiffusion >>
rect 87 67 88 68 
<< pdiffusion >>
rect 88 67 89 68 
<< pdiffusion >>
rect 89 67 90 68 
<< m1 >>
rect 92 67 93 68 
<< m1 >>
rect 100 67 101 68 
<< m2 >>
rect 100 67 101 68 
<< pdiffusion >>
rect 102 67 103 68 
<< pdiffusion >>
rect 103 67 104 68 
<< pdiffusion >>
rect 104 67 105 68 
<< pdiffusion >>
rect 105 67 106 68 
<< pdiffusion >>
rect 106 67 107 68 
<< pdiffusion >>
rect 107 67 108 68 
<< pdiffusion >>
rect 120 67 121 68 
<< pdiffusion >>
rect 121 67 122 68 
<< pdiffusion >>
rect 122 67 123 68 
<< pdiffusion >>
rect 123 67 124 68 
<< pdiffusion >>
rect 124 67 125 68 
<< pdiffusion >>
rect 125 67 126 68 
<< m1 >>
rect 129 67 130 68 
<< m1 >>
rect 131 67 132 68 
<< pdiffusion >>
rect 138 67 139 68 
<< pdiffusion >>
rect 139 67 140 68 
<< pdiffusion >>
rect 140 67 141 68 
<< pdiffusion >>
rect 141 67 142 68 
<< pdiffusion >>
rect 142 67 143 68 
<< pdiffusion >>
rect 143 67 144 68 
<< m1 >>
rect 145 67 146 68 
<< pdiffusion >>
rect 156 67 157 68 
<< pdiffusion >>
rect 157 67 158 68 
<< pdiffusion >>
rect 158 67 159 68 
<< pdiffusion >>
rect 159 67 160 68 
<< pdiffusion >>
rect 160 67 161 68 
<< pdiffusion >>
rect 161 67 162 68 
<< pdiffusion >>
rect 174 67 175 68 
<< pdiffusion >>
rect 175 67 176 68 
<< pdiffusion >>
rect 176 67 177 68 
<< pdiffusion >>
rect 177 67 178 68 
<< pdiffusion >>
rect 178 67 179 68 
<< pdiffusion >>
rect 179 67 180 68 
<< pdiffusion >>
rect 192 67 193 68 
<< pdiffusion >>
rect 193 67 194 68 
<< pdiffusion >>
rect 194 67 195 68 
<< pdiffusion >>
rect 195 67 196 68 
<< pdiffusion >>
rect 196 67 197 68 
<< pdiffusion >>
rect 197 67 198 68 
<< m1 >>
rect 199 67 200 68 
<< m1 >>
rect 201 67 202 68 
<< m2 >>
rect 202 67 203 68 
<< m1 >>
rect 203 67 204 68 
<< m2 >>
rect 203 67 204 68 
<< m2c >>
rect 203 67 204 68 
<< m1 >>
rect 203 67 204 68 
<< m2 >>
rect 203 67 204 68 
<< m1 >>
rect 204 67 205 68 
<< m1 >>
rect 205 67 206 68 
<< m1 >>
rect 206 67 207 68 
<< m1 >>
rect 207 67 208 68 
<< m1 >>
rect 208 67 209 68 
<< pdiffusion >>
rect 210 67 211 68 
<< pdiffusion >>
rect 211 67 212 68 
<< pdiffusion >>
rect 212 67 213 68 
<< pdiffusion >>
rect 213 67 214 68 
<< pdiffusion >>
rect 214 67 215 68 
<< pdiffusion >>
rect 215 67 216 68 
<< pdiffusion >>
rect 228 67 229 68 
<< pdiffusion >>
rect 229 67 230 68 
<< pdiffusion >>
rect 230 67 231 68 
<< pdiffusion >>
rect 231 67 232 68 
<< pdiffusion >>
rect 232 67 233 68 
<< pdiffusion >>
rect 233 67 234 68 
<< m1 >>
rect 235 67 236 68 
<< m2 >>
rect 235 67 236 68 
<< m2 >>
rect 236 67 237 68 
<< m1 >>
rect 237 67 238 68 
<< m2 >>
rect 237 67 238 68 
<< m2 >>
rect 238 67 239 68 
<< m1 >>
rect 239 67 240 68 
<< m2 >>
rect 239 67 240 68 
<< m2c >>
rect 239 67 240 68 
<< m1 >>
rect 239 67 240 68 
<< m2 >>
rect 239 67 240 68 
<< m1 >>
rect 240 67 241 68 
<< m1 >>
rect 241 67 242 68 
<< m1 >>
rect 242 67 243 68 
<< m1 >>
rect 243 67 244 68 
<< m1 >>
rect 244 67 245 68 
<< pdiffusion >>
rect 246 67 247 68 
<< pdiffusion >>
rect 247 67 248 68 
<< pdiffusion >>
rect 248 67 249 68 
<< pdiffusion >>
rect 249 67 250 68 
<< pdiffusion >>
rect 250 67 251 68 
<< pdiffusion >>
rect 251 67 252 68 
<< m1 >>
rect 253 67 254 68 
<< m1 >>
rect 255 67 256 68 
<< pdiffusion >>
rect 264 67 265 68 
<< pdiffusion >>
rect 265 67 266 68 
<< pdiffusion >>
rect 266 67 267 68 
<< pdiffusion >>
rect 267 67 268 68 
<< pdiffusion >>
rect 268 67 269 68 
<< pdiffusion >>
rect 269 67 270 68 
<< m1 >>
rect 280 67 281 68 
<< pdiffusion >>
rect 282 67 283 68 
<< pdiffusion >>
rect 283 67 284 68 
<< pdiffusion >>
rect 284 67 285 68 
<< pdiffusion >>
rect 285 67 286 68 
<< pdiffusion >>
rect 286 67 287 68 
<< pdiffusion >>
rect 287 67 288 68 
<< m1 >>
rect 289 67 290 68 
<< pdiffusion >>
rect 300 67 301 68 
<< pdiffusion >>
rect 301 67 302 68 
<< pdiffusion >>
rect 302 67 303 68 
<< pdiffusion >>
rect 303 67 304 68 
<< pdiffusion >>
rect 304 67 305 68 
<< pdiffusion >>
rect 305 67 306 68 
<< pdiffusion >>
rect 318 67 319 68 
<< pdiffusion >>
rect 319 67 320 68 
<< pdiffusion >>
rect 320 67 321 68 
<< pdiffusion >>
rect 321 67 322 68 
<< pdiffusion >>
rect 322 67 323 68 
<< pdiffusion >>
rect 323 67 324 68 
<< m1 >>
rect 332 67 333 68 
<< m1 >>
rect 334 67 335 68 
<< pdiffusion >>
rect 336 67 337 68 
<< pdiffusion >>
rect 337 67 338 68 
<< pdiffusion >>
rect 338 67 339 68 
<< pdiffusion >>
rect 339 67 340 68 
<< pdiffusion >>
rect 340 67 341 68 
<< pdiffusion >>
rect 341 67 342 68 
<< pdiffusion >>
rect 354 67 355 68 
<< pdiffusion >>
rect 355 67 356 68 
<< pdiffusion >>
rect 356 67 357 68 
<< pdiffusion >>
rect 357 67 358 68 
<< pdiffusion >>
rect 358 67 359 68 
<< pdiffusion >>
rect 359 67 360 68 
<< m1 >>
rect 366 67 367 68 
<< m1 >>
rect 370 67 371 68 
<< pdiffusion >>
rect 372 67 373 68 
<< pdiffusion >>
rect 373 67 374 68 
<< pdiffusion >>
rect 374 67 375 68 
<< pdiffusion >>
rect 375 67 376 68 
<< pdiffusion >>
rect 376 67 377 68 
<< pdiffusion >>
rect 377 67 378 68 
<< pdiffusion >>
rect 390 67 391 68 
<< pdiffusion >>
rect 391 67 392 68 
<< pdiffusion >>
rect 392 67 393 68 
<< pdiffusion >>
rect 393 67 394 68 
<< pdiffusion >>
rect 394 67 395 68 
<< pdiffusion >>
rect 395 67 396 68 
<< pdiffusion >>
rect 408 67 409 68 
<< pdiffusion >>
rect 409 67 410 68 
<< pdiffusion >>
rect 410 67 411 68 
<< pdiffusion >>
rect 411 67 412 68 
<< pdiffusion >>
rect 412 67 413 68 
<< pdiffusion >>
rect 413 67 414 68 
<< m1 >>
rect 415 67 416 68 
<< pdiffusion >>
rect 426 67 427 68 
<< pdiffusion >>
rect 427 67 428 68 
<< pdiffusion >>
rect 428 67 429 68 
<< pdiffusion >>
rect 429 67 430 68 
<< pdiffusion >>
rect 430 67 431 68 
<< pdiffusion >>
rect 431 67 432 68 
<< m1 >>
rect 433 67 434 68 
<< pdiffusion >>
rect 462 67 463 68 
<< pdiffusion >>
rect 463 67 464 68 
<< pdiffusion >>
rect 464 67 465 68 
<< pdiffusion >>
rect 465 67 466 68 
<< pdiffusion >>
rect 466 67 467 68 
<< pdiffusion >>
rect 467 67 468 68 
<< pdiffusion >>
rect 480 67 481 68 
<< pdiffusion >>
rect 481 67 482 68 
<< pdiffusion >>
rect 482 67 483 68 
<< pdiffusion >>
rect 483 67 484 68 
<< pdiffusion >>
rect 484 67 485 68 
<< pdiffusion >>
rect 485 67 486 68 
<< m1 >>
rect 487 67 488 68 
<< m2 >>
rect 487 67 488 68 
<< pdiffusion >>
rect 498 67 499 68 
<< pdiffusion >>
rect 499 67 500 68 
<< pdiffusion >>
rect 500 67 501 68 
<< pdiffusion >>
rect 501 67 502 68 
<< pdiffusion >>
rect 502 67 503 68 
<< pdiffusion >>
rect 503 67 504 68 
<< pdiffusion >>
rect 516 67 517 68 
<< pdiffusion >>
rect 517 67 518 68 
<< pdiffusion >>
rect 518 67 519 68 
<< pdiffusion >>
rect 519 67 520 68 
<< pdiffusion >>
rect 520 67 521 68 
<< pdiffusion >>
rect 521 67 522 68 
<< pdiffusion >>
rect 12 68 13 69 
<< pdiffusion >>
rect 13 68 14 69 
<< pdiffusion >>
rect 14 68 15 69 
<< pdiffusion >>
rect 15 68 16 69 
<< pdiffusion >>
rect 16 68 17 69 
<< pdiffusion >>
rect 17 68 18 69 
<< m1 >>
rect 28 68 29 69 
<< pdiffusion >>
rect 30 68 31 69 
<< pdiffusion >>
rect 31 68 32 69 
<< pdiffusion >>
rect 32 68 33 69 
<< pdiffusion >>
rect 33 68 34 69 
<< pdiffusion >>
rect 34 68 35 69 
<< pdiffusion >>
rect 35 68 36 69 
<< pdiffusion >>
rect 48 68 49 69 
<< pdiffusion >>
rect 49 68 50 69 
<< pdiffusion >>
rect 50 68 51 69 
<< pdiffusion >>
rect 51 68 52 69 
<< pdiffusion >>
rect 52 68 53 69 
<< pdiffusion >>
rect 53 68 54 69 
<< m1 >>
rect 64 68 65 69 
<< pdiffusion >>
rect 66 68 67 69 
<< pdiffusion >>
rect 67 68 68 69 
<< pdiffusion >>
rect 68 68 69 69 
<< pdiffusion >>
rect 69 68 70 69 
<< pdiffusion >>
rect 70 68 71 69 
<< pdiffusion >>
rect 71 68 72 69 
<< pdiffusion >>
rect 84 68 85 69 
<< pdiffusion >>
rect 85 68 86 69 
<< pdiffusion >>
rect 86 68 87 69 
<< pdiffusion >>
rect 87 68 88 69 
<< pdiffusion >>
rect 88 68 89 69 
<< pdiffusion >>
rect 89 68 90 69 
<< m1 >>
rect 92 68 93 69 
<< m1 >>
rect 100 68 101 69 
<< m2 >>
rect 100 68 101 69 
<< pdiffusion >>
rect 102 68 103 69 
<< pdiffusion >>
rect 103 68 104 69 
<< pdiffusion >>
rect 104 68 105 69 
<< pdiffusion >>
rect 105 68 106 69 
<< pdiffusion >>
rect 106 68 107 69 
<< pdiffusion >>
rect 107 68 108 69 
<< pdiffusion >>
rect 120 68 121 69 
<< pdiffusion >>
rect 121 68 122 69 
<< pdiffusion >>
rect 122 68 123 69 
<< pdiffusion >>
rect 123 68 124 69 
<< pdiffusion >>
rect 124 68 125 69 
<< pdiffusion >>
rect 125 68 126 69 
<< m1 >>
rect 129 68 130 69 
<< m1 >>
rect 131 68 132 69 
<< pdiffusion >>
rect 138 68 139 69 
<< pdiffusion >>
rect 139 68 140 69 
<< pdiffusion >>
rect 140 68 141 69 
<< pdiffusion >>
rect 141 68 142 69 
<< pdiffusion >>
rect 142 68 143 69 
<< pdiffusion >>
rect 143 68 144 69 
<< m1 >>
rect 145 68 146 69 
<< pdiffusion >>
rect 156 68 157 69 
<< pdiffusion >>
rect 157 68 158 69 
<< pdiffusion >>
rect 158 68 159 69 
<< pdiffusion >>
rect 159 68 160 69 
<< pdiffusion >>
rect 160 68 161 69 
<< pdiffusion >>
rect 161 68 162 69 
<< pdiffusion >>
rect 174 68 175 69 
<< pdiffusion >>
rect 175 68 176 69 
<< pdiffusion >>
rect 176 68 177 69 
<< pdiffusion >>
rect 177 68 178 69 
<< pdiffusion >>
rect 178 68 179 69 
<< pdiffusion >>
rect 179 68 180 69 
<< pdiffusion >>
rect 192 68 193 69 
<< pdiffusion >>
rect 193 68 194 69 
<< pdiffusion >>
rect 194 68 195 69 
<< pdiffusion >>
rect 195 68 196 69 
<< pdiffusion >>
rect 196 68 197 69 
<< pdiffusion >>
rect 197 68 198 69 
<< m1 >>
rect 199 68 200 69 
<< m1 >>
rect 201 68 202 69 
<< m2 >>
rect 202 68 203 69 
<< pdiffusion >>
rect 210 68 211 69 
<< pdiffusion >>
rect 211 68 212 69 
<< pdiffusion >>
rect 212 68 213 69 
<< pdiffusion >>
rect 213 68 214 69 
<< pdiffusion >>
rect 214 68 215 69 
<< pdiffusion >>
rect 215 68 216 69 
<< pdiffusion >>
rect 228 68 229 69 
<< pdiffusion >>
rect 229 68 230 69 
<< pdiffusion >>
rect 230 68 231 69 
<< pdiffusion >>
rect 231 68 232 69 
<< pdiffusion >>
rect 232 68 233 69 
<< pdiffusion >>
rect 233 68 234 69 
<< m1 >>
rect 235 68 236 69 
<< m2 >>
rect 235 68 236 69 
<< m1 >>
rect 237 68 238 69 
<< pdiffusion >>
rect 246 68 247 69 
<< pdiffusion >>
rect 247 68 248 69 
<< pdiffusion >>
rect 248 68 249 69 
<< pdiffusion >>
rect 249 68 250 69 
<< pdiffusion >>
rect 250 68 251 69 
<< pdiffusion >>
rect 251 68 252 69 
<< m1 >>
rect 253 68 254 69 
<< m1 >>
rect 255 68 256 69 
<< pdiffusion >>
rect 264 68 265 69 
<< pdiffusion >>
rect 265 68 266 69 
<< pdiffusion >>
rect 266 68 267 69 
<< pdiffusion >>
rect 267 68 268 69 
<< pdiffusion >>
rect 268 68 269 69 
<< pdiffusion >>
rect 269 68 270 69 
<< m1 >>
rect 280 68 281 69 
<< pdiffusion >>
rect 282 68 283 69 
<< pdiffusion >>
rect 283 68 284 69 
<< pdiffusion >>
rect 284 68 285 69 
<< pdiffusion >>
rect 285 68 286 69 
<< pdiffusion >>
rect 286 68 287 69 
<< pdiffusion >>
rect 287 68 288 69 
<< m1 >>
rect 289 68 290 69 
<< pdiffusion >>
rect 300 68 301 69 
<< pdiffusion >>
rect 301 68 302 69 
<< pdiffusion >>
rect 302 68 303 69 
<< pdiffusion >>
rect 303 68 304 69 
<< pdiffusion >>
rect 304 68 305 69 
<< pdiffusion >>
rect 305 68 306 69 
<< pdiffusion >>
rect 318 68 319 69 
<< pdiffusion >>
rect 319 68 320 69 
<< pdiffusion >>
rect 320 68 321 69 
<< pdiffusion >>
rect 321 68 322 69 
<< pdiffusion >>
rect 322 68 323 69 
<< pdiffusion >>
rect 323 68 324 69 
<< m1 >>
rect 332 68 333 69 
<< m1 >>
rect 334 68 335 69 
<< pdiffusion >>
rect 336 68 337 69 
<< pdiffusion >>
rect 337 68 338 69 
<< pdiffusion >>
rect 338 68 339 69 
<< pdiffusion >>
rect 339 68 340 69 
<< pdiffusion >>
rect 340 68 341 69 
<< pdiffusion >>
rect 341 68 342 69 
<< pdiffusion >>
rect 354 68 355 69 
<< pdiffusion >>
rect 355 68 356 69 
<< pdiffusion >>
rect 356 68 357 69 
<< pdiffusion >>
rect 357 68 358 69 
<< pdiffusion >>
rect 358 68 359 69 
<< pdiffusion >>
rect 359 68 360 69 
<< m1 >>
rect 366 68 367 69 
<< m1 >>
rect 370 68 371 69 
<< pdiffusion >>
rect 372 68 373 69 
<< pdiffusion >>
rect 373 68 374 69 
<< pdiffusion >>
rect 374 68 375 69 
<< pdiffusion >>
rect 375 68 376 69 
<< pdiffusion >>
rect 376 68 377 69 
<< pdiffusion >>
rect 377 68 378 69 
<< pdiffusion >>
rect 390 68 391 69 
<< pdiffusion >>
rect 391 68 392 69 
<< pdiffusion >>
rect 392 68 393 69 
<< pdiffusion >>
rect 393 68 394 69 
<< pdiffusion >>
rect 394 68 395 69 
<< pdiffusion >>
rect 395 68 396 69 
<< pdiffusion >>
rect 408 68 409 69 
<< pdiffusion >>
rect 409 68 410 69 
<< pdiffusion >>
rect 410 68 411 69 
<< pdiffusion >>
rect 411 68 412 69 
<< pdiffusion >>
rect 412 68 413 69 
<< pdiffusion >>
rect 413 68 414 69 
<< m1 >>
rect 415 68 416 69 
<< pdiffusion >>
rect 426 68 427 69 
<< pdiffusion >>
rect 427 68 428 69 
<< pdiffusion >>
rect 428 68 429 69 
<< pdiffusion >>
rect 429 68 430 69 
<< pdiffusion >>
rect 430 68 431 69 
<< pdiffusion >>
rect 431 68 432 69 
<< m1 >>
rect 433 68 434 69 
<< pdiffusion >>
rect 462 68 463 69 
<< pdiffusion >>
rect 463 68 464 69 
<< pdiffusion >>
rect 464 68 465 69 
<< pdiffusion >>
rect 465 68 466 69 
<< pdiffusion >>
rect 466 68 467 69 
<< pdiffusion >>
rect 467 68 468 69 
<< pdiffusion >>
rect 480 68 481 69 
<< pdiffusion >>
rect 481 68 482 69 
<< pdiffusion >>
rect 482 68 483 69 
<< pdiffusion >>
rect 483 68 484 69 
<< pdiffusion >>
rect 484 68 485 69 
<< pdiffusion >>
rect 485 68 486 69 
<< m1 >>
rect 487 68 488 69 
<< m2 >>
rect 487 68 488 69 
<< pdiffusion >>
rect 498 68 499 69 
<< pdiffusion >>
rect 499 68 500 69 
<< pdiffusion >>
rect 500 68 501 69 
<< pdiffusion >>
rect 501 68 502 69 
<< pdiffusion >>
rect 502 68 503 69 
<< pdiffusion >>
rect 503 68 504 69 
<< pdiffusion >>
rect 516 68 517 69 
<< pdiffusion >>
rect 517 68 518 69 
<< pdiffusion >>
rect 518 68 519 69 
<< pdiffusion >>
rect 519 68 520 69 
<< pdiffusion >>
rect 520 68 521 69 
<< pdiffusion >>
rect 521 68 522 69 
<< pdiffusion >>
rect 12 69 13 70 
<< pdiffusion >>
rect 13 69 14 70 
<< pdiffusion >>
rect 14 69 15 70 
<< pdiffusion >>
rect 15 69 16 70 
<< pdiffusion >>
rect 16 69 17 70 
<< pdiffusion >>
rect 17 69 18 70 
<< m1 >>
rect 28 69 29 70 
<< pdiffusion >>
rect 30 69 31 70 
<< pdiffusion >>
rect 31 69 32 70 
<< pdiffusion >>
rect 32 69 33 70 
<< pdiffusion >>
rect 33 69 34 70 
<< pdiffusion >>
rect 34 69 35 70 
<< pdiffusion >>
rect 35 69 36 70 
<< pdiffusion >>
rect 48 69 49 70 
<< pdiffusion >>
rect 49 69 50 70 
<< pdiffusion >>
rect 50 69 51 70 
<< pdiffusion >>
rect 51 69 52 70 
<< pdiffusion >>
rect 52 69 53 70 
<< pdiffusion >>
rect 53 69 54 70 
<< m1 >>
rect 64 69 65 70 
<< pdiffusion >>
rect 66 69 67 70 
<< pdiffusion >>
rect 67 69 68 70 
<< pdiffusion >>
rect 68 69 69 70 
<< pdiffusion >>
rect 69 69 70 70 
<< pdiffusion >>
rect 70 69 71 70 
<< pdiffusion >>
rect 71 69 72 70 
<< pdiffusion >>
rect 84 69 85 70 
<< pdiffusion >>
rect 85 69 86 70 
<< pdiffusion >>
rect 86 69 87 70 
<< pdiffusion >>
rect 87 69 88 70 
<< pdiffusion >>
rect 88 69 89 70 
<< pdiffusion >>
rect 89 69 90 70 
<< m1 >>
rect 92 69 93 70 
<< m1 >>
rect 100 69 101 70 
<< m2 >>
rect 100 69 101 70 
<< pdiffusion >>
rect 102 69 103 70 
<< pdiffusion >>
rect 103 69 104 70 
<< pdiffusion >>
rect 104 69 105 70 
<< pdiffusion >>
rect 105 69 106 70 
<< pdiffusion >>
rect 106 69 107 70 
<< pdiffusion >>
rect 107 69 108 70 
<< pdiffusion >>
rect 120 69 121 70 
<< pdiffusion >>
rect 121 69 122 70 
<< pdiffusion >>
rect 122 69 123 70 
<< pdiffusion >>
rect 123 69 124 70 
<< pdiffusion >>
rect 124 69 125 70 
<< pdiffusion >>
rect 125 69 126 70 
<< m1 >>
rect 129 69 130 70 
<< m1 >>
rect 131 69 132 70 
<< pdiffusion >>
rect 138 69 139 70 
<< pdiffusion >>
rect 139 69 140 70 
<< pdiffusion >>
rect 140 69 141 70 
<< pdiffusion >>
rect 141 69 142 70 
<< pdiffusion >>
rect 142 69 143 70 
<< pdiffusion >>
rect 143 69 144 70 
<< m1 >>
rect 145 69 146 70 
<< pdiffusion >>
rect 156 69 157 70 
<< pdiffusion >>
rect 157 69 158 70 
<< pdiffusion >>
rect 158 69 159 70 
<< pdiffusion >>
rect 159 69 160 70 
<< pdiffusion >>
rect 160 69 161 70 
<< pdiffusion >>
rect 161 69 162 70 
<< pdiffusion >>
rect 174 69 175 70 
<< pdiffusion >>
rect 175 69 176 70 
<< pdiffusion >>
rect 176 69 177 70 
<< pdiffusion >>
rect 177 69 178 70 
<< pdiffusion >>
rect 178 69 179 70 
<< pdiffusion >>
rect 179 69 180 70 
<< pdiffusion >>
rect 192 69 193 70 
<< pdiffusion >>
rect 193 69 194 70 
<< pdiffusion >>
rect 194 69 195 70 
<< pdiffusion >>
rect 195 69 196 70 
<< pdiffusion >>
rect 196 69 197 70 
<< pdiffusion >>
rect 197 69 198 70 
<< m1 >>
rect 199 69 200 70 
<< m1 >>
rect 201 69 202 70 
<< m2 >>
rect 202 69 203 70 
<< pdiffusion >>
rect 210 69 211 70 
<< pdiffusion >>
rect 211 69 212 70 
<< pdiffusion >>
rect 212 69 213 70 
<< pdiffusion >>
rect 213 69 214 70 
<< pdiffusion >>
rect 214 69 215 70 
<< pdiffusion >>
rect 215 69 216 70 
<< pdiffusion >>
rect 228 69 229 70 
<< pdiffusion >>
rect 229 69 230 70 
<< pdiffusion >>
rect 230 69 231 70 
<< pdiffusion >>
rect 231 69 232 70 
<< pdiffusion >>
rect 232 69 233 70 
<< pdiffusion >>
rect 233 69 234 70 
<< m1 >>
rect 235 69 236 70 
<< m2 >>
rect 235 69 236 70 
<< m1 >>
rect 237 69 238 70 
<< pdiffusion >>
rect 246 69 247 70 
<< pdiffusion >>
rect 247 69 248 70 
<< pdiffusion >>
rect 248 69 249 70 
<< pdiffusion >>
rect 249 69 250 70 
<< pdiffusion >>
rect 250 69 251 70 
<< pdiffusion >>
rect 251 69 252 70 
<< m1 >>
rect 253 69 254 70 
<< m1 >>
rect 255 69 256 70 
<< pdiffusion >>
rect 264 69 265 70 
<< pdiffusion >>
rect 265 69 266 70 
<< pdiffusion >>
rect 266 69 267 70 
<< pdiffusion >>
rect 267 69 268 70 
<< pdiffusion >>
rect 268 69 269 70 
<< pdiffusion >>
rect 269 69 270 70 
<< m1 >>
rect 280 69 281 70 
<< pdiffusion >>
rect 282 69 283 70 
<< pdiffusion >>
rect 283 69 284 70 
<< pdiffusion >>
rect 284 69 285 70 
<< pdiffusion >>
rect 285 69 286 70 
<< pdiffusion >>
rect 286 69 287 70 
<< pdiffusion >>
rect 287 69 288 70 
<< m1 >>
rect 289 69 290 70 
<< pdiffusion >>
rect 300 69 301 70 
<< pdiffusion >>
rect 301 69 302 70 
<< pdiffusion >>
rect 302 69 303 70 
<< pdiffusion >>
rect 303 69 304 70 
<< pdiffusion >>
rect 304 69 305 70 
<< pdiffusion >>
rect 305 69 306 70 
<< pdiffusion >>
rect 318 69 319 70 
<< pdiffusion >>
rect 319 69 320 70 
<< pdiffusion >>
rect 320 69 321 70 
<< pdiffusion >>
rect 321 69 322 70 
<< pdiffusion >>
rect 322 69 323 70 
<< pdiffusion >>
rect 323 69 324 70 
<< m1 >>
rect 332 69 333 70 
<< m1 >>
rect 334 69 335 70 
<< pdiffusion >>
rect 336 69 337 70 
<< pdiffusion >>
rect 337 69 338 70 
<< pdiffusion >>
rect 338 69 339 70 
<< pdiffusion >>
rect 339 69 340 70 
<< pdiffusion >>
rect 340 69 341 70 
<< pdiffusion >>
rect 341 69 342 70 
<< pdiffusion >>
rect 354 69 355 70 
<< pdiffusion >>
rect 355 69 356 70 
<< pdiffusion >>
rect 356 69 357 70 
<< pdiffusion >>
rect 357 69 358 70 
<< pdiffusion >>
rect 358 69 359 70 
<< pdiffusion >>
rect 359 69 360 70 
<< m1 >>
rect 366 69 367 70 
<< m1 >>
rect 370 69 371 70 
<< pdiffusion >>
rect 372 69 373 70 
<< pdiffusion >>
rect 373 69 374 70 
<< pdiffusion >>
rect 374 69 375 70 
<< pdiffusion >>
rect 375 69 376 70 
<< pdiffusion >>
rect 376 69 377 70 
<< pdiffusion >>
rect 377 69 378 70 
<< pdiffusion >>
rect 390 69 391 70 
<< pdiffusion >>
rect 391 69 392 70 
<< pdiffusion >>
rect 392 69 393 70 
<< pdiffusion >>
rect 393 69 394 70 
<< pdiffusion >>
rect 394 69 395 70 
<< pdiffusion >>
rect 395 69 396 70 
<< pdiffusion >>
rect 408 69 409 70 
<< pdiffusion >>
rect 409 69 410 70 
<< pdiffusion >>
rect 410 69 411 70 
<< pdiffusion >>
rect 411 69 412 70 
<< pdiffusion >>
rect 412 69 413 70 
<< pdiffusion >>
rect 413 69 414 70 
<< m1 >>
rect 415 69 416 70 
<< pdiffusion >>
rect 426 69 427 70 
<< pdiffusion >>
rect 427 69 428 70 
<< pdiffusion >>
rect 428 69 429 70 
<< pdiffusion >>
rect 429 69 430 70 
<< pdiffusion >>
rect 430 69 431 70 
<< pdiffusion >>
rect 431 69 432 70 
<< m1 >>
rect 433 69 434 70 
<< pdiffusion >>
rect 462 69 463 70 
<< pdiffusion >>
rect 463 69 464 70 
<< pdiffusion >>
rect 464 69 465 70 
<< pdiffusion >>
rect 465 69 466 70 
<< pdiffusion >>
rect 466 69 467 70 
<< pdiffusion >>
rect 467 69 468 70 
<< pdiffusion >>
rect 480 69 481 70 
<< pdiffusion >>
rect 481 69 482 70 
<< pdiffusion >>
rect 482 69 483 70 
<< pdiffusion >>
rect 483 69 484 70 
<< pdiffusion >>
rect 484 69 485 70 
<< pdiffusion >>
rect 485 69 486 70 
<< m1 >>
rect 487 69 488 70 
<< m2 >>
rect 487 69 488 70 
<< pdiffusion >>
rect 498 69 499 70 
<< pdiffusion >>
rect 499 69 500 70 
<< pdiffusion >>
rect 500 69 501 70 
<< pdiffusion >>
rect 501 69 502 70 
<< pdiffusion >>
rect 502 69 503 70 
<< pdiffusion >>
rect 503 69 504 70 
<< pdiffusion >>
rect 516 69 517 70 
<< pdiffusion >>
rect 517 69 518 70 
<< pdiffusion >>
rect 518 69 519 70 
<< pdiffusion >>
rect 519 69 520 70 
<< pdiffusion >>
rect 520 69 521 70 
<< pdiffusion >>
rect 521 69 522 70 
<< pdiffusion >>
rect 12 70 13 71 
<< pdiffusion >>
rect 13 70 14 71 
<< pdiffusion >>
rect 14 70 15 71 
<< pdiffusion >>
rect 15 70 16 71 
<< pdiffusion >>
rect 16 70 17 71 
<< pdiffusion >>
rect 17 70 18 71 
<< m1 >>
rect 28 70 29 71 
<< pdiffusion >>
rect 30 70 31 71 
<< pdiffusion >>
rect 31 70 32 71 
<< pdiffusion >>
rect 32 70 33 71 
<< pdiffusion >>
rect 33 70 34 71 
<< pdiffusion >>
rect 34 70 35 71 
<< pdiffusion >>
rect 35 70 36 71 
<< pdiffusion >>
rect 48 70 49 71 
<< pdiffusion >>
rect 49 70 50 71 
<< pdiffusion >>
rect 50 70 51 71 
<< pdiffusion >>
rect 51 70 52 71 
<< pdiffusion >>
rect 52 70 53 71 
<< pdiffusion >>
rect 53 70 54 71 
<< m1 >>
rect 64 70 65 71 
<< pdiffusion >>
rect 66 70 67 71 
<< pdiffusion >>
rect 67 70 68 71 
<< pdiffusion >>
rect 68 70 69 71 
<< pdiffusion >>
rect 69 70 70 71 
<< pdiffusion >>
rect 70 70 71 71 
<< pdiffusion >>
rect 71 70 72 71 
<< pdiffusion >>
rect 84 70 85 71 
<< pdiffusion >>
rect 85 70 86 71 
<< pdiffusion >>
rect 86 70 87 71 
<< pdiffusion >>
rect 87 70 88 71 
<< pdiffusion >>
rect 88 70 89 71 
<< pdiffusion >>
rect 89 70 90 71 
<< m1 >>
rect 92 70 93 71 
<< m1 >>
rect 100 70 101 71 
<< m2 >>
rect 100 70 101 71 
<< pdiffusion >>
rect 102 70 103 71 
<< pdiffusion >>
rect 103 70 104 71 
<< pdiffusion >>
rect 104 70 105 71 
<< pdiffusion >>
rect 105 70 106 71 
<< pdiffusion >>
rect 106 70 107 71 
<< pdiffusion >>
rect 107 70 108 71 
<< pdiffusion >>
rect 120 70 121 71 
<< pdiffusion >>
rect 121 70 122 71 
<< pdiffusion >>
rect 122 70 123 71 
<< pdiffusion >>
rect 123 70 124 71 
<< pdiffusion >>
rect 124 70 125 71 
<< pdiffusion >>
rect 125 70 126 71 
<< m1 >>
rect 129 70 130 71 
<< m1 >>
rect 131 70 132 71 
<< pdiffusion >>
rect 138 70 139 71 
<< pdiffusion >>
rect 139 70 140 71 
<< pdiffusion >>
rect 140 70 141 71 
<< pdiffusion >>
rect 141 70 142 71 
<< pdiffusion >>
rect 142 70 143 71 
<< pdiffusion >>
rect 143 70 144 71 
<< m1 >>
rect 145 70 146 71 
<< pdiffusion >>
rect 156 70 157 71 
<< pdiffusion >>
rect 157 70 158 71 
<< pdiffusion >>
rect 158 70 159 71 
<< pdiffusion >>
rect 159 70 160 71 
<< pdiffusion >>
rect 160 70 161 71 
<< pdiffusion >>
rect 161 70 162 71 
<< pdiffusion >>
rect 174 70 175 71 
<< pdiffusion >>
rect 175 70 176 71 
<< pdiffusion >>
rect 176 70 177 71 
<< pdiffusion >>
rect 177 70 178 71 
<< pdiffusion >>
rect 178 70 179 71 
<< pdiffusion >>
rect 179 70 180 71 
<< pdiffusion >>
rect 192 70 193 71 
<< pdiffusion >>
rect 193 70 194 71 
<< pdiffusion >>
rect 194 70 195 71 
<< pdiffusion >>
rect 195 70 196 71 
<< pdiffusion >>
rect 196 70 197 71 
<< pdiffusion >>
rect 197 70 198 71 
<< m1 >>
rect 199 70 200 71 
<< m1 >>
rect 201 70 202 71 
<< m2 >>
rect 202 70 203 71 
<< pdiffusion >>
rect 210 70 211 71 
<< pdiffusion >>
rect 211 70 212 71 
<< pdiffusion >>
rect 212 70 213 71 
<< pdiffusion >>
rect 213 70 214 71 
<< pdiffusion >>
rect 214 70 215 71 
<< pdiffusion >>
rect 215 70 216 71 
<< pdiffusion >>
rect 228 70 229 71 
<< pdiffusion >>
rect 229 70 230 71 
<< pdiffusion >>
rect 230 70 231 71 
<< pdiffusion >>
rect 231 70 232 71 
<< pdiffusion >>
rect 232 70 233 71 
<< pdiffusion >>
rect 233 70 234 71 
<< m1 >>
rect 235 70 236 71 
<< m2 >>
rect 235 70 236 71 
<< m1 >>
rect 237 70 238 71 
<< pdiffusion >>
rect 246 70 247 71 
<< pdiffusion >>
rect 247 70 248 71 
<< pdiffusion >>
rect 248 70 249 71 
<< pdiffusion >>
rect 249 70 250 71 
<< pdiffusion >>
rect 250 70 251 71 
<< pdiffusion >>
rect 251 70 252 71 
<< m1 >>
rect 253 70 254 71 
<< m1 >>
rect 255 70 256 71 
<< pdiffusion >>
rect 264 70 265 71 
<< pdiffusion >>
rect 265 70 266 71 
<< pdiffusion >>
rect 266 70 267 71 
<< pdiffusion >>
rect 267 70 268 71 
<< pdiffusion >>
rect 268 70 269 71 
<< pdiffusion >>
rect 269 70 270 71 
<< m1 >>
rect 280 70 281 71 
<< pdiffusion >>
rect 282 70 283 71 
<< pdiffusion >>
rect 283 70 284 71 
<< pdiffusion >>
rect 284 70 285 71 
<< pdiffusion >>
rect 285 70 286 71 
<< pdiffusion >>
rect 286 70 287 71 
<< pdiffusion >>
rect 287 70 288 71 
<< m1 >>
rect 289 70 290 71 
<< pdiffusion >>
rect 300 70 301 71 
<< pdiffusion >>
rect 301 70 302 71 
<< pdiffusion >>
rect 302 70 303 71 
<< pdiffusion >>
rect 303 70 304 71 
<< pdiffusion >>
rect 304 70 305 71 
<< pdiffusion >>
rect 305 70 306 71 
<< pdiffusion >>
rect 318 70 319 71 
<< pdiffusion >>
rect 319 70 320 71 
<< pdiffusion >>
rect 320 70 321 71 
<< pdiffusion >>
rect 321 70 322 71 
<< pdiffusion >>
rect 322 70 323 71 
<< pdiffusion >>
rect 323 70 324 71 
<< m1 >>
rect 332 70 333 71 
<< m1 >>
rect 334 70 335 71 
<< pdiffusion >>
rect 336 70 337 71 
<< pdiffusion >>
rect 337 70 338 71 
<< pdiffusion >>
rect 338 70 339 71 
<< pdiffusion >>
rect 339 70 340 71 
<< pdiffusion >>
rect 340 70 341 71 
<< pdiffusion >>
rect 341 70 342 71 
<< pdiffusion >>
rect 354 70 355 71 
<< pdiffusion >>
rect 355 70 356 71 
<< pdiffusion >>
rect 356 70 357 71 
<< pdiffusion >>
rect 357 70 358 71 
<< pdiffusion >>
rect 358 70 359 71 
<< pdiffusion >>
rect 359 70 360 71 
<< m1 >>
rect 366 70 367 71 
<< m1 >>
rect 370 70 371 71 
<< pdiffusion >>
rect 372 70 373 71 
<< pdiffusion >>
rect 373 70 374 71 
<< pdiffusion >>
rect 374 70 375 71 
<< pdiffusion >>
rect 375 70 376 71 
<< pdiffusion >>
rect 376 70 377 71 
<< pdiffusion >>
rect 377 70 378 71 
<< pdiffusion >>
rect 390 70 391 71 
<< pdiffusion >>
rect 391 70 392 71 
<< pdiffusion >>
rect 392 70 393 71 
<< pdiffusion >>
rect 393 70 394 71 
<< pdiffusion >>
rect 394 70 395 71 
<< pdiffusion >>
rect 395 70 396 71 
<< pdiffusion >>
rect 408 70 409 71 
<< pdiffusion >>
rect 409 70 410 71 
<< pdiffusion >>
rect 410 70 411 71 
<< pdiffusion >>
rect 411 70 412 71 
<< pdiffusion >>
rect 412 70 413 71 
<< pdiffusion >>
rect 413 70 414 71 
<< m1 >>
rect 415 70 416 71 
<< pdiffusion >>
rect 426 70 427 71 
<< pdiffusion >>
rect 427 70 428 71 
<< pdiffusion >>
rect 428 70 429 71 
<< pdiffusion >>
rect 429 70 430 71 
<< pdiffusion >>
rect 430 70 431 71 
<< pdiffusion >>
rect 431 70 432 71 
<< m1 >>
rect 433 70 434 71 
<< pdiffusion >>
rect 462 70 463 71 
<< pdiffusion >>
rect 463 70 464 71 
<< pdiffusion >>
rect 464 70 465 71 
<< pdiffusion >>
rect 465 70 466 71 
<< pdiffusion >>
rect 466 70 467 71 
<< pdiffusion >>
rect 467 70 468 71 
<< pdiffusion >>
rect 480 70 481 71 
<< pdiffusion >>
rect 481 70 482 71 
<< pdiffusion >>
rect 482 70 483 71 
<< pdiffusion >>
rect 483 70 484 71 
<< pdiffusion >>
rect 484 70 485 71 
<< pdiffusion >>
rect 485 70 486 71 
<< m1 >>
rect 487 70 488 71 
<< m2 >>
rect 487 70 488 71 
<< pdiffusion >>
rect 498 70 499 71 
<< pdiffusion >>
rect 499 70 500 71 
<< pdiffusion >>
rect 500 70 501 71 
<< pdiffusion >>
rect 501 70 502 71 
<< pdiffusion >>
rect 502 70 503 71 
<< pdiffusion >>
rect 503 70 504 71 
<< pdiffusion >>
rect 516 70 517 71 
<< pdiffusion >>
rect 517 70 518 71 
<< pdiffusion >>
rect 518 70 519 71 
<< pdiffusion >>
rect 519 70 520 71 
<< pdiffusion >>
rect 520 70 521 71 
<< pdiffusion >>
rect 521 70 522 71 
<< pdiffusion >>
rect 12 71 13 72 
<< pdiffusion >>
rect 13 71 14 72 
<< pdiffusion >>
rect 14 71 15 72 
<< pdiffusion >>
rect 15 71 16 72 
<< pdiffusion >>
rect 16 71 17 72 
<< pdiffusion >>
rect 17 71 18 72 
<< m1 >>
rect 28 71 29 72 
<< pdiffusion >>
rect 30 71 31 72 
<< pdiffusion >>
rect 31 71 32 72 
<< pdiffusion >>
rect 32 71 33 72 
<< pdiffusion >>
rect 33 71 34 72 
<< pdiffusion >>
rect 34 71 35 72 
<< pdiffusion >>
rect 35 71 36 72 
<< pdiffusion >>
rect 48 71 49 72 
<< pdiffusion >>
rect 49 71 50 72 
<< pdiffusion >>
rect 50 71 51 72 
<< pdiffusion >>
rect 51 71 52 72 
<< pdiffusion >>
rect 52 71 53 72 
<< pdiffusion >>
rect 53 71 54 72 
<< m1 >>
rect 64 71 65 72 
<< pdiffusion >>
rect 66 71 67 72 
<< pdiffusion >>
rect 67 71 68 72 
<< pdiffusion >>
rect 68 71 69 72 
<< pdiffusion >>
rect 69 71 70 72 
<< pdiffusion >>
rect 70 71 71 72 
<< pdiffusion >>
rect 71 71 72 72 
<< pdiffusion >>
rect 84 71 85 72 
<< pdiffusion >>
rect 85 71 86 72 
<< pdiffusion >>
rect 86 71 87 72 
<< pdiffusion >>
rect 87 71 88 72 
<< pdiffusion >>
rect 88 71 89 72 
<< pdiffusion >>
rect 89 71 90 72 
<< m1 >>
rect 92 71 93 72 
<< m1 >>
rect 100 71 101 72 
<< m2 >>
rect 100 71 101 72 
<< pdiffusion >>
rect 102 71 103 72 
<< pdiffusion >>
rect 103 71 104 72 
<< pdiffusion >>
rect 104 71 105 72 
<< pdiffusion >>
rect 105 71 106 72 
<< pdiffusion >>
rect 106 71 107 72 
<< pdiffusion >>
rect 107 71 108 72 
<< pdiffusion >>
rect 120 71 121 72 
<< pdiffusion >>
rect 121 71 122 72 
<< pdiffusion >>
rect 122 71 123 72 
<< pdiffusion >>
rect 123 71 124 72 
<< m1 >>
rect 124 71 125 72 
<< pdiffusion >>
rect 124 71 125 72 
<< pdiffusion >>
rect 125 71 126 72 
<< m1 >>
rect 129 71 130 72 
<< m1 >>
rect 131 71 132 72 
<< pdiffusion >>
rect 138 71 139 72 
<< pdiffusion >>
rect 139 71 140 72 
<< pdiffusion >>
rect 140 71 141 72 
<< pdiffusion >>
rect 141 71 142 72 
<< m1 >>
rect 142 71 143 72 
<< pdiffusion >>
rect 142 71 143 72 
<< pdiffusion >>
rect 143 71 144 72 
<< m1 >>
rect 145 71 146 72 
<< m2 >>
rect 145 71 146 72 
<< m2c >>
rect 145 71 146 72 
<< m1 >>
rect 145 71 146 72 
<< m2 >>
rect 145 71 146 72 
<< pdiffusion >>
rect 156 71 157 72 
<< pdiffusion >>
rect 157 71 158 72 
<< pdiffusion >>
rect 158 71 159 72 
<< pdiffusion >>
rect 159 71 160 72 
<< m1 >>
rect 160 71 161 72 
<< pdiffusion >>
rect 160 71 161 72 
<< pdiffusion >>
rect 161 71 162 72 
<< pdiffusion >>
rect 174 71 175 72 
<< pdiffusion >>
rect 175 71 176 72 
<< pdiffusion >>
rect 176 71 177 72 
<< pdiffusion >>
rect 177 71 178 72 
<< pdiffusion >>
rect 178 71 179 72 
<< pdiffusion >>
rect 179 71 180 72 
<< pdiffusion >>
rect 192 71 193 72 
<< pdiffusion >>
rect 193 71 194 72 
<< pdiffusion >>
rect 194 71 195 72 
<< pdiffusion >>
rect 195 71 196 72 
<< pdiffusion >>
rect 196 71 197 72 
<< pdiffusion >>
rect 197 71 198 72 
<< m1 >>
rect 199 71 200 72 
<< m1 >>
rect 201 71 202 72 
<< m2 >>
rect 202 71 203 72 
<< pdiffusion >>
rect 210 71 211 72 
<< pdiffusion >>
rect 211 71 212 72 
<< pdiffusion >>
rect 212 71 213 72 
<< pdiffusion >>
rect 213 71 214 72 
<< m1 >>
rect 214 71 215 72 
<< pdiffusion >>
rect 214 71 215 72 
<< pdiffusion >>
rect 215 71 216 72 
<< pdiffusion >>
rect 228 71 229 72 
<< pdiffusion >>
rect 229 71 230 72 
<< pdiffusion >>
rect 230 71 231 72 
<< pdiffusion >>
rect 231 71 232 72 
<< pdiffusion >>
rect 232 71 233 72 
<< pdiffusion >>
rect 233 71 234 72 
<< m1 >>
rect 235 71 236 72 
<< m2 >>
rect 235 71 236 72 
<< m1 >>
rect 237 71 238 72 
<< pdiffusion >>
rect 246 71 247 72 
<< m1 >>
rect 247 71 248 72 
<< pdiffusion >>
rect 247 71 248 72 
<< pdiffusion >>
rect 248 71 249 72 
<< pdiffusion >>
rect 249 71 250 72 
<< pdiffusion >>
rect 250 71 251 72 
<< pdiffusion >>
rect 251 71 252 72 
<< m1 >>
rect 253 71 254 72 
<< m1 >>
rect 255 71 256 72 
<< pdiffusion >>
rect 264 71 265 72 
<< pdiffusion >>
rect 265 71 266 72 
<< pdiffusion >>
rect 266 71 267 72 
<< pdiffusion >>
rect 267 71 268 72 
<< pdiffusion >>
rect 268 71 269 72 
<< pdiffusion >>
rect 269 71 270 72 
<< m1 >>
rect 280 71 281 72 
<< pdiffusion >>
rect 282 71 283 72 
<< pdiffusion >>
rect 283 71 284 72 
<< pdiffusion >>
rect 284 71 285 72 
<< pdiffusion >>
rect 285 71 286 72 
<< pdiffusion >>
rect 286 71 287 72 
<< pdiffusion >>
rect 287 71 288 72 
<< m1 >>
rect 289 71 290 72 
<< pdiffusion >>
rect 300 71 301 72 
<< pdiffusion >>
rect 301 71 302 72 
<< pdiffusion >>
rect 302 71 303 72 
<< pdiffusion >>
rect 303 71 304 72 
<< pdiffusion >>
rect 304 71 305 72 
<< pdiffusion >>
rect 305 71 306 72 
<< pdiffusion >>
rect 318 71 319 72 
<< pdiffusion >>
rect 319 71 320 72 
<< pdiffusion >>
rect 320 71 321 72 
<< pdiffusion >>
rect 321 71 322 72 
<< pdiffusion >>
rect 322 71 323 72 
<< pdiffusion >>
rect 323 71 324 72 
<< m1 >>
rect 332 71 333 72 
<< m1 >>
rect 334 71 335 72 
<< pdiffusion >>
rect 336 71 337 72 
<< pdiffusion >>
rect 337 71 338 72 
<< pdiffusion >>
rect 338 71 339 72 
<< pdiffusion >>
rect 339 71 340 72 
<< m1 >>
rect 340 71 341 72 
<< pdiffusion >>
rect 340 71 341 72 
<< pdiffusion >>
rect 341 71 342 72 
<< pdiffusion >>
rect 354 71 355 72 
<< pdiffusion >>
rect 355 71 356 72 
<< pdiffusion >>
rect 356 71 357 72 
<< pdiffusion >>
rect 357 71 358 72 
<< m1 >>
rect 358 71 359 72 
<< pdiffusion >>
rect 358 71 359 72 
<< pdiffusion >>
rect 359 71 360 72 
<< m1 >>
rect 366 71 367 72 
<< m1 >>
rect 370 71 371 72 
<< pdiffusion >>
rect 372 71 373 72 
<< pdiffusion >>
rect 373 71 374 72 
<< pdiffusion >>
rect 374 71 375 72 
<< pdiffusion >>
rect 375 71 376 72 
<< pdiffusion >>
rect 376 71 377 72 
<< pdiffusion >>
rect 377 71 378 72 
<< pdiffusion >>
rect 390 71 391 72 
<< pdiffusion >>
rect 391 71 392 72 
<< pdiffusion >>
rect 392 71 393 72 
<< pdiffusion >>
rect 393 71 394 72 
<< pdiffusion >>
rect 394 71 395 72 
<< pdiffusion >>
rect 395 71 396 72 
<< pdiffusion >>
rect 408 71 409 72 
<< pdiffusion >>
rect 409 71 410 72 
<< pdiffusion >>
rect 410 71 411 72 
<< pdiffusion >>
rect 411 71 412 72 
<< pdiffusion >>
rect 412 71 413 72 
<< pdiffusion >>
rect 413 71 414 72 
<< m1 >>
rect 415 71 416 72 
<< pdiffusion >>
rect 426 71 427 72 
<< pdiffusion >>
rect 427 71 428 72 
<< pdiffusion >>
rect 428 71 429 72 
<< pdiffusion >>
rect 429 71 430 72 
<< pdiffusion >>
rect 430 71 431 72 
<< pdiffusion >>
rect 431 71 432 72 
<< m1 >>
rect 433 71 434 72 
<< pdiffusion >>
rect 462 71 463 72 
<< pdiffusion >>
rect 463 71 464 72 
<< pdiffusion >>
rect 464 71 465 72 
<< pdiffusion >>
rect 465 71 466 72 
<< pdiffusion >>
rect 466 71 467 72 
<< pdiffusion >>
rect 467 71 468 72 
<< pdiffusion >>
rect 480 71 481 72 
<< pdiffusion >>
rect 481 71 482 72 
<< pdiffusion >>
rect 482 71 483 72 
<< pdiffusion >>
rect 483 71 484 72 
<< pdiffusion >>
rect 484 71 485 72 
<< pdiffusion >>
rect 485 71 486 72 
<< m1 >>
rect 487 71 488 72 
<< m2 >>
rect 487 71 488 72 
<< pdiffusion >>
rect 498 71 499 72 
<< pdiffusion >>
rect 499 71 500 72 
<< pdiffusion >>
rect 500 71 501 72 
<< pdiffusion >>
rect 501 71 502 72 
<< pdiffusion >>
rect 502 71 503 72 
<< pdiffusion >>
rect 503 71 504 72 
<< pdiffusion >>
rect 516 71 517 72 
<< pdiffusion >>
rect 517 71 518 72 
<< pdiffusion >>
rect 518 71 519 72 
<< pdiffusion >>
rect 519 71 520 72 
<< m1 >>
rect 520 71 521 72 
<< pdiffusion >>
rect 520 71 521 72 
<< pdiffusion >>
rect 521 71 522 72 
<< m1 >>
rect 28 72 29 73 
<< m1 >>
rect 64 72 65 73 
<< m1 >>
rect 92 72 93 73 
<< m1 >>
rect 100 72 101 73 
<< m2 >>
rect 100 72 101 73 
<< m1 >>
rect 124 72 125 73 
<< m1 >>
rect 129 72 130 73 
<< m1 >>
rect 131 72 132 73 
<< m1 >>
rect 142 72 143 73 
<< m2 >>
rect 145 72 146 73 
<< m1 >>
rect 160 72 161 73 
<< m1 >>
rect 199 72 200 73 
<< m1 >>
rect 201 72 202 73 
<< m2 >>
rect 202 72 203 73 
<< m1 >>
rect 214 72 215 73 
<< m1 >>
rect 235 72 236 73 
<< m2 >>
rect 235 72 236 73 
<< m1 >>
rect 237 72 238 73 
<< m1 >>
rect 247 72 248 73 
<< m1 >>
rect 253 72 254 73 
<< m1 >>
rect 255 72 256 73 
<< m1 >>
rect 280 72 281 73 
<< m1 >>
rect 289 72 290 73 
<< m1 >>
rect 332 72 333 73 
<< m1 >>
rect 334 72 335 73 
<< m1 >>
rect 340 72 341 73 
<< m1 >>
rect 358 72 359 73 
<< m1 >>
rect 366 72 367 73 
<< m1 >>
rect 370 72 371 73 
<< m1 >>
rect 415 72 416 73 
<< m1 >>
rect 433 72 434 73 
<< m1 >>
rect 487 72 488 73 
<< m2 >>
rect 487 72 488 73 
<< m1 >>
rect 520 72 521 73 
<< m1 >>
rect 28 73 29 74 
<< m1 >>
rect 64 73 65 74 
<< m1 >>
rect 92 73 93 74 
<< m1 >>
rect 100 73 101 74 
<< m2 >>
rect 100 73 101 74 
<< m1 >>
rect 124 73 125 74 
<< m1 >>
rect 125 73 126 74 
<< m1 >>
rect 126 73 127 74 
<< m1 >>
rect 127 73 128 74 
<< m1 >>
rect 129 73 130 74 
<< m1 >>
rect 131 73 132 74 
<< m1 >>
rect 142 73 143 74 
<< m1 >>
rect 143 73 144 74 
<< m1 >>
rect 144 73 145 74 
<< m1 >>
rect 145 73 146 74 
<< m2 >>
rect 145 73 146 74 
<< m1 >>
rect 160 73 161 74 
<< m1 >>
rect 161 73 162 74 
<< m1 >>
rect 162 73 163 74 
<< m1 >>
rect 163 73 164 74 
<< m1 >>
rect 197 73 198 74 
<< m2 >>
rect 197 73 198 74 
<< m2c >>
rect 197 73 198 74 
<< m1 >>
rect 197 73 198 74 
<< m2 >>
rect 197 73 198 74 
<< m2 >>
rect 198 73 199 74 
<< m1 >>
rect 199 73 200 74 
<< m2 >>
rect 199 73 200 74 
<< m2 >>
rect 200 73 201 74 
<< m1 >>
rect 201 73 202 74 
<< m2 >>
rect 201 73 202 74 
<< m2 >>
rect 202 73 203 74 
<< m1 >>
rect 214 73 215 74 
<< m1 >>
rect 235 73 236 74 
<< m2 >>
rect 235 73 236 74 
<< m1 >>
rect 237 73 238 74 
<< m1 >>
rect 247 73 248 74 
<< m1 >>
rect 253 73 254 74 
<< m1 >>
rect 255 73 256 74 
<< m1 >>
rect 280 73 281 74 
<< m1 >>
rect 289 73 290 74 
<< m1 >>
rect 332 73 333 74 
<< m1 >>
rect 334 73 335 74 
<< m1 >>
rect 340 73 341 74 
<< m1 >>
rect 358 73 359 74 
<< m1 >>
rect 366 73 367 74 
<< m1 >>
rect 370 73 371 74 
<< m1 >>
rect 415 73 416 74 
<< m1 >>
rect 433 73 434 74 
<< m1 >>
rect 487 73 488 74 
<< m2 >>
rect 487 73 488 74 
<< m1 >>
rect 520 73 521 74 
<< m1 >>
rect 28 74 29 75 
<< m1 >>
rect 64 74 65 75 
<< m1 >>
rect 92 74 93 75 
<< m1 >>
rect 100 74 101 75 
<< m2 >>
rect 100 74 101 75 
<< m1 >>
rect 127 74 128 75 
<< m1 >>
rect 129 74 130 75 
<< m1 >>
rect 131 74 132 75 
<< m1 >>
rect 145 74 146 75 
<< m2 >>
rect 145 74 146 75 
<< m1 >>
rect 163 74 164 75 
<< m1 >>
rect 197 74 198 75 
<< m1 >>
rect 199 74 200 75 
<< m1 >>
rect 201 74 202 75 
<< m1 >>
rect 214 74 215 75 
<< m1 >>
rect 235 74 236 75 
<< m2 >>
rect 235 74 236 75 
<< m1 >>
rect 237 74 238 75 
<< m1 >>
rect 247 74 248 75 
<< m1 >>
rect 253 74 254 75 
<< m1 >>
rect 255 74 256 75 
<< m1 >>
rect 280 74 281 75 
<< m1 >>
rect 289 74 290 75 
<< m1 >>
rect 332 74 333 75 
<< m1 >>
rect 334 74 335 75 
<< m1 >>
rect 340 74 341 75 
<< m1 >>
rect 358 74 359 75 
<< m1 >>
rect 366 74 367 75 
<< m1 >>
rect 370 74 371 75 
<< m1 >>
rect 415 74 416 75 
<< m1 >>
rect 433 74 434 75 
<< m1 >>
rect 487 74 488 75 
<< m2 >>
rect 487 74 488 75 
<< m1 >>
rect 520 74 521 75 
<< m1 >>
rect 28 75 29 76 
<< m1 >>
rect 64 75 65 76 
<< m1 >>
rect 92 75 93 76 
<< m1 >>
rect 100 75 101 76 
<< m2 >>
rect 100 75 101 76 
<< m1 >>
rect 127 75 128 76 
<< m1 >>
rect 129 75 130 76 
<< m1 >>
rect 131 75 132 76 
<< m1 >>
rect 145 75 146 76 
<< m2 >>
rect 145 75 146 76 
<< m1 >>
rect 163 75 164 76 
<< m1 >>
rect 197 75 198 76 
<< m1 >>
rect 199 75 200 76 
<< m1 >>
rect 201 75 202 76 
<< m1 >>
rect 214 75 215 76 
<< m1 >>
rect 235 75 236 76 
<< m2 >>
rect 235 75 236 76 
<< m1 >>
rect 237 75 238 76 
<< m1 >>
rect 247 75 248 76 
<< m1 >>
rect 253 75 254 76 
<< m1 >>
rect 255 75 256 76 
<< m1 >>
rect 280 75 281 76 
<< m1 >>
rect 289 75 290 76 
<< m1 >>
rect 332 75 333 76 
<< m2 >>
rect 332 75 333 76 
<< m2c >>
rect 332 75 333 76 
<< m1 >>
rect 332 75 333 76 
<< m2 >>
rect 332 75 333 76 
<< m2 >>
rect 333 75 334 76 
<< m1 >>
rect 334 75 335 76 
<< m2 >>
rect 334 75 335 76 
<< m2 >>
rect 335 75 336 76 
<< m1 >>
rect 336 75 337 76 
<< m2 >>
rect 336 75 337 76 
<< m2c >>
rect 336 75 337 76 
<< m1 >>
rect 336 75 337 76 
<< m2 >>
rect 336 75 337 76 
<< m1 >>
rect 340 75 341 76 
<< m1 >>
rect 358 75 359 76 
<< m1 >>
rect 366 75 367 76 
<< m1 >>
rect 370 75 371 76 
<< m1 >>
rect 415 75 416 76 
<< m1 >>
rect 433 75 434 76 
<< m1 >>
rect 487 75 488 76 
<< m2 >>
rect 487 75 488 76 
<< m1 >>
rect 520 75 521 76 
<< m1 >>
rect 28 76 29 77 
<< m1 >>
rect 64 76 65 77 
<< m1 >>
rect 92 76 93 77 
<< m1 >>
rect 100 76 101 77 
<< m2 >>
rect 100 76 101 77 
<< m1 >>
rect 127 76 128 77 
<< m1 >>
rect 129 76 130 77 
<< m1 >>
rect 131 76 132 77 
<< m1 >>
rect 145 76 146 77 
<< m2 >>
rect 145 76 146 77 
<< m1 >>
rect 163 76 164 77 
<< m1 >>
rect 185 76 186 77 
<< m2 >>
rect 185 76 186 77 
<< m2c >>
rect 185 76 186 77 
<< m1 >>
rect 185 76 186 77 
<< m2 >>
rect 185 76 186 77 
<< m2 >>
rect 186 76 187 77 
<< m1 >>
rect 187 76 188 77 
<< m2 >>
rect 187 76 188 77 
<< m1 >>
rect 188 76 189 77 
<< m2 >>
rect 188 76 189 77 
<< m1 >>
rect 189 76 190 77 
<< m2 >>
rect 189 76 190 77 
<< m1 >>
rect 190 76 191 77 
<< m2 >>
rect 190 76 191 77 
<< m1 >>
rect 191 76 192 77 
<< m2 >>
rect 191 76 192 77 
<< m1 >>
rect 192 76 193 77 
<< m2 >>
rect 192 76 193 77 
<< m1 >>
rect 193 76 194 77 
<< m2 >>
rect 193 76 194 77 
<< m1 >>
rect 194 76 195 77 
<< m2 >>
rect 194 76 195 77 
<< m1 >>
rect 195 76 196 77 
<< m2 >>
rect 195 76 196 77 
<< m1 >>
rect 196 76 197 77 
<< m2 >>
rect 196 76 197 77 
<< m1 >>
rect 197 76 198 77 
<< m2 >>
rect 197 76 198 77 
<< m2 >>
rect 198 76 199 77 
<< m1 >>
rect 199 76 200 77 
<< m2 >>
rect 199 76 200 77 
<< m2 >>
rect 200 76 201 77 
<< m1 >>
rect 201 76 202 77 
<< m2 >>
rect 201 76 202 77 
<< m2 >>
rect 202 76 203 77 
<< m1 >>
rect 203 76 204 77 
<< m2 >>
rect 203 76 204 77 
<< m2c >>
rect 203 76 204 77 
<< m1 >>
rect 203 76 204 77 
<< m2 >>
rect 203 76 204 77 
<< m1 >>
rect 204 76 205 77 
<< m1 >>
rect 205 76 206 77 
<< m1 >>
rect 206 76 207 77 
<< m1 >>
rect 207 76 208 77 
<< m1 >>
rect 208 76 209 77 
<< m1 >>
rect 209 76 210 77 
<< m1 >>
rect 210 76 211 77 
<< m1 >>
rect 211 76 212 77 
<< m1 >>
rect 212 76 213 77 
<< m2 >>
rect 212 76 213 77 
<< m2c >>
rect 212 76 213 77 
<< m1 >>
rect 212 76 213 77 
<< m2 >>
rect 212 76 213 77 
<< m2 >>
rect 213 76 214 77 
<< m1 >>
rect 214 76 215 77 
<< m2 >>
rect 214 76 215 77 
<< m2 >>
rect 215 76 216 77 
<< m1 >>
rect 216 76 217 77 
<< m2 >>
rect 216 76 217 77 
<< m2c >>
rect 216 76 217 77 
<< m1 >>
rect 216 76 217 77 
<< m2 >>
rect 216 76 217 77 
<< m1 >>
rect 217 76 218 77 
<< m1 >>
rect 218 76 219 77 
<< m1 >>
rect 219 76 220 77 
<< m1 >>
rect 220 76 221 77 
<< m1 >>
rect 221 76 222 77 
<< m1 >>
rect 222 76 223 77 
<< m2 >>
rect 222 76 223 77 
<< m2c >>
rect 222 76 223 77 
<< m1 >>
rect 222 76 223 77 
<< m2 >>
rect 222 76 223 77 
<< m2 >>
rect 223 76 224 77 
<< m2 >>
rect 224 76 225 77 
<< m2 >>
rect 225 76 226 77 
<< m2 >>
rect 226 76 227 77 
<< m2 >>
rect 227 76 228 77 
<< m2 >>
rect 228 76 229 77 
<< m2 >>
rect 229 76 230 77 
<< m2 >>
rect 230 76 231 77 
<< m2 >>
rect 231 76 232 77 
<< m2 >>
rect 232 76 233 77 
<< m2 >>
rect 233 76 234 77 
<< m2 >>
rect 234 76 235 77 
<< m1 >>
rect 235 76 236 77 
<< m2 >>
rect 235 76 236 77 
<< m1 >>
rect 237 76 238 77 
<< m1 >>
rect 247 76 248 77 
<< m1 >>
rect 253 76 254 77 
<< m1 >>
rect 255 76 256 77 
<< m1 >>
rect 280 76 281 77 
<< m1 >>
rect 289 76 290 77 
<< m1 >>
rect 334 76 335 77 
<< m1 >>
rect 336 76 337 77 
<< m1 >>
rect 340 76 341 77 
<< m1 >>
rect 358 76 359 77 
<< m1 >>
rect 366 76 367 77 
<< m1 >>
rect 370 76 371 77 
<< m1 >>
rect 415 76 416 77 
<< m1 >>
rect 433 76 434 77 
<< m1 >>
rect 487 76 488 77 
<< m2 >>
rect 487 76 488 77 
<< m1 >>
rect 517 76 518 77 
<< m1 >>
rect 518 76 519 77 
<< m1 >>
rect 519 76 520 77 
<< m1 >>
rect 520 76 521 77 
<< m1 >>
rect 28 77 29 78 
<< m1 >>
rect 64 77 65 78 
<< m1 >>
rect 92 77 93 78 
<< m1 >>
rect 100 77 101 78 
<< m2 >>
rect 100 77 101 78 
<< m1 >>
rect 127 77 128 78 
<< m1 >>
rect 129 77 130 78 
<< m1 >>
rect 131 77 132 78 
<< m1 >>
rect 145 77 146 78 
<< m2 >>
rect 145 77 146 78 
<< m1 >>
rect 163 77 164 78 
<< m1 >>
rect 185 77 186 78 
<< m1 >>
rect 187 77 188 78 
<< m1 >>
rect 199 77 200 78 
<< m1 >>
rect 201 77 202 78 
<< m1 >>
rect 214 77 215 78 
<< m1 >>
rect 224 77 225 78 
<< m1 >>
rect 225 77 226 78 
<< m1 >>
rect 226 77 227 78 
<< m1 >>
rect 227 77 228 78 
<< m1 >>
rect 228 77 229 78 
<< m1 >>
rect 229 77 230 78 
<< m1 >>
rect 230 77 231 78 
<< m1 >>
rect 231 77 232 78 
<< m1 >>
rect 232 77 233 78 
<< m1 >>
rect 233 77 234 78 
<< m1 >>
rect 234 77 235 78 
<< m1 >>
rect 235 77 236 78 
<< m1 >>
rect 237 77 238 78 
<< m2 >>
rect 237 77 238 78 
<< m2c >>
rect 237 77 238 78 
<< m1 >>
rect 237 77 238 78 
<< m2 >>
rect 237 77 238 78 
<< m1 >>
rect 247 77 248 78 
<< m2 >>
rect 247 77 248 78 
<< m2c >>
rect 247 77 248 78 
<< m1 >>
rect 247 77 248 78 
<< m2 >>
rect 247 77 248 78 
<< m1 >>
rect 253 77 254 78 
<< m2 >>
rect 253 77 254 78 
<< m2c >>
rect 253 77 254 78 
<< m1 >>
rect 253 77 254 78 
<< m2 >>
rect 253 77 254 78 
<< m1 >>
rect 255 77 256 78 
<< m2 >>
rect 255 77 256 78 
<< m2c >>
rect 255 77 256 78 
<< m1 >>
rect 255 77 256 78 
<< m2 >>
rect 255 77 256 78 
<< m1 >>
rect 280 77 281 78 
<< m2 >>
rect 280 77 281 78 
<< m2c >>
rect 280 77 281 78 
<< m1 >>
rect 280 77 281 78 
<< m2 >>
rect 280 77 281 78 
<< m1 >>
rect 289 77 290 78 
<< m2 >>
rect 289 77 290 78 
<< m2c >>
rect 289 77 290 78 
<< m1 >>
rect 289 77 290 78 
<< m2 >>
rect 289 77 290 78 
<< m1 >>
rect 334 77 335 78 
<< m2 >>
rect 334 77 335 78 
<< m2c >>
rect 334 77 335 78 
<< m1 >>
rect 334 77 335 78 
<< m2 >>
rect 334 77 335 78 
<< m1 >>
rect 336 77 337 78 
<< m1 >>
rect 337 77 338 78 
<< m1 >>
rect 338 77 339 78 
<< m2 >>
rect 338 77 339 78 
<< m2c >>
rect 338 77 339 78 
<< m1 >>
rect 338 77 339 78 
<< m2 >>
rect 338 77 339 78 
<< m2 >>
rect 339 77 340 78 
<< m1 >>
rect 340 77 341 78 
<< m2 >>
rect 340 77 341 78 
<< m2 >>
rect 341 77 342 78 
<< m1 >>
rect 344 77 345 78 
<< m2 >>
rect 344 77 345 78 
<< m2c >>
rect 344 77 345 78 
<< m1 >>
rect 344 77 345 78 
<< m2 >>
rect 344 77 345 78 
<< m1 >>
rect 345 77 346 78 
<< m1 >>
rect 346 77 347 78 
<< m1 >>
rect 347 77 348 78 
<< m1 >>
rect 348 77 349 78 
<< m1 >>
rect 349 77 350 78 
<< m1 >>
rect 350 77 351 78 
<< m1 >>
rect 351 77 352 78 
<< m1 >>
rect 352 77 353 78 
<< m1 >>
rect 353 77 354 78 
<< m1 >>
rect 354 77 355 78 
<< m1 >>
rect 355 77 356 78 
<< m1 >>
rect 356 77 357 78 
<< m1 >>
rect 357 77 358 78 
<< m1 >>
rect 358 77 359 78 
<< m1 >>
rect 366 77 367 78 
<< m1 >>
rect 370 77 371 78 
<< m1 >>
rect 415 77 416 78 
<< m1 >>
rect 433 77 434 78 
<< m1 >>
rect 487 77 488 78 
<< m2 >>
rect 487 77 488 78 
<< m1 >>
rect 517 77 518 78 
<< m1 >>
rect 28 78 29 79 
<< m1 >>
rect 64 78 65 79 
<< m1 >>
rect 92 78 93 79 
<< m1 >>
rect 100 78 101 79 
<< m2 >>
rect 100 78 101 79 
<< m1 >>
rect 127 78 128 79 
<< m1 >>
rect 129 78 130 79 
<< m1 >>
rect 131 78 132 79 
<< m1 >>
rect 145 78 146 79 
<< m2 >>
rect 145 78 146 79 
<< m1 >>
rect 163 78 164 79 
<< m1 >>
rect 185 78 186 79 
<< m1 >>
rect 187 78 188 79 
<< m1 >>
rect 199 78 200 79 
<< m1 >>
rect 201 78 202 79 
<< m1 >>
rect 214 78 215 79 
<< m1 >>
rect 224 78 225 79 
<< m2 >>
rect 237 78 238 79 
<< m2 >>
rect 238 78 239 79 
<< m2 >>
rect 239 78 240 79 
<< m2 >>
rect 247 78 248 79 
<< m2 >>
rect 248 78 249 79 
<< m2 >>
rect 253 78 254 79 
<< m2 >>
rect 255 78 256 79 
<< m2 >>
rect 280 78 281 79 
<< m2 >>
rect 289 78 290 79 
<< m2 >>
rect 290 78 291 79 
<< m2 >>
rect 291 78 292 79 
<< m2 >>
rect 292 78 293 79 
<< m2 >>
rect 293 78 294 79 
<< m2 >>
rect 294 78 295 79 
<< m2 >>
rect 295 78 296 79 
<< m2 >>
rect 296 78 297 79 
<< m2 >>
rect 297 78 298 79 
<< m2 >>
rect 298 78 299 79 
<< m2 >>
rect 299 78 300 79 
<< m2 >>
rect 300 78 301 79 
<< m2 >>
rect 301 78 302 79 
<< m2 >>
rect 302 78 303 79 
<< m2 >>
rect 334 78 335 79 
<< m1 >>
rect 340 78 341 79 
<< m2 >>
rect 341 78 342 79 
<< m2 >>
rect 344 78 345 79 
<< m1 >>
rect 366 78 367 79 
<< m1 >>
rect 370 78 371 79 
<< m1 >>
rect 415 78 416 79 
<< m1 >>
rect 433 78 434 79 
<< m1 >>
rect 487 78 488 79 
<< m2 >>
rect 487 78 488 79 
<< m1 >>
rect 517 78 518 79 
<< m1 >>
rect 28 79 29 80 
<< m1 >>
rect 29 79 30 80 
<< m1 >>
rect 30 79 31 80 
<< m1 >>
rect 31 79 32 80 
<< m1 >>
rect 32 79 33 80 
<< m1 >>
rect 33 79 34 80 
<< m1 >>
rect 34 79 35 80 
<< m1 >>
rect 64 79 65 80 
<< m1 >>
rect 92 79 93 80 
<< m1 >>
rect 100 79 101 80 
<< m2 >>
rect 100 79 101 80 
<< m1 >>
rect 127 79 128 80 
<< m1 >>
rect 129 79 130 80 
<< m1 >>
rect 131 79 132 80 
<< m1 >>
rect 145 79 146 80 
<< m2 >>
rect 145 79 146 80 
<< m1 >>
rect 163 79 164 80 
<< m1 >>
rect 185 79 186 80 
<< m1 >>
rect 187 79 188 80 
<< m1 >>
rect 199 79 200 80 
<< m1 >>
rect 201 79 202 80 
<< m1 >>
rect 203 79 204 80 
<< m1 >>
rect 204 79 205 80 
<< m1 >>
rect 205 79 206 80 
<< m1 >>
rect 206 79 207 80 
<< m1 >>
rect 207 79 208 80 
<< m1 >>
rect 208 79 209 80 
<< m1 >>
rect 209 79 210 80 
<< m1 >>
rect 210 79 211 80 
<< m1 >>
rect 211 79 212 80 
<< m1 >>
rect 212 79 213 80 
<< m2 >>
rect 212 79 213 80 
<< m2c >>
rect 212 79 213 80 
<< m1 >>
rect 212 79 213 80 
<< m2 >>
rect 212 79 213 80 
<< m2 >>
rect 213 79 214 80 
<< m1 >>
rect 214 79 215 80 
<< m2 >>
rect 214 79 215 80 
<< m2 >>
rect 215 79 216 80 
<< m1 >>
rect 216 79 217 80 
<< m2 >>
rect 216 79 217 80 
<< m2c >>
rect 216 79 217 80 
<< m1 >>
rect 216 79 217 80 
<< m2 >>
rect 216 79 217 80 
<< m1 >>
rect 217 79 218 80 
<< m1 >>
rect 218 79 219 80 
<< m1 >>
rect 219 79 220 80 
<< m1 >>
rect 220 79 221 80 
<< m1 >>
rect 221 79 222 80 
<< m1 >>
rect 222 79 223 80 
<< m2 >>
rect 222 79 223 80 
<< m2c >>
rect 222 79 223 80 
<< m1 >>
rect 222 79 223 80 
<< m2 >>
rect 222 79 223 80 
<< m2 >>
rect 223 79 224 80 
<< m1 >>
rect 224 79 225 80 
<< m2 >>
rect 224 79 225 80 
<< m2 >>
rect 225 79 226 80 
<< m1 >>
rect 226 79 227 80 
<< m2 >>
rect 226 79 227 80 
<< m2c >>
rect 226 79 227 80 
<< m1 >>
rect 226 79 227 80 
<< m2 >>
rect 226 79 227 80 
<< m1 >>
rect 227 79 228 80 
<< m1 >>
rect 228 79 229 80 
<< m1 >>
rect 229 79 230 80 
<< m1 >>
rect 230 79 231 80 
<< m1 >>
rect 231 79 232 80 
<< m1 >>
rect 232 79 233 80 
<< m1 >>
rect 235 79 236 80 
<< m1 >>
rect 236 79 237 80 
<< m1 >>
rect 237 79 238 80 
<< m1 >>
rect 238 79 239 80 
<< m1 >>
rect 239 79 240 80 
<< m2 >>
rect 239 79 240 80 
<< m1 >>
rect 240 79 241 80 
<< m1 >>
rect 241 79 242 80 
<< m1 >>
rect 242 79 243 80 
<< m1 >>
rect 243 79 244 80 
<< m1 >>
rect 244 79 245 80 
<< m1 >>
rect 245 79 246 80 
<< m1 >>
rect 246 79 247 80 
<< m1 >>
rect 247 79 248 80 
<< m1 >>
rect 248 79 249 80 
<< m2 >>
rect 248 79 249 80 
<< m1 >>
rect 249 79 250 80 
<< m1 >>
rect 250 79 251 80 
<< m1 >>
rect 251 79 252 80 
<< m1 >>
rect 252 79 253 80 
<< m1 >>
rect 253 79 254 80 
<< m2 >>
rect 253 79 254 80 
<< m1 >>
rect 254 79 255 80 
<< m1 >>
rect 255 79 256 80 
<< m2 >>
rect 255 79 256 80 
<< m1 >>
rect 256 79 257 80 
<< m1 >>
rect 257 79 258 80 
<< m1 >>
rect 258 79 259 80 
<< m1 >>
rect 259 79 260 80 
<< m1 >>
rect 260 79 261 80 
<< m1 >>
rect 261 79 262 80 
<< m1 >>
rect 262 79 263 80 
<< m1 >>
rect 263 79 264 80 
<< m1 >>
rect 264 79 265 80 
<< m1 >>
rect 265 79 266 80 
<< m1 >>
rect 266 79 267 80 
<< m1 >>
rect 267 79 268 80 
<< m1 >>
rect 268 79 269 80 
<< m1 >>
rect 269 79 270 80 
<< m1 >>
rect 270 79 271 80 
<< m1 >>
rect 271 79 272 80 
<< m1 >>
rect 272 79 273 80 
<< m1 >>
rect 273 79 274 80 
<< m1 >>
rect 274 79 275 80 
<< m1 >>
rect 275 79 276 80 
<< m1 >>
rect 276 79 277 80 
<< m1 >>
rect 277 79 278 80 
<< m1 >>
rect 278 79 279 80 
<< m1 >>
rect 279 79 280 80 
<< m1 >>
rect 280 79 281 80 
<< m2 >>
rect 280 79 281 80 
<< m1 >>
rect 281 79 282 80 
<< m1 >>
rect 282 79 283 80 
<< m1 >>
rect 283 79 284 80 
<< m1 >>
rect 284 79 285 80 
<< m1 >>
rect 285 79 286 80 
<< m1 >>
rect 286 79 287 80 
<< m1 >>
rect 287 79 288 80 
<< m1 >>
rect 288 79 289 80 
<< m1 >>
rect 289 79 290 80 
<< m1 >>
rect 290 79 291 80 
<< m1 >>
rect 291 79 292 80 
<< m1 >>
rect 292 79 293 80 
<< m1 >>
rect 293 79 294 80 
<< m1 >>
rect 294 79 295 80 
<< m1 >>
rect 295 79 296 80 
<< m1 >>
rect 296 79 297 80 
<< m1 >>
rect 297 79 298 80 
<< m1 >>
rect 298 79 299 80 
<< m1 >>
rect 299 79 300 80 
<< m1 >>
rect 300 79 301 80 
<< m1 >>
rect 301 79 302 80 
<< m1 >>
rect 302 79 303 80 
<< m2 >>
rect 302 79 303 80 
<< m1 >>
rect 303 79 304 80 
<< m1 >>
rect 304 79 305 80 
<< m1 >>
rect 305 79 306 80 
<< m1 >>
rect 306 79 307 80 
<< m1 >>
rect 307 79 308 80 
<< m1 >>
rect 308 79 309 80 
<< m1 >>
rect 309 79 310 80 
<< m1 >>
rect 310 79 311 80 
<< m1 >>
rect 311 79 312 80 
<< m1 >>
rect 312 79 313 80 
<< m1 >>
rect 313 79 314 80 
<< m1 >>
rect 314 79 315 80 
<< m1 >>
rect 315 79 316 80 
<< m1 >>
rect 316 79 317 80 
<< m1 >>
rect 317 79 318 80 
<< m1 >>
rect 318 79 319 80 
<< m1 >>
rect 319 79 320 80 
<< m1 >>
rect 320 79 321 80 
<< m1 >>
rect 321 79 322 80 
<< m1 >>
rect 322 79 323 80 
<< m1 >>
rect 323 79 324 80 
<< m1 >>
rect 324 79 325 80 
<< m1 >>
rect 325 79 326 80 
<< m1 >>
rect 326 79 327 80 
<< m1 >>
rect 327 79 328 80 
<< m1 >>
rect 328 79 329 80 
<< m1 >>
rect 329 79 330 80 
<< m1 >>
rect 330 79 331 80 
<< m1 >>
rect 331 79 332 80 
<< m1 >>
rect 332 79 333 80 
<< m1 >>
rect 333 79 334 80 
<< m1 >>
rect 334 79 335 80 
<< m2 >>
rect 334 79 335 80 
<< m1 >>
rect 335 79 336 80 
<< m1 >>
rect 336 79 337 80 
<< m1 >>
rect 337 79 338 80 
<< m1 >>
rect 338 79 339 80 
<< m1 >>
rect 339 79 340 80 
<< m1 >>
rect 340 79 341 80 
<< m2 >>
rect 341 79 342 80 
<< m1 >>
rect 342 79 343 80 
<< m2 >>
rect 342 79 343 80 
<< m2c >>
rect 342 79 343 80 
<< m1 >>
rect 342 79 343 80 
<< m2 >>
rect 342 79 343 80 
<< m1 >>
rect 343 79 344 80 
<< m1 >>
rect 344 79 345 80 
<< m2 >>
rect 344 79 345 80 
<< m1 >>
rect 345 79 346 80 
<< m1 >>
rect 346 79 347 80 
<< m1 >>
rect 347 79 348 80 
<< m1 >>
rect 348 79 349 80 
<< m1 >>
rect 349 79 350 80 
<< m1 >>
rect 350 79 351 80 
<< m1 >>
rect 351 79 352 80 
<< m1 >>
rect 352 79 353 80 
<< m1 >>
rect 353 79 354 80 
<< m1 >>
rect 354 79 355 80 
<< m1 >>
rect 355 79 356 80 
<< m1 >>
rect 356 79 357 80 
<< m1 >>
rect 357 79 358 80 
<< m1 >>
rect 358 79 359 80 
<< m1 >>
rect 364 79 365 80 
<< m2 >>
rect 364 79 365 80 
<< m2c >>
rect 364 79 365 80 
<< m1 >>
rect 364 79 365 80 
<< m2 >>
rect 364 79 365 80 
<< m2 >>
rect 365 79 366 80 
<< m1 >>
rect 366 79 367 80 
<< m2 >>
rect 366 79 367 80 
<< m2 >>
rect 367 79 368 80 
<< m1 >>
rect 368 79 369 80 
<< m2 >>
rect 368 79 369 80 
<< m2c >>
rect 368 79 369 80 
<< m1 >>
rect 368 79 369 80 
<< m2 >>
rect 368 79 369 80 
<< m2 >>
rect 369 79 370 80 
<< m1 >>
rect 370 79 371 80 
<< m2 >>
rect 370 79 371 80 
<< m2 >>
rect 371 79 372 80 
<< m1 >>
rect 372 79 373 80 
<< m2 >>
rect 372 79 373 80 
<< m2c >>
rect 372 79 373 80 
<< m1 >>
rect 372 79 373 80 
<< m2 >>
rect 372 79 373 80 
<< m1 >>
rect 373 79 374 80 
<< m1 >>
rect 374 79 375 80 
<< m1 >>
rect 375 79 376 80 
<< m1 >>
rect 376 79 377 80 
<< m1 >>
rect 377 79 378 80 
<< m1 >>
rect 378 79 379 80 
<< m1 >>
rect 379 79 380 80 
<< m1 >>
rect 380 79 381 80 
<< m1 >>
rect 381 79 382 80 
<< m1 >>
rect 382 79 383 80 
<< m1 >>
rect 383 79 384 80 
<< m1 >>
rect 384 79 385 80 
<< m1 >>
rect 385 79 386 80 
<< m1 >>
rect 386 79 387 80 
<< m1 >>
rect 387 79 388 80 
<< m1 >>
rect 388 79 389 80 
<< m1 >>
rect 389 79 390 80 
<< m1 >>
rect 390 79 391 80 
<< m1 >>
rect 391 79 392 80 
<< m1 >>
rect 392 79 393 80 
<< m1 >>
rect 393 79 394 80 
<< m1 >>
rect 394 79 395 80 
<< m1 >>
rect 395 79 396 80 
<< m1 >>
rect 396 79 397 80 
<< m1 >>
rect 397 79 398 80 
<< m1 >>
rect 398 79 399 80 
<< m1 >>
rect 399 79 400 80 
<< m1 >>
rect 400 79 401 80 
<< m1 >>
rect 401 79 402 80 
<< m1 >>
rect 402 79 403 80 
<< m1 >>
rect 403 79 404 80 
<< m1 >>
rect 404 79 405 80 
<< m1 >>
rect 405 79 406 80 
<< m1 >>
rect 406 79 407 80 
<< m1 >>
rect 407 79 408 80 
<< m1 >>
rect 408 79 409 80 
<< m1 >>
rect 409 79 410 80 
<< m1 >>
rect 410 79 411 80 
<< m1 >>
rect 411 79 412 80 
<< m1 >>
rect 412 79 413 80 
<< m1 >>
rect 413 79 414 80 
<< m1 >>
rect 415 79 416 80 
<< m1 >>
rect 433 79 434 80 
<< m1 >>
rect 487 79 488 80 
<< m2 >>
rect 487 79 488 80 
<< m1 >>
rect 517 79 518 80 
<< m1 >>
rect 34 80 35 81 
<< m1 >>
rect 64 80 65 81 
<< m1 >>
rect 92 80 93 81 
<< m1 >>
rect 100 80 101 81 
<< m2 >>
rect 100 80 101 81 
<< m1 >>
rect 127 80 128 81 
<< m1 >>
rect 129 80 130 81 
<< m1 >>
rect 131 80 132 81 
<< m1 >>
rect 145 80 146 81 
<< m2 >>
rect 145 80 146 81 
<< m1 >>
rect 163 80 164 81 
<< m1 >>
rect 185 80 186 81 
<< m1 >>
rect 187 80 188 81 
<< m1 >>
rect 193 80 194 81 
<< m1 >>
rect 194 80 195 81 
<< m1 >>
rect 195 80 196 81 
<< m1 >>
rect 196 80 197 81 
<< m1 >>
rect 197 80 198 81 
<< m2 >>
rect 197 80 198 81 
<< m2c >>
rect 197 80 198 81 
<< m1 >>
rect 197 80 198 81 
<< m2 >>
rect 197 80 198 81 
<< m2 >>
rect 198 80 199 81 
<< m1 >>
rect 199 80 200 81 
<< m2 >>
rect 199 80 200 81 
<< m2 >>
rect 200 80 201 81 
<< m1 >>
rect 201 80 202 81 
<< m2 >>
rect 201 80 202 81 
<< m2 >>
rect 202 80 203 81 
<< m1 >>
rect 203 80 204 81 
<< m2 >>
rect 203 80 204 81 
<< m2c >>
rect 203 80 204 81 
<< m1 >>
rect 203 80 204 81 
<< m2 >>
rect 203 80 204 81 
<< m1 >>
rect 214 80 215 81 
<< m1 >>
rect 224 80 225 81 
<< m1 >>
rect 232 80 233 81 
<< m1 >>
rect 235 80 236 81 
<< m2 >>
rect 239 80 240 81 
<< m2 >>
rect 248 80 249 81 
<< m2 >>
rect 253 80 254 81 
<< m2 >>
rect 255 80 256 81 
<< m2 >>
rect 280 80 281 81 
<< m2 >>
rect 302 80 303 81 
<< m2 >>
rect 334 80 335 81 
<< m2 >>
rect 344 80 345 81 
<< m1 >>
rect 358 80 359 81 
<< m1 >>
rect 364 80 365 81 
<< m1 >>
rect 366 80 367 81 
<< m1 >>
rect 370 80 371 81 
<< m1 >>
rect 413 80 414 81 
<< m1 >>
rect 415 80 416 81 
<< m1 >>
rect 433 80 434 81 
<< m1 >>
rect 487 80 488 81 
<< m2 >>
rect 487 80 488 81 
<< m1 >>
rect 517 80 518 81 
<< m1 >>
rect 34 81 35 82 
<< m1 >>
rect 64 81 65 82 
<< m1 >>
rect 67 81 68 82 
<< m1 >>
rect 68 81 69 82 
<< m1 >>
rect 69 81 70 82 
<< m1 >>
rect 70 81 71 82 
<< m1 >>
rect 71 81 72 82 
<< m1 >>
rect 72 81 73 82 
<< m1 >>
rect 73 81 74 82 
<< m1 >>
rect 92 81 93 82 
<< m1 >>
rect 100 81 101 82 
<< m2 >>
rect 100 81 101 82 
<< m1 >>
rect 121 81 122 82 
<< m1 >>
rect 122 81 123 82 
<< m1 >>
rect 123 81 124 82 
<< m1 >>
rect 124 81 125 82 
<< m1 >>
rect 125 81 126 82 
<< m2 >>
rect 125 81 126 82 
<< m2c >>
rect 125 81 126 82 
<< m1 >>
rect 125 81 126 82 
<< m2 >>
rect 125 81 126 82 
<< m2 >>
rect 126 81 127 82 
<< m1 >>
rect 127 81 128 82 
<< m2 >>
rect 127 81 128 82 
<< m2 >>
rect 128 81 129 82 
<< m1 >>
rect 129 81 130 82 
<< m2 >>
rect 129 81 130 82 
<< m2 >>
rect 130 81 131 82 
<< m1 >>
rect 131 81 132 82 
<< m2 >>
rect 131 81 132 82 
<< m2 >>
rect 132 81 133 82 
<< m1 >>
rect 133 81 134 82 
<< m2 >>
rect 133 81 134 82 
<< m2c >>
rect 133 81 134 82 
<< m1 >>
rect 133 81 134 82 
<< m2 >>
rect 133 81 134 82 
<< m1 >>
rect 139 81 140 82 
<< m1 >>
rect 140 81 141 82 
<< m1 >>
rect 141 81 142 82 
<< m1 >>
rect 142 81 143 82 
<< m1 >>
rect 143 81 144 82 
<< m2 >>
rect 143 81 144 82 
<< m2c >>
rect 143 81 144 82 
<< m1 >>
rect 143 81 144 82 
<< m2 >>
rect 143 81 144 82 
<< m2 >>
rect 144 81 145 82 
<< m1 >>
rect 145 81 146 82 
<< m2 >>
rect 145 81 146 82 
<< m1 >>
rect 163 81 164 82 
<< m1 >>
rect 185 81 186 82 
<< m1 >>
rect 187 81 188 82 
<< m1 >>
rect 193 81 194 82 
<< m1 >>
rect 199 81 200 82 
<< m1 >>
rect 201 81 202 82 
<< m1 >>
rect 211 81 212 82 
<< m1 >>
rect 212 81 213 82 
<< m2 >>
rect 212 81 213 82 
<< m2c >>
rect 212 81 213 82 
<< m1 >>
rect 212 81 213 82 
<< m2 >>
rect 212 81 213 82 
<< m2 >>
rect 213 81 214 82 
<< m1 >>
rect 214 81 215 82 
<< m2 >>
rect 214 81 215 82 
<< m1 >>
rect 215 81 216 82 
<< m2 >>
rect 215 81 216 82 
<< m1 >>
rect 216 81 217 82 
<< m2 >>
rect 216 81 217 82 
<< m1 >>
rect 217 81 218 82 
<< m2 >>
rect 217 81 218 82 
<< m2 >>
rect 218 81 219 82 
<< m1 >>
rect 224 81 225 82 
<< m1 >>
rect 232 81 233 82 
<< m1 >>
rect 235 81 236 82 
<< m2 >>
rect 239 81 240 82 
<< m2 >>
rect 248 81 249 82 
<< m1 >>
rect 249 81 250 82 
<< m2 >>
rect 249 81 250 82 
<< m2c >>
rect 249 81 250 82 
<< m1 >>
rect 249 81 250 82 
<< m2 >>
rect 249 81 250 82 
<< m1 >>
rect 250 81 251 82 
<< m1 >>
rect 251 81 252 82 
<< m1 >>
rect 252 81 253 82 
<< m1 >>
rect 253 81 254 82 
<< m2 >>
rect 253 81 254 82 
<< m1 >>
rect 254 81 255 82 
<< m1 >>
rect 255 81 256 82 
<< m2 >>
rect 255 81 256 82 
<< m1 >>
rect 256 81 257 82 
<< m1 >>
rect 257 81 258 82 
<< m1 >>
rect 258 81 259 82 
<< m1 >>
rect 259 81 260 82 
<< m1 >>
rect 260 81 261 82 
<< m1 >>
rect 261 81 262 82 
<< m1 >>
rect 262 81 263 82 
<< m1 >>
rect 263 81 264 82 
<< m1 >>
rect 264 81 265 82 
<< m1 >>
rect 265 81 266 82 
<< m1 >>
rect 280 81 281 82 
<< m2 >>
rect 280 81 281 82 
<< m2c >>
rect 280 81 281 82 
<< m1 >>
rect 280 81 281 82 
<< m2 >>
rect 280 81 281 82 
<< m1 >>
rect 302 81 303 82 
<< m2 >>
rect 302 81 303 82 
<< m2c >>
rect 302 81 303 82 
<< m1 >>
rect 302 81 303 82 
<< m2 >>
rect 302 81 303 82 
<< m1 >>
rect 303 81 304 82 
<< m1 >>
rect 304 81 305 82 
<< m1 >>
rect 305 81 306 82 
<< m1 >>
rect 306 81 307 82 
<< m1 >>
rect 307 81 308 82 
<< m1 >>
rect 334 81 335 82 
<< m2 >>
rect 334 81 335 82 
<< m2c >>
rect 334 81 335 82 
<< m1 >>
rect 334 81 335 82 
<< m2 >>
rect 334 81 335 82 
<< m1 >>
rect 337 81 338 82 
<< m1 >>
rect 338 81 339 82 
<< m1 >>
rect 339 81 340 82 
<< m1 >>
rect 340 81 341 82 
<< m1 >>
rect 341 81 342 82 
<< m1 >>
rect 342 81 343 82 
<< m1 >>
rect 343 81 344 82 
<< m1 >>
rect 344 81 345 82 
<< m2 >>
rect 344 81 345 82 
<< m1 >>
rect 345 81 346 82 
<< m1 >>
rect 358 81 359 82 
<< m1 >>
rect 364 81 365 82 
<< m1 >>
rect 366 81 367 82 
<< m1 >>
rect 370 81 371 82 
<< m1 >>
rect 413 81 414 82 
<< m1 >>
rect 415 81 416 82 
<< m1 >>
rect 433 81 434 82 
<< m1 >>
rect 445 81 446 82 
<< m1 >>
rect 446 81 447 82 
<< m1 >>
rect 447 81 448 82 
<< m1 >>
rect 448 81 449 82 
<< m1 >>
rect 449 81 450 82 
<< m1 >>
rect 450 81 451 82 
<< m1 >>
rect 451 81 452 82 
<< m1 >>
rect 452 81 453 82 
<< m1 >>
rect 453 81 454 82 
<< m1 >>
rect 454 81 455 82 
<< m1 >>
rect 455 81 456 82 
<< m1 >>
rect 456 81 457 82 
<< m1 >>
rect 457 81 458 82 
<< m1 >>
rect 458 81 459 82 
<< m1 >>
rect 459 81 460 82 
<< m1 >>
rect 460 81 461 82 
<< m1 >>
rect 487 81 488 82 
<< m2 >>
rect 487 81 488 82 
<< m1 >>
rect 517 81 518 82 
<< m1 >>
rect 34 82 35 83 
<< m1 >>
rect 64 82 65 83 
<< m1 >>
rect 67 82 68 83 
<< m1 >>
rect 73 82 74 83 
<< m1 >>
rect 92 82 93 83 
<< m1 >>
rect 100 82 101 83 
<< m2 >>
rect 100 82 101 83 
<< m1 >>
rect 121 82 122 83 
<< m1 >>
rect 127 82 128 83 
<< m1 >>
rect 129 82 130 83 
<< m1 >>
rect 131 82 132 83 
<< m1 >>
rect 133 82 134 83 
<< m1 >>
rect 139 82 140 83 
<< m1 >>
rect 145 82 146 83 
<< m1 >>
rect 163 82 164 83 
<< m1 >>
rect 185 82 186 83 
<< m1 >>
rect 187 82 188 83 
<< m1 >>
rect 193 82 194 83 
<< m1 >>
rect 196 82 197 83 
<< m1 >>
rect 197 82 198 83 
<< m2 >>
rect 197 82 198 83 
<< m2c >>
rect 197 82 198 83 
<< m1 >>
rect 197 82 198 83 
<< m2 >>
rect 197 82 198 83 
<< m2 >>
rect 198 82 199 83 
<< m1 >>
rect 199 82 200 83 
<< m2 >>
rect 199 82 200 83 
<< m2 >>
rect 200 82 201 83 
<< m1 >>
rect 201 82 202 83 
<< m2 >>
rect 201 82 202 83 
<< m2c >>
rect 201 82 202 83 
<< m1 >>
rect 201 82 202 83 
<< m2 >>
rect 201 82 202 83 
<< m1 >>
rect 211 82 212 83 
<< m1 >>
rect 217 82 218 83 
<< m2 >>
rect 218 82 219 83 
<< m1 >>
rect 224 82 225 83 
<< m1 >>
rect 232 82 233 83 
<< m1 >>
rect 235 82 236 83 
<< m2 >>
rect 236 82 237 83 
<< m1 >>
rect 237 82 238 83 
<< m2 >>
rect 237 82 238 83 
<< m2c >>
rect 237 82 238 83 
<< m1 >>
rect 237 82 238 83 
<< m2 >>
rect 237 82 238 83 
<< m1 >>
rect 238 82 239 83 
<< m1 >>
rect 239 82 240 83 
<< m2 >>
rect 239 82 240 83 
<< m1 >>
rect 240 82 241 83 
<< m1 >>
rect 241 82 242 83 
<< m1 >>
rect 242 82 243 83 
<< m1 >>
rect 243 82 244 83 
<< m1 >>
rect 244 82 245 83 
<< m1 >>
rect 245 82 246 83 
<< m1 >>
rect 246 82 247 83 
<< m1 >>
rect 247 82 248 83 
<< m2 >>
rect 253 82 254 83 
<< m2 >>
rect 255 82 256 83 
<< m1 >>
rect 265 82 266 83 
<< m1 >>
rect 280 82 281 83 
<< m1 >>
rect 307 82 308 83 
<< m1 >>
rect 334 82 335 83 
<< m1 >>
rect 337 82 338 83 
<< m2 >>
rect 344 82 345 83 
<< m1 >>
rect 345 82 346 83 
<< m1 >>
rect 358 82 359 83 
<< m1 >>
rect 364 82 365 83 
<< m1 >>
rect 366 82 367 83 
<< m1 >>
rect 370 82 371 83 
<< m1 >>
rect 413 82 414 83 
<< m2 >>
rect 413 82 414 83 
<< m2c >>
rect 413 82 414 83 
<< m1 >>
rect 413 82 414 83 
<< m2 >>
rect 413 82 414 83 
<< m2 >>
rect 414 82 415 83 
<< m1 >>
rect 415 82 416 83 
<< m2 >>
rect 415 82 416 83 
<< m2 >>
rect 416 82 417 83 
<< m1 >>
rect 433 82 434 83 
<< m1 >>
rect 445 82 446 83 
<< m1 >>
rect 460 82 461 83 
<< m1 >>
rect 487 82 488 83 
<< m2 >>
rect 487 82 488 83 
<< m1 >>
rect 517 82 518 83 
<< m1 >>
rect 34 83 35 84 
<< m1 >>
rect 64 83 65 84 
<< m1 >>
rect 67 83 68 84 
<< m1 >>
rect 73 83 74 84 
<< m1 >>
rect 92 83 93 84 
<< m1 >>
rect 100 83 101 84 
<< m2 >>
rect 100 83 101 84 
<< m1 >>
rect 121 83 122 84 
<< m1 >>
rect 127 83 128 84 
<< m1 >>
rect 129 83 130 84 
<< m1 >>
rect 131 83 132 84 
<< m1 >>
rect 133 83 134 84 
<< m1 >>
rect 139 83 140 84 
<< m1 >>
rect 145 83 146 84 
<< m1 >>
rect 163 83 164 84 
<< m1 >>
rect 185 83 186 84 
<< m1 >>
rect 187 83 188 84 
<< m1 >>
rect 193 83 194 84 
<< m1 >>
rect 196 83 197 84 
<< m1 >>
rect 199 83 200 84 
<< m1 >>
rect 211 83 212 84 
<< m1 >>
rect 217 83 218 84 
<< m2 >>
rect 218 83 219 84 
<< m1 >>
rect 224 83 225 84 
<< m1 >>
rect 232 83 233 84 
<< m1 >>
rect 235 83 236 84 
<< m2 >>
rect 236 83 237 84 
<< m2 >>
rect 239 83 240 84 
<< m1 >>
rect 247 83 248 84 
<< m1 >>
rect 253 83 254 84 
<< m2 >>
rect 253 83 254 84 
<< m2c >>
rect 253 83 254 84 
<< m1 >>
rect 253 83 254 84 
<< m2 >>
rect 253 83 254 84 
<< m1 >>
rect 255 83 256 84 
<< m2 >>
rect 255 83 256 84 
<< m2c >>
rect 255 83 256 84 
<< m1 >>
rect 255 83 256 84 
<< m2 >>
rect 255 83 256 84 
<< m1 >>
rect 265 83 266 84 
<< m1 >>
rect 280 83 281 84 
<< m1 >>
rect 307 83 308 84 
<< m1 >>
rect 308 83 309 84 
<< m1 >>
rect 309 83 310 84 
<< m1 >>
rect 310 83 311 84 
<< m1 >>
rect 311 83 312 84 
<< m1 >>
rect 312 83 313 84 
<< m1 >>
rect 313 83 314 84 
<< m1 >>
rect 314 83 315 84 
<< m1 >>
rect 315 83 316 84 
<< m1 >>
rect 316 83 317 84 
<< m1 >>
rect 317 83 318 84 
<< m1 >>
rect 318 83 319 84 
<< m1 >>
rect 319 83 320 84 
<< m1 >>
rect 320 83 321 84 
<< m1 >>
rect 321 83 322 84 
<< m1 >>
rect 322 83 323 84 
<< m1 >>
rect 323 83 324 84 
<< m1 >>
rect 324 83 325 84 
<< m1 >>
rect 325 83 326 84 
<< m1 >>
rect 326 83 327 84 
<< m1 >>
rect 327 83 328 84 
<< m1 >>
rect 328 83 329 84 
<< m1 >>
rect 329 83 330 84 
<< m1 >>
rect 330 83 331 84 
<< m1 >>
rect 331 83 332 84 
<< m1 >>
rect 332 83 333 84 
<< m2 >>
rect 332 83 333 84 
<< m2c >>
rect 332 83 333 84 
<< m1 >>
rect 332 83 333 84 
<< m2 >>
rect 332 83 333 84 
<< m2 >>
rect 333 83 334 84 
<< m1 >>
rect 334 83 335 84 
<< m1 >>
rect 337 83 338 84 
<< m2 >>
rect 344 83 345 84 
<< m1 >>
rect 345 83 346 84 
<< m1 >>
rect 358 83 359 84 
<< m1 >>
rect 364 83 365 84 
<< m1 >>
rect 366 83 367 84 
<< m1 >>
rect 370 83 371 84 
<< m1 >>
rect 415 83 416 84 
<< m2 >>
rect 416 83 417 84 
<< m1 >>
rect 433 83 434 84 
<< m1 >>
rect 445 83 446 84 
<< m1 >>
rect 460 83 461 84 
<< m1 >>
rect 487 83 488 84 
<< m2 >>
rect 487 83 488 84 
<< m1 >>
rect 517 83 518 84 
<< pdiffusion >>
rect 12 84 13 85 
<< pdiffusion >>
rect 13 84 14 85 
<< pdiffusion >>
rect 14 84 15 85 
<< pdiffusion >>
rect 15 84 16 85 
<< pdiffusion >>
rect 16 84 17 85 
<< pdiffusion >>
rect 17 84 18 85 
<< pdiffusion >>
rect 30 84 31 85 
<< pdiffusion >>
rect 31 84 32 85 
<< pdiffusion >>
rect 32 84 33 85 
<< pdiffusion >>
rect 33 84 34 85 
<< m1 >>
rect 34 84 35 85 
<< pdiffusion >>
rect 34 84 35 85 
<< pdiffusion >>
rect 35 84 36 85 
<< pdiffusion >>
rect 48 84 49 85 
<< pdiffusion >>
rect 49 84 50 85 
<< pdiffusion >>
rect 50 84 51 85 
<< pdiffusion >>
rect 51 84 52 85 
<< pdiffusion >>
rect 52 84 53 85 
<< pdiffusion >>
rect 53 84 54 85 
<< m1 >>
rect 64 84 65 85 
<< pdiffusion >>
rect 66 84 67 85 
<< m1 >>
rect 67 84 68 85 
<< pdiffusion >>
rect 67 84 68 85 
<< pdiffusion >>
rect 68 84 69 85 
<< pdiffusion >>
rect 69 84 70 85 
<< pdiffusion >>
rect 70 84 71 85 
<< pdiffusion >>
rect 71 84 72 85 
<< m1 >>
rect 73 84 74 85 
<< pdiffusion >>
rect 84 84 85 85 
<< pdiffusion >>
rect 85 84 86 85 
<< pdiffusion >>
rect 86 84 87 85 
<< pdiffusion >>
rect 87 84 88 85 
<< pdiffusion >>
rect 88 84 89 85 
<< pdiffusion >>
rect 89 84 90 85 
<< m1 >>
rect 92 84 93 85 
<< m1 >>
rect 100 84 101 85 
<< m2 >>
rect 100 84 101 85 
<< pdiffusion >>
rect 102 84 103 85 
<< pdiffusion >>
rect 103 84 104 85 
<< pdiffusion >>
rect 104 84 105 85 
<< pdiffusion >>
rect 105 84 106 85 
<< pdiffusion >>
rect 106 84 107 85 
<< pdiffusion >>
rect 107 84 108 85 
<< pdiffusion >>
rect 120 84 121 85 
<< m1 >>
rect 121 84 122 85 
<< pdiffusion >>
rect 121 84 122 85 
<< pdiffusion >>
rect 122 84 123 85 
<< pdiffusion >>
rect 123 84 124 85 
<< pdiffusion >>
rect 124 84 125 85 
<< pdiffusion >>
rect 125 84 126 85 
<< m1 >>
rect 127 84 128 85 
<< m1 >>
rect 129 84 130 85 
<< m1 >>
rect 131 84 132 85 
<< m1 >>
rect 133 84 134 85 
<< pdiffusion >>
rect 138 84 139 85 
<< m1 >>
rect 139 84 140 85 
<< pdiffusion >>
rect 139 84 140 85 
<< pdiffusion >>
rect 140 84 141 85 
<< pdiffusion >>
rect 141 84 142 85 
<< pdiffusion >>
rect 142 84 143 85 
<< pdiffusion >>
rect 143 84 144 85 
<< m1 >>
rect 145 84 146 85 
<< pdiffusion >>
rect 156 84 157 85 
<< pdiffusion >>
rect 157 84 158 85 
<< pdiffusion >>
rect 158 84 159 85 
<< pdiffusion >>
rect 159 84 160 85 
<< pdiffusion >>
rect 160 84 161 85 
<< pdiffusion >>
rect 161 84 162 85 
<< m1 >>
rect 163 84 164 85 
<< pdiffusion >>
rect 174 84 175 85 
<< pdiffusion >>
rect 175 84 176 85 
<< pdiffusion >>
rect 176 84 177 85 
<< pdiffusion >>
rect 177 84 178 85 
<< pdiffusion >>
rect 178 84 179 85 
<< pdiffusion >>
rect 179 84 180 85 
<< m1 >>
rect 185 84 186 85 
<< m1 >>
rect 187 84 188 85 
<< pdiffusion >>
rect 192 84 193 85 
<< m1 >>
rect 193 84 194 85 
<< pdiffusion >>
rect 193 84 194 85 
<< pdiffusion >>
rect 194 84 195 85 
<< pdiffusion >>
rect 195 84 196 85 
<< m1 >>
rect 196 84 197 85 
<< pdiffusion >>
rect 196 84 197 85 
<< pdiffusion >>
rect 197 84 198 85 
<< m1 >>
rect 199 84 200 85 
<< pdiffusion >>
rect 210 84 211 85 
<< m1 >>
rect 211 84 212 85 
<< pdiffusion >>
rect 211 84 212 85 
<< pdiffusion >>
rect 212 84 213 85 
<< pdiffusion >>
rect 213 84 214 85 
<< pdiffusion >>
rect 214 84 215 85 
<< pdiffusion >>
rect 215 84 216 85 
<< m1 >>
rect 217 84 218 85 
<< m2 >>
rect 218 84 219 85 
<< m1 >>
rect 224 84 225 85 
<< pdiffusion >>
rect 228 84 229 85 
<< pdiffusion >>
rect 229 84 230 85 
<< pdiffusion >>
rect 230 84 231 85 
<< pdiffusion >>
rect 231 84 232 85 
<< m1 >>
rect 232 84 233 85 
<< pdiffusion >>
rect 232 84 233 85 
<< pdiffusion >>
rect 233 84 234 85 
<< m1 >>
rect 235 84 236 85 
<< m2 >>
rect 236 84 237 85 
<< m1 >>
rect 239 84 240 85 
<< m2 >>
rect 239 84 240 85 
<< m2c >>
rect 239 84 240 85 
<< m1 >>
rect 239 84 240 85 
<< m2 >>
rect 239 84 240 85 
<< m1 >>
rect 240 84 241 85 
<< m1 >>
rect 241 84 242 85 
<< pdiffusion >>
rect 246 84 247 85 
<< m1 >>
rect 247 84 248 85 
<< pdiffusion >>
rect 247 84 248 85 
<< pdiffusion >>
rect 248 84 249 85 
<< pdiffusion >>
rect 249 84 250 85 
<< pdiffusion >>
rect 250 84 251 85 
<< pdiffusion >>
rect 251 84 252 85 
<< m1 >>
rect 253 84 254 85 
<< m1 >>
rect 255 84 256 85 
<< pdiffusion >>
rect 264 84 265 85 
<< m1 >>
rect 265 84 266 85 
<< pdiffusion >>
rect 265 84 266 85 
<< pdiffusion >>
rect 266 84 267 85 
<< pdiffusion >>
rect 267 84 268 85 
<< pdiffusion >>
rect 268 84 269 85 
<< pdiffusion >>
rect 269 84 270 85 
<< m1 >>
rect 280 84 281 85 
<< pdiffusion >>
rect 282 84 283 85 
<< pdiffusion >>
rect 283 84 284 85 
<< pdiffusion >>
rect 284 84 285 85 
<< pdiffusion >>
rect 285 84 286 85 
<< pdiffusion >>
rect 286 84 287 85 
<< pdiffusion >>
rect 287 84 288 85 
<< pdiffusion >>
rect 300 84 301 85 
<< pdiffusion >>
rect 301 84 302 85 
<< pdiffusion >>
rect 302 84 303 85 
<< pdiffusion >>
rect 303 84 304 85 
<< pdiffusion >>
rect 304 84 305 85 
<< pdiffusion >>
rect 305 84 306 85 
<< m2 >>
rect 333 84 334 85 
<< m1 >>
rect 334 84 335 85 
<< pdiffusion >>
rect 336 84 337 85 
<< m1 >>
rect 337 84 338 85 
<< pdiffusion >>
rect 337 84 338 85 
<< pdiffusion >>
rect 338 84 339 85 
<< pdiffusion >>
rect 339 84 340 85 
<< pdiffusion >>
rect 340 84 341 85 
<< pdiffusion >>
rect 341 84 342 85 
<< m2 >>
rect 344 84 345 85 
<< m1 >>
rect 345 84 346 85 
<< pdiffusion >>
rect 354 84 355 85 
<< pdiffusion >>
rect 355 84 356 85 
<< pdiffusion >>
rect 356 84 357 85 
<< pdiffusion >>
rect 357 84 358 85 
<< m1 >>
rect 358 84 359 85 
<< pdiffusion >>
rect 358 84 359 85 
<< pdiffusion >>
rect 359 84 360 85 
<< m1 >>
rect 364 84 365 85 
<< m1 >>
rect 366 84 367 85 
<< m1 >>
rect 370 84 371 85 
<< pdiffusion >>
rect 372 84 373 85 
<< pdiffusion >>
rect 373 84 374 85 
<< pdiffusion >>
rect 374 84 375 85 
<< pdiffusion >>
rect 375 84 376 85 
<< pdiffusion >>
rect 376 84 377 85 
<< pdiffusion >>
rect 377 84 378 85 
<< pdiffusion >>
rect 390 84 391 85 
<< pdiffusion >>
rect 391 84 392 85 
<< pdiffusion >>
rect 392 84 393 85 
<< pdiffusion >>
rect 393 84 394 85 
<< pdiffusion >>
rect 394 84 395 85 
<< pdiffusion >>
rect 395 84 396 85 
<< pdiffusion >>
rect 408 84 409 85 
<< pdiffusion >>
rect 409 84 410 85 
<< pdiffusion >>
rect 410 84 411 85 
<< pdiffusion >>
rect 411 84 412 85 
<< pdiffusion >>
rect 412 84 413 85 
<< pdiffusion >>
rect 413 84 414 85 
<< m1 >>
rect 415 84 416 85 
<< m2 >>
rect 416 84 417 85 
<< pdiffusion >>
rect 426 84 427 85 
<< pdiffusion >>
rect 427 84 428 85 
<< pdiffusion >>
rect 428 84 429 85 
<< pdiffusion >>
rect 429 84 430 85 
<< pdiffusion >>
rect 430 84 431 85 
<< pdiffusion >>
rect 431 84 432 85 
<< m1 >>
rect 433 84 434 85 
<< pdiffusion >>
rect 444 84 445 85 
<< m1 >>
rect 445 84 446 85 
<< pdiffusion >>
rect 445 84 446 85 
<< pdiffusion >>
rect 446 84 447 85 
<< pdiffusion >>
rect 447 84 448 85 
<< pdiffusion >>
rect 448 84 449 85 
<< pdiffusion >>
rect 449 84 450 85 
<< m1 >>
rect 460 84 461 85 
<< pdiffusion >>
rect 462 84 463 85 
<< pdiffusion >>
rect 463 84 464 85 
<< pdiffusion >>
rect 464 84 465 85 
<< pdiffusion >>
rect 465 84 466 85 
<< pdiffusion >>
rect 466 84 467 85 
<< pdiffusion >>
rect 467 84 468 85 
<< pdiffusion >>
rect 480 84 481 85 
<< pdiffusion >>
rect 481 84 482 85 
<< pdiffusion >>
rect 482 84 483 85 
<< pdiffusion >>
rect 483 84 484 85 
<< pdiffusion >>
rect 484 84 485 85 
<< pdiffusion >>
rect 485 84 486 85 
<< m1 >>
rect 487 84 488 85 
<< m2 >>
rect 487 84 488 85 
<< pdiffusion >>
rect 516 84 517 85 
<< m1 >>
rect 517 84 518 85 
<< pdiffusion >>
rect 517 84 518 85 
<< pdiffusion >>
rect 518 84 519 85 
<< pdiffusion >>
rect 519 84 520 85 
<< pdiffusion >>
rect 520 84 521 85 
<< pdiffusion >>
rect 521 84 522 85 
<< pdiffusion >>
rect 12 85 13 86 
<< pdiffusion >>
rect 13 85 14 86 
<< pdiffusion >>
rect 14 85 15 86 
<< pdiffusion >>
rect 15 85 16 86 
<< pdiffusion >>
rect 16 85 17 86 
<< pdiffusion >>
rect 17 85 18 86 
<< pdiffusion >>
rect 30 85 31 86 
<< pdiffusion >>
rect 31 85 32 86 
<< pdiffusion >>
rect 32 85 33 86 
<< pdiffusion >>
rect 33 85 34 86 
<< pdiffusion >>
rect 34 85 35 86 
<< pdiffusion >>
rect 35 85 36 86 
<< pdiffusion >>
rect 48 85 49 86 
<< pdiffusion >>
rect 49 85 50 86 
<< pdiffusion >>
rect 50 85 51 86 
<< pdiffusion >>
rect 51 85 52 86 
<< pdiffusion >>
rect 52 85 53 86 
<< pdiffusion >>
rect 53 85 54 86 
<< m1 >>
rect 64 85 65 86 
<< pdiffusion >>
rect 66 85 67 86 
<< pdiffusion >>
rect 67 85 68 86 
<< pdiffusion >>
rect 68 85 69 86 
<< pdiffusion >>
rect 69 85 70 86 
<< pdiffusion >>
rect 70 85 71 86 
<< pdiffusion >>
rect 71 85 72 86 
<< m1 >>
rect 73 85 74 86 
<< pdiffusion >>
rect 84 85 85 86 
<< pdiffusion >>
rect 85 85 86 86 
<< pdiffusion >>
rect 86 85 87 86 
<< pdiffusion >>
rect 87 85 88 86 
<< pdiffusion >>
rect 88 85 89 86 
<< pdiffusion >>
rect 89 85 90 86 
<< m1 >>
rect 92 85 93 86 
<< m1 >>
rect 100 85 101 86 
<< m2 >>
rect 100 85 101 86 
<< pdiffusion >>
rect 102 85 103 86 
<< pdiffusion >>
rect 103 85 104 86 
<< pdiffusion >>
rect 104 85 105 86 
<< pdiffusion >>
rect 105 85 106 86 
<< pdiffusion >>
rect 106 85 107 86 
<< pdiffusion >>
rect 107 85 108 86 
<< pdiffusion >>
rect 120 85 121 86 
<< pdiffusion >>
rect 121 85 122 86 
<< pdiffusion >>
rect 122 85 123 86 
<< pdiffusion >>
rect 123 85 124 86 
<< pdiffusion >>
rect 124 85 125 86 
<< pdiffusion >>
rect 125 85 126 86 
<< m1 >>
rect 127 85 128 86 
<< m1 >>
rect 129 85 130 86 
<< m1 >>
rect 131 85 132 86 
<< m1 >>
rect 133 85 134 86 
<< pdiffusion >>
rect 138 85 139 86 
<< pdiffusion >>
rect 139 85 140 86 
<< pdiffusion >>
rect 140 85 141 86 
<< pdiffusion >>
rect 141 85 142 86 
<< pdiffusion >>
rect 142 85 143 86 
<< pdiffusion >>
rect 143 85 144 86 
<< m1 >>
rect 145 85 146 86 
<< pdiffusion >>
rect 156 85 157 86 
<< pdiffusion >>
rect 157 85 158 86 
<< pdiffusion >>
rect 158 85 159 86 
<< pdiffusion >>
rect 159 85 160 86 
<< pdiffusion >>
rect 160 85 161 86 
<< pdiffusion >>
rect 161 85 162 86 
<< m1 >>
rect 163 85 164 86 
<< pdiffusion >>
rect 174 85 175 86 
<< pdiffusion >>
rect 175 85 176 86 
<< pdiffusion >>
rect 176 85 177 86 
<< pdiffusion >>
rect 177 85 178 86 
<< pdiffusion >>
rect 178 85 179 86 
<< pdiffusion >>
rect 179 85 180 86 
<< m1 >>
rect 185 85 186 86 
<< m1 >>
rect 187 85 188 86 
<< pdiffusion >>
rect 192 85 193 86 
<< pdiffusion >>
rect 193 85 194 86 
<< pdiffusion >>
rect 194 85 195 86 
<< pdiffusion >>
rect 195 85 196 86 
<< pdiffusion >>
rect 196 85 197 86 
<< pdiffusion >>
rect 197 85 198 86 
<< m1 >>
rect 199 85 200 86 
<< pdiffusion >>
rect 210 85 211 86 
<< pdiffusion >>
rect 211 85 212 86 
<< pdiffusion >>
rect 212 85 213 86 
<< pdiffusion >>
rect 213 85 214 86 
<< pdiffusion >>
rect 214 85 215 86 
<< pdiffusion >>
rect 215 85 216 86 
<< m1 >>
rect 217 85 218 86 
<< m2 >>
rect 218 85 219 86 
<< m1 >>
rect 224 85 225 86 
<< pdiffusion >>
rect 228 85 229 86 
<< pdiffusion >>
rect 229 85 230 86 
<< pdiffusion >>
rect 230 85 231 86 
<< pdiffusion >>
rect 231 85 232 86 
<< pdiffusion >>
rect 232 85 233 86 
<< pdiffusion >>
rect 233 85 234 86 
<< m1 >>
rect 235 85 236 86 
<< m2 >>
rect 236 85 237 86 
<< m1 >>
rect 241 85 242 86 
<< pdiffusion >>
rect 246 85 247 86 
<< pdiffusion >>
rect 247 85 248 86 
<< pdiffusion >>
rect 248 85 249 86 
<< pdiffusion >>
rect 249 85 250 86 
<< pdiffusion >>
rect 250 85 251 86 
<< pdiffusion >>
rect 251 85 252 86 
<< m1 >>
rect 253 85 254 86 
<< m1 >>
rect 255 85 256 86 
<< pdiffusion >>
rect 264 85 265 86 
<< pdiffusion >>
rect 265 85 266 86 
<< pdiffusion >>
rect 266 85 267 86 
<< pdiffusion >>
rect 267 85 268 86 
<< pdiffusion >>
rect 268 85 269 86 
<< pdiffusion >>
rect 269 85 270 86 
<< m1 >>
rect 280 85 281 86 
<< pdiffusion >>
rect 282 85 283 86 
<< pdiffusion >>
rect 283 85 284 86 
<< pdiffusion >>
rect 284 85 285 86 
<< pdiffusion >>
rect 285 85 286 86 
<< pdiffusion >>
rect 286 85 287 86 
<< pdiffusion >>
rect 287 85 288 86 
<< pdiffusion >>
rect 300 85 301 86 
<< pdiffusion >>
rect 301 85 302 86 
<< pdiffusion >>
rect 302 85 303 86 
<< pdiffusion >>
rect 303 85 304 86 
<< pdiffusion >>
rect 304 85 305 86 
<< pdiffusion >>
rect 305 85 306 86 
<< m2 >>
rect 333 85 334 86 
<< m1 >>
rect 334 85 335 86 
<< pdiffusion >>
rect 336 85 337 86 
<< pdiffusion >>
rect 337 85 338 86 
<< pdiffusion >>
rect 338 85 339 86 
<< pdiffusion >>
rect 339 85 340 86 
<< pdiffusion >>
rect 340 85 341 86 
<< pdiffusion >>
rect 341 85 342 86 
<< m2 >>
rect 344 85 345 86 
<< m1 >>
rect 345 85 346 86 
<< pdiffusion >>
rect 354 85 355 86 
<< pdiffusion >>
rect 355 85 356 86 
<< pdiffusion >>
rect 356 85 357 86 
<< pdiffusion >>
rect 357 85 358 86 
<< pdiffusion >>
rect 358 85 359 86 
<< pdiffusion >>
rect 359 85 360 86 
<< m1 >>
rect 364 85 365 86 
<< m1 >>
rect 366 85 367 86 
<< m1 >>
rect 370 85 371 86 
<< pdiffusion >>
rect 372 85 373 86 
<< pdiffusion >>
rect 373 85 374 86 
<< pdiffusion >>
rect 374 85 375 86 
<< pdiffusion >>
rect 375 85 376 86 
<< pdiffusion >>
rect 376 85 377 86 
<< pdiffusion >>
rect 377 85 378 86 
<< pdiffusion >>
rect 390 85 391 86 
<< pdiffusion >>
rect 391 85 392 86 
<< pdiffusion >>
rect 392 85 393 86 
<< pdiffusion >>
rect 393 85 394 86 
<< pdiffusion >>
rect 394 85 395 86 
<< pdiffusion >>
rect 395 85 396 86 
<< pdiffusion >>
rect 408 85 409 86 
<< pdiffusion >>
rect 409 85 410 86 
<< pdiffusion >>
rect 410 85 411 86 
<< pdiffusion >>
rect 411 85 412 86 
<< pdiffusion >>
rect 412 85 413 86 
<< pdiffusion >>
rect 413 85 414 86 
<< m1 >>
rect 415 85 416 86 
<< m2 >>
rect 416 85 417 86 
<< pdiffusion >>
rect 426 85 427 86 
<< pdiffusion >>
rect 427 85 428 86 
<< pdiffusion >>
rect 428 85 429 86 
<< pdiffusion >>
rect 429 85 430 86 
<< pdiffusion >>
rect 430 85 431 86 
<< pdiffusion >>
rect 431 85 432 86 
<< m1 >>
rect 433 85 434 86 
<< pdiffusion >>
rect 444 85 445 86 
<< pdiffusion >>
rect 445 85 446 86 
<< pdiffusion >>
rect 446 85 447 86 
<< pdiffusion >>
rect 447 85 448 86 
<< pdiffusion >>
rect 448 85 449 86 
<< pdiffusion >>
rect 449 85 450 86 
<< m1 >>
rect 460 85 461 86 
<< pdiffusion >>
rect 462 85 463 86 
<< pdiffusion >>
rect 463 85 464 86 
<< pdiffusion >>
rect 464 85 465 86 
<< pdiffusion >>
rect 465 85 466 86 
<< pdiffusion >>
rect 466 85 467 86 
<< pdiffusion >>
rect 467 85 468 86 
<< pdiffusion >>
rect 480 85 481 86 
<< pdiffusion >>
rect 481 85 482 86 
<< pdiffusion >>
rect 482 85 483 86 
<< pdiffusion >>
rect 483 85 484 86 
<< pdiffusion >>
rect 484 85 485 86 
<< pdiffusion >>
rect 485 85 486 86 
<< m1 >>
rect 487 85 488 86 
<< m2 >>
rect 487 85 488 86 
<< pdiffusion >>
rect 516 85 517 86 
<< pdiffusion >>
rect 517 85 518 86 
<< pdiffusion >>
rect 518 85 519 86 
<< pdiffusion >>
rect 519 85 520 86 
<< pdiffusion >>
rect 520 85 521 86 
<< pdiffusion >>
rect 521 85 522 86 
<< pdiffusion >>
rect 12 86 13 87 
<< pdiffusion >>
rect 13 86 14 87 
<< pdiffusion >>
rect 14 86 15 87 
<< pdiffusion >>
rect 15 86 16 87 
<< pdiffusion >>
rect 16 86 17 87 
<< pdiffusion >>
rect 17 86 18 87 
<< pdiffusion >>
rect 30 86 31 87 
<< pdiffusion >>
rect 31 86 32 87 
<< pdiffusion >>
rect 32 86 33 87 
<< pdiffusion >>
rect 33 86 34 87 
<< pdiffusion >>
rect 34 86 35 87 
<< pdiffusion >>
rect 35 86 36 87 
<< pdiffusion >>
rect 48 86 49 87 
<< pdiffusion >>
rect 49 86 50 87 
<< pdiffusion >>
rect 50 86 51 87 
<< pdiffusion >>
rect 51 86 52 87 
<< pdiffusion >>
rect 52 86 53 87 
<< pdiffusion >>
rect 53 86 54 87 
<< m1 >>
rect 64 86 65 87 
<< pdiffusion >>
rect 66 86 67 87 
<< pdiffusion >>
rect 67 86 68 87 
<< pdiffusion >>
rect 68 86 69 87 
<< pdiffusion >>
rect 69 86 70 87 
<< pdiffusion >>
rect 70 86 71 87 
<< pdiffusion >>
rect 71 86 72 87 
<< m1 >>
rect 73 86 74 87 
<< pdiffusion >>
rect 84 86 85 87 
<< pdiffusion >>
rect 85 86 86 87 
<< pdiffusion >>
rect 86 86 87 87 
<< pdiffusion >>
rect 87 86 88 87 
<< pdiffusion >>
rect 88 86 89 87 
<< pdiffusion >>
rect 89 86 90 87 
<< m1 >>
rect 92 86 93 87 
<< m1 >>
rect 100 86 101 87 
<< m2 >>
rect 100 86 101 87 
<< pdiffusion >>
rect 102 86 103 87 
<< pdiffusion >>
rect 103 86 104 87 
<< pdiffusion >>
rect 104 86 105 87 
<< pdiffusion >>
rect 105 86 106 87 
<< pdiffusion >>
rect 106 86 107 87 
<< pdiffusion >>
rect 107 86 108 87 
<< pdiffusion >>
rect 120 86 121 87 
<< pdiffusion >>
rect 121 86 122 87 
<< pdiffusion >>
rect 122 86 123 87 
<< pdiffusion >>
rect 123 86 124 87 
<< pdiffusion >>
rect 124 86 125 87 
<< pdiffusion >>
rect 125 86 126 87 
<< m1 >>
rect 127 86 128 87 
<< m1 >>
rect 129 86 130 87 
<< m1 >>
rect 131 86 132 87 
<< m1 >>
rect 133 86 134 87 
<< pdiffusion >>
rect 138 86 139 87 
<< pdiffusion >>
rect 139 86 140 87 
<< pdiffusion >>
rect 140 86 141 87 
<< pdiffusion >>
rect 141 86 142 87 
<< pdiffusion >>
rect 142 86 143 87 
<< pdiffusion >>
rect 143 86 144 87 
<< m1 >>
rect 145 86 146 87 
<< pdiffusion >>
rect 156 86 157 87 
<< pdiffusion >>
rect 157 86 158 87 
<< pdiffusion >>
rect 158 86 159 87 
<< pdiffusion >>
rect 159 86 160 87 
<< pdiffusion >>
rect 160 86 161 87 
<< pdiffusion >>
rect 161 86 162 87 
<< m1 >>
rect 163 86 164 87 
<< pdiffusion >>
rect 174 86 175 87 
<< pdiffusion >>
rect 175 86 176 87 
<< pdiffusion >>
rect 176 86 177 87 
<< pdiffusion >>
rect 177 86 178 87 
<< pdiffusion >>
rect 178 86 179 87 
<< pdiffusion >>
rect 179 86 180 87 
<< m1 >>
rect 185 86 186 87 
<< m1 >>
rect 187 86 188 87 
<< pdiffusion >>
rect 192 86 193 87 
<< pdiffusion >>
rect 193 86 194 87 
<< pdiffusion >>
rect 194 86 195 87 
<< pdiffusion >>
rect 195 86 196 87 
<< pdiffusion >>
rect 196 86 197 87 
<< pdiffusion >>
rect 197 86 198 87 
<< m1 >>
rect 199 86 200 87 
<< pdiffusion >>
rect 210 86 211 87 
<< pdiffusion >>
rect 211 86 212 87 
<< pdiffusion >>
rect 212 86 213 87 
<< pdiffusion >>
rect 213 86 214 87 
<< pdiffusion >>
rect 214 86 215 87 
<< pdiffusion >>
rect 215 86 216 87 
<< m1 >>
rect 217 86 218 87 
<< m2 >>
rect 218 86 219 87 
<< m1 >>
rect 224 86 225 87 
<< pdiffusion >>
rect 228 86 229 87 
<< pdiffusion >>
rect 229 86 230 87 
<< pdiffusion >>
rect 230 86 231 87 
<< pdiffusion >>
rect 231 86 232 87 
<< pdiffusion >>
rect 232 86 233 87 
<< pdiffusion >>
rect 233 86 234 87 
<< m1 >>
rect 235 86 236 87 
<< m2 >>
rect 236 86 237 87 
<< m1 >>
rect 241 86 242 87 
<< pdiffusion >>
rect 246 86 247 87 
<< pdiffusion >>
rect 247 86 248 87 
<< pdiffusion >>
rect 248 86 249 87 
<< pdiffusion >>
rect 249 86 250 87 
<< pdiffusion >>
rect 250 86 251 87 
<< pdiffusion >>
rect 251 86 252 87 
<< m1 >>
rect 253 86 254 87 
<< m1 >>
rect 255 86 256 87 
<< pdiffusion >>
rect 264 86 265 87 
<< pdiffusion >>
rect 265 86 266 87 
<< pdiffusion >>
rect 266 86 267 87 
<< pdiffusion >>
rect 267 86 268 87 
<< pdiffusion >>
rect 268 86 269 87 
<< pdiffusion >>
rect 269 86 270 87 
<< m1 >>
rect 280 86 281 87 
<< pdiffusion >>
rect 282 86 283 87 
<< pdiffusion >>
rect 283 86 284 87 
<< pdiffusion >>
rect 284 86 285 87 
<< pdiffusion >>
rect 285 86 286 87 
<< pdiffusion >>
rect 286 86 287 87 
<< pdiffusion >>
rect 287 86 288 87 
<< pdiffusion >>
rect 300 86 301 87 
<< pdiffusion >>
rect 301 86 302 87 
<< pdiffusion >>
rect 302 86 303 87 
<< pdiffusion >>
rect 303 86 304 87 
<< pdiffusion >>
rect 304 86 305 87 
<< pdiffusion >>
rect 305 86 306 87 
<< m2 >>
rect 333 86 334 87 
<< m1 >>
rect 334 86 335 87 
<< pdiffusion >>
rect 336 86 337 87 
<< pdiffusion >>
rect 337 86 338 87 
<< pdiffusion >>
rect 338 86 339 87 
<< pdiffusion >>
rect 339 86 340 87 
<< pdiffusion >>
rect 340 86 341 87 
<< pdiffusion >>
rect 341 86 342 87 
<< m2 >>
rect 344 86 345 87 
<< m1 >>
rect 345 86 346 87 
<< pdiffusion >>
rect 354 86 355 87 
<< pdiffusion >>
rect 355 86 356 87 
<< pdiffusion >>
rect 356 86 357 87 
<< pdiffusion >>
rect 357 86 358 87 
<< pdiffusion >>
rect 358 86 359 87 
<< pdiffusion >>
rect 359 86 360 87 
<< m1 >>
rect 364 86 365 87 
<< m1 >>
rect 366 86 367 87 
<< m1 >>
rect 370 86 371 87 
<< pdiffusion >>
rect 372 86 373 87 
<< pdiffusion >>
rect 373 86 374 87 
<< pdiffusion >>
rect 374 86 375 87 
<< pdiffusion >>
rect 375 86 376 87 
<< pdiffusion >>
rect 376 86 377 87 
<< pdiffusion >>
rect 377 86 378 87 
<< pdiffusion >>
rect 390 86 391 87 
<< pdiffusion >>
rect 391 86 392 87 
<< pdiffusion >>
rect 392 86 393 87 
<< pdiffusion >>
rect 393 86 394 87 
<< pdiffusion >>
rect 394 86 395 87 
<< pdiffusion >>
rect 395 86 396 87 
<< pdiffusion >>
rect 408 86 409 87 
<< pdiffusion >>
rect 409 86 410 87 
<< pdiffusion >>
rect 410 86 411 87 
<< pdiffusion >>
rect 411 86 412 87 
<< pdiffusion >>
rect 412 86 413 87 
<< pdiffusion >>
rect 413 86 414 87 
<< m1 >>
rect 415 86 416 87 
<< m2 >>
rect 416 86 417 87 
<< pdiffusion >>
rect 426 86 427 87 
<< pdiffusion >>
rect 427 86 428 87 
<< pdiffusion >>
rect 428 86 429 87 
<< pdiffusion >>
rect 429 86 430 87 
<< pdiffusion >>
rect 430 86 431 87 
<< pdiffusion >>
rect 431 86 432 87 
<< m1 >>
rect 433 86 434 87 
<< pdiffusion >>
rect 444 86 445 87 
<< pdiffusion >>
rect 445 86 446 87 
<< pdiffusion >>
rect 446 86 447 87 
<< pdiffusion >>
rect 447 86 448 87 
<< pdiffusion >>
rect 448 86 449 87 
<< pdiffusion >>
rect 449 86 450 87 
<< m1 >>
rect 460 86 461 87 
<< pdiffusion >>
rect 462 86 463 87 
<< pdiffusion >>
rect 463 86 464 87 
<< pdiffusion >>
rect 464 86 465 87 
<< pdiffusion >>
rect 465 86 466 87 
<< pdiffusion >>
rect 466 86 467 87 
<< pdiffusion >>
rect 467 86 468 87 
<< pdiffusion >>
rect 480 86 481 87 
<< pdiffusion >>
rect 481 86 482 87 
<< pdiffusion >>
rect 482 86 483 87 
<< pdiffusion >>
rect 483 86 484 87 
<< pdiffusion >>
rect 484 86 485 87 
<< pdiffusion >>
rect 485 86 486 87 
<< m1 >>
rect 487 86 488 87 
<< m2 >>
rect 487 86 488 87 
<< pdiffusion >>
rect 516 86 517 87 
<< pdiffusion >>
rect 517 86 518 87 
<< pdiffusion >>
rect 518 86 519 87 
<< pdiffusion >>
rect 519 86 520 87 
<< pdiffusion >>
rect 520 86 521 87 
<< pdiffusion >>
rect 521 86 522 87 
<< pdiffusion >>
rect 12 87 13 88 
<< pdiffusion >>
rect 13 87 14 88 
<< pdiffusion >>
rect 14 87 15 88 
<< pdiffusion >>
rect 15 87 16 88 
<< pdiffusion >>
rect 16 87 17 88 
<< pdiffusion >>
rect 17 87 18 88 
<< pdiffusion >>
rect 30 87 31 88 
<< pdiffusion >>
rect 31 87 32 88 
<< pdiffusion >>
rect 32 87 33 88 
<< pdiffusion >>
rect 33 87 34 88 
<< pdiffusion >>
rect 34 87 35 88 
<< pdiffusion >>
rect 35 87 36 88 
<< pdiffusion >>
rect 48 87 49 88 
<< pdiffusion >>
rect 49 87 50 88 
<< pdiffusion >>
rect 50 87 51 88 
<< pdiffusion >>
rect 51 87 52 88 
<< pdiffusion >>
rect 52 87 53 88 
<< pdiffusion >>
rect 53 87 54 88 
<< m1 >>
rect 64 87 65 88 
<< pdiffusion >>
rect 66 87 67 88 
<< pdiffusion >>
rect 67 87 68 88 
<< pdiffusion >>
rect 68 87 69 88 
<< pdiffusion >>
rect 69 87 70 88 
<< pdiffusion >>
rect 70 87 71 88 
<< pdiffusion >>
rect 71 87 72 88 
<< m1 >>
rect 73 87 74 88 
<< pdiffusion >>
rect 84 87 85 88 
<< pdiffusion >>
rect 85 87 86 88 
<< pdiffusion >>
rect 86 87 87 88 
<< pdiffusion >>
rect 87 87 88 88 
<< pdiffusion >>
rect 88 87 89 88 
<< pdiffusion >>
rect 89 87 90 88 
<< m1 >>
rect 92 87 93 88 
<< m1 >>
rect 100 87 101 88 
<< m2 >>
rect 100 87 101 88 
<< pdiffusion >>
rect 102 87 103 88 
<< pdiffusion >>
rect 103 87 104 88 
<< pdiffusion >>
rect 104 87 105 88 
<< pdiffusion >>
rect 105 87 106 88 
<< pdiffusion >>
rect 106 87 107 88 
<< pdiffusion >>
rect 107 87 108 88 
<< pdiffusion >>
rect 120 87 121 88 
<< pdiffusion >>
rect 121 87 122 88 
<< pdiffusion >>
rect 122 87 123 88 
<< pdiffusion >>
rect 123 87 124 88 
<< pdiffusion >>
rect 124 87 125 88 
<< pdiffusion >>
rect 125 87 126 88 
<< m1 >>
rect 127 87 128 88 
<< m1 >>
rect 129 87 130 88 
<< m1 >>
rect 131 87 132 88 
<< m1 >>
rect 133 87 134 88 
<< pdiffusion >>
rect 138 87 139 88 
<< pdiffusion >>
rect 139 87 140 88 
<< pdiffusion >>
rect 140 87 141 88 
<< pdiffusion >>
rect 141 87 142 88 
<< pdiffusion >>
rect 142 87 143 88 
<< pdiffusion >>
rect 143 87 144 88 
<< m1 >>
rect 145 87 146 88 
<< pdiffusion >>
rect 156 87 157 88 
<< pdiffusion >>
rect 157 87 158 88 
<< pdiffusion >>
rect 158 87 159 88 
<< pdiffusion >>
rect 159 87 160 88 
<< pdiffusion >>
rect 160 87 161 88 
<< pdiffusion >>
rect 161 87 162 88 
<< m1 >>
rect 163 87 164 88 
<< pdiffusion >>
rect 174 87 175 88 
<< pdiffusion >>
rect 175 87 176 88 
<< pdiffusion >>
rect 176 87 177 88 
<< pdiffusion >>
rect 177 87 178 88 
<< pdiffusion >>
rect 178 87 179 88 
<< pdiffusion >>
rect 179 87 180 88 
<< m1 >>
rect 185 87 186 88 
<< m1 >>
rect 187 87 188 88 
<< pdiffusion >>
rect 192 87 193 88 
<< pdiffusion >>
rect 193 87 194 88 
<< pdiffusion >>
rect 194 87 195 88 
<< pdiffusion >>
rect 195 87 196 88 
<< pdiffusion >>
rect 196 87 197 88 
<< pdiffusion >>
rect 197 87 198 88 
<< m1 >>
rect 199 87 200 88 
<< pdiffusion >>
rect 210 87 211 88 
<< pdiffusion >>
rect 211 87 212 88 
<< pdiffusion >>
rect 212 87 213 88 
<< pdiffusion >>
rect 213 87 214 88 
<< pdiffusion >>
rect 214 87 215 88 
<< pdiffusion >>
rect 215 87 216 88 
<< m1 >>
rect 217 87 218 88 
<< m2 >>
rect 218 87 219 88 
<< m1 >>
rect 224 87 225 88 
<< pdiffusion >>
rect 228 87 229 88 
<< pdiffusion >>
rect 229 87 230 88 
<< pdiffusion >>
rect 230 87 231 88 
<< pdiffusion >>
rect 231 87 232 88 
<< pdiffusion >>
rect 232 87 233 88 
<< pdiffusion >>
rect 233 87 234 88 
<< m1 >>
rect 235 87 236 88 
<< m2 >>
rect 236 87 237 88 
<< m1 >>
rect 241 87 242 88 
<< pdiffusion >>
rect 246 87 247 88 
<< pdiffusion >>
rect 247 87 248 88 
<< pdiffusion >>
rect 248 87 249 88 
<< pdiffusion >>
rect 249 87 250 88 
<< pdiffusion >>
rect 250 87 251 88 
<< pdiffusion >>
rect 251 87 252 88 
<< m1 >>
rect 253 87 254 88 
<< m1 >>
rect 255 87 256 88 
<< pdiffusion >>
rect 264 87 265 88 
<< pdiffusion >>
rect 265 87 266 88 
<< pdiffusion >>
rect 266 87 267 88 
<< pdiffusion >>
rect 267 87 268 88 
<< pdiffusion >>
rect 268 87 269 88 
<< pdiffusion >>
rect 269 87 270 88 
<< m1 >>
rect 280 87 281 88 
<< pdiffusion >>
rect 282 87 283 88 
<< pdiffusion >>
rect 283 87 284 88 
<< pdiffusion >>
rect 284 87 285 88 
<< pdiffusion >>
rect 285 87 286 88 
<< pdiffusion >>
rect 286 87 287 88 
<< pdiffusion >>
rect 287 87 288 88 
<< pdiffusion >>
rect 300 87 301 88 
<< pdiffusion >>
rect 301 87 302 88 
<< pdiffusion >>
rect 302 87 303 88 
<< pdiffusion >>
rect 303 87 304 88 
<< pdiffusion >>
rect 304 87 305 88 
<< pdiffusion >>
rect 305 87 306 88 
<< m2 >>
rect 333 87 334 88 
<< m1 >>
rect 334 87 335 88 
<< pdiffusion >>
rect 336 87 337 88 
<< pdiffusion >>
rect 337 87 338 88 
<< pdiffusion >>
rect 338 87 339 88 
<< pdiffusion >>
rect 339 87 340 88 
<< pdiffusion >>
rect 340 87 341 88 
<< pdiffusion >>
rect 341 87 342 88 
<< m2 >>
rect 344 87 345 88 
<< m1 >>
rect 345 87 346 88 
<< pdiffusion >>
rect 354 87 355 88 
<< pdiffusion >>
rect 355 87 356 88 
<< pdiffusion >>
rect 356 87 357 88 
<< pdiffusion >>
rect 357 87 358 88 
<< pdiffusion >>
rect 358 87 359 88 
<< pdiffusion >>
rect 359 87 360 88 
<< m1 >>
rect 364 87 365 88 
<< m1 >>
rect 366 87 367 88 
<< m1 >>
rect 370 87 371 88 
<< pdiffusion >>
rect 372 87 373 88 
<< pdiffusion >>
rect 373 87 374 88 
<< pdiffusion >>
rect 374 87 375 88 
<< pdiffusion >>
rect 375 87 376 88 
<< pdiffusion >>
rect 376 87 377 88 
<< pdiffusion >>
rect 377 87 378 88 
<< pdiffusion >>
rect 390 87 391 88 
<< pdiffusion >>
rect 391 87 392 88 
<< pdiffusion >>
rect 392 87 393 88 
<< pdiffusion >>
rect 393 87 394 88 
<< pdiffusion >>
rect 394 87 395 88 
<< pdiffusion >>
rect 395 87 396 88 
<< pdiffusion >>
rect 408 87 409 88 
<< pdiffusion >>
rect 409 87 410 88 
<< pdiffusion >>
rect 410 87 411 88 
<< pdiffusion >>
rect 411 87 412 88 
<< pdiffusion >>
rect 412 87 413 88 
<< pdiffusion >>
rect 413 87 414 88 
<< m1 >>
rect 415 87 416 88 
<< m2 >>
rect 416 87 417 88 
<< pdiffusion >>
rect 426 87 427 88 
<< pdiffusion >>
rect 427 87 428 88 
<< pdiffusion >>
rect 428 87 429 88 
<< pdiffusion >>
rect 429 87 430 88 
<< pdiffusion >>
rect 430 87 431 88 
<< pdiffusion >>
rect 431 87 432 88 
<< m1 >>
rect 433 87 434 88 
<< pdiffusion >>
rect 444 87 445 88 
<< pdiffusion >>
rect 445 87 446 88 
<< pdiffusion >>
rect 446 87 447 88 
<< pdiffusion >>
rect 447 87 448 88 
<< pdiffusion >>
rect 448 87 449 88 
<< pdiffusion >>
rect 449 87 450 88 
<< m1 >>
rect 460 87 461 88 
<< pdiffusion >>
rect 462 87 463 88 
<< pdiffusion >>
rect 463 87 464 88 
<< pdiffusion >>
rect 464 87 465 88 
<< pdiffusion >>
rect 465 87 466 88 
<< pdiffusion >>
rect 466 87 467 88 
<< pdiffusion >>
rect 467 87 468 88 
<< pdiffusion >>
rect 480 87 481 88 
<< pdiffusion >>
rect 481 87 482 88 
<< pdiffusion >>
rect 482 87 483 88 
<< pdiffusion >>
rect 483 87 484 88 
<< pdiffusion >>
rect 484 87 485 88 
<< pdiffusion >>
rect 485 87 486 88 
<< m1 >>
rect 487 87 488 88 
<< m2 >>
rect 487 87 488 88 
<< pdiffusion >>
rect 516 87 517 88 
<< pdiffusion >>
rect 517 87 518 88 
<< pdiffusion >>
rect 518 87 519 88 
<< pdiffusion >>
rect 519 87 520 88 
<< pdiffusion >>
rect 520 87 521 88 
<< pdiffusion >>
rect 521 87 522 88 
<< pdiffusion >>
rect 12 88 13 89 
<< pdiffusion >>
rect 13 88 14 89 
<< pdiffusion >>
rect 14 88 15 89 
<< pdiffusion >>
rect 15 88 16 89 
<< pdiffusion >>
rect 16 88 17 89 
<< pdiffusion >>
rect 17 88 18 89 
<< pdiffusion >>
rect 30 88 31 89 
<< pdiffusion >>
rect 31 88 32 89 
<< pdiffusion >>
rect 32 88 33 89 
<< pdiffusion >>
rect 33 88 34 89 
<< pdiffusion >>
rect 34 88 35 89 
<< pdiffusion >>
rect 35 88 36 89 
<< pdiffusion >>
rect 48 88 49 89 
<< pdiffusion >>
rect 49 88 50 89 
<< pdiffusion >>
rect 50 88 51 89 
<< pdiffusion >>
rect 51 88 52 89 
<< pdiffusion >>
rect 52 88 53 89 
<< pdiffusion >>
rect 53 88 54 89 
<< m1 >>
rect 64 88 65 89 
<< pdiffusion >>
rect 66 88 67 89 
<< pdiffusion >>
rect 67 88 68 89 
<< pdiffusion >>
rect 68 88 69 89 
<< pdiffusion >>
rect 69 88 70 89 
<< pdiffusion >>
rect 70 88 71 89 
<< pdiffusion >>
rect 71 88 72 89 
<< m1 >>
rect 73 88 74 89 
<< pdiffusion >>
rect 84 88 85 89 
<< pdiffusion >>
rect 85 88 86 89 
<< pdiffusion >>
rect 86 88 87 89 
<< pdiffusion >>
rect 87 88 88 89 
<< pdiffusion >>
rect 88 88 89 89 
<< pdiffusion >>
rect 89 88 90 89 
<< m1 >>
rect 92 88 93 89 
<< m1 >>
rect 100 88 101 89 
<< m2 >>
rect 100 88 101 89 
<< pdiffusion >>
rect 102 88 103 89 
<< pdiffusion >>
rect 103 88 104 89 
<< pdiffusion >>
rect 104 88 105 89 
<< pdiffusion >>
rect 105 88 106 89 
<< pdiffusion >>
rect 106 88 107 89 
<< pdiffusion >>
rect 107 88 108 89 
<< pdiffusion >>
rect 120 88 121 89 
<< pdiffusion >>
rect 121 88 122 89 
<< pdiffusion >>
rect 122 88 123 89 
<< pdiffusion >>
rect 123 88 124 89 
<< pdiffusion >>
rect 124 88 125 89 
<< pdiffusion >>
rect 125 88 126 89 
<< m1 >>
rect 127 88 128 89 
<< m1 >>
rect 129 88 130 89 
<< m1 >>
rect 131 88 132 89 
<< m1 >>
rect 133 88 134 89 
<< pdiffusion >>
rect 138 88 139 89 
<< pdiffusion >>
rect 139 88 140 89 
<< pdiffusion >>
rect 140 88 141 89 
<< pdiffusion >>
rect 141 88 142 89 
<< pdiffusion >>
rect 142 88 143 89 
<< pdiffusion >>
rect 143 88 144 89 
<< m1 >>
rect 145 88 146 89 
<< pdiffusion >>
rect 156 88 157 89 
<< pdiffusion >>
rect 157 88 158 89 
<< pdiffusion >>
rect 158 88 159 89 
<< pdiffusion >>
rect 159 88 160 89 
<< pdiffusion >>
rect 160 88 161 89 
<< pdiffusion >>
rect 161 88 162 89 
<< m1 >>
rect 163 88 164 89 
<< pdiffusion >>
rect 174 88 175 89 
<< pdiffusion >>
rect 175 88 176 89 
<< pdiffusion >>
rect 176 88 177 89 
<< pdiffusion >>
rect 177 88 178 89 
<< pdiffusion >>
rect 178 88 179 89 
<< pdiffusion >>
rect 179 88 180 89 
<< m1 >>
rect 185 88 186 89 
<< m1 >>
rect 187 88 188 89 
<< pdiffusion >>
rect 192 88 193 89 
<< pdiffusion >>
rect 193 88 194 89 
<< pdiffusion >>
rect 194 88 195 89 
<< pdiffusion >>
rect 195 88 196 89 
<< pdiffusion >>
rect 196 88 197 89 
<< pdiffusion >>
rect 197 88 198 89 
<< m1 >>
rect 199 88 200 89 
<< pdiffusion >>
rect 210 88 211 89 
<< pdiffusion >>
rect 211 88 212 89 
<< pdiffusion >>
rect 212 88 213 89 
<< pdiffusion >>
rect 213 88 214 89 
<< pdiffusion >>
rect 214 88 215 89 
<< pdiffusion >>
rect 215 88 216 89 
<< m1 >>
rect 217 88 218 89 
<< m2 >>
rect 218 88 219 89 
<< m1 >>
rect 224 88 225 89 
<< pdiffusion >>
rect 228 88 229 89 
<< pdiffusion >>
rect 229 88 230 89 
<< pdiffusion >>
rect 230 88 231 89 
<< pdiffusion >>
rect 231 88 232 89 
<< pdiffusion >>
rect 232 88 233 89 
<< pdiffusion >>
rect 233 88 234 89 
<< m1 >>
rect 235 88 236 89 
<< m2 >>
rect 236 88 237 89 
<< m1 >>
rect 241 88 242 89 
<< pdiffusion >>
rect 246 88 247 89 
<< pdiffusion >>
rect 247 88 248 89 
<< pdiffusion >>
rect 248 88 249 89 
<< pdiffusion >>
rect 249 88 250 89 
<< pdiffusion >>
rect 250 88 251 89 
<< pdiffusion >>
rect 251 88 252 89 
<< m1 >>
rect 253 88 254 89 
<< m1 >>
rect 255 88 256 89 
<< pdiffusion >>
rect 264 88 265 89 
<< pdiffusion >>
rect 265 88 266 89 
<< pdiffusion >>
rect 266 88 267 89 
<< pdiffusion >>
rect 267 88 268 89 
<< pdiffusion >>
rect 268 88 269 89 
<< pdiffusion >>
rect 269 88 270 89 
<< m1 >>
rect 280 88 281 89 
<< pdiffusion >>
rect 282 88 283 89 
<< pdiffusion >>
rect 283 88 284 89 
<< pdiffusion >>
rect 284 88 285 89 
<< pdiffusion >>
rect 285 88 286 89 
<< pdiffusion >>
rect 286 88 287 89 
<< pdiffusion >>
rect 287 88 288 89 
<< pdiffusion >>
rect 300 88 301 89 
<< pdiffusion >>
rect 301 88 302 89 
<< pdiffusion >>
rect 302 88 303 89 
<< pdiffusion >>
rect 303 88 304 89 
<< pdiffusion >>
rect 304 88 305 89 
<< pdiffusion >>
rect 305 88 306 89 
<< m2 >>
rect 333 88 334 89 
<< m1 >>
rect 334 88 335 89 
<< pdiffusion >>
rect 336 88 337 89 
<< pdiffusion >>
rect 337 88 338 89 
<< pdiffusion >>
rect 338 88 339 89 
<< pdiffusion >>
rect 339 88 340 89 
<< pdiffusion >>
rect 340 88 341 89 
<< pdiffusion >>
rect 341 88 342 89 
<< m2 >>
rect 344 88 345 89 
<< m1 >>
rect 345 88 346 89 
<< pdiffusion >>
rect 354 88 355 89 
<< pdiffusion >>
rect 355 88 356 89 
<< pdiffusion >>
rect 356 88 357 89 
<< pdiffusion >>
rect 357 88 358 89 
<< pdiffusion >>
rect 358 88 359 89 
<< pdiffusion >>
rect 359 88 360 89 
<< m1 >>
rect 364 88 365 89 
<< m1 >>
rect 366 88 367 89 
<< m1 >>
rect 370 88 371 89 
<< pdiffusion >>
rect 372 88 373 89 
<< pdiffusion >>
rect 373 88 374 89 
<< pdiffusion >>
rect 374 88 375 89 
<< pdiffusion >>
rect 375 88 376 89 
<< pdiffusion >>
rect 376 88 377 89 
<< pdiffusion >>
rect 377 88 378 89 
<< pdiffusion >>
rect 390 88 391 89 
<< pdiffusion >>
rect 391 88 392 89 
<< pdiffusion >>
rect 392 88 393 89 
<< pdiffusion >>
rect 393 88 394 89 
<< pdiffusion >>
rect 394 88 395 89 
<< pdiffusion >>
rect 395 88 396 89 
<< pdiffusion >>
rect 408 88 409 89 
<< pdiffusion >>
rect 409 88 410 89 
<< pdiffusion >>
rect 410 88 411 89 
<< pdiffusion >>
rect 411 88 412 89 
<< pdiffusion >>
rect 412 88 413 89 
<< pdiffusion >>
rect 413 88 414 89 
<< m1 >>
rect 415 88 416 89 
<< m2 >>
rect 416 88 417 89 
<< pdiffusion >>
rect 426 88 427 89 
<< pdiffusion >>
rect 427 88 428 89 
<< pdiffusion >>
rect 428 88 429 89 
<< pdiffusion >>
rect 429 88 430 89 
<< pdiffusion >>
rect 430 88 431 89 
<< pdiffusion >>
rect 431 88 432 89 
<< m1 >>
rect 433 88 434 89 
<< pdiffusion >>
rect 444 88 445 89 
<< pdiffusion >>
rect 445 88 446 89 
<< pdiffusion >>
rect 446 88 447 89 
<< pdiffusion >>
rect 447 88 448 89 
<< pdiffusion >>
rect 448 88 449 89 
<< pdiffusion >>
rect 449 88 450 89 
<< m1 >>
rect 460 88 461 89 
<< pdiffusion >>
rect 462 88 463 89 
<< pdiffusion >>
rect 463 88 464 89 
<< pdiffusion >>
rect 464 88 465 89 
<< pdiffusion >>
rect 465 88 466 89 
<< pdiffusion >>
rect 466 88 467 89 
<< pdiffusion >>
rect 467 88 468 89 
<< pdiffusion >>
rect 480 88 481 89 
<< pdiffusion >>
rect 481 88 482 89 
<< pdiffusion >>
rect 482 88 483 89 
<< pdiffusion >>
rect 483 88 484 89 
<< pdiffusion >>
rect 484 88 485 89 
<< pdiffusion >>
rect 485 88 486 89 
<< m1 >>
rect 487 88 488 89 
<< m2 >>
rect 487 88 488 89 
<< pdiffusion >>
rect 516 88 517 89 
<< pdiffusion >>
rect 517 88 518 89 
<< pdiffusion >>
rect 518 88 519 89 
<< pdiffusion >>
rect 519 88 520 89 
<< pdiffusion >>
rect 520 88 521 89 
<< pdiffusion >>
rect 521 88 522 89 
<< pdiffusion >>
rect 12 89 13 90 
<< pdiffusion >>
rect 13 89 14 90 
<< pdiffusion >>
rect 14 89 15 90 
<< pdiffusion >>
rect 15 89 16 90 
<< pdiffusion >>
rect 16 89 17 90 
<< pdiffusion >>
rect 17 89 18 90 
<< pdiffusion >>
rect 30 89 31 90 
<< pdiffusion >>
rect 31 89 32 90 
<< pdiffusion >>
rect 32 89 33 90 
<< pdiffusion >>
rect 33 89 34 90 
<< pdiffusion >>
rect 34 89 35 90 
<< pdiffusion >>
rect 35 89 36 90 
<< pdiffusion >>
rect 48 89 49 90 
<< m1 >>
rect 49 89 50 90 
<< pdiffusion >>
rect 49 89 50 90 
<< pdiffusion >>
rect 50 89 51 90 
<< pdiffusion >>
rect 51 89 52 90 
<< pdiffusion >>
rect 52 89 53 90 
<< pdiffusion >>
rect 53 89 54 90 
<< m1 >>
rect 64 89 65 90 
<< pdiffusion >>
rect 66 89 67 90 
<< pdiffusion >>
rect 67 89 68 90 
<< pdiffusion >>
rect 68 89 69 90 
<< pdiffusion >>
rect 69 89 70 90 
<< pdiffusion >>
rect 70 89 71 90 
<< pdiffusion >>
rect 71 89 72 90 
<< m1 >>
rect 73 89 74 90 
<< pdiffusion >>
rect 84 89 85 90 
<< pdiffusion >>
rect 85 89 86 90 
<< pdiffusion >>
rect 86 89 87 90 
<< pdiffusion >>
rect 87 89 88 90 
<< m1 >>
rect 88 89 89 90 
<< pdiffusion >>
rect 88 89 89 90 
<< pdiffusion >>
rect 89 89 90 90 
<< m1 >>
rect 92 89 93 90 
<< m1 >>
rect 100 89 101 90 
<< m2 >>
rect 100 89 101 90 
<< pdiffusion >>
rect 102 89 103 90 
<< pdiffusion >>
rect 103 89 104 90 
<< pdiffusion >>
rect 104 89 105 90 
<< pdiffusion >>
rect 105 89 106 90 
<< pdiffusion >>
rect 106 89 107 90 
<< pdiffusion >>
rect 107 89 108 90 
<< pdiffusion >>
rect 120 89 121 90 
<< pdiffusion >>
rect 121 89 122 90 
<< pdiffusion >>
rect 122 89 123 90 
<< pdiffusion >>
rect 123 89 124 90 
<< pdiffusion >>
rect 124 89 125 90 
<< pdiffusion >>
rect 125 89 126 90 
<< m1 >>
rect 127 89 128 90 
<< m1 >>
rect 129 89 130 90 
<< m1 >>
rect 131 89 132 90 
<< m1 >>
rect 133 89 134 90 
<< pdiffusion >>
rect 138 89 139 90 
<< pdiffusion >>
rect 139 89 140 90 
<< pdiffusion >>
rect 140 89 141 90 
<< pdiffusion >>
rect 141 89 142 90 
<< pdiffusion >>
rect 142 89 143 90 
<< pdiffusion >>
rect 143 89 144 90 
<< m1 >>
rect 145 89 146 90 
<< pdiffusion >>
rect 156 89 157 90 
<< pdiffusion >>
rect 157 89 158 90 
<< pdiffusion >>
rect 158 89 159 90 
<< pdiffusion >>
rect 159 89 160 90 
<< pdiffusion >>
rect 160 89 161 90 
<< pdiffusion >>
rect 161 89 162 90 
<< m1 >>
rect 163 89 164 90 
<< pdiffusion >>
rect 174 89 175 90 
<< pdiffusion >>
rect 175 89 176 90 
<< pdiffusion >>
rect 176 89 177 90 
<< pdiffusion >>
rect 177 89 178 90 
<< m1 >>
rect 178 89 179 90 
<< pdiffusion >>
rect 178 89 179 90 
<< pdiffusion >>
rect 179 89 180 90 
<< m1 >>
rect 185 89 186 90 
<< m1 >>
rect 187 89 188 90 
<< pdiffusion >>
rect 192 89 193 90 
<< pdiffusion >>
rect 193 89 194 90 
<< pdiffusion >>
rect 194 89 195 90 
<< pdiffusion >>
rect 195 89 196 90 
<< pdiffusion >>
rect 196 89 197 90 
<< pdiffusion >>
rect 197 89 198 90 
<< m1 >>
rect 199 89 200 90 
<< pdiffusion >>
rect 210 89 211 90 
<< pdiffusion >>
rect 211 89 212 90 
<< pdiffusion >>
rect 212 89 213 90 
<< pdiffusion >>
rect 213 89 214 90 
<< m1 >>
rect 214 89 215 90 
<< pdiffusion >>
rect 214 89 215 90 
<< pdiffusion >>
rect 215 89 216 90 
<< m1 >>
rect 217 89 218 90 
<< m2 >>
rect 218 89 219 90 
<< m1 >>
rect 224 89 225 90 
<< pdiffusion >>
rect 228 89 229 90 
<< pdiffusion >>
rect 229 89 230 90 
<< pdiffusion >>
rect 230 89 231 90 
<< pdiffusion >>
rect 231 89 232 90 
<< pdiffusion >>
rect 232 89 233 90 
<< pdiffusion >>
rect 233 89 234 90 
<< m1 >>
rect 235 89 236 90 
<< m2 >>
rect 236 89 237 90 
<< m1 >>
rect 241 89 242 90 
<< pdiffusion >>
rect 246 89 247 90 
<< m1 >>
rect 247 89 248 90 
<< pdiffusion >>
rect 247 89 248 90 
<< pdiffusion >>
rect 248 89 249 90 
<< pdiffusion >>
rect 249 89 250 90 
<< pdiffusion >>
rect 250 89 251 90 
<< pdiffusion >>
rect 251 89 252 90 
<< m1 >>
rect 253 89 254 90 
<< m1 >>
rect 255 89 256 90 
<< pdiffusion >>
rect 264 89 265 90 
<< pdiffusion >>
rect 265 89 266 90 
<< pdiffusion >>
rect 266 89 267 90 
<< pdiffusion >>
rect 267 89 268 90 
<< pdiffusion >>
rect 268 89 269 90 
<< pdiffusion >>
rect 269 89 270 90 
<< m1 >>
rect 280 89 281 90 
<< pdiffusion >>
rect 282 89 283 90 
<< pdiffusion >>
rect 283 89 284 90 
<< pdiffusion >>
rect 284 89 285 90 
<< pdiffusion >>
rect 285 89 286 90 
<< m1 >>
rect 286 89 287 90 
<< pdiffusion >>
rect 286 89 287 90 
<< pdiffusion >>
rect 287 89 288 90 
<< pdiffusion >>
rect 300 89 301 90 
<< pdiffusion >>
rect 301 89 302 90 
<< pdiffusion >>
rect 302 89 303 90 
<< pdiffusion >>
rect 303 89 304 90 
<< m1 >>
rect 304 89 305 90 
<< pdiffusion >>
rect 304 89 305 90 
<< pdiffusion >>
rect 305 89 306 90 
<< m2 >>
rect 333 89 334 90 
<< m1 >>
rect 334 89 335 90 
<< pdiffusion >>
rect 336 89 337 90 
<< m1 >>
rect 337 89 338 90 
<< pdiffusion >>
rect 337 89 338 90 
<< pdiffusion >>
rect 338 89 339 90 
<< pdiffusion >>
rect 339 89 340 90 
<< pdiffusion >>
rect 340 89 341 90 
<< pdiffusion >>
rect 341 89 342 90 
<< m2 >>
rect 344 89 345 90 
<< m1 >>
rect 345 89 346 90 
<< pdiffusion >>
rect 354 89 355 90 
<< pdiffusion >>
rect 355 89 356 90 
<< pdiffusion >>
rect 356 89 357 90 
<< pdiffusion >>
rect 357 89 358 90 
<< m1 >>
rect 358 89 359 90 
<< pdiffusion >>
rect 358 89 359 90 
<< pdiffusion >>
rect 359 89 360 90 
<< m1 >>
rect 364 89 365 90 
<< m1 >>
rect 366 89 367 90 
<< m1 >>
rect 370 89 371 90 
<< pdiffusion >>
rect 372 89 373 90 
<< pdiffusion >>
rect 373 89 374 90 
<< pdiffusion >>
rect 374 89 375 90 
<< pdiffusion >>
rect 375 89 376 90 
<< pdiffusion >>
rect 376 89 377 90 
<< pdiffusion >>
rect 377 89 378 90 
<< pdiffusion >>
rect 390 89 391 90 
<< pdiffusion >>
rect 391 89 392 90 
<< pdiffusion >>
rect 392 89 393 90 
<< pdiffusion >>
rect 393 89 394 90 
<< m1 >>
rect 394 89 395 90 
<< pdiffusion >>
rect 394 89 395 90 
<< pdiffusion >>
rect 395 89 396 90 
<< pdiffusion >>
rect 408 89 409 90 
<< pdiffusion >>
rect 409 89 410 90 
<< pdiffusion >>
rect 410 89 411 90 
<< pdiffusion >>
rect 411 89 412 90 
<< pdiffusion >>
rect 412 89 413 90 
<< pdiffusion >>
rect 413 89 414 90 
<< m1 >>
rect 415 89 416 90 
<< m2 >>
rect 416 89 417 90 
<< pdiffusion >>
rect 426 89 427 90 
<< pdiffusion >>
rect 427 89 428 90 
<< pdiffusion >>
rect 428 89 429 90 
<< pdiffusion >>
rect 429 89 430 90 
<< pdiffusion >>
rect 430 89 431 90 
<< pdiffusion >>
rect 431 89 432 90 
<< m1 >>
rect 433 89 434 90 
<< pdiffusion >>
rect 444 89 445 90 
<< pdiffusion >>
rect 445 89 446 90 
<< pdiffusion >>
rect 446 89 447 90 
<< pdiffusion >>
rect 447 89 448 90 
<< m1 >>
rect 448 89 449 90 
<< pdiffusion >>
rect 448 89 449 90 
<< pdiffusion >>
rect 449 89 450 90 
<< m1 >>
rect 460 89 461 90 
<< pdiffusion >>
rect 462 89 463 90 
<< pdiffusion >>
rect 463 89 464 90 
<< pdiffusion >>
rect 464 89 465 90 
<< pdiffusion >>
rect 465 89 466 90 
<< m1 >>
rect 466 89 467 90 
<< pdiffusion >>
rect 466 89 467 90 
<< pdiffusion >>
rect 467 89 468 90 
<< pdiffusion >>
rect 480 89 481 90 
<< m1 >>
rect 481 89 482 90 
<< pdiffusion >>
rect 481 89 482 90 
<< pdiffusion >>
rect 482 89 483 90 
<< pdiffusion >>
rect 483 89 484 90 
<< pdiffusion >>
rect 484 89 485 90 
<< pdiffusion >>
rect 485 89 486 90 
<< m1 >>
rect 487 89 488 90 
<< m2 >>
rect 487 89 488 90 
<< pdiffusion >>
rect 516 89 517 90 
<< pdiffusion >>
rect 517 89 518 90 
<< pdiffusion >>
rect 518 89 519 90 
<< pdiffusion >>
rect 519 89 520 90 
<< pdiffusion >>
rect 520 89 521 90 
<< pdiffusion >>
rect 521 89 522 90 
<< m1 >>
rect 49 90 50 91 
<< m1 >>
rect 64 90 65 91 
<< m1 >>
rect 73 90 74 91 
<< m1 >>
rect 88 90 89 91 
<< m1 >>
rect 92 90 93 91 
<< m1 >>
rect 100 90 101 91 
<< m2 >>
rect 100 90 101 91 
<< m1 >>
rect 127 90 128 91 
<< m1 >>
rect 129 90 130 91 
<< m1 >>
rect 131 90 132 91 
<< m1 >>
rect 133 90 134 91 
<< m1 >>
rect 145 90 146 91 
<< m1 >>
rect 163 90 164 91 
<< m1 >>
rect 178 90 179 91 
<< m1 >>
rect 185 90 186 91 
<< m1 >>
rect 187 90 188 91 
<< m1 >>
rect 199 90 200 91 
<< m1 >>
rect 214 90 215 91 
<< m1 >>
rect 217 90 218 91 
<< m2 >>
rect 218 90 219 91 
<< m1 >>
rect 224 90 225 91 
<< m2 >>
rect 224 90 225 91 
<< m2c >>
rect 224 90 225 91 
<< m1 >>
rect 224 90 225 91 
<< m2 >>
rect 224 90 225 91 
<< m1 >>
rect 235 90 236 91 
<< m2 >>
rect 236 90 237 91 
<< m1 >>
rect 241 90 242 91 
<< m1 >>
rect 247 90 248 91 
<< m1 >>
rect 253 90 254 91 
<< m1 >>
rect 255 90 256 91 
<< m1 >>
rect 280 90 281 91 
<< m1 >>
rect 286 90 287 91 
<< m1 >>
rect 304 90 305 91 
<< m2 >>
rect 333 90 334 91 
<< m1 >>
rect 334 90 335 91 
<< m1 >>
rect 337 90 338 91 
<< m2 >>
rect 344 90 345 91 
<< m1 >>
rect 345 90 346 91 
<< m1 >>
rect 358 90 359 91 
<< m2 >>
rect 362 90 363 91 
<< m1 >>
rect 363 90 364 91 
<< m2 >>
rect 363 90 364 91 
<< m2c >>
rect 363 90 364 91 
<< m1 >>
rect 363 90 364 91 
<< m2 >>
rect 363 90 364 91 
<< m1 >>
rect 364 90 365 91 
<< m1 >>
rect 366 90 367 91 
<< m1 >>
rect 370 90 371 91 
<< m1 >>
rect 394 90 395 91 
<< m1 >>
rect 415 90 416 91 
<< m2 >>
rect 416 90 417 91 
<< m1 >>
rect 433 90 434 91 
<< m1 >>
rect 448 90 449 91 
<< m1 >>
rect 460 90 461 91 
<< m1 >>
rect 466 90 467 91 
<< m1 >>
rect 481 90 482 91 
<< m1 >>
rect 487 90 488 91 
<< m2 >>
rect 487 90 488 91 
<< m1 >>
rect 49 91 50 92 
<< m1 >>
rect 64 91 65 92 
<< m1 >>
rect 73 91 74 92 
<< m1 >>
rect 88 91 89 92 
<< m1 >>
rect 92 91 93 92 
<< m1 >>
rect 100 91 101 92 
<< m2 >>
rect 100 91 101 92 
<< m1 >>
rect 127 91 128 92 
<< m1 >>
rect 129 91 130 92 
<< m1 >>
rect 131 91 132 92 
<< m1 >>
rect 133 91 134 92 
<< m1 >>
rect 145 91 146 92 
<< m1 >>
rect 163 91 164 92 
<< m1 >>
rect 178 91 179 92 
<< m2 >>
rect 179 91 180 92 
<< m1 >>
rect 180 91 181 92 
<< m2 >>
rect 180 91 181 92 
<< m2c >>
rect 180 91 181 92 
<< m1 >>
rect 180 91 181 92 
<< m2 >>
rect 180 91 181 92 
<< m1 >>
rect 181 91 182 92 
<< m1 >>
rect 182 91 183 92 
<< m1 >>
rect 183 91 184 92 
<< m1 >>
rect 184 91 185 92 
<< m1 >>
rect 185 91 186 92 
<< m1 >>
rect 187 91 188 92 
<< m1 >>
rect 199 91 200 92 
<< m1 >>
rect 214 91 215 92 
<< m1 >>
rect 215 91 216 92 
<< m1 >>
rect 216 91 217 92 
<< m1 >>
rect 217 91 218 92 
<< m2 >>
rect 218 91 219 92 
<< m2 >>
rect 224 91 225 92 
<< m1 >>
rect 233 91 234 92 
<< m2 >>
rect 233 91 234 92 
<< m2c >>
rect 233 91 234 92 
<< m1 >>
rect 233 91 234 92 
<< m2 >>
rect 233 91 234 92 
<< m2 >>
rect 234 91 235 92 
<< m1 >>
rect 235 91 236 92 
<< m2 >>
rect 235 91 236 92 
<< m2 >>
rect 236 91 237 92 
<< m1 >>
rect 241 91 242 92 
<< m1 >>
rect 247 91 248 92 
<< m1 >>
rect 251 91 252 92 
<< m2 >>
rect 251 91 252 92 
<< m2c >>
rect 251 91 252 92 
<< m1 >>
rect 251 91 252 92 
<< m2 >>
rect 251 91 252 92 
<< m1 >>
rect 252 91 253 92 
<< m1 >>
rect 253 91 254 92 
<< m1 >>
rect 255 91 256 92 
<< m1 >>
rect 280 91 281 92 
<< m1 >>
rect 286 91 287 92 
<< m1 >>
rect 304 91 305 92 
<< m2 >>
rect 333 91 334 92 
<< m1 >>
rect 334 91 335 92 
<< m2 >>
rect 334 91 335 92 
<< m2 >>
rect 335 91 336 92 
<< m1 >>
rect 336 91 337 92 
<< m2 >>
rect 336 91 337 92 
<< m2c >>
rect 336 91 337 92 
<< m1 >>
rect 336 91 337 92 
<< m2 >>
rect 336 91 337 92 
<< m1 >>
rect 337 91 338 92 
<< m2 >>
rect 344 91 345 92 
<< m1 >>
rect 345 91 346 92 
<< m1 >>
rect 358 91 359 92 
<< m1 >>
rect 359 91 360 92 
<< m1 >>
rect 360 91 361 92 
<< m1 >>
rect 361 91 362 92 
<< m2 >>
rect 362 91 363 92 
<< m1 >>
rect 366 91 367 92 
<< m1 >>
rect 370 91 371 92 
<< m1 >>
rect 394 91 395 92 
<< m1 >>
rect 415 91 416 92 
<< m2 >>
rect 416 91 417 92 
<< m1 >>
rect 417 91 418 92 
<< m2 >>
rect 417 91 418 92 
<< m2c >>
rect 417 91 418 92 
<< m1 >>
rect 417 91 418 92 
<< m2 >>
rect 417 91 418 92 
<< m1 >>
rect 418 91 419 92 
<< m1 >>
rect 419 91 420 92 
<< m1 >>
rect 420 91 421 92 
<< m1 >>
rect 421 91 422 92 
<< m1 >>
rect 422 91 423 92 
<< m1 >>
rect 423 91 424 92 
<< m1 >>
rect 424 91 425 92 
<< m1 >>
rect 425 91 426 92 
<< m1 >>
rect 426 91 427 92 
<< m2 >>
rect 426 91 427 92 
<< m2c >>
rect 426 91 427 92 
<< m1 >>
rect 426 91 427 92 
<< m2 >>
rect 426 91 427 92 
<< m1 >>
rect 433 91 434 92 
<< m1 >>
rect 448 91 449 92 
<< m1 >>
rect 460 91 461 92 
<< m1 >>
rect 466 91 467 92 
<< m2 >>
rect 467 91 468 92 
<< m1 >>
rect 468 91 469 92 
<< m2 >>
rect 468 91 469 92 
<< m2c >>
rect 468 91 469 92 
<< m1 >>
rect 468 91 469 92 
<< m2 >>
rect 468 91 469 92 
<< m1 >>
rect 469 91 470 92 
<< m1 >>
rect 470 91 471 92 
<< m1 >>
rect 471 91 472 92 
<< m1 >>
rect 472 91 473 92 
<< m1 >>
rect 473 91 474 92 
<< m1 >>
rect 474 91 475 92 
<< m1 >>
rect 475 91 476 92 
<< m1 >>
rect 476 91 477 92 
<< m1 >>
rect 477 91 478 92 
<< m1 >>
rect 478 91 479 92 
<< m1 >>
rect 479 91 480 92 
<< m1 >>
rect 480 91 481 92 
<< m1 >>
rect 481 91 482 92 
<< m1 >>
rect 485 91 486 92 
<< m2 >>
rect 485 91 486 92 
<< m2c >>
rect 485 91 486 92 
<< m1 >>
rect 485 91 486 92 
<< m2 >>
rect 485 91 486 92 
<< m2 >>
rect 486 91 487 92 
<< m1 >>
rect 487 91 488 92 
<< m2 >>
rect 487 91 488 92 
<< m1 >>
rect 49 92 50 93 
<< m1 >>
rect 64 92 65 93 
<< m1 >>
rect 73 92 74 93 
<< m1 >>
rect 88 92 89 93 
<< m1 >>
rect 92 92 93 93 
<< m1 >>
rect 100 92 101 93 
<< m2 >>
rect 100 92 101 93 
<< m1 >>
rect 127 92 128 93 
<< m1 >>
rect 129 92 130 93 
<< m1 >>
rect 131 92 132 93 
<< m1 >>
rect 133 92 134 93 
<< m1 >>
rect 145 92 146 93 
<< m1 >>
rect 163 92 164 93 
<< m1 >>
rect 178 92 179 93 
<< m2 >>
rect 179 92 180 93 
<< m1 >>
rect 187 92 188 93 
<< m1 >>
rect 194 92 195 93 
<< m2 >>
rect 194 92 195 93 
<< m2c >>
rect 194 92 195 93 
<< m1 >>
rect 194 92 195 93 
<< m2 >>
rect 194 92 195 93 
<< m1 >>
rect 195 92 196 93 
<< m1 >>
rect 196 92 197 93 
<< m1 >>
rect 197 92 198 93 
<< m1 >>
rect 198 92 199 93 
<< m1 >>
rect 199 92 200 93 
<< m2 >>
rect 218 92 219 93 
<< m1 >>
rect 219 92 220 93 
<< m2 >>
rect 219 92 220 93 
<< m2c >>
rect 219 92 220 93 
<< m1 >>
rect 219 92 220 93 
<< m2 >>
rect 219 92 220 93 
<< m1 >>
rect 220 92 221 93 
<< m1 >>
rect 221 92 222 93 
<< m1 >>
rect 222 92 223 93 
<< m1 >>
rect 223 92 224 93 
<< m1 >>
rect 224 92 225 93 
<< m2 >>
rect 224 92 225 93 
<< m1 >>
rect 225 92 226 93 
<< m1 >>
rect 226 92 227 93 
<< m1 >>
rect 227 92 228 93 
<< m1 >>
rect 228 92 229 93 
<< m1 >>
rect 233 92 234 93 
<< m1 >>
rect 235 92 236 93 
<< m1 >>
rect 241 92 242 93 
<< m1 >>
rect 247 92 248 93 
<< m2 >>
rect 247 92 248 93 
<< m2c >>
rect 247 92 248 93 
<< m1 >>
rect 247 92 248 93 
<< m2 >>
rect 247 92 248 93 
<< m2 >>
rect 248 92 249 93 
<< m2 >>
rect 249 92 250 93 
<< m2 >>
rect 250 92 251 93 
<< m2 >>
rect 251 92 252 93 
<< m1 >>
rect 255 92 256 93 
<< m1 >>
rect 280 92 281 93 
<< m2 >>
rect 280 92 281 93 
<< m2c >>
rect 280 92 281 93 
<< m1 >>
rect 280 92 281 93 
<< m2 >>
rect 280 92 281 93 
<< m1 >>
rect 286 92 287 93 
<< m1 >>
rect 304 92 305 93 
<< m1 >>
rect 334 92 335 93 
<< m2 >>
rect 344 92 345 93 
<< m1 >>
rect 345 92 346 93 
<< m2 >>
rect 357 92 358 93 
<< m2 >>
rect 358 92 359 93 
<< m2 >>
rect 359 92 360 93 
<< m2 >>
rect 360 92 361 93 
<< m1 >>
rect 361 92 362 93 
<< m2 >>
rect 361 92 362 93 
<< m2 >>
rect 362 92 363 93 
<< m1 >>
rect 366 92 367 93 
<< m2 >>
rect 366 92 367 93 
<< m2c >>
rect 366 92 367 93 
<< m1 >>
rect 366 92 367 93 
<< m2 >>
rect 366 92 367 93 
<< m1 >>
rect 370 92 371 93 
<< m1 >>
rect 394 92 395 93 
<< m1 >>
rect 415 92 416 93 
<< m2 >>
rect 426 92 427 93 
<< m1 >>
rect 433 92 434 93 
<< m1 >>
rect 448 92 449 93 
<< m1 >>
rect 460 92 461 93 
<< m1 >>
rect 464 92 465 93 
<< m2 >>
rect 464 92 465 93 
<< m2c >>
rect 464 92 465 93 
<< m1 >>
rect 464 92 465 93 
<< m2 >>
rect 464 92 465 93 
<< m2 >>
rect 465 92 466 93 
<< m1 >>
rect 466 92 467 93 
<< m2 >>
rect 466 92 467 93 
<< m2 >>
rect 467 92 468 93 
<< m1 >>
rect 485 92 486 93 
<< m1 >>
rect 487 92 488 93 
<< m1 >>
rect 49 93 50 94 
<< m1 >>
rect 64 93 65 94 
<< m2 >>
rect 64 93 65 94 
<< m2c >>
rect 64 93 65 94 
<< m1 >>
rect 64 93 65 94 
<< m2 >>
rect 64 93 65 94 
<< m1 >>
rect 73 93 74 94 
<< m1 >>
rect 88 93 89 94 
<< m1 >>
rect 92 93 93 94 
<< m1 >>
rect 100 93 101 94 
<< m2 >>
rect 100 93 101 94 
<< m1 >>
rect 127 93 128 94 
<< m1 >>
rect 129 93 130 94 
<< m1 >>
rect 131 93 132 94 
<< m1 >>
rect 133 93 134 94 
<< m1 >>
rect 145 93 146 94 
<< m1 >>
rect 163 93 164 94 
<< m1 >>
rect 178 93 179 94 
<< m2 >>
rect 179 93 180 94 
<< m1 >>
rect 187 93 188 94 
<< m2 >>
rect 194 93 195 94 
<< m2 >>
rect 224 93 225 94 
<< m1 >>
rect 228 93 229 94 
<< m1 >>
rect 233 93 234 94 
<< m1 >>
rect 235 93 236 94 
<< m1 >>
rect 241 93 242 94 
<< m2 >>
rect 241 93 242 94 
<< m2c >>
rect 241 93 242 94 
<< m1 >>
rect 241 93 242 94 
<< m2 >>
rect 241 93 242 94 
<< m1 >>
rect 248 93 249 94 
<< m1 >>
rect 249 93 250 94 
<< m1 >>
rect 250 93 251 94 
<< m1 >>
rect 251 93 252 94 
<< m1 >>
rect 252 93 253 94 
<< m1 >>
rect 253 93 254 94 
<< m2 >>
rect 253 93 254 94 
<< m2c >>
rect 253 93 254 94 
<< m1 >>
rect 253 93 254 94 
<< m2 >>
rect 253 93 254 94 
<< m2 >>
rect 254 93 255 94 
<< m1 >>
rect 255 93 256 94 
<< m2 >>
rect 255 93 256 94 
<< m2 >>
rect 256 93 257 94 
<< m1 >>
rect 257 93 258 94 
<< m2 >>
rect 257 93 258 94 
<< m2c >>
rect 257 93 258 94 
<< m1 >>
rect 257 93 258 94 
<< m2 >>
rect 257 93 258 94 
<< m2 >>
rect 280 93 281 94 
<< m1 >>
rect 286 93 287 94 
<< m1 >>
rect 304 93 305 94 
<< m1 >>
rect 334 93 335 94 
<< m2 >>
rect 344 93 345 94 
<< m1 >>
rect 345 93 346 94 
<< m2 >>
rect 357 93 358 94 
<< m1 >>
rect 361 93 362 94 
<< m2 >>
rect 366 93 367 94 
<< m1 >>
rect 370 93 371 94 
<< m1 >>
rect 394 93 395 94 
<< m1 >>
rect 413 93 414 94 
<< m2 >>
rect 413 93 414 94 
<< m2c >>
rect 413 93 414 94 
<< m1 >>
rect 413 93 414 94 
<< m2 >>
rect 413 93 414 94 
<< m2 >>
rect 414 93 415 94 
<< m1 >>
rect 415 93 416 94 
<< m2 >>
rect 415 93 416 94 
<< m2 >>
rect 416 93 417 94 
<< m1 >>
rect 417 93 418 94 
<< m2 >>
rect 417 93 418 94 
<< m2c >>
rect 417 93 418 94 
<< m1 >>
rect 417 93 418 94 
<< m2 >>
rect 417 93 418 94 
<< m1 >>
rect 418 93 419 94 
<< m1 >>
rect 419 93 420 94 
<< m1 >>
rect 420 93 421 94 
<< m1 >>
rect 421 93 422 94 
<< m1 >>
rect 422 93 423 94 
<< m1 >>
rect 423 93 424 94 
<< m1 >>
rect 424 93 425 94 
<< m1 >>
rect 425 93 426 94 
<< m1 >>
rect 426 93 427 94 
<< m2 >>
rect 426 93 427 94 
<< m1 >>
rect 433 93 434 94 
<< m1 >>
rect 448 93 449 94 
<< m2 >>
rect 449 93 450 94 
<< m1 >>
rect 450 93 451 94 
<< m2 >>
rect 450 93 451 94 
<< m2c >>
rect 450 93 451 94 
<< m1 >>
rect 450 93 451 94 
<< m2 >>
rect 450 93 451 94 
<< m1 >>
rect 451 93 452 94 
<< m1 >>
rect 452 93 453 94 
<< m1 >>
rect 453 93 454 94 
<< m1 >>
rect 454 93 455 94 
<< m1 >>
rect 455 93 456 94 
<< m1 >>
rect 456 93 457 94 
<< m1 >>
rect 457 93 458 94 
<< m1 >>
rect 458 93 459 94 
<< m2 >>
rect 458 93 459 94 
<< m2c >>
rect 458 93 459 94 
<< m1 >>
rect 458 93 459 94 
<< m2 >>
rect 458 93 459 94 
<< m2 >>
rect 459 93 460 94 
<< m1 >>
rect 460 93 461 94 
<< m2 >>
rect 460 93 461 94 
<< m2 >>
rect 461 93 462 94 
<< m1 >>
rect 462 93 463 94 
<< m2 >>
rect 462 93 463 94 
<< m2c >>
rect 462 93 463 94 
<< m1 >>
rect 462 93 463 94 
<< m2 >>
rect 462 93 463 94 
<< m1 >>
rect 464 93 465 94 
<< m1 >>
rect 466 93 467 94 
<< m1 >>
rect 485 93 486 94 
<< m1 >>
rect 487 93 488 94 
<< m1 >>
rect 49 94 50 95 
<< m2 >>
rect 64 94 65 95 
<< m1 >>
rect 73 94 74 95 
<< m1 >>
rect 88 94 89 95 
<< m1 >>
rect 92 94 93 95 
<< m1 >>
rect 100 94 101 95 
<< m2 >>
rect 100 94 101 95 
<< m1 >>
rect 127 94 128 95 
<< m1 >>
rect 129 94 130 95 
<< m1 >>
rect 131 94 132 95 
<< m1 >>
rect 133 94 134 95 
<< m1 >>
rect 134 94 135 95 
<< m1 >>
rect 135 94 136 95 
<< m1 >>
rect 136 94 137 95 
<< m1 >>
rect 137 94 138 95 
<< m1 >>
rect 138 94 139 95 
<< m1 >>
rect 139 94 140 95 
<< m1 >>
rect 140 94 141 95 
<< m1 >>
rect 141 94 142 95 
<< m1 >>
rect 142 94 143 95 
<< m1 >>
rect 143 94 144 95 
<< m2 >>
rect 143 94 144 95 
<< m2c >>
rect 143 94 144 95 
<< m1 >>
rect 143 94 144 95 
<< m2 >>
rect 143 94 144 95 
<< m2 >>
rect 144 94 145 95 
<< m1 >>
rect 145 94 146 95 
<< m2 >>
rect 145 94 146 95 
<< m2 >>
rect 146 94 147 95 
<< m1 >>
rect 147 94 148 95 
<< m2 >>
rect 147 94 148 95 
<< m2c >>
rect 147 94 148 95 
<< m1 >>
rect 147 94 148 95 
<< m2 >>
rect 147 94 148 95 
<< m1 >>
rect 148 94 149 95 
<< m1 >>
rect 149 94 150 95 
<< m1 >>
rect 163 94 164 95 
<< m1 >>
rect 164 94 165 95 
<< m1 >>
rect 165 94 166 95 
<< m1 >>
rect 166 94 167 95 
<< m1 >>
rect 167 94 168 95 
<< m1 >>
rect 168 94 169 95 
<< m1 >>
rect 169 94 170 95 
<< m1 >>
rect 170 94 171 95 
<< m1 >>
rect 171 94 172 95 
<< m1 >>
rect 172 94 173 95 
<< m1 >>
rect 173 94 174 95 
<< m1 >>
rect 174 94 175 95 
<< m2 >>
rect 174 94 175 95 
<< m1 >>
rect 175 94 176 95 
<< m2 >>
rect 175 94 176 95 
<< m1 >>
rect 176 94 177 95 
<< m2 >>
rect 176 94 177 95 
<< m1 >>
rect 177 94 178 95 
<< m2 >>
rect 177 94 178 95 
<< m1 >>
rect 178 94 179 95 
<< m2 >>
rect 178 94 179 95 
<< m2 >>
rect 179 94 180 95 
<< m1 >>
rect 187 94 188 95 
<< m1 >>
rect 190 94 191 95 
<< m1 >>
rect 191 94 192 95 
<< m1 >>
rect 192 94 193 95 
<< m1 >>
rect 193 94 194 95 
<< m1 >>
rect 194 94 195 95 
<< m2 >>
rect 194 94 195 95 
<< m1 >>
rect 195 94 196 95 
<< m1 >>
rect 196 94 197 95 
<< m1 >>
rect 197 94 198 95 
<< m1 >>
rect 198 94 199 95 
<< m1 >>
rect 199 94 200 95 
<< m1 >>
rect 200 94 201 95 
<< m1 >>
rect 201 94 202 95 
<< m1 >>
rect 202 94 203 95 
<< m1 >>
rect 203 94 204 95 
<< m1 >>
rect 204 94 205 95 
<< m1 >>
rect 205 94 206 95 
<< m1 >>
rect 206 94 207 95 
<< m1 >>
rect 207 94 208 95 
<< m1 >>
rect 208 94 209 95 
<< m1 >>
rect 209 94 210 95 
<< m1 >>
rect 210 94 211 95 
<< m1 >>
rect 211 94 212 95 
<< m1 >>
rect 212 94 213 95 
<< m1 >>
rect 213 94 214 95 
<< m1 >>
rect 214 94 215 95 
<< m1 >>
rect 215 94 216 95 
<< m1 >>
rect 216 94 217 95 
<< m1 >>
rect 217 94 218 95 
<< m1 >>
rect 218 94 219 95 
<< m1 >>
rect 219 94 220 95 
<< m1 >>
rect 220 94 221 95 
<< m1 >>
rect 221 94 222 95 
<< m1 >>
rect 222 94 223 95 
<< m1 >>
rect 223 94 224 95 
<< m1 >>
rect 224 94 225 95 
<< m2 >>
rect 224 94 225 95 
<< m1 >>
rect 225 94 226 95 
<< m1 >>
rect 226 94 227 95 
<< m2 >>
rect 226 94 227 95 
<< m2c >>
rect 226 94 227 95 
<< m1 >>
rect 226 94 227 95 
<< m2 >>
rect 226 94 227 95 
<< m2 >>
rect 227 94 228 95 
<< m1 >>
rect 228 94 229 95 
<< m2 >>
rect 228 94 229 95 
<< m2 >>
rect 229 94 230 95 
<< m1 >>
rect 230 94 231 95 
<< m2 >>
rect 230 94 231 95 
<< m2c >>
rect 230 94 231 95 
<< m1 >>
rect 230 94 231 95 
<< m2 >>
rect 230 94 231 95 
<< m1 >>
rect 231 94 232 95 
<< m1 >>
rect 232 94 233 95 
<< m1 >>
rect 233 94 234 95 
<< m1 >>
rect 235 94 236 95 
<< m2 >>
rect 241 94 242 95 
<< m1 >>
rect 248 94 249 95 
<< m1 >>
rect 255 94 256 95 
<< m1 >>
rect 257 94 258 95 
<< m1 >>
rect 258 94 259 95 
<< m1 >>
rect 259 94 260 95 
<< m1 >>
rect 260 94 261 95 
<< m1 >>
rect 261 94 262 95 
<< m1 >>
rect 262 94 263 95 
<< m1 >>
rect 263 94 264 95 
<< m1 >>
rect 264 94 265 95 
<< m1 >>
rect 265 94 266 95 
<< m1 >>
rect 266 94 267 95 
<< m1 >>
rect 267 94 268 95 
<< m1 >>
rect 268 94 269 95 
<< m1 >>
rect 269 94 270 95 
<< m1 >>
rect 270 94 271 95 
<< m1 >>
rect 271 94 272 95 
<< m1 >>
rect 272 94 273 95 
<< m1 >>
rect 273 94 274 95 
<< m1 >>
rect 274 94 275 95 
<< m1 >>
rect 275 94 276 95 
<< m1 >>
rect 276 94 277 95 
<< m1 >>
rect 277 94 278 95 
<< m1 >>
rect 278 94 279 95 
<< m1 >>
rect 279 94 280 95 
<< m1 >>
rect 280 94 281 95 
<< m2 >>
rect 280 94 281 95 
<< m1 >>
rect 281 94 282 95 
<< m1 >>
rect 282 94 283 95 
<< m1 >>
rect 283 94 284 95 
<< m1 >>
rect 284 94 285 95 
<< m1 >>
rect 285 94 286 95 
<< m1 >>
rect 286 94 287 95 
<< m1 >>
rect 304 94 305 95 
<< m1 >>
rect 334 94 335 95 
<< m2 >>
rect 344 94 345 95 
<< m1 >>
rect 345 94 346 95 
<< m2 >>
rect 346 94 347 95 
<< m1 >>
rect 347 94 348 95 
<< m2 >>
rect 347 94 348 95 
<< m2c >>
rect 347 94 348 95 
<< m1 >>
rect 347 94 348 95 
<< m2 >>
rect 347 94 348 95 
<< m1 >>
rect 348 94 349 95 
<< m1 >>
rect 349 94 350 95 
<< m1 >>
rect 350 94 351 95 
<< m1 >>
rect 351 94 352 95 
<< m1 >>
rect 352 94 353 95 
<< m1 >>
rect 353 94 354 95 
<< m1 >>
rect 354 94 355 95 
<< m1 >>
rect 355 94 356 95 
<< m1 >>
rect 356 94 357 95 
<< m1 >>
rect 357 94 358 95 
<< m2 >>
rect 357 94 358 95 
<< m1 >>
rect 358 94 359 95 
<< m1 >>
rect 359 94 360 95 
<< m2 >>
rect 359 94 360 95 
<< m2c >>
rect 359 94 360 95 
<< m1 >>
rect 359 94 360 95 
<< m2 >>
rect 359 94 360 95 
<< m2 >>
rect 360 94 361 95 
<< m1 >>
rect 361 94 362 95 
<< m2 >>
rect 361 94 362 95 
<< m2 >>
rect 362 94 363 95 
<< m1 >>
rect 363 94 364 95 
<< m2 >>
rect 363 94 364 95 
<< m2c >>
rect 363 94 364 95 
<< m1 >>
rect 363 94 364 95 
<< m2 >>
rect 363 94 364 95 
<< m1 >>
rect 364 94 365 95 
<< m1 >>
rect 365 94 366 95 
<< m1 >>
rect 366 94 367 95 
<< m2 >>
rect 366 94 367 95 
<< m1 >>
rect 367 94 368 95 
<< m1 >>
rect 368 94 369 95 
<< m2 >>
rect 368 94 369 95 
<< m2c >>
rect 368 94 369 95 
<< m1 >>
rect 368 94 369 95 
<< m2 >>
rect 368 94 369 95 
<< m2 >>
rect 369 94 370 95 
<< m1 >>
rect 370 94 371 95 
<< m2 >>
rect 370 94 371 95 
<< m2 >>
rect 371 94 372 95 
<< m1 >>
rect 372 94 373 95 
<< m2 >>
rect 372 94 373 95 
<< m2c >>
rect 372 94 373 95 
<< m1 >>
rect 372 94 373 95 
<< m2 >>
rect 372 94 373 95 
<< m1 >>
rect 373 94 374 95 
<< m1 >>
rect 374 94 375 95 
<< m1 >>
rect 375 94 376 95 
<< m1 >>
rect 376 94 377 95 
<< m1 >>
rect 377 94 378 95 
<< m1 >>
rect 378 94 379 95 
<< m1 >>
rect 379 94 380 95 
<< m1 >>
rect 380 94 381 95 
<< m1 >>
rect 381 94 382 95 
<< m1 >>
rect 382 94 383 95 
<< m1 >>
rect 383 94 384 95 
<< m1 >>
rect 384 94 385 95 
<< m1 >>
rect 385 94 386 95 
<< m1 >>
rect 386 94 387 95 
<< m1 >>
rect 387 94 388 95 
<< m1 >>
rect 388 94 389 95 
<< m1 >>
rect 389 94 390 95 
<< m1 >>
rect 390 94 391 95 
<< m1 >>
rect 391 94 392 95 
<< m1 >>
rect 392 94 393 95 
<< m2 >>
rect 392 94 393 95 
<< m2c >>
rect 392 94 393 95 
<< m1 >>
rect 392 94 393 95 
<< m2 >>
rect 392 94 393 95 
<< m2 >>
rect 393 94 394 95 
<< m1 >>
rect 394 94 395 95 
<< m2 >>
rect 394 94 395 95 
<< m2 >>
rect 395 94 396 95 
<< m1 >>
rect 396 94 397 95 
<< m2 >>
rect 396 94 397 95 
<< m2c >>
rect 396 94 397 95 
<< m1 >>
rect 396 94 397 95 
<< m2 >>
rect 396 94 397 95 
<< m1 >>
rect 397 94 398 95 
<< m1 >>
rect 398 94 399 95 
<< m1 >>
rect 399 94 400 95 
<< m1 >>
rect 400 94 401 95 
<< m1 >>
rect 401 94 402 95 
<< m1 >>
rect 402 94 403 95 
<< m1 >>
rect 403 94 404 95 
<< m1 >>
rect 404 94 405 95 
<< m1 >>
rect 405 94 406 95 
<< m1 >>
rect 406 94 407 95 
<< m1 >>
rect 407 94 408 95 
<< m1 >>
rect 408 94 409 95 
<< m1 >>
rect 409 94 410 95 
<< m1 >>
rect 410 94 411 95 
<< m1 >>
rect 411 94 412 95 
<< m1 >>
rect 412 94 413 95 
<< m1 >>
rect 413 94 414 95 
<< m1 >>
rect 415 94 416 95 
<< m1 >>
rect 426 94 427 95 
<< m2 >>
rect 426 94 427 95 
<< m1 >>
rect 427 94 428 95 
<< m1 >>
rect 428 94 429 95 
<< m1 >>
rect 429 94 430 95 
<< m1 >>
rect 430 94 431 95 
<< m1 >>
rect 431 94 432 95 
<< m2 >>
rect 431 94 432 95 
<< m2c >>
rect 431 94 432 95 
<< m1 >>
rect 431 94 432 95 
<< m2 >>
rect 431 94 432 95 
<< m2 >>
rect 432 94 433 95 
<< m1 >>
rect 433 94 434 95 
<< m2 >>
rect 433 94 434 95 
<< m1 >>
rect 434 94 435 95 
<< m2 >>
rect 434 94 435 95 
<< m1 >>
rect 435 94 436 95 
<< m2 >>
rect 435 94 436 95 
<< m1 >>
rect 436 94 437 95 
<< m2 >>
rect 436 94 437 95 
<< m1 >>
rect 437 94 438 95 
<< m2 >>
rect 437 94 438 95 
<< m1 >>
rect 438 94 439 95 
<< m2 >>
rect 438 94 439 95 
<< m1 >>
rect 439 94 440 95 
<< m2 >>
rect 439 94 440 95 
<< m1 >>
rect 440 94 441 95 
<< m2 >>
rect 440 94 441 95 
<< m1 >>
rect 441 94 442 95 
<< m2 >>
rect 441 94 442 95 
<< m1 >>
rect 442 94 443 95 
<< m2 >>
rect 442 94 443 95 
<< m1 >>
rect 443 94 444 95 
<< m2 >>
rect 443 94 444 95 
<< m1 >>
rect 444 94 445 95 
<< m2 >>
rect 444 94 445 95 
<< m1 >>
rect 445 94 446 95 
<< m2 >>
rect 445 94 446 95 
<< m1 >>
rect 446 94 447 95 
<< m2 >>
rect 446 94 447 95 
<< m1 >>
rect 447 94 448 95 
<< m2 >>
rect 447 94 448 95 
<< m1 >>
rect 448 94 449 95 
<< m2 >>
rect 448 94 449 95 
<< m2 >>
rect 449 94 450 95 
<< m1 >>
rect 460 94 461 95 
<< m1 >>
rect 462 94 463 95 
<< m1 >>
rect 463 94 464 95 
<< m1 >>
rect 464 94 465 95 
<< m1 >>
rect 466 94 467 95 
<< m1 >>
rect 485 94 486 95 
<< m1 >>
rect 487 94 488 95 
<< m1 >>
rect 49 95 50 96 
<< m1 >>
rect 50 95 51 96 
<< m1 >>
rect 51 95 52 96 
<< m1 >>
rect 52 95 53 96 
<< m1 >>
rect 53 95 54 96 
<< m1 >>
rect 54 95 55 96 
<< m1 >>
rect 55 95 56 96 
<< m1 >>
rect 56 95 57 96 
<< m1 >>
rect 57 95 58 96 
<< m1 >>
rect 58 95 59 96 
<< m1 >>
rect 59 95 60 96 
<< m1 >>
rect 60 95 61 96 
<< m1 >>
rect 61 95 62 96 
<< m1 >>
rect 62 95 63 96 
<< m1 >>
rect 63 95 64 96 
<< m1 >>
rect 64 95 65 96 
<< m2 >>
rect 64 95 65 96 
<< m1 >>
rect 65 95 66 96 
<< m1 >>
rect 66 95 67 96 
<< m1 >>
rect 67 95 68 96 
<< m1 >>
rect 68 95 69 96 
<< m1 >>
rect 69 95 70 96 
<< m1 >>
rect 70 95 71 96 
<< m1 >>
rect 71 95 72 96 
<< m2 >>
rect 71 95 72 96 
<< m2c >>
rect 71 95 72 96 
<< m1 >>
rect 71 95 72 96 
<< m2 >>
rect 71 95 72 96 
<< m2 >>
rect 72 95 73 96 
<< m1 >>
rect 73 95 74 96 
<< m2 >>
rect 73 95 74 96 
<< m2 >>
rect 74 95 75 96 
<< m1 >>
rect 75 95 76 96 
<< m2 >>
rect 75 95 76 96 
<< m2c >>
rect 75 95 76 96 
<< m1 >>
rect 75 95 76 96 
<< m2 >>
rect 75 95 76 96 
<< m1 >>
rect 76 95 77 96 
<< m1 >>
rect 77 95 78 96 
<< m1 >>
rect 78 95 79 96 
<< m1 >>
rect 79 95 80 96 
<< m1 >>
rect 80 95 81 96 
<< m1 >>
rect 81 95 82 96 
<< m1 >>
rect 82 95 83 96 
<< m1 >>
rect 83 95 84 96 
<< m1 >>
rect 84 95 85 96 
<< m1 >>
rect 85 95 86 96 
<< m1 >>
rect 86 95 87 96 
<< m2 >>
rect 86 95 87 96 
<< m2c >>
rect 86 95 87 96 
<< m1 >>
rect 86 95 87 96 
<< m2 >>
rect 86 95 87 96 
<< m2 >>
rect 87 95 88 96 
<< m1 >>
rect 88 95 89 96 
<< m2 >>
rect 88 95 89 96 
<< m2 >>
rect 89 95 90 96 
<< m1 >>
rect 92 95 93 96 
<< m1 >>
rect 100 95 101 96 
<< m2 >>
rect 100 95 101 96 
<< m1 >>
rect 127 95 128 96 
<< m1 >>
rect 129 95 130 96 
<< m1 >>
rect 131 95 132 96 
<< m1 >>
rect 145 95 146 96 
<< m1 >>
rect 149 95 150 96 
<< m2 >>
rect 149 95 150 96 
<< m2c >>
rect 149 95 150 96 
<< m1 >>
rect 149 95 150 96 
<< m2 >>
rect 149 95 150 96 
<< m2 >>
rect 174 95 175 96 
<< m1 >>
rect 187 95 188 96 
<< m2 >>
rect 189 95 190 96 
<< m1 >>
rect 190 95 191 96 
<< m2 >>
rect 190 95 191 96 
<< m2 >>
rect 191 95 192 96 
<< m2 >>
rect 192 95 193 96 
<< m2 >>
rect 193 95 194 96 
<< m2 >>
rect 194 95 195 96 
<< m2 >>
rect 224 95 225 96 
<< m1 >>
rect 228 95 229 96 
<< m1 >>
rect 235 95 236 96 
<< m1 >>
rect 239 95 240 96 
<< m2 >>
rect 239 95 240 96 
<< m2c >>
rect 239 95 240 96 
<< m1 >>
rect 239 95 240 96 
<< m2 >>
rect 239 95 240 96 
<< m1 >>
rect 240 95 241 96 
<< m1 >>
rect 241 95 242 96 
<< m2 >>
rect 241 95 242 96 
<< m1 >>
rect 242 95 243 96 
<< m1 >>
rect 243 95 244 96 
<< m1 >>
rect 244 95 245 96 
<< m1 >>
rect 245 95 246 96 
<< m1 >>
rect 246 95 247 96 
<< m1 >>
rect 247 95 248 96 
<< m1 >>
rect 248 95 249 96 
<< m1 >>
rect 255 95 256 96 
<< m2 >>
rect 255 95 256 96 
<< m2c >>
rect 255 95 256 96 
<< m1 >>
rect 255 95 256 96 
<< m2 >>
rect 255 95 256 96 
<< m2 >>
rect 280 95 281 96 
<< m1 >>
rect 304 95 305 96 
<< m1 >>
rect 334 95 335 96 
<< m2 >>
rect 344 95 345 96 
<< m1 >>
rect 345 95 346 96 
<< m2 >>
rect 346 95 347 96 
<< m2 >>
rect 357 95 358 96 
<< m1 >>
rect 361 95 362 96 
<< m2 >>
rect 366 95 367 96 
<< m1 >>
rect 370 95 371 96 
<< m1 >>
rect 394 95 395 96 
<< m1 >>
rect 415 95 416 96 
<< m2 >>
rect 415 95 416 96 
<< m2c >>
rect 415 95 416 96 
<< m1 >>
rect 415 95 416 96 
<< m2 >>
rect 415 95 416 96 
<< m2 >>
rect 426 95 427 96 
<< m1 >>
rect 460 95 461 96 
<< m2 >>
rect 460 95 461 96 
<< m2c >>
rect 460 95 461 96 
<< m1 >>
rect 460 95 461 96 
<< m2 >>
rect 460 95 461 96 
<< m1 >>
rect 466 95 467 96 
<< m2 >>
rect 466 95 467 96 
<< m2c >>
rect 466 95 467 96 
<< m1 >>
rect 466 95 467 96 
<< m2 >>
rect 466 95 467 96 
<< m1 >>
rect 485 95 486 96 
<< m2 >>
rect 485 95 486 96 
<< m2c >>
rect 485 95 486 96 
<< m1 >>
rect 485 95 486 96 
<< m2 >>
rect 485 95 486 96 
<< m1 >>
rect 487 95 488 96 
<< m2 >>
rect 487 95 488 96 
<< m2c >>
rect 487 95 488 96 
<< m1 >>
rect 487 95 488 96 
<< m2 >>
rect 487 95 488 96 
<< m2 >>
rect 64 96 65 97 
<< m1 >>
rect 73 96 74 97 
<< m1 >>
rect 88 96 89 97 
<< m2 >>
rect 89 96 90 97 
<< m1 >>
rect 92 96 93 97 
<< m2 >>
rect 92 96 93 97 
<< m2c >>
rect 92 96 93 97 
<< m1 >>
rect 92 96 93 97 
<< m2 >>
rect 92 96 93 97 
<< m1 >>
rect 100 96 101 97 
<< m2 >>
rect 100 96 101 97 
<< m1 >>
rect 127 96 128 97 
<< m1 >>
rect 129 96 130 97 
<< m1 >>
rect 131 96 132 97 
<< m1 >>
rect 145 96 146 97 
<< m2 >>
rect 149 96 150 97 
<< m2 >>
rect 150 96 151 97 
<< m2 >>
rect 151 96 152 97 
<< m2 >>
rect 152 96 153 97 
<< m2 >>
rect 153 96 154 97 
<< m2 >>
rect 154 96 155 97 
<< m2 >>
rect 155 96 156 97 
<< m2 >>
rect 156 96 157 97 
<< m2 >>
rect 157 96 158 97 
<< m2 >>
rect 158 96 159 97 
<< m2 >>
rect 174 96 175 97 
<< m1 >>
rect 187 96 188 97 
<< m2 >>
rect 189 96 190 97 
<< m1 >>
rect 190 96 191 97 
<< m1 >>
rect 224 96 225 97 
<< m2 >>
rect 224 96 225 97 
<< m2c >>
rect 224 96 225 97 
<< m1 >>
rect 224 96 225 97 
<< m2 >>
rect 224 96 225 97 
<< m1 >>
rect 228 96 229 97 
<< m1 >>
rect 235 96 236 97 
<< m2 >>
rect 239 96 240 97 
<< m2 >>
rect 241 96 242 97 
<< m2 >>
rect 255 96 256 97 
<< m1 >>
rect 280 96 281 97 
<< m2 >>
rect 280 96 281 97 
<< m2c >>
rect 280 96 281 97 
<< m1 >>
rect 280 96 281 97 
<< m2 >>
rect 280 96 281 97 
<< m1 >>
rect 304 96 305 97 
<< m1 >>
rect 334 96 335 97 
<< m2 >>
rect 344 96 345 97 
<< m1 >>
rect 345 96 346 97 
<< m2 >>
rect 346 96 347 97 
<< m1 >>
rect 352 96 353 97 
<< m1 >>
rect 353 96 354 97 
<< m1 >>
rect 354 96 355 97 
<< m1 >>
rect 355 96 356 97 
<< m1 >>
rect 356 96 357 97 
<< m1 >>
rect 357 96 358 97 
<< m2 >>
rect 357 96 358 97 
<< m2c >>
rect 357 96 358 97 
<< m1 >>
rect 357 96 358 97 
<< m2 >>
rect 357 96 358 97 
<< m1 >>
rect 361 96 362 97 
<< m1 >>
rect 366 96 367 97 
<< m2 >>
rect 366 96 367 97 
<< m2c >>
rect 366 96 367 97 
<< m1 >>
rect 366 96 367 97 
<< m2 >>
rect 366 96 367 97 
<< m1 >>
rect 370 96 371 97 
<< m2 >>
rect 390 96 391 97 
<< m2 >>
rect 391 96 392 97 
<< m2 >>
rect 392 96 393 97 
<< m2 >>
rect 393 96 394 97 
<< m1 >>
rect 394 96 395 97 
<< m2 >>
rect 394 96 395 97 
<< m2 >>
rect 395 96 396 97 
<< m2 >>
rect 396 96 397 97 
<< m2 >>
rect 397 96 398 97 
<< m2 >>
rect 398 96 399 97 
<< m2 >>
rect 399 96 400 97 
<< m2 >>
rect 400 96 401 97 
<< m2 >>
rect 401 96 402 97 
<< m2 >>
rect 402 96 403 97 
<< m2 >>
rect 403 96 404 97 
<< m2 >>
rect 404 96 405 97 
<< m2 >>
rect 405 96 406 97 
<< m2 >>
rect 406 96 407 97 
<< m2 >>
rect 407 96 408 97 
<< m2 >>
rect 408 96 409 97 
<< m2 >>
rect 409 96 410 97 
<< m2 >>
rect 410 96 411 97 
<< m2 >>
rect 411 96 412 97 
<< m2 >>
rect 412 96 413 97 
<< m2 >>
rect 413 96 414 97 
<< m2 >>
rect 414 96 415 97 
<< m2 >>
rect 415 96 416 97 
<< m2 >>
rect 426 96 427 97 
<< m2 >>
rect 460 96 461 97 
<< m2 >>
rect 466 96 467 97 
<< m2 >>
rect 480 96 481 97 
<< m2 >>
rect 481 96 482 97 
<< m2 >>
rect 482 96 483 97 
<< m2 >>
rect 483 96 484 97 
<< m2 >>
rect 484 96 485 97 
<< m2 >>
rect 485 96 486 97 
<< m2 >>
rect 487 96 488 97 
<< m1 >>
rect 46 97 47 98 
<< m1 >>
rect 47 97 48 98 
<< m2 >>
rect 47 97 48 98 
<< m2c >>
rect 47 97 48 98 
<< m1 >>
rect 47 97 48 98 
<< m2 >>
rect 47 97 48 98 
<< m2 >>
rect 48 97 49 98 
<< m1 >>
rect 49 97 50 98 
<< m2 >>
rect 49 97 50 98 
<< m1 >>
rect 50 97 51 98 
<< m2 >>
rect 50 97 51 98 
<< m1 >>
rect 51 97 52 98 
<< m2 >>
rect 51 97 52 98 
<< m1 >>
rect 52 97 53 98 
<< m2 >>
rect 52 97 53 98 
<< m1 >>
rect 53 97 54 98 
<< m1 >>
rect 54 97 55 98 
<< m1 >>
rect 55 97 56 98 
<< m1 >>
rect 56 97 57 98 
<< m1 >>
rect 57 97 58 98 
<< m1 >>
rect 58 97 59 98 
<< m1 >>
rect 59 97 60 98 
<< m1 >>
rect 60 97 61 98 
<< m1 >>
rect 61 97 62 98 
<< m1 >>
rect 62 97 63 98 
<< m1 >>
rect 63 97 64 98 
<< m1 >>
rect 64 97 65 98 
<< m2 >>
rect 64 97 65 98 
<< m1 >>
rect 65 97 66 98 
<< m1 >>
rect 66 97 67 98 
<< m1 >>
rect 67 97 68 98 
<< m1 >>
rect 68 97 69 98 
<< m1 >>
rect 69 97 70 98 
<< m1 >>
rect 70 97 71 98 
<< m1 >>
rect 71 97 72 98 
<< m2 >>
rect 71 97 72 98 
<< m2c >>
rect 71 97 72 98 
<< m1 >>
rect 71 97 72 98 
<< m2 >>
rect 71 97 72 98 
<< m2 >>
rect 72 97 73 98 
<< m1 >>
rect 73 97 74 98 
<< m2 >>
rect 73 97 74 98 
<< m2 >>
rect 74 97 75 98 
<< m1 >>
rect 75 97 76 98 
<< m2 >>
rect 75 97 76 98 
<< m2c >>
rect 75 97 76 98 
<< m1 >>
rect 75 97 76 98 
<< m2 >>
rect 75 97 76 98 
<< m1 >>
rect 76 97 77 98 
<< m1 >>
rect 77 97 78 98 
<< m1 >>
rect 78 97 79 98 
<< m1 >>
rect 79 97 80 98 
<< m1 >>
rect 80 97 81 98 
<< m1 >>
rect 81 97 82 98 
<< m1 >>
rect 82 97 83 98 
<< m1 >>
rect 83 97 84 98 
<< m1 >>
rect 84 97 85 98 
<< m1 >>
rect 85 97 86 98 
<< m1 >>
rect 86 97 87 98 
<< m1 >>
rect 87 97 88 98 
<< m1 >>
rect 88 97 89 98 
<< m2 >>
rect 89 97 90 98 
<< m2 >>
rect 92 97 93 98 
<< m1 >>
rect 100 97 101 98 
<< m2 >>
rect 100 97 101 98 
<< m1 >>
rect 127 97 128 98 
<< m1 >>
rect 129 97 130 98 
<< m1 >>
rect 131 97 132 98 
<< m1 >>
rect 138 97 139 98 
<< m1 >>
rect 139 97 140 98 
<< m1 >>
rect 140 97 141 98 
<< m1 >>
rect 141 97 142 98 
<< m1 >>
rect 142 97 143 98 
<< m1 >>
rect 143 97 144 98 
<< m2 >>
rect 143 97 144 98 
<< m2c >>
rect 143 97 144 98 
<< m1 >>
rect 143 97 144 98 
<< m2 >>
rect 143 97 144 98 
<< m2 >>
rect 144 97 145 98 
<< m1 >>
rect 145 97 146 98 
<< m2 >>
rect 145 97 146 98 
<< m2 >>
rect 146 97 147 98 
<< m1 >>
rect 147 97 148 98 
<< m2 >>
rect 147 97 148 98 
<< m2c >>
rect 147 97 148 98 
<< m1 >>
rect 147 97 148 98 
<< m2 >>
rect 147 97 148 98 
<< m1 >>
rect 148 97 149 98 
<< m1 >>
rect 149 97 150 98 
<< m1 >>
rect 150 97 151 98 
<< m1 >>
rect 151 97 152 98 
<< m1 >>
rect 152 97 153 98 
<< m1 >>
rect 153 97 154 98 
<< m1 >>
rect 154 97 155 98 
<< m1 >>
rect 155 97 156 98 
<< m1 >>
rect 156 97 157 98 
<< m1 >>
rect 157 97 158 98 
<< m1 >>
rect 158 97 159 98 
<< m2 >>
rect 158 97 159 98 
<< m1 >>
rect 159 97 160 98 
<< m1 >>
rect 160 97 161 98 
<< m1 >>
rect 161 97 162 98 
<< m1 >>
rect 162 97 163 98 
<< m1 >>
rect 163 97 164 98 
<< m1 >>
rect 164 97 165 98 
<< m1 >>
rect 165 97 166 98 
<< m1 >>
rect 166 97 167 98 
<< m1 >>
rect 167 97 168 98 
<< m1 >>
rect 168 97 169 98 
<< m1 >>
rect 169 97 170 98 
<< m1 >>
rect 170 97 171 98 
<< m1 >>
rect 171 97 172 98 
<< m1 >>
rect 172 97 173 98 
<< m1 >>
rect 173 97 174 98 
<< m1 >>
rect 174 97 175 98 
<< m2 >>
rect 174 97 175 98 
<< m1 >>
rect 175 97 176 98 
<< m1 >>
rect 176 97 177 98 
<< m1 >>
rect 177 97 178 98 
<< m1 >>
rect 178 97 179 98 
<< m1 >>
rect 187 97 188 98 
<< m2 >>
rect 189 97 190 98 
<< m1 >>
rect 190 97 191 98 
<< m1 >>
rect 224 97 225 98 
<< m1 >>
rect 228 97 229 98 
<< m1 >>
rect 229 97 230 98 
<< m1 >>
rect 230 97 231 98 
<< m1 >>
rect 231 97 232 98 
<< m1 >>
rect 232 97 233 98 
<< m1 >>
rect 233 97 234 98 
<< m2 >>
rect 233 97 234 98 
<< m2c >>
rect 233 97 234 98 
<< m1 >>
rect 233 97 234 98 
<< m2 >>
rect 233 97 234 98 
<< m2 >>
rect 234 97 235 98 
<< m1 >>
rect 235 97 236 98 
<< m2 >>
rect 235 97 236 98 
<< m2 >>
rect 236 97 237 98 
<< m1 >>
rect 237 97 238 98 
<< m2 >>
rect 237 97 238 98 
<< m2c >>
rect 237 97 238 98 
<< m1 >>
rect 237 97 238 98 
<< m2 >>
rect 237 97 238 98 
<< m1 >>
rect 238 97 239 98 
<< m1 >>
rect 239 97 240 98 
<< m2 >>
rect 239 97 240 98 
<< m1 >>
rect 240 97 241 98 
<< m1 >>
rect 241 97 242 98 
<< m2 >>
rect 241 97 242 98 
<< m1 >>
rect 242 97 243 98 
<< m1 >>
rect 243 97 244 98 
<< m1 >>
rect 244 97 245 98 
<< m1 >>
rect 245 97 246 98 
<< m1 >>
rect 246 97 247 98 
<< m1 >>
rect 247 97 248 98 
<< m1 >>
rect 248 97 249 98 
<< m1 >>
rect 249 97 250 98 
<< m1 >>
rect 250 97 251 98 
<< m1 >>
rect 251 97 252 98 
<< m1 >>
rect 252 97 253 98 
<< m1 >>
rect 253 97 254 98 
<< m1 >>
rect 254 97 255 98 
<< m1 >>
rect 255 97 256 98 
<< m2 >>
rect 255 97 256 98 
<< m1 >>
rect 256 97 257 98 
<< m1 >>
rect 257 97 258 98 
<< m1 >>
rect 258 97 259 98 
<< m1 >>
rect 259 97 260 98 
<< m1 >>
rect 260 97 261 98 
<< m1 >>
rect 261 97 262 98 
<< m1 >>
rect 262 97 263 98 
<< m1 >>
rect 263 97 264 98 
<< m1 >>
rect 264 97 265 98 
<< m1 >>
rect 265 97 266 98 
<< m1 >>
rect 280 97 281 98 
<< m1 >>
rect 283 97 284 98 
<< m1 >>
rect 284 97 285 98 
<< m1 >>
rect 285 97 286 98 
<< m1 >>
rect 286 97 287 98 
<< m1 >>
rect 287 97 288 98 
<< m1 >>
rect 288 97 289 98 
<< m1 >>
rect 289 97 290 98 
<< m1 >>
rect 290 97 291 98 
<< m1 >>
rect 291 97 292 98 
<< m1 >>
rect 292 97 293 98 
<< m1 >>
rect 293 97 294 98 
<< m1 >>
rect 294 97 295 98 
<< m1 >>
rect 295 97 296 98 
<< m1 >>
rect 296 97 297 98 
<< m1 >>
rect 297 97 298 98 
<< m1 >>
rect 298 97 299 98 
<< m1 >>
rect 299 97 300 98 
<< m1 >>
rect 300 97 301 98 
<< m1 >>
rect 301 97 302 98 
<< m1 >>
rect 302 97 303 98 
<< m1 >>
rect 303 97 304 98 
<< m1 >>
rect 304 97 305 98 
<< m1 >>
rect 307 97 308 98 
<< m1 >>
rect 308 97 309 98 
<< m1 >>
rect 309 97 310 98 
<< m1 >>
rect 310 97 311 98 
<< m1 >>
rect 311 97 312 98 
<< m1 >>
rect 312 97 313 98 
<< m1 >>
rect 313 97 314 98 
<< m1 >>
rect 314 97 315 98 
<< m1 >>
rect 315 97 316 98 
<< m1 >>
rect 316 97 317 98 
<< m1 >>
rect 317 97 318 98 
<< m1 >>
rect 318 97 319 98 
<< m1 >>
rect 319 97 320 98 
<< m1 >>
rect 320 97 321 98 
<< m1 >>
rect 321 97 322 98 
<< m1 >>
rect 322 97 323 98 
<< m1 >>
rect 323 97 324 98 
<< m1 >>
rect 324 97 325 98 
<< m1 >>
rect 325 97 326 98 
<< m1 >>
rect 326 97 327 98 
<< m1 >>
rect 327 97 328 98 
<< m1 >>
rect 328 97 329 98 
<< m1 >>
rect 329 97 330 98 
<< m1 >>
rect 330 97 331 98 
<< m1 >>
rect 331 97 332 98 
<< m1 >>
rect 332 97 333 98 
<< m2 >>
rect 332 97 333 98 
<< m2c >>
rect 332 97 333 98 
<< m1 >>
rect 332 97 333 98 
<< m2 >>
rect 332 97 333 98 
<< m2 >>
rect 333 97 334 98 
<< m1 >>
rect 334 97 335 98 
<< m2 >>
rect 334 97 335 98 
<< m2 >>
rect 335 97 336 98 
<< m1 >>
rect 336 97 337 98 
<< m2 >>
rect 336 97 337 98 
<< m2c >>
rect 336 97 337 98 
<< m1 >>
rect 336 97 337 98 
<< m2 >>
rect 336 97 337 98 
<< m1 >>
rect 337 97 338 98 
<< m1 >>
rect 338 97 339 98 
<< m1 >>
rect 339 97 340 98 
<< m1 >>
rect 340 97 341 98 
<< m1 >>
rect 341 97 342 98 
<< m1 >>
rect 342 97 343 98 
<< m1 >>
rect 343 97 344 98 
<< m2 >>
rect 343 97 344 98 
<< m2c >>
rect 343 97 344 98 
<< m1 >>
rect 343 97 344 98 
<< m2 >>
rect 343 97 344 98 
<< m2 >>
rect 344 97 345 98 
<< m1 >>
rect 345 97 346 98 
<< m2 >>
rect 346 97 347 98 
<< m1 >>
rect 352 97 353 98 
<< m1 >>
rect 361 97 362 98 
<< m1 >>
rect 366 97 367 98 
<< m2 >>
rect 369 97 370 98 
<< m1 >>
rect 370 97 371 98 
<< m2 >>
rect 370 97 371 98 
<< m2 >>
rect 371 97 372 98 
<< m2 >>
rect 372 97 373 98 
<< m1 >>
rect 373 97 374 98 
<< m2 >>
rect 373 97 374 98 
<< m1 >>
rect 374 97 375 98 
<< m2 >>
rect 374 97 375 98 
<< m1 >>
rect 375 97 376 98 
<< m1 >>
rect 376 97 377 98 
<< m1 >>
rect 377 97 378 98 
<< m1 >>
rect 378 97 379 98 
<< m1 >>
rect 379 97 380 98 
<< m1 >>
rect 380 97 381 98 
<< m1 >>
rect 381 97 382 98 
<< m1 >>
rect 382 97 383 98 
<< m1 >>
rect 383 97 384 98 
<< m1 >>
rect 384 97 385 98 
<< m1 >>
rect 385 97 386 98 
<< m1 >>
rect 386 97 387 98 
<< m1 >>
rect 387 97 388 98 
<< m1 >>
rect 388 97 389 98 
<< m1 >>
rect 389 97 390 98 
<< m1 >>
rect 390 97 391 98 
<< m2 >>
rect 390 97 391 98 
<< m1 >>
rect 391 97 392 98 
<< m1 >>
rect 392 97 393 98 
<< m1 >>
rect 393 97 394 98 
<< m1 >>
rect 394 97 395 98 
<< m1 >>
rect 397 97 398 98 
<< m1 >>
rect 398 97 399 98 
<< m1 >>
rect 399 97 400 98 
<< m1 >>
rect 400 97 401 98 
<< m1 >>
rect 401 97 402 98 
<< m1 >>
rect 402 97 403 98 
<< m1 >>
rect 403 97 404 98 
<< m1 >>
rect 404 97 405 98 
<< m1 >>
rect 405 97 406 98 
<< m1 >>
rect 406 97 407 98 
<< m1 >>
rect 407 97 408 98 
<< m1 >>
rect 408 97 409 98 
<< m1 >>
rect 409 97 410 98 
<< m1 >>
rect 410 97 411 98 
<< m1 >>
rect 411 97 412 98 
<< m1 >>
rect 412 97 413 98 
<< m1 >>
rect 413 97 414 98 
<< m1 >>
rect 414 97 415 98 
<< m1 >>
rect 415 97 416 98 
<< m1 >>
rect 416 97 417 98 
<< m1 >>
rect 417 97 418 98 
<< m1 >>
rect 418 97 419 98 
<< m1 >>
rect 419 97 420 98 
<< m1 >>
rect 420 97 421 98 
<< m1 >>
rect 421 97 422 98 
<< m1 >>
rect 422 97 423 98 
<< m1 >>
rect 423 97 424 98 
<< m1 >>
rect 424 97 425 98 
<< m1 >>
rect 425 97 426 98 
<< m1 >>
rect 426 97 427 98 
<< m2 >>
rect 426 97 427 98 
<< m1 >>
rect 427 97 428 98 
<< m2 >>
rect 427 97 428 98 
<< m1 >>
rect 428 97 429 98 
<< m2 >>
rect 428 97 429 98 
<< m1 >>
rect 429 97 430 98 
<< m2 >>
rect 429 97 430 98 
<< m1 >>
rect 430 97 431 98 
<< m2 >>
rect 430 97 431 98 
<< m1 >>
rect 431 97 432 98 
<< m2 >>
rect 431 97 432 98 
<< m1 >>
rect 432 97 433 98 
<< m2 >>
rect 432 97 433 98 
<< m1 >>
rect 433 97 434 98 
<< m2 >>
rect 433 97 434 98 
<< m1 >>
rect 434 97 435 98 
<< m2 >>
rect 434 97 435 98 
<< m1 >>
rect 435 97 436 98 
<< m2 >>
rect 435 97 436 98 
<< m1 >>
rect 436 97 437 98 
<< m2 >>
rect 436 97 437 98 
<< m1 >>
rect 437 97 438 98 
<< m2 >>
rect 437 97 438 98 
<< m1 >>
rect 438 97 439 98 
<< m2 >>
rect 438 97 439 98 
<< m1 >>
rect 439 97 440 98 
<< m2 >>
rect 439 97 440 98 
<< m1 >>
rect 440 97 441 98 
<< m2 >>
rect 440 97 441 98 
<< m1 >>
rect 441 97 442 98 
<< m2 >>
rect 441 97 442 98 
<< m1 >>
rect 442 97 443 98 
<< m2 >>
rect 442 97 443 98 
<< m1 >>
rect 443 97 444 98 
<< m2 >>
rect 443 97 444 98 
<< m1 >>
rect 444 97 445 98 
<< m2 >>
rect 444 97 445 98 
<< m1 >>
rect 445 97 446 98 
<< m2 >>
rect 445 97 446 98 
<< m1 >>
rect 446 97 447 98 
<< m2 >>
rect 446 97 447 98 
<< m1 >>
rect 447 97 448 98 
<< m2 >>
rect 447 97 448 98 
<< m1 >>
rect 448 97 449 98 
<< m2 >>
rect 448 97 449 98 
<< m1 >>
rect 449 97 450 98 
<< m2 >>
rect 449 97 450 98 
<< m1 >>
rect 450 97 451 98 
<< m2 >>
rect 450 97 451 98 
<< m1 >>
rect 451 97 452 98 
<< m2 >>
rect 451 97 452 98 
<< m1 >>
rect 452 97 453 98 
<< m2 >>
rect 452 97 453 98 
<< m1 >>
rect 453 97 454 98 
<< m2 >>
rect 453 97 454 98 
<< m1 >>
rect 454 97 455 98 
<< m2 >>
rect 454 97 455 98 
<< m1 >>
rect 455 97 456 98 
<< m2 >>
rect 455 97 456 98 
<< m1 >>
rect 456 97 457 98 
<< m2 >>
rect 456 97 457 98 
<< m1 >>
rect 457 97 458 98 
<< m1 >>
rect 458 97 459 98 
<< m1 >>
rect 459 97 460 98 
<< m1 >>
rect 460 97 461 98 
<< m2 >>
rect 460 97 461 98 
<< m1 >>
rect 461 97 462 98 
<< m1 >>
rect 462 97 463 98 
<< m1 >>
rect 463 97 464 98 
<< m1 >>
rect 464 97 465 98 
<< m1 >>
rect 465 97 466 98 
<< m1 >>
rect 466 97 467 98 
<< m2 >>
rect 466 97 467 98 
<< m1 >>
rect 467 97 468 98 
<< m1 >>
rect 468 97 469 98 
<< m1 >>
rect 469 97 470 98 
<< m1 >>
rect 470 97 471 98 
<< m1 >>
rect 471 97 472 98 
<< m1 >>
rect 472 97 473 98 
<< m1 >>
rect 473 97 474 98 
<< m1 >>
rect 474 97 475 98 
<< m1 >>
rect 475 97 476 98 
<< m1 >>
rect 476 97 477 98 
<< m1 >>
rect 477 97 478 98 
<< m1 >>
rect 478 97 479 98 
<< m1 >>
rect 479 97 480 98 
<< m1 >>
rect 480 97 481 98 
<< m2 >>
rect 480 97 481 98 
<< m1 >>
rect 481 97 482 98 
<< m1 >>
rect 482 97 483 98 
<< m1 >>
rect 483 97 484 98 
<< m1 >>
rect 484 97 485 98 
<< m1 >>
rect 485 97 486 98 
<< m1 >>
rect 486 97 487 98 
<< m1 >>
rect 487 97 488 98 
<< m2 >>
rect 487 97 488 98 
<< m1 >>
rect 488 97 489 98 
<< m1 >>
rect 489 97 490 98 
<< m1 >>
rect 490 97 491 98 
<< m1 >>
rect 491 97 492 98 
<< m1 >>
rect 492 97 493 98 
<< m1 >>
rect 493 97 494 98 
<< m1 >>
rect 494 97 495 98 
<< m1 >>
rect 495 97 496 98 
<< m1 >>
rect 496 97 497 98 
<< m1 >>
rect 497 97 498 98 
<< m1 >>
rect 498 97 499 98 
<< m1 >>
rect 499 97 500 98 
<< m1 >>
rect 500 97 501 98 
<< m1 >>
rect 501 97 502 98 
<< m1 >>
rect 502 97 503 98 
<< m1 >>
rect 46 98 47 99 
<< m1 >>
rect 49 98 50 99 
<< m2 >>
rect 52 98 53 99 
<< m2 >>
rect 64 98 65 99 
<< m1 >>
rect 73 98 74 99 
<< m2 >>
rect 89 98 90 99 
<< m1 >>
rect 90 98 91 99 
<< m2 >>
rect 90 98 91 99 
<< m2c >>
rect 90 98 91 99 
<< m1 >>
rect 90 98 91 99 
<< m2 >>
rect 90 98 91 99 
<< m1 >>
rect 91 98 92 99 
<< m1 >>
rect 92 98 93 99 
<< m2 >>
rect 92 98 93 99 
<< m1 >>
rect 93 98 94 99 
<< m1 >>
rect 94 98 95 99 
<< m1 >>
rect 95 98 96 99 
<< m1 >>
rect 96 98 97 99 
<< m1 >>
rect 97 98 98 99 
<< m1 >>
rect 98 98 99 99 
<< m1 >>
rect 100 98 101 99 
<< m2 >>
rect 100 98 101 99 
<< m1 >>
rect 127 98 128 99 
<< m1 >>
rect 129 98 130 99 
<< m1 >>
rect 131 98 132 99 
<< m1 >>
rect 138 98 139 99 
<< m2 >>
rect 138 98 139 99 
<< m2c >>
rect 138 98 139 99 
<< m1 >>
rect 138 98 139 99 
<< m2 >>
rect 138 98 139 99 
<< m1 >>
rect 145 98 146 99 
<< m2 >>
rect 158 98 159 99 
<< m2 >>
rect 174 98 175 99 
<< m1 >>
rect 178 98 179 99 
<< m1 >>
rect 187 98 188 99 
<< m2 >>
rect 189 98 190 99 
<< m1 >>
rect 190 98 191 99 
<< m1 >>
rect 224 98 225 99 
<< m1 >>
rect 235 98 236 99 
<< m2 >>
rect 239 98 240 99 
<< m2 >>
rect 241 98 242 99 
<< m2 >>
rect 255 98 256 99 
<< m1 >>
rect 265 98 266 99 
<< m1 >>
rect 280 98 281 99 
<< m1 >>
rect 283 98 284 99 
<< m1 >>
rect 307 98 308 99 
<< m1 >>
rect 334 98 335 99 
<< m1 >>
rect 345 98 346 99 
<< m2 >>
rect 346 98 347 99 
<< m1 >>
rect 352 98 353 99 
<< m1 >>
rect 361 98 362 99 
<< m1 >>
rect 366 98 367 99 
<< m2 >>
rect 369 98 370 99 
<< m1 >>
rect 370 98 371 99 
<< m1 >>
rect 373 98 374 99 
<< m2 >>
rect 374 98 375 99 
<< m2 >>
rect 390 98 391 99 
<< m1 >>
rect 397 98 398 99 
<< m2 >>
rect 456 98 457 99 
<< m2 >>
rect 460 98 461 99 
<< m2 >>
rect 466 98 467 99 
<< m2 >>
rect 480 98 481 99 
<< m2 >>
rect 487 98 488 99 
<< m1 >>
rect 502 98 503 99 
<< m1 >>
rect 46 99 47 100 
<< m1 >>
rect 49 99 50 100 
<< m1 >>
rect 52 99 53 100 
<< m2 >>
rect 52 99 53 100 
<< m2c >>
rect 52 99 53 100 
<< m1 >>
rect 52 99 53 100 
<< m2 >>
rect 52 99 53 100 
<< m1 >>
rect 64 99 65 100 
<< m2 >>
rect 64 99 65 100 
<< m2c >>
rect 64 99 65 100 
<< m1 >>
rect 64 99 65 100 
<< m2 >>
rect 64 99 65 100 
<< m1 >>
rect 73 99 74 100 
<< m2 >>
rect 92 99 93 100 
<< m1 >>
rect 98 99 99 100 
<< m1 >>
rect 100 99 101 100 
<< m2 >>
rect 100 99 101 100 
<< m1 >>
rect 127 99 128 100 
<< m1 >>
rect 129 99 130 100 
<< m1 >>
rect 131 99 132 100 
<< m2 >>
rect 136 99 137 100 
<< m2 >>
rect 137 99 138 100 
<< m2 >>
rect 138 99 139 100 
<< m1 >>
rect 145 99 146 100 
<< m2 >>
rect 158 99 159 100 
<< m2 >>
rect 159 99 160 100 
<< m2 >>
rect 160 99 161 100 
<< m2 >>
rect 161 99 162 100 
<< m2 >>
rect 162 99 163 100 
<< m2 >>
rect 163 99 164 100 
<< m2 >>
rect 164 99 165 100 
<< m1 >>
rect 165 99 166 100 
<< m2 >>
rect 165 99 166 100 
<< m2c >>
rect 165 99 166 100 
<< m1 >>
rect 165 99 166 100 
<< m2 >>
rect 165 99 166 100 
<< m1 >>
rect 172 99 173 100 
<< m1 >>
rect 173 99 174 100 
<< m1 >>
rect 174 99 175 100 
<< m2 >>
rect 174 99 175 100 
<< m2c >>
rect 174 99 175 100 
<< m1 >>
rect 174 99 175 100 
<< m2 >>
rect 174 99 175 100 
<< m1 >>
rect 178 99 179 100 
<< m1 >>
rect 187 99 188 100 
<< m2 >>
rect 189 99 190 100 
<< m1 >>
rect 190 99 191 100 
<< m1 >>
rect 224 99 225 100 
<< m1 >>
rect 229 99 230 100 
<< m1 >>
rect 230 99 231 100 
<< m1 >>
rect 231 99 232 100 
<< m1 >>
rect 232 99 233 100 
<< m1 >>
rect 233 99 234 100 
<< m2 >>
rect 233 99 234 100 
<< m2c >>
rect 233 99 234 100 
<< m1 >>
rect 233 99 234 100 
<< m2 >>
rect 233 99 234 100 
<< m2 >>
rect 234 99 235 100 
<< m1 >>
rect 235 99 236 100 
<< m2 >>
rect 235 99 236 100 
<< m2 >>
rect 236 99 237 100 
<< m1 >>
rect 237 99 238 100 
<< m2 >>
rect 237 99 238 100 
<< m2c >>
rect 237 99 238 100 
<< m1 >>
rect 237 99 238 100 
<< m2 >>
rect 237 99 238 100 
<< m1 >>
rect 238 99 239 100 
<< m1 >>
rect 239 99 240 100 
<< m2 >>
rect 239 99 240 100 
<< m2c >>
rect 239 99 240 100 
<< m1 >>
rect 239 99 240 100 
<< m2 >>
rect 239 99 240 100 
<< m1 >>
rect 241 99 242 100 
<< m2 >>
rect 241 99 242 100 
<< m2c >>
rect 241 99 242 100 
<< m1 >>
rect 241 99 242 100 
<< m2 >>
rect 241 99 242 100 
<< m1 >>
rect 255 99 256 100 
<< m2 >>
rect 255 99 256 100 
<< m2c >>
rect 255 99 256 100 
<< m1 >>
rect 255 99 256 100 
<< m2 >>
rect 255 99 256 100 
<< m1 >>
rect 265 99 266 100 
<< m1 >>
rect 280 99 281 100 
<< m1 >>
rect 283 99 284 100 
<< m1 >>
rect 307 99 308 100 
<< m1 >>
rect 334 99 335 100 
<< m1 >>
rect 343 99 344 100 
<< m2 >>
rect 343 99 344 100 
<< m2c >>
rect 343 99 344 100 
<< m1 >>
rect 343 99 344 100 
<< m2 >>
rect 343 99 344 100 
<< m2 >>
rect 344 99 345 100 
<< m1 >>
rect 345 99 346 100 
<< m2 >>
rect 345 99 346 100 
<< m2 >>
rect 346 99 347 100 
<< m1 >>
rect 352 99 353 100 
<< m1 >>
rect 361 99 362 100 
<< m1 >>
rect 366 99 367 100 
<< m2 >>
rect 369 99 370 100 
<< m1 >>
rect 370 99 371 100 
<< m1 >>
rect 373 99 374 100 
<< m2 >>
rect 374 99 375 100 
<< m1 >>
rect 375 99 376 100 
<< m2 >>
rect 375 99 376 100 
<< m2c >>
rect 375 99 376 100 
<< m1 >>
rect 375 99 376 100 
<< m2 >>
rect 375 99 376 100 
<< m1 >>
rect 376 99 377 100 
<< m1 >>
rect 377 99 378 100 
<< m1 >>
rect 378 99 379 100 
<< m1 >>
rect 379 99 380 100 
<< m1 >>
rect 388 99 389 100 
<< m1 >>
rect 389 99 390 100 
<< m1 >>
rect 390 99 391 100 
<< m2 >>
rect 390 99 391 100 
<< m2c >>
rect 390 99 391 100 
<< m1 >>
rect 390 99 391 100 
<< m2 >>
rect 390 99 391 100 
<< m1 >>
rect 397 99 398 100 
<< m1 >>
rect 456 99 457 100 
<< m2 >>
rect 456 99 457 100 
<< m2c >>
rect 456 99 457 100 
<< m1 >>
rect 456 99 457 100 
<< m2 >>
rect 456 99 457 100 
<< m1 >>
rect 460 99 461 100 
<< m2 >>
rect 460 99 461 100 
<< m2c >>
rect 460 99 461 100 
<< m1 >>
rect 460 99 461 100 
<< m2 >>
rect 460 99 461 100 
<< m1 >>
rect 466 99 467 100 
<< m2 >>
rect 466 99 467 100 
<< m2c >>
rect 466 99 467 100 
<< m1 >>
rect 466 99 467 100 
<< m2 >>
rect 466 99 467 100 
<< m1 >>
rect 478 99 479 100 
<< m1 >>
rect 479 99 480 100 
<< m1 >>
rect 480 99 481 100 
<< m2 >>
rect 480 99 481 100 
<< m2c >>
rect 480 99 481 100 
<< m1 >>
rect 480 99 481 100 
<< m2 >>
rect 480 99 481 100 
<< m1 >>
rect 487 99 488 100 
<< m2 >>
rect 487 99 488 100 
<< m2c >>
rect 487 99 488 100 
<< m1 >>
rect 487 99 488 100 
<< m2 >>
rect 487 99 488 100 
<< m1 >>
rect 502 99 503 100 
<< m1 >>
rect 46 100 47 101 
<< m1 >>
rect 49 100 50 101 
<< m1 >>
rect 52 100 53 101 
<< m1 >>
rect 64 100 65 101 
<< m1 >>
rect 73 100 74 101 
<< m1 >>
rect 92 100 93 101 
<< m2 >>
rect 92 100 93 101 
<< m2c >>
rect 92 100 93 101 
<< m1 >>
rect 92 100 93 101 
<< m2 >>
rect 92 100 93 101 
<< m1 >>
rect 96 100 97 101 
<< m2 >>
rect 96 100 97 101 
<< m2c >>
rect 96 100 97 101 
<< m1 >>
rect 96 100 97 101 
<< m2 >>
rect 96 100 97 101 
<< m2 >>
rect 97 100 98 101 
<< m1 >>
rect 98 100 99 101 
<< m2 >>
rect 98 100 99 101 
<< m2 >>
rect 99 100 100 101 
<< m1 >>
rect 100 100 101 101 
<< m2 >>
rect 100 100 101 101 
<< m1 >>
rect 127 100 128 101 
<< m1 >>
rect 129 100 130 101 
<< m1 >>
rect 131 100 132 101 
<< m1 >>
rect 133 100 134 101 
<< m1 >>
rect 134 100 135 101 
<< m1 >>
rect 135 100 136 101 
<< m1 >>
rect 136 100 137 101 
<< m2 >>
rect 136 100 137 101 
<< m1 >>
rect 137 100 138 101 
<< m1 >>
rect 138 100 139 101 
<< m1 >>
rect 139 100 140 101 
<< m1 >>
rect 145 100 146 101 
<< m1 >>
rect 154 100 155 101 
<< m1 >>
rect 155 100 156 101 
<< m1 >>
rect 156 100 157 101 
<< m1 >>
rect 157 100 158 101 
<< m1 >>
rect 160 100 161 101 
<< m1 >>
rect 161 100 162 101 
<< m1 >>
rect 162 100 163 101 
<< m1 >>
rect 163 100 164 101 
<< m1 >>
rect 165 100 166 101 
<< m1 >>
rect 172 100 173 101 
<< m1 >>
rect 178 100 179 101 
<< m1 >>
rect 187 100 188 101 
<< m2 >>
rect 189 100 190 101 
<< m1 >>
rect 190 100 191 101 
<< m1 >>
rect 214 100 215 101 
<< m1 >>
rect 215 100 216 101 
<< m1 >>
rect 216 100 217 101 
<< m1 >>
rect 217 100 218 101 
<< m1 >>
rect 224 100 225 101 
<< m1 >>
rect 229 100 230 101 
<< m1 >>
rect 235 100 236 101 
<< m1 >>
rect 241 100 242 101 
<< m1 >>
rect 250 100 251 101 
<< m1 >>
rect 251 100 252 101 
<< m1 >>
rect 252 100 253 101 
<< m1 >>
rect 253 100 254 101 
<< m1 >>
rect 255 100 256 101 
<< m1 >>
rect 265 100 266 101 
<< m1 >>
rect 268 100 269 101 
<< m1 >>
rect 269 100 270 101 
<< m1 >>
rect 270 100 271 101 
<< m1 >>
rect 271 100 272 101 
<< m1 >>
rect 280 100 281 101 
<< m1 >>
rect 283 100 284 101 
<< m1 >>
rect 307 100 308 101 
<< m1 >>
rect 332 100 333 101 
<< m2 >>
rect 332 100 333 101 
<< m2c >>
rect 332 100 333 101 
<< m1 >>
rect 332 100 333 101 
<< m2 >>
rect 332 100 333 101 
<< m2 >>
rect 333 100 334 101 
<< m1 >>
rect 334 100 335 101 
<< m2 >>
rect 334 100 335 101 
<< m2 >>
rect 335 100 336 101 
<< m1 >>
rect 336 100 337 101 
<< m2 >>
rect 336 100 337 101 
<< m2c >>
rect 336 100 337 101 
<< m1 >>
rect 336 100 337 101 
<< m2 >>
rect 336 100 337 101 
<< m1 >>
rect 337 100 338 101 
<< m1 >>
rect 343 100 344 101 
<< m1 >>
rect 345 100 346 101 
<< m1 >>
rect 352 100 353 101 
<< m1 >>
rect 361 100 362 101 
<< m1 >>
rect 366 100 367 101 
<< m2 >>
rect 369 100 370 101 
<< m1 >>
rect 370 100 371 101 
<< m1 >>
rect 373 100 374 101 
<< m1 >>
rect 379 100 380 101 
<< m1 >>
rect 388 100 389 101 
<< m1 >>
rect 397 100 398 101 
<< m1 >>
rect 430 100 431 101 
<< m1 >>
rect 431 100 432 101 
<< m1 >>
rect 432 100 433 101 
<< m1 >>
rect 433 100 434 101 
<< m1 >>
rect 456 100 457 101 
<< m1 >>
rect 460 100 461 101 
<< m1 >>
rect 466 100 467 101 
<< m1 >>
rect 478 100 479 101 
<< m1 >>
rect 487 100 488 101 
<< m1 >>
rect 502 100 503 101 
<< m1 >>
rect 46 101 47 102 
<< m1 >>
rect 49 101 50 102 
<< m1 >>
rect 52 101 53 102 
<< m1 >>
rect 64 101 65 102 
<< m1 >>
rect 73 101 74 102 
<< m1 >>
rect 92 101 93 102 
<< m1 >>
rect 96 101 97 102 
<< m1 >>
rect 98 101 99 102 
<< m1 >>
rect 100 101 101 102 
<< m1 >>
rect 127 101 128 102 
<< m1 >>
rect 129 101 130 102 
<< m1 >>
rect 131 101 132 102 
<< m1 >>
rect 133 101 134 102 
<< m2 >>
rect 136 101 137 102 
<< m1 >>
rect 139 101 140 102 
<< m1 >>
rect 145 101 146 102 
<< m1 >>
rect 154 101 155 102 
<< m1 >>
rect 157 101 158 102 
<< m1 >>
rect 160 101 161 102 
<< m1 >>
rect 163 101 164 102 
<< m1 >>
rect 165 101 166 102 
<< m1 >>
rect 172 101 173 102 
<< m1 >>
rect 178 101 179 102 
<< m1 >>
rect 187 101 188 102 
<< m2 >>
rect 189 101 190 102 
<< m1 >>
rect 190 101 191 102 
<< m1 >>
rect 214 101 215 102 
<< m1 >>
rect 217 101 218 102 
<< m1 >>
rect 224 101 225 102 
<< m1 >>
rect 229 101 230 102 
<< m1 >>
rect 235 101 236 102 
<< m1 >>
rect 241 101 242 102 
<< m1 >>
rect 250 101 251 102 
<< m1 >>
rect 253 101 254 102 
<< m1 >>
rect 255 101 256 102 
<< m1 >>
rect 265 101 266 102 
<< m1 >>
rect 268 101 269 102 
<< m1 >>
rect 271 101 272 102 
<< m1 >>
rect 280 101 281 102 
<< m1 >>
rect 283 101 284 102 
<< m1 >>
rect 307 101 308 102 
<< m1 >>
rect 332 101 333 102 
<< m1 >>
rect 334 101 335 102 
<< m1 >>
rect 337 101 338 102 
<< m1 >>
rect 343 101 344 102 
<< m1 >>
rect 345 101 346 102 
<< m2 >>
rect 346 101 347 102 
<< m1 >>
rect 347 101 348 102 
<< m2 >>
rect 347 101 348 102 
<< m2c >>
rect 347 101 348 102 
<< m1 >>
rect 347 101 348 102 
<< m2 >>
rect 347 101 348 102 
<< m1 >>
rect 348 101 349 102 
<< m1 >>
rect 349 101 350 102 
<< m1 >>
rect 350 101 351 102 
<< m1 >>
rect 351 101 352 102 
<< m1 >>
rect 352 101 353 102 
<< m1 >>
rect 361 101 362 102 
<< m1 >>
rect 366 101 367 102 
<< m2 >>
rect 369 101 370 102 
<< m1 >>
rect 370 101 371 102 
<< m1 >>
rect 373 101 374 102 
<< m1 >>
rect 379 101 380 102 
<< m1 >>
rect 388 101 389 102 
<< m1 >>
rect 397 101 398 102 
<< m1 >>
rect 430 101 431 102 
<< m1 >>
rect 433 101 434 102 
<< m1 >>
rect 456 101 457 102 
<< m1 >>
rect 460 101 461 102 
<< m1 >>
rect 466 101 467 102 
<< m1 >>
rect 478 101 479 102 
<< m1 >>
rect 487 101 488 102 
<< m1 >>
rect 502 101 503 102 
<< pdiffusion >>
rect 12 102 13 103 
<< pdiffusion >>
rect 13 102 14 103 
<< pdiffusion >>
rect 14 102 15 103 
<< pdiffusion >>
rect 15 102 16 103 
<< pdiffusion >>
rect 16 102 17 103 
<< pdiffusion >>
rect 17 102 18 103 
<< pdiffusion >>
rect 30 102 31 103 
<< pdiffusion >>
rect 31 102 32 103 
<< pdiffusion >>
rect 32 102 33 103 
<< pdiffusion >>
rect 33 102 34 103 
<< pdiffusion >>
rect 34 102 35 103 
<< pdiffusion >>
rect 35 102 36 103 
<< m1 >>
rect 46 102 47 103 
<< pdiffusion >>
rect 48 102 49 103 
<< m1 >>
rect 49 102 50 103 
<< pdiffusion >>
rect 49 102 50 103 
<< pdiffusion >>
rect 50 102 51 103 
<< pdiffusion >>
rect 51 102 52 103 
<< m1 >>
rect 52 102 53 103 
<< pdiffusion >>
rect 52 102 53 103 
<< pdiffusion >>
rect 53 102 54 103 
<< m1 >>
rect 64 102 65 103 
<< pdiffusion >>
rect 66 102 67 103 
<< pdiffusion >>
rect 67 102 68 103 
<< pdiffusion >>
rect 68 102 69 103 
<< pdiffusion >>
rect 69 102 70 103 
<< pdiffusion >>
rect 70 102 71 103 
<< pdiffusion >>
rect 71 102 72 103 
<< m1 >>
rect 73 102 74 103 
<< pdiffusion >>
rect 84 102 85 103 
<< pdiffusion >>
rect 85 102 86 103 
<< pdiffusion >>
rect 86 102 87 103 
<< pdiffusion >>
rect 87 102 88 103 
<< pdiffusion >>
rect 88 102 89 103 
<< pdiffusion >>
rect 89 102 90 103 
<< m1 >>
rect 92 102 93 103 
<< m1 >>
rect 96 102 97 103 
<< m1 >>
rect 98 102 99 103 
<< m1 >>
rect 100 102 101 103 
<< pdiffusion >>
rect 102 102 103 103 
<< pdiffusion >>
rect 103 102 104 103 
<< pdiffusion >>
rect 104 102 105 103 
<< pdiffusion >>
rect 105 102 106 103 
<< pdiffusion >>
rect 106 102 107 103 
<< pdiffusion >>
rect 107 102 108 103 
<< m1 >>
rect 127 102 128 103 
<< m1 >>
rect 129 102 130 103 
<< m1 >>
rect 131 102 132 103 
<< m1 >>
rect 133 102 134 103 
<< m1 >>
rect 136 102 137 103 
<< m2 >>
rect 136 102 137 103 
<< m2c >>
rect 136 102 137 103 
<< m1 >>
rect 136 102 137 103 
<< m2 >>
rect 136 102 137 103 
<< pdiffusion >>
rect 138 102 139 103 
<< m1 >>
rect 139 102 140 103 
<< pdiffusion >>
rect 139 102 140 103 
<< pdiffusion >>
rect 140 102 141 103 
<< pdiffusion >>
rect 141 102 142 103 
<< pdiffusion >>
rect 142 102 143 103 
<< pdiffusion >>
rect 143 102 144 103 
<< m1 >>
rect 145 102 146 103 
<< m1 >>
rect 154 102 155 103 
<< pdiffusion >>
rect 156 102 157 103 
<< m1 >>
rect 157 102 158 103 
<< pdiffusion >>
rect 157 102 158 103 
<< pdiffusion >>
rect 158 102 159 103 
<< pdiffusion >>
rect 159 102 160 103 
<< m1 >>
rect 160 102 161 103 
<< pdiffusion >>
rect 160 102 161 103 
<< pdiffusion >>
rect 161 102 162 103 
<< m1 >>
rect 163 102 164 103 
<< m1 >>
rect 165 102 166 103 
<< m1 >>
rect 172 102 173 103 
<< pdiffusion >>
rect 174 102 175 103 
<< pdiffusion >>
rect 175 102 176 103 
<< pdiffusion >>
rect 176 102 177 103 
<< pdiffusion >>
rect 177 102 178 103 
<< m1 >>
rect 178 102 179 103 
<< pdiffusion >>
rect 178 102 179 103 
<< pdiffusion >>
rect 179 102 180 103 
<< m1 >>
rect 187 102 188 103 
<< m2 >>
rect 189 102 190 103 
<< m1 >>
rect 190 102 191 103 
<< pdiffusion >>
rect 192 102 193 103 
<< pdiffusion >>
rect 193 102 194 103 
<< pdiffusion >>
rect 194 102 195 103 
<< pdiffusion >>
rect 195 102 196 103 
<< pdiffusion >>
rect 196 102 197 103 
<< pdiffusion >>
rect 197 102 198 103 
<< pdiffusion >>
rect 210 102 211 103 
<< pdiffusion >>
rect 211 102 212 103 
<< pdiffusion >>
rect 212 102 213 103 
<< pdiffusion >>
rect 213 102 214 103 
<< m1 >>
rect 214 102 215 103 
<< pdiffusion >>
rect 214 102 215 103 
<< pdiffusion >>
rect 215 102 216 103 
<< m1 >>
rect 217 102 218 103 
<< m1 >>
rect 224 102 225 103 
<< pdiffusion >>
rect 228 102 229 103 
<< m1 >>
rect 229 102 230 103 
<< pdiffusion >>
rect 229 102 230 103 
<< pdiffusion >>
rect 230 102 231 103 
<< pdiffusion >>
rect 231 102 232 103 
<< pdiffusion >>
rect 232 102 233 103 
<< pdiffusion >>
rect 233 102 234 103 
<< m1 >>
rect 235 102 236 103 
<< m1 >>
rect 241 102 242 103 
<< pdiffusion >>
rect 246 102 247 103 
<< pdiffusion >>
rect 247 102 248 103 
<< pdiffusion >>
rect 248 102 249 103 
<< pdiffusion >>
rect 249 102 250 103 
<< m1 >>
rect 250 102 251 103 
<< pdiffusion >>
rect 250 102 251 103 
<< pdiffusion >>
rect 251 102 252 103 
<< m1 >>
rect 253 102 254 103 
<< m1 >>
rect 255 102 256 103 
<< pdiffusion >>
rect 264 102 265 103 
<< m1 >>
rect 265 102 266 103 
<< pdiffusion >>
rect 265 102 266 103 
<< pdiffusion >>
rect 266 102 267 103 
<< pdiffusion >>
rect 267 102 268 103 
<< m1 >>
rect 268 102 269 103 
<< pdiffusion >>
rect 268 102 269 103 
<< pdiffusion >>
rect 269 102 270 103 
<< m1 >>
rect 271 102 272 103 
<< m1 >>
rect 280 102 281 103 
<< m1 >>
rect 283 102 284 103 
<< pdiffusion >>
rect 300 102 301 103 
<< pdiffusion >>
rect 301 102 302 103 
<< pdiffusion >>
rect 302 102 303 103 
<< pdiffusion >>
rect 303 102 304 103 
<< pdiffusion >>
rect 304 102 305 103 
<< pdiffusion >>
rect 305 102 306 103 
<< m1 >>
rect 307 102 308 103 
<< pdiffusion >>
rect 318 102 319 103 
<< pdiffusion >>
rect 319 102 320 103 
<< pdiffusion >>
rect 320 102 321 103 
<< pdiffusion >>
rect 321 102 322 103 
<< pdiffusion >>
rect 322 102 323 103 
<< pdiffusion >>
rect 323 102 324 103 
<< m1 >>
rect 332 102 333 103 
<< m1 >>
rect 334 102 335 103 
<< pdiffusion >>
rect 336 102 337 103 
<< m1 >>
rect 337 102 338 103 
<< pdiffusion >>
rect 337 102 338 103 
<< pdiffusion >>
rect 338 102 339 103 
<< pdiffusion >>
rect 339 102 340 103 
<< pdiffusion >>
rect 340 102 341 103 
<< pdiffusion >>
rect 341 102 342 103 
<< m1 >>
rect 343 102 344 103 
<< m1 >>
rect 345 102 346 103 
<< m2 >>
rect 346 102 347 103 
<< pdiffusion >>
rect 354 102 355 103 
<< pdiffusion >>
rect 355 102 356 103 
<< pdiffusion >>
rect 356 102 357 103 
<< pdiffusion >>
rect 357 102 358 103 
<< pdiffusion >>
rect 358 102 359 103 
<< pdiffusion >>
rect 359 102 360 103 
<< m1 >>
rect 361 102 362 103 
<< m1 >>
rect 366 102 367 103 
<< m2 >>
rect 369 102 370 103 
<< m1 >>
rect 370 102 371 103 
<< pdiffusion >>
rect 372 102 373 103 
<< m1 >>
rect 373 102 374 103 
<< pdiffusion >>
rect 373 102 374 103 
<< pdiffusion >>
rect 374 102 375 103 
<< pdiffusion >>
rect 375 102 376 103 
<< pdiffusion >>
rect 376 102 377 103 
<< pdiffusion >>
rect 377 102 378 103 
<< m1 >>
rect 379 102 380 103 
<< m1 >>
rect 388 102 389 103 
<< pdiffusion >>
rect 390 102 391 103 
<< pdiffusion >>
rect 391 102 392 103 
<< pdiffusion >>
rect 392 102 393 103 
<< pdiffusion >>
rect 393 102 394 103 
<< pdiffusion >>
rect 394 102 395 103 
<< pdiffusion >>
rect 395 102 396 103 
<< m1 >>
rect 397 102 398 103 
<< pdiffusion >>
rect 408 102 409 103 
<< pdiffusion >>
rect 409 102 410 103 
<< pdiffusion >>
rect 410 102 411 103 
<< pdiffusion >>
rect 411 102 412 103 
<< pdiffusion >>
rect 412 102 413 103 
<< pdiffusion >>
rect 413 102 414 103 
<< pdiffusion >>
rect 426 102 427 103 
<< pdiffusion >>
rect 427 102 428 103 
<< pdiffusion >>
rect 428 102 429 103 
<< pdiffusion >>
rect 429 102 430 103 
<< m1 >>
rect 430 102 431 103 
<< pdiffusion >>
rect 430 102 431 103 
<< pdiffusion >>
rect 431 102 432 103 
<< m1 >>
rect 433 102 434 103 
<< pdiffusion >>
rect 444 102 445 103 
<< pdiffusion >>
rect 445 102 446 103 
<< pdiffusion >>
rect 446 102 447 103 
<< pdiffusion >>
rect 447 102 448 103 
<< pdiffusion >>
rect 448 102 449 103 
<< pdiffusion >>
rect 449 102 450 103 
<< m1 >>
rect 456 102 457 103 
<< m1 >>
rect 460 102 461 103 
<< pdiffusion >>
rect 462 102 463 103 
<< pdiffusion >>
rect 463 102 464 103 
<< pdiffusion >>
rect 464 102 465 103 
<< pdiffusion >>
rect 465 102 466 103 
<< m1 >>
rect 466 102 467 103 
<< pdiffusion >>
rect 466 102 467 103 
<< pdiffusion >>
rect 467 102 468 103 
<< m1 >>
rect 478 102 479 103 
<< pdiffusion >>
rect 480 102 481 103 
<< pdiffusion >>
rect 481 102 482 103 
<< pdiffusion >>
rect 482 102 483 103 
<< pdiffusion >>
rect 483 102 484 103 
<< pdiffusion >>
rect 484 102 485 103 
<< pdiffusion >>
rect 485 102 486 103 
<< m1 >>
rect 487 102 488 103 
<< pdiffusion >>
rect 498 102 499 103 
<< pdiffusion >>
rect 499 102 500 103 
<< pdiffusion >>
rect 500 102 501 103 
<< pdiffusion >>
rect 501 102 502 103 
<< m1 >>
rect 502 102 503 103 
<< pdiffusion >>
rect 502 102 503 103 
<< pdiffusion >>
rect 503 102 504 103 
<< pdiffusion >>
rect 516 102 517 103 
<< pdiffusion >>
rect 517 102 518 103 
<< pdiffusion >>
rect 518 102 519 103 
<< pdiffusion >>
rect 519 102 520 103 
<< pdiffusion >>
rect 520 102 521 103 
<< pdiffusion >>
rect 521 102 522 103 
<< pdiffusion >>
rect 12 103 13 104 
<< pdiffusion >>
rect 13 103 14 104 
<< pdiffusion >>
rect 14 103 15 104 
<< pdiffusion >>
rect 15 103 16 104 
<< pdiffusion >>
rect 16 103 17 104 
<< pdiffusion >>
rect 17 103 18 104 
<< pdiffusion >>
rect 30 103 31 104 
<< pdiffusion >>
rect 31 103 32 104 
<< pdiffusion >>
rect 32 103 33 104 
<< pdiffusion >>
rect 33 103 34 104 
<< pdiffusion >>
rect 34 103 35 104 
<< pdiffusion >>
rect 35 103 36 104 
<< m1 >>
rect 46 103 47 104 
<< pdiffusion >>
rect 48 103 49 104 
<< pdiffusion >>
rect 49 103 50 104 
<< pdiffusion >>
rect 50 103 51 104 
<< pdiffusion >>
rect 51 103 52 104 
<< pdiffusion >>
rect 52 103 53 104 
<< pdiffusion >>
rect 53 103 54 104 
<< m1 >>
rect 64 103 65 104 
<< pdiffusion >>
rect 66 103 67 104 
<< pdiffusion >>
rect 67 103 68 104 
<< pdiffusion >>
rect 68 103 69 104 
<< pdiffusion >>
rect 69 103 70 104 
<< pdiffusion >>
rect 70 103 71 104 
<< pdiffusion >>
rect 71 103 72 104 
<< m1 >>
rect 73 103 74 104 
<< pdiffusion >>
rect 84 103 85 104 
<< pdiffusion >>
rect 85 103 86 104 
<< pdiffusion >>
rect 86 103 87 104 
<< pdiffusion >>
rect 87 103 88 104 
<< pdiffusion >>
rect 88 103 89 104 
<< pdiffusion >>
rect 89 103 90 104 
<< m1 >>
rect 92 103 93 104 
<< m1 >>
rect 96 103 97 104 
<< m1 >>
rect 98 103 99 104 
<< m1 >>
rect 100 103 101 104 
<< pdiffusion >>
rect 102 103 103 104 
<< pdiffusion >>
rect 103 103 104 104 
<< pdiffusion >>
rect 104 103 105 104 
<< pdiffusion >>
rect 105 103 106 104 
<< pdiffusion >>
rect 106 103 107 104 
<< pdiffusion >>
rect 107 103 108 104 
<< m1 >>
rect 127 103 128 104 
<< m1 >>
rect 129 103 130 104 
<< m1 >>
rect 131 103 132 104 
<< m1 >>
rect 133 103 134 104 
<< m1 >>
rect 136 103 137 104 
<< pdiffusion >>
rect 138 103 139 104 
<< pdiffusion >>
rect 139 103 140 104 
<< pdiffusion >>
rect 140 103 141 104 
<< pdiffusion >>
rect 141 103 142 104 
<< pdiffusion >>
rect 142 103 143 104 
<< pdiffusion >>
rect 143 103 144 104 
<< m1 >>
rect 145 103 146 104 
<< m1 >>
rect 154 103 155 104 
<< pdiffusion >>
rect 156 103 157 104 
<< pdiffusion >>
rect 157 103 158 104 
<< pdiffusion >>
rect 158 103 159 104 
<< pdiffusion >>
rect 159 103 160 104 
<< pdiffusion >>
rect 160 103 161 104 
<< pdiffusion >>
rect 161 103 162 104 
<< m1 >>
rect 163 103 164 104 
<< m1 >>
rect 165 103 166 104 
<< m1 >>
rect 172 103 173 104 
<< pdiffusion >>
rect 174 103 175 104 
<< pdiffusion >>
rect 175 103 176 104 
<< pdiffusion >>
rect 176 103 177 104 
<< pdiffusion >>
rect 177 103 178 104 
<< pdiffusion >>
rect 178 103 179 104 
<< pdiffusion >>
rect 179 103 180 104 
<< m1 >>
rect 187 103 188 104 
<< m2 >>
rect 189 103 190 104 
<< m1 >>
rect 190 103 191 104 
<< pdiffusion >>
rect 192 103 193 104 
<< pdiffusion >>
rect 193 103 194 104 
<< pdiffusion >>
rect 194 103 195 104 
<< pdiffusion >>
rect 195 103 196 104 
<< pdiffusion >>
rect 196 103 197 104 
<< pdiffusion >>
rect 197 103 198 104 
<< pdiffusion >>
rect 210 103 211 104 
<< pdiffusion >>
rect 211 103 212 104 
<< pdiffusion >>
rect 212 103 213 104 
<< pdiffusion >>
rect 213 103 214 104 
<< pdiffusion >>
rect 214 103 215 104 
<< pdiffusion >>
rect 215 103 216 104 
<< m1 >>
rect 217 103 218 104 
<< m1 >>
rect 224 103 225 104 
<< pdiffusion >>
rect 228 103 229 104 
<< pdiffusion >>
rect 229 103 230 104 
<< pdiffusion >>
rect 230 103 231 104 
<< pdiffusion >>
rect 231 103 232 104 
<< pdiffusion >>
rect 232 103 233 104 
<< pdiffusion >>
rect 233 103 234 104 
<< m1 >>
rect 235 103 236 104 
<< m1 >>
rect 241 103 242 104 
<< pdiffusion >>
rect 246 103 247 104 
<< pdiffusion >>
rect 247 103 248 104 
<< pdiffusion >>
rect 248 103 249 104 
<< pdiffusion >>
rect 249 103 250 104 
<< pdiffusion >>
rect 250 103 251 104 
<< pdiffusion >>
rect 251 103 252 104 
<< m1 >>
rect 253 103 254 104 
<< m1 >>
rect 255 103 256 104 
<< pdiffusion >>
rect 264 103 265 104 
<< pdiffusion >>
rect 265 103 266 104 
<< pdiffusion >>
rect 266 103 267 104 
<< pdiffusion >>
rect 267 103 268 104 
<< pdiffusion >>
rect 268 103 269 104 
<< pdiffusion >>
rect 269 103 270 104 
<< m1 >>
rect 271 103 272 104 
<< m1 >>
rect 280 103 281 104 
<< m1 >>
rect 283 103 284 104 
<< pdiffusion >>
rect 300 103 301 104 
<< pdiffusion >>
rect 301 103 302 104 
<< pdiffusion >>
rect 302 103 303 104 
<< pdiffusion >>
rect 303 103 304 104 
<< pdiffusion >>
rect 304 103 305 104 
<< pdiffusion >>
rect 305 103 306 104 
<< m1 >>
rect 307 103 308 104 
<< pdiffusion >>
rect 318 103 319 104 
<< pdiffusion >>
rect 319 103 320 104 
<< pdiffusion >>
rect 320 103 321 104 
<< pdiffusion >>
rect 321 103 322 104 
<< pdiffusion >>
rect 322 103 323 104 
<< pdiffusion >>
rect 323 103 324 104 
<< m1 >>
rect 332 103 333 104 
<< m1 >>
rect 334 103 335 104 
<< pdiffusion >>
rect 336 103 337 104 
<< pdiffusion >>
rect 337 103 338 104 
<< pdiffusion >>
rect 338 103 339 104 
<< pdiffusion >>
rect 339 103 340 104 
<< pdiffusion >>
rect 340 103 341 104 
<< pdiffusion >>
rect 341 103 342 104 
<< m1 >>
rect 343 103 344 104 
<< m1 >>
rect 345 103 346 104 
<< m2 >>
rect 346 103 347 104 
<< pdiffusion >>
rect 354 103 355 104 
<< pdiffusion >>
rect 355 103 356 104 
<< pdiffusion >>
rect 356 103 357 104 
<< pdiffusion >>
rect 357 103 358 104 
<< pdiffusion >>
rect 358 103 359 104 
<< pdiffusion >>
rect 359 103 360 104 
<< m1 >>
rect 361 103 362 104 
<< m1 >>
rect 366 103 367 104 
<< m2 >>
rect 369 103 370 104 
<< m1 >>
rect 370 103 371 104 
<< pdiffusion >>
rect 372 103 373 104 
<< pdiffusion >>
rect 373 103 374 104 
<< pdiffusion >>
rect 374 103 375 104 
<< pdiffusion >>
rect 375 103 376 104 
<< pdiffusion >>
rect 376 103 377 104 
<< pdiffusion >>
rect 377 103 378 104 
<< m1 >>
rect 379 103 380 104 
<< m1 >>
rect 388 103 389 104 
<< pdiffusion >>
rect 390 103 391 104 
<< pdiffusion >>
rect 391 103 392 104 
<< pdiffusion >>
rect 392 103 393 104 
<< pdiffusion >>
rect 393 103 394 104 
<< pdiffusion >>
rect 394 103 395 104 
<< pdiffusion >>
rect 395 103 396 104 
<< m1 >>
rect 397 103 398 104 
<< pdiffusion >>
rect 408 103 409 104 
<< pdiffusion >>
rect 409 103 410 104 
<< pdiffusion >>
rect 410 103 411 104 
<< pdiffusion >>
rect 411 103 412 104 
<< pdiffusion >>
rect 412 103 413 104 
<< pdiffusion >>
rect 413 103 414 104 
<< pdiffusion >>
rect 426 103 427 104 
<< pdiffusion >>
rect 427 103 428 104 
<< pdiffusion >>
rect 428 103 429 104 
<< pdiffusion >>
rect 429 103 430 104 
<< pdiffusion >>
rect 430 103 431 104 
<< pdiffusion >>
rect 431 103 432 104 
<< m1 >>
rect 433 103 434 104 
<< pdiffusion >>
rect 444 103 445 104 
<< pdiffusion >>
rect 445 103 446 104 
<< pdiffusion >>
rect 446 103 447 104 
<< pdiffusion >>
rect 447 103 448 104 
<< pdiffusion >>
rect 448 103 449 104 
<< pdiffusion >>
rect 449 103 450 104 
<< m1 >>
rect 456 103 457 104 
<< m1 >>
rect 460 103 461 104 
<< pdiffusion >>
rect 462 103 463 104 
<< pdiffusion >>
rect 463 103 464 104 
<< pdiffusion >>
rect 464 103 465 104 
<< pdiffusion >>
rect 465 103 466 104 
<< pdiffusion >>
rect 466 103 467 104 
<< pdiffusion >>
rect 467 103 468 104 
<< m1 >>
rect 478 103 479 104 
<< pdiffusion >>
rect 480 103 481 104 
<< pdiffusion >>
rect 481 103 482 104 
<< pdiffusion >>
rect 482 103 483 104 
<< pdiffusion >>
rect 483 103 484 104 
<< pdiffusion >>
rect 484 103 485 104 
<< pdiffusion >>
rect 485 103 486 104 
<< m1 >>
rect 487 103 488 104 
<< pdiffusion >>
rect 498 103 499 104 
<< pdiffusion >>
rect 499 103 500 104 
<< pdiffusion >>
rect 500 103 501 104 
<< pdiffusion >>
rect 501 103 502 104 
<< pdiffusion >>
rect 502 103 503 104 
<< pdiffusion >>
rect 503 103 504 104 
<< pdiffusion >>
rect 516 103 517 104 
<< pdiffusion >>
rect 517 103 518 104 
<< pdiffusion >>
rect 518 103 519 104 
<< pdiffusion >>
rect 519 103 520 104 
<< pdiffusion >>
rect 520 103 521 104 
<< pdiffusion >>
rect 521 103 522 104 
<< pdiffusion >>
rect 12 104 13 105 
<< pdiffusion >>
rect 13 104 14 105 
<< pdiffusion >>
rect 14 104 15 105 
<< pdiffusion >>
rect 15 104 16 105 
<< pdiffusion >>
rect 16 104 17 105 
<< pdiffusion >>
rect 17 104 18 105 
<< pdiffusion >>
rect 30 104 31 105 
<< pdiffusion >>
rect 31 104 32 105 
<< pdiffusion >>
rect 32 104 33 105 
<< pdiffusion >>
rect 33 104 34 105 
<< pdiffusion >>
rect 34 104 35 105 
<< pdiffusion >>
rect 35 104 36 105 
<< m1 >>
rect 46 104 47 105 
<< pdiffusion >>
rect 48 104 49 105 
<< pdiffusion >>
rect 49 104 50 105 
<< pdiffusion >>
rect 50 104 51 105 
<< pdiffusion >>
rect 51 104 52 105 
<< pdiffusion >>
rect 52 104 53 105 
<< pdiffusion >>
rect 53 104 54 105 
<< m1 >>
rect 64 104 65 105 
<< pdiffusion >>
rect 66 104 67 105 
<< pdiffusion >>
rect 67 104 68 105 
<< pdiffusion >>
rect 68 104 69 105 
<< pdiffusion >>
rect 69 104 70 105 
<< pdiffusion >>
rect 70 104 71 105 
<< pdiffusion >>
rect 71 104 72 105 
<< m1 >>
rect 73 104 74 105 
<< pdiffusion >>
rect 84 104 85 105 
<< pdiffusion >>
rect 85 104 86 105 
<< pdiffusion >>
rect 86 104 87 105 
<< pdiffusion >>
rect 87 104 88 105 
<< pdiffusion >>
rect 88 104 89 105 
<< pdiffusion >>
rect 89 104 90 105 
<< m1 >>
rect 92 104 93 105 
<< m1 >>
rect 96 104 97 105 
<< m1 >>
rect 98 104 99 105 
<< m1 >>
rect 100 104 101 105 
<< pdiffusion >>
rect 102 104 103 105 
<< pdiffusion >>
rect 103 104 104 105 
<< pdiffusion >>
rect 104 104 105 105 
<< pdiffusion >>
rect 105 104 106 105 
<< pdiffusion >>
rect 106 104 107 105 
<< pdiffusion >>
rect 107 104 108 105 
<< m1 >>
rect 127 104 128 105 
<< m1 >>
rect 129 104 130 105 
<< m1 >>
rect 131 104 132 105 
<< m1 >>
rect 133 104 134 105 
<< m1 >>
rect 136 104 137 105 
<< pdiffusion >>
rect 138 104 139 105 
<< pdiffusion >>
rect 139 104 140 105 
<< pdiffusion >>
rect 140 104 141 105 
<< pdiffusion >>
rect 141 104 142 105 
<< pdiffusion >>
rect 142 104 143 105 
<< pdiffusion >>
rect 143 104 144 105 
<< m1 >>
rect 145 104 146 105 
<< m1 >>
rect 154 104 155 105 
<< pdiffusion >>
rect 156 104 157 105 
<< pdiffusion >>
rect 157 104 158 105 
<< pdiffusion >>
rect 158 104 159 105 
<< pdiffusion >>
rect 159 104 160 105 
<< pdiffusion >>
rect 160 104 161 105 
<< pdiffusion >>
rect 161 104 162 105 
<< m1 >>
rect 163 104 164 105 
<< m1 >>
rect 165 104 166 105 
<< m1 >>
rect 172 104 173 105 
<< pdiffusion >>
rect 174 104 175 105 
<< pdiffusion >>
rect 175 104 176 105 
<< pdiffusion >>
rect 176 104 177 105 
<< pdiffusion >>
rect 177 104 178 105 
<< pdiffusion >>
rect 178 104 179 105 
<< pdiffusion >>
rect 179 104 180 105 
<< m1 >>
rect 187 104 188 105 
<< m2 >>
rect 189 104 190 105 
<< m1 >>
rect 190 104 191 105 
<< pdiffusion >>
rect 192 104 193 105 
<< pdiffusion >>
rect 193 104 194 105 
<< pdiffusion >>
rect 194 104 195 105 
<< pdiffusion >>
rect 195 104 196 105 
<< pdiffusion >>
rect 196 104 197 105 
<< pdiffusion >>
rect 197 104 198 105 
<< pdiffusion >>
rect 210 104 211 105 
<< pdiffusion >>
rect 211 104 212 105 
<< pdiffusion >>
rect 212 104 213 105 
<< pdiffusion >>
rect 213 104 214 105 
<< pdiffusion >>
rect 214 104 215 105 
<< pdiffusion >>
rect 215 104 216 105 
<< m1 >>
rect 217 104 218 105 
<< m1 >>
rect 224 104 225 105 
<< pdiffusion >>
rect 228 104 229 105 
<< pdiffusion >>
rect 229 104 230 105 
<< pdiffusion >>
rect 230 104 231 105 
<< pdiffusion >>
rect 231 104 232 105 
<< pdiffusion >>
rect 232 104 233 105 
<< pdiffusion >>
rect 233 104 234 105 
<< m1 >>
rect 235 104 236 105 
<< m1 >>
rect 241 104 242 105 
<< pdiffusion >>
rect 246 104 247 105 
<< pdiffusion >>
rect 247 104 248 105 
<< pdiffusion >>
rect 248 104 249 105 
<< pdiffusion >>
rect 249 104 250 105 
<< pdiffusion >>
rect 250 104 251 105 
<< pdiffusion >>
rect 251 104 252 105 
<< m1 >>
rect 253 104 254 105 
<< m1 >>
rect 255 104 256 105 
<< pdiffusion >>
rect 264 104 265 105 
<< pdiffusion >>
rect 265 104 266 105 
<< pdiffusion >>
rect 266 104 267 105 
<< pdiffusion >>
rect 267 104 268 105 
<< pdiffusion >>
rect 268 104 269 105 
<< pdiffusion >>
rect 269 104 270 105 
<< m1 >>
rect 271 104 272 105 
<< m1 >>
rect 280 104 281 105 
<< m1 >>
rect 283 104 284 105 
<< pdiffusion >>
rect 300 104 301 105 
<< pdiffusion >>
rect 301 104 302 105 
<< pdiffusion >>
rect 302 104 303 105 
<< pdiffusion >>
rect 303 104 304 105 
<< pdiffusion >>
rect 304 104 305 105 
<< pdiffusion >>
rect 305 104 306 105 
<< m1 >>
rect 307 104 308 105 
<< pdiffusion >>
rect 318 104 319 105 
<< pdiffusion >>
rect 319 104 320 105 
<< pdiffusion >>
rect 320 104 321 105 
<< pdiffusion >>
rect 321 104 322 105 
<< pdiffusion >>
rect 322 104 323 105 
<< pdiffusion >>
rect 323 104 324 105 
<< m1 >>
rect 332 104 333 105 
<< m1 >>
rect 334 104 335 105 
<< pdiffusion >>
rect 336 104 337 105 
<< pdiffusion >>
rect 337 104 338 105 
<< pdiffusion >>
rect 338 104 339 105 
<< pdiffusion >>
rect 339 104 340 105 
<< pdiffusion >>
rect 340 104 341 105 
<< pdiffusion >>
rect 341 104 342 105 
<< m1 >>
rect 343 104 344 105 
<< m1 >>
rect 345 104 346 105 
<< m2 >>
rect 346 104 347 105 
<< pdiffusion >>
rect 354 104 355 105 
<< pdiffusion >>
rect 355 104 356 105 
<< pdiffusion >>
rect 356 104 357 105 
<< pdiffusion >>
rect 357 104 358 105 
<< pdiffusion >>
rect 358 104 359 105 
<< pdiffusion >>
rect 359 104 360 105 
<< m1 >>
rect 361 104 362 105 
<< m1 >>
rect 366 104 367 105 
<< m2 >>
rect 369 104 370 105 
<< m1 >>
rect 370 104 371 105 
<< pdiffusion >>
rect 372 104 373 105 
<< pdiffusion >>
rect 373 104 374 105 
<< pdiffusion >>
rect 374 104 375 105 
<< pdiffusion >>
rect 375 104 376 105 
<< pdiffusion >>
rect 376 104 377 105 
<< pdiffusion >>
rect 377 104 378 105 
<< m1 >>
rect 379 104 380 105 
<< m1 >>
rect 388 104 389 105 
<< pdiffusion >>
rect 390 104 391 105 
<< pdiffusion >>
rect 391 104 392 105 
<< pdiffusion >>
rect 392 104 393 105 
<< pdiffusion >>
rect 393 104 394 105 
<< pdiffusion >>
rect 394 104 395 105 
<< pdiffusion >>
rect 395 104 396 105 
<< m1 >>
rect 397 104 398 105 
<< pdiffusion >>
rect 408 104 409 105 
<< pdiffusion >>
rect 409 104 410 105 
<< pdiffusion >>
rect 410 104 411 105 
<< pdiffusion >>
rect 411 104 412 105 
<< pdiffusion >>
rect 412 104 413 105 
<< pdiffusion >>
rect 413 104 414 105 
<< pdiffusion >>
rect 426 104 427 105 
<< pdiffusion >>
rect 427 104 428 105 
<< pdiffusion >>
rect 428 104 429 105 
<< pdiffusion >>
rect 429 104 430 105 
<< pdiffusion >>
rect 430 104 431 105 
<< pdiffusion >>
rect 431 104 432 105 
<< m1 >>
rect 433 104 434 105 
<< pdiffusion >>
rect 444 104 445 105 
<< pdiffusion >>
rect 445 104 446 105 
<< pdiffusion >>
rect 446 104 447 105 
<< pdiffusion >>
rect 447 104 448 105 
<< pdiffusion >>
rect 448 104 449 105 
<< pdiffusion >>
rect 449 104 450 105 
<< m1 >>
rect 456 104 457 105 
<< m1 >>
rect 460 104 461 105 
<< pdiffusion >>
rect 462 104 463 105 
<< pdiffusion >>
rect 463 104 464 105 
<< pdiffusion >>
rect 464 104 465 105 
<< pdiffusion >>
rect 465 104 466 105 
<< pdiffusion >>
rect 466 104 467 105 
<< pdiffusion >>
rect 467 104 468 105 
<< m1 >>
rect 478 104 479 105 
<< pdiffusion >>
rect 480 104 481 105 
<< pdiffusion >>
rect 481 104 482 105 
<< pdiffusion >>
rect 482 104 483 105 
<< pdiffusion >>
rect 483 104 484 105 
<< pdiffusion >>
rect 484 104 485 105 
<< pdiffusion >>
rect 485 104 486 105 
<< m1 >>
rect 487 104 488 105 
<< pdiffusion >>
rect 498 104 499 105 
<< pdiffusion >>
rect 499 104 500 105 
<< pdiffusion >>
rect 500 104 501 105 
<< pdiffusion >>
rect 501 104 502 105 
<< pdiffusion >>
rect 502 104 503 105 
<< pdiffusion >>
rect 503 104 504 105 
<< pdiffusion >>
rect 516 104 517 105 
<< pdiffusion >>
rect 517 104 518 105 
<< pdiffusion >>
rect 518 104 519 105 
<< pdiffusion >>
rect 519 104 520 105 
<< pdiffusion >>
rect 520 104 521 105 
<< pdiffusion >>
rect 521 104 522 105 
<< pdiffusion >>
rect 12 105 13 106 
<< pdiffusion >>
rect 13 105 14 106 
<< pdiffusion >>
rect 14 105 15 106 
<< pdiffusion >>
rect 15 105 16 106 
<< pdiffusion >>
rect 16 105 17 106 
<< pdiffusion >>
rect 17 105 18 106 
<< pdiffusion >>
rect 30 105 31 106 
<< pdiffusion >>
rect 31 105 32 106 
<< pdiffusion >>
rect 32 105 33 106 
<< pdiffusion >>
rect 33 105 34 106 
<< pdiffusion >>
rect 34 105 35 106 
<< pdiffusion >>
rect 35 105 36 106 
<< m1 >>
rect 46 105 47 106 
<< pdiffusion >>
rect 48 105 49 106 
<< pdiffusion >>
rect 49 105 50 106 
<< pdiffusion >>
rect 50 105 51 106 
<< pdiffusion >>
rect 51 105 52 106 
<< pdiffusion >>
rect 52 105 53 106 
<< pdiffusion >>
rect 53 105 54 106 
<< m1 >>
rect 64 105 65 106 
<< pdiffusion >>
rect 66 105 67 106 
<< pdiffusion >>
rect 67 105 68 106 
<< pdiffusion >>
rect 68 105 69 106 
<< pdiffusion >>
rect 69 105 70 106 
<< pdiffusion >>
rect 70 105 71 106 
<< pdiffusion >>
rect 71 105 72 106 
<< m1 >>
rect 73 105 74 106 
<< pdiffusion >>
rect 84 105 85 106 
<< pdiffusion >>
rect 85 105 86 106 
<< pdiffusion >>
rect 86 105 87 106 
<< pdiffusion >>
rect 87 105 88 106 
<< pdiffusion >>
rect 88 105 89 106 
<< pdiffusion >>
rect 89 105 90 106 
<< m1 >>
rect 92 105 93 106 
<< m1 >>
rect 96 105 97 106 
<< m1 >>
rect 98 105 99 106 
<< m1 >>
rect 100 105 101 106 
<< pdiffusion >>
rect 102 105 103 106 
<< pdiffusion >>
rect 103 105 104 106 
<< pdiffusion >>
rect 104 105 105 106 
<< pdiffusion >>
rect 105 105 106 106 
<< pdiffusion >>
rect 106 105 107 106 
<< pdiffusion >>
rect 107 105 108 106 
<< m1 >>
rect 127 105 128 106 
<< m1 >>
rect 129 105 130 106 
<< m1 >>
rect 131 105 132 106 
<< m1 >>
rect 133 105 134 106 
<< m1 >>
rect 136 105 137 106 
<< pdiffusion >>
rect 138 105 139 106 
<< pdiffusion >>
rect 139 105 140 106 
<< pdiffusion >>
rect 140 105 141 106 
<< pdiffusion >>
rect 141 105 142 106 
<< pdiffusion >>
rect 142 105 143 106 
<< pdiffusion >>
rect 143 105 144 106 
<< m1 >>
rect 145 105 146 106 
<< m1 >>
rect 154 105 155 106 
<< pdiffusion >>
rect 156 105 157 106 
<< pdiffusion >>
rect 157 105 158 106 
<< pdiffusion >>
rect 158 105 159 106 
<< pdiffusion >>
rect 159 105 160 106 
<< pdiffusion >>
rect 160 105 161 106 
<< pdiffusion >>
rect 161 105 162 106 
<< m1 >>
rect 163 105 164 106 
<< m1 >>
rect 165 105 166 106 
<< m1 >>
rect 172 105 173 106 
<< pdiffusion >>
rect 174 105 175 106 
<< pdiffusion >>
rect 175 105 176 106 
<< pdiffusion >>
rect 176 105 177 106 
<< pdiffusion >>
rect 177 105 178 106 
<< pdiffusion >>
rect 178 105 179 106 
<< pdiffusion >>
rect 179 105 180 106 
<< m1 >>
rect 187 105 188 106 
<< m2 >>
rect 189 105 190 106 
<< m1 >>
rect 190 105 191 106 
<< pdiffusion >>
rect 192 105 193 106 
<< pdiffusion >>
rect 193 105 194 106 
<< pdiffusion >>
rect 194 105 195 106 
<< pdiffusion >>
rect 195 105 196 106 
<< pdiffusion >>
rect 196 105 197 106 
<< pdiffusion >>
rect 197 105 198 106 
<< pdiffusion >>
rect 210 105 211 106 
<< pdiffusion >>
rect 211 105 212 106 
<< pdiffusion >>
rect 212 105 213 106 
<< pdiffusion >>
rect 213 105 214 106 
<< pdiffusion >>
rect 214 105 215 106 
<< pdiffusion >>
rect 215 105 216 106 
<< m1 >>
rect 217 105 218 106 
<< m1 >>
rect 224 105 225 106 
<< pdiffusion >>
rect 228 105 229 106 
<< pdiffusion >>
rect 229 105 230 106 
<< pdiffusion >>
rect 230 105 231 106 
<< pdiffusion >>
rect 231 105 232 106 
<< pdiffusion >>
rect 232 105 233 106 
<< pdiffusion >>
rect 233 105 234 106 
<< m1 >>
rect 235 105 236 106 
<< m1 >>
rect 241 105 242 106 
<< pdiffusion >>
rect 246 105 247 106 
<< pdiffusion >>
rect 247 105 248 106 
<< pdiffusion >>
rect 248 105 249 106 
<< pdiffusion >>
rect 249 105 250 106 
<< pdiffusion >>
rect 250 105 251 106 
<< pdiffusion >>
rect 251 105 252 106 
<< m1 >>
rect 253 105 254 106 
<< m1 >>
rect 255 105 256 106 
<< pdiffusion >>
rect 264 105 265 106 
<< pdiffusion >>
rect 265 105 266 106 
<< pdiffusion >>
rect 266 105 267 106 
<< pdiffusion >>
rect 267 105 268 106 
<< pdiffusion >>
rect 268 105 269 106 
<< pdiffusion >>
rect 269 105 270 106 
<< m1 >>
rect 271 105 272 106 
<< m1 >>
rect 280 105 281 106 
<< m1 >>
rect 283 105 284 106 
<< pdiffusion >>
rect 300 105 301 106 
<< pdiffusion >>
rect 301 105 302 106 
<< pdiffusion >>
rect 302 105 303 106 
<< pdiffusion >>
rect 303 105 304 106 
<< pdiffusion >>
rect 304 105 305 106 
<< pdiffusion >>
rect 305 105 306 106 
<< m1 >>
rect 307 105 308 106 
<< pdiffusion >>
rect 318 105 319 106 
<< pdiffusion >>
rect 319 105 320 106 
<< pdiffusion >>
rect 320 105 321 106 
<< pdiffusion >>
rect 321 105 322 106 
<< pdiffusion >>
rect 322 105 323 106 
<< pdiffusion >>
rect 323 105 324 106 
<< m1 >>
rect 332 105 333 106 
<< m1 >>
rect 334 105 335 106 
<< pdiffusion >>
rect 336 105 337 106 
<< pdiffusion >>
rect 337 105 338 106 
<< pdiffusion >>
rect 338 105 339 106 
<< pdiffusion >>
rect 339 105 340 106 
<< pdiffusion >>
rect 340 105 341 106 
<< pdiffusion >>
rect 341 105 342 106 
<< m1 >>
rect 343 105 344 106 
<< m1 >>
rect 345 105 346 106 
<< m2 >>
rect 346 105 347 106 
<< pdiffusion >>
rect 354 105 355 106 
<< pdiffusion >>
rect 355 105 356 106 
<< pdiffusion >>
rect 356 105 357 106 
<< pdiffusion >>
rect 357 105 358 106 
<< pdiffusion >>
rect 358 105 359 106 
<< pdiffusion >>
rect 359 105 360 106 
<< m1 >>
rect 361 105 362 106 
<< m1 >>
rect 366 105 367 106 
<< m2 >>
rect 369 105 370 106 
<< m1 >>
rect 370 105 371 106 
<< pdiffusion >>
rect 372 105 373 106 
<< pdiffusion >>
rect 373 105 374 106 
<< pdiffusion >>
rect 374 105 375 106 
<< pdiffusion >>
rect 375 105 376 106 
<< pdiffusion >>
rect 376 105 377 106 
<< pdiffusion >>
rect 377 105 378 106 
<< m1 >>
rect 379 105 380 106 
<< m1 >>
rect 388 105 389 106 
<< pdiffusion >>
rect 390 105 391 106 
<< pdiffusion >>
rect 391 105 392 106 
<< pdiffusion >>
rect 392 105 393 106 
<< pdiffusion >>
rect 393 105 394 106 
<< pdiffusion >>
rect 394 105 395 106 
<< pdiffusion >>
rect 395 105 396 106 
<< m1 >>
rect 397 105 398 106 
<< pdiffusion >>
rect 408 105 409 106 
<< pdiffusion >>
rect 409 105 410 106 
<< pdiffusion >>
rect 410 105 411 106 
<< pdiffusion >>
rect 411 105 412 106 
<< pdiffusion >>
rect 412 105 413 106 
<< pdiffusion >>
rect 413 105 414 106 
<< pdiffusion >>
rect 426 105 427 106 
<< pdiffusion >>
rect 427 105 428 106 
<< pdiffusion >>
rect 428 105 429 106 
<< pdiffusion >>
rect 429 105 430 106 
<< pdiffusion >>
rect 430 105 431 106 
<< pdiffusion >>
rect 431 105 432 106 
<< m1 >>
rect 433 105 434 106 
<< pdiffusion >>
rect 444 105 445 106 
<< pdiffusion >>
rect 445 105 446 106 
<< pdiffusion >>
rect 446 105 447 106 
<< pdiffusion >>
rect 447 105 448 106 
<< pdiffusion >>
rect 448 105 449 106 
<< pdiffusion >>
rect 449 105 450 106 
<< m1 >>
rect 456 105 457 106 
<< m1 >>
rect 460 105 461 106 
<< pdiffusion >>
rect 462 105 463 106 
<< pdiffusion >>
rect 463 105 464 106 
<< pdiffusion >>
rect 464 105 465 106 
<< pdiffusion >>
rect 465 105 466 106 
<< pdiffusion >>
rect 466 105 467 106 
<< pdiffusion >>
rect 467 105 468 106 
<< m1 >>
rect 478 105 479 106 
<< pdiffusion >>
rect 480 105 481 106 
<< pdiffusion >>
rect 481 105 482 106 
<< pdiffusion >>
rect 482 105 483 106 
<< pdiffusion >>
rect 483 105 484 106 
<< pdiffusion >>
rect 484 105 485 106 
<< pdiffusion >>
rect 485 105 486 106 
<< m1 >>
rect 487 105 488 106 
<< pdiffusion >>
rect 498 105 499 106 
<< pdiffusion >>
rect 499 105 500 106 
<< pdiffusion >>
rect 500 105 501 106 
<< pdiffusion >>
rect 501 105 502 106 
<< pdiffusion >>
rect 502 105 503 106 
<< pdiffusion >>
rect 503 105 504 106 
<< pdiffusion >>
rect 516 105 517 106 
<< pdiffusion >>
rect 517 105 518 106 
<< pdiffusion >>
rect 518 105 519 106 
<< pdiffusion >>
rect 519 105 520 106 
<< pdiffusion >>
rect 520 105 521 106 
<< pdiffusion >>
rect 521 105 522 106 
<< pdiffusion >>
rect 12 106 13 107 
<< pdiffusion >>
rect 13 106 14 107 
<< pdiffusion >>
rect 14 106 15 107 
<< pdiffusion >>
rect 15 106 16 107 
<< pdiffusion >>
rect 16 106 17 107 
<< pdiffusion >>
rect 17 106 18 107 
<< pdiffusion >>
rect 30 106 31 107 
<< pdiffusion >>
rect 31 106 32 107 
<< pdiffusion >>
rect 32 106 33 107 
<< pdiffusion >>
rect 33 106 34 107 
<< pdiffusion >>
rect 34 106 35 107 
<< pdiffusion >>
rect 35 106 36 107 
<< m1 >>
rect 46 106 47 107 
<< pdiffusion >>
rect 48 106 49 107 
<< pdiffusion >>
rect 49 106 50 107 
<< pdiffusion >>
rect 50 106 51 107 
<< pdiffusion >>
rect 51 106 52 107 
<< pdiffusion >>
rect 52 106 53 107 
<< pdiffusion >>
rect 53 106 54 107 
<< m1 >>
rect 64 106 65 107 
<< pdiffusion >>
rect 66 106 67 107 
<< pdiffusion >>
rect 67 106 68 107 
<< pdiffusion >>
rect 68 106 69 107 
<< pdiffusion >>
rect 69 106 70 107 
<< pdiffusion >>
rect 70 106 71 107 
<< pdiffusion >>
rect 71 106 72 107 
<< m1 >>
rect 73 106 74 107 
<< pdiffusion >>
rect 84 106 85 107 
<< pdiffusion >>
rect 85 106 86 107 
<< pdiffusion >>
rect 86 106 87 107 
<< pdiffusion >>
rect 87 106 88 107 
<< pdiffusion >>
rect 88 106 89 107 
<< pdiffusion >>
rect 89 106 90 107 
<< m1 >>
rect 92 106 93 107 
<< m1 >>
rect 96 106 97 107 
<< m1 >>
rect 98 106 99 107 
<< m1 >>
rect 100 106 101 107 
<< pdiffusion >>
rect 102 106 103 107 
<< pdiffusion >>
rect 103 106 104 107 
<< pdiffusion >>
rect 104 106 105 107 
<< pdiffusion >>
rect 105 106 106 107 
<< pdiffusion >>
rect 106 106 107 107 
<< pdiffusion >>
rect 107 106 108 107 
<< m1 >>
rect 127 106 128 107 
<< m1 >>
rect 129 106 130 107 
<< m1 >>
rect 131 106 132 107 
<< m1 >>
rect 133 106 134 107 
<< m1 >>
rect 136 106 137 107 
<< pdiffusion >>
rect 138 106 139 107 
<< pdiffusion >>
rect 139 106 140 107 
<< pdiffusion >>
rect 140 106 141 107 
<< pdiffusion >>
rect 141 106 142 107 
<< pdiffusion >>
rect 142 106 143 107 
<< pdiffusion >>
rect 143 106 144 107 
<< m1 >>
rect 145 106 146 107 
<< m1 >>
rect 154 106 155 107 
<< pdiffusion >>
rect 156 106 157 107 
<< pdiffusion >>
rect 157 106 158 107 
<< pdiffusion >>
rect 158 106 159 107 
<< pdiffusion >>
rect 159 106 160 107 
<< pdiffusion >>
rect 160 106 161 107 
<< pdiffusion >>
rect 161 106 162 107 
<< m1 >>
rect 163 106 164 107 
<< m1 >>
rect 165 106 166 107 
<< m1 >>
rect 172 106 173 107 
<< pdiffusion >>
rect 174 106 175 107 
<< pdiffusion >>
rect 175 106 176 107 
<< pdiffusion >>
rect 176 106 177 107 
<< pdiffusion >>
rect 177 106 178 107 
<< pdiffusion >>
rect 178 106 179 107 
<< pdiffusion >>
rect 179 106 180 107 
<< m1 >>
rect 187 106 188 107 
<< m2 >>
rect 189 106 190 107 
<< m1 >>
rect 190 106 191 107 
<< pdiffusion >>
rect 192 106 193 107 
<< pdiffusion >>
rect 193 106 194 107 
<< pdiffusion >>
rect 194 106 195 107 
<< pdiffusion >>
rect 195 106 196 107 
<< pdiffusion >>
rect 196 106 197 107 
<< pdiffusion >>
rect 197 106 198 107 
<< pdiffusion >>
rect 210 106 211 107 
<< pdiffusion >>
rect 211 106 212 107 
<< pdiffusion >>
rect 212 106 213 107 
<< pdiffusion >>
rect 213 106 214 107 
<< pdiffusion >>
rect 214 106 215 107 
<< pdiffusion >>
rect 215 106 216 107 
<< m1 >>
rect 217 106 218 107 
<< m1 >>
rect 224 106 225 107 
<< pdiffusion >>
rect 228 106 229 107 
<< pdiffusion >>
rect 229 106 230 107 
<< pdiffusion >>
rect 230 106 231 107 
<< pdiffusion >>
rect 231 106 232 107 
<< pdiffusion >>
rect 232 106 233 107 
<< pdiffusion >>
rect 233 106 234 107 
<< m1 >>
rect 235 106 236 107 
<< m1 >>
rect 241 106 242 107 
<< pdiffusion >>
rect 246 106 247 107 
<< pdiffusion >>
rect 247 106 248 107 
<< pdiffusion >>
rect 248 106 249 107 
<< pdiffusion >>
rect 249 106 250 107 
<< pdiffusion >>
rect 250 106 251 107 
<< pdiffusion >>
rect 251 106 252 107 
<< m1 >>
rect 253 106 254 107 
<< m1 >>
rect 255 106 256 107 
<< pdiffusion >>
rect 264 106 265 107 
<< pdiffusion >>
rect 265 106 266 107 
<< pdiffusion >>
rect 266 106 267 107 
<< pdiffusion >>
rect 267 106 268 107 
<< pdiffusion >>
rect 268 106 269 107 
<< pdiffusion >>
rect 269 106 270 107 
<< m1 >>
rect 271 106 272 107 
<< m1 >>
rect 280 106 281 107 
<< m1 >>
rect 283 106 284 107 
<< pdiffusion >>
rect 300 106 301 107 
<< pdiffusion >>
rect 301 106 302 107 
<< pdiffusion >>
rect 302 106 303 107 
<< pdiffusion >>
rect 303 106 304 107 
<< pdiffusion >>
rect 304 106 305 107 
<< pdiffusion >>
rect 305 106 306 107 
<< m1 >>
rect 307 106 308 107 
<< pdiffusion >>
rect 318 106 319 107 
<< pdiffusion >>
rect 319 106 320 107 
<< pdiffusion >>
rect 320 106 321 107 
<< pdiffusion >>
rect 321 106 322 107 
<< pdiffusion >>
rect 322 106 323 107 
<< pdiffusion >>
rect 323 106 324 107 
<< m1 >>
rect 332 106 333 107 
<< m1 >>
rect 334 106 335 107 
<< pdiffusion >>
rect 336 106 337 107 
<< pdiffusion >>
rect 337 106 338 107 
<< pdiffusion >>
rect 338 106 339 107 
<< pdiffusion >>
rect 339 106 340 107 
<< pdiffusion >>
rect 340 106 341 107 
<< pdiffusion >>
rect 341 106 342 107 
<< m1 >>
rect 343 106 344 107 
<< m1 >>
rect 345 106 346 107 
<< m2 >>
rect 346 106 347 107 
<< pdiffusion >>
rect 354 106 355 107 
<< pdiffusion >>
rect 355 106 356 107 
<< pdiffusion >>
rect 356 106 357 107 
<< pdiffusion >>
rect 357 106 358 107 
<< pdiffusion >>
rect 358 106 359 107 
<< pdiffusion >>
rect 359 106 360 107 
<< m1 >>
rect 361 106 362 107 
<< m1 >>
rect 366 106 367 107 
<< m2 >>
rect 366 106 367 107 
<< m2c >>
rect 366 106 367 107 
<< m1 >>
rect 366 106 367 107 
<< m2 >>
rect 366 106 367 107 
<< m2 >>
rect 369 106 370 107 
<< m1 >>
rect 370 106 371 107 
<< pdiffusion >>
rect 372 106 373 107 
<< pdiffusion >>
rect 373 106 374 107 
<< pdiffusion >>
rect 374 106 375 107 
<< pdiffusion >>
rect 375 106 376 107 
<< pdiffusion >>
rect 376 106 377 107 
<< pdiffusion >>
rect 377 106 378 107 
<< m1 >>
rect 379 106 380 107 
<< m1 >>
rect 388 106 389 107 
<< pdiffusion >>
rect 390 106 391 107 
<< pdiffusion >>
rect 391 106 392 107 
<< pdiffusion >>
rect 392 106 393 107 
<< pdiffusion >>
rect 393 106 394 107 
<< pdiffusion >>
rect 394 106 395 107 
<< pdiffusion >>
rect 395 106 396 107 
<< m1 >>
rect 397 106 398 107 
<< pdiffusion >>
rect 408 106 409 107 
<< pdiffusion >>
rect 409 106 410 107 
<< pdiffusion >>
rect 410 106 411 107 
<< pdiffusion >>
rect 411 106 412 107 
<< pdiffusion >>
rect 412 106 413 107 
<< pdiffusion >>
rect 413 106 414 107 
<< pdiffusion >>
rect 426 106 427 107 
<< pdiffusion >>
rect 427 106 428 107 
<< pdiffusion >>
rect 428 106 429 107 
<< pdiffusion >>
rect 429 106 430 107 
<< pdiffusion >>
rect 430 106 431 107 
<< pdiffusion >>
rect 431 106 432 107 
<< m1 >>
rect 433 106 434 107 
<< pdiffusion >>
rect 444 106 445 107 
<< pdiffusion >>
rect 445 106 446 107 
<< pdiffusion >>
rect 446 106 447 107 
<< pdiffusion >>
rect 447 106 448 107 
<< pdiffusion >>
rect 448 106 449 107 
<< pdiffusion >>
rect 449 106 450 107 
<< m1 >>
rect 456 106 457 107 
<< m1 >>
rect 460 106 461 107 
<< pdiffusion >>
rect 462 106 463 107 
<< pdiffusion >>
rect 463 106 464 107 
<< pdiffusion >>
rect 464 106 465 107 
<< pdiffusion >>
rect 465 106 466 107 
<< pdiffusion >>
rect 466 106 467 107 
<< pdiffusion >>
rect 467 106 468 107 
<< m1 >>
rect 478 106 479 107 
<< pdiffusion >>
rect 480 106 481 107 
<< pdiffusion >>
rect 481 106 482 107 
<< pdiffusion >>
rect 482 106 483 107 
<< pdiffusion >>
rect 483 106 484 107 
<< pdiffusion >>
rect 484 106 485 107 
<< pdiffusion >>
rect 485 106 486 107 
<< m1 >>
rect 487 106 488 107 
<< pdiffusion >>
rect 498 106 499 107 
<< pdiffusion >>
rect 499 106 500 107 
<< pdiffusion >>
rect 500 106 501 107 
<< pdiffusion >>
rect 501 106 502 107 
<< pdiffusion >>
rect 502 106 503 107 
<< pdiffusion >>
rect 503 106 504 107 
<< pdiffusion >>
rect 516 106 517 107 
<< pdiffusion >>
rect 517 106 518 107 
<< pdiffusion >>
rect 518 106 519 107 
<< pdiffusion >>
rect 519 106 520 107 
<< pdiffusion >>
rect 520 106 521 107 
<< pdiffusion >>
rect 521 106 522 107 
<< pdiffusion >>
rect 12 107 13 108 
<< pdiffusion >>
rect 13 107 14 108 
<< pdiffusion >>
rect 14 107 15 108 
<< pdiffusion >>
rect 15 107 16 108 
<< pdiffusion >>
rect 16 107 17 108 
<< pdiffusion >>
rect 17 107 18 108 
<< pdiffusion >>
rect 30 107 31 108 
<< pdiffusion >>
rect 31 107 32 108 
<< pdiffusion >>
rect 32 107 33 108 
<< pdiffusion >>
rect 33 107 34 108 
<< pdiffusion >>
rect 34 107 35 108 
<< pdiffusion >>
rect 35 107 36 108 
<< m1 >>
rect 46 107 47 108 
<< pdiffusion >>
rect 48 107 49 108 
<< pdiffusion >>
rect 49 107 50 108 
<< pdiffusion >>
rect 50 107 51 108 
<< pdiffusion >>
rect 51 107 52 108 
<< pdiffusion >>
rect 52 107 53 108 
<< pdiffusion >>
rect 53 107 54 108 
<< m1 >>
rect 64 107 65 108 
<< pdiffusion >>
rect 66 107 67 108 
<< pdiffusion >>
rect 67 107 68 108 
<< pdiffusion >>
rect 68 107 69 108 
<< pdiffusion >>
rect 69 107 70 108 
<< pdiffusion >>
rect 70 107 71 108 
<< pdiffusion >>
rect 71 107 72 108 
<< m1 >>
rect 73 107 74 108 
<< pdiffusion >>
rect 84 107 85 108 
<< pdiffusion >>
rect 85 107 86 108 
<< pdiffusion >>
rect 86 107 87 108 
<< pdiffusion >>
rect 87 107 88 108 
<< m1 >>
rect 88 107 89 108 
<< pdiffusion >>
rect 88 107 89 108 
<< pdiffusion >>
rect 89 107 90 108 
<< m1 >>
rect 92 107 93 108 
<< m1 >>
rect 96 107 97 108 
<< m1 >>
rect 98 107 99 108 
<< m1 >>
rect 100 107 101 108 
<< pdiffusion >>
rect 102 107 103 108 
<< pdiffusion >>
rect 103 107 104 108 
<< pdiffusion >>
rect 104 107 105 108 
<< pdiffusion >>
rect 105 107 106 108 
<< pdiffusion >>
rect 106 107 107 108 
<< pdiffusion >>
rect 107 107 108 108 
<< m1 >>
rect 127 107 128 108 
<< m1 >>
rect 129 107 130 108 
<< m1 >>
rect 131 107 132 108 
<< m1 >>
rect 133 107 134 108 
<< m1 >>
rect 136 107 137 108 
<< pdiffusion >>
rect 138 107 139 108 
<< pdiffusion >>
rect 139 107 140 108 
<< pdiffusion >>
rect 140 107 141 108 
<< pdiffusion >>
rect 141 107 142 108 
<< pdiffusion >>
rect 142 107 143 108 
<< pdiffusion >>
rect 143 107 144 108 
<< m1 >>
rect 145 107 146 108 
<< m1 >>
rect 154 107 155 108 
<< pdiffusion >>
rect 156 107 157 108 
<< pdiffusion >>
rect 157 107 158 108 
<< pdiffusion >>
rect 158 107 159 108 
<< pdiffusion >>
rect 159 107 160 108 
<< pdiffusion >>
rect 160 107 161 108 
<< pdiffusion >>
rect 161 107 162 108 
<< m1 >>
rect 163 107 164 108 
<< m1 >>
rect 165 107 166 108 
<< m1 >>
rect 172 107 173 108 
<< pdiffusion >>
rect 174 107 175 108 
<< m1 >>
rect 175 107 176 108 
<< pdiffusion >>
rect 175 107 176 108 
<< pdiffusion >>
rect 176 107 177 108 
<< pdiffusion >>
rect 177 107 178 108 
<< m1 >>
rect 178 107 179 108 
<< pdiffusion >>
rect 178 107 179 108 
<< pdiffusion >>
rect 179 107 180 108 
<< m1 >>
rect 187 107 188 108 
<< m2 >>
rect 189 107 190 108 
<< m1 >>
rect 190 107 191 108 
<< pdiffusion >>
rect 192 107 193 108 
<< pdiffusion >>
rect 193 107 194 108 
<< pdiffusion >>
rect 194 107 195 108 
<< pdiffusion >>
rect 195 107 196 108 
<< pdiffusion >>
rect 196 107 197 108 
<< pdiffusion >>
rect 197 107 198 108 
<< pdiffusion >>
rect 210 107 211 108 
<< pdiffusion >>
rect 211 107 212 108 
<< pdiffusion >>
rect 212 107 213 108 
<< pdiffusion >>
rect 213 107 214 108 
<< m1 >>
rect 214 107 215 108 
<< pdiffusion >>
rect 214 107 215 108 
<< pdiffusion >>
rect 215 107 216 108 
<< m1 >>
rect 217 107 218 108 
<< m1 >>
rect 224 107 225 108 
<< pdiffusion >>
rect 228 107 229 108 
<< m1 >>
rect 229 107 230 108 
<< pdiffusion >>
rect 229 107 230 108 
<< pdiffusion >>
rect 230 107 231 108 
<< pdiffusion >>
rect 231 107 232 108 
<< pdiffusion >>
rect 232 107 233 108 
<< pdiffusion >>
rect 233 107 234 108 
<< m1 >>
rect 235 107 236 108 
<< m1 >>
rect 241 107 242 108 
<< pdiffusion >>
rect 246 107 247 108 
<< pdiffusion >>
rect 247 107 248 108 
<< pdiffusion >>
rect 248 107 249 108 
<< pdiffusion >>
rect 249 107 250 108 
<< m1 >>
rect 250 107 251 108 
<< pdiffusion >>
rect 250 107 251 108 
<< pdiffusion >>
rect 251 107 252 108 
<< m1 >>
rect 253 107 254 108 
<< m1 >>
rect 255 107 256 108 
<< pdiffusion >>
rect 264 107 265 108 
<< pdiffusion >>
rect 265 107 266 108 
<< pdiffusion >>
rect 266 107 267 108 
<< pdiffusion >>
rect 267 107 268 108 
<< pdiffusion >>
rect 268 107 269 108 
<< pdiffusion >>
rect 269 107 270 108 
<< m1 >>
rect 271 107 272 108 
<< m1 >>
rect 280 107 281 108 
<< m1 >>
rect 283 107 284 108 
<< pdiffusion >>
rect 300 107 301 108 
<< m1 >>
rect 301 107 302 108 
<< pdiffusion >>
rect 301 107 302 108 
<< pdiffusion >>
rect 302 107 303 108 
<< pdiffusion >>
rect 303 107 304 108 
<< pdiffusion >>
rect 304 107 305 108 
<< pdiffusion >>
rect 305 107 306 108 
<< m1 >>
rect 307 107 308 108 
<< pdiffusion >>
rect 318 107 319 108 
<< m1 >>
rect 319 107 320 108 
<< pdiffusion >>
rect 319 107 320 108 
<< pdiffusion >>
rect 320 107 321 108 
<< pdiffusion >>
rect 321 107 322 108 
<< pdiffusion >>
rect 322 107 323 108 
<< pdiffusion >>
rect 323 107 324 108 
<< m1 >>
rect 332 107 333 108 
<< m1 >>
rect 334 107 335 108 
<< pdiffusion >>
rect 336 107 337 108 
<< pdiffusion >>
rect 337 107 338 108 
<< pdiffusion >>
rect 338 107 339 108 
<< pdiffusion >>
rect 339 107 340 108 
<< pdiffusion >>
rect 340 107 341 108 
<< pdiffusion >>
rect 341 107 342 108 
<< m1 >>
rect 343 107 344 108 
<< m1 >>
rect 345 107 346 108 
<< m2 >>
rect 346 107 347 108 
<< pdiffusion >>
rect 354 107 355 108 
<< m1 >>
rect 355 107 356 108 
<< pdiffusion >>
rect 355 107 356 108 
<< pdiffusion >>
rect 356 107 357 108 
<< pdiffusion >>
rect 357 107 358 108 
<< pdiffusion >>
rect 358 107 359 108 
<< pdiffusion >>
rect 359 107 360 108 
<< m1 >>
rect 361 107 362 108 
<< m2 >>
rect 366 107 367 108 
<< m2 >>
rect 369 107 370 108 
<< m1 >>
rect 370 107 371 108 
<< pdiffusion >>
rect 372 107 373 108 
<< pdiffusion >>
rect 373 107 374 108 
<< pdiffusion >>
rect 374 107 375 108 
<< pdiffusion >>
rect 375 107 376 108 
<< pdiffusion >>
rect 376 107 377 108 
<< pdiffusion >>
rect 377 107 378 108 
<< m1 >>
rect 379 107 380 108 
<< m1 >>
rect 388 107 389 108 
<< pdiffusion >>
rect 390 107 391 108 
<< pdiffusion >>
rect 391 107 392 108 
<< pdiffusion >>
rect 392 107 393 108 
<< pdiffusion >>
rect 393 107 394 108 
<< pdiffusion >>
rect 394 107 395 108 
<< pdiffusion >>
rect 395 107 396 108 
<< m1 >>
rect 397 107 398 108 
<< pdiffusion >>
rect 408 107 409 108 
<< pdiffusion >>
rect 409 107 410 108 
<< pdiffusion >>
rect 410 107 411 108 
<< pdiffusion >>
rect 411 107 412 108 
<< pdiffusion >>
rect 412 107 413 108 
<< pdiffusion >>
rect 413 107 414 108 
<< pdiffusion >>
rect 426 107 427 108 
<< pdiffusion >>
rect 427 107 428 108 
<< pdiffusion >>
rect 428 107 429 108 
<< pdiffusion >>
rect 429 107 430 108 
<< m1 >>
rect 430 107 431 108 
<< pdiffusion >>
rect 430 107 431 108 
<< pdiffusion >>
rect 431 107 432 108 
<< m1 >>
rect 433 107 434 108 
<< pdiffusion >>
rect 444 107 445 108 
<< pdiffusion >>
rect 445 107 446 108 
<< pdiffusion >>
rect 446 107 447 108 
<< pdiffusion >>
rect 447 107 448 108 
<< pdiffusion >>
rect 448 107 449 108 
<< pdiffusion >>
rect 449 107 450 108 
<< m1 >>
rect 456 107 457 108 
<< m1 >>
rect 460 107 461 108 
<< pdiffusion >>
rect 462 107 463 108 
<< pdiffusion >>
rect 463 107 464 108 
<< pdiffusion >>
rect 464 107 465 108 
<< pdiffusion >>
rect 465 107 466 108 
<< pdiffusion >>
rect 466 107 467 108 
<< pdiffusion >>
rect 467 107 468 108 
<< m1 >>
rect 478 107 479 108 
<< pdiffusion >>
rect 480 107 481 108 
<< m1 >>
rect 481 107 482 108 
<< pdiffusion >>
rect 481 107 482 108 
<< pdiffusion >>
rect 482 107 483 108 
<< pdiffusion >>
rect 483 107 484 108 
<< m1 >>
rect 484 107 485 108 
<< pdiffusion >>
rect 484 107 485 108 
<< pdiffusion >>
rect 485 107 486 108 
<< m1 >>
rect 487 107 488 108 
<< pdiffusion >>
rect 498 107 499 108 
<< pdiffusion >>
rect 499 107 500 108 
<< pdiffusion >>
rect 500 107 501 108 
<< pdiffusion >>
rect 501 107 502 108 
<< pdiffusion >>
rect 502 107 503 108 
<< pdiffusion >>
rect 503 107 504 108 
<< pdiffusion >>
rect 516 107 517 108 
<< pdiffusion >>
rect 517 107 518 108 
<< pdiffusion >>
rect 518 107 519 108 
<< pdiffusion >>
rect 519 107 520 108 
<< pdiffusion >>
rect 520 107 521 108 
<< pdiffusion >>
rect 521 107 522 108 
<< m1 >>
rect 46 108 47 109 
<< m1 >>
rect 64 108 65 109 
<< m1 >>
rect 73 108 74 109 
<< m1 >>
rect 88 108 89 109 
<< m1 >>
rect 92 108 93 109 
<< m1 >>
rect 96 108 97 109 
<< m1 >>
rect 98 108 99 109 
<< m1 >>
rect 100 108 101 109 
<< m1 >>
rect 127 108 128 109 
<< m1 >>
rect 129 108 130 109 
<< m1 >>
rect 131 108 132 109 
<< m1 >>
rect 133 108 134 109 
<< m1 >>
rect 136 108 137 109 
<< m1 >>
rect 145 108 146 109 
<< m1 >>
rect 154 108 155 109 
<< m1 >>
rect 163 108 164 109 
<< m1 >>
rect 165 108 166 109 
<< m1 >>
rect 172 108 173 109 
<< m1 >>
rect 175 108 176 109 
<< m1 >>
rect 178 108 179 109 
<< m2 >>
rect 178 108 179 109 
<< m2c >>
rect 178 108 179 109 
<< m1 >>
rect 178 108 179 109 
<< m2 >>
rect 178 108 179 109 
<< m1 >>
rect 187 108 188 109 
<< m2 >>
rect 187 108 188 109 
<< m2c >>
rect 187 108 188 109 
<< m1 >>
rect 187 108 188 109 
<< m2 >>
rect 187 108 188 109 
<< m2 >>
rect 189 108 190 109 
<< m1 >>
rect 190 108 191 109 
<< m1 >>
rect 214 108 215 109 
<< m1 >>
rect 217 108 218 109 
<< m1 >>
rect 224 108 225 109 
<< m1 >>
rect 229 108 230 109 
<< m1 >>
rect 235 108 236 109 
<< m1 >>
rect 241 108 242 109 
<< m1 >>
rect 250 108 251 109 
<< m1 >>
rect 253 108 254 109 
<< m1 >>
rect 255 108 256 109 
<< m1 >>
rect 271 108 272 109 
<< m1 >>
rect 280 108 281 109 
<< m1 >>
rect 283 108 284 109 
<< m1 >>
rect 301 108 302 109 
<< m1 >>
rect 307 108 308 109 
<< m1 >>
rect 319 108 320 109 
<< m1 >>
rect 332 108 333 109 
<< m1 >>
rect 334 108 335 109 
<< m1 >>
rect 343 108 344 109 
<< m1 >>
rect 345 108 346 109 
<< m2 >>
rect 346 108 347 109 
<< m1 >>
rect 355 108 356 109 
<< m1 >>
rect 361 108 362 109 
<< m1 >>
rect 363 108 364 109 
<< m1 >>
rect 364 108 365 109 
<< m1 >>
rect 365 108 366 109 
<< m1 >>
rect 366 108 367 109 
<< m2 >>
rect 366 108 367 109 
<< m1 >>
rect 367 108 368 109 
<< m1 >>
rect 368 108 369 109 
<< m2 >>
rect 368 108 369 109 
<< m2c >>
rect 368 108 369 109 
<< m1 >>
rect 368 108 369 109 
<< m2 >>
rect 368 108 369 109 
<< m2 >>
rect 369 108 370 109 
<< m1 >>
rect 370 108 371 109 
<< m1 >>
rect 379 108 380 109 
<< m1 >>
rect 388 108 389 109 
<< m1 >>
rect 397 108 398 109 
<< m1 >>
rect 430 108 431 109 
<< m1 >>
rect 433 108 434 109 
<< m1 >>
rect 456 108 457 109 
<< m1 >>
rect 460 108 461 109 
<< m1 >>
rect 478 108 479 109 
<< m1 >>
rect 481 108 482 109 
<< m1 >>
rect 484 108 485 109 
<< m1 >>
rect 487 108 488 109 
<< m1 >>
rect 46 109 47 110 
<< m1 >>
rect 64 109 65 110 
<< m1 >>
rect 73 109 74 110 
<< m1 >>
rect 88 109 89 110 
<< m1 >>
rect 92 109 93 110 
<< m1 >>
rect 96 109 97 110 
<< m1 >>
rect 98 109 99 110 
<< m1 >>
rect 100 109 101 110 
<< m1 >>
rect 127 109 128 110 
<< m1 >>
rect 129 109 130 110 
<< m1 >>
rect 131 109 132 110 
<< m1 >>
rect 133 109 134 110 
<< m1 >>
rect 136 109 137 110 
<< m1 >>
rect 145 109 146 110 
<< m1 >>
rect 154 109 155 110 
<< m1 >>
rect 163 109 164 110 
<< m1 >>
rect 165 109 166 110 
<< m1 >>
rect 172 109 173 110 
<< m1 >>
rect 175 109 176 110 
<< m2 >>
rect 178 109 179 110 
<< m2 >>
rect 179 109 180 110 
<< m2 >>
rect 180 109 181 110 
<< m2 >>
rect 181 109 182 110 
<< m2 >>
rect 182 109 183 110 
<< m2 >>
rect 183 109 184 110 
<< m2 >>
rect 184 109 185 110 
<< m2 >>
rect 185 109 186 110 
<< m2 >>
rect 186 109 187 110 
<< m2 >>
rect 187 109 188 110 
<< m2 >>
rect 189 109 190 110 
<< m1 >>
rect 190 109 191 110 
<< m1 >>
rect 214 109 215 110 
<< m1 >>
rect 217 109 218 110 
<< m1 >>
rect 224 109 225 110 
<< m1 >>
rect 225 109 226 110 
<< m1 >>
rect 226 109 227 110 
<< m1 >>
rect 227 109 228 110 
<< m1 >>
rect 228 109 229 110 
<< m1 >>
rect 229 109 230 110 
<< m1 >>
rect 235 109 236 110 
<< m1 >>
rect 241 109 242 110 
<< m1 >>
rect 250 109 251 110 
<< m1 >>
rect 253 109 254 110 
<< m1 >>
rect 255 109 256 110 
<< m1 >>
rect 271 109 272 110 
<< m1 >>
rect 280 109 281 110 
<< m1 >>
rect 283 109 284 110 
<< m1 >>
rect 301 109 302 110 
<< m1 >>
rect 307 109 308 110 
<< m1 >>
rect 319 109 320 110 
<< m1 >>
rect 332 109 333 110 
<< m1 >>
rect 334 109 335 110 
<< m1 >>
rect 343 109 344 110 
<< m1 >>
rect 345 109 346 110 
<< m2 >>
rect 346 109 347 110 
<< m1 >>
rect 355 109 356 110 
<< m1 >>
rect 361 109 362 110 
<< m1 >>
rect 363 109 364 110 
<< m2 >>
rect 366 109 367 110 
<< m1 >>
rect 370 109 371 110 
<< m1 >>
rect 379 109 380 110 
<< m2 >>
rect 379 109 380 110 
<< m2c >>
rect 379 109 380 110 
<< m1 >>
rect 379 109 380 110 
<< m2 >>
rect 379 109 380 110 
<< m1 >>
rect 388 109 389 110 
<< m1 >>
rect 397 109 398 110 
<< m1 >>
rect 430 109 431 110 
<< m2 >>
rect 431 109 432 110 
<< m1 >>
rect 432 109 433 110 
<< m2 >>
rect 432 109 433 110 
<< m2c >>
rect 432 109 433 110 
<< m1 >>
rect 432 109 433 110 
<< m2 >>
rect 432 109 433 110 
<< m1 >>
rect 433 109 434 110 
<< m1 >>
rect 456 109 457 110 
<< m1 >>
rect 460 109 461 110 
<< m1 >>
rect 478 109 479 110 
<< m1 >>
rect 481 109 482 110 
<< m1 >>
rect 482 109 483 110 
<< m2 >>
rect 482 109 483 110 
<< m2c >>
rect 482 109 483 110 
<< m1 >>
rect 482 109 483 110 
<< m2 >>
rect 482 109 483 110 
<< m2 >>
rect 483 109 484 110 
<< m1 >>
rect 484 109 485 110 
<< m1 >>
rect 487 109 488 110 
<< m1 >>
rect 46 110 47 111 
<< m1 >>
rect 64 110 65 111 
<< m1 >>
rect 73 110 74 111 
<< m1 >>
rect 86 110 87 111 
<< m2 >>
rect 86 110 87 111 
<< m2c >>
rect 86 110 87 111 
<< m1 >>
rect 86 110 87 111 
<< m2 >>
rect 86 110 87 111 
<< m1 >>
rect 87 110 88 111 
<< m1 >>
rect 88 110 89 111 
<< m1 >>
rect 92 110 93 111 
<< m2 >>
rect 92 110 93 111 
<< m2c >>
rect 92 110 93 111 
<< m1 >>
rect 92 110 93 111 
<< m2 >>
rect 92 110 93 111 
<< m1 >>
rect 96 110 97 111 
<< m2 >>
rect 96 110 97 111 
<< m2c >>
rect 96 110 97 111 
<< m1 >>
rect 96 110 97 111 
<< m2 >>
rect 96 110 97 111 
<< m1 >>
rect 98 110 99 111 
<< m2 >>
rect 98 110 99 111 
<< m2c >>
rect 98 110 99 111 
<< m1 >>
rect 98 110 99 111 
<< m2 >>
rect 98 110 99 111 
<< m2 >>
rect 99 110 100 111 
<< m1 >>
rect 100 110 101 111 
<< m2 >>
rect 100 110 101 111 
<< m1 >>
rect 101 110 102 111 
<< m1 >>
rect 102 110 103 111 
<< m2 >>
rect 102 110 103 111 
<< m2c >>
rect 102 110 103 111 
<< m1 >>
rect 102 110 103 111 
<< m2 >>
rect 102 110 103 111 
<< m1 >>
rect 127 110 128 111 
<< m2 >>
rect 127 110 128 111 
<< m2c >>
rect 127 110 128 111 
<< m1 >>
rect 127 110 128 111 
<< m2 >>
rect 127 110 128 111 
<< m1 >>
rect 129 110 130 111 
<< m2 >>
rect 129 110 130 111 
<< m2c >>
rect 129 110 130 111 
<< m1 >>
rect 129 110 130 111 
<< m2 >>
rect 129 110 130 111 
<< m1 >>
rect 131 110 132 111 
<< m2 >>
rect 131 110 132 111 
<< m2c >>
rect 131 110 132 111 
<< m1 >>
rect 131 110 132 111 
<< m2 >>
rect 131 110 132 111 
<< m1 >>
rect 133 110 134 111 
<< m2 >>
rect 133 110 134 111 
<< m2c >>
rect 133 110 134 111 
<< m1 >>
rect 133 110 134 111 
<< m2 >>
rect 133 110 134 111 
<< m1 >>
rect 136 110 137 111 
<< m2 >>
rect 136 110 137 111 
<< m2c >>
rect 136 110 137 111 
<< m1 >>
rect 136 110 137 111 
<< m2 >>
rect 136 110 137 111 
<< m1 >>
rect 145 110 146 111 
<< m2 >>
rect 145 110 146 111 
<< m2c >>
rect 145 110 146 111 
<< m1 >>
rect 145 110 146 111 
<< m2 >>
rect 145 110 146 111 
<< m1 >>
rect 154 110 155 111 
<< m2 >>
rect 154 110 155 111 
<< m2c >>
rect 154 110 155 111 
<< m1 >>
rect 154 110 155 111 
<< m2 >>
rect 154 110 155 111 
<< m1 >>
rect 163 110 164 111 
<< m2 >>
rect 163 110 164 111 
<< m2c >>
rect 163 110 164 111 
<< m1 >>
rect 163 110 164 111 
<< m2 >>
rect 163 110 164 111 
<< m1 >>
rect 165 110 166 111 
<< m2 >>
rect 165 110 166 111 
<< m2c >>
rect 165 110 166 111 
<< m1 >>
rect 165 110 166 111 
<< m2 >>
rect 165 110 166 111 
<< m1 >>
rect 172 110 173 111 
<< m2 >>
rect 172 110 173 111 
<< m2c >>
rect 172 110 173 111 
<< m1 >>
rect 172 110 173 111 
<< m2 >>
rect 172 110 173 111 
<< m1 >>
rect 175 110 176 111 
<< m1 >>
rect 176 110 177 111 
<< m1 >>
rect 177 110 178 111 
<< m1 >>
rect 178 110 179 111 
<< m1 >>
rect 179 110 180 111 
<< m1 >>
rect 180 110 181 111 
<< m1 >>
rect 181 110 182 111 
<< m1 >>
rect 182 110 183 111 
<< m1 >>
rect 183 110 184 111 
<< m1 >>
rect 184 110 185 111 
<< m1 >>
rect 185 110 186 111 
<< m1 >>
rect 186 110 187 111 
<< m1 >>
rect 187 110 188 111 
<< m1 >>
rect 188 110 189 111 
<< m1 >>
rect 189 110 190 111 
<< m2 >>
rect 189 110 190 111 
<< m1 >>
rect 190 110 191 111 
<< m1 >>
rect 214 110 215 111 
<< m2 >>
rect 214 110 215 111 
<< m2c >>
rect 214 110 215 111 
<< m1 >>
rect 214 110 215 111 
<< m2 >>
rect 214 110 215 111 
<< m1 >>
rect 217 110 218 111 
<< m2 >>
rect 217 110 218 111 
<< m2c >>
rect 217 110 218 111 
<< m1 >>
rect 217 110 218 111 
<< m2 >>
rect 217 110 218 111 
<< m1 >>
rect 235 110 236 111 
<< m2 >>
rect 235 110 236 111 
<< m2c >>
rect 235 110 236 111 
<< m1 >>
rect 235 110 236 111 
<< m2 >>
rect 235 110 236 111 
<< m1 >>
rect 241 110 242 111 
<< m2 >>
rect 241 110 242 111 
<< m2c >>
rect 241 110 242 111 
<< m1 >>
rect 241 110 242 111 
<< m2 >>
rect 241 110 242 111 
<< m1 >>
rect 248 110 249 111 
<< m2 >>
rect 248 110 249 111 
<< m2c >>
rect 248 110 249 111 
<< m1 >>
rect 248 110 249 111 
<< m2 >>
rect 248 110 249 111 
<< m1 >>
rect 249 110 250 111 
<< m1 >>
rect 250 110 251 111 
<< m1 >>
rect 253 110 254 111 
<< m2 >>
rect 253 110 254 111 
<< m2c >>
rect 253 110 254 111 
<< m1 >>
rect 253 110 254 111 
<< m2 >>
rect 253 110 254 111 
<< m1 >>
rect 255 110 256 111 
<< m2 >>
rect 255 110 256 111 
<< m2c >>
rect 255 110 256 111 
<< m1 >>
rect 255 110 256 111 
<< m2 >>
rect 255 110 256 111 
<< m1 >>
rect 271 110 272 111 
<< m1 >>
rect 280 110 281 111 
<< m1 >>
rect 283 110 284 111 
<< m1 >>
rect 301 110 302 111 
<< m1 >>
rect 302 110 303 111 
<< m1 >>
rect 303 110 304 111 
<< m1 >>
rect 304 110 305 111 
<< m1 >>
rect 305 110 306 111 
<< m1 >>
rect 306 110 307 111 
<< m1 >>
rect 307 110 308 111 
<< m1 >>
rect 319 110 320 111 
<< m1 >>
rect 320 110 321 111 
<< m1 >>
rect 321 110 322 111 
<< m1 >>
rect 322 110 323 111 
<< m1 >>
rect 323 110 324 111 
<< m1 >>
rect 324 110 325 111 
<< m1 >>
rect 325 110 326 111 
<< m1 >>
rect 326 110 327 111 
<< m1 >>
rect 327 110 328 111 
<< m1 >>
rect 328 110 329 111 
<< m1 >>
rect 329 110 330 111 
<< m1 >>
rect 330 110 331 111 
<< m1 >>
rect 331 110 332 111 
<< m1 >>
rect 332 110 333 111 
<< m1 >>
rect 334 110 335 111 
<< m1 >>
rect 343 110 344 111 
<< m1 >>
rect 345 110 346 111 
<< m2 >>
rect 346 110 347 111 
<< m1 >>
rect 355 110 356 111 
<< m1 >>
rect 361 110 362 111 
<< m2 >>
rect 361 110 362 111 
<< m2 >>
rect 362 110 363 111 
<< m1 >>
rect 363 110 364 111 
<< m2 >>
rect 363 110 364 111 
<< m2c >>
rect 363 110 364 111 
<< m1 >>
rect 363 110 364 111 
<< m2 >>
rect 363 110 364 111 
<< m1 >>
rect 366 110 367 111 
<< m2 >>
rect 366 110 367 111 
<< m2c >>
rect 366 110 367 111 
<< m1 >>
rect 366 110 367 111 
<< m2 >>
rect 366 110 367 111 
<< m1 >>
rect 370 110 371 111 
<< m2 >>
rect 370 110 371 111 
<< m2c >>
rect 370 110 371 111 
<< m1 >>
rect 370 110 371 111 
<< m2 >>
rect 370 110 371 111 
<< m2 >>
rect 379 110 380 111 
<< m1 >>
rect 388 110 389 111 
<< m1 >>
rect 397 110 398 111 
<< m1 >>
rect 430 110 431 111 
<< m2 >>
rect 431 110 432 111 
<< m1 >>
rect 456 110 457 111 
<< m1 >>
rect 460 110 461 111 
<< m1 >>
rect 478 110 479 111 
<< m2 >>
rect 483 110 484 111 
<< m1 >>
rect 484 110 485 111 
<< m2 >>
rect 484 110 485 111 
<< m2 >>
rect 485 110 486 111 
<< m1 >>
rect 486 110 487 111 
<< m2 >>
rect 486 110 487 111 
<< m2c >>
rect 486 110 487 111 
<< m1 >>
rect 486 110 487 111 
<< m2 >>
rect 486 110 487 111 
<< m1 >>
rect 487 110 488 111 
<< m1 >>
rect 46 111 47 112 
<< m1 >>
rect 64 111 65 112 
<< m1 >>
rect 73 111 74 112 
<< m2 >>
rect 86 111 87 112 
<< m2 >>
rect 92 111 93 112 
<< m2 >>
rect 96 111 97 112 
<< m2 >>
rect 100 111 101 112 
<< m2 >>
rect 102 111 103 112 
<< m2 >>
rect 127 111 128 112 
<< m2 >>
rect 129 111 130 112 
<< m2 >>
rect 131 111 132 112 
<< m2 >>
rect 133 111 134 112 
<< m2 >>
rect 136 111 137 112 
<< m2 >>
rect 145 111 146 112 
<< m2 >>
rect 154 111 155 112 
<< m2 >>
rect 163 111 164 112 
<< m2 >>
rect 165 111 166 112 
<< m2 >>
rect 172 111 173 112 
<< m2 >>
rect 189 111 190 112 
<< m2 >>
rect 214 111 215 112 
<< m2 >>
rect 217 111 218 112 
<< m2 >>
rect 235 111 236 112 
<< m2 >>
rect 241 111 242 112 
<< m2 >>
rect 248 111 249 112 
<< m2 >>
rect 253 111 254 112 
<< m2 >>
rect 255 111 256 112 
<< m1 >>
rect 271 111 272 112 
<< m1 >>
rect 280 111 281 112 
<< m1 >>
rect 283 111 284 112 
<< m1 >>
rect 334 111 335 112 
<< m1 >>
rect 343 111 344 112 
<< m1 >>
rect 345 111 346 112 
<< m2 >>
rect 346 111 347 112 
<< m1 >>
rect 355 111 356 112 
<< m1 >>
rect 361 111 362 112 
<< m2 >>
rect 361 111 362 112 
<< m2 >>
rect 366 111 367 112 
<< m2 >>
rect 370 111 371 112 
<< m2 >>
rect 375 111 376 112 
<< m1 >>
rect 376 111 377 112 
<< m2 >>
rect 376 111 377 112 
<< m2c >>
rect 376 111 377 112 
<< m1 >>
rect 376 111 377 112 
<< m2 >>
rect 376 111 377 112 
<< m1 >>
rect 377 111 378 112 
<< m1 >>
rect 378 111 379 112 
<< m1 >>
rect 379 111 380 112 
<< m2 >>
rect 379 111 380 112 
<< m1 >>
rect 380 111 381 112 
<< m1 >>
rect 381 111 382 112 
<< m1 >>
rect 382 111 383 112 
<< m1 >>
rect 383 111 384 112 
<< m1 >>
rect 384 111 385 112 
<< m1 >>
rect 385 111 386 112 
<< m1 >>
rect 386 111 387 112 
<< m1 >>
rect 387 111 388 112 
<< m1 >>
rect 388 111 389 112 
<< m1 >>
rect 397 111 398 112 
<< m1 >>
rect 430 111 431 112 
<< m2 >>
rect 431 111 432 112 
<< m1 >>
rect 456 111 457 112 
<< m1 >>
rect 460 111 461 112 
<< m1 >>
rect 478 111 479 112 
<< m1 >>
rect 484 111 485 112 
<< m1 >>
rect 46 112 47 113 
<< m1 >>
rect 64 112 65 113 
<< m1 >>
rect 73 112 74 113 
<< m1 >>
rect 74 112 75 113 
<< m1 >>
rect 75 112 76 113 
<< m1 >>
rect 76 112 77 113 
<< m1 >>
rect 77 112 78 113 
<< m1 >>
rect 78 112 79 113 
<< m1 >>
rect 79 112 80 113 
<< m1 >>
rect 80 112 81 113 
<< m1 >>
rect 81 112 82 113 
<< m1 >>
rect 82 112 83 113 
<< m1 >>
rect 83 112 84 113 
<< m1 >>
rect 84 112 85 113 
<< m1 >>
rect 85 112 86 113 
<< m1 >>
rect 86 112 87 113 
<< m2 >>
rect 86 112 87 113 
<< m1 >>
rect 87 112 88 113 
<< m1 >>
rect 88 112 89 113 
<< m1 >>
rect 89 112 90 113 
<< m1 >>
rect 90 112 91 113 
<< m1 >>
rect 91 112 92 113 
<< m1 >>
rect 92 112 93 113 
<< m2 >>
rect 92 112 93 113 
<< m1 >>
rect 93 112 94 113 
<< m1 >>
rect 94 112 95 113 
<< m1 >>
rect 95 112 96 113 
<< m1 >>
rect 96 112 97 113 
<< m2 >>
rect 96 112 97 113 
<< m1 >>
rect 97 112 98 113 
<< m1 >>
rect 98 112 99 113 
<< m1 >>
rect 99 112 100 113 
<< m1 >>
rect 100 112 101 113 
<< m2 >>
rect 100 112 101 113 
<< m1 >>
rect 101 112 102 113 
<< m1 >>
rect 102 112 103 113 
<< m2 >>
rect 102 112 103 113 
<< m1 >>
rect 103 112 104 113 
<< m1 >>
rect 104 112 105 113 
<< m1 >>
rect 105 112 106 113 
<< m1 >>
rect 106 112 107 113 
<< m1 >>
rect 107 112 108 113 
<< m1 >>
rect 108 112 109 113 
<< m1 >>
rect 109 112 110 113 
<< m1 >>
rect 110 112 111 113 
<< m1 >>
rect 111 112 112 113 
<< m1 >>
rect 112 112 113 113 
<< m1 >>
rect 113 112 114 113 
<< m1 >>
rect 114 112 115 113 
<< m1 >>
rect 115 112 116 113 
<< m1 >>
rect 116 112 117 113 
<< m1 >>
rect 117 112 118 113 
<< m1 >>
rect 118 112 119 113 
<< m1 >>
rect 119 112 120 113 
<< m1 >>
rect 120 112 121 113 
<< m1 >>
rect 121 112 122 113 
<< m1 >>
rect 122 112 123 113 
<< m1 >>
rect 123 112 124 113 
<< m1 >>
rect 124 112 125 113 
<< m1 >>
rect 125 112 126 113 
<< m1 >>
rect 126 112 127 113 
<< m1 >>
rect 127 112 128 113 
<< m2 >>
rect 127 112 128 113 
<< m1 >>
rect 128 112 129 113 
<< m1 >>
rect 129 112 130 113 
<< m2 >>
rect 129 112 130 113 
<< m1 >>
rect 130 112 131 113 
<< m1 >>
rect 131 112 132 113 
<< m2 >>
rect 131 112 132 113 
<< m1 >>
rect 132 112 133 113 
<< m1 >>
rect 133 112 134 113 
<< m2 >>
rect 133 112 134 113 
<< m1 >>
rect 134 112 135 113 
<< m1 >>
rect 135 112 136 113 
<< m1 >>
rect 136 112 137 113 
<< m2 >>
rect 136 112 137 113 
<< m1 >>
rect 137 112 138 113 
<< m1 >>
rect 138 112 139 113 
<< m1 >>
rect 139 112 140 113 
<< m1 >>
rect 140 112 141 113 
<< m1 >>
rect 141 112 142 113 
<< m1 >>
rect 142 112 143 113 
<< m1 >>
rect 143 112 144 113 
<< m1 >>
rect 144 112 145 113 
<< m1 >>
rect 145 112 146 113 
<< m2 >>
rect 145 112 146 113 
<< m1 >>
rect 146 112 147 113 
<< m1 >>
rect 147 112 148 113 
<< m1 >>
rect 148 112 149 113 
<< m1 >>
rect 149 112 150 113 
<< m1 >>
rect 150 112 151 113 
<< m1 >>
rect 151 112 152 113 
<< m1 >>
rect 152 112 153 113 
<< m1 >>
rect 153 112 154 113 
<< m1 >>
rect 154 112 155 113 
<< m2 >>
rect 154 112 155 113 
<< m1 >>
rect 155 112 156 113 
<< m1 >>
rect 156 112 157 113 
<< m1 >>
rect 157 112 158 113 
<< m1 >>
rect 158 112 159 113 
<< m1 >>
rect 159 112 160 113 
<< m1 >>
rect 160 112 161 113 
<< m1 >>
rect 161 112 162 113 
<< m1 >>
rect 162 112 163 113 
<< m1 >>
rect 163 112 164 113 
<< m2 >>
rect 163 112 164 113 
<< m1 >>
rect 164 112 165 113 
<< m1 >>
rect 165 112 166 113 
<< m2 >>
rect 165 112 166 113 
<< m1 >>
rect 166 112 167 113 
<< m1 >>
rect 167 112 168 113 
<< m1 >>
rect 168 112 169 113 
<< m1 >>
rect 169 112 170 113 
<< m1 >>
rect 170 112 171 113 
<< m1 >>
rect 171 112 172 113 
<< m1 >>
rect 172 112 173 113 
<< m2 >>
rect 172 112 173 113 
<< m1 >>
rect 173 112 174 113 
<< m1 >>
rect 174 112 175 113 
<< m1 >>
rect 175 112 176 113 
<< m1 >>
rect 176 112 177 113 
<< m1 >>
rect 177 112 178 113 
<< m1 >>
rect 178 112 179 113 
<< m1 >>
rect 179 112 180 113 
<< m1 >>
rect 180 112 181 113 
<< m1 >>
rect 181 112 182 113 
<< m1 >>
rect 182 112 183 113 
<< m1 >>
rect 183 112 184 113 
<< m1 >>
rect 184 112 185 113 
<< m1 >>
rect 185 112 186 113 
<< m1 >>
rect 186 112 187 113 
<< m1 >>
rect 187 112 188 113 
<< m1 >>
rect 188 112 189 113 
<< m1 >>
rect 189 112 190 113 
<< m2 >>
rect 189 112 190 113 
<< m1 >>
rect 190 112 191 113 
<< m1 >>
rect 191 112 192 113 
<< m1 >>
rect 192 112 193 113 
<< m1 >>
rect 193 112 194 113 
<< m1 >>
rect 194 112 195 113 
<< m1 >>
rect 195 112 196 113 
<< m1 >>
rect 196 112 197 113 
<< m1 >>
rect 197 112 198 113 
<< m1 >>
rect 198 112 199 113 
<< m1 >>
rect 199 112 200 113 
<< m1 >>
rect 200 112 201 113 
<< m1 >>
rect 201 112 202 113 
<< m1 >>
rect 202 112 203 113 
<< m1 >>
rect 203 112 204 113 
<< m1 >>
rect 204 112 205 113 
<< m1 >>
rect 205 112 206 113 
<< m1 >>
rect 206 112 207 113 
<< m1 >>
rect 207 112 208 113 
<< m1 >>
rect 208 112 209 113 
<< m1 >>
rect 209 112 210 113 
<< m1 >>
rect 210 112 211 113 
<< m1 >>
rect 211 112 212 113 
<< m1 >>
rect 212 112 213 113 
<< m1 >>
rect 213 112 214 113 
<< m1 >>
rect 214 112 215 113 
<< m2 >>
rect 214 112 215 113 
<< m1 >>
rect 215 112 216 113 
<< m1 >>
rect 216 112 217 113 
<< m1 >>
rect 217 112 218 113 
<< m2 >>
rect 217 112 218 113 
<< m1 >>
rect 218 112 219 113 
<< m1 >>
rect 219 112 220 113 
<< m1 >>
rect 220 112 221 113 
<< m1 >>
rect 221 112 222 113 
<< m1 >>
rect 222 112 223 113 
<< m1 >>
rect 223 112 224 113 
<< m1 >>
rect 224 112 225 113 
<< m1 >>
rect 225 112 226 113 
<< m1 >>
rect 226 112 227 113 
<< m1 >>
rect 227 112 228 113 
<< m1 >>
rect 228 112 229 113 
<< m1 >>
rect 229 112 230 113 
<< m1 >>
rect 230 112 231 113 
<< m1 >>
rect 231 112 232 113 
<< m1 >>
rect 232 112 233 113 
<< m1 >>
rect 233 112 234 113 
<< m1 >>
rect 234 112 235 113 
<< m1 >>
rect 235 112 236 113 
<< m2 >>
rect 235 112 236 113 
<< m1 >>
rect 236 112 237 113 
<< m1 >>
rect 237 112 238 113 
<< m1 >>
rect 238 112 239 113 
<< m1 >>
rect 239 112 240 113 
<< m1 >>
rect 240 112 241 113 
<< m1 >>
rect 241 112 242 113 
<< m2 >>
rect 241 112 242 113 
<< m1 >>
rect 242 112 243 113 
<< m2 >>
rect 242 112 243 113 
<< m1 >>
rect 243 112 244 113 
<< m2 >>
rect 243 112 244 113 
<< m1 >>
rect 244 112 245 113 
<< m2 >>
rect 244 112 245 113 
<< m1 >>
rect 245 112 246 113 
<< m2 >>
rect 245 112 246 113 
<< m1 >>
rect 246 112 247 113 
<< m2 >>
rect 246 112 247 113 
<< m1 >>
rect 247 112 248 113 
<< m2 >>
rect 247 112 248 113 
<< m1 >>
rect 248 112 249 113 
<< m2 >>
rect 248 112 249 113 
<< m1 >>
rect 249 112 250 113 
<< m1 >>
rect 250 112 251 113 
<< m1 >>
rect 251 112 252 113 
<< m1 >>
rect 252 112 253 113 
<< m1 >>
rect 253 112 254 113 
<< m2 >>
rect 253 112 254 113 
<< m1 >>
rect 254 112 255 113 
<< m1 >>
rect 255 112 256 113 
<< m2 >>
rect 255 112 256 113 
<< m1 >>
rect 256 112 257 113 
<< m1 >>
rect 257 112 258 113 
<< m1 >>
rect 258 112 259 113 
<< m1 >>
rect 259 112 260 113 
<< m1 >>
rect 260 112 261 113 
<< m1 >>
rect 261 112 262 113 
<< m1 >>
rect 262 112 263 113 
<< m1 >>
rect 263 112 264 113 
<< m1 >>
rect 264 112 265 113 
<< m1 >>
rect 265 112 266 113 
<< m1 >>
rect 266 112 267 113 
<< m1 >>
rect 267 112 268 113 
<< m1 >>
rect 268 112 269 113 
<< m1 >>
rect 271 112 272 113 
<< m1 >>
rect 280 112 281 113 
<< m1 >>
rect 283 112 284 113 
<< m1 >>
rect 298 112 299 113 
<< m1 >>
rect 299 112 300 113 
<< m1 >>
rect 300 112 301 113 
<< m1 >>
rect 301 112 302 113 
<< m1 >>
rect 302 112 303 113 
<< m1 >>
rect 303 112 304 113 
<< m1 >>
rect 304 112 305 113 
<< m1 >>
rect 305 112 306 113 
<< m1 >>
rect 306 112 307 113 
<< m1 >>
rect 307 112 308 113 
<< m1 >>
rect 308 112 309 113 
<< m1 >>
rect 309 112 310 113 
<< m1 >>
rect 310 112 311 113 
<< m1 >>
rect 311 112 312 113 
<< m1 >>
rect 312 112 313 113 
<< m1 >>
rect 313 112 314 113 
<< m1 >>
rect 314 112 315 113 
<< m1 >>
rect 315 112 316 113 
<< m1 >>
rect 316 112 317 113 
<< m1 >>
rect 317 112 318 113 
<< m1 >>
rect 318 112 319 113 
<< m1 >>
rect 319 112 320 113 
<< m1 >>
rect 320 112 321 113 
<< m1 >>
rect 321 112 322 113 
<< m1 >>
rect 322 112 323 113 
<< m1 >>
rect 323 112 324 113 
<< m1 >>
rect 324 112 325 113 
<< m1 >>
rect 325 112 326 113 
<< m1 >>
rect 326 112 327 113 
<< m1 >>
rect 327 112 328 113 
<< m1 >>
rect 328 112 329 113 
<< m1 >>
rect 329 112 330 113 
<< m1 >>
rect 330 112 331 113 
<< m1 >>
rect 331 112 332 113 
<< m1 >>
rect 332 112 333 113 
<< m2 >>
rect 332 112 333 113 
<< m2c >>
rect 332 112 333 113 
<< m1 >>
rect 332 112 333 113 
<< m2 >>
rect 332 112 333 113 
<< m2 >>
rect 333 112 334 113 
<< m1 >>
rect 334 112 335 113 
<< m2 >>
rect 334 112 335 113 
<< m2 >>
rect 335 112 336 113 
<< m1 >>
rect 336 112 337 113 
<< m2 >>
rect 336 112 337 113 
<< m2c >>
rect 336 112 337 113 
<< m1 >>
rect 336 112 337 113 
<< m2 >>
rect 336 112 337 113 
<< m1 >>
rect 337 112 338 113 
<< m1 >>
rect 338 112 339 113 
<< m1 >>
rect 339 112 340 113 
<< m1 >>
rect 340 112 341 113 
<< m1 >>
rect 341 112 342 113 
<< m1 >>
rect 342 112 343 113 
<< m1 >>
rect 343 112 344 113 
<< m1 >>
rect 345 112 346 113 
<< m2 >>
rect 346 112 347 113 
<< m1 >>
rect 355 112 356 113 
<< m1 >>
rect 361 112 362 113 
<< m2 >>
rect 361 112 362 113 
<< m1 >>
rect 362 112 363 113 
<< m1 >>
rect 363 112 364 113 
<< m1 >>
rect 364 112 365 113 
<< m1 >>
rect 365 112 366 113 
<< m1 >>
rect 366 112 367 113 
<< m2 >>
rect 366 112 367 113 
<< m1 >>
rect 367 112 368 113 
<< m1 >>
rect 368 112 369 113 
<< m1 >>
rect 369 112 370 113 
<< m1 >>
rect 370 112 371 113 
<< m2 >>
rect 370 112 371 113 
<< m1 >>
rect 371 112 372 113 
<< m1 >>
rect 372 112 373 113 
<< m2 >>
rect 372 112 373 113 
<< m1 >>
rect 373 112 374 113 
<< m2 >>
rect 373 112 374 113 
<< m1 >>
rect 374 112 375 113 
<< m2 >>
rect 374 112 375 113 
<< m2 >>
rect 375 112 376 113 
<< m2 >>
rect 379 112 380 113 
<< m1 >>
rect 397 112 398 113 
<< m1 >>
rect 430 112 431 113 
<< m2 >>
rect 431 112 432 113 
<< m1 >>
rect 456 112 457 113 
<< m1 >>
rect 460 112 461 113 
<< m1 >>
rect 478 112 479 113 
<< m1 >>
rect 484 112 485 113 
<< m1 >>
rect 46 113 47 114 
<< m1 >>
rect 64 113 65 114 
<< m2 >>
rect 72 113 73 114 
<< m2 >>
rect 73 113 74 114 
<< m2 >>
rect 74 113 75 114 
<< m2 >>
rect 75 113 76 114 
<< m2 >>
rect 76 113 77 114 
<< m2 >>
rect 77 113 78 114 
<< m2 >>
rect 78 113 79 114 
<< m2 >>
rect 79 113 80 114 
<< m2 >>
rect 80 113 81 114 
<< m2 >>
rect 81 113 82 114 
<< m2 >>
rect 82 113 83 114 
<< m2 >>
rect 83 113 84 114 
<< m2 >>
rect 84 113 85 114 
<< m2 >>
rect 85 113 86 114 
<< m2 >>
rect 86 113 87 114 
<< m2 >>
rect 92 113 93 114 
<< m2 >>
rect 96 113 97 114 
<< m2 >>
rect 100 113 101 114 
<< m2 >>
rect 102 113 103 114 
<< m2 >>
rect 103 113 104 114 
<< m2 >>
rect 104 113 105 114 
<< m2 >>
rect 105 113 106 114 
<< m2 >>
rect 106 113 107 114 
<< m2 >>
rect 107 113 108 114 
<< m2 >>
rect 108 113 109 114 
<< m2 >>
rect 109 113 110 114 
<< m2 >>
rect 110 113 111 114 
<< m2 >>
rect 111 113 112 114 
<< m2 >>
rect 112 113 113 114 
<< m2 >>
rect 113 113 114 114 
<< m2 >>
rect 114 113 115 114 
<< m2 >>
rect 115 113 116 114 
<< m2 >>
rect 116 113 117 114 
<< m2 >>
rect 117 113 118 114 
<< m2 >>
rect 118 113 119 114 
<< m2 >>
rect 119 113 120 114 
<< m2 >>
rect 120 113 121 114 
<< m2 >>
rect 121 113 122 114 
<< m2 >>
rect 122 113 123 114 
<< m2 >>
rect 123 113 124 114 
<< m2 >>
rect 124 113 125 114 
<< m2 >>
rect 125 113 126 114 
<< m2 >>
rect 127 113 128 114 
<< m2 >>
rect 129 113 130 114 
<< m2 >>
rect 131 113 132 114 
<< m2 >>
rect 133 113 134 114 
<< m2 >>
rect 136 113 137 114 
<< m2 >>
rect 145 113 146 114 
<< m2 >>
rect 154 113 155 114 
<< m2 >>
rect 163 113 164 114 
<< m2 >>
rect 165 113 166 114 
<< m2 >>
rect 172 113 173 114 
<< m2 >>
rect 181 113 182 114 
<< m2 >>
rect 182 113 183 114 
<< m2 >>
rect 183 113 184 114 
<< m2 >>
rect 184 113 185 114 
<< m2 >>
rect 185 113 186 114 
<< m2 >>
rect 186 113 187 114 
<< m2 >>
rect 187 113 188 114 
<< m2 >>
rect 188 113 189 114 
<< m2 >>
rect 189 113 190 114 
<< m2 >>
rect 214 113 215 114 
<< m2 >>
rect 217 113 218 114 
<< m2 >>
rect 235 113 236 114 
<< m2 >>
rect 253 113 254 114 
<< m2 >>
rect 255 113 256 114 
<< m1 >>
rect 268 113 269 114 
<< m1 >>
rect 271 113 272 114 
<< m2 >>
rect 272 113 273 114 
<< m1 >>
rect 273 113 274 114 
<< m2 >>
rect 273 113 274 114 
<< m2c >>
rect 273 113 274 114 
<< m1 >>
rect 273 113 274 114 
<< m2 >>
rect 273 113 274 114 
<< m1 >>
rect 274 113 275 114 
<< m1 >>
rect 275 113 276 114 
<< m1 >>
rect 276 113 277 114 
<< m1 >>
rect 277 113 278 114 
<< m1 >>
rect 278 113 279 114 
<< m2 >>
rect 278 113 279 114 
<< m2c >>
rect 278 113 279 114 
<< m1 >>
rect 278 113 279 114 
<< m2 >>
rect 278 113 279 114 
<< m2 >>
rect 279 113 280 114 
<< m1 >>
rect 280 113 281 114 
<< m2 >>
rect 280 113 281 114 
<< m2 >>
rect 281 113 282 114 
<< m2 >>
rect 282 113 283 114 
<< m1 >>
rect 283 113 284 114 
<< m2 >>
rect 283 113 284 114 
<< m2 >>
rect 284 113 285 114 
<< m1 >>
rect 285 113 286 114 
<< m2 >>
rect 285 113 286 114 
<< m2c >>
rect 285 113 286 114 
<< m1 >>
rect 285 113 286 114 
<< m2 >>
rect 285 113 286 114 
<< m1 >>
rect 286 113 287 114 
<< m1 >>
rect 287 113 288 114 
<< m1 >>
rect 288 113 289 114 
<< m1 >>
rect 289 113 290 114 
<< m1 >>
rect 290 113 291 114 
<< m1 >>
rect 291 113 292 114 
<< m1 >>
rect 292 113 293 114 
<< m1 >>
rect 293 113 294 114 
<< m1 >>
rect 294 113 295 114 
<< m1 >>
rect 295 113 296 114 
<< m1 >>
rect 296 113 297 114 
<< m1 >>
rect 298 113 299 114 
<< m1 >>
rect 334 113 335 114 
<< m1 >>
rect 345 113 346 114 
<< m2 >>
rect 346 113 347 114 
<< m1 >>
rect 355 113 356 114 
<< m2 >>
rect 361 113 362 114 
<< m2 >>
rect 366 113 367 114 
<< m2 >>
rect 370 113 371 114 
<< m2 >>
rect 372 113 373 114 
<< m1 >>
rect 374 113 375 114 
<< m1 >>
rect 379 113 380 114 
<< m2 >>
rect 379 113 380 114 
<< m2c >>
rect 379 113 380 114 
<< m1 >>
rect 379 113 380 114 
<< m2 >>
rect 379 113 380 114 
<< m1 >>
rect 380 113 381 114 
<< m1 >>
rect 381 113 382 114 
<< m1 >>
rect 397 113 398 114 
<< m1 >>
rect 430 113 431 114 
<< m2 >>
rect 431 113 432 114 
<< m1 >>
rect 456 113 457 114 
<< m1 >>
rect 460 113 461 114 
<< m1 >>
rect 478 113 479 114 
<< m1 >>
rect 484 113 485 114 
<< m1 >>
rect 46 114 47 115 
<< m1 >>
rect 64 114 65 115 
<< m1 >>
rect 72 114 73 115 
<< m2 >>
rect 72 114 73 115 
<< m2c >>
rect 72 114 73 115 
<< m1 >>
rect 72 114 73 115 
<< m2 >>
rect 72 114 73 115 
<< m1 >>
rect 92 114 93 115 
<< m2 >>
rect 92 114 93 115 
<< m2c >>
rect 92 114 93 115 
<< m1 >>
rect 92 114 93 115 
<< m2 >>
rect 92 114 93 115 
<< m1 >>
rect 96 114 97 115 
<< m2 >>
rect 96 114 97 115 
<< m2c >>
rect 96 114 97 115 
<< m1 >>
rect 96 114 97 115 
<< m2 >>
rect 96 114 97 115 
<< m1 >>
rect 100 114 101 115 
<< m2 >>
rect 100 114 101 115 
<< m2c >>
rect 100 114 101 115 
<< m1 >>
rect 100 114 101 115 
<< m2 >>
rect 100 114 101 115 
<< m1 >>
rect 124 114 125 115 
<< m1 >>
rect 125 114 126 115 
<< m2 >>
rect 125 114 126 115 
<< m1 >>
rect 126 114 127 115 
<< m1 >>
rect 127 114 128 115 
<< m2 >>
rect 127 114 128 115 
<< m2c >>
rect 127 114 128 115 
<< m1 >>
rect 127 114 128 115 
<< m2 >>
rect 127 114 128 115 
<< m1 >>
rect 129 114 130 115 
<< m2 >>
rect 129 114 130 115 
<< m2c >>
rect 129 114 130 115 
<< m1 >>
rect 129 114 130 115 
<< m2 >>
rect 129 114 130 115 
<< m1 >>
rect 130 114 131 115 
<< m1 >>
rect 131 114 132 115 
<< m2 >>
rect 131 114 132 115 
<< m1 >>
rect 132 114 133 115 
<< m1 >>
rect 133 114 134 115 
<< m2 >>
rect 133 114 134 115 
<< m1 >>
rect 134 114 135 115 
<< m1 >>
rect 135 114 136 115 
<< m1 >>
rect 136 114 137 115 
<< m2 >>
rect 136 114 137 115 
<< m1 >>
rect 137 114 138 115 
<< m1 >>
rect 138 114 139 115 
<< m1 >>
rect 139 114 140 115 
<< m1 >>
rect 140 114 141 115 
<< m1 >>
rect 141 114 142 115 
<< m1 >>
rect 142 114 143 115 
<< m1 >>
rect 143 114 144 115 
<< m1 >>
rect 144 114 145 115 
<< m1 >>
rect 145 114 146 115 
<< m2 >>
rect 145 114 146 115 
<< m1 >>
rect 146 114 147 115 
<< m1 >>
rect 147 114 148 115 
<< m1 >>
rect 148 114 149 115 
<< m1 >>
rect 149 114 150 115 
<< m1 >>
rect 150 114 151 115 
<< m1 >>
rect 151 114 152 115 
<< m1 >>
rect 152 114 153 115 
<< m1 >>
rect 153 114 154 115 
<< m1 >>
rect 154 114 155 115 
<< m2 >>
rect 154 114 155 115 
<< m1 >>
rect 155 114 156 115 
<< m1 >>
rect 156 114 157 115 
<< m1 >>
rect 157 114 158 115 
<< m1 >>
rect 158 114 159 115 
<< m1 >>
rect 159 114 160 115 
<< m1 >>
rect 160 114 161 115 
<< m1 >>
rect 163 114 164 115 
<< m2 >>
rect 163 114 164 115 
<< m2c >>
rect 163 114 164 115 
<< m1 >>
rect 163 114 164 115 
<< m2 >>
rect 163 114 164 115 
<< m1 >>
rect 165 114 166 115 
<< m2 >>
rect 165 114 166 115 
<< m2c >>
rect 165 114 166 115 
<< m1 >>
rect 165 114 166 115 
<< m2 >>
rect 165 114 166 115 
<< m1 >>
rect 172 114 173 115 
<< m2 >>
rect 172 114 173 115 
<< m2c >>
rect 172 114 173 115 
<< m1 >>
rect 172 114 173 115 
<< m2 >>
rect 172 114 173 115 
<< m1 >>
rect 181 114 182 115 
<< m2 >>
rect 181 114 182 115 
<< m2c >>
rect 181 114 182 115 
<< m1 >>
rect 181 114 182 115 
<< m2 >>
rect 181 114 182 115 
<< m1 >>
rect 210 114 211 115 
<< m1 >>
rect 211 114 212 115 
<< m1 >>
rect 212 114 213 115 
<< m1 >>
rect 213 114 214 115 
<< m1 >>
rect 214 114 215 115 
<< m2 >>
rect 214 114 215 115 
<< m2c >>
rect 214 114 215 115 
<< m1 >>
rect 214 114 215 115 
<< m2 >>
rect 214 114 215 115 
<< m1 >>
rect 217 114 218 115 
<< m2 >>
rect 217 114 218 115 
<< m2c >>
rect 217 114 218 115 
<< m1 >>
rect 217 114 218 115 
<< m2 >>
rect 217 114 218 115 
<< m1 >>
rect 235 114 236 115 
<< m2 >>
rect 235 114 236 115 
<< m2c >>
rect 235 114 236 115 
<< m1 >>
rect 235 114 236 115 
<< m2 >>
rect 235 114 236 115 
<< m1 >>
rect 253 114 254 115 
<< m2 >>
rect 253 114 254 115 
<< m2c >>
rect 253 114 254 115 
<< m1 >>
rect 253 114 254 115 
<< m2 >>
rect 253 114 254 115 
<< m1 >>
rect 255 114 256 115 
<< m2 >>
rect 255 114 256 115 
<< m2c >>
rect 255 114 256 115 
<< m1 >>
rect 255 114 256 115 
<< m2 >>
rect 255 114 256 115 
<< m1 >>
rect 268 114 269 115 
<< m1 >>
rect 271 114 272 115 
<< m2 >>
rect 272 114 273 115 
<< m1 >>
rect 280 114 281 115 
<< m1 >>
rect 283 114 284 115 
<< m1 >>
rect 296 114 297 115 
<< m2 >>
rect 296 114 297 115 
<< m2c >>
rect 296 114 297 115 
<< m1 >>
rect 296 114 297 115 
<< m2 >>
rect 296 114 297 115 
<< m2 >>
rect 297 114 298 115 
<< m1 >>
rect 298 114 299 115 
<< m2 >>
rect 298 114 299 115 
<< m2 >>
rect 299 114 300 115 
<< m1 >>
rect 300 114 301 115 
<< m2 >>
rect 300 114 301 115 
<< m2c >>
rect 300 114 301 115 
<< m1 >>
rect 300 114 301 115 
<< m2 >>
rect 300 114 301 115 
<< m1 >>
rect 301 114 302 115 
<< m1 >>
rect 302 114 303 115 
<< m1 >>
rect 303 114 304 115 
<< m1 >>
rect 304 114 305 115 
<< m1 >>
rect 305 114 306 115 
<< m1 >>
rect 306 114 307 115 
<< m1 >>
rect 307 114 308 115 
<< m1 >>
rect 308 114 309 115 
<< m1 >>
rect 309 114 310 115 
<< m1 >>
rect 310 114 311 115 
<< m1 >>
rect 311 114 312 115 
<< m1 >>
rect 312 114 313 115 
<< m1 >>
rect 313 114 314 115 
<< m1 >>
rect 314 114 315 115 
<< m1 >>
rect 315 114 316 115 
<< m1 >>
rect 316 114 317 115 
<< m1 >>
rect 317 114 318 115 
<< m1 >>
rect 318 114 319 115 
<< m1 >>
rect 319 114 320 115 
<< m1 >>
rect 320 114 321 115 
<< m1 >>
rect 321 114 322 115 
<< m1 >>
rect 322 114 323 115 
<< m1 >>
rect 323 114 324 115 
<< m1 >>
rect 324 114 325 115 
<< m1 >>
rect 325 114 326 115 
<< m1 >>
rect 326 114 327 115 
<< m1 >>
rect 327 114 328 115 
<< m1 >>
rect 328 114 329 115 
<< m1 >>
rect 329 114 330 115 
<< m1 >>
rect 330 114 331 115 
<< m1 >>
rect 331 114 332 115 
<< m1 >>
rect 332 114 333 115 
<< m2 >>
rect 332 114 333 115 
<< m2c >>
rect 332 114 333 115 
<< m1 >>
rect 332 114 333 115 
<< m2 >>
rect 332 114 333 115 
<< m2 >>
rect 333 114 334 115 
<< m1 >>
rect 334 114 335 115 
<< m2 >>
rect 334 114 335 115 
<< m2 >>
rect 335 114 336 115 
<< m1 >>
rect 336 114 337 115 
<< m2 >>
rect 336 114 337 115 
<< m2c >>
rect 336 114 337 115 
<< m1 >>
rect 336 114 337 115 
<< m2 >>
rect 336 114 337 115 
<< m1 >>
rect 337 114 338 115 
<< m1 >>
rect 338 114 339 115 
<< m1 >>
rect 339 114 340 115 
<< m1 >>
rect 340 114 341 115 
<< m1 >>
rect 341 114 342 115 
<< m1 >>
rect 342 114 343 115 
<< m1 >>
rect 343 114 344 115 
<< m2 >>
rect 343 114 344 115 
<< m2c >>
rect 343 114 344 115 
<< m1 >>
rect 343 114 344 115 
<< m2 >>
rect 343 114 344 115 
<< m2 >>
rect 344 114 345 115 
<< m1 >>
rect 345 114 346 115 
<< m2 >>
rect 345 114 346 115 
<< m2 >>
rect 346 114 347 115 
<< m1 >>
rect 355 114 356 115 
<< m1 >>
rect 356 114 357 115 
<< m1 >>
rect 357 114 358 115 
<< m1 >>
rect 358 114 359 115 
<< m1 >>
rect 359 114 360 115 
<< m1 >>
rect 360 114 361 115 
<< m1 >>
rect 361 114 362 115 
<< m2 >>
rect 361 114 362 115 
<< m1 >>
rect 366 114 367 115 
<< m2 >>
rect 366 114 367 115 
<< m2c >>
rect 366 114 367 115 
<< m1 >>
rect 366 114 367 115 
<< m2 >>
rect 366 114 367 115 
<< m1 >>
rect 370 114 371 115 
<< m2 >>
rect 370 114 371 115 
<< m2c >>
rect 370 114 371 115 
<< m1 >>
rect 370 114 371 115 
<< m2 >>
rect 370 114 371 115 
<< m1 >>
rect 372 114 373 115 
<< m2 >>
rect 372 114 373 115 
<< m2c >>
rect 372 114 373 115 
<< m1 >>
rect 372 114 373 115 
<< m2 >>
rect 372 114 373 115 
<< m1 >>
rect 374 114 375 115 
<< m1 >>
rect 381 114 382 115 
<< m1 >>
rect 397 114 398 115 
<< m1 >>
rect 430 114 431 115 
<< m2 >>
rect 431 114 432 115 
<< m1 >>
rect 456 114 457 115 
<< m1 >>
rect 460 114 461 115 
<< m1 >>
rect 478 114 479 115 
<< m1 >>
rect 484 114 485 115 
<< m1 >>
rect 46 115 47 116 
<< m1 >>
rect 64 115 65 116 
<< m1 >>
rect 72 115 73 116 
<< m1 >>
rect 92 115 93 116 
<< m1 >>
rect 96 115 97 116 
<< m1 >>
rect 100 115 101 116 
<< m1 >>
rect 124 115 125 116 
<< m2 >>
rect 125 115 126 116 
<< m2 >>
rect 131 115 132 116 
<< m2 >>
rect 133 115 134 116 
<< m2 >>
rect 136 115 137 116 
<< m2 >>
rect 145 115 146 116 
<< m2 >>
rect 154 115 155 116 
<< m1 >>
rect 160 115 161 116 
<< m1 >>
rect 163 115 164 116 
<< m1 >>
rect 165 115 166 116 
<< m1 >>
rect 172 115 173 116 
<< m1 >>
rect 181 115 182 116 
<< m1 >>
rect 210 115 211 116 
<< m1 >>
rect 217 115 218 116 
<< m1 >>
rect 235 115 236 116 
<< m1 >>
rect 253 115 254 116 
<< m1 >>
rect 255 115 256 116 
<< m1 >>
rect 268 115 269 116 
<< m1 >>
rect 271 115 272 116 
<< m2 >>
rect 272 115 273 116 
<< m1 >>
rect 278 115 279 116 
<< m2 >>
rect 278 115 279 116 
<< m2c >>
rect 278 115 279 116 
<< m1 >>
rect 278 115 279 116 
<< m2 >>
rect 278 115 279 116 
<< m2 >>
rect 279 115 280 116 
<< m1 >>
rect 280 115 281 116 
<< m2 >>
rect 280 115 281 116 
<< m2 >>
rect 281 115 282 116 
<< m2 >>
rect 282 115 283 116 
<< m1 >>
rect 283 115 284 116 
<< m2 >>
rect 283 115 284 116 
<< m2 >>
rect 284 115 285 116 
<< m1 >>
rect 298 115 299 116 
<< m1 >>
rect 334 115 335 116 
<< m1 >>
rect 345 115 346 116 
<< m1 >>
rect 361 115 362 116 
<< m2 >>
rect 361 115 362 116 
<< m1 >>
rect 366 115 367 116 
<< m1 >>
rect 370 115 371 116 
<< m1 >>
rect 372 115 373 116 
<< m2 >>
rect 372 115 373 116 
<< m1 >>
rect 374 115 375 116 
<< m2 >>
rect 374 115 375 116 
<< m2c >>
rect 374 115 375 116 
<< m1 >>
rect 374 115 375 116 
<< m2 >>
rect 374 115 375 116 
<< m1 >>
rect 381 115 382 116 
<< m1 >>
rect 397 115 398 116 
<< m1 >>
rect 430 115 431 116 
<< m2 >>
rect 431 115 432 116 
<< m1 >>
rect 456 115 457 116 
<< m1 >>
rect 460 115 461 116 
<< m1 >>
rect 478 115 479 116 
<< m1 >>
rect 484 115 485 116 
<< m1 >>
rect 46 116 47 117 
<< m1 >>
rect 64 116 65 117 
<< m1 >>
rect 72 116 73 117 
<< m1 >>
rect 92 116 93 117 
<< m1 >>
rect 96 116 97 117 
<< m1 >>
rect 97 116 98 117 
<< m1 >>
rect 98 116 99 117 
<< m2 >>
rect 98 116 99 117 
<< m2c >>
rect 98 116 99 117 
<< m1 >>
rect 98 116 99 117 
<< m2 >>
rect 98 116 99 117 
<< m2 >>
rect 99 116 100 117 
<< m1 >>
rect 100 116 101 117 
<< m1 >>
rect 124 116 125 117 
<< m2 >>
rect 125 116 126 117 
<< m1 >>
rect 131 116 132 117 
<< m2 >>
rect 131 116 132 117 
<< m2c >>
rect 131 116 132 117 
<< m1 >>
rect 131 116 132 117 
<< m2 >>
rect 131 116 132 117 
<< m1 >>
rect 133 116 134 117 
<< m2 >>
rect 133 116 134 117 
<< m2c >>
rect 133 116 134 117 
<< m1 >>
rect 133 116 134 117 
<< m2 >>
rect 133 116 134 117 
<< m1 >>
rect 136 116 137 117 
<< m2 >>
rect 136 116 137 117 
<< m2c >>
rect 136 116 137 117 
<< m1 >>
rect 136 116 137 117 
<< m2 >>
rect 136 116 137 117 
<< m1 >>
rect 145 116 146 117 
<< m2 >>
rect 145 116 146 117 
<< m2c >>
rect 145 116 146 117 
<< m1 >>
rect 145 116 146 117 
<< m2 >>
rect 145 116 146 117 
<< m1 >>
rect 154 116 155 117 
<< m2 >>
rect 154 116 155 117 
<< m2c >>
rect 154 116 155 117 
<< m1 >>
rect 154 116 155 117 
<< m2 >>
rect 154 116 155 117 
<< m1 >>
rect 160 116 161 117 
<< m1 >>
rect 163 116 164 117 
<< m1 >>
rect 165 116 166 117 
<< m2 >>
rect 166 116 167 117 
<< m1 >>
rect 167 116 168 117 
<< m2 >>
rect 167 116 168 117 
<< m2c >>
rect 167 116 168 117 
<< m1 >>
rect 167 116 168 117 
<< m2 >>
rect 167 116 168 117 
<< m1 >>
rect 168 116 169 117 
<< m1 >>
rect 169 116 170 117 
<< m1 >>
rect 170 116 171 117 
<< m1 >>
rect 171 116 172 117 
<< m1 >>
rect 172 116 173 117 
<< m1 >>
rect 181 116 182 117 
<< m1 >>
rect 210 116 211 117 
<< m2 >>
rect 210 116 211 117 
<< m2c >>
rect 210 116 211 117 
<< m1 >>
rect 210 116 211 117 
<< m2 >>
rect 210 116 211 117 
<< m1 >>
rect 217 116 218 117 
<< m1 >>
rect 235 116 236 117 
<< m1 >>
rect 253 116 254 117 
<< m1 >>
rect 255 116 256 117 
<< m1 >>
rect 268 116 269 117 
<< m1 >>
rect 271 116 272 117 
<< m2 >>
rect 272 116 273 117 
<< m1 >>
rect 278 116 279 117 
<< m1 >>
rect 280 116 281 117 
<< m1 >>
rect 283 116 284 117 
<< m2 >>
rect 284 116 285 117 
<< m1 >>
rect 298 116 299 117 
<< m1 >>
rect 334 116 335 117 
<< m1 >>
rect 345 116 346 117 
<< m1 >>
rect 361 116 362 117 
<< m2 >>
rect 361 116 362 117 
<< m1 >>
rect 366 116 367 117 
<< m1 >>
rect 370 116 371 117 
<< m2 >>
rect 370 116 371 117 
<< m2 >>
rect 371 116 372 117 
<< m2 >>
rect 372 116 373 117 
<< m2 >>
rect 374 116 375 117 
<< m2 >>
rect 375 116 376 117 
<< m2 >>
rect 376 116 377 117 
<< m2 >>
rect 377 116 378 117 
<< m2 >>
rect 378 116 379 117 
<< m2 >>
rect 379 116 380 117 
<< m1 >>
rect 381 116 382 117 
<< m1 >>
rect 397 116 398 117 
<< m1 >>
rect 430 116 431 117 
<< m2 >>
rect 431 116 432 117 
<< m1 >>
rect 456 116 457 117 
<< m1 >>
rect 460 116 461 117 
<< m1 >>
rect 478 116 479 117 
<< m1 >>
rect 484 116 485 117 
<< m1 >>
rect 46 117 47 118 
<< m1 >>
rect 64 117 65 118 
<< m1 >>
rect 72 117 73 118 
<< m1 >>
rect 92 117 93 118 
<< m2 >>
rect 99 117 100 118 
<< m1 >>
rect 100 117 101 118 
<< m1 >>
rect 103 117 104 118 
<< m1 >>
rect 104 117 105 118 
<< m1 >>
rect 105 117 106 118 
<< m1 >>
rect 106 117 107 118 
<< m1 >>
rect 107 117 108 118 
<< m1 >>
rect 108 117 109 118 
<< m1 >>
rect 109 117 110 118 
<< m1 >>
rect 110 117 111 118 
<< m1 >>
rect 111 117 112 118 
<< m1 >>
rect 112 117 113 118 
<< m1 >>
rect 113 117 114 118 
<< m1 >>
rect 114 117 115 118 
<< m1 >>
rect 115 117 116 118 
<< m1 >>
rect 116 117 117 118 
<< m1 >>
rect 117 117 118 118 
<< m1 >>
rect 118 117 119 118 
<< m1 >>
rect 124 117 125 118 
<< m2 >>
rect 125 117 126 118 
<< m1 >>
rect 131 117 132 118 
<< m1 >>
rect 133 117 134 118 
<< m1 >>
rect 136 117 137 118 
<< m1 >>
rect 145 117 146 118 
<< m1 >>
rect 154 117 155 118 
<< m1 >>
rect 160 117 161 118 
<< m1 >>
rect 163 117 164 118 
<< m1 >>
rect 165 117 166 118 
<< m2 >>
rect 166 117 167 118 
<< m1 >>
rect 181 117 182 118 
<< m2 >>
rect 208 117 209 118 
<< m2 >>
rect 209 117 210 118 
<< m2 >>
rect 210 117 211 118 
<< m1 >>
rect 217 117 218 118 
<< m1 >>
rect 235 117 236 118 
<< m1 >>
rect 253 117 254 118 
<< m1 >>
rect 255 117 256 118 
<< m1 >>
rect 268 117 269 118 
<< m1 >>
rect 271 117 272 118 
<< m2 >>
rect 272 117 273 118 
<< m1 >>
rect 278 117 279 118 
<< m1 >>
rect 280 117 281 118 
<< m1 >>
rect 283 117 284 118 
<< m2 >>
rect 284 117 285 118 
<< m1 >>
rect 298 117 299 118 
<< m1 >>
rect 334 117 335 118 
<< m1 >>
rect 337 117 338 118 
<< m1 >>
rect 338 117 339 118 
<< m1 >>
rect 339 117 340 118 
<< m1 >>
rect 340 117 341 118 
<< m1 >>
rect 341 117 342 118 
<< m1 >>
rect 342 117 343 118 
<< m1 >>
rect 343 117 344 118 
<< m1 >>
rect 345 117 346 118 
<< m1 >>
rect 361 117 362 118 
<< m2 >>
rect 361 117 362 118 
<< m1 >>
rect 366 117 367 118 
<< m1 >>
rect 370 117 371 118 
<< m2 >>
rect 370 117 371 118 
<< m1 >>
rect 373 117 374 118 
<< m1 >>
rect 374 117 375 118 
<< m1 >>
rect 375 117 376 118 
<< m1 >>
rect 376 117 377 118 
<< m1 >>
rect 377 117 378 118 
<< m1 >>
rect 378 117 379 118 
<< m1 >>
rect 379 117 380 118 
<< m2 >>
rect 379 117 380 118 
<< m1 >>
rect 381 117 382 118 
<< m1 >>
rect 397 117 398 118 
<< m1 >>
rect 430 117 431 118 
<< m2 >>
rect 431 117 432 118 
<< m1 >>
rect 456 117 457 118 
<< m1 >>
rect 460 117 461 118 
<< m1 >>
rect 478 117 479 118 
<< m1 >>
rect 484 117 485 118 
<< m1 >>
rect 16 118 17 119 
<< m1 >>
rect 17 118 18 119 
<< m1 >>
rect 18 118 19 119 
<< m1 >>
rect 19 118 20 119 
<< m1 >>
rect 46 118 47 119 
<< m1 >>
rect 64 118 65 119 
<< m1 >>
rect 70 118 71 119 
<< m1 >>
rect 71 118 72 119 
<< m1 >>
rect 72 118 73 119 
<< m1 >>
rect 92 118 93 119 
<< m2 >>
rect 99 118 100 119 
<< m1 >>
rect 100 118 101 119 
<< m1 >>
rect 103 118 104 119 
<< m2 >>
rect 106 118 107 119 
<< m2 >>
rect 107 118 108 119 
<< m2 >>
rect 108 118 109 119 
<< m2 >>
rect 109 118 110 119 
<< m1 >>
rect 118 118 119 119 
<< m1 >>
rect 124 118 125 119 
<< m2 >>
rect 125 118 126 119 
<< m1 >>
rect 126 118 127 119 
<< m2 >>
rect 126 118 127 119 
<< m2c >>
rect 126 118 127 119 
<< m1 >>
rect 126 118 127 119 
<< m2 >>
rect 126 118 127 119 
<< m1 >>
rect 127 118 128 119 
<< m1 >>
rect 128 118 129 119 
<< m1 >>
rect 129 118 130 119 
<< m1 >>
rect 131 118 132 119 
<< m1 >>
rect 133 118 134 119 
<< m1 >>
rect 136 118 137 119 
<< m1 >>
rect 145 118 146 119 
<< m1 >>
rect 154 118 155 119 
<< m1 >>
rect 160 118 161 119 
<< m1 >>
rect 163 118 164 119 
<< m1 >>
rect 165 118 166 119 
<< m2 >>
rect 166 118 167 119 
<< m1 >>
rect 181 118 182 119 
<< m1 >>
rect 199 118 200 119 
<< m1 >>
rect 200 118 201 119 
<< m1 >>
rect 201 118 202 119 
<< m1 >>
rect 202 118 203 119 
<< m1 >>
rect 203 118 204 119 
<< m1 >>
rect 204 118 205 119 
<< m1 >>
rect 205 118 206 119 
<< m1 >>
rect 206 118 207 119 
<< m1 >>
rect 207 118 208 119 
<< m1 >>
rect 208 118 209 119 
<< m2 >>
rect 208 118 209 119 
<< m1 >>
rect 209 118 210 119 
<< m1 >>
rect 210 118 211 119 
<< m1 >>
rect 211 118 212 119 
<< m1 >>
rect 217 118 218 119 
<< m1 >>
rect 235 118 236 119 
<< m1 >>
rect 244 118 245 119 
<< m1 >>
rect 245 118 246 119 
<< m1 >>
rect 246 118 247 119 
<< m1 >>
rect 247 118 248 119 
<< m1 >>
rect 253 118 254 119 
<< m1 >>
rect 255 118 256 119 
<< m1 >>
rect 268 118 269 119 
<< m1 >>
rect 271 118 272 119 
<< m2 >>
rect 272 118 273 119 
<< m1 >>
rect 278 118 279 119 
<< m1 >>
rect 280 118 281 119 
<< m1 >>
rect 283 118 284 119 
<< m2 >>
rect 284 118 285 119 
<< m1 >>
rect 285 118 286 119 
<< m2 >>
rect 285 118 286 119 
<< m2c >>
rect 285 118 286 119 
<< m1 >>
rect 285 118 286 119 
<< m2 >>
rect 285 118 286 119 
<< m1 >>
rect 286 118 287 119 
<< m1 >>
rect 298 118 299 119 
<< m1 >>
rect 334 118 335 119 
<< m1 >>
rect 337 118 338 119 
<< m1 >>
rect 343 118 344 119 
<< m1 >>
rect 345 118 346 119 
<< m1 >>
rect 361 118 362 119 
<< m2 >>
rect 361 118 362 119 
<< m1 >>
rect 366 118 367 119 
<< m1 >>
rect 370 118 371 119 
<< m2 >>
rect 370 118 371 119 
<< m1 >>
rect 373 118 374 119 
<< m1 >>
rect 379 118 380 119 
<< m2 >>
rect 379 118 380 119 
<< m1 >>
rect 381 118 382 119 
<< m1 >>
rect 394 118 395 119 
<< m1 >>
rect 395 118 396 119 
<< m1 >>
rect 396 118 397 119 
<< m1 >>
rect 397 118 398 119 
<< m1 >>
rect 430 118 431 119 
<< m2 >>
rect 431 118 432 119 
<< m1 >>
rect 456 118 457 119 
<< m1 >>
rect 460 118 461 119 
<< m1 >>
rect 461 118 462 119 
<< m1 >>
rect 462 118 463 119 
<< m1 >>
rect 463 118 464 119 
<< m1 >>
rect 478 118 479 119 
<< m1 >>
rect 484 118 485 119 
<< m1 >>
rect 16 119 17 120 
<< m1 >>
rect 19 119 20 120 
<< m1 >>
rect 46 119 47 120 
<< m1 >>
rect 64 119 65 120 
<< m1 >>
rect 70 119 71 120 
<< m1 >>
rect 92 119 93 120 
<< m2 >>
rect 99 119 100 120 
<< m1 >>
rect 100 119 101 120 
<< m1 >>
rect 103 119 104 120 
<< m1 >>
rect 106 119 107 120 
<< m2 >>
rect 106 119 107 120 
<< m2c >>
rect 106 119 107 120 
<< m1 >>
rect 106 119 107 120 
<< m2 >>
rect 106 119 107 120 
<< m1 >>
rect 109 119 110 120 
<< m2 >>
rect 109 119 110 120 
<< m2c >>
rect 109 119 110 120 
<< m1 >>
rect 109 119 110 120 
<< m2 >>
rect 109 119 110 120 
<< m1 >>
rect 118 119 119 120 
<< m1 >>
rect 124 119 125 120 
<< m1 >>
rect 129 119 130 120 
<< m1 >>
rect 131 119 132 120 
<< m1 >>
rect 133 119 134 120 
<< m1 >>
rect 136 119 137 120 
<< m1 >>
rect 145 119 146 120 
<< m1 >>
rect 154 119 155 120 
<< m1 >>
rect 160 119 161 120 
<< m1 >>
rect 163 119 164 120 
<< m1 >>
rect 165 119 166 120 
<< m2 >>
rect 166 119 167 120 
<< m1 >>
rect 181 119 182 120 
<< m1 >>
rect 199 119 200 120 
<< m2 >>
rect 208 119 209 120 
<< m1 >>
rect 211 119 212 120 
<< m1 >>
rect 217 119 218 120 
<< m1 >>
rect 235 119 236 120 
<< m1 >>
rect 244 119 245 120 
<< m1 >>
rect 247 119 248 120 
<< m1 >>
rect 253 119 254 120 
<< m1 >>
rect 255 119 256 120 
<< m1 >>
rect 268 119 269 120 
<< m1 >>
rect 271 119 272 120 
<< m2 >>
rect 272 119 273 120 
<< m1 >>
rect 278 119 279 120 
<< m1 >>
rect 280 119 281 120 
<< m1 >>
rect 283 119 284 120 
<< m1 >>
rect 286 119 287 120 
<< m1 >>
rect 298 119 299 120 
<< m1 >>
rect 334 119 335 120 
<< m1 >>
rect 337 119 338 120 
<< m1 >>
rect 343 119 344 120 
<< m1 >>
rect 345 119 346 120 
<< m1 >>
rect 361 119 362 120 
<< m2 >>
rect 361 119 362 120 
<< m1 >>
rect 366 119 367 120 
<< m1 >>
rect 370 119 371 120 
<< m2 >>
rect 370 119 371 120 
<< m1 >>
rect 373 119 374 120 
<< m1 >>
rect 379 119 380 120 
<< m2 >>
rect 379 119 380 120 
<< m1 >>
rect 381 119 382 120 
<< m1 >>
rect 394 119 395 120 
<< m1 >>
rect 430 119 431 120 
<< m2 >>
rect 431 119 432 120 
<< m1 >>
rect 456 119 457 120 
<< m1 >>
rect 463 119 464 120 
<< m1 >>
rect 478 119 479 120 
<< m1 >>
rect 484 119 485 120 
<< pdiffusion >>
rect 12 120 13 121 
<< pdiffusion >>
rect 13 120 14 121 
<< pdiffusion >>
rect 14 120 15 121 
<< pdiffusion >>
rect 15 120 16 121 
<< m1 >>
rect 16 120 17 121 
<< pdiffusion >>
rect 16 120 17 121 
<< pdiffusion >>
rect 17 120 18 121 
<< m1 >>
rect 19 120 20 121 
<< pdiffusion >>
rect 30 120 31 121 
<< pdiffusion >>
rect 31 120 32 121 
<< pdiffusion >>
rect 32 120 33 121 
<< pdiffusion >>
rect 33 120 34 121 
<< pdiffusion >>
rect 34 120 35 121 
<< pdiffusion >>
rect 35 120 36 121 
<< m1 >>
rect 46 120 47 121 
<< pdiffusion >>
rect 48 120 49 121 
<< pdiffusion >>
rect 49 120 50 121 
<< pdiffusion >>
rect 50 120 51 121 
<< pdiffusion >>
rect 51 120 52 121 
<< pdiffusion >>
rect 52 120 53 121 
<< pdiffusion >>
rect 53 120 54 121 
<< m1 >>
rect 64 120 65 121 
<< pdiffusion >>
rect 66 120 67 121 
<< pdiffusion >>
rect 67 120 68 121 
<< pdiffusion >>
rect 68 120 69 121 
<< pdiffusion >>
rect 69 120 70 121 
<< m1 >>
rect 70 120 71 121 
<< pdiffusion >>
rect 70 120 71 121 
<< pdiffusion >>
rect 71 120 72 121 
<< pdiffusion >>
rect 84 120 85 121 
<< pdiffusion >>
rect 85 120 86 121 
<< pdiffusion >>
rect 86 120 87 121 
<< pdiffusion >>
rect 87 120 88 121 
<< pdiffusion >>
rect 88 120 89 121 
<< pdiffusion >>
rect 89 120 90 121 
<< m1 >>
rect 92 120 93 121 
<< m2 >>
rect 99 120 100 121 
<< m1 >>
rect 100 120 101 121 
<< pdiffusion >>
rect 102 120 103 121 
<< m1 >>
rect 103 120 104 121 
<< pdiffusion >>
rect 103 120 104 121 
<< pdiffusion >>
rect 104 120 105 121 
<< pdiffusion >>
rect 105 120 106 121 
<< m1 >>
rect 106 120 107 121 
<< pdiffusion >>
rect 106 120 107 121 
<< pdiffusion >>
rect 107 120 108 121 
<< m1 >>
rect 109 120 110 121 
<< m1 >>
rect 118 120 119 121 
<< pdiffusion >>
rect 120 120 121 121 
<< pdiffusion >>
rect 121 120 122 121 
<< pdiffusion >>
rect 122 120 123 121 
<< pdiffusion >>
rect 123 120 124 121 
<< m1 >>
rect 124 120 125 121 
<< pdiffusion >>
rect 124 120 125 121 
<< pdiffusion >>
rect 125 120 126 121 
<< m1 >>
rect 129 120 130 121 
<< m1 >>
rect 131 120 132 121 
<< m1 >>
rect 133 120 134 121 
<< m1 >>
rect 136 120 137 121 
<< pdiffusion >>
rect 138 120 139 121 
<< pdiffusion >>
rect 139 120 140 121 
<< pdiffusion >>
rect 140 120 141 121 
<< pdiffusion >>
rect 141 120 142 121 
<< pdiffusion >>
rect 142 120 143 121 
<< pdiffusion >>
rect 143 120 144 121 
<< m1 >>
rect 145 120 146 121 
<< m1 >>
rect 154 120 155 121 
<< pdiffusion >>
rect 156 120 157 121 
<< pdiffusion >>
rect 157 120 158 121 
<< pdiffusion >>
rect 158 120 159 121 
<< pdiffusion >>
rect 159 120 160 121 
<< m1 >>
rect 160 120 161 121 
<< pdiffusion >>
rect 160 120 161 121 
<< pdiffusion >>
rect 161 120 162 121 
<< m1 >>
rect 163 120 164 121 
<< m1 >>
rect 165 120 166 121 
<< m2 >>
rect 166 120 167 121 
<< pdiffusion >>
rect 174 120 175 121 
<< pdiffusion >>
rect 175 120 176 121 
<< pdiffusion >>
rect 176 120 177 121 
<< pdiffusion >>
rect 177 120 178 121 
<< pdiffusion >>
rect 178 120 179 121 
<< pdiffusion >>
rect 179 120 180 121 
<< m1 >>
rect 181 120 182 121 
<< pdiffusion >>
rect 192 120 193 121 
<< pdiffusion >>
rect 193 120 194 121 
<< pdiffusion >>
rect 194 120 195 121 
<< pdiffusion >>
rect 195 120 196 121 
<< pdiffusion >>
rect 196 120 197 121 
<< pdiffusion >>
rect 197 120 198 121 
<< m1 >>
rect 199 120 200 121 
<< m1 >>
rect 208 120 209 121 
<< m2 >>
rect 208 120 209 121 
<< m2c >>
rect 208 120 209 121 
<< m1 >>
rect 208 120 209 121 
<< m2 >>
rect 208 120 209 121 
<< pdiffusion >>
rect 210 120 211 121 
<< m1 >>
rect 211 120 212 121 
<< pdiffusion >>
rect 211 120 212 121 
<< pdiffusion >>
rect 212 120 213 121 
<< pdiffusion >>
rect 213 120 214 121 
<< pdiffusion >>
rect 214 120 215 121 
<< pdiffusion >>
rect 215 120 216 121 
<< m1 >>
rect 217 120 218 121 
<< pdiffusion >>
rect 228 120 229 121 
<< pdiffusion >>
rect 229 120 230 121 
<< pdiffusion >>
rect 230 120 231 121 
<< pdiffusion >>
rect 231 120 232 121 
<< pdiffusion >>
rect 232 120 233 121 
<< pdiffusion >>
rect 233 120 234 121 
<< m1 >>
rect 235 120 236 121 
<< m1 >>
rect 244 120 245 121 
<< pdiffusion >>
rect 246 120 247 121 
<< m1 >>
rect 247 120 248 121 
<< pdiffusion >>
rect 247 120 248 121 
<< pdiffusion >>
rect 248 120 249 121 
<< pdiffusion >>
rect 249 120 250 121 
<< pdiffusion >>
rect 250 120 251 121 
<< pdiffusion >>
rect 251 120 252 121 
<< m1 >>
rect 253 120 254 121 
<< m1 >>
rect 255 120 256 121 
<< pdiffusion >>
rect 264 120 265 121 
<< pdiffusion >>
rect 265 120 266 121 
<< pdiffusion >>
rect 266 120 267 121 
<< pdiffusion >>
rect 267 120 268 121 
<< m1 >>
rect 268 120 269 121 
<< pdiffusion >>
rect 268 120 269 121 
<< pdiffusion >>
rect 269 120 270 121 
<< m1 >>
rect 271 120 272 121 
<< m2 >>
rect 272 120 273 121 
<< m1 >>
rect 278 120 279 121 
<< m1 >>
rect 280 120 281 121 
<< pdiffusion >>
rect 282 120 283 121 
<< m1 >>
rect 283 120 284 121 
<< pdiffusion >>
rect 283 120 284 121 
<< pdiffusion >>
rect 284 120 285 121 
<< pdiffusion >>
rect 285 120 286 121 
<< m1 >>
rect 286 120 287 121 
<< pdiffusion >>
rect 286 120 287 121 
<< pdiffusion >>
rect 287 120 288 121 
<< m1 >>
rect 298 120 299 121 
<< pdiffusion >>
rect 300 120 301 121 
<< pdiffusion >>
rect 301 120 302 121 
<< pdiffusion >>
rect 302 120 303 121 
<< pdiffusion >>
rect 303 120 304 121 
<< pdiffusion >>
rect 304 120 305 121 
<< pdiffusion >>
rect 305 120 306 121 
<< pdiffusion >>
rect 318 120 319 121 
<< pdiffusion >>
rect 319 120 320 121 
<< pdiffusion >>
rect 320 120 321 121 
<< pdiffusion >>
rect 321 120 322 121 
<< pdiffusion >>
rect 322 120 323 121 
<< pdiffusion >>
rect 323 120 324 121 
<< m1 >>
rect 334 120 335 121 
<< pdiffusion >>
rect 336 120 337 121 
<< m1 >>
rect 337 120 338 121 
<< pdiffusion >>
rect 337 120 338 121 
<< pdiffusion >>
rect 338 120 339 121 
<< pdiffusion >>
rect 339 120 340 121 
<< pdiffusion >>
rect 340 120 341 121 
<< pdiffusion >>
rect 341 120 342 121 
<< m1 >>
rect 343 120 344 121 
<< m1 >>
rect 345 120 346 121 
<< pdiffusion >>
rect 354 120 355 121 
<< pdiffusion >>
rect 355 120 356 121 
<< pdiffusion >>
rect 356 120 357 121 
<< pdiffusion >>
rect 357 120 358 121 
<< pdiffusion >>
rect 358 120 359 121 
<< pdiffusion >>
rect 359 120 360 121 
<< m1 >>
rect 361 120 362 121 
<< m2 >>
rect 361 120 362 121 
<< m1 >>
rect 366 120 367 121 
<< m1 >>
rect 370 120 371 121 
<< m2 >>
rect 370 120 371 121 
<< pdiffusion >>
rect 372 120 373 121 
<< m1 >>
rect 373 120 374 121 
<< pdiffusion >>
rect 373 120 374 121 
<< pdiffusion >>
rect 374 120 375 121 
<< pdiffusion >>
rect 375 120 376 121 
<< pdiffusion >>
rect 376 120 377 121 
<< pdiffusion >>
rect 377 120 378 121 
<< m1 >>
rect 379 120 380 121 
<< m2 >>
rect 379 120 380 121 
<< m1 >>
rect 381 120 382 121 
<< pdiffusion >>
rect 390 120 391 121 
<< pdiffusion >>
rect 391 120 392 121 
<< pdiffusion >>
rect 392 120 393 121 
<< pdiffusion >>
rect 393 120 394 121 
<< m1 >>
rect 394 120 395 121 
<< pdiffusion >>
rect 394 120 395 121 
<< pdiffusion >>
rect 395 120 396 121 
<< pdiffusion >>
rect 408 120 409 121 
<< pdiffusion >>
rect 409 120 410 121 
<< pdiffusion >>
rect 410 120 411 121 
<< pdiffusion >>
rect 411 120 412 121 
<< pdiffusion >>
rect 412 120 413 121 
<< pdiffusion >>
rect 413 120 414 121 
<< m1 >>
rect 430 120 431 121 
<< m2 >>
rect 431 120 432 121 
<< pdiffusion >>
rect 444 120 445 121 
<< pdiffusion >>
rect 445 120 446 121 
<< pdiffusion >>
rect 446 120 447 121 
<< pdiffusion >>
rect 447 120 448 121 
<< pdiffusion >>
rect 448 120 449 121 
<< pdiffusion >>
rect 449 120 450 121 
<< m1 >>
rect 456 120 457 121 
<< pdiffusion >>
rect 462 120 463 121 
<< m1 >>
rect 463 120 464 121 
<< pdiffusion >>
rect 463 120 464 121 
<< pdiffusion >>
rect 464 120 465 121 
<< pdiffusion >>
rect 465 120 466 121 
<< pdiffusion >>
rect 466 120 467 121 
<< pdiffusion >>
rect 467 120 468 121 
<< m1 >>
rect 478 120 479 121 
<< m1 >>
rect 484 120 485 121 
<< pdiffusion >>
rect 498 120 499 121 
<< pdiffusion >>
rect 499 120 500 121 
<< pdiffusion >>
rect 500 120 501 121 
<< pdiffusion >>
rect 501 120 502 121 
<< pdiffusion >>
rect 502 120 503 121 
<< pdiffusion >>
rect 503 120 504 121 
<< pdiffusion >>
rect 516 120 517 121 
<< pdiffusion >>
rect 517 120 518 121 
<< pdiffusion >>
rect 518 120 519 121 
<< pdiffusion >>
rect 519 120 520 121 
<< pdiffusion >>
rect 520 120 521 121 
<< pdiffusion >>
rect 521 120 522 121 
<< pdiffusion >>
rect 12 121 13 122 
<< pdiffusion >>
rect 13 121 14 122 
<< pdiffusion >>
rect 14 121 15 122 
<< pdiffusion >>
rect 15 121 16 122 
<< pdiffusion >>
rect 16 121 17 122 
<< pdiffusion >>
rect 17 121 18 122 
<< m1 >>
rect 19 121 20 122 
<< pdiffusion >>
rect 30 121 31 122 
<< pdiffusion >>
rect 31 121 32 122 
<< pdiffusion >>
rect 32 121 33 122 
<< pdiffusion >>
rect 33 121 34 122 
<< pdiffusion >>
rect 34 121 35 122 
<< pdiffusion >>
rect 35 121 36 122 
<< m1 >>
rect 46 121 47 122 
<< pdiffusion >>
rect 48 121 49 122 
<< pdiffusion >>
rect 49 121 50 122 
<< pdiffusion >>
rect 50 121 51 122 
<< pdiffusion >>
rect 51 121 52 122 
<< pdiffusion >>
rect 52 121 53 122 
<< pdiffusion >>
rect 53 121 54 122 
<< m1 >>
rect 64 121 65 122 
<< pdiffusion >>
rect 66 121 67 122 
<< pdiffusion >>
rect 67 121 68 122 
<< pdiffusion >>
rect 68 121 69 122 
<< pdiffusion >>
rect 69 121 70 122 
<< pdiffusion >>
rect 70 121 71 122 
<< pdiffusion >>
rect 71 121 72 122 
<< pdiffusion >>
rect 84 121 85 122 
<< pdiffusion >>
rect 85 121 86 122 
<< pdiffusion >>
rect 86 121 87 122 
<< pdiffusion >>
rect 87 121 88 122 
<< pdiffusion >>
rect 88 121 89 122 
<< pdiffusion >>
rect 89 121 90 122 
<< m1 >>
rect 92 121 93 122 
<< m2 >>
rect 99 121 100 122 
<< m1 >>
rect 100 121 101 122 
<< pdiffusion >>
rect 102 121 103 122 
<< pdiffusion >>
rect 103 121 104 122 
<< pdiffusion >>
rect 104 121 105 122 
<< pdiffusion >>
rect 105 121 106 122 
<< pdiffusion >>
rect 106 121 107 122 
<< pdiffusion >>
rect 107 121 108 122 
<< m1 >>
rect 109 121 110 122 
<< m1 >>
rect 118 121 119 122 
<< pdiffusion >>
rect 120 121 121 122 
<< pdiffusion >>
rect 121 121 122 122 
<< pdiffusion >>
rect 122 121 123 122 
<< pdiffusion >>
rect 123 121 124 122 
<< pdiffusion >>
rect 124 121 125 122 
<< pdiffusion >>
rect 125 121 126 122 
<< m1 >>
rect 129 121 130 122 
<< m1 >>
rect 131 121 132 122 
<< m1 >>
rect 133 121 134 122 
<< m1 >>
rect 136 121 137 122 
<< pdiffusion >>
rect 138 121 139 122 
<< pdiffusion >>
rect 139 121 140 122 
<< pdiffusion >>
rect 140 121 141 122 
<< pdiffusion >>
rect 141 121 142 122 
<< pdiffusion >>
rect 142 121 143 122 
<< pdiffusion >>
rect 143 121 144 122 
<< m1 >>
rect 145 121 146 122 
<< m1 >>
rect 154 121 155 122 
<< pdiffusion >>
rect 156 121 157 122 
<< pdiffusion >>
rect 157 121 158 122 
<< pdiffusion >>
rect 158 121 159 122 
<< pdiffusion >>
rect 159 121 160 122 
<< pdiffusion >>
rect 160 121 161 122 
<< pdiffusion >>
rect 161 121 162 122 
<< m1 >>
rect 163 121 164 122 
<< m1 >>
rect 165 121 166 122 
<< m2 >>
rect 166 121 167 122 
<< pdiffusion >>
rect 174 121 175 122 
<< pdiffusion >>
rect 175 121 176 122 
<< pdiffusion >>
rect 176 121 177 122 
<< pdiffusion >>
rect 177 121 178 122 
<< pdiffusion >>
rect 178 121 179 122 
<< pdiffusion >>
rect 179 121 180 122 
<< m1 >>
rect 181 121 182 122 
<< pdiffusion >>
rect 192 121 193 122 
<< pdiffusion >>
rect 193 121 194 122 
<< pdiffusion >>
rect 194 121 195 122 
<< pdiffusion >>
rect 195 121 196 122 
<< pdiffusion >>
rect 196 121 197 122 
<< pdiffusion >>
rect 197 121 198 122 
<< m1 >>
rect 199 121 200 122 
<< m1 >>
rect 208 121 209 122 
<< pdiffusion >>
rect 210 121 211 122 
<< pdiffusion >>
rect 211 121 212 122 
<< pdiffusion >>
rect 212 121 213 122 
<< pdiffusion >>
rect 213 121 214 122 
<< pdiffusion >>
rect 214 121 215 122 
<< pdiffusion >>
rect 215 121 216 122 
<< m1 >>
rect 217 121 218 122 
<< pdiffusion >>
rect 228 121 229 122 
<< pdiffusion >>
rect 229 121 230 122 
<< pdiffusion >>
rect 230 121 231 122 
<< pdiffusion >>
rect 231 121 232 122 
<< pdiffusion >>
rect 232 121 233 122 
<< pdiffusion >>
rect 233 121 234 122 
<< m1 >>
rect 235 121 236 122 
<< m1 >>
rect 244 121 245 122 
<< pdiffusion >>
rect 246 121 247 122 
<< pdiffusion >>
rect 247 121 248 122 
<< pdiffusion >>
rect 248 121 249 122 
<< pdiffusion >>
rect 249 121 250 122 
<< pdiffusion >>
rect 250 121 251 122 
<< pdiffusion >>
rect 251 121 252 122 
<< m1 >>
rect 253 121 254 122 
<< m1 >>
rect 255 121 256 122 
<< pdiffusion >>
rect 264 121 265 122 
<< pdiffusion >>
rect 265 121 266 122 
<< pdiffusion >>
rect 266 121 267 122 
<< pdiffusion >>
rect 267 121 268 122 
<< pdiffusion >>
rect 268 121 269 122 
<< pdiffusion >>
rect 269 121 270 122 
<< m1 >>
rect 271 121 272 122 
<< m2 >>
rect 272 121 273 122 
<< m1 >>
rect 278 121 279 122 
<< m1 >>
rect 280 121 281 122 
<< pdiffusion >>
rect 282 121 283 122 
<< pdiffusion >>
rect 283 121 284 122 
<< pdiffusion >>
rect 284 121 285 122 
<< pdiffusion >>
rect 285 121 286 122 
<< pdiffusion >>
rect 286 121 287 122 
<< pdiffusion >>
rect 287 121 288 122 
<< m1 >>
rect 298 121 299 122 
<< pdiffusion >>
rect 300 121 301 122 
<< pdiffusion >>
rect 301 121 302 122 
<< pdiffusion >>
rect 302 121 303 122 
<< pdiffusion >>
rect 303 121 304 122 
<< pdiffusion >>
rect 304 121 305 122 
<< pdiffusion >>
rect 305 121 306 122 
<< pdiffusion >>
rect 318 121 319 122 
<< pdiffusion >>
rect 319 121 320 122 
<< pdiffusion >>
rect 320 121 321 122 
<< pdiffusion >>
rect 321 121 322 122 
<< pdiffusion >>
rect 322 121 323 122 
<< pdiffusion >>
rect 323 121 324 122 
<< m1 >>
rect 334 121 335 122 
<< pdiffusion >>
rect 336 121 337 122 
<< pdiffusion >>
rect 337 121 338 122 
<< pdiffusion >>
rect 338 121 339 122 
<< pdiffusion >>
rect 339 121 340 122 
<< pdiffusion >>
rect 340 121 341 122 
<< pdiffusion >>
rect 341 121 342 122 
<< m1 >>
rect 343 121 344 122 
<< m1 >>
rect 345 121 346 122 
<< pdiffusion >>
rect 354 121 355 122 
<< pdiffusion >>
rect 355 121 356 122 
<< pdiffusion >>
rect 356 121 357 122 
<< pdiffusion >>
rect 357 121 358 122 
<< pdiffusion >>
rect 358 121 359 122 
<< pdiffusion >>
rect 359 121 360 122 
<< m1 >>
rect 361 121 362 122 
<< m2 >>
rect 361 121 362 122 
<< m1 >>
rect 366 121 367 122 
<< m1 >>
rect 370 121 371 122 
<< m2 >>
rect 370 121 371 122 
<< pdiffusion >>
rect 372 121 373 122 
<< pdiffusion >>
rect 373 121 374 122 
<< pdiffusion >>
rect 374 121 375 122 
<< pdiffusion >>
rect 375 121 376 122 
<< pdiffusion >>
rect 376 121 377 122 
<< pdiffusion >>
rect 377 121 378 122 
<< m1 >>
rect 379 121 380 122 
<< m2 >>
rect 379 121 380 122 
<< m1 >>
rect 381 121 382 122 
<< pdiffusion >>
rect 390 121 391 122 
<< pdiffusion >>
rect 391 121 392 122 
<< pdiffusion >>
rect 392 121 393 122 
<< pdiffusion >>
rect 393 121 394 122 
<< pdiffusion >>
rect 394 121 395 122 
<< pdiffusion >>
rect 395 121 396 122 
<< pdiffusion >>
rect 408 121 409 122 
<< pdiffusion >>
rect 409 121 410 122 
<< pdiffusion >>
rect 410 121 411 122 
<< pdiffusion >>
rect 411 121 412 122 
<< pdiffusion >>
rect 412 121 413 122 
<< pdiffusion >>
rect 413 121 414 122 
<< m1 >>
rect 430 121 431 122 
<< m2 >>
rect 431 121 432 122 
<< pdiffusion >>
rect 444 121 445 122 
<< pdiffusion >>
rect 445 121 446 122 
<< pdiffusion >>
rect 446 121 447 122 
<< pdiffusion >>
rect 447 121 448 122 
<< pdiffusion >>
rect 448 121 449 122 
<< pdiffusion >>
rect 449 121 450 122 
<< m1 >>
rect 456 121 457 122 
<< pdiffusion >>
rect 462 121 463 122 
<< pdiffusion >>
rect 463 121 464 122 
<< pdiffusion >>
rect 464 121 465 122 
<< pdiffusion >>
rect 465 121 466 122 
<< pdiffusion >>
rect 466 121 467 122 
<< pdiffusion >>
rect 467 121 468 122 
<< m1 >>
rect 478 121 479 122 
<< m1 >>
rect 484 121 485 122 
<< pdiffusion >>
rect 498 121 499 122 
<< pdiffusion >>
rect 499 121 500 122 
<< pdiffusion >>
rect 500 121 501 122 
<< pdiffusion >>
rect 501 121 502 122 
<< pdiffusion >>
rect 502 121 503 122 
<< pdiffusion >>
rect 503 121 504 122 
<< pdiffusion >>
rect 516 121 517 122 
<< pdiffusion >>
rect 517 121 518 122 
<< pdiffusion >>
rect 518 121 519 122 
<< pdiffusion >>
rect 519 121 520 122 
<< pdiffusion >>
rect 520 121 521 122 
<< pdiffusion >>
rect 521 121 522 122 
<< pdiffusion >>
rect 12 122 13 123 
<< pdiffusion >>
rect 13 122 14 123 
<< pdiffusion >>
rect 14 122 15 123 
<< pdiffusion >>
rect 15 122 16 123 
<< pdiffusion >>
rect 16 122 17 123 
<< pdiffusion >>
rect 17 122 18 123 
<< m1 >>
rect 19 122 20 123 
<< pdiffusion >>
rect 30 122 31 123 
<< pdiffusion >>
rect 31 122 32 123 
<< pdiffusion >>
rect 32 122 33 123 
<< pdiffusion >>
rect 33 122 34 123 
<< pdiffusion >>
rect 34 122 35 123 
<< pdiffusion >>
rect 35 122 36 123 
<< m1 >>
rect 46 122 47 123 
<< pdiffusion >>
rect 48 122 49 123 
<< pdiffusion >>
rect 49 122 50 123 
<< pdiffusion >>
rect 50 122 51 123 
<< pdiffusion >>
rect 51 122 52 123 
<< pdiffusion >>
rect 52 122 53 123 
<< pdiffusion >>
rect 53 122 54 123 
<< m1 >>
rect 64 122 65 123 
<< pdiffusion >>
rect 66 122 67 123 
<< pdiffusion >>
rect 67 122 68 123 
<< pdiffusion >>
rect 68 122 69 123 
<< pdiffusion >>
rect 69 122 70 123 
<< pdiffusion >>
rect 70 122 71 123 
<< pdiffusion >>
rect 71 122 72 123 
<< pdiffusion >>
rect 84 122 85 123 
<< pdiffusion >>
rect 85 122 86 123 
<< pdiffusion >>
rect 86 122 87 123 
<< pdiffusion >>
rect 87 122 88 123 
<< pdiffusion >>
rect 88 122 89 123 
<< pdiffusion >>
rect 89 122 90 123 
<< m1 >>
rect 92 122 93 123 
<< m2 >>
rect 99 122 100 123 
<< m1 >>
rect 100 122 101 123 
<< pdiffusion >>
rect 102 122 103 123 
<< pdiffusion >>
rect 103 122 104 123 
<< pdiffusion >>
rect 104 122 105 123 
<< pdiffusion >>
rect 105 122 106 123 
<< pdiffusion >>
rect 106 122 107 123 
<< pdiffusion >>
rect 107 122 108 123 
<< m1 >>
rect 109 122 110 123 
<< m1 >>
rect 118 122 119 123 
<< pdiffusion >>
rect 120 122 121 123 
<< pdiffusion >>
rect 121 122 122 123 
<< pdiffusion >>
rect 122 122 123 123 
<< pdiffusion >>
rect 123 122 124 123 
<< pdiffusion >>
rect 124 122 125 123 
<< pdiffusion >>
rect 125 122 126 123 
<< m1 >>
rect 129 122 130 123 
<< m1 >>
rect 131 122 132 123 
<< m1 >>
rect 133 122 134 123 
<< m1 >>
rect 136 122 137 123 
<< pdiffusion >>
rect 138 122 139 123 
<< pdiffusion >>
rect 139 122 140 123 
<< pdiffusion >>
rect 140 122 141 123 
<< pdiffusion >>
rect 141 122 142 123 
<< pdiffusion >>
rect 142 122 143 123 
<< pdiffusion >>
rect 143 122 144 123 
<< m1 >>
rect 145 122 146 123 
<< m1 >>
rect 154 122 155 123 
<< pdiffusion >>
rect 156 122 157 123 
<< pdiffusion >>
rect 157 122 158 123 
<< pdiffusion >>
rect 158 122 159 123 
<< pdiffusion >>
rect 159 122 160 123 
<< pdiffusion >>
rect 160 122 161 123 
<< pdiffusion >>
rect 161 122 162 123 
<< m1 >>
rect 163 122 164 123 
<< m1 >>
rect 165 122 166 123 
<< m2 >>
rect 166 122 167 123 
<< pdiffusion >>
rect 174 122 175 123 
<< pdiffusion >>
rect 175 122 176 123 
<< pdiffusion >>
rect 176 122 177 123 
<< pdiffusion >>
rect 177 122 178 123 
<< pdiffusion >>
rect 178 122 179 123 
<< pdiffusion >>
rect 179 122 180 123 
<< m1 >>
rect 181 122 182 123 
<< pdiffusion >>
rect 192 122 193 123 
<< pdiffusion >>
rect 193 122 194 123 
<< pdiffusion >>
rect 194 122 195 123 
<< pdiffusion >>
rect 195 122 196 123 
<< pdiffusion >>
rect 196 122 197 123 
<< pdiffusion >>
rect 197 122 198 123 
<< m1 >>
rect 199 122 200 123 
<< m1 >>
rect 208 122 209 123 
<< pdiffusion >>
rect 210 122 211 123 
<< pdiffusion >>
rect 211 122 212 123 
<< pdiffusion >>
rect 212 122 213 123 
<< pdiffusion >>
rect 213 122 214 123 
<< pdiffusion >>
rect 214 122 215 123 
<< pdiffusion >>
rect 215 122 216 123 
<< m1 >>
rect 217 122 218 123 
<< pdiffusion >>
rect 228 122 229 123 
<< pdiffusion >>
rect 229 122 230 123 
<< pdiffusion >>
rect 230 122 231 123 
<< pdiffusion >>
rect 231 122 232 123 
<< pdiffusion >>
rect 232 122 233 123 
<< pdiffusion >>
rect 233 122 234 123 
<< m1 >>
rect 235 122 236 123 
<< m1 >>
rect 244 122 245 123 
<< pdiffusion >>
rect 246 122 247 123 
<< pdiffusion >>
rect 247 122 248 123 
<< pdiffusion >>
rect 248 122 249 123 
<< pdiffusion >>
rect 249 122 250 123 
<< pdiffusion >>
rect 250 122 251 123 
<< pdiffusion >>
rect 251 122 252 123 
<< m1 >>
rect 253 122 254 123 
<< m1 >>
rect 255 122 256 123 
<< pdiffusion >>
rect 264 122 265 123 
<< pdiffusion >>
rect 265 122 266 123 
<< pdiffusion >>
rect 266 122 267 123 
<< pdiffusion >>
rect 267 122 268 123 
<< pdiffusion >>
rect 268 122 269 123 
<< pdiffusion >>
rect 269 122 270 123 
<< m1 >>
rect 271 122 272 123 
<< m2 >>
rect 272 122 273 123 
<< m1 >>
rect 278 122 279 123 
<< m1 >>
rect 280 122 281 123 
<< pdiffusion >>
rect 282 122 283 123 
<< pdiffusion >>
rect 283 122 284 123 
<< pdiffusion >>
rect 284 122 285 123 
<< pdiffusion >>
rect 285 122 286 123 
<< pdiffusion >>
rect 286 122 287 123 
<< pdiffusion >>
rect 287 122 288 123 
<< m1 >>
rect 298 122 299 123 
<< pdiffusion >>
rect 300 122 301 123 
<< pdiffusion >>
rect 301 122 302 123 
<< pdiffusion >>
rect 302 122 303 123 
<< pdiffusion >>
rect 303 122 304 123 
<< pdiffusion >>
rect 304 122 305 123 
<< pdiffusion >>
rect 305 122 306 123 
<< pdiffusion >>
rect 318 122 319 123 
<< pdiffusion >>
rect 319 122 320 123 
<< pdiffusion >>
rect 320 122 321 123 
<< pdiffusion >>
rect 321 122 322 123 
<< pdiffusion >>
rect 322 122 323 123 
<< pdiffusion >>
rect 323 122 324 123 
<< m1 >>
rect 334 122 335 123 
<< pdiffusion >>
rect 336 122 337 123 
<< pdiffusion >>
rect 337 122 338 123 
<< pdiffusion >>
rect 338 122 339 123 
<< pdiffusion >>
rect 339 122 340 123 
<< pdiffusion >>
rect 340 122 341 123 
<< pdiffusion >>
rect 341 122 342 123 
<< m1 >>
rect 343 122 344 123 
<< m1 >>
rect 345 122 346 123 
<< pdiffusion >>
rect 354 122 355 123 
<< pdiffusion >>
rect 355 122 356 123 
<< pdiffusion >>
rect 356 122 357 123 
<< pdiffusion >>
rect 357 122 358 123 
<< pdiffusion >>
rect 358 122 359 123 
<< pdiffusion >>
rect 359 122 360 123 
<< m1 >>
rect 361 122 362 123 
<< m2 >>
rect 361 122 362 123 
<< m1 >>
rect 366 122 367 123 
<< m1 >>
rect 370 122 371 123 
<< m2 >>
rect 370 122 371 123 
<< pdiffusion >>
rect 372 122 373 123 
<< pdiffusion >>
rect 373 122 374 123 
<< pdiffusion >>
rect 374 122 375 123 
<< pdiffusion >>
rect 375 122 376 123 
<< pdiffusion >>
rect 376 122 377 123 
<< pdiffusion >>
rect 377 122 378 123 
<< m1 >>
rect 379 122 380 123 
<< m2 >>
rect 379 122 380 123 
<< m1 >>
rect 381 122 382 123 
<< pdiffusion >>
rect 390 122 391 123 
<< pdiffusion >>
rect 391 122 392 123 
<< pdiffusion >>
rect 392 122 393 123 
<< pdiffusion >>
rect 393 122 394 123 
<< pdiffusion >>
rect 394 122 395 123 
<< pdiffusion >>
rect 395 122 396 123 
<< pdiffusion >>
rect 408 122 409 123 
<< pdiffusion >>
rect 409 122 410 123 
<< pdiffusion >>
rect 410 122 411 123 
<< pdiffusion >>
rect 411 122 412 123 
<< pdiffusion >>
rect 412 122 413 123 
<< pdiffusion >>
rect 413 122 414 123 
<< m1 >>
rect 430 122 431 123 
<< m2 >>
rect 431 122 432 123 
<< pdiffusion >>
rect 444 122 445 123 
<< pdiffusion >>
rect 445 122 446 123 
<< pdiffusion >>
rect 446 122 447 123 
<< pdiffusion >>
rect 447 122 448 123 
<< pdiffusion >>
rect 448 122 449 123 
<< pdiffusion >>
rect 449 122 450 123 
<< m1 >>
rect 456 122 457 123 
<< pdiffusion >>
rect 462 122 463 123 
<< pdiffusion >>
rect 463 122 464 123 
<< pdiffusion >>
rect 464 122 465 123 
<< pdiffusion >>
rect 465 122 466 123 
<< pdiffusion >>
rect 466 122 467 123 
<< pdiffusion >>
rect 467 122 468 123 
<< m1 >>
rect 478 122 479 123 
<< m1 >>
rect 484 122 485 123 
<< pdiffusion >>
rect 498 122 499 123 
<< pdiffusion >>
rect 499 122 500 123 
<< pdiffusion >>
rect 500 122 501 123 
<< pdiffusion >>
rect 501 122 502 123 
<< pdiffusion >>
rect 502 122 503 123 
<< pdiffusion >>
rect 503 122 504 123 
<< pdiffusion >>
rect 516 122 517 123 
<< pdiffusion >>
rect 517 122 518 123 
<< pdiffusion >>
rect 518 122 519 123 
<< pdiffusion >>
rect 519 122 520 123 
<< pdiffusion >>
rect 520 122 521 123 
<< pdiffusion >>
rect 521 122 522 123 
<< pdiffusion >>
rect 12 123 13 124 
<< pdiffusion >>
rect 13 123 14 124 
<< pdiffusion >>
rect 14 123 15 124 
<< pdiffusion >>
rect 15 123 16 124 
<< pdiffusion >>
rect 16 123 17 124 
<< pdiffusion >>
rect 17 123 18 124 
<< m1 >>
rect 19 123 20 124 
<< pdiffusion >>
rect 30 123 31 124 
<< pdiffusion >>
rect 31 123 32 124 
<< pdiffusion >>
rect 32 123 33 124 
<< pdiffusion >>
rect 33 123 34 124 
<< pdiffusion >>
rect 34 123 35 124 
<< pdiffusion >>
rect 35 123 36 124 
<< m1 >>
rect 46 123 47 124 
<< pdiffusion >>
rect 48 123 49 124 
<< pdiffusion >>
rect 49 123 50 124 
<< pdiffusion >>
rect 50 123 51 124 
<< pdiffusion >>
rect 51 123 52 124 
<< pdiffusion >>
rect 52 123 53 124 
<< pdiffusion >>
rect 53 123 54 124 
<< m1 >>
rect 64 123 65 124 
<< pdiffusion >>
rect 66 123 67 124 
<< pdiffusion >>
rect 67 123 68 124 
<< pdiffusion >>
rect 68 123 69 124 
<< pdiffusion >>
rect 69 123 70 124 
<< pdiffusion >>
rect 70 123 71 124 
<< pdiffusion >>
rect 71 123 72 124 
<< pdiffusion >>
rect 84 123 85 124 
<< pdiffusion >>
rect 85 123 86 124 
<< pdiffusion >>
rect 86 123 87 124 
<< pdiffusion >>
rect 87 123 88 124 
<< pdiffusion >>
rect 88 123 89 124 
<< pdiffusion >>
rect 89 123 90 124 
<< m1 >>
rect 92 123 93 124 
<< m2 >>
rect 99 123 100 124 
<< m1 >>
rect 100 123 101 124 
<< pdiffusion >>
rect 102 123 103 124 
<< pdiffusion >>
rect 103 123 104 124 
<< pdiffusion >>
rect 104 123 105 124 
<< pdiffusion >>
rect 105 123 106 124 
<< pdiffusion >>
rect 106 123 107 124 
<< pdiffusion >>
rect 107 123 108 124 
<< m1 >>
rect 109 123 110 124 
<< m1 >>
rect 118 123 119 124 
<< pdiffusion >>
rect 120 123 121 124 
<< pdiffusion >>
rect 121 123 122 124 
<< pdiffusion >>
rect 122 123 123 124 
<< pdiffusion >>
rect 123 123 124 124 
<< pdiffusion >>
rect 124 123 125 124 
<< pdiffusion >>
rect 125 123 126 124 
<< m1 >>
rect 129 123 130 124 
<< m1 >>
rect 131 123 132 124 
<< m1 >>
rect 133 123 134 124 
<< m1 >>
rect 136 123 137 124 
<< pdiffusion >>
rect 138 123 139 124 
<< pdiffusion >>
rect 139 123 140 124 
<< pdiffusion >>
rect 140 123 141 124 
<< pdiffusion >>
rect 141 123 142 124 
<< pdiffusion >>
rect 142 123 143 124 
<< pdiffusion >>
rect 143 123 144 124 
<< m1 >>
rect 145 123 146 124 
<< m1 >>
rect 154 123 155 124 
<< pdiffusion >>
rect 156 123 157 124 
<< pdiffusion >>
rect 157 123 158 124 
<< pdiffusion >>
rect 158 123 159 124 
<< pdiffusion >>
rect 159 123 160 124 
<< pdiffusion >>
rect 160 123 161 124 
<< pdiffusion >>
rect 161 123 162 124 
<< m1 >>
rect 163 123 164 124 
<< m1 >>
rect 165 123 166 124 
<< m2 >>
rect 166 123 167 124 
<< pdiffusion >>
rect 174 123 175 124 
<< pdiffusion >>
rect 175 123 176 124 
<< pdiffusion >>
rect 176 123 177 124 
<< pdiffusion >>
rect 177 123 178 124 
<< pdiffusion >>
rect 178 123 179 124 
<< pdiffusion >>
rect 179 123 180 124 
<< m1 >>
rect 181 123 182 124 
<< pdiffusion >>
rect 192 123 193 124 
<< pdiffusion >>
rect 193 123 194 124 
<< pdiffusion >>
rect 194 123 195 124 
<< pdiffusion >>
rect 195 123 196 124 
<< pdiffusion >>
rect 196 123 197 124 
<< pdiffusion >>
rect 197 123 198 124 
<< m1 >>
rect 199 123 200 124 
<< m1 >>
rect 208 123 209 124 
<< pdiffusion >>
rect 210 123 211 124 
<< pdiffusion >>
rect 211 123 212 124 
<< pdiffusion >>
rect 212 123 213 124 
<< pdiffusion >>
rect 213 123 214 124 
<< pdiffusion >>
rect 214 123 215 124 
<< pdiffusion >>
rect 215 123 216 124 
<< m1 >>
rect 217 123 218 124 
<< pdiffusion >>
rect 228 123 229 124 
<< pdiffusion >>
rect 229 123 230 124 
<< pdiffusion >>
rect 230 123 231 124 
<< pdiffusion >>
rect 231 123 232 124 
<< pdiffusion >>
rect 232 123 233 124 
<< pdiffusion >>
rect 233 123 234 124 
<< m1 >>
rect 235 123 236 124 
<< m1 >>
rect 244 123 245 124 
<< pdiffusion >>
rect 246 123 247 124 
<< pdiffusion >>
rect 247 123 248 124 
<< pdiffusion >>
rect 248 123 249 124 
<< pdiffusion >>
rect 249 123 250 124 
<< pdiffusion >>
rect 250 123 251 124 
<< pdiffusion >>
rect 251 123 252 124 
<< m1 >>
rect 253 123 254 124 
<< m1 >>
rect 255 123 256 124 
<< pdiffusion >>
rect 264 123 265 124 
<< pdiffusion >>
rect 265 123 266 124 
<< pdiffusion >>
rect 266 123 267 124 
<< pdiffusion >>
rect 267 123 268 124 
<< pdiffusion >>
rect 268 123 269 124 
<< pdiffusion >>
rect 269 123 270 124 
<< m1 >>
rect 271 123 272 124 
<< m2 >>
rect 272 123 273 124 
<< m1 >>
rect 278 123 279 124 
<< m1 >>
rect 280 123 281 124 
<< pdiffusion >>
rect 282 123 283 124 
<< pdiffusion >>
rect 283 123 284 124 
<< pdiffusion >>
rect 284 123 285 124 
<< pdiffusion >>
rect 285 123 286 124 
<< pdiffusion >>
rect 286 123 287 124 
<< pdiffusion >>
rect 287 123 288 124 
<< m1 >>
rect 298 123 299 124 
<< pdiffusion >>
rect 300 123 301 124 
<< pdiffusion >>
rect 301 123 302 124 
<< pdiffusion >>
rect 302 123 303 124 
<< pdiffusion >>
rect 303 123 304 124 
<< pdiffusion >>
rect 304 123 305 124 
<< pdiffusion >>
rect 305 123 306 124 
<< pdiffusion >>
rect 318 123 319 124 
<< pdiffusion >>
rect 319 123 320 124 
<< pdiffusion >>
rect 320 123 321 124 
<< pdiffusion >>
rect 321 123 322 124 
<< pdiffusion >>
rect 322 123 323 124 
<< pdiffusion >>
rect 323 123 324 124 
<< m1 >>
rect 334 123 335 124 
<< pdiffusion >>
rect 336 123 337 124 
<< pdiffusion >>
rect 337 123 338 124 
<< pdiffusion >>
rect 338 123 339 124 
<< pdiffusion >>
rect 339 123 340 124 
<< pdiffusion >>
rect 340 123 341 124 
<< pdiffusion >>
rect 341 123 342 124 
<< m1 >>
rect 343 123 344 124 
<< m1 >>
rect 345 123 346 124 
<< pdiffusion >>
rect 354 123 355 124 
<< pdiffusion >>
rect 355 123 356 124 
<< pdiffusion >>
rect 356 123 357 124 
<< pdiffusion >>
rect 357 123 358 124 
<< pdiffusion >>
rect 358 123 359 124 
<< pdiffusion >>
rect 359 123 360 124 
<< m1 >>
rect 361 123 362 124 
<< m2 >>
rect 361 123 362 124 
<< m1 >>
rect 366 123 367 124 
<< m1 >>
rect 370 123 371 124 
<< m2 >>
rect 370 123 371 124 
<< pdiffusion >>
rect 372 123 373 124 
<< pdiffusion >>
rect 373 123 374 124 
<< pdiffusion >>
rect 374 123 375 124 
<< pdiffusion >>
rect 375 123 376 124 
<< pdiffusion >>
rect 376 123 377 124 
<< pdiffusion >>
rect 377 123 378 124 
<< m1 >>
rect 379 123 380 124 
<< m2 >>
rect 379 123 380 124 
<< m1 >>
rect 381 123 382 124 
<< pdiffusion >>
rect 390 123 391 124 
<< pdiffusion >>
rect 391 123 392 124 
<< pdiffusion >>
rect 392 123 393 124 
<< pdiffusion >>
rect 393 123 394 124 
<< pdiffusion >>
rect 394 123 395 124 
<< pdiffusion >>
rect 395 123 396 124 
<< pdiffusion >>
rect 408 123 409 124 
<< pdiffusion >>
rect 409 123 410 124 
<< pdiffusion >>
rect 410 123 411 124 
<< pdiffusion >>
rect 411 123 412 124 
<< pdiffusion >>
rect 412 123 413 124 
<< pdiffusion >>
rect 413 123 414 124 
<< m1 >>
rect 430 123 431 124 
<< m2 >>
rect 431 123 432 124 
<< pdiffusion >>
rect 444 123 445 124 
<< pdiffusion >>
rect 445 123 446 124 
<< pdiffusion >>
rect 446 123 447 124 
<< pdiffusion >>
rect 447 123 448 124 
<< pdiffusion >>
rect 448 123 449 124 
<< pdiffusion >>
rect 449 123 450 124 
<< m1 >>
rect 456 123 457 124 
<< pdiffusion >>
rect 462 123 463 124 
<< pdiffusion >>
rect 463 123 464 124 
<< pdiffusion >>
rect 464 123 465 124 
<< pdiffusion >>
rect 465 123 466 124 
<< pdiffusion >>
rect 466 123 467 124 
<< pdiffusion >>
rect 467 123 468 124 
<< m1 >>
rect 478 123 479 124 
<< m1 >>
rect 484 123 485 124 
<< pdiffusion >>
rect 498 123 499 124 
<< pdiffusion >>
rect 499 123 500 124 
<< pdiffusion >>
rect 500 123 501 124 
<< pdiffusion >>
rect 501 123 502 124 
<< pdiffusion >>
rect 502 123 503 124 
<< pdiffusion >>
rect 503 123 504 124 
<< pdiffusion >>
rect 516 123 517 124 
<< pdiffusion >>
rect 517 123 518 124 
<< pdiffusion >>
rect 518 123 519 124 
<< pdiffusion >>
rect 519 123 520 124 
<< pdiffusion >>
rect 520 123 521 124 
<< pdiffusion >>
rect 521 123 522 124 
<< pdiffusion >>
rect 12 124 13 125 
<< pdiffusion >>
rect 13 124 14 125 
<< pdiffusion >>
rect 14 124 15 125 
<< pdiffusion >>
rect 15 124 16 125 
<< pdiffusion >>
rect 16 124 17 125 
<< pdiffusion >>
rect 17 124 18 125 
<< m1 >>
rect 19 124 20 125 
<< pdiffusion >>
rect 30 124 31 125 
<< pdiffusion >>
rect 31 124 32 125 
<< pdiffusion >>
rect 32 124 33 125 
<< pdiffusion >>
rect 33 124 34 125 
<< pdiffusion >>
rect 34 124 35 125 
<< pdiffusion >>
rect 35 124 36 125 
<< m1 >>
rect 46 124 47 125 
<< pdiffusion >>
rect 48 124 49 125 
<< pdiffusion >>
rect 49 124 50 125 
<< pdiffusion >>
rect 50 124 51 125 
<< pdiffusion >>
rect 51 124 52 125 
<< pdiffusion >>
rect 52 124 53 125 
<< pdiffusion >>
rect 53 124 54 125 
<< m1 >>
rect 64 124 65 125 
<< pdiffusion >>
rect 66 124 67 125 
<< pdiffusion >>
rect 67 124 68 125 
<< pdiffusion >>
rect 68 124 69 125 
<< pdiffusion >>
rect 69 124 70 125 
<< pdiffusion >>
rect 70 124 71 125 
<< pdiffusion >>
rect 71 124 72 125 
<< pdiffusion >>
rect 84 124 85 125 
<< pdiffusion >>
rect 85 124 86 125 
<< pdiffusion >>
rect 86 124 87 125 
<< pdiffusion >>
rect 87 124 88 125 
<< pdiffusion >>
rect 88 124 89 125 
<< pdiffusion >>
rect 89 124 90 125 
<< m1 >>
rect 92 124 93 125 
<< m2 >>
rect 99 124 100 125 
<< m1 >>
rect 100 124 101 125 
<< pdiffusion >>
rect 102 124 103 125 
<< pdiffusion >>
rect 103 124 104 125 
<< pdiffusion >>
rect 104 124 105 125 
<< pdiffusion >>
rect 105 124 106 125 
<< pdiffusion >>
rect 106 124 107 125 
<< pdiffusion >>
rect 107 124 108 125 
<< m1 >>
rect 109 124 110 125 
<< m1 >>
rect 118 124 119 125 
<< pdiffusion >>
rect 120 124 121 125 
<< pdiffusion >>
rect 121 124 122 125 
<< pdiffusion >>
rect 122 124 123 125 
<< pdiffusion >>
rect 123 124 124 125 
<< pdiffusion >>
rect 124 124 125 125 
<< pdiffusion >>
rect 125 124 126 125 
<< m1 >>
rect 129 124 130 125 
<< m1 >>
rect 131 124 132 125 
<< m1 >>
rect 133 124 134 125 
<< m1 >>
rect 136 124 137 125 
<< pdiffusion >>
rect 138 124 139 125 
<< pdiffusion >>
rect 139 124 140 125 
<< pdiffusion >>
rect 140 124 141 125 
<< pdiffusion >>
rect 141 124 142 125 
<< pdiffusion >>
rect 142 124 143 125 
<< pdiffusion >>
rect 143 124 144 125 
<< m1 >>
rect 145 124 146 125 
<< m1 >>
rect 154 124 155 125 
<< pdiffusion >>
rect 156 124 157 125 
<< pdiffusion >>
rect 157 124 158 125 
<< pdiffusion >>
rect 158 124 159 125 
<< pdiffusion >>
rect 159 124 160 125 
<< pdiffusion >>
rect 160 124 161 125 
<< pdiffusion >>
rect 161 124 162 125 
<< m1 >>
rect 163 124 164 125 
<< m1 >>
rect 165 124 166 125 
<< m2 >>
rect 166 124 167 125 
<< pdiffusion >>
rect 174 124 175 125 
<< pdiffusion >>
rect 175 124 176 125 
<< pdiffusion >>
rect 176 124 177 125 
<< pdiffusion >>
rect 177 124 178 125 
<< pdiffusion >>
rect 178 124 179 125 
<< pdiffusion >>
rect 179 124 180 125 
<< m1 >>
rect 181 124 182 125 
<< pdiffusion >>
rect 192 124 193 125 
<< pdiffusion >>
rect 193 124 194 125 
<< pdiffusion >>
rect 194 124 195 125 
<< pdiffusion >>
rect 195 124 196 125 
<< pdiffusion >>
rect 196 124 197 125 
<< pdiffusion >>
rect 197 124 198 125 
<< m1 >>
rect 199 124 200 125 
<< m1 >>
rect 208 124 209 125 
<< pdiffusion >>
rect 210 124 211 125 
<< pdiffusion >>
rect 211 124 212 125 
<< pdiffusion >>
rect 212 124 213 125 
<< pdiffusion >>
rect 213 124 214 125 
<< pdiffusion >>
rect 214 124 215 125 
<< pdiffusion >>
rect 215 124 216 125 
<< m1 >>
rect 217 124 218 125 
<< pdiffusion >>
rect 228 124 229 125 
<< pdiffusion >>
rect 229 124 230 125 
<< pdiffusion >>
rect 230 124 231 125 
<< pdiffusion >>
rect 231 124 232 125 
<< pdiffusion >>
rect 232 124 233 125 
<< pdiffusion >>
rect 233 124 234 125 
<< m1 >>
rect 235 124 236 125 
<< m1 >>
rect 244 124 245 125 
<< pdiffusion >>
rect 246 124 247 125 
<< pdiffusion >>
rect 247 124 248 125 
<< pdiffusion >>
rect 248 124 249 125 
<< pdiffusion >>
rect 249 124 250 125 
<< pdiffusion >>
rect 250 124 251 125 
<< pdiffusion >>
rect 251 124 252 125 
<< m1 >>
rect 253 124 254 125 
<< m1 >>
rect 255 124 256 125 
<< pdiffusion >>
rect 264 124 265 125 
<< pdiffusion >>
rect 265 124 266 125 
<< pdiffusion >>
rect 266 124 267 125 
<< pdiffusion >>
rect 267 124 268 125 
<< pdiffusion >>
rect 268 124 269 125 
<< pdiffusion >>
rect 269 124 270 125 
<< m1 >>
rect 271 124 272 125 
<< m2 >>
rect 272 124 273 125 
<< m1 >>
rect 278 124 279 125 
<< m1 >>
rect 280 124 281 125 
<< pdiffusion >>
rect 282 124 283 125 
<< pdiffusion >>
rect 283 124 284 125 
<< pdiffusion >>
rect 284 124 285 125 
<< pdiffusion >>
rect 285 124 286 125 
<< pdiffusion >>
rect 286 124 287 125 
<< pdiffusion >>
rect 287 124 288 125 
<< m1 >>
rect 298 124 299 125 
<< pdiffusion >>
rect 300 124 301 125 
<< pdiffusion >>
rect 301 124 302 125 
<< pdiffusion >>
rect 302 124 303 125 
<< pdiffusion >>
rect 303 124 304 125 
<< pdiffusion >>
rect 304 124 305 125 
<< pdiffusion >>
rect 305 124 306 125 
<< pdiffusion >>
rect 318 124 319 125 
<< pdiffusion >>
rect 319 124 320 125 
<< pdiffusion >>
rect 320 124 321 125 
<< pdiffusion >>
rect 321 124 322 125 
<< pdiffusion >>
rect 322 124 323 125 
<< pdiffusion >>
rect 323 124 324 125 
<< m1 >>
rect 334 124 335 125 
<< pdiffusion >>
rect 336 124 337 125 
<< pdiffusion >>
rect 337 124 338 125 
<< pdiffusion >>
rect 338 124 339 125 
<< pdiffusion >>
rect 339 124 340 125 
<< pdiffusion >>
rect 340 124 341 125 
<< pdiffusion >>
rect 341 124 342 125 
<< m1 >>
rect 343 124 344 125 
<< m1 >>
rect 345 124 346 125 
<< pdiffusion >>
rect 354 124 355 125 
<< pdiffusion >>
rect 355 124 356 125 
<< pdiffusion >>
rect 356 124 357 125 
<< pdiffusion >>
rect 357 124 358 125 
<< pdiffusion >>
rect 358 124 359 125 
<< pdiffusion >>
rect 359 124 360 125 
<< m1 >>
rect 361 124 362 125 
<< m2 >>
rect 361 124 362 125 
<< m1 >>
rect 366 124 367 125 
<< m1 >>
rect 370 124 371 125 
<< m2 >>
rect 370 124 371 125 
<< pdiffusion >>
rect 372 124 373 125 
<< pdiffusion >>
rect 373 124 374 125 
<< pdiffusion >>
rect 374 124 375 125 
<< pdiffusion >>
rect 375 124 376 125 
<< pdiffusion >>
rect 376 124 377 125 
<< pdiffusion >>
rect 377 124 378 125 
<< m1 >>
rect 379 124 380 125 
<< m2 >>
rect 379 124 380 125 
<< m1 >>
rect 381 124 382 125 
<< pdiffusion >>
rect 390 124 391 125 
<< pdiffusion >>
rect 391 124 392 125 
<< pdiffusion >>
rect 392 124 393 125 
<< pdiffusion >>
rect 393 124 394 125 
<< pdiffusion >>
rect 394 124 395 125 
<< pdiffusion >>
rect 395 124 396 125 
<< pdiffusion >>
rect 408 124 409 125 
<< pdiffusion >>
rect 409 124 410 125 
<< pdiffusion >>
rect 410 124 411 125 
<< pdiffusion >>
rect 411 124 412 125 
<< pdiffusion >>
rect 412 124 413 125 
<< pdiffusion >>
rect 413 124 414 125 
<< m1 >>
rect 430 124 431 125 
<< m2 >>
rect 431 124 432 125 
<< pdiffusion >>
rect 444 124 445 125 
<< pdiffusion >>
rect 445 124 446 125 
<< pdiffusion >>
rect 446 124 447 125 
<< pdiffusion >>
rect 447 124 448 125 
<< pdiffusion >>
rect 448 124 449 125 
<< pdiffusion >>
rect 449 124 450 125 
<< m1 >>
rect 456 124 457 125 
<< pdiffusion >>
rect 462 124 463 125 
<< pdiffusion >>
rect 463 124 464 125 
<< pdiffusion >>
rect 464 124 465 125 
<< pdiffusion >>
rect 465 124 466 125 
<< pdiffusion >>
rect 466 124 467 125 
<< pdiffusion >>
rect 467 124 468 125 
<< m1 >>
rect 478 124 479 125 
<< m1 >>
rect 484 124 485 125 
<< pdiffusion >>
rect 498 124 499 125 
<< pdiffusion >>
rect 499 124 500 125 
<< pdiffusion >>
rect 500 124 501 125 
<< pdiffusion >>
rect 501 124 502 125 
<< pdiffusion >>
rect 502 124 503 125 
<< pdiffusion >>
rect 503 124 504 125 
<< pdiffusion >>
rect 516 124 517 125 
<< pdiffusion >>
rect 517 124 518 125 
<< pdiffusion >>
rect 518 124 519 125 
<< pdiffusion >>
rect 519 124 520 125 
<< pdiffusion >>
rect 520 124 521 125 
<< pdiffusion >>
rect 521 124 522 125 
<< pdiffusion >>
rect 12 125 13 126 
<< pdiffusion >>
rect 13 125 14 126 
<< pdiffusion >>
rect 14 125 15 126 
<< pdiffusion >>
rect 15 125 16 126 
<< pdiffusion >>
rect 16 125 17 126 
<< pdiffusion >>
rect 17 125 18 126 
<< m1 >>
rect 19 125 20 126 
<< pdiffusion >>
rect 30 125 31 126 
<< pdiffusion >>
rect 31 125 32 126 
<< pdiffusion >>
rect 32 125 33 126 
<< pdiffusion >>
rect 33 125 34 126 
<< pdiffusion >>
rect 34 125 35 126 
<< pdiffusion >>
rect 35 125 36 126 
<< m1 >>
rect 46 125 47 126 
<< pdiffusion >>
rect 48 125 49 126 
<< pdiffusion >>
rect 49 125 50 126 
<< pdiffusion >>
rect 50 125 51 126 
<< pdiffusion >>
rect 51 125 52 126 
<< pdiffusion >>
rect 52 125 53 126 
<< pdiffusion >>
rect 53 125 54 126 
<< m1 >>
rect 64 125 65 126 
<< pdiffusion >>
rect 66 125 67 126 
<< pdiffusion >>
rect 67 125 68 126 
<< pdiffusion >>
rect 68 125 69 126 
<< pdiffusion >>
rect 69 125 70 126 
<< pdiffusion >>
rect 70 125 71 126 
<< pdiffusion >>
rect 71 125 72 126 
<< pdiffusion >>
rect 84 125 85 126 
<< m1 >>
rect 85 125 86 126 
<< pdiffusion >>
rect 85 125 86 126 
<< pdiffusion >>
rect 86 125 87 126 
<< m1 >>
rect 87 125 88 126 
<< m2 >>
rect 87 125 88 126 
<< m2c >>
rect 87 125 88 126 
<< m1 >>
rect 87 125 88 126 
<< m2 >>
rect 87 125 88 126 
<< pdiffusion >>
rect 87 125 88 126 
<< m1 >>
rect 88 125 89 126 
<< pdiffusion >>
rect 88 125 89 126 
<< pdiffusion >>
rect 89 125 90 126 
<< m1 >>
rect 92 125 93 126 
<< m2 >>
rect 99 125 100 126 
<< m1 >>
rect 100 125 101 126 
<< pdiffusion >>
rect 102 125 103 126 
<< pdiffusion >>
rect 103 125 104 126 
<< pdiffusion >>
rect 104 125 105 126 
<< pdiffusion >>
rect 105 125 106 126 
<< pdiffusion >>
rect 106 125 107 126 
<< pdiffusion >>
rect 107 125 108 126 
<< m1 >>
rect 109 125 110 126 
<< m1 >>
rect 118 125 119 126 
<< pdiffusion >>
rect 120 125 121 126 
<< pdiffusion >>
rect 121 125 122 126 
<< pdiffusion >>
rect 122 125 123 126 
<< pdiffusion >>
rect 123 125 124 126 
<< m1 >>
rect 124 125 125 126 
<< pdiffusion >>
rect 124 125 125 126 
<< pdiffusion >>
rect 125 125 126 126 
<< m1 >>
rect 129 125 130 126 
<< m1 >>
rect 131 125 132 126 
<< m1 >>
rect 133 125 134 126 
<< m1 >>
rect 136 125 137 126 
<< pdiffusion >>
rect 138 125 139 126 
<< pdiffusion >>
rect 139 125 140 126 
<< pdiffusion >>
rect 140 125 141 126 
<< pdiffusion >>
rect 141 125 142 126 
<< m1 >>
rect 142 125 143 126 
<< pdiffusion >>
rect 142 125 143 126 
<< pdiffusion >>
rect 143 125 144 126 
<< m1 >>
rect 145 125 146 126 
<< m2 >>
rect 145 125 146 126 
<< m2c >>
rect 145 125 146 126 
<< m1 >>
rect 145 125 146 126 
<< m2 >>
rect 145 125 146 126 
<< m1 >>
rect 154 125 155 126 
<< pdiffusion >>
rect 156 125 157 126 
<< pdiffusion >>
rect 157 125 158 126 
<< pdiffusion >>
rect 158 125 159 126 
<< pdiffusion >>
rect 159 125 160 126 
<< pdiffusion >>
rect 160 125 161 126 
<< pdiffusion >>
rect 161 125 162 126 
<< m1 >>
rect 163 125 164 126 
<< m1 >>
rect 165 125 166 126 
<< m2 >>
rect 166 125 167 126 
<< pdiffusion >>
rect 174 125 175 126 
<< m1 >>
rect 175 125 176 126 
<< pdiffusion >>
rect 175 125 176 126 
<< pdiffusion >>
rect 176 125 177 126 
<< pdiffusion >>
rect 177 125 178 126 
<< pdiffusion >>
rect 178 125 179 126 
<< pdiffusion >>
rect 179 125 180 126 
<< m1 >>
rect 181 125 182 126 
<< pdiffusion >>
rect 192 125 193 126 
<< pdiffusion >>
rect 193 125 194 126 
<< pdiffusion >>
rect 194 125 195 126 
<< pdiffusion >>
rect 195 125 196 126 
<< pdiffusion >>
rect 196 125 197 126 
<< pdiffusion >>
rect 197 125 198 126 
<< m1 >>
rect 199 125 200 126 
<< m1 >>
rect 208 125 209 126 
<< pdiffusion >>
rect 210 125 211 126 
<< m1 >>
rect 211 125 212 126 
<< pdiffusion >>
rect 211 125 212 126 
<< pdiffusion >>
rect 212 125 213 126 
<< pdiffusion >>
rect 213 125 214 126 
<< pdiffusion >>
rect 214 125 215 126 
<< pdiffusion >>
rect 215 125 216 126 
<< m1 >>
rect 217 125 218 126 
<< pdiffusion >>
rect 228 125 229 126 
<< pdiffusion >>
rect 229 125 230 126 
<< pdiffusion >>
rect 230 125 231 126 
<< pdiffusion >>
rect 231 125 232 126 
<< m1 >>
rect 232 125 233 126 
<< pdiffusion >>
rect 232 125 233 126 
<< pdiffusion >>
rect 233 125 234 126 
<< m1 >>
rect 235 125 236 126 
<< m1 >>
rect 244 125 245 126 
<< pdiffusion >>
rect 246 125 247 126 
<< pdiffusion >>
rect 247 125 248 126 
<< pdiffusion >>
rect 248 125 249 126 
<< pdiffusion >>
rect 249 125 250 126 
<< m1 >>
rect 250 125 251 126 
<< pdiffusion >>
rect 250 125 251 126 
<< pdiffusion >>
rect 251 125 252 126 
<< m1 >>
rect 253 125 254 126 
<< m1 >>
rect 255 125 256 126 
<< pdiffusion >>
rect 264 125 265 126 
<< pdiffusion >>
rect 265 125 266 126 
<< pdiffusion >>
rect 266 125 267 126 
<< pdiffusion >>
rect 267 125 268 126 
<< m1 >>
rect 268 125 269 126 
<< pdiffusion >>
rect 268 125 269 126 
<< pdiffusion >>
rect 269 125 270 126 
<< m1 >>
rect 271 125 272 126 
<< m2 >>
rect 272 125 273 126 
<< m1 >>
rect 278 125 279 126 
<< m1 >>
rect 280 125 281 126 
<< pdiffusion >>
rect 282 125 283 126 
<< pdiffusion >>
rect 283 125 284 126 
<< pdiffusion >>
rect 284 125 285 126 
<< pdiffusion >>
rect 285 125 286 126 
<< pdiffusion >>
rect 286 125 287 126 
<< pdiffusion >>
rect 287 125 288 126 
<< m1 >>
rect 298 125 299 126 
<< pdiffusion >>
rect 300 125 301 126 
<< pdiffusion >>
rect 301 125 302 126 
<< pdiffusion >>
rect 302 125 303 126 
<< pdiffusion >>
rect 303 125 304 126 
<< pdiffusion >>
rect 304 125 305 126 
<< pdiffusion >>
rect 305 125 306 126 
<< pdiffusion >>
rect 318 125 319 126 
<< pdiffusion >>
rect 319 125 320 126 
<< pdiffusion >>
rect 320 125 321 126 
<< pdiffusion >>
rect 321 125 322 126 
<< pdiffusion >>
rect 322 125 323 126 
<< pdiffusion >>
rect 323 125 324 126 
<< m1 >>
rect 334 125 335 126 
<< pdiffusion >>
rect 336 125 337 126 
<< pdiffusion >>
rect 337 125 338 126 
<< pdiffusion >>
rect 338 125 339 126 
<< pdiffusion >>
rect 339 125 340 126 
<< pdiffusion >>
rect 340 125 341 126 
<< pdiffusion >>
rect 341 125 342 126 
<< m1 >>
rect 343 125 344 126 
<< m1 >>
rect 345 125 346 126 
<< pdiffusion >>
rect 354 125 355 126 
<< pdiffusion >>
rect 355 125 356 126 
<< pdiffusion >>
rect 356 125 357 126 
<< pdiffusion >>
rect 357 125 358 126 
<< pdiffusion >>
rect 358 125 359 126 
<< pdiffusion >>
rect 359 125 360 126 
<< m1 >>
rect 361 125 362 126 
<< m2 >>
rect 361 125 362 126 
<< m1 >>
rect 366 125 367 126 
<< m1 >>
rect 370 125 371 126 
<< m2 >>
rect 370 125 371 126 
<< pdiffusion >>
rect 372 125 373 126 
<< m1 >>
rect 373 125 374 126 
<< pdiffusion >>
rect 373 125 374 126 
<< pdiffusion >>
rect 374 125 375 126 
<< pdiffusion >>
rect 375 125 376 126 
<< pdiffusion >>
rect 376 125 377 126 
<< pdiffusion >>
rect 377 125 378 126 
<< m1 >>
rect 379 125 380 126 
<< m2 >>
rect 379 125 380 126 
<< m1 >>
rect 381 125 382 126 
<< pdiffusion >>
rect 390 125 391 126 
<< pdiffusion >>
rect 391 125 392 126 
<< pdiffusion >>
rect 392 125 393 126 
<< pdiffusion >>
rect 393 125 394 126 
<< m1 >>
rect 394 125 395 126 
<< pdiffusion >>
rect 394 125 395 126 
<< pdiffusion >>
rect 395 125 396 126 
<< pdiffusion >>
rect 408 125 409 126 
<< m1 >>
rect 409 125 410 126 
<< pdiffusion >>
rect 409 125 410 126 
<< pdiffusion >>
rect 410 125 411 126 
<< pdiffusion >>
rect 411 125 412 126 
<< m1 >>
rect 412 125 413 126 
<< pdiffusion >>
rect 412 125 413 126 
<< pdiffusion >>
rect 413 125 414 126 
<< m1 >>
rect 430 125 431 126 
<< m2 >>
rect 431 125 432 126 
<< pdiffusion >>
rect 444 125 445 126 
<< pdiffusion >>
rect 445 125 446 126 
<< pdiffusion >>
rect 446 125 447 126 
<< pdiffusion >>
rect 447 125 448 126 
<< pdiffusion >>
rect 448 125 449 126 
<< pdiffusion >>
rect 449 125 450 126 
<< m1 >>
rect 456 125 457 126 
<< pdiffusion >>
rect 462 125 463 126 
<< pdiffusion >>
rect 463 125 464 126 
<< pdiffusion >>
rect 464 125 465 126 
<< pdiffusion >>
rect 465 125 466 126 
<< m1 >>
rect 466 125 467 126 
<< pdiffusion >>
rect 466 125 467 126 
<< pdiffusion >>
rect 467 125 468 126 
<< m1 >>
rect 478 125 479 126 
<< m1 >>
rect 484 125 485 126 
<< pdiffusion >>
rect 498 125 499 126 
<< pdiffusion >>
rect 499 125 500 126 
<< pdiffusion >>
rect 500 125 501 126 
<< pdiffusion >>
rect 501 125 502 126 
<< m1 >>
rect 502 125 503 126 
<< pdiffusion >>
rect 502 125 503 126 
<< pdiffusion >>
rect 503 125 504 126 
<< pdiffusion >>
rect 516 125 517 126 
<< pdiffusion >>
rect 517 125 518 126 
<< pdiffusion >>
rect 518 125 519 126 
<< pdiffusion >>
rect 519 125 520 126 
<< pdiffusion >>
rect 520 125 521 126 
<< pdiffusion >>
rect 521 125 522 126 
<< m1 >>
rect 19 126 20 127 
<< m1 >>
rect 46 126 47 127 
<< m1 >>
rect 64 126 65 127 
<< m1 >>
rect 85 126 86 127 
<< m1 >>
rect 88 126 89 127 
<< m2 >>
rect 88 126 89 127 
<< m1 >>
rect 92 126 93 127 
<< m2 >>
rect 99 126 100 127 
<< m1 >>
rect 100 126 101 127 
<< m1 >>
rect 109 126 110 127 
<< m1 >>
rect 118 126 119 127 
<< m1 >>
rect 124 126 125 127 
<< m1 >>
rect 129 126 130 127 
<< m1 >>
rect 131 126 132 127 
<< m1 >>
rect 133 126 134 127 
<< m1 >>
rect 136 126 137 127 
<< m1 >>
rect 142 126 143 127 
<< m2 >>
rect 145 126 146 127 
<< m1 >>
rect 154 126 155 127 
<< m1 >>
rect 163 126 164 127 
<< m1 >>
rect 165 126 166 127 
<< m2 >>
rect 166 126 167 127 
<< m1 >>
rect 175 126 176 127 
<< m1 >>
rect 181 126 182 127 
<< m1 >>
rect 199 126 200 127 
<< m1 >>
rect 208 126 209 127 
<< m1 >>
rect 211 126 212 127 
<< m1 >>
rect 217 126 218 127 
<< m1 >>
rect 232 126 233 127 
<< m1 >>
rect 235 126 236 127 
<< m1 >>
rect 244 126 245 127 
<< m1 >>
rect 250 126 251 127 
<< m1 >>
rect 253 126 254 127 
<< m1 >>
rect 255 126 256 127 
<< m1 >>
rect 268 126 269 127 
<< m1 >>
rect 271 126 272 127 
<< m2 >>
rect 272 126 273 127 
<< m1 >>
rect 278 126 279 127 
<< m1 >>
rect 280 126 281 127 
<< m1 >>
rect 298 126 299 127 
<< m1 >>
rect 334 126 335 127 
<< m1 >>
rect 343 126 344 127 
<< m1 >>
rect 345 126 346 127 
<< m1 >>
rect 361 126 362 127 
<< m2 >>
rect 361 126 362 127 
<< m1 >>
rect 366 126 367 127 
<< m1 >>
rect 370 126 371 127 
<< m2 >>
rect 370 126 371 127 
<< m1 >>
rect 373 126 374 127 
<< m1 >>
rect 379 126 380 127 
<< m2 >>
rect 379 126 380 127 
<< m1 >>
rect 381 126 382 127 
<< m1 >>
rect 394 126 395 127 
<< m1 >>
rect 409 126 410 127 
<< m1 >>
rect 412 126 413 127 
<< m1 >>
rect 430 126 431 127 
<< m2 >>
rect 431 126 432 127 
<< m1 >>
rect 456 126 457 127 
<< m1 >>
rect 466 126 467 127 
<< m1 >>
rect 478 126 479 127 
<< m1 >>
rect 484 126 485 127 
<< m1 >>
rect 502 126 503 127 
<< m1 >>
rect 19 127 20 128 
<< m1 >>
rect 46 127 47 128 
<< m1 >>
rect 64 127 65 128 
<< m1 >>
rect 85 127 86 128 
<< m2 >>
rect 88 127 89 128 
<< m1 >>
rect 92 127 93 128 
<< m2 >>
rect 99 127 100 128 
<< m1 >>
rect 100 127 101 128 
<< m2 >>
rect 100 127 101 128 
<< m2 >>
rect 101 127 102 128 
<< m1 >>
rect 102 127 103 128 
<< m2 >>
rect 102 127 103 128 
<< m2c >>
rect 102 127 103 128 
<< m1 >>
rect 102 127 103 128 
<< m2 >>
rect 102 127 103 128 
<< m1 >>
rect 109 127 110 128 
<< m1 >>
rect 118 127 119 128 
<< m1 >>
rect 124 127 125 128 
<< m1 >>
rect 129 127 130 128 
<< m1 >>
rect 131 127 132 128 
<< m1 >>
rect 133 127 134 128 
<< m1 >>
rect 136 127 137 128 
<< m1 >>
rect 142 127 143 128 
<< m1 >>
rect 143 127 144 128 
<< m1 >>
rect 144 127 145 128 
<< m1 >>
rect 145 127 146 128 
<< m2 >>
rect 145 127 146 128 
<< m1 >>
rect 146 127 147 128 
<< m1 >>
rect 147 127 148 128 
<< m1 >>
rect 148 127 149 128 
<< m1 >>
rect 149 127 150 128 
<< m1 >>
rect 150 127 151 128 
<< m1 >>
rect 151 127 152 128 
<< m1 >>
rect 152 127 153 128 
<< m1 >>
rect 153 127 154 128 
<< m1 >>
rect 154 127 155 128 
<< m1 >>
rect 161 127 162 128 
<< m2 >>
rect 161 127 162 128 
<< m2c >>
rect 161 127 162 128 
<< m1 >>
rect 161 127 162 128 
<< m2 >>
rect 161 127 162 128 
<< m2 >>
rect 162 127 163 128 
<< m1 >>
rect 163 127 164 128 
<< m2 >>
rect 163 127 164 128 
<< m2 >>
rect 164 127 165 128 
<< m1 >>
rect 165 127 166 128 
<< m2 >>
rect 165 127 166 128 
<< m2 >>
rect 166 127 167 128 
<< m1 >>
rect 175 127 176 128 
<< m1 >>
rect 181 127 182 128 
<< m1 >>
rect 199 127 200 128 
<< m1 >>
rect 208 127 209 128 
<< m1 >>
rect 209 127 210 128 
<< m1 >>
rect 210 127 211 128 
<< m1 >>
rect 211 127 212 128 
<< m1 >>
rect 217 127 218 128 
<< m1 >>
rect 232 127 233 128 
<< m1 >>
rect 235 127 236 128 
<< m1 >>
rect 244 127 245 128 
<< m1 >>
rect 250 127 251 128 
<< m1 >>
rect 251 127 252 128 
<< m2 >>
rect 251 127 252 128 
<< m2c >>
rect 251 127 252 128 
<< m1 >>
rect 251 127 252 128 
<< m2 >>
rect 251 127 252 128 
<< m2 >>
rect 252 127 253 128 
<< m1 >>
rect 253 127 254 128 
<< m2 >>
rect 253 127 254 128 
<< m2 >>
rect 254 127 255 128 
<< m1 >>
rect 255 127 256 128 
<< m2 >>
rect 255 127 256 128 
<< m2c >>
rect 255 127 256 128 
<< m1 >>
rect 255 127 256 128 
<< m2 >>
rect 255 127 256 128 
<< m1 >>
rect 268 127 269 128 
<< m1 >>
rect 269 127 270 128 
<< m2 >>
rect 269 127 270 128 
<< m2c >>
rect 269 127 270 128 
<< m1 >>
rect 269 127 270 128 
<< m2 >>
rect 269 127 270 128 
<< m2 >>
rect 270 127 271 128 
<< m1 >>
rect 271 127 272 128 
<< m2 >>
rect 271 127 272 128 
<< m2 >>
rect 272 127 273 128 
<< m1 >>
rect 278 127 279 128 
<< m1 >>
rect 280 127 281 128 
<< m1 >>
rect 298 127 299 128 
<< m1 >>
rect 334 127 335 128 
<< m1 >>
rect 343 127 344 128 
<< m1 >>
rect 345 127 346 128 
<< m1 >>
rect 361 127 362 128 
<< m2 >>
rect 361 127 362 128 
<< m1 >>
rect 366 127 367 128 
<< m1 >>
rect 370 127 371 128 
<< m2 >>
rect 370 127 371 128 
<< m1 >>
rect 371 127 372 128 
<< m1 >>
rect 372 127 373 128 
<< m1 >>
rect 373 127 374 128 
<< m1 >>
rect 379 127 380 128 
<< m2 >>
rect 379 127 380 128 
<< m1 >>
rect 381 127 382 128 
<< m1 >>
rect 394 127 395 128 
<< m1 >>
rect 395 127 396 128 
<< m1 >>
rect 396 127 397 128 
<< m1 >>
rect 397 127 398 128 
<< m1 >>
rect 398 127 399 128 
<< m1 >>
rect 399 127 400 128 
<< m1 >>
rect 400 127 401 128 
<< m1 >>
rect 401 127 402 128 
<< m1 >>
rect 402 127 403 128 
<< m1 >>
rect 403 127 404 128 
<< m1 >>
rect 404 127 405 128 
<< m1 >>
rect 405 127 406 128 
<< m1 >>
rect 406 127 407 128 
<< m1 >>
rect 407 127 408 128 
<< m1 >>
rect 408 127 409 128 
<< m1 >>
rect 409 127 410 128 
<< m1 >>
rect 412 127 413 128 
<< m2 >>
rect 420 127 421 128 
<< m2 >>
rect 421 127 422 128 
<< m2 >>
rect 422 127 423 128 
<< m2 >>
rect 423 127 424 128 
<< m2 >>
rect 424 127 425 128 
<< m2 >>
rect 425 127 426 128 
<< m2 >>
rect 426 127 427 128 
<< m2 >>
rect 427 127 428 128 
<< m2 >>
rect 428 127 429 128 
<< m2 >>
rect 429 127 430 128 
<< m1 >>
rect 430 127 431 128 
<< m2 >>
rect 430 127 431 128 
<< m2 >>
rect 431 127 432 128 
<< m1 >>
rect 456 127 457 128 
<< m1 >>
rect 466 127 467 128 
<< m1 >>
rect 467 127 468 128 
<< m1 >>
rect 468 127 469 128 
<< m1 >>
rect 469 127 470 128 
<< m1 >>
rect 478 127 479 128 
<< m1 >>
rect 484 127 485 128 
<< m1 >>
rect 502 127 503 128 
<< m1 >>
rect 19 128 20 129 
<< m1 >>
rect 46 128 47 129 
<< m1 >>
rect 64 128 65 129 
<< m1 >>
rect 85 128 86 129 
<< m1 >>
rect 86 128 87 129 
<< m1 >>
rect 87 128 88 129 
<< m1 >>
rect 88 128 89 129 
<< m2 >>
rect 88 128 89 129 
<< m1 >>
rect 89 128 90 129 
<< m1 >>
rect 90 128 91 129 
<< m2 >>
rect 90 128 91 129 
<< m2c >>
rect 90 128 91 129 
<< m1 >>
rect 90 128 91 129 
<< m2 >>
rect 90 128 91 129 
<< m2 >>
rect 91 128 92 129 
<< m1 >>
rect 92 128 93 129 
<< m2 >>
rect 92 128 93 129 
<< m2 >>
rect 93 128 94 129 
<< m1 >>
rect 94 128 95 129 
<< m2 >>
rect 94 128 95 129 
<< m2c >>
rect 94 128 95 129 
<< m1 >>
rect 94 128 95 129 
<< m2 >>
rect 94 128 95 129 
<< m1 >>
rect 100 128 101 129 
<< m1 >>
rect 102 128 103 129 
<< m1 >>
rect 104 128 105 129 
<< m2 >>
rect 104 128 105 129 
<< m2c >>
rect 104 128 105 129 
<< m1 >>
rect 104 128 105 129 
<< m2 >>
rect 104 128 105 129 
<< m1 >>
rect 105 128 106 129 
<< m1 >>
rect 106 128 107 129 
<< m1 >>
rect 107 128 108 129 
<< m1 >>
rect 108 128 109 129 
<< m1 >>
rect 109 128 110 129 
<< m1 >>
rect 118 128 119 129 
<< m1 >>
rect 124 128 125 129 
<< m1 >>
rect 129 128 130 129 
<< m1 >>
rect 131 128 132 129 
<< m1 >>
rect 133 128 134 129 
<< m1 >>
rect 136 128 137 129 
<< m2 >>
rect 145 128 146 129 
<< m1 >>
rect 161 128 162 129 
<< m1 >>
rect 163 128 164 129 
<< m1 >>
rect 165 128 166 129 
<< m1 >>
rect 175 128 176 129 
<< m1 >>
rect 176 128 177 129 
<< m1 >>
rect 177 128 178 129 
<< m1 >>
rect 178 128 179 129 
<< m1 >>
rect 179 128 180 129 
<< m1 >>
rect 180 128 181 129 
<< m1 >>
rect 181 128 182 129 
<< m1 >>
rect 199 128 200 129 
<< m1 >>
rect 217 128 218 129 
<< m1 >>
rect 232 128 233 129 
<< m1 >>
rect 235 128 236 129 
<< m1 >>
rect 244 128 245 129 
<< m1 >>
rect 253 128 254 129 
<< m1 >>
rect 271 128 272 129 
<< m1 >>
rect 278 128 279 129 
<< m2 >>
rect 278 128 279 129 
<< m2c >>
rect 278 128 279 129 
<< m1 >>
rect 278 128 279 129 
<< m2 >>
rect 278 128 279 129 
<< m1 >>
rect 280 128 281 129 
<< m2 >>
rect 280 128 281 129 
<< m2c >>
rect 280 128 281 129 
<< m1 >>
rect 280 128 281 129 
<< m2 >>
rect 280 128 281 129 
<< m1 >>
rect 298 128 299 129 
<< m1 >>
rect 334 128 335 129 
<< m1 >>
rect 343 128 344 129 
<< m1 >>
rect 345 128 346 129 
<< m1 >>
rect 358 128 359 129 
<< m1 >>
rect 359 128 360 129 
<< m2 >>
rect 359 128 360 129 
<< m2c >>
rect 359 128 360 129 
<< m1 >>
rect 359 128 360 129 
<< m2 >>
rect 359 128 360 129 
<< m2 >>
rect 360 128 361 129 
<< m1 >>
rect 361 128 362 129 
<< m2 >>
rect 361 128 362 129 
<< m1 >>
rect 366 128 367 129 
<< m2 >>
rect 370 128 371 129 
<< m1 >>
rect 379 128 380 129 
<< m2 >>
rect 379 128 380 129 
<< m1 >>
rect 381 128 382 129 
<< m2 >>
rect 381 128 382 129 
<< m2c >>
rect 381 128 382 129 
<< m1 >>
rect 381 128 382 129 
<< m2 >>
rect 381 128 382 129 
<< m1 >>
rect 412 128 413 129 
<< m1 >>
rect 413 128 414 129 
<< m1 >>
rect 414 128 415 129 
<< m1 >>
rect 415 128 416 129 
<< m1 >>
rect 416 128 417 129 
<< m1 >>
rect 417 128 418 129 
<< m1 >>
rect 418 128 419 129 
<< m1 >>
rect 419 128 420 129 
<< m1 >>
rect 420 128 421 129 
<< m2 >>
rect 420 128 421 129 
<< m1 >>
rect 421 128 422 129 
<< m1 >>
rect 422 128 423 129 
<< m1 >>
rect 423 128 424 129 
<< m1 >>
rect 424 128 425 129 
<< m1 >>
rect 425 128 426 129 
<< m1 >>
rect 426 128 427 129 
<< m1 >>
rect 427 128 428 129 
<< m1 >>
rect 430 128 431 129 
<< m1 >>
rect 456 128 457 129 
<< m1 >>
rect 469 128 470 129 
<< m1 >>
rect 478 128 479 129 
<< m1 >>
rect 484 128 485 129 
<< m1 >>
rect 502 128 503 129 
<< m1 >>
rect 19 129 20 130 
<< m1 >>
rect 46 129 47 130 
<< m1 >>
rect 64 129 65 130 
<< m2 >>
rect 88 129 89 130 
<< m1 >>
rect 92 129 93 130 
<< m1 >>
rect 94 129 95 130 
<< m1 >>
rect 95 129 96 130 
<< m1 >>
rect 96 129 97 130 
<< m1 >>
rect 97 129 98 130 
<< m1 >>
rect 98 129 99 130 
<< m2 >>
rect 98 129 99 130 
<< m2c >>
rect 98 129 99 130 
<< m1 >>
rect 98 129 99 130 
<< m2 >>
rect 98 129 99 130 
<< m2 >>
rect 99 129 100 130 
<< m1 >>
rect 100 129 101 130 
<< m1 >>
rect 102 129 103 130 
<< m2 >>
rect 104 129 105 130 
<< m1 >>
rect 118 129 119 130 
<< m1 >>
rect 124 129 125 130 
<< m1 >>
rect 129 129 130 130 
<< m1 >>
rect 131 129 132 130 
<< m1 >>
rect 133 129 134 130 
<< m1 >>
rect 136 129 137 130 
<< m1 >>
rect 145 129 146 130 
<< m2 >>
rect 145 129 146 130 
<< m2c >>
rect 145 129 146 130 
<< m1 >>
rect 145 129 146 130 
<< m2 >>
rect 145 129 146 130 
<< m1 >>
rect 161 129 162 130 
<< m1 >>
rect 163 129 164 130 
<< m1 >>
rect 165 129 166 130 
<< m1 >>
rect 199 129 200 130 
<< m1 >>
rect 217 129 218 130 
<< m1 >>
rect 232 129 233 130 
<< m1 >>
rect 235 129 236 130 
<< m1 >>
rect 244 129 245 130 
<< m1 >>
rect 253 129 254 130 
<< m1 >>
rect 271 129 272 130 
<< m2 >>
rect 278 129 279 130 
<< m2 >>
rect 280 129 281 130 
<< m2 >>
rect 284 129 285 130 
<< m1 >>
rect 285 129 286 130 
<< m2 >>
rect 285 129 286 130 
<< m2c >>
rect 285 129 286 130 
<< m1 >>
rect 285 129 286 130 
<< m2 >>
rect 285 129 286 130 
<< m1 >>
rect 286 129 287 130 
<< m1 >>
rect 287 129 288 130 
<< m1 >>
rect 288 129 289 130 
<< m1 >>
rect 289 129 290 130 
<< m1 >>
rect 290 129 291 130 
<< m1 >>
rect 291 129 292 130 
<< m1 >>
rect 292 129 293 130 
<< m1 >>
rect 293 129 294 130 
<< m1 >>
rect 294 129 295 130 
<< m1 >>
rect 295 129 296 130 
<< m1 >>
rect 296 129 297 130 
<< m1 >>
rect 297 129 298 130 
<< m1 >>
rect 298 129 299 130 
<< m1 >>
rect 334 129 335 130 
<< m1 >>
rect 343 129 344 130 
<< m1 >>
rect 345 129 346 130 
<< m1 >>
rect 358 129 359 130 
<< m1 >>
rect 361 129 362 130 
<< m1 >>
rect 366 129 367 130 
<< m1 >>
rect 370 129 371 130 
<< m2 >>
rect 370 129 371 130 
<< m2c >>
rect 370 129 371 130 
<< m1 >>
rect 370 129 371 130 
<< m2 >>
rect 370 129 371 130 
<< m1 >>
rect 379 129 380 130 
<< m2 >>
rect 379 129 380 130 
<< m2 >>
rect 381 129 382 130 
<< m2 >>
rect 420 129 421 130 
<< m1 >>
rect 427 129 428 130 
<< m1 >>
rect 430 129 431 130 
<< m1 >>
rect 456 129 457 130 
<< m1 >>
rect 469 129 470 130 
<< m1 >>
rect 478 129 479 130 
<< m1 >>
rect 484 129 485 130 
<< m1 >>
rect 502 129 503 130 
<< m1 >>
rect 19 130 20 131 
<< m1 >>
rect 46 130 47 131 
<< m1 >>
rect 64 130 65 131 
<< m1 >>
rect 88 130 89 131 
<< m2 >>
rect 88 130 89 131 
<< m2c >>
rect 88 130 89 131 
<< m1 >>
rect 88 130 89 131 
<< m2 >>
rect 88 130 89 131 
<< m1 >>
rect 92 130 93 131 
<< m2 >>
rect 99 130 100 131 
<< m1 >>
rect 100 130 101 131 
<< m2 >>
rect 100 130 101 131 
<< m2 >>
rect 101 130 102 131 
<< m1 >>
rect 102 130 103 131 
<< m2 >>
rect 102 130 103 131 
<< m1 >>
rect 103 130 104 131 
<< m2 >>
rect 103 130 104 131 
<< m1 >>
rect 104 130 105 131 
<< m2 >>
rect 104 130 105 131 
<< m1 >>
rect 105 130 106 131 
<< m1 >>
rect 106 130 107 131 
<< m1 >>
rect 107 130 108 131 
<< m1 >>
rect 108 130 109 131 
<< m1 >>
rect 109 130 110 131 
<< m1 >>
rect 118 130 119 131 
<< m1 >>
rect 124 130 125 131 
<< m1 >>
rect 129 130 130 131 
<< m1 >>
rect 131 130 132 131 
<< m1 >>
rect 133 130 134 131 
<< m1 >>
rect 136 130 137 131 
<< m1 >>
rect 145 130 146 131 
<< m1 >>
rect 161 130 162 131 
<< m1 >>
rect 163 130 164 131 
<< m1 >>
rect 165 130 166 131 
<< m1 >>
rect 166 130 167 131 
<< m1 >>
rect 167 130 168 131 
<< m1 >>
rect 168 130 169 131 
<< m1 >>
rect 169 130 170 131 
<< m1 >>
rect 170 130 171 131 
<< m1 >>
rect 171 130 172 131 
<< m1 >>
rect 172 130 173 131 
<< m1 >>
rect 173 130 174 131 
<< m1 >>
rect 174 130 175 131 
<< m1 >>
rect 175 130 176 131 
<< m1 >>
rect 176 130 177 131 
<< m1 >>
rect 177 130 178 131 
<< m1 >>
rect 178 130 179 131 
<< m1 >>
rect 179 130 180 131 
<< m1 >>
rect 180 130 181 131 
<< m1 >>
rect 181 130 182 131 
<< m1 >>
rect 182 130 183 131 
<< m1 >>
rect 183 130 184 131 
<< m1 >>
rect 184 130 185 131 
<< m1 >>
rect 185 130 186 131 
<< m1 >>
rect 186 130 187 131 
<< m1 >>
rect 187 130 188 131 
<< m1 >>
rect 188 130 189 131 
<< m1 >>
rect 189 130 190 131 
<< m1 >>
rect 190 130 191 131 
<< m1 >>
rect 191 130 192 131 
<< m1 >>
rect 192 130 193 131 
<< m1 >>
rect 193 130 194 131 
<< m1 >>
rect 194 130 195 131 
<< m1 >>
rect 195 130 196 131 
<< m1 >>
rect 196 130 197 131 
<< m1 >>
rect 197 130 198 131 
<< m2 >>
rect 197 130 198 131 
<< m2c >>
rect 197 130 198 131 
<< m1 >>
rect 197 130 198 131 
<< m2 >>
rect 197 130 198 131 
<< m2 >>
rect 198 130 199 131 
<< m1 >>
rect 199 130 200 131 
<< m2 >>
rect 199 130 200 131 
<< m2 >>
rect 200 130 201 131 
<< m1 >>
rect 201 130 202 131 
<< m2 >>
rect 201 130 202 131 
<< m2c >>
rect 201 130 202 131 
<< m1 >>
rect 201 130 202 131 
<< m2 >>
rect 201 130 202 131 
<< m1 >>
rect 202 130 203 131 
<< m1 >>
rect 203 130 204 131 
<< m1 >>
rect 204 130 205 131 
<< m1 >>
rect 205 130 206 131 
<< m1 >>
rect 206 130 207 131 
<< m1 >>
rect 207 130 208 131 
<< m1 >>
rect 208 130 209 131 
<< m1 >>
rect 209 130 210 131 
<< m1 >>
rect 210 130 211 131 
<< m1 >>
rect 211 130 212 131 
<< m1 >>
rect 212 130 213 131 
<< m1 >>
rect 213 130 214 131 
<< m1 >>
rect 214 130 215 131 
<< m1 >>
rect 215 130 216 131 
<< m2 >>
rect 215 130 216 131 
<< m2c >>
rect 215 130 216 131 
<< m1 >>
rect 215 130 216 131 
<< m2 >>
rect 215 130 216 131 
<< m2 >>
rect 216 130 217 131 
<< m1 >>
rect 217 130 218 131 
<< m2 >>
rect 217 130 218 131 
<< m1 >>
rect 226 130 227 131 
<< m1 >>
rect 227 130 228 131 
<< m1 >>
rect 228 130 229 131 
<< m1 >>
rect 229 130 230 131 
<< m1 >>
rect 230 130 231 131 
<< m1 >>
rect 231 130 232 131 
<< m1 >>
rect 232 130 233 131 
<< m1 >>
rect 235 130 236 131 
<< m1 >>
rect 244 130 245 131 
<< m1 >>
rect 253 130 254 131 
<< m1 >>
rect 254 130 255 131 
<< m1 >>
rect 255 130 256 131 
<< m1 >>
rect 256 130 257 131 
<< m1 >>
rect 257 130 258 131 
<< m1 >>
rect 258 130 259 131 
<< m1 >>
rect 259 130 260 131 
<< m1 >>
rect 260 130 261 131 
<< m1 >>
rect 261 130 262 131 
<< m1 >>
rect 262 130 263 131 
<< m1 >>
rect 263 130 264 131 
<< m1 >>
rect 264 130 265 131 
<< m1 >>
rect 265 130 266 131 
<< m1 >>
rect 271 130 272 131 
<< m1 >>
rect 272 130 273 131 
<< m1 >>
rect 273 130 274 131 
<< m1 >>
rect 274 130 275 131 
<< m1 >>
rect 275 130 276 131 
<< m1 >>
rect 276 130 277 131 
<< m1 >>
rect 277 130 278 131 
<< m1 >>
rect 278 130 279 131 
<< m2 >>
rect 278 130 279 131 
<< m1 >>
rect 279 130 280 131 
<< m1 >>
rect 280 130 281 131 
<< m2 >>
rect 280 130 281 131 
<< m1 >>
rect 281 130 282 131 
<< m1 >>
rect 282 130 283 131 
<< m2 >>
rect 282 130 283 131 
<< m1 >>
rect 283 130 284 131 
<< m2 >>
rect 283 130 284 131 
<< m2 >>
rect 284 130 285 131 
<< m1 >>
rect 334 130 335 131 
<< m1 >>
rect 343 130 344 131 
<< m1 >>
rect 345 130 346 131 
<< m1 >>
rect 358 130 359 131 
<< m2 >>
rect 358 130 359 131 
<< m2c >>
rect 358 130 359 131 
<< m1 >>
rect 358 130 359 131 
<< m2 >>
rect 358 130 359 131 
<< m1 >>
rect 361 130 362 131 
<< m2 >>
rect 361 130 362 131 
<< m2c >>
rect 361 130 362 131 
<< m1 >>
rect 361 130 362 131 
<< m2 >>
rect 361 130 362 131 
<< m1 >>
rect 366 130 367 131 
<< m2 >>
rect 366 130 367 131 
<< m2c >>
rect 366 130 367 131 
<< m1 >>
rect 366 130 367 131 
<< m2 >>
rect 366 130 367 131 
<< m1 >>
rect 370 130 371 131 
<< m2 >>
rect 370 130 371 131 
<< m1 >>
rect 379 130 380 131 
<< m2 >>
rect 379 130 380 131 
<< m1 >>
rect 380 130 381 131 
<< m1 >>
rect 381 130 382 131 
<< m2 >>
rect 381 130 382 131 
<< m1 >>
rect 382 130 383 131 
<< m2 >>
rect 382 130 383 131 
<< m1 >>
rect 383 130 384 131 
<< m2 >>
rect 383 130 384 131 
<< m1 >>
rect 384 130 385 131 
<< m2 >>
rect 384 130 385 131 
<< m1 >>
rect 385 130 386 131 
<< m2 >>
rect 385 130 386 131 
<< m1 >>
rect 386 130 387 131 
<< m2 >>
rect 386 130 387 131 
<< m1 >>
rect 387 130 388 131 
<< m2 >>
rect 387 130 388 131 
<< m1 >>
rect 388 130 389 131 
<< m2 >>
rect 388 130 389 131 
<< m1 >>
rect 389 130 390 131 
<< m2 >>
rect 389 130 390 131 
<< m1 >>
rect 390 130 391 131 
<< m2 >>
rect 390 130 391 131 
<< m1 >>
rect 391 130 392 131 
<< m2 >>
rect 391 130 392 131 
<< m1 >>
rect 392 130 393 131 
<< m2 >>
rect 392 130 393 131 
<< m1 >>
rect 393 130 394 131 
<< m2 >>
rect 393 130 394 131 
<< m1 >>
rect 394 130 395 131 
<< m2 >>
rect 394 130 395 131 
<< m1 >>
rect 395 130 396 131 
<< m2 >>
rect 395 130 396 131 
<< m1 >>
rect 396 130 397 131 
<< m2 >>
rect 396 130 397 131 
<< m1 >>
rect 397 130 398 131 
<< m2 >>
rect 397 130 398 131 
<< m1 >>
rect 398 130 399 131 
<< m2 >>
rect 398 130 399 131 
<< m1 >>
rect 399 130 400 131 
<< m2 >>
rect 399 130 400 131 
<< m1 >>
rect 400 130 401 131 
<< m2 >>
rect 400 130 401 131 
<< m1 >>
rect 401 130 402 131 
<< m2 >>
rect 401 130 402 131 
<< m1 >>
rect 402 130 403 131 
<< m2 >>
rect 402 130 403 131 
<< m1 >>
rect 403 130 404 131 
<< m2 >>
rect 403 130 404 131 
<< m1 >>
rect 404 130 405 131 
<< m2 >>
rect 404 130 405 131 
<< m1 >>
rect 405 130 406 131 
<< m2 >>
rect 405 130 406 131 
<< m1 >>
rect 406 130 407 131 
<< m2 >>
rect 406 130 407 131 
<< m1 >>
rect 407 130 408 131 
<< m2 >>
rect 407 130 408 131 
<< m1 >>
rect 408 130 409 131 
<< m2 >>
rect 408 130 409 131 
<< m1 >>
rect 409 130 410 131 
<< m2 >>
rect 409 130 410 131 
<< m1 >>
rect 410 130 411 131 
<< m2 >>
rect 410 130 411 131 
<< m1 >>
rect 411 130 412 131 
<< m2 >>
rect 411 130 412 131 
<< m1 >>
rect 412 130 413 131 
<< m2 >>
rect 412 130 413 131 
<< m1 >>
rect 413 130 414 131 
<< m2 >>
rect 413 130 414 131 
<< m1 >>
rect 414 130 415 131 
<< m2 >>
rect 414 130 415 131 
<< m1 >>
rect 415 130 416 131 
<< m2 >>
rect 415 130 416 131 
<< m2 >>
rect 416 130 417 131 
<< m1 >>
rect 417 130 418 131 
<< m2 >>
rect 417 130 418 131 
<< m2c >>
rect 417 130 418 131 
<< m1 >>
rect 417 130 418 131 
<< m2 >>
rect 417 130 418 131 
<< m1 >>
rect 418 130 419 131 
<< m1 >>
rect 419 130 420 131 
<< m2 >>
rect 420 130 421 131 
<< m1 >>
rect 427 130 428 131 
<< m1 >>
rect 430 130 431 131 
<< m1 >>
rect 456 130 457 131 
<< m1 >>
rect 469 130 470 131 
<< m1 >>
rect 478 130 479 131 
<< m1 >>
rect 484 130 485 131 
<< m1 >>
rect 485 130 486 131 
<< m1 >>
rect 486 130 487 131 
<< m1 >>
rect 487 130 488 131 
<< m1 >>
rect 488 130 489 131 
<< m1 >>
rect 489 130 490 131 
<< m1 >>
rect 490 130 491 131 
<< m1 >>
rect 491 130 492 131 
<< m1 >>
rect 492 130 493 131 
<< m1 >>
rect 493 130 494 131 
<< m1 >>
rect 494 130 495 131 
<< m1 >>
rect 495 130 496 131 
<< m1 >>
rect 496 130 497 131 
<< m1 >>
rect 497 130 498 131 
<< m1 >>
rect 498 130 499 131 
<< m1 >>
rect 499 130 500 131 
<< m1 >>
rect 500 130 501 131 
<< m1 >>
rect 501 130 502 131 
<< m1 >>
rect 502 130 503 131 
<< m1 >>
rect 19 131 20 132 
<< m1 >>
rect 46 131 47 132 
<< m1 >>
rect 64 131 65 132 
<< m1 >>
rect 88 131 89 132 
<< m1 >>
rect 92 131 93 132 
<< m1 >>
rect 100 131 101 132 
<< m1 >>
rect 109 131 110 132 
<< m1 >>
rect 114 131 115 132 
<< m1 >>
rect 115 131 116 132 
<< m1 >>
rect 116 131 117 132 
<< m2 >>
rect 116 131 117 132 
<< m2c >>
rect 116 131 117 132 
<< m1 >>
rect 116 131 117 132 
<< m2 >>
rect 116 131 117 132 
<< m2 >>
rect 117 131 118 132 
<< m1 >>
rect 118 131 119 132 
<< m2 >>
rect 118 131 119 132 
<< m2 >>
rect 119 131 120 132 
<< m1 >>
rect 120 131 121 132 
<< m2 >>
rect 120 131 121 132 
<< m2c >>
rect 120 131 121 132 
<< m1 >>
rect 120 131 121 132 
<< m2 >>
rect 120 131 121 132 
<< m1 >>
rect 121 131 122 132 
<< m1 >>
rect 122 131 123 132 
<< m2 >>
rect 122 131 123 132 
<< m2c >>
rect 122 131 123 132 
<< m1 >>
rect 122 131 123 132 
<< m2 >>
rect 122 131 123 132 
<< m2 >>
rect 123 131 124 132 
<< m1 >>
rect 124 131 125 132 
<< m2 >>
rect 124 131 125 132 
<< m2 >>
rect 125 131 126 132 
<< m1 >>
rect 126 131 127 132 
<< m2 >>
rect 126 131 127 132 
<< m1 >>
rect 127 131 128 132 
<< m2 >>
rect 127 131 128 132 
<< m2c >>
rect 127 131 128 132 
<< m1 >>
rect 127 131 128 132 
<< m2 >>
rect 127 131 128 132 
<< m2 >>
rect 128 131 129 132 
<< m1 >>
rect 129 131 130 132 
<< m2 >>
rect 129 131 130 132 
<< m2 >>
rect 130 131 131 132 
<< m1 >>
rect 131 131 132 132 
<< m2 >>
rect 131 131 132 132 
<< m2 >>
rect 132 131 133 132 
<< m1 >>
rect 133 131 134 132 
<< m2 >>
rect 133 131 134 132 
<< m2 >>
rect 134 131 135 132 
<< m2 >>
rect 135 131 136 132 
<< m1 >>
rect 136 131 137 132 
<< m2 >>
rect 136 131 137 132 
<< m2 >>
rect 137 131 138 132 
<< m1 >>
rect 138 131 139 132 
<< m2 >>
rect 138 131 139 132 
<< m2c >>
rect 138 131 139 132 
<< m1 >>
rect 138 131 139 132 
<< m2 >>
rect 138 131 139 132 
<< m1 >>
rect 139 131 140 132 
<< m1 >>
rect 140 131 141 132 
<< m1 >>
rect 141 131 142 132 
<< m1 >>
rect 142 131 143 132 
<< m1 >>
rect 143 131 144 132 
<< m2 >>
rect 143 131 144 132 
<< m2c >>
rect 143 131 144 132 
<< m1 >>
rect 143 131 144 132 
<< m2 >>
rect 143 131 144 132 
<< m2 >>
rect 144 131 145 132 
<< m1 >>
rect 145 131 146 132 
<< m2 >>
rect 145 131 146 132 
<< m2 >>
rect 146 131 147 132 
<< m1 >>
rect 147 131 148 132 
<< m2 >>
rect 147 131 148 132 
<< m2c >>
rect 147 131 148 132 
<< m1 >>
rect 147 131 148 132 
<< m2 >>
rect 147 131 148 132 
<< m1 >>
rect 148 131 149 132 
<< m1 >>
rect 149 131 150 132 
<< m1 >>
rect 150 131 151 132 
<< m1 >>
rect 151 131 152 132 
<< m1 >>
rect 152 131 153 132 
<< m1 >>
rect 153 131 154 132 
<< m1 >>
rect 154 131 155 132 
<< m1 >>
rect 155 131 156 132 
<< m1 >>
rect 156 131 157 132 
<< m1 >>
rect 157 131 158 132 
<< m1 >>
rect 158 131 159 132 
<< m1 >>
rect 159 131 160 132 
<< m1 >>
rect 160 131 161 132 
<< m1 >>
rect 161 131 162 132 
<< m1 >>
rect 163 131 164 132 
<< m1 >>
rect 199 131 200 132 
<< m1 >>
rect 217 131 218 132 
<< m2 >>
rect 217 131 218 132 
<< m1 >>
rect 226 131 227 132 
<< m1 >>
rect 235 131 236 132 
<< m1 >>
rect 244 131 245 132 
<< m1 >>
rect 265 131 266 132 
<< m2 >>
rect 278 131 279 132 
<< m2 >>
rect 280 131 281 132 
<< m2 >>
rect 282 131 283 132 
<< m1 >>
rect 283 131 284 132 
<< m1 >>
rect 334 131 335 132 
<< m1 >>
rect 343 131 344 132 
<< m1 >>
rect 345 131 346 132 
<< m2 >>
rect 358 131 359 132 
<< m2 >>
rect 361 131 362 132 
<< m2 >>
rect 366 131 367 132 
<< m2 >>
rect 370 131 371 132 
<< m2 >>
rect 379 131 380 132 
<< m1 >>
rect 415 131 416 132 
<< m1 >>
rect 419 131 420 132 
<< m2 >>
rect 420 131 421 132 
<< m1 >>
rect 427 131 428 132 
<< m1 >>
rect 430 131 431 132 
<< m1 >>
rect 456 131 457 132 
<< m1 >>
rect 469 131 470 132 
<< m1 >>
rect 478 131 479 132 
<< m1 >>
rect 19 132 20 133 
<< m1 >>
rect 46 132 47 133 
<< m1 >>
rect 64 132 65 133 
<< m1 >>
rect 88 132 89 133 
<< m1 >>
rect 92 132 93 133 
<< m1 >>
rect 100 132 101 133 
<< m1 >>
rect 109 132 110 133 
<< m1 >>
rect 114 132 115 133 
<< m1 >>
rect 118 132 119 133 
<< m1 >>
rect 124 132 125 133 
<< m1 >>
rect 129 132 130 133 
<< m1 >>
rect 131 132 132 133 
<< m1 >>
rect 133 132 134 133 
<< m1 >>
rect 136 132 137 133 
<< m1 >>
rect 145 132 146 133 
<< m1 >>
rect 163 132 164 133 
<< m1 >>
rect 199 132 200 133 
<< m1 >>
rect 217 132 218 133 
<< m2 >>
rect 217 132 218 133 
<< m1 >>
rect 226 132 227 133 
<< m1 >>
rect 235 132 236 133 
<< m1 >>
rect 244 132 245 133 
<< m1 >>
rect 265 132 266 133 
<< m1 >>
rect 278 132 279 133 
<< m2 >>
rect 278 132 279 133 
<< m2c >>
rect 278 132 279 133 
<< m1 >>
rect 278 132 279 133 
<< m2 >>
rect 278 132 279 133 
<< m1 >>
rect 280 132 281 133 
<< m2 >>
rect 280 132 281 133 
<< m2c >>
rect 280 132 281 133 
<< m1 >>
rect 280 132 281 133 
<< m2 >>
rect 280 132 281 133 
<< m2 >>
rect 282 132 283 133 
<< m1 >>
rect 283 132 284 133 
<< m1 >>
rect 334 132 335 133 
<< m1 >>
rect 343 132 344 133 
<< m1 >>
rect 345 132 346 133 
<< m1 >>
rect 346 132 347 133 
<< m1 >>
rect 347 132 348 133 
<< m1 >>
rect 348 132 349 133 
<< m1 >>
rect 349 132 350 133 
<< m1 >>
rect 350 132 351 133 
<< m1 >>
rect 351 132 352 133 
<< m1 >>
rect 352 132 353 133 
<< m1 >>
rect 353 132 354 133 
<< m1 >>
rect 354 132 355 133 
<< m1 >>
rect 355 132 356 133 
<< m1 >>
rect 356 132 357 133 
<< m1 >>
rect 357 132 358 133 
<< m1 >>
rect 358 132 359 133 
<< m2 >>
rect 358 132 359 133 
<< m1 >>
rect 359 132 360 133 
<< m1 >>
rect 360 132 361 133 
<< m1 >>
rect 361 132 362 133 
<< m2 >>
rect 361 132 362 133 
<< m1 >>
rect 362 132 363 133 
<< m1 >>
rect 363 132 364 133 
<< m1 >>
rect 364 132 365 133 
<< m1 >>
rect 365 132 366 133 
<< m1 >>
rect 366 132 367 133 
<< m2 >>
rect 366 132 367 133 
<< m1 >>
rect 367 132 368 133 
<< m1 >>
rect 368 132 369 133 
<< m1 >>
rect 369 132 370 133 
<< m1 >>
rect 370 132 371 133 
<< m2 >>
rect 370 132 371 133 
<< m1 >>
rect 371 132 372 133 
<< m1 >>
rect 372 132 373 133 
<< m1 >>
rect 373 132 374 133 
<< m1 >>
rect 374 132 375 133 
<< m1 >>
rect 375 132 376 133 
<< m1 >>
rect 376 132 377 133 
<< m1 >>
rect 377 132 378 133 
<< m1 >>
rect 378 132 379 133 
<< m1 >>
rect 379 132 380 133 
<< m2 >>
rect 379 132 380 133 
<< m1 >>
rect 415 132 416 133 
<< m1 >>
rect 419 132 420 133 
<< m2 >>
rect 420 132 421 133 
<< m1 >>
rect 427 132 428 133 
<< m1 >>
rect 430 132 431 133 
<< m1 >>
rect 456 132 457 133 
<< m1 >>
rect 469 132 470 133 
<< m1 >>
rect 478 132 479 133 
<< m1 >>
rect 19 133 20 134 
<< m1 >>
rect 46 133 47 134 
<< m1 >>
rect 64 133 65 134 
<< m1 >>
rect 88 133 89 134 
<< m2 >>
rect 88 133 89 134 
<< m2c >>
rect 88 133 89 134 
<< m1 >>
rect 88 133 89 134 
<< m2 >>
rect 88 133 89 134 
<< m1 >>
rect 92 133 93 134 
<< m2 >>
rect 92 133 93 134 
<< m2c >>
rect 92 133 93 134 
<< m1 >>
rect 92 133 93 134 
<< m2 >>
rect 92 133 93 134 
<< m1 >>
rect 100 133 101 134 
<< m1 >>
rect 109 133 110 134 
<< m1 >>
rect 114 133 115 134 
<< m1 >>
rect 118 133 119 134 
<< m1 >>
rect 124 133 125 134 
<< m1 >>
rect 129 133 130 134 
<< m1 >>
rect 131 133 132 134 
<< m1 >>
rect 133 133 134 134 
<< m1 >>
rect 136 133 137 134 
<< m1 >>
rect 145 133 146 134 
<< m1 >>
rect 163 133 164 134 
<< m1 >>
rect 199 133 200 134 
<< m1 >>
rect 217 133 218 134 
<< m2 >>
rect 217 133 218 134 
<< m1 >>
rect 226 133 227 134 
<< m1 >>
rect 235 133 236 134 
<< m1 >>
rect 244 133 245 134 
<< m1 >>
rect 265 133 266 134 
<< m1 >>
rect 278 133 279 134 
<< m1 >>
rect 280 133 281 134 
<< m2 >>
rect 282 133 283 134 
<< m1 >>
rect 283 133 284 134 
<< m1 >>
rect 334 133 335 134 
<< m1 >>
rect 343 133 344 134 
<< m2 >>
rect 358 133 359 134 
<< m2 >>
rect 361 133 362 134 
<< m2 >>
rect 366 133 367 134 
<< m2 >>
rect 370 133 371 134 
<< m1 >>
rect 379 133 380 134 
<< m2 >>
rect 379 133 380 134 
<< m1 >>
rect 415 133 416 134 
<< m1 >>
rect 419 133 420 134 
<< m2 >>
rect 420 133 421 134 
<< m1 >>
rect 427 133 428 134 
<< m1 >>
rect 430 133 431 134 
<< m1 >>
rect 456 133 457 134 
<< m1 >>
rect 469 133 470 134 
<< m1 >>
rect 478 133 479 134 
<< m1 >>
rect 19 134 20 135 
<< m1 >>
rect 46 134 47 135 
<< m1 >>
rect 64 134 65 135 
<< m2 >>
rect 88 134 89 135 
<< m2 >>
rect 92 134 93 135 
<< m2 >>
rect 93 134 94 135 
<< m2 >>
rect 94 134 95 135 
<< m2 >>
rect 95 134 96 135 
<< m2 >>
rect 96 134 97 135 
<< m2 >>
rect 97 134 98 135 
<< m1 >>
rect 100 134 101 135 
<< m1 >>
rect 109 134 110 135 
<< m1 >>
rect 114 134 115 135 
<< m1 >>
rect 118 134 119 135 
<< m1 >>
rect 124 134 125 135 
<< m1 >>
rect 129 134 130 135 
<< m1 >>
rect 131 134 132 135 
<< m1 >>
rect 133 134 134 135 
<< m1 >>
rect 136 134 137 135 
<< m1 >>
rect 145 134 146 135 
<< m1 >>
rect 163 134 164 135 
<< m1 >>
rect 199 134 200 135 
<< m1 >>
rect 217 134 218 135 
<< m2 >>
rect 217 134 218 135 
<< m1 >>
rect 226 134 227 135 
<< m1 >>
rect 235 134 236 135 
<< m1 >>
rect 244 134 245 135 
<< m1 >>
rect 265 134 266 135 
<< m1 >>
rect 278 134 279 135 
<< m1 >>
rect 280 134 281 135 
<< m2 >>
rect 280 134 281 135 
<< m2 >>
rect 281 134 282 135 
<< m2 >>
rect 282 134 283 135 
<< m1 >>
rect 283 134 284 135 
<< m1 >>
rect 334 134 335 135 
<< m1 >>
rect 343 134 344 135 
<< m1 >>
rect 358 134 359 135 
<< m2 >>
rect 358 134 359 135 
<< m2c >>
rect 358 134 359 135 
<< m1 >>
rect 358 134 359 135 
<< m2 >>
rect 358 134 359 135 
<< m1 >>
rect 361 134 362 135 
<< m2 >>
rect 361 134 362 135 
<< m2c >>
rect 361 134 362 135 
<< m1 >>
rect 361 134 362 135 
<< m2 >>
rect 361 134 362 135 
<< m1 >>
rect 366 134 367 135 
<< m2 >>
rect 366 134 367 135 
<< m2c >>
rect 366 134 367 135 
<< m1 >>
rect 366 134 367 135 
<< m2 >>
rect 366 134 367 135 
<< m1 >>
rect 370 134 371 135 
<< m2 >>
rect 370 134 371 135 
<< m2c >>
rect 370 134 371 135 
<< m1 >>
rect 370 134 371 135 
<< m2 >>
rect 370 134 371 135 
<< m1 >>
rect 379 134 380 135 
<< m2 >>
rect 379 134 380 135 
<< m1 >>
rect 415 134 416 135 
<< m1 >>
rect 419 134 420 135 
<< m2 >>
rect 420 134 421 135 
<< m1 >>
rect 427 134 428 135 
<< m1 >>
rect 430 134 431 135 
<< m1 >>
rect 456 134 457 135 
<< m1 >>
rect 469 134 470 135 
<< m1 >>
rect 478 134 479 135 
<< m1 >>
rect 13 135 14 136 
<< m1 >>
rect 14 135 15 136 
<< m1 >>
rect 15 135 16 136 
<< m1 >>
rect 16 135 17 136 
<< m1 >>
rect 17 135 18 136 
<< m1 >>
rect 18 135 19 136 
<< m1 >>
rect 19 135 20 136 
<< m1 >>
rect 46 135 47 136 
<< m1 >>
rect 64 135 65 136 
<< m1 >>
rect 67 135 68 136 
<< m1 >>
rect 68 135 69 136 
<< m1 >>
rect 69 135 70 136 
<< m1 >>
rect 70 135 71 136 
<< m1 >>
rect 71 135 72 136 
<< m1 >>
rect 72 135 73 136 
<< m1 >>
rect 73 135 74 136 
<< m1 >>
rect 74 135 75 136 
<< m1 >>
rect 75 135 76 136 
<< m1 >>
rect 76 135 77 136 
<< m1 >>
rect 77 135 78 136 
<< m1 >>
rect 78 135 79 136 
<< m1 >>
rect 79 135 80 136 
<< m1 >>
rect 80 135 81 136 
<< m1 >>
rect 81 135 82 136 
<< m1 >>
rect 82 135 83 136 
<< m1 >>
rect 83 135 84 136 
<< m1 >>
rect 84 135 85 136 
<< m1 >>
rect 85 135 86 136 
<< m1 >>
rect 86 135 87 136 
<< m1 >>
rect 87 135 88 136 
<< m1 >>
rect 88 135 89 136 
<< m2 >>
rect 88 135 89 136 
<< m1 >>
rect 89 135 90 136 
<< m1 >>
rect 90 135 91 136 
<< m1 >>
rect 91 135 92 136 
<< m1 >>
rect 92 135 93 136 
<< m1 >>
rect 93 135 94 136 
<< m1 >>
rect 94 135 95 136 
<< m1 >>
rect 95 135 96 136 
<< m1 >>
rect 96 135 97 136 
<< m1 >>
rect 97 135 98 136 
<< m2 >>
rect 97 135 98 136 
<< m1 >>
rect 98 135 99 136 
<< m1 >>
rect 100 135 101 136 
<< m1 >>
rect 109 135 110 136 
<< m1 >>
rect 114 135 115 136 
<< m1 >>
rect 118 135 119 136 
<< m1 >>
rect 124 135 125 136 
<< m1 >>
rect 125 135 126 136 
<< m1 >>
rect 126 135 127 136 
<< m1 >>
rect 127 135 128 136 
<< m1 >>
rect 129 135 130 136 
<< m1 >>
rect 131 135 132 136 
<< m1 >>
rect 133 135 134 136 
<< m1 >>
rect 136 135 137 136 
<< m1 >>
rect 145 135 146 136 
<< m1 >>
rect 163 135 164 136 
<< m1 >>
rect 199 135 200 136 
<< m1 >>
rect 217 135 218 136 
<< m2 >>
rect 217 135 218 136 
<< m1 >>
rect 226 135 227 136 
<< m1 >>
rect 235 135 236 136 
<< m1 >>
rect 244 135 245 136 
<< m1 >>
rect 265 135 266 136 
<< m1 >>
rect 278 135 279 136 
<< m1 >>
rect 280 135 281 136 
<< m2 >>
rect 280 135 281 136 
<< m1 >>
rect 283 135 284 136 
<< m1 >>
rect 334 135 335 136 
<< m1 >>
rect 343 135 344 136 
<< m1 >>
rect 358 135 359 136 
<< m1 >>
rect 361 135 362 136 
<< m1 >>
rect 366 135 367 136 
<< m1 >>
rect 370 135 371 136 
<< m1 >>
rect 379 135 380 136 
<< m2 >>
rect 379 135 380 136 
<< m1 >>
rect 415 135 416 136 
<< m1 >>
rect 419 135 420 136 
<< m2 >>
rect 420 135 421 136 
<< m1 >>
rect 427 135 428 136 
<< m1 >>
rect 430 135 431 136 
<< m1 >>
rect 431 135 432 136 
<< m1 >>
rect 432 135 433 136 
<< m1 >>
rect 433 135 434 136 
<< m1 >>
rect 434 135 435 136 
<< m1 >>
rect 435 135 436 136 
<< m1 >>
rect 436 135 437 136 
<< m1 >>
rect 437 135 438 136 
<< m1 >>
rect 438 135 439 136 
<< m1 >>
rect 439 135 440 136 
<< m1 >>
rect 440 135 441 136 
<< m1 >>
rect 441 135 442 136 
<< m1 >>
rect 442 135 443 136 
<< m1 >>
rect 456 135 457 136 
<< m1 >>
rect 469 135 470 136 
<< m1 >>
rect 478 135 479 136 
<< m1 >>
rect 13 136 14 137 
<< m1 >>
rect 34 136 35 137 
<< m1 >>
rect 35 136 36 137 
<< m1 >>
rect 36 136 37 137 
<< m1 >>
rect 37 136 38 137 
<< m1 >>
rect 46 136 47 137 
<< m1 >>
rect 64 136 65 137 
<< m1 >>
rect 67 136 68 137 
<< m2 >>
rect 88 136 89 137 
<< m2 >>
rect 97 136 98 137 
<< m1 >>
rect 98 136 99 137 
<< m1 >>
rect 100 136 101 137 
<< m1 >>
rect 109 136 110 137 
<< m1 >>
rect 114 136 115 137 
<< m1 >>
rect 118 136 119 137 
<< m2 >>
rect 118 136 119 137 
<< m2 >>
rect 119 136 120 137 
<< m1 >>
rect 120 136 121 137 
<< m2 >>
rect 120 136 121 137 
<< m2c >>
rect 120 136 121 137 
<< m1 >>
rect 120 136 121 137 
<< m2 >>
rect 120 136 121 137 
<< m1 >>
rect 121 136 122 137 
<< m1 >>
rect 127 136 128 137 
<< m1 >>
rect 129 136 130 137 
<< m1 >>
rect 131 136 132 137 
<< m1 >>
rect 133 136 134 137 
<< m1 >>
rect 136 136 137 137 
<< m1 >>
rect 145 136 146 137 
<< m1 >>
rect 163 136 164 137 
<< m1 >>
rect 199 136 200 137 
<< m1 >>
rect 217 136 218 137 
<< m2 >>
rect 217 136 218 137 
<< m1 >>
rect 226 136 227 137 
<< m1 >>
rect 235 136 236 137 
<< m1 >>
rect 244 136 245 137 
<< m1 >>
rect 265 136 266 137 
<< m1 >>
rect 278 136 279 137 
<< m1 >>
rect 280 136 281 137 
<< m2 >>
rect 280 136 281 137 
<< m1 >>
rect 283 136 284 137 
<< m1 >>
rect 334 136 335 137 
<< m1 >>
rect 343 136 344 137 
<< m1 >>
rect 358 136 359 137 
<< m1 >>
rect 361 136 362 137 
<< m1 >>
rect 366 136 367 137 
<< m1 >>
rect 370 136 371 137 
<< m1 >>
rect 379 136 380 137 
<< m2 >>
rect 379 136 380 137 
<< m1 >>
rect 415 136 416 137 
<< m1 >>
rect 419 136 420 137 
<< m2 >>
rect 420 136 421 137 
<< m1 >>
rect 427 136 428 137 
<< m1 >>
rect 442 136 443 137 
<< m1 >>
rect 456 136 457 137 
<< m1 >>
rect 469 136 470 137 
<< m1 >>
rect 478 136 479 137 
<< m1 >>
rect 13 137 14 138 
<< m1 >>
rect 34 137 35 138 
<< m1 >>
rect 37 137 38 138 
<< m1 >>
rect 46 137 47 138 
<< m1 >>
rect 64 137 65 138 
<< m1 >>
rect 67 137 68 138 
<< m1 >>
rect 88 137 89 138 
<< m2 >>
rect 88 137 89 138 
<< m2c >>
rect 88 137 89 138 
<< m1 >>
rect 88 137 89 138 
<< m2 >>
rect 88 137 89 138 
<< m2 >>
rect 97 137 98 138 
<< m1 >>
rect 98 137 99 138 
<< m1 >>
rect 100 137 101 138 
<< m1 >>
rect 109 137 110 138 
<< m1 >>
rect 114 137 115 138 
<< m1 >>
rect 118 137 119 138 
<< m2 >>
rect 118 137 119 138 
<< m1 >>
rect 121 137 122 138 
<< m1 >>
rect 127 137 128 138 
<< m1 >>
rect 129 137 130 138 
<< m1 >>
rect 131 137 132 138 
<< m1 >>
rect 133 137 134 138 
<< m1 >>
rect 136 137 137 138 
<< m1 >>
rect 145 137 146 138 
<< m1 >>
rect 163 137 164 138 
<< m1 >>
rect 199 137 200 138 
<< m1 >>
rect 217 137 218 138 
<< m2 >>
rect 217 137 218 138 
<< m1 >>
rect 226 137 227 138 
<< m1 >>
rect 235 137 236 138 
<< m1 >>
rect 244 137 245 138 
<< m1 >>
rect 265 137 266 138 
<< m1 >>
rect 278 137 279 138 
<< m1 >>
rect 280 137 281 138 
<< m2 >>
rect 280 137 281 138 
<< m1 >>
rect 283 137 284 138 
<< m1 >>
rect 334 137 335 138 
<< m1 >>
rect 343 137 344 138 
<< m1 >>
rect 358 137 359 138 
<< m1 >>
rect 361 137 362 138 
<< m1 >>
rect 366 137 367 138 
<< m1 >>
rect 370 137 371 138 
<< m1 >>
rect 379 137 380 138 
<< m2 >>
rect 379 137 380 138 
<< m1 >>
rect 415 137 416 138 
<< m1 >>
rect 419 137 420 138 
<< m2 >>
rect 420 137 421 138 
<< m1 >>
rect 427 137 428 138 
<< m1 >>
rect 442 137 443 138 
<< m1 >>
rect 456 137 457 138 
<< m1 >>
rect 469 137 470 138 
<< m1 >>
rect 478 137 479 138 
<< pdiffusion >>
rect 12 138 13 139 
<< m1 >>
rect 13 138 14 139 
<< pdiffusion >>
rect 13 138 14 139 
<< pdiffusion >>
rect 14 138 15 139 
<< pdiffusion >>
rect 15 138 16 139 
<< pdiffusion >>
rect 16 138 17 139 
<< pdiffusion >>
rect 17 138 18 139 
<< pdiffusion >>
rect 30 138 31 139 
<< pdiffusion >>
rect 31 138 32 139 
<< pdiffusion >>
rect 32 138 33 139 
<< pdiffusion >>
rect 33 138 34 139 
<< m1 >>
rect 34 138 35 139 
<< pdiffusion >>
rect 34 138 35 139 
<< pdiffusion >>
rect 35 138 36 139 
<< m1 >>
rect 37 138 38 139 
<< m1 >>
rect 46 138 47 139 
<< pdiffusion >>
rect 48 138 49 139 
<< pdiffusion >>
rect 49 138 50 139 
<< pdiffusion >>
rect 50 138 51 139 
<< pdiffusion >>
rect 51 138 52 139 
<< pdiffusion >>
rect 52 138 53 139 
<< pdiffusion >>
rect 53 138 54 139 
<< m1 >>
rect 64 138 65 139 
<< pdiffusion >>
rect 66 138 67 139 
<< m1 >>
rect 67 138 68 139 
<< pdiffusion >>
rect 67 138 68 139 
<< pdiffusion >>
rect 68 138 69 139 
<< pdiffusion >>
rect 69 138 70 139 
<< pdiffusion >>
rect 70 138 71 139 
<< pdiffusion >>
rect 71 138 72 139 
<< m1 >>
rect 88 138 89 139 
<< m2 >>
rect 97 138 98 139 
<< m1 >>
rect 98 138 99 139 
<< m1 >>
rect 100 138 101 139 
<< pdiffusion >>
rect 102 138 103 139 
<< pdiffusion >>
rect 103 138 104 139 
<< pdiffusion >>
rect 104 138 105 139 
<< pdiffusion >>
rect 105 138 106 139 
<< pdiffusion >>
rect 106 138 107 139 
<< pdiffusion >>
rect 107 138 108 139 
<< m1 >>
rect 109 138 110 139 
<< m1 >>
rect 114 138 115 139 
<< m1 >>
rect 118 138 119 139 
<< m2 >>
rect 118 138 119 139 
<< pdiffusion >>
rect 120 138 121 139 
<< m1 >>
rect 121 138 122 139 
<< pdiffusion >>
rect 121 138 122 139 
<< pdiffusion >>
rect 122 138 123 139 
<< pdiffusion >>
rect 123 138 124 139 
<< pdiffusion >>
rect 124 138 125 139 
<< pdiffusion >>
rect 125 138 126 139 
<< m1 >>
rect 127 138 128 139 
<< m1 >>
rect 129 138 130 139 
<< m1 >>
rect 131 138 132 139 
<< m1 >>
rect 133 138 134 139 
<< m1 >>
rect 136 138 137 139 
<< pdiffusion >>
rect 138 138 139 139 
<< pdiffusion >>
rect 139 138 140 139 
<< pdiffusion >>
rect 140 138 141 139 
<< pdiffusion >>
rect 141 138 142 139 
<< pdiffusion >>
rect 142 138 143 139 
<< pdiffusion >>
rect 143 138 144 139 
<< m1 >>
rect 145 138 146 139 
<< pdiffusion >>
rect 156 138 157 139 
<< pdiffusion >>
rect 157 138 158 139 
<< pdiffusion >>
rect 158 138 159 139 
<< pdiffusion >>
rect 159 138 160 139 
<< pdiffusion >>
rect 160 138 161 139 
<< pdiffusion >>
rect 161 138 162 139 
<< m1 >>
rect 163 138 164 139 
<< pdiffusion >>
rect 174 138 175 139 
<< pdiffusion >>
rect 175 138 176 139 
<< pdiffusion >>
rect 176 138 177 139 
<< pdiffusion >>
rect 177 138 178 139 
<< pdiffusion >>
rect 178 138 179 139 
<< pdiffusion >>
rect 179 138 180 139 
<< pdiffusion >>
rect 192 138 193 139 
<< pdiffusion >>
rect 193 138 194 139 
<< pdiffusion >>
rect 194 138 195 139 
<< pdiffusion >>
rect 195 138 196 139 
<< pdiffusion >>
rect 196 138 197 139 
<< pdiffusion >>
rect 197 138 198 139 
<< m1 >>
rect 199 138 200 139 
<< pdiffusion >>
rect 210 138 211 139 
<< pdiffusion >>
rect 211 138 212 139 
<< pdiffusion >>
rect 212 138 213 139 
<< pdiffusion >>
rect 213 138 214 139 
<< pdiffusion >>
rect 214 138 215 139 
<< pdiffusion >>
rect 215 138 216 139 
<< m1 >>
rect 217 138 218 139 
<< m2 >>
rect 217 138 218 139 
<< m1 >>
rect 226 138 227 139 
<< pdiffusion >>
rect 228 138 229 139 
<< pdiffusion >>
rect 229 138 230 139 
<< pdiffusion >>
rect 230 138 231 139 
<< pdiffusion >>
rect 231 138 232 139 
<< pdiffusion >>
rect 232 138 233 139 
<< pdiffusion >>
rect 233 138 234 139 
<< m1 >>
rect 235 138 236 139 
<< m1 >>
rect 244 138 245 139 
<< pdiffusion >>
rect 246 138 247 139 
<< pdiffusion >>
rect 247 138 248 139 
<< pdiffusion >>
rect 248 138 249 139 
<< pdiffusion >>
rect 249 138 250 139 
<< pdiffusion >>
rect 250 138 251 139 
<< pdiffusion >>
rect 251 138 252 139 
<< pdiffusion >>
rect 264 138 265 139 
<< m1 >>
rect 265 138 266 139 
<< pdiffusion >>
rect 265 138 266 139 
<< pdiffusion >>
rect 266 138 267 139 
<< pdiffusion >>
rect 267 138 268 139 
<< pdiffusion >>
rect 268 138 269 139 
<< pdiffusion >>
rect 269 138 270 139 
<< m1 >>
rect 278 138 279 139 
<< m1 >>
rect 280 138 281 139 
<< m2 >>
rect 280 138 281 139 
<< pdiffusion >>
rect 282 138 283 139 
<< m1 >>
rect 283 138 284 139 
<< pdiffusion >>
rect 283 138 284 139 
<< pdiffusion >>
rect 284 138 285 139 
<< pdiffusion >>
rect 285 138 286 139 
<< pdiffusion >>
rect 286 138 287 139 
<< pdiffusion >>
rect 287 138 288 139 
<< pdiffusion >>
rect 300 138 301 139 
<< pdiffusion >>
rect 301 138 302 139 
<< pdiffusion >>
rect 302 138 303 139 
<< pdiffusion >>
rect 303 138 304 139 
<< pdiffusion >>
rect 304 138 305 139 
<< pdiffusion >>
rect 305 138 306 139 
<< m1 >>
rect 334 138 335 139 
<< m1 >>
rect 343 138 344 139 
<< pdiffusion >>
rect 354 138 355 139 
<< pdiffusion >>
rect 355 138 356 139 
<< pdiffusion >>
rect 356 138 357 139 
<< pdiffusion >>
rect 357 138 358 139 
<< m1 >>
rect 358 138 359 139 
<< pdiffusion >>
rect 358 138 359 139 
<< pdiffusion >>
rect 359 138 360 139 
<< m1 >>
rect 361 138 362 139 
<< m1 >>
rect 366 138 367 139 
<< m1 >>
rect 370 138 371 139 
<< pdiffusion >>
rect 372 138 373 139 
<< pdiffusion >>
rect 373 138 374 139 
<< pdiffusion >>
rect 374 138 375 139 
<< pdiffusion >>
rect 375 138 376 139 
<< pdiffusion >>
rect 376 138 377 139 
<< pdiffusion >>
rect 377 138 378 139 
<< m1 >>
rect 379 138 380 139 
<< m2 >>
rect 379 138 380 139 
<< pdiffusion >>
rect 390 138 391 139 
<< pdiffusion >>
rect 391 138 392 139 
<< pdiffusion >>
rect 392 138 393 139 
<< pdiffusion >>
rect 393 138 394 139 
<< pdiffusion >>
rect 394 138 395 139 
<< pdiffusion >>
rect 395 138 396 139 
<< pdiffusion >>
rect 408 138 409 139 
<< pdiffusion >>
rect 409 138 410 139 
<< pdiffusion >>
rect 410 138 411 139 
<< pdiffusion >>
rect 411 138 412 139 
<< pdiffusion >>
rect 412 138 413 139 
<< pdiffusion >>
rect 413 138 414 139 
<< m1 >>
rect 415 138 416 139 
<< m1 >>
rect 419 138 420 139 
<< m2 >>
rect 420 138 421 139 
<< pdiffusion >>
rect 426 138 427 139 
<< m1 >>
rect 427 138 428 139 
<< pdiffusion >>
rect 427 138 428 139 
<< pdiffusion >>
rect 428 138 429 139 
<< pdiffusion >>
rect 429 138 430 139 
<< pdiffusion >>
rect 430 138 431 139 
<< pdiffusion >>
rect 431 138 432 139 
<< m1 >>
rect 442 138 443 139 
<< pdiffusion >>
rect 444 138 445 139 
<< pdiffusion >>
rect 445 138 446 139 
<< pdiffusion >>
rect 446 138 447 139 
<< pdiffusion >>
rect 447 138 448 139 
<< pdiffusion >>
rect 448 138 449 139 
<< pdiffusion >>
rect 449 138 450 139 
<< m1 >>
rect 456 138 457 139 
<< pdiffusion >>
rect 462 138 463 139 
<< pdiffusion >>
rect 463 138 464 139 
<< pdiffusion >>
rect 464 138 465 139 
<< pdiffusion >>
rect 465 138 466 139 
<< pdiffusion >>
rect 466 138 467 139 
<< pdiffusion >>
rect 467 138 468 139 
<< m1 >>
rect 469 138 470 139 
<< m1 >>
rect 478 138 479 139 
<< pdiffusion >>
rect 498 138 499 139 
<< pdiffusion >>
rect 499 138 500 139 
<< pdiffusion >>
rect 500 138 501 139 
<< pdiffusion >>
rect 501 138 502 139 
<< pdiffusion >>
rect 502 138 503 139 
<< pdiffusion >>
rect 503 138 504 139 
<< pdiffusion >>
rect 516 138 517 139 
<< pdiffusion >>
rect 517 138 518 139 
<< pdiffusion >>
rect 518 138 519 139 
<< pdiffusion >>
rect 519 138 520 139 
<< pdiffusion >>
rect 520 138 521 139 
<< pdiffusion >>
rect 521 138 522 139 
<< pdiffusion >>
rect 12 139 13 140 
<< pdiffusion >>
rect 13 139 14 140 
<< pdiffusion >>
rect 14 139 15 140 
<< pdiffusion >>
rect 15 139 16 140 
<< pdiffusion >>
rect 16 139 17 140 
<< pdiffusion >>
rect 17 139 18 140 
<< pdiffusion >>
rect 30 139 31 140 
<< pdiffusion >>
rect 31 139 32 140 
<< pdiffusion >>
rect 32 139 33 140 
<< pdiffusion >>
rect 33 139 34 140 
<< pdiffusion >>
rect 34 139 35 140 
<< pdiffusion >>
rect 35 139 36 140 
<< m1 >>
rect 37 139 38 140 
<< m1 >>
rect 46 139 47 140 
<< pdiffusion >>
rect 48 139 49 140 
<< pdiffusion >>
rect 49 139 50 140 
<< pdiffusion >>
rect 50 139 51 140 
<< pdiffusion >>
rect 51 139 52 140 
<< pdiffusion >>
rect 52 139 53 140 
<< pdiffusion >>
rect 53 139 54 140 
<< m1 >>
rect 64 139 65 140 
<< pdiffusion >>
rect 66 139 67 140 
<< pdiffusion >>
rect 67 139 68 140 
<< pdiffusion >>
rect 68 139 69 140 
<< pdiffusion >>
rect 69 139 70 140 
<< pdiffusion >>
rect 70 139 71 140 
<< pdiffusion >>
rect 71 139 72 140 
<< m1 >>
rect 88 139 89 140 
<< m2 >>
rect 97 139 98 140 
<< m1 >>
rect 98 139 99 140 
<< m1 >>
rect 100 139 101 140 
<< pdiffusion >>
rect 102 139 103 140 
<< pdiffusion >>
rect 103 139 104 140 
<< pdiffusion >>
rect 104 139 105 140 
<< pdiffusion >>
rect 105 139 106 140 
<< pdiffusion >>
rect 106 139 107 140 
<< pdiffusion >>
rect 107 139 108 140 
<< m1 >>
rect 109 139 110 140 
<< m1 >>
rect 114 139 115 140 
<< m1 >>
rect 118 139 119 140 
<< m2 >>
rect 118 139 119 140 
<< pdiffusion >>
rect 120 139 121 140 
<< pdiffusion >>
rect 121 139 122 140 
<< pdiffusion >>
rect 122 139 123 140 
<< pdiffusion >>
rect 123 139 124 140 
<< pdiffusion >>
rect 124 139 125 140 
<< pdiffusion >>
rect 125 139 126 140 
<< m1 >>
rect 127 139 128 140 
<< m1 >>
rect 129 139 130 140 
<< m1 >>
rect 131 139 132 140 
<< m1 >>
rect 133 139 134 140 
<< m1 >>
rect 136 139 137 140 
<< pdiffusion >>
rect 138 139 139 140 
<< pdiffusion >>
rect 139 139 140 140 
<< pdiffusion >>
rect 140 139 141 140 
<< pdiffusion >>
rect 141 139 142 140 
<< pdiffusion >>
rect 142 139 143 140 
<< pdiffusion >>
rect 143 139 144 140 
<< m1 >>
rect 145 139 146 140 
<< pdiffusion >>
rect 156 139 157 140 
<< pdiffusion >>
rect 157 139 158 140 
<< pdiffusion >>
rect 158 139 159 140 
<< pdiffusion >>
rect 159 139 160 140 
<< pdiffusion >>
rect 160 139 161 140 
<< pdiffusion >>
rect 161 139 162 140 
<< m1 >>
rect 163 139 164 140 
<< pdiffusion >>
rect 174 139 175 140 
<< pdiffusion >>
rect 175 139 176 140 
<< pdiffusion >>
rect 176 139 177 140 
<< pdiffusion >>
rect 177 139 178 140 
<< pdiffusion >>
rect 178 139 179 140 
<< pdiffusion >>
rect 179 139 180 140 
<< pdiffusion >>
rect 192 139 193 140 
<< pdiffusion >>
rect 193 139 194 140 
<< pdiffusion >>
rect 194 139 195 140 
<< pdiffusion >>
rect 195 139 196 140 
<< pdiffusion >>
rect 196 139 197 140 
<< pdiffusion >>
rect 197 139 198 140 
<< m1 >>
rect 199 139 200 140 
<< pdiffusion >>
rect 210 139 211 140 
<< pdiffusion >>
rect 211 139 212 140 
<< pdiffusion >>
rect 212 139 213 140 
<< pdiffusion >>
rect 213 139 214 140 
<< pdiffusion >>
rect 214 139 215 140 
<< pdiffusion >>
rect 215 139 216 140 
<< m1 >>
rect 217 139 218 140 
<< m2 >>
rect 217 139 218 140 
<< m1 >>
rect 226 139 227 140 
<< pdiffusion >>
rect 228 139 229 140 
<< pdiffusion >>
rect 229 139 230 140 
<< pdiffusion >>
rect 230 139 231 140 
<< pdiffusion >>
rect 231 139 232 140 
<< pdiffusion >>
rect 232 139 233 140 
<< pdiffusion >>
rect 233 139 234 140 
<< m1 >>
rect 235 139 236 140 
<< m1 >>
rect 244 139 245 140 
<< pdiffusion >>
rect 246 139 247 140 
<< pdiffusion >>
rect 247 139 248 140 
<< pdiffusion >>
rect 248 139 249 140 
<< pdiffusion >>
rect 249 139 250 140 
<< pdiffusion >>
rect 250 139 251 140 
<< pdiffusion >>
rect 251 139 252 140 
<< pdiffusion >>
rect 264 139 265 140 
<< pdiffusion >>
rect 265 139 266 140 
<< pdiffusion >>
rect 266 139 267 140 
<< pdiffusion >>
rect 267 139 268 140 
<< pdiffusion >>
rect 268 139 269 140 
<< pdiffusion >>
rect 269 139 270 140 
<< m1 >>
rect 278 139 279 140 
<< m1 >>
rect 280 139 281 140 
<< m2 >>
rect 280 139 281 140 
<< pdiffusion >>
rect 282 139 283 140 
<< pdiffusion >>
rect 283 139 284 140 
<< pdiffusion >>
rect 284 139 285 140 
<< pdiffusion >>
rect 285 139 286 140 
<< pdiffusion >>
rect 286 139 287 140 
<< pdiffusion >>
rect 287 139 288 140 
<< pdiffusion >>
rect 300 139 301 140 
<< pdiffusion >>
rect 301 139 302 140 
<< pdiffusion >>
rect 302 139 303 140 
<< pdiffusion >>
rect 303 139 304 140 
<< pdiffusion >>
rect 304 139 305 140 
<< pdiffusion >>
rect 305 139 306 140 
<< m1 >>
rect 334 139 335 140 
<< m1 >>
rect 343 139 344 140 
<< pdiffusion >>
rect 354 139 355 140 
<< pdiffusion >>
rect 355 139 356 140 
<< pdiffusion >>
rect 356 139 357 140 
<< pdiffusion >>
rect 357 139 358 140 
<< pdiffusion >>
rect 358 139 359 140 
<< pdiffusion >>
rect 359 139 360 140 
<< m1 >>
rect 361 139 362 140 
<< m1 >>
rect 366 139 367 140 
<< m1 >>
rect 370 139 371 140 
<< pdiffusion >>
rect 372 139 373 140 
<< pdiffusion >>
rect 373 139 374 140 
<< pdiffusion >>
rect 374 139 375 140 
<< pdiffusion >>
rect 375 139 376 140 
<< pdiffusion >>
rect 376 139 377 140 
<< pdiffusion >>
rect 377 139 378 140 
<< m1 >>
rect 379 139 380 140 
<< m2 >>
rect 379 139 380 140 
<< pdiffusion >>
rect 390 139 391 140 
<< pdiffusion >>
rect 391 139 392 140 
<< pdiffusion >>
rect 392 139 393 140 
<< pdiffusion >>
rect 393 139 394 140 
<< pdiffusion >>
rect 394 139 395 140 
<< pdiffusion >>
rect 395 139 396 140 
<< pdiffusion >>
rect 408 139 409 140 
<< pdiffusion >>
rect 409 139 410 140 
<< pdiffusion >>
rect 410 139 411 140 
<< pdiffusion >>
rect 411 139 412 140 
<< pdiffusion >>
rect 412 139 413 140 
<< pdiffusion >>
rect 413 139 414 140 
<< m1 >>
rect 415 139 416 140 
<< m1 >>
rect 419 139 420 140 
<< m2 >>
rect 420 139 421 140 
<< pdiffusion >>
rect 426 139 427 140 
<< pdiffusion >>
rect 427 139 428 140 
<< pdiffusion >>
rect 428 139 429 140 
<< pdiffusion >>
rect 429 139 430 140 
<< pdiffusion >>
rect 430 139 431 140 
<< pdiffusion >>
rect 431 139 432 140 
<< m1 >>
rect 442 139 443 140 
<< pdiffusion >>
rect 444 139 445 140 
<< pdiffusion >>
rect 445 139 446 140 
<< pdiffusion >>
rect 446 139 447 140 
<< pdiffusion >>
rect 447 139 448 140 
<< pdiffusion >>
rect 448 139 449 140 
<< pdiffusion >>
rect 449 139 450 140 
<< m1 >>
rect 456 139 457 140 
<< pdiffusion >>
rect 462 139 463 140 
<< pdiffusion >>
rect 463 139 464 140 
<< pdiffusion >>
rect 464 139 465 140 
<< pdiffusion >>
rect 465 139 466 140 
<< pdiffusion >>
rect 466 139 467 140 
<< pdiffusion >>
rect 467 139 468 140 
<< m1 >>
rect 469 139 470 140 
<< m1 >>
rect 478 139 479 140 
<< pdiffusion >>
rect 498 139 499 140 
<< pdiffusion >>
rect 499 139 500 140 
<< pdiffusion >>
rect 500 139 501 140 
<< pdiffusion >>
rect 501 139 502 140 
<< pdiffusion >>
rect 502 139 503 140 
<< pdiffusion >>
rect 503 139 504 140 
<< pdiffusion >>
rect 516 139 517 140 
<< pdiffusion >>
rect 517 139 518 140 
<< pdiffusion >>
rect 518 139 519 140 
<< pdiffusion >>
rect 519 139 520 140 
<< pdiffusion >>
rect 520 139 521 140 
<< pdiffusion >>
rect 521 139 522 140 
<< pdiffusion >>
rect 12 140 13 141 
<< pdiffusion >>
rect 13 140 14 141 
<< pdiffusion >>
rect 14 140 15 141 
<< pdiffusion >>
rect 15 140 16 141 
<< pdiffusion >>
rect 16 140 17 141 
<< pdiffusion >>
rect 17 140 18 141 
<< pdiffusion >>
rect 30 140 31 141 
<< pdiffusion >>
rect 31 140 32 141 
<< pdiffusion >>
rect 32 140 33 141 
<< pdiffusion >>
rect 33 140 34 141 
<< pdiffusion >>
rect 34 140 35 141 
<< pdiffusion >>
rect 35 140 36 141 
<< m1 >>
rect 37 140 38 141 
<< m1 >>
rect 46 140 47 141 
<< pdiffusion >>
rect 48 140 49 141 
<< pdiffusion >>
rect 49 140 50 141 
<< pdiffusion >>
rect 50 140 51 141 
<< pdiffusion >>
rect 51 140 52 141 
<< pdiffusion >>
rect 52 140 53 141 
<< pdiffusion >>
rect 53 140 54 141 
<< m1 >>
rect 64 140 65 141 
<< pdiffusion >>
rect 66 140 67 141 
<< pdiffusion >>
rect 67 140 68 141 
<< pdiffusion >>
rect 68 140 69 141 
<< pdiffusion >>
rect 69 140 70 141 
<< pdiffusion >>
rect 70 140 71 141 
<< pdiffusion >>
rect 71 140 72 141 
<< m1 >>
rect 88 140 89 141 
<< m2 >>
rect 97 140 98 141 
<< m1 >>
rect 98 140 99 141 
<< m1 >>
rect 100 140 101 141 
<< pdiffusion >>
rect 102 140 103 141 
<< pdiffusion >>
rect 103 140 104 141 
<< pdiffusion >>
rect 104 140 105 141 
<< pdiffusion >>
rect 105 140 106 141 
<< pdiffusion >>
rect 106 140 107 141 
<< pdiffusion >>
rect 107 140 108 141 
<< m1 >>
rect 109 140 110 141 
<< m1 >>
rect 114 140 115 141 
<< m1 >>
rect 118 140 119 141 
<< m2 >>
rect 118 140 119 141 
<< pdiffusion >>
rect 120 140 121 141 
<< pdiffusion >>
rect 121 140 122 141 
<< pdiffusion >>
rect 122 140 123 141 
<< pdiffusion >>
rect 123 140 124 141 
<< pdiffusion >>
rect 124 140 125 141 
<< pdiffusion >>
rect 125 140 126 141 
<< m1 >>
rect 127 140 128 141 
<< m1 >>
rect 129 140 130 141 
<< m1 >>
rect 131 140 132 141 
<< m1 >>
rect 133 140 134 141 
<< m1 >>
rect 136 140 137 141 
<< pdiffusion >>
rect 138 140 139 141 
<< pdiffusion >>
rect 139 140 140 141 
<< pdiffusion >>
rect 140 140 141 141 
<< pdiffusion >>
rect 141 140 142 141 
<< pdiffusion >>
rect 142 140 143 141 
<< pdiffusion >>
rect 143 140 144 141 
<< m1 >>
rect 145 140 146 141 
<< pdiffusion >>
rect 156 140 157 141 
<< pdiffusion >>
rect 157 140 158 141 
<< pdiffusion >>
rect 158 140 159 141 
<< pdiffusion >>
rect 159 140 160 141 
<< pdiffusion >>
rect 160 140 161 141 
<< pdiffusion >>
rect 161 140 162 141 
<< m1 >>
rect 163 140 164 141 
<< pdiffusion >>
rect 174 140 175 141 
<< pdiffusion >>
rect 175 140 176 141 
<< pdiffusion >>
rect 176 140 177 141 
<< pdiffusion >>
rect 177 140 178 141 
<< pdiffusion >>
rect 178 140 179 141 
<< pdiffusion >>
rect 179 140 180 141 
<< pdiffusion >>
rect 192 140 193 141 
<< pdiffusion >>
rect 193 140 194 141 
<< pdiffusion >>
rect 194 140 195 141 
<< pdiffusion >>
rect 195 140 196 141 
<< pdiffusion >>
rect 196 140 197 141 
<< pdiffusion >>
rect 197 140 198 141 
<< m1 >>
rect 199 140 200 141 
<< pdiffusion >>
rect 210 140 211 141 
<< pdiffusion >>
rect 211 140 212 141 
<< pdiffusion >>
rect 212 140 213 141 
<< pdiffusion >>
rect 213 140 214 141 
<< pdiffusion >>
rect 214 140 215 141 
<< pdiffusion >>
rect 215 140 216 141 
<< m1 >>
rect 217 140 218 141 
<< m2 >>
rect 217 140 218 141 
<< m1 >>
rect 226 140 227 141 
<< pdiffusion >>
rect 228 140 229 141 
<< pdiffusion >>
rect 229 140 230 141 
<< pdiffusion >>
rect 230 140 231 141 
<< pdiffusion >>
rect 231 140 232 141 
<< pdiffusion >>
rect 232 140 233 141 
<< pdiffusion >>
rect 233 140 234 141 
<< m1 >>
rect 235 140 236 141 
<< m1 >>
rect 244 140 245 141 
<< pdiffusion >>
rect 246 140 247 141 
<< pdiffusion >>
rect 247 140 248 141 
<< pdiffusion >>
rect 248 140 249 141 
<< pdiffusion >>
rect 249 140 250 141 
<< pdiffusion >>
rect 250 140 251 141 
<< pdiffusion >>
rect 251 140 252 141 
<< pdiffusion >>
rect 264 140 265 141 
<< pdiffusion >>
rect 265 140 266 141 
<< pdiffusion >>
rect 266 140 267 141 
<< pdiffusion >>
rect 267 140 268 141 
<< pdiffusion >>
rect 268 140 269 141 
<< pdiffusion >>
rect 269 140 270 141 
<< m1 >>
rect 278 140 279 141 
<< m1 >>
rect 280 140 281 141 
<< m2 >>
rect 280 140 281 141 
<< pdiffusion >>
rect 282 140 283 141 
<< pdiffusion >>
rect 283 140 284 141 
<< pdiffusion >>
rect 284 140 285 141 
<< pdiffusion >>
rect 285 140 286 141 
<< pdiffusion >>
rect 286 140 287 141 
<< pdiffusion >>
rect 287 140 288 141 
<< pdiffusion >>
rect 300 140 301 141 
<< pdiffusion >>
rect 301 140 302 141 
<< pdiffusion >>
rect 302 140 303 141 
<< pdiffusion >>
rect 303 140 304 141 
<< pdiffusion >>
rect 304 140 305 141 
<< pdiffusion >>
rect 305 140 306 141 
<< m1 >>
rect 334 140 335 141 
<< m1 >>
rect 343 140 344 141 
<< pdiffusion >>
rect 354 140 355 141 
<< pdiffusion >>
rect 355 140 356 141 
<< pdiffusion >>
rect 356 140 357 141 
<< pdiffusion >>
rect 357 140 358 141 
<< pdiffusion >>
rect 358 140 359 141 
<< pdiffusion >>
rect 359 140 360 141 
<< m1 >>
rect 361 140 362 141 
<< m1 >>
rect 366 140 367 141 
<< m1 >>
rect 370 140 371 141 
<< pdiffusion >>
rect 372 140 373 141 
<< pdiffusion >>
rect 373 140 374 141 
<< pdiffusion >>
rect 374 140 375 141 
<< pdiffusion >>
rect 375 140 376 141 
<< pdiffusion >>
rect 376 140 377 141 
<< pdiffusion >>
rect 377 140 378 141 
<< m1 >>
rect 379 140 380 141 
<< m2 >>
rect 379 140 380 141 
<< pdiffusion >>
rect 390 140 391 141 
<< pdiffusion >>
rect 391 140 392 141 
<< pdiffusion >>
rect 392 140 393 141 
<< pdiffusion >>
rect 393 140 394 141 
<< pdiffusion >>
rect 394 140 395 141 
<< pdiffusion >>
rect 395 140 396 141 
<< pdiffusion >>
rect 408 140 409 141 
<< pdiffusion >>
rect 409 140 410 141 
<< pdiffusion >>
rect 410 140 411 141 
<< pdiffusion >>
rect 411 140 412 141 
<< pdiffusion >>
rect 412 140 413 141 
<< pdiffusion >>
rect 413 140 414 141 
<< m1 >>
rect 415 140 416 141 
<< m1 >>
rect 419 140 420 141 
<< m2 >>
rect 420 140 421 141 
<< pdiffusion >>
rect 426 140 427 141 
<< pdiffusion >>
rect 427 140 428 141 
<< pdiffusion >>
rect 428 140 429 141 
<< pdiffusion >>
rect 429 140 430 141 
<< pdiffusion >>
rect 430 140 431 141 
<< pdiffusion >>
rect 431 140 432 141 
<< m1 >>
rect 442 140 443 141 
<< pdiffusion >>
rect 444 140 445 141 
<< pdiffusion >>
rect 445 140 446 141 
<< pdiffusion >>
rect 446 140 447 141 
<< pdiffusion >>
rect 447 140 448 141 
<< pdiffusion >>
rect 448 140 449 141 
<< pdiffusion >>
rect 449 140 450 141 
<< m1 >>
rect 456 140 457 141 
<< pdiffusion >>
rect 462 140 463 141 
<< pdiffusion >>
rect 463 140 464 141 
<< pdiffusion >>
rect 464 140 465 141 
<< pdiffusion >>
rect 465 140 466 141 
<< pdiffusion >>
rect 466 140 467 141 
<< pdiffusion >>
rect 467 140 468 141 
<< m1 >>
rect 469 140 470 141 
<< m1 >>
rect 478 140 479 141 
<< pdiffusion >>
rect 498 140 499 141 
<< pdiffusion >>
rect 499 140 500 141 
<< pdiffusion >>
rect 500 140 501 141 
<< pdiffusion >>
rect 501 140 502 141 
<< pdiffusion >>
rect 502 140 503 141 
<< pdiffusion >>
rect 503 140 504 141 
<< pdiffusion >>
rect 516 140 517 141 
<< pdiffusion >>
rect 517 140 518 141 
<< pdiffusion >>
rect 518 140 519 141 
<< pdiffusion >>
rect 519 140 520 141 
<< pdiffusion >>
rect 520 140 521 141 
<< pdiffusion >>
rect 521 140 522 141 
<< pdiffusion >>
rect 12 141 13 142 
<< pdiffusion >>
rect 13 141 14 142 
<< pdiffusion >>
rect 14 141 15 142 
<< pdiffusion >>
rect 15 141 16 142 
<< pdiffusion >>
rect 16 141 17 142 
<< pdiffusion >>
rect 17 141 18 142 
<< pdiffusion >>
rect 30 141 31 142 
<< pdiffusion >>
rect 31 141 32 142 
<< pdiffusion >>
rect 32 141 33 142 
<< pdiffusion >>
rect 33 141 34 142 
<< pdiffusion >>
rect 34 141 35 142 
<< pdiffusion >>
rect 35 141 36 142 
<< m1 >>
rect 37 141 38 142 
<< m1 >>
rect 46 141 47 142 
<< pdiffusion >>
rect 48 141 49 142 
<< pdiffusion >>
rect 49 141 50 142 
<< pdiffusion >>
rect 50 141 51 142 
<< pdiffusion >>
rect 51 141 52 142 
<< pdiffusion >>
rect 52 141 53 142 
<< pdiffusion >>
rect 53 141 54 142 
<< m1 >>
rect 64 141 65 142 
<< pdiffusion >>
rect 66 141 67 142 
<< pdiffusion >>
rect 67 141 68 142 
<< pdiffusion >>
rect 68 141 69 142 
<< pdiffusion >>
rect 69 141 70 142 
<< pdiffusion >>
rect 70 141 71 142 
<< pdiffusion >>
rect 71 141 72 142 
<< m1 >>
rect 88 141 89 142 
<< m2 >>
rect 97 141 98 142 
<< m1 >>
rect 98 141 99 142 
<< m1 >>
rect 100 141 101 142 
<< pdiffusion >>
rect 102 141 103 142 
<< pdiffusion >>
rect 103 141 104 142 
<< pdiffusion >>
rect 104 141 105 142 
<< pdiffusion >>
rect 105 141 106 142 
<< pdiffusion >>
rect 106 141 107 142 
<< pdiffusion >>
rect 107 141 108 142 
<< m1 >>
rect 109 141 110 142 
<< m1 >>
rect 114 141 115 142 
<< m1 >>
rect 118 141 119 142 
<< m2 >>
rect 118 141 119 142 
<< pdiffusion >>
rect 120 141 121 142 
<< pdiffusion >>
rect 121 141 122 142 
<< pdiffusion >>
rect 122 141 123 142 
<< pdiffusion >>
rect 123 141 124 142 
<< pdiffusion >>
rect 124 141 125 142 
<< pdiffusion >>
rect 125 141 126 142 
<< m1 >>
rect 127 141 128 142 
<< m1 >>
rect 129 141 130 142 
<< m1 >>
rect 131 141 132 142 
<< m1 >>
rect 133 141 134 142 
<< m1 >>
rect 136 141 137 142 
<< pdiffusion >>
rect 138 141 139 142 
<< pdiffusion >>
rect 139 141 140 142 
<< pdiffusion >>
rect 140 141 141 142 
<< pdiffusion >>
rect 141 141 142 142 
<< pdiffusion >>
rect 142 141 143 142 
<< pdiffusion >>
rect 143 141 144 142 
<< m1 >>
rect 145 141 146 142 
<< pdiffusion >>
rect 156 141 157 142 
<< pdiffusion >>
rect 157 141 158 142 
<< pdiffusion >>
rect 158 141 159 142 
<< pdiffusion >>
rect 159 141 160 142 
<< pdiffusion >>
rect 160 141 161 142 
<< pdiffusion >>
rect 161 141 162 142 
<< m1 >>
rect 163 141 164 142 
<< pdiffusion >>
rect 174 141 175 142 
<< pdiffusion >>
rect 175 141 176 142 
<< pdiffusion >>
rect 176 141 177 142 
<< pdiffusion >>
rect 177 141 178 142 
<< pdiffusion >>
rect 178 141 179 142 
<< pdiffusion >>
rect 179 141 180 142 
<< pdiffusion >>
rect 192 141 193 142 
<< pdiffusion >>
rect 193 141 194 142 
<< pdiffusion >>
rect 194 141 195 142 
<< pdiffusion >>
rect 195 141 196 142 
<< pdiffusion >>
rect 196 141 197 142 
<< pdiffusion >>
rect 197 141 198 142 
<< m1 >>
rect 199 141 200 142 
<< pdiffusion >>
rect 210 141 211 142 
<< pdiffusion >>
rect 211 141 212 142 
<< pdiffusion >>
rect 212 141 213 142 
<< pdiffusion >>
rect 213 141 214 142 
<< pdiffusion >>
rect 214 141 215 142 
<< pdiffusion >>
rect 215 141 216 142 
<< m1 >>
rect 217 141 218 142 
<< m2 >>
rect 217 141 218 142 
<< m1 >>
rect 226 141 227 142 
<< pdiffusion >>
rect 228 141 229 142 
<< pdiffusion >>
rect 229 141 230 142 
<< pdiffusion >>
rect 230 141 231 142 
<< pdiffusion >>
rect 231 141 232 142 
<< pdiffusion >>
rect 232 141 233 142 
<< pdiffusion >>
rect 233 141 234 142 
<< m1 >>
rect 235 141 236 142 
<< m1 >>
rect 244 141 245 142 
<< pdiffusion >>
rect 246 141 247 142 
<< pdiffusion >>
rect 247 141 248 142 
<< pdiffusion >>
rect 248 141 249 142 
<< pdiffusion >>
rect 249 141 250 142 
<< pdiffusion >>
rect 250 141 251 142 
<< pdiffusion >>
rect 251 141 252 142 
<< pdiffusion >>
rect 264 141 265 142 
<< pdiffusion >>
rect 265 141 266 142 
<< pdiffusion >>
rect 266 141 267 142 
<< pdiffusion >>
rect 267 141 268 142 
<< pdiffusion >>
rect 268 141 269 142 
<< pdiffusion >>
rect 269 141 270 142 
<< m1 >>
rect 278 141 279 142 
<< m1 >>
rect 280 141 281 142 
<< m2 >>
rect 280 141 281 142 
<< pdiffusion >>
rect 282 141 283 142 
<< pdiffusion >>
rect 283 141 284 142 
<< pdiffusion >>
rect 284 141 285 142 
<< pdiffusion >>
rect 285 141 286 142 
<< pdiffusion >>
rect 286 141 287 142 
<< pdiffusion >>
rect 287 141 288 142 
<< pdiffusion >>
rect 300 141 301 142 
<< pdiffusion >>
rect 301 141 302 142 
<< pdiffusion >>
rect 302 141 303 142 
<< pdiffusion >>
rect 303 141 304 142 
<< pdiffusion >>
rect 304 141 305 142 
<< pdiffusion >>
rect 305 141 306 142 
<< m1 >>
rect 334 141 335 142 
<< m1 >>
rect 343 141 344 142 
<< pdiffusion >>
rect 354 141 355 142 
<< pdiffusion >>
rect 355 141 356 142 
<< pdiffusion >>
rect 356 141 357 142 
<< pdiffusion >>
rect 357 141 358 142 
<< pdiffusion >>
rect 358 141 359 142 
<< pdiffusion >>
rect 359 141 360 142 
<< m1 >>
rect 361 141 362 142 
<< m1 >>
rect 366 141 367 142 
<< m1 >>
rect 370 141 371 142 
<< pdiffusion >>
rect 372 141 373 142 
<< pdiffusion >>
rect 373 141 374 142 
<< pdiffusion >>
rect 374 141 375 142 
<< pdiffusion >>
rect 375 141 376 142 
<< pdiffusion >>
rect 376 141 377 142 
<< pdiffusion >>
rect 377 141 378 142 
<< m1 >>
rect 379 141 380 142 
<< m2 >>
rect 379 141 380 142 
<< pdiffusion >>
rect 390 141 391 142 
<< pdiffusion >>
rect 391 141 392 142 
<< pdiffusion >>
rect 392 141 393 142 
<< pdiffusion >>
rect 393 141 394 142 
<< pdiffusion >>
rect 394 141 395 142 
<< pdiffusion >>
rect 395 141 396 142 
<< pdiffusion >>
rect 408 141 409 142 
<< pdiffusion >>
rect 409 141 410 142 
<< pdiffusion >>
rect 410 141 411 142 
<< pdiffusion >>
rect 411 141 412 142 
<< pdiffusion >>
rect 412 141 413 142 
<< pdiffusion >>
rect 413 141 414 142 
<< m1 >>
rect 415 141 416 142 
<< m1 >>
rect 419 141 420 142 
<< m2 >>
rect 420 141 421 142 
<< pdiffusion >>
rect 426 141 427 142 
<< pdiffusion >>
rect 427 141 428 142 
<< pdiffusion >>
rect 428 141 429 142 
<< pdiffusion >>
rect 429 141 430 142 
<< pdiffusion >>
rect 430 141 431 142 
<< pdiffusion >>
rect 431 141 432 142 
<< m1 >>
rect 442 141 443 142 
<< pdiffusion >>
rect 444 141 445 142 
<< pdiffusion >>
rect 445 141 446 142 
<< pdiffusion >>
rect 446 141 447 142 
<< pdiffusion >>
rect 447 141 448 142 
<< pdiffusion >>
rect 448 141 449 142 
<< pdiffusion >>
rect 449 141 450 142 
<< m1 >>
rect 456 141 457 142 
<< pdiffusion >>
rect 462 141 463 142 
<< pdiffusion >>
rect 463 141 464 142 
<< pdiffusion >>
rect 464 141 465 142 
<< pdiffusion >>
rect 465 141 466 142 
<< pdiffusion >>
rect 466 141 467 142 
<< pdiffusion >>
rect 467 141 468 142 
<< m1 >>
rect 469 141 470 142 
<< m1 >>
rect 478 141 479 142 
<< pdiffusion >>
rect 498 141 499 142 
<< pdiffusion >>
rect 499 141 500 142 
<< pdiffusion >>
rect 500 141 501 142 
<< pdiffusion >>
rect 501 141 502 142 
<< pdiffusion >>
rect 502 141 503 142 
<< pdiffusion >>
rect 503 141 504 142 
<< pdiffusion >>
rect 516 141 517 142 
<< pdiffusion >>
rect 517 141 518 142 
<< pdiffusion >>
rect 518 141 519 142 
<< pdiffusion >>
rect 519 141 520 142 
<< pdiffusion >>
rect 520 141 521 142 
<< pdiffusion >>
rect 521 141 522 142 
<< pdiffusion >>
rect 12 142 13 143 
<< pdiffusion >>
rect 13 142 14 143 
<< pdiffusion >>
rect 14 142 15 143 
<< pdiffusion >>
rect 15 142 16 143 
<< pdiffusion >>
rect 16 142 17 143 
<< pdiffusion >>
rect 17 142 18 143 
<< pdiffusion >>
rect 30 142 31 143 
<< pdiffusion >>
rect 31 142 32 143 
<< pdiffusion >>
rect 32 142 33 143 
<< pdiffusion >>
rect 33 142 34 143 
<< pdiffusion >>
rect 34 142 35 143 
<< pdiffusion >>
rect 35 142 36 143 
<< m1 >>
rect 37 142 38 143 
<< m1 >>
rect 46 142 47 143 
<< pdiffusion >>
rect 48 142 49 143 
<< pdiffusion >>
rect 49 142 50 143 
<< pdiffusion >>
rect 50 142 51 143 
<< pdiffusion >>
rect 51 142 52 143 
<< pdiffusion >>
rect 52 142 53 143 
<< pdiffusion >>
rect 53 142 54 143 
<< m1 >>
rect 64 142 65 143 
<< pdiffusion >>
rect 66 142 67 143 
<< pdiffusion >>
rect 67 142 68 143 
<< pdiffusion >>
rect 68 142 69 143 
<< pdiffusion >>
rect 69 142 70 143 
<< pdiffusion >>
rect 70 142 71 143 
<< pdiffusion >>
rect 71 142 72 143 
<< m1 >>
rect 88 142 89 143 
<< m2 >>
rect 97 142 98 143 
<< m1 >>
rect 98 142 99 143 
<< m1 >>
rect 100 142 101 143 
<< pdiffusion >>
rect 102 142 103 143 
<< pdiffusion >>
rect 103 142 104 143 
<< pdiffusion >>
rect 104 142 105 143 
<< pdiffusion >>
rect 105 142 106 143 
<< pdiffusion >>
rect 106 142 107 143 
<< pdiffusion >>
rect 107 142 108 143 
<< m1 >>
rect 109 142 110 143 
<< m1 >>
rect 114 142 115 143 
<< m1 >>
rect 118 142 119 143 
<< m2 >>
rect 118 142 119 143 
<< pdiffusion >>
rect 120 142 121 143 
<< pdiffusion >>
rect 121 142 122 143 
<< pdiffusion >>
rect 122 142 123 143 
<< pdiffusion >>
rect 123 142 124 143 
<< pdiffusion >>
rect 124 142 125 143 
<< pdiffusion >>
rect 125 142 126 143 
<< m1 >>
rect 127 142 128 143 
<< m1 >>
rect 129 142 130 143 
<< m1 >>
rect 131 142 132 143 
<< m1 >>
rect 133 142 134 143 
<< m1 >>
rect 136 142 137 143 
<< pdiffusion >>
rect 138 142 139 143 
<< pdiffusion >>
rect 139 142 140 143 
<< pdiffusion >>
rect 140 142 141 143 
<< pdiffusion >>
rect 141 142 142 143 
<< pdiffusion >>
rect 142 142 143 143 
<< pdiffusion >>
rect 143 142 144 143 
<< m1 >>
rect 145 142 146 143 
<< pdiffusion >>
rect 156 142 157 143 
<< pdiffusion >>
rect 157 142 158 143 
<< pdiffusion >>
rect 158 142 159 143 
<< pdiffusion >>
rect 159 142 160 143 
<< pdiffusion >>
rect 160 142 161 143 
<< pdiffusion >>
rect 161 142 162 143 
<< m1 >>
rect 163 142 164 143 
<< pdiffusion >>
rect 174 142 175 143 
<< pdiffusion >>
rect 175 142 176 143 
<< pdiffusion >>
rect 176 142 177 143 
<< pdiffusion >>
rect 177 142 178 143 
<< pdiffusion >>
rect 178 142 179 143 
<< pdiffusion >>
rect 179 142 180 143 
<< pdiffusion >>
rect 192 142 193 143 
<< pdiffusion >>
rect 193 142 194 143 
<< pdiffusion >>
rect 194 142 195 143 
<< pdiffusion >>
rect 195 142 196 143 
<< pdiffusion >>
rect 196 142 197 143 
<< pdiffusion >>
rect 197 142 198 143 
<< m1 >>
rect 199 142 200 143 
<< pdiffusion >>
rect 210 142 211 143 
<< pdiffusion >>
rect 211 142 212 143 
<< pdiffusion >>
rect 212 142 213 143 
<< pdiffusion >>
rect 213 142 214 143 
<< pdiffusion >>
rect 214 142 215 143 
<< pdiffusion >>
rect 215 142 216 143 
<< m1 >>
rect 217 142 218 143 
<< m2 >>
rect 217 142 218 143 
<< m1 >>
rect 226 142 227 143 
<< pdiffusion >>
rect 228 142 229 143 
<< pdiffusion >>
rect 229 142 230 143 
<< pdiffusion >>
rect 230 142 231 143 
<< pdiffusion >>
rect 231 142 232 143 
<< pdiffusion >>
rect 232 142 233 143 
<< pdiffusion >>
rect 233 142 234 143 
<< m1 >>
rect 235 142 236 143 
<< m1 >>
rect 244 142 245 143 
<< pdiffusion >>
rect 246 142 247 143 
<< pdiffusion >>
rect 247 142 248 143 
<< pdiffusion >>
rect 248 142 249 143 
<< pdiffusion >>
rect 249 142 250 143 
<< pdiffusion >>
rect 250 142 251 143 
<< pdiffusion >>
rect 251 142 252 143 
<< pdiffusion >>
rect 264 142 265 143 
<< pdiffusion >>
rect 265 142 266 143 
<< pdiffusion >>
rect 266 142 267 143 
<< pdiffusion >>
rect 267 142 268 143 
<< pdiffusion >>
rect 268 142 269 143 
<< pdiffusion >>
rect 269 142 270 143 
<< m1 >>
rect 278 142 279 143 
<< m1 >>
rect 280 142 281 143 
<< m2 >>
rect 280 142 281 143 
<< pdiffusion >>
rect 282 142 283 143 
<< pdiffusion >>
rect 283 142 284 143 
<< pdiffusion >>
rect 284 142 285 143 
<< pdiffusion >>
rect 285 142 286 143 
<< pdiffusion >>
rect 286 142 287 143 
<< pdiffusion >>
rect 287 142 288 143 
<< pdiffusion >>
rect 300 142 301 143 
<< pdiffusion >>
rect 301 142 302 143 
<< pdiffusion >>
rect 302 142 303 143 
<< pdiffusion >>
rect 303 142 304 143 
<< pdiffusion >>
rect 304 142 305 143 
<< pdiffusion >>
rect 305 142 306 143 
<< m1 >>
rect 334 142 335 143 
<< m1 >>
rect 343 142 344 143 
<< pdiffusion >>
rect 354 142 355 143 
<< pdiffusion >>
rect 355 142 356 143 
<< pdiffusion >>
rect 356 142 357 143 
<< pdiffusion >>
rect 357 142 358 143 
<< pdiffusion >>
rect 358 142 359 143 
<< pdiffusion >>
rect 359 142 360 143 
<< m1 >>
rect 361 142 362 143 
<< m1 >>
rect 366 142 367 143 
<< m1 >>
rect 370 142 371 143 
<< pdiffusion >>
rect 372 142 373 143 
<< pdiffusion >>
rect 373 142 374 143 
<< pdiffusion >>
rect 374 142 375 143 
<< pdiffusion >>
rect 375 142 376 143 
<< pdiffusion >>
rect 376 142 377 143 
<< pdiffusion >>
rect 377 142 378 143 
<< m1 >>
rect 379 142 380 143 
<< m2 >>
rect 379 142 380 143 
<< pdiffusion >>
rect 390 142 391 143 
<< pdiffusion >>
rect 391 142 392 143 
<< pdiffusion >>
rect 392 142 393 143 
<< pdiffusion >>
rect 393 142 394 143 
<< pdiffusion >>
rect 394 142 395 143 
<< pdiffusion >>
rect 395 142 396 143 
<< pdiffusion >>
rect 408 142 409 143 
<< pdiffusion >>
rect 409 142 410 143 
<< pdiffusion >>
rect 410 142 411 143 
<< pdiffusion >>
rect 411 142 412 143 
<< pdiffusion >>
rect 412 142 413 143 
<< pdiffusion >>
rect 413 142 414 143 
<< m1 >>
rect 415 142 416 143 
<< m1 >>
rect 419 142 420 143 
<< m2 >>
rect 420 142 421 143 
<< pdiffusion >>
rect 426 142 427 143 
<< pdiffusion >>
rect 427 142 428 143 
<< pdiffusion >>
rect 428 142 429 143 
<< pdiffusion >>
rect 429 142 430 143 
<< pdiffusion >>
rect 430 142 431 143 
<< pdiffusion >>
rect 431 142 432 143 
<< m1 >>
rect 442 142 443 143 
<< pdiffusion >>
rect 444 142 445 143 
<< pdiffusion >>
rect 445 142 446 143 
<< pdiffusion >>
rect 446 142 447 143 
<< pdiffusion >>
rect 447 142 448 143 
<< pdiffusion >>
rect 448 142 449 143 
<< pdiffusion >>
rect 449 142 450 143 
<< m1 >>
rect 456 142 457 143 
<< pdiffusion >>
rect 462 142 463 143 
<< pdiffusion >>
rect 463 142 464 143 
<< pdiffusion >>
rect 464 142 465 143 
<< pdiffusion >>
rect 465 142 466 143 
<< pdiffusion >>
rect 466 142 467 143 
<< pdiffusion >>
rect 467 142 468 143 
<< m1 >>
rect 469 142 470 143 
<< m1 >>
rect 478 142 479 143 
<< pdiffusion >>
rect 498 142 499 143 
<< pdiffusion >>
rect 499 142 500 143 
<< pdiffusion >>
rect 500 142 501 143 
<< pdiffusion >>
rect 501 142 502 143 
<< pdiffusion >>
rect 502 142 503 143 
<< pdiffusion >>
rect 503 142 504 143 
<< pdiffusion >>
rect 516 142 517 143 
<< pdiffusion >>
rect 517 142 518 143 
<< pdiffusion >>
rect 518 142 519 143 
<< pdiffusion >>
rect 519 142 520 143 
<< pdiffusion >>
rect 520 142 521 143 
<< pdiffusion >>
rect 521 142 522 143 
<< pdiffusion >>
rect 12 143 13 144 
<< pdiffusion >>
rect 13 143 14 144 
<< pdiffusion >>
rect 14 143 15 144 
<< pdiffusion >>
rect 15 143 16 144 
<< pdiffusion >>
rect 16 143 17 144 
<< pdiffusion >>
rect 17 143 18 144 
<< pdiffusion >>
rect 30 143 31 144 
<< pdiffusion >>
rect 31 143 32 144 
<< pdiffusion >>
rect 32 143 33 144 
<< pdiffusion >>
rect 33 143 34 144 
<< m1 >>
rect 34 143 35 144 
<< pdiffusion >>
rect 34 143 35 144 
<< pdiffusion >>
rect 35 143 36 144 
<< m1 >>
rect 37 143 38 144 
<< m2 >>
rect 37 143 38 144 
<< m2c >>
rect 37 143 38 144 
<< m1 >>
rect 37 143 38 144 
<< m2 >>
rect 37 143 38 144 
<< m1 >>
rect 46 143 47 144 
<< pdiffusion >>
rect 48 143 49 144 
<< pdiffusion >>
rect 49 143 50 144 
<< pdiffusion >>
rect 50 143 51 144 
<< pdiffusion >>
rect 51 143 52 144 
<< pdiffusion >>
rect 52 143 53 144 
<< pdiffusion >>
rect 53 143 54 144 
<< m1 >>
rect 64 143 65 144 
<< pdiffusion >>
rect 66 143 67 144 
<< pdiffusion >>
rect 67 143 68 144 
<< pdiffusion >>
rect 68 143 69 144 
<< pdiffusion >>
rect 69 143 70 144 
<< m1 >>
rect 70 143 71 144 
<< pdiffusion >>
rect 70 143 71 144 
<< pdiffusion >>
rect 71 143 72 144 
<< m1 >>
rect 88 143 89 144 
<< m2 >>
rect 97 143 98 144 
<< m1 >>
rect 98 143 99 144 
<< m1 >>
rect 100 143 101 144 
<< pdiffusion >>
rect 102 143 103 144 
<< pdiffusion >>
rect 103 143 104 144 
<< pdiffusion >>
rect 104 143 105 144 
<< pdiffusion >>
rect 105 143 106 144 
<< pdiffusion >>
rect 106 143 107 144 
<< pdiffusion >>
rect 107 143 108 144 
<< m1 >>
rect 109 143 110 144 
<< m1 >>
rect 114 143 115 144 
<< m1 >>
rect 118 143 119 144 
<< m2 >>
rect 118 143 119 144 
<< pdiffusion >>
rect 120 143 121 144 
<< pdiffusion >>
rect 121 143 122 144 
<< pdiffusion >>
rect 122 143 123 144 
<< pdiffusion >>
rect 123 143 124 144 
<< m1 >>
rect 124 143 125 144 
<< pdiffusion >>
rect 124 143 125 144 
<< pdiffusion >>
rect 125 143 126 144 
<< m1 >>
rect 127 143 128 144 
<< m1 >>
rect 129 143 130 144 
<< m1 >>
rect 131 143 132 144 
<< m1 >>
rect 133 143 134 144 
<< m1 >>
rect 136 143 137 144 
<< pdiffusion >>
rect 138 143 139 144 
<< pdiffusion >>
rect 139 143 140 144 
<< pdiffusion >>
rect 140 143 141 144 
<< pdiffusion >>
rect 141 143 142 144 
<< m1 >>
rect 142 143 143 144 
<< pdiffusion >>
rect 142 143 143 144 
<< pdiffusion >>
rect 143 143 144 144 
<< m1 >>
rect 145 143 146 144 
<< pdiffusion >>
rect 156 143 157 144 
<< pdiffusion >>
rect 157 143 158 144 
<< pdiffusion >>
rect 158 143 159 144 
<< pdiffusion >>
rect 159 143 160 144 
<< pdiffusion >>
rect 160 143 161 144 
<< pdiffusion >>
rect 161 143 162 144 
<< m1 >>
rect 163 143 164 144 
<< pdiffusion >>
rect 174 143 175 144 
<< pdiffusion >>
rect 175 143 176 144 
<< pdiffusion >>
rect 176 143 177 144 
<< pdiffusion >>
rect 177 143 178 144 
<< pdiffusion >>
rect 178 143 179 144 
<< pdiffusion >>
rect 179 143 180 144 
<< pdiffusion >>
rect 192 143 193 144 
<< m1 >>
rect 193 143 194 144 
<< pdiffusion >>
rect 193 143 194 144 
<< pdiffusion >>
rect 194 143 195 144 
<< pdiffusion >>
rect 195 143 196 144 
<< pdiffusion >>
rect 196 143 197 144 
<< pdiffusion >>
rect 197 143 198 144 
<< m1 >>
rect 199 143 200 144 
<< pdiffusion >>
rect 210 143 211 144 
<< m1 >>
rect 211 143 212 144 
<< pdiffusion >>
rect 211 143 212 144 
<< pdiffusion >>
rect 212 143 213 144 
<< pdiffusion >>
rect 213 143 214 144 
<< pdiffusion >>
rect 214 143 215 144 
<< pdiffusion >>
rect 215 143 216 144 
<< m1 >>
rect 217 143 218 144 
<< m2 >>
rect 217 143 218 144 
<< m1 >>
rect 226 143 227 144 
<< pdiffusion >>
rect 228 143 229 144 
<< pdiffusion >>
rect 229 143 230 144 
<< pdiffusion >>
rect 230 143 231 144 
<< pdiffusion >>
rect 231 143 232 144 
<< m1 >>
rect 232 143 233 144 
<< pdiffusion >>
rect 232 143 233 144 
<< pdiffusion >>
rect 233 143 234 144 
<< m1 >>
rect 235 143 236 144 
<< m1 >>
rect 244 143 245 144 
<< pdiffusion >>
rect 246 143 247 144 
<< pdiffusion >>
rect 247 143 248 144 
<< pdiffusion >>
rect 248 143 249 144 
<< pdiffusion >>
rect 249 143 250 144 
<< pdiffusion >>
rect 250 143 251 144 
<< pdiffusion >>
rect 251 143 252 144 
<< pdiffusion >>
rect 264 143 265 144 
<< pdiffusion >>
rect 265 143 266 144 
<< pdiffusion >>
rect 266 143 267 144 
<< pdiffusion >>
rect 267 143 268 144 
<< pdiffusion >>
rect 268 143 269 144 
<< pdiffusion >>
rect 269 143 270 144 
<< m1 >>
rect 278 143 279 144 
<< m1 >>
rect 280 143 281 144 
<< m2 >>
rect 280 143 281 144 
<< pdiffusion >>
rect 282 143 283 144 
<< pdiffusion >>
rect 283 143 284 144 
<< pdiffusion >>
rect 284 143 285 144 
<< pdiffusion >>
rect 285 143 286 144 
<< pdiffusion >>
rect 286 143 287 144 
<< pdiffusion >>
rect 287 143 288 144 
<< pdiffusion >>
rect 300 143 301 144 
<< pdiffusion >>
rect 301 143 302 144 
<< pdiffusion >>
rect 302 143 303 144 
<< pdiffusion >>
rect 303 143 304 144 
<< pdiffusion >>
rect 304 143 305 144 
<< pdiffusion >>
rect 305 143 306 144 
<< m1 >>
rect 334 143 335 144 
<< m1 >>
rect 343 143 344 144 
<< pdiffusion >>
rect 354 143 355 144 
<< pdiffusion >>
rect 355 143 356 144 
<< pdiffusion >>
rect 356 143 357 144 
<< pdiffusion >>
rect 357 143 358 144 
<< pdiffusion >>
rect 358 143 359 144 
<< pdiffusion >>
rect 359 143 360 144 
<< m1 >>
rect 361 143 362 144 
<< m1 >>
rect 366 143 367 144 
<< m1 >>
rect 370 143 371 144 
<< pdiffusion >>
rect 372 143 373 144 
<< pdiffusion >>
rect 373 143 374 144 
<< pdiffusion >>
rect 374 143 375 144 
<< pdiffusion >>
rect 375 143 376 144 
<< pdiffusion >>
rect 376 143 377 144 
<< pdiffusion >>
rect 377 143 378 144 
<< m1 >>
rect 379 143 380 144 
<< m2 >>
rect 379 143 380 144 
<< pdiffusion >>
rect 390 143 391 144 
<< pdiffusion >>
rect 391 143 392 144 
<< pdiffusion >>
rect 392 143 393 144 
<< pdiffusion >>
rect 393 143 394 144 
<< pdiffusion >>
rect 394 143 395 144 
<< pdiffusion >>
rect 395 143 396 144 
<< pdiffusion >>
rect 408 143 409 144 
<< pdiffusion >>
rect 409 143 410 144 
<< pdiffusion >>
rect 410 143 411 144 
<< pdiffusion >>
rect 411 143 412 144 
<< m1 >>
rect 412 143 413 144 
<< pdiffusion >>
rect 412 143 413 144 
<< pdiffusion >>
rect 413 143 414 144 
<< m1 >>
rect 415 143 416 144 
<< m1 >>
rect 419 143 420 144 
<< m2 >>
rect 420 143 421 144 
<< pdiffusion >>
rect 426 143 427 144 
<< m1 >>
rect 427 143 428 144 
<< pdiffusion >>
rect 427 143 428 144 
<< pdiffusion >>
rect 428 143 429 144 
<< pdiffusion >>
rect 429 143 430 144 
<< pdiffusion >>
rect 430 143 431 144 
<< pdiffusion >>
rect 431 143 432 144 
<< m1 >>
rect 442 143 443 144 
<< pdiffusion >>
rect 444 143 445 144 
<< pdiffusion >>
rect 445 143 446 144 
<< pdiffusion >>
rect 446 143 447 144 
<< pdiffusion >>
rect 447 143 448 144 
<< pdiffusion >>
rect 448 143 449 144 
<< pdiffusion >>
rect 449 143 450 144 
<< m1 >>
rect 456 143 457 144 
<< pdiffusion >>
rect 462 143 463 144 
<< pdiffusion >>
rect 463 143 464 144 
<< pdiffusion >>
rect 464 143 465 144 
<< pdiffusion >>
rect 465 143 466 144 
<< pdiffusion >>
rect 466 143 467 144 
<< pdiffusion >>
rect 467 143 468 144 
<< m1 >>
rect 469 143 470 144 
<< m1 >>
rect 478 143 479 144 
<< pdiffusion >>
rect 498 143 499 144 
<< pdiffusion >>
rect 499 143 500 144 
<< pdiffusion >>
rect 500 143 501 144 
<< pdiffusion >>
rect 501 143 502 144 
<< pdiffusion >>
rect 502 143 503 144 
<< pdiffusion >>
rect 503 143 504 144 
<< pdiffusion >>
rect 516 143 517 144 
<< pdiffusion >>
rect 517 143 518 144 
<< pdiffusion >>
rect 518 143 519 144 
<< pdiffusion >>
rect 519 143 520 144 
<< pdiffusion >>
rect 520 143 521 144 
<< pdiffusion >>
rect 521 143 522 144 
<< m1 >>
rect 34 144 35 145 
<< m2 >>
rect 37 144 38 145 
<< m1 >>
rect 46 144 47 145 
<< m1 >>
rect 64 144 65 145 
<< m1 >>
rect 70 144 71 145 
<< m1 >>
rect 88 144 89 145 
<< m2 >>
rect 97 144 98 145 
<< m1 >>
rect 98 144 99 145 
<< m1 >>
rect 100 144 101 145 
<< m1 >>
rect 109 144 110 145 
<< m1 >>
rect 114 144 115 145 
<< m1 >>
rect 118 144 119 145 
<< m2 >>
rect 118 144 119 145 
<< m1 >>
rect 124 144 125 145 
<< m1 >>
rect 127 144 128 145 
<< m1 >>
rect 129 144 130 145 
<< m1 >>
rect 131 144 132 145 
<< m1 >>
rect 133 144 134 145 
<< m1 >>
rect 136 144 137 145 
<< m1 >>
rect 142 144 143 145 
<< m1 >>
rect 145 144 146 145 
<< m1 >>
rect 163 144 164 145 
<< m1 >>
rect 193 144 194 145 
<< m1 >>
rect 199 144 200 145 
<< m1 >>
rect 211 144 212 145 
<< m1 >>
rect 217 144 218 145 
<< m2 >>
rect 217 144 218 145 
<< m1 >>
rect 226 144 227 145 
<< m1 >>
rect 232 144 233 145 
<< m1 >>
rect 235 144 236 145 
<< m1 >>
rect 244 144 245 145 
<< m1 >>
rect 278 144 279 145 
<< m1 >>
rect 280 144 281 145 
<< m2 >>
rect 280 144 281 145 
<< m1 >>
rect 334 144 335 145 
<< m1 >>
rect 343 144 344 145 
<< m1 >>
rect 361 144 362 145 
<< m1 >>
rect 366 144 367 145 
<< m1 >>
rect 370 144 371 145 
<< m1 >>
rect 379 144 380 145 
<< m2 >>
rect 379 144 380 145 
<< m1 >>
rect 412 144 413 145 
<< m1 >>
rect 415 144 416 145 
<< m1 >>
rect 419 144 420 145 
<< m2 >>
rect 420 144 421 145 
<< m1 >>
rect 427 144 428 145 
<< m1 >>
rect 442 144 443 145 
<< m1 >>
rect 456 144 457 145 
<< m1 >>
rect 469 144 470 145 
<< m1 >>
rect 478 144 479 145 
<< m1 >>
rect 34 145 35 146 
<< m1 >>
rect 35 145 36 146 
<< m1 >>
rect 36 145 37 146 
<< m1 >>
rect 37 145 38 146 
<< m2 >>
rect 37 145 38 146 
<< m1 >>
rect 38 145 39 146 
<< m1 >>
rect 39 145 40 146 
<< m1 >>
rect 40 145 41 146 
<< m1 >>
rect 41 145 42 146 
<< m1 >>
rect 42 145 43 146 
<< m1 >>
rect 43 145 44 146 
<< m1 >>
rect 44 145 45 146 
<< m1 >>
rect 45 145 46 146 
<< m1 >>
rect 46 145 47 146 
<< m1 >>
rect 64 145 65 146 
<< m1 >>
rect 70 145 71 146 
<< m1 >>
rect 71 145 72 146 
<< m1 >>
rect 72 145 73 146 
<< m1 >>
rect 73 145 74 146 
<< m1 >>
rect 74 145 75 146 
<< m1 >>
rect 75 145 76 146 
<< m1 >>
rect 76 145 77 146 
<< m1 >>
rect 77 145 78 146 
<< m1 >>
rect 78 145 79 146 
<< m1 >>
rect 79 145 80 146 
<< m1 >>
rect 80 145 81 146 
<< m1 >>
rect 81 145 82 146 
<< m1 >>
rect 82 145 83 146 
<< m1 >>
rect 83 145 84 146 
<< m1 >>
rect 84 145 85 146 
<< m1 >>
rect 85 145 86 146 
<< m1 >>
rect 86 145 87 146 
<< m1 >>
rect 87 145 88 146 
<< m1 >>
rect 88 145 89 146 
<< m2 >>
rect 97 145 98 146 
<< m1 >>
rect 98 145 99 146 
<< m1 >>
rect 100 145 101 146 
<< m1 >>
rect 109 145 110 146 
<< m1 >>
rect 114 145 115 146 
<< m1 >>
rect 118 145 119 146 
<< m2 >>
rect 118 145 119 146 
<< m1 >>
rect 124 145 125 146 
<< m1 >>
rect 125 145 126 146 
<< m2 >>
rect 125 145 126 146 
<< m2c >>
rect 125 145 126 146 
<< m1 >>
rect 125 145 126 146 
<< m2 >>
rect 125 145 126 146 
<< m2 >>
rect 126 145 127 146 
<< m1 >>
rect 127 145 128 146 
<< m2 >>
rect 127 145 128 146 
<< m2 >>
rect 128 145 129 146 
<< m1 >>
rect 129 145 130 146 
<< m2 >>
rect 129 145 130 146 
<< m2 >>
rect 130 145 131 146 
<< m1 >>
rect 131 145 132 146 
<< m2 >>
rect 131 145 132 146 
<< m2 >>
rect 132 145 133 146 
<< m1 >>
rect 133 145 134 146 
<< m2 >>
rect 133 145 134 146 
<< m2c >>
rect 133 145 134 146 
<< m1 >>
rect 133 145 134 146 
<< m2 >>
rect 133 145 134 146 
<< m1 >>
rect 136 145 137 146 
<< m1 >>
rect 142 145 143 146 
<< m1 >>
rect 143 145 144 146 
<< m2 >>
rect 143 145 144 146 
<< m2c >>
rect 143 145 144 146 
<< m1 >>
rect 143 145 144 146 
<< m2 >>
rect 143 145 144 146 
<< m2 >>
rect 144 145 145 146 
<< m1 >>
rect 145 145 146 146 
<< m2 >>
rect 145 145 146 146 
<< m2 >>
rect 146 145 147 146 
<< m1 >>
rect 147 145 148 146 
<< m2 >>
rect 147 145 148 146 
<< m2c >>
rect 147 145 148 146 
<< m1 >>
rect 147 145 148 146 
<< m2 >>
rect 147 145 148 146 
<< m1 >>
rect 163 145 164 146 
<< m1 >>
rect 193 145 194 146 
<< m1 >>
rect 199 145 200 146 
<< m1 >>
rect 211 145 212 146 
<< m1 >>
rect 217 145 218 146 
<< m2 >>
rect 217 145 218 146 
<< m1 >>
rect 226 145 227 146 
<< m1 >>
rect 232 145 233 146 
<< m1 >>
rect 235 145 236 146 
<< m1 >>
rect 244 145 245 146 
<< m1 >>
rect 278 145 279 146 
<< m1 >>
rect 280 145 281 146 
<< m2 >>
rect 280 145 281 146 
<< m1 >>
rect 334 145 335 146 
<< m1 >>
rect 343 145 344 146 
<< m1 >>
rect 361 145 362 146 
<< m1 >>
rect 366 145 367 146 
<< m1 >>
rect 370 145 371 146 
<< m1 >>
rect 379 145 380 146 
<< m2 >>
rect 379 145 380 146 
<< m1 >>
rect 412 145 413 146 
<< m1 >>
rect 413 145 414 146 
<< m2 >>
rect 413 145 414 146 
<< m2c >>
rect 413 145 414 146 
<< m1 >>
rect 413 145 414 146 
<< m2 >>
rect 413 145 414 146 
<< m2 >>
rect 414 145 415 146 
<< m1 >>
rect 415 145 416 146 
<< m2 >>
rect 415 145 416 146 
<< m2 >>
rect 416 145 417 146 
<< m1 >>
rect 417 145 418 146 
<< m2 >>
rect 417 145 418 146 
<< m2c >>
rect 417 145 418 146 
<< m1 >>
rect 417 145 418 146 
<< m2 >>
rect 417 145 418 146 
<< m1 >>
rect 419 145 420 146 
<< m2 >>
rect 420 145 421 146 
<< m1 >>
rect 427 145 428 146 
<< m1 >>
rect 442 145 443 146 
<< m1 >>
rect 456 145 457 146 
<< m1 >>
rect 469 145 470 146 
<< m1 >>
rect 478 145 479 146 
<< m2 >>
rect 37 146 38 147 
<< m1 >>
rect 64 146 65 147 
<< m2 >>
rect 97 146 98 147 
<< m1 >>
rect 98 146 99 147 
<< m1 >>
rect 100 146 101 147 
<< m1 >>
rect 109 146 110 147 
<< m1 >>
rect 114 146 115 147 
<< m1 >>
rect 118 146 119 147 
<< m2 >>
rect 118 146 119 147 
<< m1 >>
rect 127 146 128 147 
<< m1 >>
rect 129 146 130 147 
<< m1 >>
rect 131 146 132 147 
<< m1 >>
rect 136 146 137 147 
<< m1 >>
rect 145 146 146 147 
<< m1 >>
rect 147 146 148 147 
<< m1 >>
rect 158 146 159 147 
<< m1 >>
rect 159 146 160 147 
<< m1 >>
rect 160 146 161 147 
<< m1 >>
rect 161 146 162 147 
<< m2 >>
rect 161 146 162 147 
<< m2c >>
rect 161 146 162 147 
<< m1 >>
rect 161 146 162 147 
<< m2 >>
rect 161 146 162 147 
<< m2 >>
rect 162 146 163 147 
<< m1 >>
rect 163 146 164 147 
<< m2 >>
rect 163 146 164 147 
<< m2 >>
rect 164 146 165 147 
<< m1 >>
rect 165 146 166 147 
<< m2 >>
rect 165 146 166 147 
<< m2c >>
rect 165 146 166 147 
<< m1 >>
rect 165 146 166 147 
<< m2 >>
rect 165 146 166 147 
<< m1 >>
rect 193 146 194 147 
<< m1 >>
rect 194 146 195 147 
<< m1 >>
rect 195 146 196 147 
<< m1 >>
rect 196 146 197 147 
<< m1 >>
rect 197 146 198 147 
<< m1 >>
rect 198 146 199 147 
<< m1 >>
rect 199 146 200 147 
<< m1 >>
rect 211 146 212 147 
<< m1 >>
rect 217 146 218 147 
<< m2 >>
rect 217 146 218 147 
<< m1 >>
rect 226 146 227 147 
<< m2 >>
rect 226 146 227 147 
<< m2c >>
rect 226 146 227 147 
<< m1 >>
rect 226 146 227 147 
<< m2 >>
rect 226 146 227 147 
<< m1 >>
rect 232 146 233 147 
<< m1 >>
rect 235 146 236 147 
<< m1 >>
rect 244 146 245 147 
<< m1 >>
rect 278 146 279 147 
<< m1 >>
rect 280 146 281 147 
<< m2 >>
rect 280 146 281 147 
<< m1 >>
rect 334 146 335 147 
<< m1 >>
rect 343 146 344 147 
<< m1 >>
rect 361 146 362 147 
<< m1 >>
rect 366 146 367 147 
<< m1 >>
rect 370 146 371 147 
<< m1 >>
rect 379 146 380 147 
<< m2 >>
rect 379 146 380 147 
<< m1 >>
rect 415 146 416 147 
<< m1 >>
rect 417 146 418 147 
<< m1 >>
rect 419 146 420 147 
<< m2 >>
rect 420 146 421 147 
<< m1 >>
rect 427 146 428 147 
<< m1 >>
rect 428 146 429 147 
<< m1 >>
rect 429 146 430 147 
<< m1 >>
rect 430 146 431 147 
<< m1 >>
rect 431 146 432 147 
<< m1 >>
rect 432 146 433 147 
<< m1 >>
rect 433 146 434 147 
<< m1 >>
rect 442 146 443 147 
<< m1 >>
rect 456 146 457 147 
<< m1 >>
rect 469 146 470 147 
<< m1 >>
rect 478 146 479 147 
<< m2 >>
rect 478 146 479 147 
<< m2c >>
rect 478 146 479 147 
<< m1 >>
rect 478 146 479 147 
<< m2 >>
rect 478 146 479 147 
<< m1 >>
rect 37 147 38 148 
<< m2 >>
rect 37 147 38 148 
<< m2c >>
rect 37 147 38 148 
<< m1 >>
rect 37 147 38 148 
<< m2 >>
rect 37 147 38 148 
<< m1 >>
rect 64 147 65 148 
<< m2 >>
rect 97 147 98 148 
<< m1 >>
rect 98 147 99 148 
<< m1 >>
rect 100 147 101 148 
<< m1 >>
rect 109 147 110 148 
<< m1 >>
rect 114 147 115 148 
<< m1 >>
rect 118 147 119 148 
<< m2 >>
rect 118 147 119 148 
<< m1 >>
rect 127 147 128 148 
<< m2 >>
rect 127 147 128 148 
<< m2 >>
rect 128 147 129 148 
<< m1 >>
rect 129 147 130 148 
<< m2 >>
rect 129 147 130 148 
<< m2 >>
rect 130 147 131 148 
<< m1 >>
rect 131 147 132 148 
<< m2 >>
rect 131 147 132 148 
<< m2 >>
rect 132 147 133 148 
<< m1 >>
rect 133 147 134 148 
<< m2 >>
rect 133 147 134 148 
<< m2c >>
rect 133 147 134 148 
<< m1 >>
rect 133 147 134 148 
<< m2 >>
rect 133 147 134 148 
<< m1 >>
rect 134 147 135 148 
<< m1 >>
rect 135 147 136 148 
<< m1 >>
rect 136 147 137 148 
<< m1 >>
rect 145 147 146 148 
<< m1 >>
rect 147 147 148 148 
<< m1 >>
rect 158 147 159 148 
<< m1 >>
rect 163 147 164 148 
<< m1 >>
rect 165 147 166 148 
<< m1 >>
rect 211 147 212 148 
<< m1 >>
rect 217 147 218 148 
<< m2 >>
rect 217 147 218 148 
<< m2 >>
rect 218 147 219 148 
<< m2 >>
rect 219 147 220 148 
<< m2 >>
rect 220 147 221 148 
<< m2 >>
rect 221 147 222 148 
<< m2 >>
rect 226 147 227 148 
<< m1 >>
rect 232 147 233 148 
<< m1 >>
rect 235 147 236 148 
<< m1 >>
rect 244 147 245 148 
<< m1 >>
rect 278 147 279 148 
<< m1 >>
rect 280 147 281 148 
<< m2 >>
rect 280 147 281 148 
<< m1 >>
rect 334 147 335 148 
<< m1 >>
rect 343 147 344 148 
<< m1 >>
rect 361 147 362 148 
<< m1 >>
rect 366 147 367 148 
<< m1 >>
rect 370 147 371 148 
<< m1 >>
rect 379 147 380 148 
<< m2 >>
rect 379 147 380 148 
<< m1 >>
rect 412 147 413 148 
<< m1 >>
rect 413 147 414 148 
<< m2 >>
rect 413 147 414 148 
<< m2c >>
rect 413 147 414 148 
<< m1 >>
rect 413 147 414 148 
<< m2 >>
rect 413 147 414 148 
<< m2 >>
rect 414 147 415 148 
<< m1 >>
rect 415 147 416 148 
<< m2 >>
rect 415 147 416 148 
<< m2 >>
rect 416 147 417 148 
<< m1 >>
rect 417 147 418 148 
<< m2 >>
rect 417 147 418 148 
<< m2 >>
rect 418 147 419 148 
<< m1 >>
rect 419 147 420 148 
<< m2 >>
rect 419 147 420 148 
<< m2 >>
rect 420 147 421 148 
<< m1 >>
rect 433 147 434 148 
<< m1 >>
rect 442 147 443 148 
<< m1 >>
rect 456 147 457 148 
<< m1 >>
rect 469 147 470 148 
<< m2 >>
rect 478 147 479 148 
<< m1 >>
rect 37 148 38 149 
<< m1 >>
rect 64 148 65 149 
<< m2 >>
rect 97 148 98 149 
<< m1 >>
rect 98 148 99 149 
<< m1 >>
rect 100 148 101 149 
<< m1 >>
rect 109 148 110 149 
<< m1 >>
rect 114 148 115 149 
<< m1 >>
rect 118 148 119 149 
<< m2 >>
rect 118 148 119 149 
<< m1 >>
rect 127 148 128 149 
<< m2 >>
rect 127 148 128 149 
<< m1 >>
rect 129 148 130 149 
<< m1 >>
rect 131 148 132 149 
<< m1 >>
rect 145 148 146 149 
<< m2 >>
rect 145 148 146 149 
<< m2c >>
rect 145 148 146 149 
<< m1 >>
rect 145 148 146 149 
<< m2 >>
rect 145 148 146 149 
<< m1 >>
rect 147 148 148 149 
<< m1 >>
rect 148 148 149 149 
<< m1 >>
rect 149 148 150 149 
<< m1 >>
rect 150 148 151 149 
<< m1 >>
rect 151 148 152 149 
<< m1 >>
rect 152 148 153 149 
<< m1 >>
rect 153 148 154 149 
<< m1 >>
rect 154 148 155 149 
<< m1 >>
rect 155 148 156 149 
<< m1 >>
rect 156 148 157 149 
<< m1 >>
rect 157 148 158 149 
<< m1 >>
rect 158 148 159 149 
<< m1 >>
rect 163 148 164 149 
<< m2 >>
rect 163 148 164 149 
<< m2c >>
rect 163 148 164 149 
<< m1 >>
rect 163 148 164 149 
<< m2 >>
rect 163 148 164 149 
<< m1 >>
rect 165 148 166 149 
<< m1 >>
rect 166 148 167 149 
<< m1 >>
rect 167 148 168 149 
<< m1 >>
rect 168 148 169 149 
<< m1 >>
rect 169 148 170 149 
<< m1 >>
rect 170 148 171 149 
<< m1 >>
rect 171 148 172 149 
<< m1 >>
rect 172 148 173 149 
<< m1 >>
rect 173 148 174 149 
<< m1 >>
rect 174 148 175 149 
<< m1 >>
rect 175 148 176 149 
<< m1 >>
rect 176 148 177 149 
<< m1 >>
rect 177 148 178 149 
<< m1 >>
rect 178 148 179 149 
<< m1 >>
rect 179 148 180 149 
<< m1 >>
rect 180 148 181 149 
<< m1 >>
rect 181 148 182 149 
<< m1 >>
rect 182 148 183 149 
<< m1 >>
rect 183 148 184 149 
<< m1 >>
rect 184 148 185 149 
<< m1 >>
rect 185 148 186 149 
<< m1 >>
rect 186 148 187 149 
<< m1 >>
rect 187 148 188 149 
<< m1 >>
rect 188 148 189 149 
<< m1 >>
rect 189 148 190 149 
<< m1 >>
rect 190 148 191 149 
<< m1 >>
rect 191 148 192 149 
<< m1 >>
rect 192 148 193 149 
<< m1 >>
rect 193 148 194 149 
<< m1 >>
rect 194 148 195 149 
<< m1 >>
rect 195 148 196 149 
<< m1 >>
rect 196 148 197 149 
<< m2 >>
rect 196 148 197 149 
<< m2c >>
rect 196 148 197 149 
<< m1 >>
rect 196 148 197 149 
<< m2 >>
rect 196 148 197 149 
<< m1 >>
rect 211 148 212 149 
<< m2 >>
rect 211 148 212 149 
<< m2c >>
rect 211 148 212 149 
<< m1 >>
rect 211 148 212 149 
<< m2 >>
rect 211 148 212 149 
<< m1 >>
rect 217 148 218 149 
<< m1 >>
rect 218 148 219 149 
<< m1 >>
rect 219 148 220 149 
<< m1 >>
rect 220 148 221 149 
<< m1 >>
rect 221 148 222 149 
<< m2 >>
rect 221 148 222 149 
<< m1 >>
rect 222 148 223 149 
<< m1 >>
rect 223 148 224 149 
<< m1 >>
rect 224 148 225 149 
<< m1 >>
rect 225 148 226 149 
<< m1 >>
rect 226 148 227 149 
<< m2 >>
rect 226 148 227 149 
<< m1 >>
rect 227 148 228 149 
<< m1 >>
rect 228 148 229 149 
<< m1 >>
rect 229 148 230 149 
<< m1 >>
rect 230 148 231 149 
<< m1 >>
rect 231 148 232 149 
<< m1 >>
rect 232 148 233 149 
<< m1 >>
rect 235 148 236 149 
<< m1 >>
rect 244 148 245 149 
<< m1 >>
rect 278 148 279 149 
<< m1 >>
rect 280 148 281 149 
<< m2 >>
rect 280 148 281 149 
<< m1 >>
rect 334 148 335 149 
<< m1 >>
rect 343 148 344 149 
<< m1 >>
rect 361 148 362 149 
<< m1 >>
rect 366 148 367 149 
<< m1 >>
rect 370 148 371 149 
<< m1 >>
rect 379 148 380 149 
<< m2 >>
rect 379 148 380 149 
<< m1 >>
rect 412 148 413 149 
<< m1 >>
rect 415 148 416 149 
<< m1 >>
rect 417 148 418 149 
<< m1 >>
rect 419 148 420 149 
<< m1 >>
rect 433 148 434 149 
<< m1 >>
rect 442 148 443 149 
<< m1 >>
rect 456 148 457 149 
<< m1 >>
rect 469 148 470 149 
<< m1 >>
rect 470 148 471 149 
<< m1 >>
rect 471 148 472 149 
<< m1 >>
rect 472 148 473 149 
<< m1 >>
rect 473 148 474 149 
<< m1 >>
rect 474 148 475 149 
<< m1 >>
rect 475 148 476 149 
<< m1 >>
rect 476 148 477 149 
<< m1 >>
rect 477 148 478 149 
<< m1 >>
rect 478 148 479 149 
<< m2 >>
rect 478 148 479 149 
<< m1 >>
rect 479 148 480 149 
<< m1 >>
rect 480 148 481 149 
<< m1 >>
rect 481 148 482 149 
<< m1 >>
rect 482 148 483 149 
<< m1 >>
rect 483 148 484 149 
<< m1 >>
rect 484 148 485 149 
<< m1 >>
rect 485 148 486 149 
<< m1 >>
rect 486 148 487 149 
<< m1 >>
rect 487 148 488 149 
<< m1 >>
rect 488 148 489 149 
<< m1 >>
rect 489 148 490 149 
<< m1 >>
rect 490 148 491 149 
<< m1 >>
rect 491 148 492 149 
<< m1 >>
rect 492 148 493 149 
<< m1 >>
rect 493 148 494 149 
<< m1 >>
rect 494 148 495 149 
<< m1 >>
rect 495 148 496 149 
<< m1 >>
rect 496 148 497 149 
<< m1 >>
rect 497 148 498 149 
<< m1 >>
rect 498 148 499 149 
<< m1 >>
rect 499 148 500 149 
<< m1 >>
rect 500 148 501 149 
<< m1 >>
rect 501 148 502 149 
<< m1 >>
rect 502 148 503 149 
<< m1 >>
rect 503 148 504 149 
<< m1 >>
rect 504 148 505 149 
<< m1 >>
rect 505 148 506 149 
<< m1 >>
rect 506 148 507 149 
<< m1 >>
rect 507 148 508 149 
<< m1 >>
rect 508 148 509 149 
<< m1 >>
rect 509 148 510 149 
<< m1 >>
rect 510 148 511 149 
<< m1 >>
rect 511 148 512 149 
<< m1 >>
rect 512 148 513 149 
<< m1 >>
rect 513 148 514 149 
<< m1 >>
rect 514 148 515 149 
<< m1 >>
rect 515 148 516 149 
<< m1 >>
rect 516 148 517 149 
<< m1 >>
rect 517 148 518 149 
<< m1 >>
rect 518 148 519 149 
<< m1 >>
rect 519 148 520 149 
<< m1 >>
rect 520 148 521 149 
<< m1 >>
rect 37 149 38 150 
<< m1 >>
rect 64 149 65 150 
<< m2 >>
rect 97 149 98 150 
<< m1 >>
rect 98 149 99 150 
<< m1 >>
rect 100 149 101 150 
<< m1 >>
rect 109 149 110 150 
<< m1 >>
rect 114 149 115 150 
<< m1 >>
rect 118 149 119 150 
<< m2 >>
rect 118 149 119 150 
<< m1 >>
rect 127 149 128 150 
<< m2 >>
rect 127 149 128 150 
<< m1 >>
rect 129 149 130 150 
<< m1 >>
rect 131 149 132 150 
<< m2 >>
rect 145 149 146 150 
<< m2 >>
rect 146 149 147 150 
<< m2 >>
rect 147 149 148 150 
<< m2 >>
rect 148 149 149 150 
<< m2 >>
rect 149 149 150 150 
<< m2 >>
rect 150 149 151 150 
<< m2 >>
rect 151 149 152 150 
<< m2 >>
rect 152 149 153 150 
<< m2 >>
rect 153 149 154 150 
<< m2 >>
rect 154 149 155 150 
<< m2 >>
rect 155 149 156 150 
<< m2 >>
rect 156 149 157 150 
<< m2 >>
rect 157 149 158 150 
<< m2 >>
rect 158 149 159 150 
<< m2 >>
rect 159 149 160 150 
<< m2 >>
rect 163 149 164 150 
<< m2 >>
rect 164 149 165 150 
<< m2 >>
rect 165 149 166 150 
<< m2 >>
rect 166 149 167 150 
<< m2 >>
rect 167 149 168 150 
<< m2 >>
rect 168 149 169 150 
<< m2 >>
rect 169 149 170 150 
<< m2 >>
rect 170 149 171 150 
<< m2 >>
rect 171 149 172 150 
<< m2 >>
rect 172 149 173 150 
<< m2 >>
rect 173 149 174 150 
<< m2 >>
rect 174 149 175 150 
<< m2 >>
rect 175 149 176 150 
<< m2 >>
rect 176 149 177 150 
<< m2 >>
rect 177 149 178 150 
<< m2 >>
rect 178 149 179 150 
<< m2 >>
rect 179 149 180 150 
<< m2 >>
rect 180 149 181 150 
<< m2 >>
rect 181 149 182 150 
<< m2 >>
rect 182 149 183 150 
<< m2 >>
rect 183 149 184 150 
<< m2 >>
rect 184 149 185 150 
<< m2 >>
rect 185 149 186 150 
<< m2 >>
rect 186 149 187 150 
<< m2 >>
rect 187 149 188 150 
<< m2 >>
rect 188 149 189 150 
<< m2 >>
rect 189 149 190 150 
<< m2 >>
rect 190 149 191 150 
<< m2 >>
rect 191 149 192 150 
<< m2 >>
rect 192 149 193 150 
<< m2 >>
rect 193 149 194 150 
<< m2 >>
rect 194 149 195 150 
<< m2 >>
rect 196 149 197 150 
<< m2 >>
rect 197 149 198 150 
<< m2 >>
rect 211 149 212 150 
<< m2 >>
rect 212 149 213 150 
<< m2 >>
rect 213 149 214 150 
<< m2 >>
rect 214 149 215 150 
<< m2 >>
rect 221 149 222 150 
<< m2 >>
rect 226 149 227 150 
<< m1 >>
rect 235 149 236 150 
<< m1 >>
rect 244 149 245 150 
<< m1 >>
rect 278 149 279 150 
<< m1 >>
rect 280 149 281 150 
<< m2 >>
rect 280 149 281 150 
<< m1 >>
rect 334 149 335 150 
<< m1 >>
rect 343 149 344 150 
<< m2 >>
rect 343 149 344 150 
<< m2c >>
rect 343 149 344 150 
<< m1 >>
rect 343 149 344 150 
<< m2 >>
rect 343 149 344 150 
<< m1 >>
rect 361 149 362 150 
<< m2 >>
rect 361 149 362 150 
<< m2c >>
rect 361 149 362 150 
<< m1 >>
rect 361 149 362 150 
<< m2 >>
rect 361 149 362 150 
<< m1 >>
rect 366 149 367 150 
<< m2 >>
rect 366 149 367 150 
<< m2c >>
rect 366 149 367 150 
<< m1 >>
rect 366 149 367 150 
<< m2 >>
rect 366 149 367 150 
<< m1 >>
rect 370 149 371 150 
<< m2 >>
rect 370 149 371 150 
<< m2c >>
rect 370 149 371 150 
<< m1 >>
rect 370 149 371 150 
<< m2 >>
rect 370 149 371 150 
<< m1 >>
rect 379 149 380 150 
<< m2 >>
rect 379 149 380 150 
<< m1 >>
rect 412 149 413 150 
<< m1 >>
rect 415 149 416 150 
<< m1 >>
rect 417 149 418 150 
<< m1 >>
rect 419 149 420 150 
<< m1 >>
rect 433 149 434 150 
<< m1 >>
rect 442 149 443 150 
<< m1 >>
rect 456 149 457 150 
<< m2 >>
rect 478 149 479 150 
<< m1 >>
rect 520 149 521 150 
<< m1 >>
rect 37 150 38 151 
<< m1 >>
rect 64 150 65 151 
<< m2 >>
rect 97 150 98 151 
<< m1 >>
rect 98 150 99 151 
<< m1 >>
rect 100 150 101 151 
<< m1 >>
rect 109 150 110 151 
<< m1 >>
rect 114 150 115 151 
<< m1 >>
rect 118 150 119 151 
<< m2 >>
rect 118 150 119 151 
<< m2 >>
rect 120 150 121 151 
<< m2 >>
rect 121 150 122 151 
<< m2 >>
rect 122 150 123 151 
<< m2 >>
rect 123 150 124 151 
<< m2 >>
rect 124 150 125 151 
<< m2 >>
rect 125 150 126 151 
<< m2 >>
rect 126 150 127 151 
<< m1 >>
rect 127 150 128 151 
<< m2 >>
rect 127 150 128 151 
<< m1 >>
rect 129 150 130 151 
<< m1 >>
rect 131 150 132 151 
<< m1 >>
rect 132 150 133 151 
<< m1 >>
rect 133 150 134 151 
<< m1 >>
rect 134 150 135 151 
<< m1 >>
rect 135 150 136 151 
<< m1 >>
rect 136 150 137 151 
<< m1 >>
rect 137 150 138 151 
<< m1 >>
rect 138 150 139 151 
<< m1 >>
rect 139 150 140 151 
<< m1 >>
rect 140 150 141 151 
<< m1 >>
rect 141 150 142 151 
<< m1 >>
rect 142 150 143 151 
<< m1 >>
rect 143 150 144 151 
<< m1 >>
rect 144 150 145 151 
<< m1 >>
rect 145 150 146 151 
<< m1 >>
rect 146 150 147 151 
<< m1 >>
rect 147 150 148 151 
<< m1 >>
rect 148 150 149 151 
<< m1 >>
rect 149 150 150 151 
<< m1 >>
rect 150 150 151 151 
<< m1 >>
rect 151 150 152 151 
<< m1 >>
rect 152 150 153 151 
<< m1 >>
rect 153 150 154 151 
<< m1 >>
rect 154 150 155 151 
<< m1 >>
rect 155 150 156 151 
<< m1 >>
rect 156 150 157 151 
<< m1 >>
rect 157 150 158 151 
<< m1 >>
rect 158 150 159 151 
<< m1 >>
rect 159 150 160 151 
<< m2 >>
rect 159 150 160 151 
<< m1 >>
rect 160 150 161 151 
<< m1 >>
rect 161 150 162 151 
<< m1 >>
rect 162 150 163 151 
<< m1 >>
rect 163 150 164 151 
<< m1 >>
rect 164 150 165 151 
<< m1 >>
rect 165 150 166 151 
<< m1 >>
rect 166 150 167 151 
<< m1 >>
rect 167 150 168 151 
<< m1 >>
rect 168 150 169 151 
<< m1 >>
rect 169 150 170 151 
<< m1 >>
rect 170 150 171 151 
<< m1 >>
rect 171 150 172 151 
<< m1 >>
rect 172 150 173 151 
<< m1 >>
rect 173 150 174 151 
<< m1 >>
rect 174 150 175 151 
<< m1 >>
rect 175 150 176 151 
<< m1 >>
rect 176 150 177 151 
<< m1 >>
rect 177 150 178 151 
<< m1 >>
rect 178 150 179 151 
<< m1 >>
rect 179 150 180 151 
<< m1 >>
rect 180 150 181 151 
<< m1 >>
rect 181 150 182 151 
<< m1 >>
rect 182 150 183 151 
<< m1 >>
rect 183 150 184 151 
<< m1 >>
rect 184 150 185 151 
<< m1 >>
rect 185 150 186 151 
<< m1 >>
rect 186 150 187 151 
<< m1 >>
rect 187 150 188 151 
<< m1 >>
rect 188 150 189 151 
<< m1 >>
rect 189 150 190 151 
<< m1 >>
rect 190 150 191 151 
<< m1 >>
rect 191 150 192 151 
<< m1 >>
rect 192 150 193 151 
<< m1 >>
rect 193 150 194 151 
<< m1 >>
rect 194 150 195 151 
<< m2 >>
rect 194 150 195 151 
<< m1 >>
rect 195 150 196 151 
<< m1 >>
rect 196 150 197 151 
<< m1 >>
rect 197 150 198 151 
<< m2 >>
rect 197 150 198 151 
<< m1 >>
rect 198 150 199 151 
<< m1 >>
rect 199 150 200 151 
<< m1 >>
rect 200 150 201 151 
<< m1 >>
rect 201 150 202 151 
<< m1 >>
rect 202 150 203 151 
<< m1 >>
rect 203 150 204 151 
<< m1 >>
rect 204 150 205 151 
<< m1 >>
rect 205 150 206 151 
<< m1 >>
rect 206 150 207 151 
<< m1 >>
rect 207 150 208 151 
<< m1 >>
rect 208 150 209 151 
<< m1 >>
rect 209 150 210 151 
<< m1 >>
rect 210 150 211 151 
<< m1 >>
rect 211 150 212 151 
<< m1 >>
rect 212 150 213 151 
<< m1 >>
rect 213 150 214 151 
<< m1 >>
rect 214 150 215 151 
<< m2 >>
rect 214 150 215 151 
<< m1 >>
rect 215 150 216 151 
<< m2 >>
rect 215 150 216 151 
<< m1 >>
rect 216 150 217 151 
<< m2 >>
rect 216 150 217 151 
<< m1 >>
rect 217 150 218 151 
<< m2 >>
rect 217 150 218 151 
<< m2 >>
rect 218 150 219 151 
<< m1 >>
rect 219 150 220 151 
<< m2 >>
rect 219 150 220 151 
<< m2c >>
rect 219 150 220 151 
<< m1 >>
rect 219 150 220 151 
<< m2 >>
rect 219 150 220 151 
<< m1 >>
rect 221 150 222 151 
<< m2 >>
rect 221 150 222 151 
<< m2c >>
rect 221 150 222 151 
<< m1 >>
rect 221 150 222 151 
<< m2 >>
rect 221 150 222 151 
<< m1 >>
rect 226 150 227 151 
<< m2 >>
rect 226 150 227 151 
<< m2c >>
rect 226 150 227 151 
<< m1 >>
rect 226 150 227 151 
<< m2 >>
rect 226 150 227 151 
<< m1 >>
rect 235 150 236 151 
<< m1 >>
rect 244 150 245 151 
<< m1 >>
rect 278 150 279 151 
<< m1 >>
rect 280 150 281 151 
<< m2 >>
rect 280 150 281 151 
<< m1 >>
rect 334 150 335 151 
<< m2 >>
rect 343 150 344 151 
<< m2 >>
rect 361 150 362 151 
<< m2 >>
rect 366 150 367 151 
<< m2 >>
rect 370 150 371 151 
<< m1 >>
rect 379 150 380 151 
<< m2 >>
rect 379 150 380 151 
<< m1 >>
rect 412 150 413 151 
<< m1 >>
rect 415 150 416 151 
<< m1 >>
rect 417 150 418 151 
<< m1 >>
rect 419 150 420 151 
<< m1 >>
rect 433 150 434 151 
<< m1 >>
rect 442 150 443 151 
<< m1 >>
rect 456 150 457 151 
<< m1 >>
rect 478 150 479 151 
<< m2 >>
rect 478 150 479 151 
<< m2c >>
rect 478 150 479 151 
<< m1 >>
rect 478 150 479 151 
<< m2 >>
rect 478 150 479 151 
<< m1 >>
rect 520 150 521 151 
<< m1 >>
rect 37 151 38 152 
<< m1 >>
rect 64 151 65 152 
<< m2 >>
rect 97 151 98 152 
<< m1 >>
rect 98 151 99 152 
<< m1 >>
rect 100 151 101 152 
<< m1 >>
rect 109 151 110 152 
<< m1 >>
rect 114 151 115 152 
<< m1 >>
rect 118 151 119 152 
<< m2 >>
rect 118 151 119 152 
<< m1 >>
rect 119 151 120 152 
<< m1 >>
rect 120 151 121 152 
<< m2 >>
rect 120 151 121 152 
<< m1 >>
rect 121 151 122 152 
<< m1 >>
rect 122 151 123 152 
<< m1 >>
rect 123 151 124 152 
<< m1 >>
rect 124 151 125 152 
<< m1 >>
rect 125 151 126 152 
<< m1 >>
rect 127 151 128 152 
<< m1 >>
rect 129 151 130 152 
<< m2 >>
rect 129 151 130 152 
<< m2c >>
rect 129 151 130 152 
<< m1 >>
rect 129 151 130 152 
<< m2 >>
rect 129 151 130 152 
<< m2 >>
rect 130 151 131 152 
<< m2 >>
rect 131 151 132 152 
<< m2 >>
rect 132 151 133 152 
<< m2 >>
rect 133 151 134 152 
<< m2 >>
rect 134 151 135 152 
<< m2 >>
rect 135 151 136 152 
<< m2 >>
rect 136 151 137 152 
<< m2 >>
rect 137 151 138 152 
<< m2 >>
rect 138 151 139 152 
<< m2 >>
rect 139 151 140 152 
<< m2 >>
rect 140 151 141 152 
<< m2 >>
rect 141 151 142 152 
<< m2 >>
rect 142 151 143 152 
<< m2 >>
rect 143 151 144 152 
<< m2 >>
rect 144 151 145 152 
<< m2 >>
rect 145 151 146 152 
<< m2 >>
rect 146 151 147 152 
<< m2 >>
rect 147 151 148 152 
<< m2 >>
rect 148 151 149 152 
<< m2 >>
rect 149 151 150 152 
<< m2 >>
rect 150 151 151 152 
<< m2 >>
rect 151 151 152 152 
<< m2 >>
rect 152 151 153 152 
<< m2 >>
rect 153 151 154 152 
<< m2 >>
rect 154 151 155 152 
<< m2 >>
rect 155 151 156 152 
<< m2 >>
rect 156 151 157 152 
<< m2 >>
rect 157 151 158 152 
<< m2 >>
rect 159 151 160 152 
<< m2 >>
rect 160 151 161 152 
<< m2 >>
rect 161 151 162 152 
<< m2 >>
rect 162 151 163 152 
<< m2 >>
rect 163 151 164 152 
<< m2 >>
rect 164 151 165 152 
<< m2 >>
rect 165 151 166 152 
<< m2 >>
rect 166 151 167 152 
<< m2 >>
rect 167 151 168 152 
<< m2 >>
rect 168 151 169 152 
<< m2 >>
rect 169 151 170 152 
<< m2 >>
rect 170 151 171 152 
<< m2 >>
rect 171 151 172 152 
<< m2 >>
rect 172 151 173 152 
<< m2 >>
rect 173 151 174 152 
<< m2 >>
rect 174 151 175 152 
<< m2 >>
rect 175 151 176 152 
<< m2 >>
rect 176 151 177 152 
<< m2 >>
rect 194 151 195 152 
<< m2 >>
rect 197 151 198 152 
<< m2 >>
rect 199 151 200 152 
<< m2 >>
rect 200 151 201 152 
<< m2 >>
rect 201 151 202 152 
<< m2 >>
rect 202 151 203 152 
<< m2 >>
rect 203 151 204 152 
<< m2 >>
rect 204 151 205 152 
<< m2 >>
rect 205 151 206 152 
<< m2 >>
rect 206 151 207 152 
<< m2 >>
rect 207 151 208 152 
<< m2 >>
rect 208 151 209 152 
<< m2 >>
rect 209 151 210 152 
<< m2 >>
rect 210 151 211 152 
<< m2 >>
rect 211 151 212 152 
<< m2 >>
rect 212 151 213 152 
<< m1 >>
rect 217 151 218 152 
<< m1 >>
rect 219 151 220 152 
<< m2 >>
rect 221 151 222 152 
<< m1 >>
rect 226 151 227 152 
<< m1 >>
rect 228 151 229 152 
<< m1 >>
rect 229 151 230 152 
<< m1 >>
rect 230 151 231 152 
<< m1 >>
rect 231 151 232 152 
<< m1 >>
rect 232 151 233 152 
<< m1 >>
rect 233 151 234 152 
<< m2 >>
rect 233 151 234 152 
<< m2c >>
rect 233 151 234 152 
<< m1 >>
rect 233 151 234 152 
<< m2 >>
rect 233 151 234 152 
<< m2 >>
rect 234 151 235 152 
<< m1 >>
rect 235 151 236 152 
<< m2 >>
rect 235 151 236 152 
<< m2 >>
rect 236 151 237 152 
<< m1 >>
rect 237 151 238 152 
<< m2 >>
rect 237 151 238 152 
<< m2c >>
rect 237 151 238 152 
<< m1 >>
rect 237 151 238 152 
<< m2 >>
rect 237 151 238 152 
<< m1 >>
rect 244 151 245 152 
<< m1 >>
rect 278 151 279 152 
<< m1 >>
rect 280 151 281 152 
<< m2 >>
rect 280 151 281 152 
<< m1 >>
rect 283 151 284 152 
<< m1 >>
rect 284 151 285 152 
<< m1 >>
rect 285 151 286 152 
<< m1 >>
rect 286 151 287 152 
<< m1 >>
rect 287 151 288 152 
<< m1 >>
rect 288 151 289 152 
<< m1 >>
rect 289 151 290 152 
<< m1 >>
rect 290 151 291 152 
<< m1 >>
rect 291 151 292 152 
<< m1 >>
rect 292 151 293 152 
<< m1 >>
rect 293 151 294 152 
<< m1 >>
rect 294 151 295 152 
<< m1 >>
rect 295 151 296 152 
<< m1 >>
rect 296 151 297 152 
<< m1 >>
rect 297 151 298 152 
<< m1 >>
rect 298 151 299 152 
<< m1 >>
rect 299 151 300 152 
<< m1 >>
rect 300 151 301 152 
<< m1 >>
rect 301 151 302 152 
<< m1 >>
rect 302 151 303 152 
<< m1 >>
rect 303 151 304 152 
<< m1 >>
rect 304 151 305 152 
<< m1 >>
rect 305 151 306 152 
<< m1 >>
rect 306 151 307 152 
<< m1 >>
rect 307 151 308 152 
<< m1 >>
rect 308 151 309 152 
<< m1 >>
rect 309 151 310 152 
<< m1 >>
rect 310 151 311 152 
<< m1 >>
rect 311 151 312 152 
<< m1 >>
rect 312 151 313 152 
<< m1 >>
rect 313 151 314 152 
<< m1 >>
rect 314 151 315 152 
<< m1 >>
rect 315 151 316 152 
<< m1 >>
rect 316 151 317 152 
<< m1 >>
rect 317 151 318 152 
<< m1 >>
rect 318 151 319 152 
<< m1 >>
rect 319 151 320 152 
<< m1 >>
rect 320 151 321 152 
<< m1 >>
rect 321 151 322 152 
<< m1 >>
rect 322 151 323 152 
<< m1 >>
rect 334 151 335 152 
<< m1 >>
rect 336 151 337 152 
<< m1 >>
rect 337 151 338 152 
<< m1 >>
rect 338 151 339 152 
<< m1 >>
rect 339 151 340 152 
<< m1 >>
rect 340 151 341 152 
<< m1 >>
rect 341 151 342 152 
<< m1 >>
rect 342 151 343 152 
<< m1 >>
rect 343 151 344 152 
<< m2 >>
rect 343 151 344 152 
<< m1 >>
rect 344 151 345 152 
<< m1 >>
rect 345 151 346 152 
<< m1 >>
rect 346 151 347 152 
<< m1 >>
rect 347 151 348 152 
<< m1 >>
rect 348 151 349 152 
<< m1 >>
rect 349 151 350 152 
<< m1 >>
rect 350 151 351 152 
<< m1 >>
rect 351 151 352 152 
<< m1 >>
rect 352 151 353 152 
<< m1 >>
rect 353 151 354 152 
<< m1 >>
rect 354 151 355 152 
<< m1 >>
rect 355 151 356 152 
<< m1 >>
rect 356 151 357 152 
<< m1 >>
rect 357 151 358 152 
<< m1 >>
rect 358 151 359 152 
<< m1 >>
rect 359 151 360 152 
<< m1 >>
rect 360 151 361 152 
<< m1 >>
rect 361 151 362 152 
<< m2 >>
rect 361 151 362 152 
<< m1 >>
rect 362 151 363 152 
<< m1 >>
rect 363 151 364 152 
<< m1 >>
rect 364 151 365 152 
<< m1 >>
rect 365 151 366 152 
<< m1 >>
rect 366 151 367 152 
<< m2 >>
rect 366 151 367 152 
<< m1 >>
rect 367 151 368 152 
<< m1 >>
rect 368 151 369 152 
<< m1 >>
rect 369 151 370 152 
<< m1 >>
rect 370 151 371 152 
<< m2 >>
rect 370 151 371 152 
<< m1 >>
rect 371 151 372 152 
<< m1 >>
rect 372 151 373 152 
<< m1 >>
rect 373 151 374 152 
<< m1 >>
rect 374 151 375 152 
<< m1 >>
rect 375 151 376 152 
<< m1 >>
rect 376 151 377 152 
<< m1 >>
rect 379 151 380 152 
<< m2 >>
rect 379 151 380 152 
<< m1 >>
rect 412 151 413 152 
<< m1 >>
rect 415 151 416 152 
<< m1 >>
rect 417 151 418 152 
<< m1 >>
rect 419 151 420 152 
<< m1 >>
rect 433 151 434 152 
<< m1 >>
rect 442 151 443 152 
<< m1 >>
rect 456 151 457 152 
<< m1 >>
rect 478 151 479 152 
<< m1 >>
rect 520 151 521 152 
<< m1 >>
rect 37 152 38 153 
<< m1 >>
rect 64 152 65 153 
<< m2 >>
rect 97 152 98 153 
<< m1 >>
rect 98 152 99 153 
<< m1 >>
rect 100 152 101 153 
<< m1 >>
rect 109 152 110 153 
<< m1 >>
rect 114 152 115 153 
<< m2 >>
rect 118 152 119 153 
<< m2 >>
rect 120 152 121 153 
<< m1 >>
rect 125 152 126 153 
<< m1 >>
rect 127 152 128 153 
<< m1 >>
rect 157 152 158 153 
<< m2 >>
rect 157 152 158 153 
<< m2c >>
rect 157 152 158 153 
<< m1 >>
rect 157 152 158 153 
<< m2 >>
rect 157 152 158 153 
<< m1 >>
rect 176 152 177 153 
<< m2 >>
rect 176 152 177 153 
<< m2c >>
rect 176 152 177 153 
<< m1 >>
rect 176 152 177 153 
<< m2 >>
rect 176 152 177 153 
<< m1 >>
rect 177 152 178 153 
<< m1 >>
rect 178 152 179 153 
<< m1 >>
rect 194 152 195 153 
<< m2 >>
rect 194 152 195 153 
<< m2c >>
rect 194 152 195 153 
<< m1 >>
rect 194 152 195 153 
<< m2 >>
rect 194 152 195 153 
<< m1 >>
rect 195 152 196 153 
<< m1 >>
rect 196 152 197 153 
<< m2 >>
rect 197 152 198 153 
<< m1 >>
rect 199 152 200 153 
<< m2 >>
rect 199 152 200 153 
<< m2c >>
rect 199 152 200 153 
<< m1 >>
rect 199 152 200 153 
<< m2 >>
rect 199 152 200 153 
<< m1 >>
rect 212 152 213 153 
<< m2 >>
rect 212 152 213 153 
<< m2c >>
rect 212 152 213 153 
<< m1 >>
rect 212 152 213 153 
<< m2 >>
rect 212 152 213 153 
<< m1 >>
rect 213 152 214 153 
<< m1 >>
rect 214 152 215 153 
<< m1 >>
rect 217 152 218 153 
<< m1 >>
rect 219 152 220 153 
<< m1 >>
rect 220 152 221 153 
<< m1 >>
rect 221 152 222 153 
<< m2 >>
rect 221 152 222 153 
<< m1 >>
rect 222 152 223 153 
<< m1 >>
rect 223 152 224 153 
<< m1 >>
rect 224 152 225 153 
<< m2 >>
rect 224 152 225 153 
<< m2c >>
rect 224 152 225 153 
<< m1 >>
rect 224 152 225 153 
<< m2 >>
rect 224 152 225 153 
<< m2 >>
rect 225 152 226 153 
<< m1 >>
rect 226 152 227 153 
<< m2 >>
rect 226 152 227 153 
<< m2 >>
rect 227 152 228 153 
<< m1 >>
rect 228 152 229 153 
<< m2 >>
rect 228 152 229 153 
<< m2c >>
rect 228 152 229 153 
<< m1 >>
rect 228 152 229 153 
<< m2 >>
rect 228 152 229 153 
<< m1 >>
rect 235 152 236 153 
<< m1 >>
rect 237 152 238 153 
<< m1 >>
rect 244 152 245 153 
<< m1 >>
rect 278 152 279 153 
<< m1 >>
rect 280 152 281 153 
<< m2 >>
rect 280 152 281 153 
<< m1 >>
rect 283 152 284 153 
<< m1 >>
rect 322 152 323 153 
<< m1 >>
rect 334 152 335 153 
<< m1 >>
rect 336 152 337 153 
<< m2 >>
rect 343 152 344 153 
<< m2 >>
rect 361 152 362 153 
<< m2 >>
rect 366 152 367 153 
<< m2 >>
rect 370 152 371 153 
<< m1 >>
rect 376 152 377 153 
<< m1 >>
rect 379 152 380 153 
<< m2 >>
rect 379 152 380 153 
<< m1 >>
rect 412 152 413 153 
<< m1 >>
rect 415 152 416 153 
<< m1 >>
rect 417 152 418 153 
<< m1 >>
rect 419 152 420 153 
<< m1 >>
rect 433 152 434 153 
<< m1 >>
rect 442 152 443 153 
<< m1 >>
rect 456 152 457 153 
<< m1 >>
rect 478 152 479 153 
<< m1 >>
rect 520 152 521 153 
<< m1 >>
rect 37 153 38 154 
<< m1 >>
rect 64 153 65 154 
<< m2 >>
rect 97 153 98 154 
<< m1 >>
rect 98 153 99 154 
<< m1 >>
rect 100 153 101 154 
<< m1 >>
rect 109 153 110 154 
<< m1 >>
rect 114 153 115 154 
<< m1 >>
rect 118 153 119 154 
<< m2 >>
rect 118 153 119 154 
<< m1 >>
rect 119 153 120 154 
<< m1 >>
rect 120 153 121 154 
<< m2 >>
rect 120 153 121 154 
<< m2c >>
rect 120 153 121 154 
<< m1 >>
rect 120 153 121 154 
<< m2 >>
rect 120 153 121 154 
<< m1 >>
rect 125 153 126 154 
<< m1 >>
rect 127 153 128 154 
<< m1 >>
rect 157 153 158 154 
<< m1 >>
rect 178 153 179 154 
<< m1 >>
rect 196 153 197 154 
<< m2 >>
rect 197 153 198 154 
<< m1 >>
rect 199 153 200 154 
<< m1 >>
rect 214 153 215 154 
<< m1 >>
rect 217 153 218 154 
<< m2 >>
rect 221 153 222 154 
<< m1 >>
rect 226 153 227 154 
<< m1 >>
rect 235 153 236 154 
<< m1 >>
rect 237 153 238 154 
<< m1 >>
rect 244 153 245 154 
<< m1 >>
rect 278 153 279 154 
<< m1 >>
rect 280 153 281 154 
<< m2 >>
rect 280 153 281 154 
<< m1 >>
rect 283 153 284 154 
<< m1 >>
rect 322 153 323 154 
<< m1 >>
rect 334 153 335 154 
<< m1 >>
rect 336 153 337 154 
<< m1 >>
rect 343 153 344 154 
<< m2 >>
rect 343 153 344 154 
<< m2c >>
rect 343 153 344 154 
<< m1 >>
rect 343 153 344 154 
<< m2 >>
rect 343 153 344 154 
<< m1 >>
rect 361 153 362 154 
<< m2 >>
rect 361 153 362 154 
<< m2c >>
rect 361 153 362 154 
<< m1 >>
rect 361 153 362 154 
<< m2 >>
rect 361 153 362 154 
<< m1 >>
rect 366 153 367 154 
<< m2 >>
rect 366 153 367 154 
<< m2c >>
rect 366 153 367 154 
<< m1 >>
rect 366 153 367 154 
<< m2 >>
rect 366 153 367 154 
<< m1 >>
rect 370 153 371 154 
<< m2 >>
rect 370 153 371 154 
<< m2c >>
rect 370 153 371 154 
<< m1 >>
rect 370 153 371 154 
<< m2 >>
rect 370 153 371 154 
<< m1 >>
rect 376 153 377 154 
<< m1 >>
rect 379 153 380 154 
<< m2 >>
rect 379 153 380 154 
<< m1 >>
rect 391 153 392 154 
<< m1 >>
rect 392 153 393 154 
<< m1 >>
rect 393 153 394 154 
<< m1 >>
rect 394 153 395 154 
<< m1 >>
rect 395 153 396 154 
<< m1 >>
rect 396 153 397 154 
<< m1 >>
rect 397 153 398 154 
<< m1 >>
rect 398 153 399 154 
<< m1 >>
rect 399 153 400 154 
<< m1 >>
rect 400 153 401 154 
<< m1 >>
rect 401 153 402 154 
<< m1 >>
rect 402 153 403 154 
<< m1 >>
rect 403 153 404 154 
<< m1 >>
rect 404 153 405 154 
<< m1 >>
rect 405 153 406 154 
<< m1 >>
rect 406 153 407 154 
<< m1 >>
rect 412 153 413 154 
<< m1 >>
rect 415 153 416 154 
<< m1 >>
rect 417 153 418 154 
<< m1 >>
rect 419 153 420 154 
<< m1 >>
rect 433 153 434 154 
<< m1 >>
rect 442 153 443 154 
<< m1 >>
rect 456 153 457 154 
<< m1 >>
rect 478 153 479 154 
<< m1 >>
rect 520 153 521 154 
<< m1 >>
rect 37 154 38 155 
<< m1 >>
rect 64 154 65 155 
<< m2 >>
rect 97 154 98 155 
<< m1 >>
rect 98 154 99 155 
<< m1 >>
rect 100 154 101 155 
<< m1 >>
rect 109 154 110 155 
<< m1 >>
rect 114 154 115 155 
<< m1 >>
rect 118 154 119 155 
<< m2 >>
rect 118 154 119 155 
<< m1 >>
rect 125 154 126 155 
<< m2 >>
rect 125 154 126 155 
<< m2c >>
rect 125 154 126 155 
<< m1 >>
rect 125 154 126 155 
<< m2 >>
rect 125 154 126 155 
<< m2 >>
rect 126 154 127 155 
<< m1 >>
rect 127 154 128 155 
<< m2 >>
rect 127 154 128 155 
<< m2 >>
rect 128 154 129 155 
<< m1 >>
rect 129 154 130 155 
<< m2 >>
rect 129 154 130 155 
<< m2c >>
rect 129 154 130 155 
<< m1 >>
rect 129 154 130 155 
<< m2 >>
rect 129 154 130 155 
<< m1 >>
rect 130 154 131 155 
<< m1 >>
rect 131 154 132 155 
<< m1 >>
rect 132 154 133 155 
<< m1 >>
rect 133 154 134 155 
<< m1 >>
rect 134 154 135 155 
<< m1 >>
rect 135 154 136 155 
<< m1 >>
rect 136 154 137 155 
<< m1 >>
rect 137 154 138 155 
<< m1 >>
rect 138 154 139 155 
<< m1 >>
rect 139 154 140 155 
<< m1 >>
rect 157 154 158 155 
<< m1 >>
rect 178 154 179 155 
<< m1 >>
rect 196 154 197 155 
<< m2 >>
rect 197 154 198 155 
<< m2 >>
rect 198 154 199 155 
<< m1 >>
rect 199 154 200 155 
<< m2 >>
rect 199 154 200 155 
<< m1 >>
rect 214 154 215 155 
<< m1 >>
rect 217 154 218 155 
<< m1 >>
rect 221 154 222 155 
<< m2 >>
rect 221 154 222 155 
<< m2c >>
rect 221 154 222 155 
<< m1 >>
rect 221 154 222 155 
<< m2 >>
rect 221 154 222 155 
<< m1 >>
rect 226 154 227 155 
<< m1 >>
rect 235 154 236 155 
<< m1 >>
rect 237 154 238 155 
<< m1 >>
rect 244 154 245 155 
<< m1 >>
rect 250 154 251 155 
<< m1 >>
rect 251 154 252 155 
<< m1 >>
rect 252 154 253 155 
<< m1 >>
rect 253 154 254 155 
<< m1 >>
rect 278 154 279 155 
<< m1 >>
rect 280 154 281 155 
<< m2 >>
rect 280 154 281 155 
<< m1 >>
rect 283 154 284 155 
<< m1 >>
rect 322 154 323 155 
<< m1 >>
rect 334 154 335 155 
<< m1 >>
rect 336 154 337 155 
<< m1 >>
rect 343 154 344 155 
<< m1 >>
rect 345 154 346 155 
<< m1 >>
rect 346 154 347 155 
<< m1 >>
rect 347 154 348 155 
<< m1 >>
rect 348 154 349 155 
<< m1 >>
rect 349 154 350 155 
<< m1 >>
rect 350 154 351 155 
<< m1 >>
rect 351 154 352 155 
<< m1 >>
rect 352 154 353 155 
<< m1 >>
rect 353 154 354 155 
<< m1 >>
rect 354 154 355 155 
<< m1 >>
rect 355 154 356 155 
<< m1 >>
rect 361 154 362 155 
<< m2 >>
rect 366 154 367 155 
<< m1 >>
rect 370 154 371 155 
<< m1 >>
rect 376 154 377 155 
<< m1 >>
rect 379 154 380 155 
<< m2 >>
rect 379 154 380 155 
<< m1 >>
rect 391 154 392 155 
<< m1 >>
rect 406 154 407 155 
<< m1 >>
rect 412 154 413 155 
<< m1 >>
rect 415 154 416 155 
<< m1 >>
rect 417 154 418 155 
<< m1 >>
rect 419 154 420 155 
<< m1 >>
rect 433 154 434 155 
<< m1 >>
rect 442 154 443 155 
<< m1 >>
rect 456 154 457 155 
<< m1 >>
rect 478 154 479 155 
<< m1 >>
rect 520 154 521 155 
<< m1 >>
rect 37 155 38 156 
<< m1 >>
rect 64 155 65 156 
<< m2 >>
rect 97 155 98 156 
<< m1 >>
rect 98 155 99 156 
<< m1 >>
rect 100 155 101 156 
<< m1 >>
rect 109 155 110 156 
<< m1 >>
rect 114 155 115 156 
<< m1 >>
rect 118 155 119 156 
<< m2 >>
rect 118 155 119 156 
<< m1 >>
rect 127 155 128 156 
<< m1 >>
rect 139 155 140 156 
<< m1 >>
rect 157 155 158 156 
<< m1 >>
rect 178 155 179 156 
<< m1 >>
rect 196 155 197 156 
<< m1 >>
rect 199 155 200 156 
<< m2 >>
rect 199 155 200 156 
<< m1 >>
rect 214 155 215 156 
<< m1 >>
rect 217 155 218 156 
<< m1 >>
rect 221 155 222 156 
<< m1 >>
rect 226 155 227 156 
<< m1 >>
rect 235 155 236 156 
<< m1 >>
rect 237 155 238 156 
<< m1 >>
rect 244 155 245 156 
<< m1 >>
rect 250 155 251 156 
<< m1 >>
rect 253 155 254 156 
<< m1 >>
rect 278 155 279 156 
<< m1 >>
rect 280 155 281 156 
<< m2 >>
rect 280 155 281 156 
<< m1 >>
rect 283 155 284 156 
<< m1 >>
rect 322 155 323 156 
<< m1 >>
rect 334 155 335 156 
<< m1 >>
rect 336 155 337 156 
<< m1 >>
rect 343 155 344 156 
<< m1 >>
rect 345 155 346 156 
<< m1 >>
rect 355 155 356 156 
<< m1 >>
rect 361 155 362 156 
<< m1 >>
rect 362 155 363 156 
<< m1 >>
rect 363 155 364 156 
<< m1 >>
rect 364 155 365 156 
<< m1 >>
rect 365 155 366 156 
<< m1 >>
rect 366 155 367 156 
<< m2 >>
rect 366 155 367 156 
<< m1 >>
rect 367 155 368 156 
<< m1 >>
rect 368 155 369 156 
<< m2 >>
rect 368 155 369 156 
<< m2c >>
rect 368 155 369 156 
<< m1 >>
rect 368 155 369 156 
<< m2 >>
rect 368 155 369 156 
<< m2 >>
rect 369 155 370 156 
<< m1 >>
rect 370 155 371 156 
<< m1 >>
rect 376 155 377 156 
<< m1 >>
rect 379 155 380 156 
<< m2 >>
rect 379 155 380 156 
<< m1 >>
rect 391 155 392 156 
<< m1 >>
rect 406 155 407 156 
<< m1 >>
rect 412 155 413 156 
<< m1 >>
rect 415 155 416 156 
<< m1 >>
rect 417 155 418 156 
<< m1 >>
rect 419 155 420 156 
<< m1 >>
rect 433 155 434 156 
<< m1 >>
rect 442 155 443 156 
<< m1 >>
rect 456 155 457 156 
<< m1 >>
rect 478 155 479 156 
<< m1 >>
rect 520 155 521 156 
<< pdiffusion >>
rect 12 156 13 157 
<< pdiffusion >>
rect 13 156 14 157 
<< pdiffusion >>
rect 14 156 15 157 
<< pdiffusion >>
rect 15 156 16 157 
<< pdiffusion >>
rect 16 156 17 157 
<< pdiffusion >>
rect 17 156 18 157 
<< pdiffusion >>
rect 30 156 31 157 
<< pdiffusion >>
rect 31 156 32 157 
<< pdiffusion >>
rect 32 156 33 157 
<< pdiffusion >>
rect 33 156 34 157 
<< pdiffusion >>
rect 34 156 35 157 
<< pdiffusion >>
rect 35 156 36 157 
<< m1 >>
rect 37 156 38 157 
<< pdiffusion >>
rect 48 156 49 157 
<< pdiffusion >>
rect 49 156 50 157 
<< pdiffusion >>
rect 50 156 51 157 
<< pdiffusion >>
rect 51 156 52 157 
<< pdiffusion >>
rect 52 156 53 157 
<< pdiffusion >>
rect 53 156 54 157 
<< m1 >>
rect 64 156 65 157 
<< pdiffusion >>
rect 66 156 67 157 
<< pdiffusion >>
rect 67 156 68 157 
<< pdiffusion >>
rect 68 156 69 157 
<< pdiffusion >>
rect 69 156 70 157 
<< pdiffusion >>
rect 70 156 71 157 
<< pdiffusion >>
rect 71 156 72 157 
<< pdiffusion >>
rect 84 156 85 157 
<< pdiffusion >>
rect 85 156 86 157 
<< pdiffusion >>
rect 86 156 87 157 
<< pdiffusion >>
rect 87 156 88 157 
<< pdiffusion >>
rect 88 156 89 157 
<< pdiffusion >>
rect 89 156 90 157 
<< m2 >>
rect 97 156 98 157 
<< m1 >>
rect 98 156 99 157 
<< m1 >>
rect 100 156 101 157 
<< pdiffusion >>
rect 102 156 103 157 
<< pdiffusion >>
rect 103 156 104 157 
<< pdiffusion >>
rect 104 156 105 157 
<< pdiffusion >>
rect 105 156 106 157 
<< pdiffusion >>
rect 106 156 107 157 
<< pdiffusion >>
rect 107 156 108 157 
<< m1 >>
rect 109 156 110 157 
<< m1 >>
rect 114 156 115 157 
<< m1 >>
rect 118 156 119 157 
<< m2 >>
rect 118 156 119 157 
<< pdiffusion >>
rect 120 156 121 157 
<< pdiffusion >>
rect 121 156 122 157 
<< pdiffusion >>
rect 122 156 123 157 
<< pdiffusion >>
rect 123 156 124 157 
<< pdiffusion >>
rect 124 156 125 157 
<< pdiffusion >>
rect 125 156 126 157 
<< m1 >>
rect 127 156 128 157 
<< pdiffusion >>
rect 138 156 139 157 
<< m1 >>
rect 139 156 140 157 
<< pdiffusion >>
rect 139 156 140 157 
<< pdiffusion >>
rect 140 156 141 157 
<< pdiffusion >>
rect 141 156 142 157 
<< pdiffusion >>
rect 142 156 143 157 
<< pdiffusion >>
rect 143 156 144 157 
<< pdiffusion >>
rect 156 156 157 157 
<< m1 >>
rect 157 156 158 157 
<< pdiffusion >>
rect 157 156 158 157 
<< pdiffusion >>
rect 158 156 159 157 
<< pdiffusion >>
rect 159 156 160 157 
<< pdiffusion >>
rect 160 156 161 157 
<< pdiffusion >>
rect 161 156 162 157 
<< pdiffusion >>
rect 174 156 175 157 
<< pdiffusion >>
rect 175 156 176 157 
<< pdiffusion >>
rect 176 156 177 157 
<< pdiffusion >>
rect 177 156 178 157 
<< m1 >>
rect 178 156 179 157 
<< pdiffusion >>
rect 178 156 179 157 
<< pdiffusion >>
rect 179 156 180 157 
<< pdiffusion >>
rect 192 156 193 157 
<< pdiffusion >>
rect 193 156 194 157 
<< pdiffusion >>
rect 194 156 195 157 
<< pdiffusion >>
rect 195 156 196 157 
<< m1 >>
rect 196 156 197 157 
<< pdiffusion >>
rect 196 156 197 157 
<< pdiffusion >>
rect 197 156 198 157 
<< m1 >>
rect 199 156 200 157 
<< m2 >>
rect 199 156 200 157 
<< pdiffusion >>
rect 210 156 211 157 
<< pdiffusion >>
rect 211 156 212 157 
<< pdiffusion >>
rect 212 156 213 157 
<< pdiffusion >>
rect 213 156 214 157 
<< m1 >>
rect 214 156 215 157 
<< pdiffusion >>
rect 214 156 215 157 
<< pdiffusion >>
rect 215 156 216 157 
<< m1 >>
rect 217 156 218 157 
<< m1 >>
rect 221 156 222 157 
<< m1 >>
rect 226 156 227 157 
<< pdiffusion >>
rect 228 156 229 157 
<< pdiffusion >>
rect 229 156 230 157 
<< pdiffusion >>
rect 230 156 231 157 
<< pdiffusion >>
rect 231 156 232 157 
<< pdiffusion >>
rect 232 156 233 157 
<< pdiffusion >>
rect 233 156 234 157 
<< m1 >>
rect 235 156 236 157 
<< m1 >>
rect 237 156 238 157 
<< m1 >>
rect 244 156 245 157 
<< pdiffusion >>
rect 246 156 247 157 
<< pdiffusion >>
rect 247 156 248 157 
<< pdiffusion >>
rect 248 156 249 157 
<< pdiffusion >>
rect 249 156 250 157 
<< m1 >>
rect 250 156 251 157 
<< pdiffusion >>
rect 250 156 251 157 
<< pdiffusion >>
rect 251 156 252 157 
<< m1 >>
rect 253 156 254 157 
<< pdiffusion >>
rect 264 156 265 157 
<< pdiffusion >>
rect 265 156 266 157 
<< pdiffusion >>
rect 266 156 267 157 
<< pdiffusion >>
rect 267 156 268 157 
<< pdiffusion >>
rect 268 156 269 157 
<< pdiffusion >>
rect 269 156 270 157 
<< m1 >>
rect 278 156 279 157 
<< m1 >>
rect 280 156 281 157 
<< m2 >>
rect 280 156 281 157 
<< pdiffusion >>
rect 282 156 283 157 
<< m1 >>
rect 283 156 284 157 
<< pdiffusion >>
rect 283 156 284 157 
<< pdiffusion >>
rect 284 156 285 157 
<< pdiffusion >>
rect 285 156 286 157 
<< pdiffusion >>
rect 286 156 287 157 
<< pdiffusion >>
rect 287 156 288 157 
<< pdiffusion >>
rect 300 156 301 157 
<< pdiffusion >>
rect 301 156 302 157 
<< pdiffusion >>
rect 302 156 303 157 
<< pdiffusion >>
rect 303 156 304 157 
<< pdiffusion >>
rect 304 156 305 157 
<< pdiffusion >>
rect 305 156 306 157 
<< pdiffusion >>
rect 318 156 319 157 
<< pdiffusion >>
rect 319 156 320 157 
<< pdiffusion >>
rect 320 156 321 157 
<< pdiffusion >>
rect 321 156 322 157 
<< m1 >>
rect 322 156 323 157 
<< pdiffusion >>
rect 322 156 323 157 
<< pdiffusion >>
rect 323 156 324 157 
<< m1 >>
rect 334 156 335 157 
<< m1 >>
rect 336 156 337 157 
<< m1 >>
rect 343 156 344 157 
<< m1 >>
rect 345 156 346 157 
<< pdiffusion >>
rect 354 156 355 157 
<< m1 >>
rect 355 156 356 157 
<< pdiffusion >>
rect 355 156 356 157 
<< pdiffusion >>
rect 356 156 357 157 
<< pdiffusion >>
rect 357 156 358 157 
<< pdiffusion >>
rect 358 156 359 157 
<< pdiffusion >>
rect 359 156 360 157 
<< m2 >>
rect 366 156 367 157 
<< m2 >>
rect 369 156 370 157 
<< m1 >>
rect 370 156 371 157 
<< pdiffusion >>
rect 372 156 373 157 
<< pdiffusion >>
rect 373 156 374 157 
<< pdiffusion >>
rect 374 156 375 157 
<< pdiffusion >>
rect 375 156 376 157 
<< m1 >>
rect 376 156 377 157 
<< pdiffusion >>
rect 376 156 377 157 
<< pdiffusion >>
rect 377 156 378 157 
<< m1 >>
rect 379 156 380 157 
<< m2 >>
rect 379 156 380 157 
<< pdiffusion >>
rect 390 156 391 157 
<< m1 >>
rect 391 156 392 157 
<< pdiffusion >>
rect 391 156 392 157 
<< pdiffusion >>
rect 392 156 393 157 
<< pdiffusion >>
rect 393 156 394 157 
<< pdiffusion >>
rect 394 156 395 157 
<< pdiffusion >>
rect 395 156 396 157 
<< m1 >>
rect 406 156 407 157 
<< pdiffusion >>
rect 408 156 409 157 
<< pdiffusion >>
rect 409 156 410 157 
<< pdiffusion >>
rect 410 156 411 157 
<< pdiffusion >>
rect 411 156 412 157 
<< m1 >>
rect 412 156 413 157 
<< pdiffusion >>
rect 412 156 413 157 
<< pdiffusion >>
rect 413 156 414 157 
<< m1 >>
rect 415 156 416 157 
<< m1 >>
rect 417 156 418 157 
<< m1 >>
rect 419 156 420 157 
<< pdiffusion >>
rect 426 156 427 157 
<< pdiffusion >>
rect 427 156 428 157 
<< pdiffusion >>
rect 428 156 429 157 
<< pdiffusion >>
rect 429 156 430 157 
<< pdiffusion >>
rect 430 156 431 157 
<< pdiffusion >>
rect 431 156 432 157 
<< m1 >>
rect 433 156 434 157 
<< m1 >>
rect 442 156 443 157 
<< pdiffusion >>
rect 444 156 445 157 
<< pdiffusion >>
rect 445 156 446 157 
<< pdiffusion >>
rect 446 156 447 157 
<< pdiffusion >>
rect 447 156 448 157 
<< pdiffusion >>
rect 448 156 449 157 
<< pdiffusion >>
rect 449 156 450 157 
<< m1 >>
rect 456 156 457 157 
<< pdiffusion >>
rect 462 156 463 157 
<< pdiffusion >>
rect 463 156 464 157 
<< pdiffusion >>
rect 464 156 465 157 
<< pdiffusion >>
rect 465 156 466 157 
<< pdiffusion >>
rect 466 156 467 157 
<< pdiffusion >>
rect 467 156 468 157 
<< m1 >>
rect 478 156 479 157 
<< pdiffusion >>
rect 480 156 481 157 
<< pdiffusion >>
rect 481 156 482 157 
<< pdiffusion >>
rect 482 156 483 157 
<< pdiffusion >>
rect 483 156 484 157 
<< pdiffusion >>
rect 484 156 485 157 
<< pdiffusion >>
rect 485 156 486 157 
<< pdiffusion >>
rect 498 156 499 157 
<< pdiffusion >>
rect 499 156 500 157 
<< pdiffusion >>
rect 500 156 501 157 
<< pdiffusion >>
rect 501 156 502 157 
<< pdiffusion >>
rect 502 156 503 157 
<< pdiffusion >>
rect 503 156 504 157 
<< pdiffusion >>
rect 516 156 517 157 
<< pdiffusion >>
rect 517 156 518 157 
<< pdiffusion >>
rect 518 156 519 157 
<< pdiffusion >>
rect 519 156 520 157 
<< m1 >>
rect 520 156 521 157 
<< pdiffusion >>
rect 520 156 521 157 
<< pdiffusion >>
rect 521 156 522 157 
<< pdiffusion >>
rect 12 157 13 158 
<< pdiffusion >>
rect 13 157 14 158 
<< pdiffusion >>
rect 14 157 15 158 
<< pdiffusion >>
rect 15 157 16 158 
<< pdiffusion >>
rect 16 157 17 158 
<< pdiffusion >>
rect 17 157 18 158 
<< pdiffusion >>
rect 30 157 31 158 
<< pdiffusion >>
rect 31 157 32 158 
<< pdiffusion >>
rect 32 157 33 158 
<< pdiffusion >>
rect 33 157 34 158 
<< pdiffusion >>
rect 34 157 35 158 
<< pdiffusion >>
rect 35 157 36 158 
<< m1 >>
rect 37 157 38 158 
<< pdiffusion >>
rect 48 157 49 158 
<< pdiffusion >>
rect 49 157 50 158 
<< pdiffusion >>
rect 50 157 51 158 
<< pdiffusion >>
rect 51 157 52 158 
<< pdiffusion >>
rect 52 157 53 158 
<< pdiffusion >>
rect 53 157 54 158 
<< m1 >>
rect 64 157 65 158 
<< pdiffusion >>
rect 66 157 67 158 
<< pdiffusion >>
rect 67 157 68 158 
<< pdiffusion >>
rect 68 157 69 158 
<< pdiffusion >>
rect 69 157 70 158 
<< pdiffusion >>
rect 70 157 71 158 
<< pdiffusion >>
rect 71 157 72 158 
<< pdiffusion >>
rect 84 157 85 158 
<< pdiffusion >>
rect 85 157 86 158 
<< pdiffusion >>
rect 86 157 87 158 
<< pdiffusion >>
rect 87 157 88 158 
<< pdiffusion >>
rect 88 157 89 158 
<< pdiffusion >>
rect 89 157 90 158 
<< m2 >>
rect 97 157 98 158 
<< m1 >>
rect 98 157 99 158 
<< m1 >>
rect 100 157 101 158 
<< pdiffusion >>
rect 102 157 103 158 
<< pdiffusion >>
rect 103 157 104 158 
<< pdiffusion >>
rect 104 157 105 158 
<< pdiffusion >>
rect 105 157 106 158 
<< pdiffusion >>
rect 106 157 107 158 
<< pdiffusion >>
rect 107 157 108 158 
<< m1 >>
rect 109 157 110 158 
<< m1 >>
rect 114 157 115 158 
<< m1 >>
rect 118 157 119 158 
<< m2 >>
rect 118 157 119 158 
<< pdiffusion >>
rect 120 157 121 158 
<< pdiffusion >>
rect 121 157 122 158 
<< pdiffusion >>
rect 122 157 123 158 
<< pdiffusion >>
rect 123 157 124 158 
<< pdiffusion >>
rect 124 157 125 158 
<< pdiffusion >>
rect 125 157 126 158 
<< m1 >>
rect 127 157 128 158 
<< pdiffusion >>
rect 138 157 139 158 
<< pdiffusion >>
rect 139 157 140 158 
<< pdiffusion >>
rect 140 157 141 158 
<< pdiffusion >>
rect 141 157 142 158 
<< pdiffusion >>
rect 142 157 143 158 
<< pdiffusion >>
rect 143 157 144 158 
<< pdiffusion >>
rect 156 157 157 158 
<< pdiffusion >>
rect 157 157 158 158 
<< pdiffusion >>
rect 158 157 159 158 
<< pdiffusion >>
rect 159 157 160 158 
<< pdiffusion >>
rect 160 157 161 158 
<< pdiffusion >>
rect 161 157 162 158 
<< pdiffusion >>
rect 174 157 175 158 
<< pdiffusion >>
rect 175 157 176 158 
<< pdiffusion >>
rect 176 157 177 158 
<< pdiffusion >>
rect 177 157 178 158 
<< pdiffusion >>
rect 178 157 179 158 
<< pdiffusion >>
rect 179 157 180 158 
<< pdiffusion >>
rect 192 157 193 158 
<< pdiffusion >>
rect 193 157 194 158 
<< pdiffusion >>
rect 194 157 195 158 
<< pdiffusion >>
rect 195 157 196 158 
<< pdiffusion >>
rect 196 157 197 158 
<< pdiffusion >>
rect 197 157 198 158 
<< m1 >>
rect 199 157 200 158 
<< m2 >>
rect 199 157 200 158 
<< pdiffusion >>
rect 210 157 211 158 
<< pdiffusion >>
rect 211 157 212 158 
<< pdiffusion >>
rect 212 157 213 158 
<< pdiffusion >>
rect 213 157 214 158 
<< pdiffusion >>
rect 214 157 215 158 
<< pdiffusion >>
rect 215 157 216 158 
<< m1 >>
rect 217 157 218 158 
<< m1 >>
rect 221 157 222 158 
<< m1 >>
rect 226 157 227 158 
<< pdiffusion >>
rect 228 157 229 158 
<< pdiffusion >>
rect 229 157 230 158 
<< pdiffusion >>
rect 230 157 231 158 
<< pdiffusion >>
rect 231 157 232 158 
<< pdiffusion >>
rect 232 157 233 158 
<< pdiffusion >>
rect 233 157 234 158 
<< m1 >>
rect 235 157 236 158 
<< m1 >>
rect 237 157 238 158 
<< m1 >>
rect 244 157 245 158 
<< pdiffusion >>
rect 246 157 247 158 
<< pdiffusion >>
rect 247 157 248 158 
<< pdiffusion >>
rect 248 157 249 158 
<< pdiffusion >>
rect 249 157 250 158 
<< pdiffusion >>
rect 250 157 251 158 
<< pdiffusion >>
rect 251 157 252 158 
<< m1 >>
rect 253 157 254 158 
<< pdiffusion >>
rect 264 157 265 158 
<< pdiffusion >>
rect 265 157 266 158 
<< pdiffusion >>
rect 266 157 267 158 
<< pdiffusion >>
rect 267 157 268 158 
<< pdiffusion >>
rect 268 157 269 158 
<< pdiffusion >>
rect 269 157 270 158 
<< m1 >>
rect 278 157 279 158 
<< m1 >>
rect 280 157 281 158 
<< m2 >>
rect 280 157 281 158 
<< pdiffusion >>
rect 282 157 283 158 
<< pdiffusion >>
rect 283 157 284 158 
<< pdiffusion >>
rect 284 157 285 158 
<< pdiffusion >>
rect 285 157 286 158 
<< pdiffusion >>
rect 286 157 287 158 
<< pdiffusion >>
rect 287 157 288 158 
<< pdiffusion >>
rect 300 157 301 158 
<< pdiffusion >>
rect 301 157 302 158 
<< pdiffusion >>
rect 302 157 303 158 
<< pdiffusion >>
rect 303 157 304 158 
<< pdiffusion >>
rect 304 157 305 158 
<< pdiffusion >>
rect 305 157 306 158 
<< pdiffusion >>
rect 318 157 319 158 
<< pdiffusion >>
rect 319 157 320 158 
<< pdiffusion >>
rect 320 157 321 158 
<< pdiffusion >>
rect 321 157 322 158 
<< pdiffusion >>
rect 322 157 323 158 
<< pdiffusion >>
rect 323 157 324 158 
<< m1 >>
rect 334 157 335 158 
<< m1 >>
rect 336 157 337 158 
<< m1 >>
rect 343 157 344 158 
<< m1 >>
rect 345 157 346 158 
<< pdiffusion >>
rect 354 157 355 158 
<< pdiffusion >>
rect 355 157 356 158 
<< pdiffusion >>
rect 356 157 357 158 
<< pdiffusion >>
rect 357 157 358 158 
<< pdiffusion >>
rect 358 157 359 158 
<< pdiffusion >>
rect 359 157 360 158 
<< m1 >>
rect 366 157 367 158 
<< m2 >>
rect 366 157 367 158 
<< m2c >>
rect 366 157 367 158 
<< m1 >>
rect 366 157 367 158 
<< m2 >>
rect 366 157 367 158 
<< m2 >>
rect 369 157 370 158 
<< m1 >>
rect 370 157 371 158 
<< pdiffusion >>
rect 372 157 373 158 
<< pdiffusion >>
rect 373 157 374 158 
<< pdiffusion >>
rect 374 157 375 158 
<< pdiffusion >>
rect 375 157 376 158 
<< pdiffusion >>
rect 376 157 377 158 
<< pdiffusion >>
rect 377 157 378 158 
<< m1 >>
rect 379 157 380 158 
<< m2 >>
rect 379 157 380 158 
<< pdiffusion >>
rect 390 157 391 158 
<< pdiffusion >>
rect 391 157 392 158 
<< pdiffusion >>
rect 392 157 393 158 
<< pdiffusion >>
rect 393 157 394 158 
<< pdiffusion >>
rect 394 157 395 158 
<< pdiffusion >>
rect 395 157 396 158 
<< m1 >>
rect 406 157 407 158 
<< pdiffusion >>
rect 408 157 409 158 
<< pdiffusion >>
rect 409 157 410 158 
<< pdiffusion >>
rect 410 157 411 158 
<< pdiffusion >>
rect 411 157 412 158 
<< pdiffusion >>
rect 412 157 413 158 
<< pdiffusion >>
rect 413 157 414 158 
<< m1 >>
rect 415 157 416 158 
<< m1 >>
rect 417 157 418 158 
<< m1 >>
rect 419 157 420 158 
<< pdiffusion >>
rect 426 157 427 158 
<< pdiffusion >>
rect 427 157 428 158 
<< pdiffusion >>
rect 428 157 429 158 
<< pdiffusion >>
rect 429 157 430 158 
<< pdiffusion >>
rect 430 157 431 158 
<< pdiffusion >>
rect 431 157 432 158 
<< m1 >>
rect 433 157 434 158 
<< m1 >>
rect 442 157 443 158 
<< pdiffusion >>
rect 444 157 445 158 
<< pdiffusion >>
rect 445 157 446 158 
<< pdiffusion >>
rect 446 157 447 158 
<< pdiffusion >>
rect 447 157 448 158 
<< pdiffusion >>
rect 448 157 449 158 
<< pdiffusion >>
rect 449 157 450 158 
<< m1 >>
rect 456 157 457 158 
<< pdiffusion >>
rect 462 157 463 158 
<< pdiffusion >>
rect 463 157 464 158 
<< pdiffusion >>
rect 464 157 465 158 
<< pdiffusion >>
rect 465 157 466 158 
<< pdiffusion >>
rect 466 157 467 158 
<< pdiffusion >>
rect 467 157 468 158 
<< m1 >>
rect 478 157 479 158 
<< pdiffusion >>
rect 480 157 481 158 
<< pdiffusion >>
rect 481 157 482 158 
<< pdiffusion >>
rect 482 157 483 158 
<< pdiffusion >>
rect 483 157 484 158 
<< pdiffusion >>
rect 484 157 485 158 
<< pdiffusion >>
rect 485 157 486 158 
<< pdiffusion >>
rect 498 157 499 158 
<< pdiffusion >>
rect 499 157 500 158 
<< pdiffusion >>
rect 500 157 501 158 
<< pdiffusion >>
rect 501 157 502 158 
<< pdiffusion >>
rect 502 157 503 158 
<< pdiffusion >>
rect 503 157 504 158 
<< pdiffusion >>
rect 516 157 517 158 
<< pdiffusion >>
rect 517 157 518 158 
<< pdiffusion >>
rect 518 157 519 158 
<< pdiffusion >>
rect 519 157 520 158 
<< pdiffusion >>
rect 520 157 521 158 
<< pdiffusion >>
rect 521 157 522 158 
<< pdiffusion >>
rect 12 158 13 159 
<< pdiffusion >>
rect 13 158 14 159 
<< pdiffusion >>
rect 14 158 15 159 
<< pdiffusion >>
rect 15 158 16 159 
<< pdiffusion >>
rect 16 158 17 159 
<< pdiffusion >>
rect 17 158 18 159 
<< pdiffusion >>
rect 30 158 31 159 
<< pdiffusion >>
rect 31 158 32 159 
<< pdiffusion >>
rect 32 158 33 159 
<< pdiffusion >>
rect 33 158 34 159 
<< pdiffusion >>
rect 34 158 35 159 
<< pdiffusion >>
rect 35 158 36 159 
<< m1 >>
rect 37 158 38 159 
<< pdiffusion >>
rect 48 158 49 159 
<< pdiffusion >>
rect 49 158 50 159 
<< pdiffusion >>
rect 50 158 51 159 
<< pdiffusion >>
rect 51 158 52 159 
<< pdiffusion >>
rect 52 158 53 159 
<< pdiffusion >>
rect 53 158 54 159 
<< m1 >>
rect 64 158 65 159 
<< pdiffusion >>
rect 66 158 67 159 
<< pdiffusion >>
rect 67 158 68 159 
<< pdiffusion >>
rect 68 158 69 159 
<< pdiffusion >>
rect 69 158 70 159 
<< pdiffusion >>
rect 70 158 71 159 
<< pdiffusion >>
rect 71 158 72 159 
<< pdiffusion >>
rect 84 158 85 159 
<< pdiffusion >>
rect 85 158 86 159 
<< pdiffusion >>
rect 86 158 87 159 
<< pdiffusion >>
rect 87 158 88 159 
<< pdiffusion >>
rect 88 158 89 159 
<< pdiffusion >>
rect 89 158 90 159 
<< m2 >>
rect 97 158 98 159 
<< m1 >>
rect 98 158 99 159 
<< m1 >>
rect 100 158 101 159 
<< pdiffusion >>
rect 102 158 103 159 
<< pdiffusion >>
rect 103 158 104 159 
<< pdiffusion >>
rect 104 158 105 159 
<< pdiffusion >>
rect 105 158 106 159 
<< pdiffusion >>
rect 106 158 107 159 
<< pdiffusion >>
rect 107 158 108 159 
<< m1 >>
rect 109 158 110 159 
<< m1 >>
rect 114 158 115 159 
<< m1 >>
rect 118 158 119 159 
<< m2 >>
rect 118 158 119 159 
<< pdiffusion >>
rect 120 158 121 159 
<< pdiffusion >>
rect 121 158 122 159 
<< pdiffusion >>
rect 122 158 123 159 
<< pdiffusion >>
rect 123 158 124 159 
<< pdiffusion >>
rect 124 158 125 159 
<< pdiffusion >>
rect 125 158 126 159 
<< m1 >>
rect 127 158 128 159 
<< pdiffusion >>
rect 138 158 139 159 
<< pdiffusion >>
rect 139 158 140 159 
<< pdiffusion >>
rect 140 158 141 159 
<< pdiffusion >>
rect 141 158 142 159 
<< pdiffusion >>
rect 142 158 143 159 
<< pdiffusion >>
rect 143 158 144 159 
<< pdiffusion >>
rect 156 158 157 159 
<< pdiffusion >>
rect 157 158 158 159 
<< pdiffusion >>
rect 158 158 159 159 
<< pdiffusion >>
rect 159 158 160 159 
<< pdiffusion >>
rect 160 158 161 159 
<< pdiffusion >>
rect 161 158 162 159 
<< pdiffusion >>
rect 174 158 175 159 
<< pdiffusion >>
rect 175 158 176 159 
<< pdiffusion >>
rect 176 158 177 159 
<< pdiffusion >>
rect 177 158 178 159 
<< pdiffusion >>
rect 178 158 179 159 
<< pdiffusion >>
rect 179 158 180 159 
<< pdiffusion >>
rect 192 158 193 159 
<< pdiffusion >>
rect 193 158 194 159 
<< pdiffusion >>
rect 194 158 195 159 
<< pdiffusion >>
rect 195 158 196 159 
<< pdiffusion >>
rect 196 158 197 159 
<< pdiffusion >>
rect 197 158 198 159 
<< m1 >>
rect 199 158 200 159 
<< m2 >>
rect 199 158 200 159 
<< pdiffusion >>
rect 210 158 211 159 
<< pdiffusion >>
rect 211 158 212 159 
<< pdiffusion >>
rect 212 158 213 159 
<< pdiffusion >>
rect 213 158 214 159 
<< pdiffusion >>
rect 214 158 215 159 
<< pdiffusion >>
rect 215 158 216 159 
<< m1 >>
rect 217 158 218 159 
<< m1 >>
rect 221 158 222 159 
<< m1 >>
rect 226 158 227 159 
<< pdiffusion >>
rect 228 158 229 159 
<< pdiffusion >>
rect 229 158 230 159 
<< pdiffusion >>
rect 230 158 231 159 
<< pdiffusion >>
rect 231 158 232 159 
<< pdiffusion >>
rect 232 158 233 159 
<< pdiffusion >>
rect 233 158 234 159 
<< m1 >>
rect 235 158 236 159 
<< m1 >>
rect 237 158 238 159 
<< m1 >>
rect 244 158 245 159 
<< pdiffusion >>
rect 246 158 247 159 
<< pdiffusion >>
rect 247 158 248 159 
<< pdiffusion >>
rect 248 158 249 159 
<< pdiffusion >>
rect 249 158 250 159 
<< pdiffusion >>
rect 250 158 251 159 
<< pdiffusion >>
rect 251 158 252 159 
<< m1 >>
rect 253 158 254 159 
<< pdiffusion >>
rect 264 158 265 159 
<< pdiffusion >>
rect 265 158 266 159 
<< pdiffusion >>
rect 266 158 267 159 
<< pdiffusion >>
rect 267 158 268 159 
<< pdiffusion >>
rect 268 158 269 159 
<< pdiffusion >>
rect 269 158 270 159 
<< m1 >>
rect 278 158 279 159 
<< m1 >>
rect 280 158 281 159 
<< m2 >>
rect 280 158 281 159 
<< pdiffusion >>
rect 282 158 283 159 
<< pdiffusion >>
rect 283 158 284 159 
<< pdiffusion >>
rect 284 158 285 159 
<< pdiffusion >>
rect 285 158 286 159 
<< pdiffusion >>
rect 286 158 287 159 
<< pdiffusion >>
rect 287 158 288 159 
<< pdiffusion >>
rect 300 158 301 159 
<< pdiffusion >>
rect 301 158 302 159 
<< pdiffusion >>
rect 302 158 303 159 
<< pdiffusion >>
rect 303 158 304 159 
<< pdiffusion >>
rect 304 158 305 159 
<< pdiffusion >>
rect 305 158 306 159 
<< pdiffusion >>
rect 318 158 319 159 
<< pdiffusion >>
rect 319 158 320 159 
<< pdiffusion >>
rect 320 158 321 159 
<< pdiffusion >>
rect 321 158 322 159 
<< pdiffusion >>
rect 322 158 323 159 
<< pdiffusion >>
rect 323 158 324 159 
<< m1 >>
rect 334 158 335 159 
<< m1 >>
rect 336 158 337 159 
<< m1 >>
rect 343 158 344 159 
<< m1 >>
rect 345 158 346 159 
<< pdiffusion >>
rect 354 158 355 159 
<< pdiffusion >>
rect 355 158 356 159 
<< pdiffusion >>
rect 356 158 357 159 
<< pdiffusion >>
rect 357 158 358 159 
<< pdiffusion >>
rect 358 158 359 159 
<< pdiffusion >>
rect 359 158 360 159 
<< m1 >>
rect 366 158 367 159 
<< m2 >>
rect 369 158 370 159 
<< m1 >>
rect 370 158 371 159 
<< pdiffusion >>
rect 372 158 373 159 
<< pdiffusion >>
rect 373 158 374 159 
<< pdiffusion >>
rect 374 158 375 159 
<< pdiffusion >>
rect 375 158 376 159 
<< pdiffusion >>
rect 376 158 377 159 
<< pdiffusion >>
rect 377 158 378 159 
<< m1 >>
rect 379 158 380 159 
<< m2 >>
rect 379 158 380 159 
<< pdiffusion >>
rect 390 158 391 159 
<< pdiffusion >>
rect 391 158 392 159 
<< pdiffusion >>
rect 392 158 393 159 
<< pdiffusion >>
rect 393 158 394 159 
<< pdiffusion >>
rect 394 158 395 159 
<< pdiffusion >>
rect 395 158 396 159 
<< m1 >>
rect 406 158 407 159 
<< pdiffusion >>
rect 408 158 409 159 
<< pdiffusion >>
rect 409 158 410 159 
<< pdiffusion >>
rect 410 158 411 159 
<< pdiffusion >>
rect 411 158 412 159 
<< pdiffusion >>
rect 412 158 413 159 
<< pdiffusion >>
rect 413 158 414 159 
<< m1 >>
rect 415 158 416 159 
<< m1 >>
rect 417 158 418 159 
<< m1 >>
rect 419 158 420 159 
<< pdiffusion >>
rect 426 158 427 159 
<< pdiffusion >>
rect 427 158 428 159 
<< pdiffusion >>
rect 428 158 429 159 
<< pdiffusion >>
rect 429 158 430 159 
<< pdiffusion >>
rect 430 158 431 159 
<< pdiffusion >>
rect 431 158 432 159 
<< m1 >>
rect 433 158 434 159 
<< m1 >>
rect 442 158 443 159 
<< pdiffusion >>
rect 444 158 445 159 
<< pdiffusion >>
rect 445 158 446 159 
<< pdiffusion >>
rect 446 158 447 159 
<< pdiffusion >>
rect 447 158 448 159 
<< pdiffusion >>
rect 448 158 449 159 
<< pdiffusion >>
rect 449 158 450 159 
<< m1 >>
rect 456 158 457 159 
<< pdiffusion >>
rect 462 158 463 159 
<< pdiffusion >>
rect 463 158 464 159 
<< pdiffusion >>
rect 464 158 465 159 
<< pdiffusion >>
rect 465 158 466 159 
<< pdiffusion >>
rect 466 158 467 159 
<< pdiffusion >>
rect 467 158 468 159 
<< m1 >>
rect 478 158 479 159 
<< pdiffusion >>
rect 480 158 481 159 
<< pdiffusion >>
rect 481 158 482 159 
<< pdiffusion >>
rect 482 158 483 159 
<< pdiffusion >>
rect 483 158 484 159 
<< pdiffusion >>
rect 484 158 485 159 
<< pdiffusion >>
rect 485 158 486 159 
<< pdiffusion >>
rect 498 158 499 159 
<< pdiffusion >>
rect 499 158 500 159 
<< pdiffusion >>
rect 500 158 501 159 
<< pdiffusion >>
rect 501 158 502 159 
<< pdiffusion >>
rect 502 158 503 159 
<< pdiffusion >>
rect 503 158 504 159 
<< pdiffusion >>
rect 516 158 517 159 
<< pdiffusion >>
rect 517 158 518 159 
<< pdiffusion >>
rect 518 158 519 159 
<< pdiffusion >>
rect 519 158 520 159 
<< pdiffusion >>
rect 520 158 521 159 
<< pdiffusion >>
rect 521 158 522 159 
<< pdiffusion >>
rect 12 159 13 160 
<< pdiffusion >>
rect 13 159 14 160 
<< pdiffusion >>
rect 14 159 15 160 
<< pdiffusion >>
rect 15 159 16 160 
<< pdiffusion >>
rect 16 159 17 160 
<< pdiffusion >>
rect 17 159 18 160 
<< pdiffusion >>
rect 30 159 31 160 
<< pdiffusion >>
rect 31 159 32 160 
<< pdiffusion >>
rect 32 159 33 160 
<< pdiffusion >>
rect 33 159 34 160 
<< pdiffusion >>
rect 34 159 35 160 
<< pdiffusion >>
rect 35 159 36 160 
<< m1 >>
rect 37 159 38 160 
<< pdiffusion >>
rect 48 159 49 160 
<< pdiffusion >>
rect 49 159 50 160 
<< pdiffusion >>
rect 50 159 51 160 
<< pdiffusion >>
rect 51 159 52 160 
<< pdiffusion >>
rect 52 159 53 160 
<< pdiffusion >>
rect 53 159 54 160 
<< m1 >>
rect 64 159 65 160 
<< pdiffusion >>
rect 66 159 67 160 
<< pdiffusion >>
rect 67 159 68 160 
<< pdiffusion >>
rect 68 159 69 160 
<< pdiffusion >>
rect 69 159 70 160 
<< pdiffusion >>
rect 70 159 71 160 
<< pdiffusion >>
rect 71 159 72 160 
<< pdiffusion >>
rect 84 159 85 160 
<< pdiffusion >>
rect 85 159 86 160 
<< pdiffusion >>
rect 86 159 87 160 
<< pdiffusion >>
rect 87 159 88 160 
<< pdiffusion >>
rect 88 159 89 160 
<< pdiffusion >>
rect 89 159 90 160 
<< m2 >>
rect 97 159 98 160 
<< m1 >>
rect 98 159 99 160 
<< m1 >>
rect 100 159 101 160 
<< pdiffusion >>
rect 102 159 103 160 
<< pdiffusion >>
rect 103 159 104 160 
<< pdiffusion >>
rect 104 159 105 160 
<< pdiffusion >>
rect 105 159 106 160 
<< pdiffusion >>
rect 106 159 107 160 
<< pdiffusion >>
rect 107 159 108 160 
<< m1 >>
rect 109 159 110 160 
<< m1 >>
rect 114 159 115 160 
<< m1 >>
rect 118 159 119 160 
<< m2 >>
rect 118 159 119 160 
<< pdiffusion >>
rect 120 159 121 160 
<< pdiffusion >>
rect 121 159 122 160 
<< pdiffusion >>
rect 122 159 123 160 
<< pdiffusion >>
rect 123 159 124 160 
<< pdiffusion >>
rect 124 159 125 160 
<< pdiffusion >>
rect 125 159 126 160 
<< m1 >>
rect 127 159 128 160 
<< pdiffusion >>
rect 138 159 139 160 
<< pdiffusion >>
rect 139 159 140 160 
<< pdiffusion >>
rect 140 159 141 160 
<< pdiffusion >>
rect 141 159 142 160 
<< pdiffusion >>
rect 142 159 143 160 
<< pdiffusion >>
rect 143 159 144 160 
<< pdiffusion >>
rect 156 159 157 160 
<< pdiffusion >>
rect 157 159 158 160 
<< pdiffusion >>
rect 158 159 159 160 
<< pdiffusion >>
rect 159 159 160 160 
<< pdiffusion >>
rect 160 159 161 160 
<< pdiffusion >>
rect 161 159 162 160 
<< pdiffusion >>
rect 174 159 175 160 
<< pdiffusion >>
rect 175 159 176 160 
<< pdiffusion >>
rect 176 159 177 160 
<< pdiffusion >>
rect 177 159 178 160 
<< pdiffusion >>
rect 178 159 179 160 
<< pdiffusion >>
rect 179 159 180 160 
<< pdiffusion >>
rect 192 159 193 160 
<< pdiffusion >>
rect 193 159 194 160 
<< pdiffusion >>
rect 194 159 195 160 
<< pdiffusion >>
rect 195 159 196 160 
<< pdiffusion >>
rect 196 159 197 160 
<< pdiffusion >>
rect 197 159 198 160 
<< m1 >>
rect 199 159 200 160 
<< m2 >>
rect 199 159 200 160 
<< pdiffusion >>
rect 210 159 211 160 
<< pdiffusion >>
rect 211 159 212 160 
<< pdiffusion >>
rect 212 159 213 160 
<< pdiffusion >>
rect 213 159 214 160 
<< pdiffusion >>
rect 214 159 215 160 
<< pdiffusion >>
rect 215 159 216 160 
<< m1 >>
rect 217 159 218 160 
<< m1 >>
rect 221 159 222 160 
<< m1 >>
rect 226 159 227 160 
<< pdiffusion >>
rect 228 159 229 160 
<< pdiffusion >>
rect 229 159 230 160 
<< pdiffusion >>
rect 230 159 231 160 
<< pdiffusion >>
rect 231 159 232 160 
<< pdiffusion >>
rect 232 159 233 160 
<< pdiffusion >>
rect 233 159 234 160 
<< m1 >>
rect 235 159 236 160 
<< m1 >>
rect 237 159 238 160 
<< m1 >>
rect 244 159 245 160 
<< pdiffusion >>
rect 246 159 247 160 
<< pdiffusion >>
rect 247 159 248 160 
<< pdiffusion >>
rect 248 159 249 160 
<< pdiffusion >>
rect 249 159 250 160 
<< pdiffusion >>
rect 250 159 251 160 
<< pdiffusion >>
rect 251 159 252 160 
<< m1 >>
rect 253 159 254 160 
<< pdiffusion >>
rect 264 159 265 160 
<< pdiffusion >>
rect 265 159 266 160 
<< pdiffusion >>
rect 266 159 267 160 
<< pdiffusion >>
rect 267 159 268 160 
<< pdiffusion >>
rect 268 159 269 160 
<< pdiffusion >>
rect 269 159 270 160 
<< m1 >>
rect 278 159 279 160 
<< m1 >>
rect 280 159 281 160 
<< m2 >>
rect 280 159 281 160 
<< pdiffusion >>
rect 282 159 283 160 
<< pdiffusion >>
rect 283 159 284 160 
<< pdiffusion >>
rect 284 159 285 160 
<< pdiffusion >>
rect 285 159 286 160 
<< pdiffusion >>
rect 286 159 287 160 
<< pdiffusion >>
rect 287 159 288 160 
<< pdiffusion >>
rect 300 159 301 160 
<< pdiffusion >>
rect 301 159 302 160 
<< pdiffusion >>
rect 302 159 303 160 
<< pdiffusion >>
rect 303 159 304 160 
<< pdiffusion >>
rect 304 159 305 160 
<< pdiffusion >>
rect 305 159 306 160 
<< pdiffusion >>
rect 318 159 319 160 
<< pdiffusion >>
rect 319 159 320 160 
<< pdiffusion >>
rect 320 159 321 160 
<< pdiffusion >>
rect 321 159 322 160 
<< pdiffusion >>
rect 322 159 323 160 
<< pdiffusion >>
rect 323 159 324 160 
<< m1 >>
rect 334 159 335 160 
<< m1 >>
rect 336 159 337 160 
<< m1 >>
rect 343 159 344 160 
<< m1 >>
rect 345 159 346 160 
<< pdiffusion >>
rect 354 159 355 160 
<< pdiffusion >>
rect 355 159 356 160 
<< pdiffusion >>
rect 356 159 357 160 
<< pdiffusion >>
rect 357 159 358 160 
<< pdiffusion >>
rect 358 159 359 160 
<< pdiffusion >>
rect 359 159 360 160 
<< m1 >>
rect 366 159 367 160 
<< m2 >>
rect 369 159 370 160 
<< m1 >>
rect 370 159 371 160 
<< pdiffusion >>
rect 372 159 373 160 
<< pdiffusion >>
rect 373 159 374 160 
<< pdiffusion >>
rect 374 159 375 160 
<< pdiffusion >>
rect 375 159 376 160 
<< pdiffusion >>
rect 376 159 377 160 
<< pdiffusion >>
rect 377 159 378 160 
<< m1 >>
rect 379 159 380 160 
<< m2 >>
rect 379 159 380 160 
<< pdiffusion >>
rect 390 159 391 160 
<< pdiffusion >>
rect 391 159 392 160 
<< pdiffusion >>
rect 392 159 393 160 
<< pdiffusion >>
rect 393 159 394 160 
<< pdiffusion >>
rect 394 159 395 160 
<< pdiffusion >>
rect 395 159 396 160 
<< m1 >>
rect 406 159 407 160 
<< pdiffusion >>
rect 408 159 409 160 
<< pdiffusion >>
rect 409 159 410 160 
<< pdiffusion >>
rect 410 159 411 160 
<< pdiffusion >>
rect 411 159 412 160 
<< pdiffusion >>
rect 412 159 413 160 
<< pdiffusion >>
rect 413 159 414 160 
<< m1 >>
rect 415 159 416 160 
<< m1 >>
rect 417 159 418 160 
<< m1 >>
rect 419 159 420 160 
<< pdiffusion >>
rect 426 159 427 160 
<< pdiffusion >>
rect 427 159 428 160 
<< pdiffusion >>
rect 428 159 429 160 
<< pdiffusion >>
rect 429 159 430 160 
<< pdiffusion >>
rect 430 159 431 160 
<< pdiffusion >>
rect 431 159 432 160 
<< m1 >>
rect 433 159 434 160 
<< m1 >>
rect 442 159 443 160 
<< pdiffusion >>
rect 444 159 445 160 
<< pdiffusion >>
rect 445 159 446 160 
<< pdiffusion >>
rect 446 159 447 160 
<< pdiffusion >>
rect 447 159 448 160 
<< pdiffusion >>
rect 448 159 449 160 
<< pdiffusion >>
rect 449 159 450 160 
<< m1 >>
rect 456 159 457 160 
<< pdiffusion >>
rect 462 159 463 160 
<< pdiffusion >>
rect 463 159 464 160 
<< pdiffusion >>
rect 464 159 465 160 
<< pdiffusion >>
rect 465 159 466 160 
<< pdiffusion >>
rect 466 159 467 160 
<< pdiffusion >>
rect 467 159 468 160 
<< m1 >>
rect 478 159 479 160 
<< pdiffusion >>
rect 480 159 481 160 
<< pdiffusion >>
rect 481 159 482 160 
<< pdiffusion >>
rect 482 159 483 160 
<< pdiffusion >>
rect 483 159 484 160 
<< pdiffusion >>
rect 484 159 485 160 
<< pdiffusion >>
rect 485 159 486 160 
<< pdiffusion >>
rect 498 159 499 160 
<< pdiffusion >>
rect 499 159 500 160 
<< pdiffusion >>
rect 500 159 501 160 
<< pdiffusion >>
rect 501 159 502 160 
<< pdiffusion >>
rect 502 159 503 160 
<< pdiffusion >>
rect 503 159 504 160 
<< pdiffusion >>
rect 516 159 517 160 
<< pdiffusion >>
rect 517 159 518 160 
<< pdiffusion >>
rect 518 159 519 160 
<< pdiffusion >>
rect 519 159 520 160 
<< pdiffusion >>
rect 520 159 521 160 
<< pdiffusion >>
rect 521 159 522 160 
<< pdiffusion >>
rect 12 160 13 161 
<< pdiffusion >>
rect 13 160 14 161 
<< pdiffusion >>
rect 14 160 15 161 
<< pdiffusion >>
rect 15 160 16 161 
<< pdiffusion >>
rect 16 160 17 161 
<< pdiffusion >>
rect 17 160 18 161 
<< pdiffusion >>
rect 30 160 31 161 
<< pdiffusion >>
rect 31 160 32 161 
<< pdiffusion >>
rect 32 160 33 161 
<< pdiffusion >>
rect 33 160 34 161 
<< pdiffusion >>
rect 34 160 35 161 
<< pdiffusion >>
rect 35 160 36 161 
<< m1 >>
rect 37 160 38 161 
<< pdiffusion >>
rect 48 160 49 161 
<< pdiffusion >>
rect 49 160 50 161 
<< pdiffusion >>
rect 50 160 51 161 
<< pdiffusion >>
rect 51 160 52 161 
<< pdiffusion >>
rect 52 160 53 161 
<< pdiffusion >>
rect 53 160 54 161 
<< m1 >>
rect 64 160 65 161 
<< pdiffusion >>
rect 66 160 67 161 
<< pdiffusion >>
rect 67 160 68 161 
<< pdiffusion >>
rect 68 160 69 161 
<< pdiffusion >>
rect 69 160 70 161 
<< pdiffusion >>
rect 70 160 71 161 
<< pdiffusion >>
rect 71 160 72 161 
<< pdiffusion >>
rect 84 160 85 161 
<< pdiffusion >>
rect 85 160 86 161 
<< pdiffusion >>
rect 86 160 87 161 
<< pdiffusion >>
rect 87 160 88 161 
<< pdiffusion >>
rect 88 160 89 161 
<< pdiffusion >>
rect 89 160 90 161 
<< m2 >>
rect 97 160 98 161 
<< m1 >>
rect 98 160 99 161 
<< m1 >>
rect 100 160 101 161 
<< pdiffusion >>
rect 102 160 103 161 
<< pdiffusion >>
rect 103 160 104 161 
<< pdiffusion >>
rect 104 160 105 161 
<< pdiffusion >>
rect 105 160 106 161 
<< pdiffusion >>
rect 106 160 107 161 
<< pdiffusion >>
rect 107 160 108 161 
<< m1 >>
rect 109 160 110 161 
<< m1 >>
rect 114 160 115 161 
<< m1 >>
rect 118 160 119 161 
<< m2 >>
rect 118 160 119 161 
<< pdiffusion >>
rect 120 160 121 161 
<< pdiffusion >>
rect 121 160 122 161 
<< pdiffusion >>
rect 122 160 123 161 
<< pdiffusion >>
rect 123 160 124 161 
<< pdiffusion >>
rect 124 160 125 161 
<< pdiffusion >>
rect 125 160 126 161 
<< m1 >>
rect 127 160 128 161 
<< pdiffusion >>
rect 138 160 139 161 
<< pdiffusion >>
rect 139 160 140 161 
<< pdiffusion >>
rect 140 160 141 161 
<< pdiffusion >>
rect 141 160 142 161 
<< pdiffusion >>
rect 142 160 143 161 
<< pdiffusion >>
rect 143 160 144 161 
<< pdiffusion >>
rect 156 160 157 161 
<< pdiffusion >>
rect 157 160 158 161 
<< pdiffusion >>
rect 158 160 159 161 
<< pdiffusion >>
rect 159 160 160 161 
<< pdiffusion >>
rect 160 160 161 161 
<< pdiffusion >>
rect 161 160 162 161 
<< pdiffusion >>
rect 174 160 175 161 
<< pdiffusion >>
rect 175 160 176 161 
<< pdiffusion >>
rect 176 160 177 161 
<< pdiffusion >>
rect 177 160 178 161 
<< pdiffusion >>
rect 178 160 179 161 
<< pdiffusion >>
rect 179 160 180 161 
<< pdiffusion >>
rect 192 160 193 161 
<< pdiffusion >>
rect 193 160 194 161 
<< pdiffusion >>
rect 194 160 195 161 
<< pdiffusion >>
rect 195 160 196 161 
<< pdiffusion >>
rect 196 160 197 161 
<< pdiffusion >>
rect 197 160 198 161 
<< m1 >>
rect 199 160 200 161 
<< m2 >>
rect 199 160 200 161 
<< pdiffusion >>
rect 210 160 211 161 
<< pdiffusion >>
rect 211 160 212 161 
<< pdiffusion >>
rect 212 160 213 161 
<< pdiffusion >>
rect 213 160 214 161 
<< pdiffusion >>
rect 214 160 215 161 
<< pdiffusion >>
rect 215 160 216 161 
<< m1 >>
rect 217 160 218 161 
<< m1 >>
rect 221 160 222 161 
<< m1 >>
rect 226 160 227 161 
<< pdiffusion >>
rect 228 160 229 161 
<< pdiffusion >>
rect 229 160 230 161 
<< pdiffusion >>
rect 230 160 231 161 
<< pdiffusion >>
rect 231 160 232 161 
<< pdiffusion >>
rect 232 160 233 161 
<< pdiffusion >>
rect 233 160 234 161 
<< m1 >>
rect 235 160 236 161 
<< m1 >>
rect 237 160 238 161 
<< m1 >>
rect 244 160 245 161 
<< pdiffusion >>
rect 246 160 247 161 
<< pdiffusion >>
rect 247 160 248 161 
<< pdiffusion >>
rect 248 160 249 161 
<< pdiffusion >>
rect 249 160 250 161 
<< pdiffusion >>
rect 250 160 251 161 
<< pdiffusion >>
rect 251 160 252 161 
<< m1 >>
rect 253 160 254 161 
<< pdiffusion >>
rect 264 160 265 161 
<< pdiffusion >>
rect 265 160 266 161 
<< pdiffusion >>
rect 266 160 267 161 
<< pdiffusion >>
rect 267 160 268 161 
<< pdiffusion >>
rect 268 160 269 161 
<< pdiffusion >>
rect 269 160 270 161 
<< m1 >>
rect 278 160 279 161 
<< m1 >>
rect 280 160 281 161 
<< m2 >>
rect 280 160 281 161 
<< pdiffusion >>
rect 282 160 283 161 
<< pdiffusion >>
rect 283 160 284 161 
<< pdiffusion >>
rect 284 160 285 161 
<< pdiffusion >>
rect 285 160 286 161 
<< pdiffusion >>
rect 286 160 287 161 
<< pdiffusion >>
rect 287 160 288 161 
<< pdiffusion >>
rect 300 160 301 161 
<< pdiffusion >>
rect 301 160 302 161 
<< pdiffusion >>
rect 302 160 303 161 
<< pdiffusion >>
rect 303 160 304 161 
<< pdiffusion >>
rect 304 160 305 161 
<< pdiffusion >>
rect 305 160 306 161 
<< pdiffusion >>
rect 318 160 319 161 
<< pdiffusion >>
rect 319 160 320 161 
<< pdiffusion >>
rect 320 160 321 161 
<< pdiffusion >>
rect 321 160 322 161 
<< pdiffusion >>
rect 322 160 323 161 
<< pdiffusion >>
rect 323 160 324 161 
<< m1 >>
rect 334 160 335 161 
<< m1 >>
rect 336 160 337 161 
<< m1 >>
rect 343 160 344 161 
<< m1 >>
rect 345 160 346 161 
<< pdiffusion >>
rect 354 160 355 161 
<< pdiffusion >>
rect 355 160 356 161 
<< pdiffusion >>
rect 356 160 357 161 
<< pdiffusion >>
rect 357 160 358 161 
<< pdiffusion >>
rect 358 160 359 161 
<< pdiffusion >>
rect 359 160 360 161 
<< m1 >>
rect 366 160 367 161 
<< m2 >>
rect 369 160 370 161 
<< m1 >>
rect 370 160 371 161 
<< pdiffusion >>
rect 372 160 373 161 
<< pdiffusion >>
rect 373 160 374 161 
<< pdiffusion >>
rect 374 160 375 161 
<< pdiffusion >>
rect 375 160 376 161 
<< pdiffusion >>
rect 376 160 377 161 
<< pdiffusion >>
rect 377 160 378 161 
<< m1 >>
rect 379 160 380 161 
<< m2 >>
rect 379 160 380 161 
<< pdiffusion >>
rect 390 160 391 161 
<< pdiffusion >>
rect 391 160 392 161 
<< pdiffusion >>
rect 392 160 393 161 
<< pdiffusion >>
rect 393 160 394 161 
<< pdiffusion >>
rect 394 160 395 161 
<< pdiffusion >>
rect 395 160 396 161 
<< m1 >>
rect 406 160 407 161 
<< pdiffusion >>
rect 408 160 409 161 
<< pdiffusion >>
rect 409 160 410 161 
<< pdiffusion >>
rect 410 160 411 161 
<< pdiffusion >>
rect 411 160 412 161 
<< pdiffusion >>
rect 412 160 413 161 
<< pdiffusion >>
rect 413 160 414 161 
<< m1 >>
rect 415 160 416 161 
<< m1 >>
rect 417 160 418 161 
<< m1 >>
rect 419 160 420 161 
<< pdiffusion >>
rect 426 160 427 161 
<< pdiffusion >>
rect 427 160 428 161 
<< pdiffusion >>
rect 428 160 429 161 
<< pdiffusion >>
rect 429 160 430 161 
<< pdiffusion >>
rect 430 160 431 161 
<< pdiffusion >>
rect 431 160 432 161 
<< m1 >>
rect 433 160 434 161 
<< m1 >>
rect 442 160 443 161 
<< pdiffusion >>
rect 444 160 445 161 
<< pdiffusion >>
rect 445 160 446 161 
<< pdiffusion >>
rect 446 160 447 161 
<< pdiffusion >>
rect 447 160 448 161 
<< pdiffusion >>
rect 448 160 449 161 
<< pdiffusion >>
rect 449 160 450 161 
<< m1 >>
rect 456 160 457 161 
<< pdiffusion >>
rect 462 160 463 161 
<< pdiffusion >>
rect 463 160 464 161 
<< pdiffusion >>
rect 464 160 465 161 
<< pdiffusion >>
rect 465 160 466 161 
<< pdiffusion >>
rect 466 160 467 161 
<< pdiffusion >>
rect 467 160 468 161 
<< m1 >>
rect 478 160 479 161 
<< pdiffusion >>
rect 480 160 481 161 
<< pdiffusion >>
rect 481 160 482 161 
<< pdiffusion >>
rect 482 160 483 161 
<< pdiffusion >>
rect 483 160 484 161 
<< pdiffusion >>
rect 484 160 485 161 
<< pdiffusion >>
rect 485 160 486 161 
<< pdiffusion >>
rect 498 160 499 161 
<< pdiffusion >>
rect 499 160 500 161 
<< pdiffusion >>
rect 500 160 501 161 
<< pdiffusion >>
rect 501 160 502 161 
<< pdiffusion >>
rect 502 160 503 161 
<< pdiffusion >>
rect 503 160 504 161 
<< pdiffusion >>
rect 516 160 517 161 
<< pdiffusion >>
rect 517 160 518 161 
<< pdiffusion >>
rect 518 160 519 161 
<< pdiffusion >>
rect 519 160 520 161 
<< pdiffusion >>
rect 520 160 521 161 
<< pdiffusion >>
rect 521 160 522 161 
<< pdiffusion >>
rect 12 161 13 162 
<< pdiffusion >>
rect 13 161 14 162 
<< pdiffusion >>
rect 14 161 15 162 
<< pdiffusion >>
rect 15 161 16 162 
<< pdiffusion >>
rect 16 161 17 162 
<< pdiffusion >>
rect 17 161 18 162 
<< pdiffusion >>
rect 30 161 31 162 
<< pdiffusion >>
rect 31 161 32 162 
<< pdiffusion >>
rect 32 161 33 162 
<< pdiffusion >>
rect 33 161 34 162 
<< pdiffusion >>
rect 34 161 35 162 
<< pdiffusion >>
rect 35 161 36 162 
<< m1 >>
rect 37 161 38 162 
<< pdiffusion >>
rect 48 161 49 162 
<< pdiffusion >>
rect 49 161 50 162 
<< pdiffusion >>
rect 50 161 51 162 
<< pdiffusion >>
rect 51 161 52 162 
<< pdiffusion >>
rect 52 161 53 162 
<< pdiffusion >>
rect 53 161 54 162 
<< m1 >>
rect 64 161 65 162 
<< pdiffusion >>
rect 66 161 67 162 
<< pdiffusion >>
rect 67 161 68 162 
<< pdiffusion >>
rect 68 161 69 162 
<< pdiffusion >>
rect 69 161 70 162 
<< pdiffusion >>
rect 70 161 71 162 
<< pdiffusion >>
rect 71 161 72 162 
<< pdiffusion >>
rect 84 161 85 162 
<< pdiffusion >>
rect 85 161 86 162 
<< pdiffusion >>
rect 86 161 87 162 
<< pdiffusion >>
rect 87 161 88 162 
<< pdiffusion >>
rect 88 161 89 162 
<< pdiffusion >>
rect 89 161 90 162 
<< m2 >>
rect 97 161 98 162 
<< m1 >>
rect 98 161 99 162 
<< m1 >>
rect 100 161 101 162 
<< pdiffusion >>
rect 102 161 103 162 
<< pdiffusion >>
rect 103 161 104 162 
<< pdiffusion >>
rect 104 161 105 162 
<< pdiffusion >>
rect 105 161 106 162 
<< pdiffusion >>
rect 106 161 107 162 
<< pdiffusion >>
rect 107 161 108 162 
<< m1 >>
rect 109 161 110 162 
<< m1 >>
rect 114 161 115 162 
<< m1 >>
rect 118 161 119 162 
<< m2 >>
rect 118 161 119 162 
<< pdiffusion >>
rect 120 161 121 162 
<< pdiffusion >>
rect 121 161 122 162 
<< pdiffusion >>
rect 122 161 123 162 
<< pdiffusion >>
rect 123 161 124 162 
<< pdiffusion >>
rect 124 161 125 162 
<< pdiffusion >>
rect 125 161 126 162 
<< m1 >>
rect 127 161 128 162 
<< pdiffusion >>
rect 138 161 139 162 
<< pdiffusion >>
rect 139 161 140 162 
<< pdiffusion >>
rect 140 161 141 162 
<< pdiffusion >>
rect 141 161 142 162 
<< pdiffusion >>
rect 142 161 143 162 
<< pdiffusion >>
rect 143 161 144 162 
<< pdiffusion >>
rect 156 161 157 162 
<< pdiffusion >>
rect 157 161 158 162 
<< pdiffusion >>
rect 158 161 159 162 
<< pdiffusion >>
rect 159 161 160 162 
<< m1 >>
rect 160 161 161 162 
<< pdiffusion >>
rect 160 161 161 162 
<< pdiffusion >>
rect 161 161 162 162 
<< pdiffusion >>
rect 174 161 175 162 
<< m1 >>
rect 175 161 176 162 
<< pdiffusion >>
rect 175 161 176 162 
<< pdiffusion >>
rect 176 161 177 162 
<< pdiffusion >>
rect 177 161 178 162 
<< pdiffusion >>
rect 178 161 179 162 
<< pdiffusion >>
rect 179 161 180 162 
<< pdiffusion >>
rect 192 161 193 162 
<< m1 >>
rect 193 161 194 162 
<< pdiffusion >>
rect 193 161 194 162 
<< pdiffusion >>
rect 194 161 195 162 
<< pdiffusion >>
rect 195 161 196 162 
<< pdiffusion >>
rect 196 161 197 162 
<< pdiffusion >>
rect 197 161 198 162 
<< m1 >>
rect 199 161 200 162 
<< m2 >>
rect 199 161 200 162 
<< pdiffusion >>
rect 210 161 211 162 
<< pdiffusion >>
rect 211 161 212 162 
<< pdiffusion >>
rect 212 161 213 162 
<< pdiffusion >>
rect 213 161 214 162 
<< pdiffusion >>
rect 214 161 215 162 
<< pdiffusion >>
rect 215 161 216 162 
<< m1 >>
rect 217 161 218 162 
<< m1 >>
rect 221 161 222 162 
<< m2 >>
rect 221 161 222 162 
<< m2c >>
rect 221 161 222 162 
<< m1 >>
rect 221 161 222 162 
<< m2 >>
rect 221 161 222 162 
<< m1 >>
rect 226 161 227 162 
<< m2 >>
rect 226 161 227 162 
<< m2c >>
rect 226 161 227 162 
<< m1 >>
rect 226 161 227 162 
<< m2 >>
rect 226 161 227 162 
<< pdiffusion >>
rect 228 161 229 162 
<< m1 >>
rect 229 161 230 162 
<< pdiffusion >>
rect 229 161 230 162 
<< pdiffusion >>
rect 230 161 231 162 
<< pdiffusion >>
rect 231 161 232 162 
<< pdiffusion >>
rect 232 161 233 162 
<< pdiffusion >>
rect 233 161 234 162 
<< m1 >>
rect 235 161 236 162 
<< m1 >>
rect 237 161 238 162 
<< m1 >>
rect 244 161 245 162 
<< m2 >>
rect 244 161 245 162 
<< m2c >>
rect 244 161 245 162 
<< m1 >>
rect 244 161 245 162 
<< m2 >>
rect 244 161 245 162 
<< pdiffusion >>
rect 246 161 247 162 
<< m1 >>
rect 247 161 248 162 
<< pdiffusion >>
rect 247 161 248 162 
<< pdiffusion >>
rect 248 161 249 162 
<< pdiffusion >>
rect 249 161 250 162 
<< pdiffusion >>
rect 250 161 251 162 
<< pdiffusion >>
rect 251 161 252 162 
<< m1 >>
rect 253 161 254 162 
<< pdiffusion >>
rect 264 161 265 162 
<< pdiffusion >>
rect 265 161 266 162 
<< pdiffusion >>
rect 266 161 267 162 
<< pdiffusion >>
rect 267 161 268 162 
<< pdiffusion >>
rect 268 161 269 162 
<< pdiffusion >>
rect 269 161 270 162 
<< m1 >>
rect 278 161 279 162 
<< m1 >>
rect 280 161 281 162 
<< m2 >>
rect 280 161 281 162 
<< pdiffusion >>
rect 282 161 283 162 
<< pdiffusion >>
rect 283 161 284 162 
<< pdiffusion >>
rect 284 161 285 162 
<< pdiffusion >>
rect 285 161 286 162 
<< m1 >>
rect 286 161 287 162 
<< pdiffusion >>
rect 286 161 287 162 
<< pdiffusion >>
rect 287 161 288 162 
<< pdiffusion >>
rect 300 161 301 162 
<< pdiffusion >>
rect 301 161 302 162 
<< pdiffusion >>
rect 302 161 303 162 
<< pdiffusion >>
rect 303 161 304 162 
<< pdiffusion >>
rect 304 161 305 162 
<< pdiffusion >>
rect 305 161 306 162 
<< pdiffusion >>
rect 318 161 319 162 
<< m1 >>
rect 319 161 320 162 
<< pdiffusion >>
rect 319 161 320 162 
<< pdiffusion >>
rect 320 161 321 162 
<< pdiffusion >>
rect 321 161 322 162 
<< pdiffusion >>
rect 322 161 323 162 
<< pdiffusion >>
rect 323 161 324 162 
<< m1 >>
rect 334 161 335 162 
<< m1 >>
rect 336 161 337 162 
<< m1 >>
rect 343 161 344 162 
<< m1 >>
rect 345 161 346 162 
<< pdiffusion >>
rect 354 161 355 162 
<< pdiffusion >>
rect 355 161 356 162 
<< pdiffusion >>
rect 356 161 357 162 
<< pdiffusion >>
rect 357 161 358 162 
<< pdiffusion >>
rect 358 161 359 162 
<< pdiffusion >>
rect 359 161 360 162 
<< m1 >>
rect 366 161 367 162 
<< m2 >>
rect 369 161 370 162 
<< m1 >>
rect 370 161 371 162 
<< pdiffusion >>
rect 372 161 373 162 
<< pdiffusion >>
rect 373 161 374 162 
<< pdiffusion >>
rect 374 161 375 162 
<< pdiffusion >>
rect 375 161 376 162 
<< pdiffusion >>
rect 376 161 377 162 
<< pdiffusion >>
rect 377 161 378 162 
<< m1 >>
rect 379 161 380 162 
<< m2 >>
rect 379 161 380 162 
<< pdiffusion >>
rect 390 161 391 162 
<< m1 >>
rect 391 161 392 162 
<< pdiffusion >>
rect 391 161 392 162 
<< pdiffusion >>
rect 392 161 393 162 
<< pdiffusion >>
rect 393 161 394 162 
<< pdiffusion >>
rect 394 161 395 162 
<< pdiffusion >>
rect 395 161 396 162 
<< m1 >>
rect 406 161 407 162 
<< pdiffusion >>
rect 408 161 409 162 
<< m1 >>
rect 409 161 410 162 
<< pdiffusion >>
rect 409 161 410 162 
<< pdiffusion >>
rect 410 161 411 162 
<< pdiffusion >>
rect 411 161 412 162 
<< m1 >>
rect 412 161 413 162 
<< pdiffusion >>
rect 412 161 413 162 
<< pdiffusion >>
rect 413 161 414 162 
<< m1 >>
rect 415 161 416 162 
<< m1 >>
rect 417 161 418 162 
<< m1 >>
rect 419 161 420 162 
<< pdiffusion >>
rect 426 161 427 162 
<< pdiffusion >>
rect 427 161 428 162 
<< pdiffusion >>
rect 428 161 429 162 
<< pdiffusion >>
rect 429 161 430 162 
<< pdiffusion >>
rect 430 161 431 162 
<< pdiffusion >>
rect 431 161 432 162 
<< m1 >>
rect 433 161 434 162 
<< m1 >>
rect 442 161 443 162 
<< pdiffusion >>
rect 444 161 445 162 
<< pdiffusion >>
rect 445 161 446 162 
<< pdiffusion >>
rect 446 161 447 162 
<< pdiffusion >>
rect 447 161 448 162 
<< m1 >>
rect 448 161 449 162 
<< pdiffusion >>
rect 448 161 449 162 
<< pdiffusion >>
rect 449 161 450 162 
<< m1 >>
rect 456 161 457 162 
<< pdiffusion >>
rect 462 161 463 162 
<< pdiffusion >>
rect 463 161 464 162 
<< pdiffusion >>
rect 464 161 465 162 
<< pdiffusion >>
rect 465 161 466 162 
<< pdiffusion >>
rect 466 161 467 162 
<< pdiffusion >>
rect 467 161 468 162 
<< m1 >>
rect 478 161 479 162 
<< pdiffusion >>
rect 480 161 481 162 
<< pdiffusion >>
rect 481 161 482 162 
<< pdiffusion >>
rect 482 161 483 162 
<< pdiffusion >>
rect 483 161 484 162 
<< pdiffusion >>
rect 484 161 485 162 
<< pdiffusion >>
rect 485 161 486 162 
<< pdiffusion >>
rect 498 161 499 162 
<< pdiffusion >>
rect 499 161 500 162 
<< pdiffusion >>
rect 500 161 501 162 
<< pdiffusion >>
rect 501 161 502 162 
<< pdiffusion >>
rect 502 161 503 162 
<< pdiffusion >>
rect 503 161 504 162 
<< pdiffusion >>
rect 516 161 517 162 
<< pdiffusion >>
rect 517 161 518 162 
<< pdiffusion >>
rect 518 161 519 162 
<< pdiffusion >>
rect 519 161 520 162 
<< pdiffusion >>
rect 520 161 521 162 
<< pdiffusion >>
rect 521 161 522 162 
<< m1 >>
rect 37 162 38 163 
<< m1 >>
rect 64 162 65 163 
<< m2 >>
rect 97 162 98 163 
<< m1 >>
rect 98 162 99 163 
<< m1 >>
rect 100 162 101 163 
<< m1 >>
rect 109 162 110 163 
<< m1 >>
rect 114 162 115 163 
<< m1 >>
rect 118 162 119 163 
<< m2 >>
rect 118 162 119 163 
<< m1 >>
rect 127 162 128 163 
<< m1 >>
rect 160 162 161 163 
<< m1 >>
rect 175 162 176 163 
<< m1 >>
rect 193 162 194 163 
<< m1 >>
rect 199 162 200 163 
<< m2 >>
rect 199 162 200 163 
<< m1 >>
rect 217 162 218 163 
<< m2 >>
rect 221 162 222 163 
<< m2 >>
rect 226 162 227 163 
<< m1 >>
rect 229 162 230 163 
<< m1 >>
rect 235 162 236 163 
<< m1 >>
rect 237 162 238 163 
<< m2 >>
rect 244 162 245 163 
<< m1 >>
rect 247 162 248 163 
<< m1 >>
rect 253 162 254 163 
<< m1 >>
rect 278 162 279 163 
<< m1 >>
rect 280 162 281 163 
<< m2 >>
rect 280 162 281 163 
<< m1 >>
rect 286 162 287 163 
<< m1 >>
rect 319 162 320 163 
<< m1 >>
rect 334 162 335 163 
<< m1 >>
rect 336 162 337 163 
<< m1 >>
rect 343 162 344 163 
<< m1 >>
rect 345 162 346 163 
<< m1 >>
rect 366 162 367 163 
<< m2 >>
rect 369 162 370 163 
<< m1 >>
rect 370 162 371 163 
<< m1 >>
rect 379 162 380 163 
<< m2 >>
rect 379 162 380 163 
<< m1 >>
rect 391 162 392 163 
<< m1 >>
rect 406 162 407 163 
<< m1 >>
rect 409 162 410 163 
<< m1 >>
rect 412 162 413 163 
<< m1 >>
rect 415 162 416 163 
<< m1 >>
rect 417 162 418 163 
<< m1 >>
rect 419 162 420 163 
<< m1 >>
rect 433 162 434 163 
<< m1 >>
rect 442 162 443 163 
<< m1 >>
rect 448 162 449 163 
<< m1 >>
rect 456 162 457 163 
<< m1 >>
rect 478 162 479 163 
<< m1 >>
rect 37 163 38 164 
<< m1 >>
rect 64 163 65 164 
<< m2 >>
rect 97 163 98 164 
<< m1 >>
rect 98 163 99 164 
<< m1 >>
rect 100 163 101 164 
<< m1 >>
rect 109 163 110 164 
<< m1 >>
rect 114 163 115 164 
<< m2 >>
rect 114 163 115 164 
<< m2c >>
rect 114 163 115 164 
<< m1 >>
rect 114 163 115 164 
<< m2 >>
rect 114 163 115 164 
<< m1 >>
rect 118 163 119 164 
<< m2 >>
rect 118 163 119 164 
<< m2 >>
rect 119 163 120 164 
<< m1 >>
rect 120 163 121 164 
<< m2 >>
rect 120 163 121 164 
<< m2c >>
rect 120 163 121 164 
<< m1 >>
rect 120 163 121 164 
<< m2 >>
rect 120 163 121 164 
<< m1 >>
rect 127 163 128 164 
<< m1 >>
rect 160 163 161 164 
<< m1 >>
rect 175 163 176 164 
<< m1 >>
rect 193 163 194 164 
<< m1 >>
rect 199 163 200 164 
<< m2 >>
rect 199 163 200 164 
<< m1 >>
rect 217 163 218 164 
<< m1 >>
rect 218 163 219 164 
<< m1 >>
rect 219 163 220 164 
<< m1 >>
rect 220 163 221 164 
<< m1 >>
rect 221 163 222 164 
<< m2 >>
rect 221 163 222 164 
<< m1 >>
rect 222 163 223 164 
<< m1 >>
rect 223 163 224 164 
<< m1 >>
rect 224 163 225 164 
<< m1 >>
rect 225 163 226 164 
<< m1 >>
rect 226 163 227 164 
<< m2 >>
rect 226 163 227 164 
<< m1 >>
rect 227 163 228 164 
<< m1 >>
rect 228 163 229 164 
<< m1 >>
rect 229 163 230 164 
<< m1 >>
rect 235 163 236 164 
<< m1 >>
rect 237 163 238 164 
<< m1 >>
rect 238 163 239 164 
<< m1 >>
rect 239 163 240 164 
<< m1 >>
rect 240 163 241 164 
<< m1 >>
rect 241 163 242 164 
<< m1 >>
rect 242 163 243 164 
<< m1 >>
rect 243 163 244 164 
<< m1 >>
rect 244 163 245 164 
<< m2 >>
rect 244 163 245 164 
<< m1 >>
rect 245 163 246 164 
<< m1 >>
rect 246 163 247 164 
<< m1 >>
rect 247 163 248 164 
<< m1 >>
rect 253 163 254 164 
<< m1 >>
rect 278 163 279 164 
<< m1 >>
rect 280 163 281 164 
<< m2 >>
rect 280 163 281 164 
<< m1 >>
rect 286 163 287 164 
<< m1 >>
rect 287 163 288 164 
<< m1 >>
rect 288 163 289 164 
<< m1 >>
rect 319 163 320 164 
<< m1 >>
rect 334 163 335 164 
<< m1 >>
rect 336 163 337 164 
<< m1 >>
rect 343 163 344 164 
<< m1 >>
rect 345 163 346 164 
<< m1 >>
rect 366 163 367 164 
<< m2 >>
rect 369 163 370 164 
<< m1 >>
rect 370 163 371 164 
<< m2 >>
rect 370 163 371 164 
<< m2 >>
rect 371 163 372 164 
<< m1 >>
rect 372 163 373 164 
<< m2 >>
rect 372 163 373 164 
<< m2c >>
rect 372 163 373 164 
<< m1 >>
rect 372 163 373 164 
<< m2 >>
rect 372 163 373 164 
<< m1 >>
rect 379 163 380 164 
<< m2 >>
rect 379 163 380 164 
<< m1 >>
rect 380 163 381 164 
<< m1 >>
rect 381 163 382 164 
<< m1 >>
rect 382 163 383 164 
<< m1 >>
rect 383 163 384 164 
<< m1 >>
rect 384 163 385 164 
<< m1 >>
rect 385 163 386 164 
<< m1 >>
rect 386 163 387 164 
<< m1 >>
rect 387 163 388 164 
<< m1 >>
rect 388 163 389 164 
<< m1 >>
rect 389 163 390 164 
<< m1 >>
rect 390 163 391 164 
<< m1 >>
rect 391 163 392 164 
<< m1 >>
rect 402 163 403 164 
<< m1 >>
rect 403 163 404 164 
<< m1 >>
rect 404 163 405 164 
<< m2 >>
rect 404 163 405 164 
<< m2c >>
rect 404 163 405 164 
<< m1 >>
rect 404 163 405 164 
<< m2 >>
rect 404 163 405 164 
<< m2 >>
rect 405 163 406 164 
<< m1 >>
rect 406 163 407 164 
<< m2 >>
rect 406 163 407 164 
<< m2 >>
rect 407 163 408 164 
<< m1 >>
rect 408 163 409 164 
<< m2 >>
rect 408 163 409 164 
<< m2c >>
rect 408 163 409 164 
<< m1 >>
rect 408 163 409 164 
<< m2 >>
rect 408 163 409 164 
<< m1 >>
rect 409 163 410 164 
<< m1 >>
rect 412 163 413 164 
<< m1 >>
rect 415 163 416 164 
<< m1 >>
rect 417 163 418 164 
<< m1 >>
rect 419 163 420 164 
<< m1 >>
rect 420 163 421 164 
<< m1 >>
rect 421 163 422 164 
<< m1 >>
rect 422 163 423 164 
<< m1 >>
rect 423 163 424 164 
<< m1 >>
rect 424 163 425 164 
<< m1 >>
rect 425 163 426 164 
<< m1 >>
rect 433 163 434 164 
<< m1 >>
rect 442 163 443 164 
<< m1 >>
rect 448 163 449 164 
<< m1 >>
rect 456 163 457 164 
<< m1 >>
rect 478 163 479 164 
<< m1 >>
rect 34 164 35 165 
<< m1 >>
rect 35 164 36 165 
<< m1 >>
rect 36 164 37 165 
<< m1 >>
rect 37 164 38 165 
<< m1 >>
rect 64 164 65 165 
<< m2 >>
rect 97 164 98 165 
<< m1 >>
rect 98 164 99 165 
<< m1 >>
rect 100 164 101 165 
<< m1 >>
rect 109 164 110 165 
<< m2 >>
rect 114 164 115 165 
<< m1 >>
rect 118 164 119 165 
<< m1 >>
rect 120 164 121 165 
<< m1 >>
rect 127 164 128 165 
<< m1 >>
rect 160 164 161 165 
<< m1 >>
rect 175 164 176 165 
<< m1 >>
rect 193 164 194 165 
<< m1 >>
rect 199 164 200 165 
<< m2 >>
rect 199 164 200 165 
<< m2 >>
rect 221 164 222 165 
<< m2 >>
rect 226 164 227 165 
<< m1 >>
rect 235 164 236 165 
<< m2 >>
rect 244 164 245 165 
<< m1 >>
rect 253 164 254 165 
<< m1 >>
rect 278 164 279 165 
<< m1 >>
rect 280 164 281 165 
<< m2 >>
rect 280 164 281 165 
<< m1 >>
rect 288 164 289 165 
<< m1 >>
rect 319 164 320 165 
<< m1 >>
rect 322 164 323 165 
<< m1 >>
rect 323 164 324 165 
<< m1 >>
rect 324 164 325 165 
<< m1 >>
rect 325 164 326 165 
<< m1 >>
rect 326 164 327 165 
<< m1 >>
rect 327 164 328 165 
<< m1 >>
rect 328 164 329 165 
<< m1 >>
rect 329 164 330 165 
<< m1 >>
rect 330 164 331 165 
<< m1 >>
rect 331 164 332 165 
<< m1 >>
rect 332 164 333 165 
<< m1 >>
rect 333 164 334 165 
<< m1 >>
rect 334 164 335 165 
<< m1 >>
rect 336 164 337 165 
<< m1 >>
rect 343 164 344 165 
<< m1 >>
rect 345 164 346 165 
<< m1 >>
rect 366 164 367 165 
<< m2 >>
rect 366 164 367 165 
<< m2c >>
rect 366 164 367 165 
<< m1 >>
rect 366 164 367 165 
<< m2 >>
rect 366 164 367 165 
<< m1 >>
rect 370 164 371 165 
<< m1 >>
rect 372 164 373 165 
<< m2 >>
rect 379 164 380 165 
<< m1 >>
rect 402 164 403 165 
<< m1 >>
rect 406 164 407 165 
<< m1 >>
rect 412 164 413 165 
<< m1 >>
rect 415 164 416 165 
<< m1 >>
rect 417 164 418 165 
<< m1 >>
rect 425 164 426 165 
<< m1 >>
rect 433 164 434 165 
<< m1 >>
rect 442 164 443 165 
<< m1 >>
rect 443 164 444 165 
<< m1 >>
rect 444 164 445 165 
<< m2 >>
rect 444 164 445 165 
<< m2c >>
rect 444 164 445 165 
<< m1 >>
rect 444 164 445 165 
<< m2 >>
rect 444 164 445 165 
<< m1 >>
rect 448 164 449 165 
<< m1 >>
rect 456 164 457 165 
<< m1 >>
rect 478 164 479 165 
<< m1 >>
rect 34 165 35 166 
<< m1 >>
rect 64 165 65 166 
<< m2 >>
rect 97 165 98 166 
<< m1 >>
rect 98 165 99 166 
<< m1 >>
rect 100 165 101 166 
<< m1 >>
rect 109 165 110 166 
<< m1 >>
rect 110 165 111 166 
<< m1 >>
rect 111 165 112 166 
<< m1 >>
rect 112 165 113 166 
<< m1 >>
rect 113 165 114 166 
<< m1 >>
rect 114 165 115 166 
<< m2 >>
rect 114 165 115 166 
<< m1 >>
rect 115 165 116 166 
<< m1 >>
rect 116 165 117 166 
<< m2 >>
rect 116 165 117 166 
<< m2c >>
rect 116 165 117 166 
<< m1 >>
rect 116 165 117 166 
<< m2 >>
rect 116 165 117 166 
<< m2 >>
rect 117 165 118 166 
<< m1 >>
rect 118 165 119 166 
<< m1 >>
rect 120 165 121 166 
<< m1 >>
rect 127 165 128 166 
<< m1 >>
rect 160 165 161 166 
<< m1 >>
rect 175 165 176 166 
<< m1 >>
rect 193 165 194 166 
<< m1 >>
rect 199 165 200 166 
<< m2 >>
rect 199 165 200 166 
<< m1 >>
rect 221 165 222 166 
<< m2 >>
rect 221 165 222 166 
<< m2c >>
rect 221 165 222 166 
<< m1 >>
rect 221 165 222 166 
<< m2 >>
rect 221 165 222 166 
<< m1 >>
rect 226 165 227 166 
<< m2 >>
rect 226 165 227 166 
<< m2c >>
rect 226 165 227 166 
<< m1 >>
rect 226 165 227 166 
<< m2 >>
rect 226 165 227 166 
<< m1 >>
rect 235 165 236 166 
<< m1 >>
rect 244 165 245 166 
<< m2 >>
rect 244 165 245 166 
<< m2c >>
rect 244 165 245 166 
<< m1 >>
rect 244 165 245 166 
<< m2 >>
rect 244 165 245 166 
<< m1 >>
rect 253 165 254 166 
<< m1 >>
rect 278 165 279 166 
<< m1 >>
rect 280 165 281 166 
<< m2 >>
rect 280 165 281 166 
<< m1 >>
rect 288 165 289 166 
<< m1 >>
rect 319 165 320 166 
<< m1 >>
rect 322 165 323 166 
<< m1 >>
rect 336 165 337 166 
<< m1 >>
rect 343 165 344 166 
<< m1 >>
rect 345 165 346 166 
<< m2 >>
rect 366 165 367 166 
<< m1 >>
rect 370 165 371 166 
<< m1 >>
rect 372 165 373 166 
<< m1 >>
rect 379 165 380 166 
<< m2 >>
rect 379 165 380 166 
<< m2c >>
rect 379 165 380 166 
<< m1 >>
rect 379 165 380 166 
<< m2 >>
rect 379 165 380 166 
<< m1 >>
rect 380 165 381 166 
<< m1 >>
rect 381 165 382 166 
<< m1 >>
rect 382 165 383 166 
<< m1 >>
rect 383 165 384 166 
<< m1 >>
rect 402 165 403 166 
<< m1 >>
rect 406 165 407 166 
<< m2 >>
rect 411 165 412 166 
<< m1 >>
rect 412 165 413 166 
<< m2 >>
rect 412 165 413 166 
<< m2 >>
rect 413 165 414 166 
<< m2 >>
rect 414 165 415 166 
<< m1 >>
rect 415 165 416 166 
<< m2 >>
rect 415 165 416 166 
<< m2 >>
rect 416 165 417 166 
<< m1 >>
rect 417 165 418 166 
<< m2 >>
rect 417 165 418 166 
<< m2 >>
rect 418 165 419 166 
<< m1 >>
rect 419 165 420 166 
<< m2 >>
rect 419 165 420 166 
<< m2c >>
rect 419 165 420 166 
<< m1 >>
rect 419 165 420 166 
<< m2 >>
rect 419 165 420 166 
<< m1 >>
rect 420 165 421 166 
<< m1 >>
rect 421 165 422 166 
<< m1 >>
rect 422 165 423 166 
<< m1 >>
rect 423 165 424 166 
<< m1 >>
rect 425 165 426 166 
<< m1 >>
rect 433 165 434 166 
<< m2 >>
rect 444 165 445 166 
<< m1 >>
rect 448 165 449 166 
<< m1 >>
rect 456 165 457 166 
<< m2 >>
rect 456 165 457 166 
<< m2c >>
rect 456 165 457 166 
<< m1 >>
rect 456 165 457 166 
<< m2 >>
rect 456 165 457 166 
<< m1 >>
rect 478 165 479 166 
<< m1 >>
rect 34 166 35 167 
<< m1 >>
rect 64 166 65 167 
<< m2 >>
rect 97 166 98 167 
<< m1 >>
rect 98 166 99 167 
<< m1 >>
rect 100 166 101 167 
<< m2 >>
rect 114 166 115 167 
<< m2 >>
rect 117 166 118 167 
<< m1 >>
rect 118 166 119 167 
<< m1 >>
rect 120 166 121 167 
<< m1 >>
rect 121 166 122 167 
<< m1 >>
rect 122 166 123 167 
<< m1 >>
rect 123 166 124 167 
<< m1 >>
rect 124 166 125 167 
<< m1 >>
rect 125 166 126 167 
<< m2 >>
rect 125 166 126 167 
<< m2c >>
rect 125 166 126 167 
<< m1 >>
rect 125 166 126 167 
<< m2 >>
rect 125 166 126 167 
<< m2 >>
rect 126 166 127 167 
<< m1 >>
rect 127 166 128 167 
<< m2 >>
rect 127 166 128 167 
<< m2 >>
rect 128 166 129 167 
<< m1 >>
rect 129 166 130 167 
<< m2 >>
rect 129 166 130 167 
<< m2c >>
rect 129 166 130 167 
<< m1 >>
rect 129 166 130 167 
<< m2 >>
rect 129 166 130 167 
<< m1 >>
rect 160 166 161 167 
<< m1 >>
rect 175 166 176 167 
<< m1 >>
rect 193 166 194 167 
<< m1 >>
rect 199 166 200 167 
<< m2 >>
rect 199 166 200 167 
<< m1 >>
rect 221 166 222 167 
<< m1 >>
rect 226 166 227 167 
<< m1 >>
rect 235 166 236 167 
<< m1 >>
rect 244 166 245 167 
<< m1 >>
rect 253 166 254 167 
<< m1 >>
rect 278 166 279 167 
<< m1 >>
rect 280 166 281 167 
<< m2 >>
rect 280 166 281 167 
<< m1 >>
rect 288 166 289 167 
<< m1 >>
rect 319 166 320 167 
<< m1 >>
rect 322 166 323 167 
<< m1 >>
rect 336 166 337 167 
<< m1 >>
rect 343 166 344 167 
<< m1 >>
rect 345 166 346 167 
<< m1 >>
rect 354 166 355 167 
<< m1 >>
rect 355 166 356 167 
<< m1 >>
rect 356 166 357 167 
<< m1 >>
rect 357 166 358 167 
<< m1 >>
rect 358 166 359 167 
<< m1 >>
rect 359 166 360 167 
<< m1 >>
rect 360 166 361 167 
<< m1 >>
rect 361 166 362 167 
<< m1 >>
rect 362 166 363 167 
<< m1 >>
rect 363 166 364 167 
<< m1 >>
rect 364 166 365 167 
<< m1 >>
rect 365 166 366 167 
<< m1 >>
rect 366 166 367 167 
<< m2 >>
rect 366 166 367 167 
<< m1 >>
rect 367 166 368 167 
<< m1 >>
rect 368 166 369 167 
<< m1 >>
rect 369 166 370 167 
<< m1 >>
rect 370 166 371 167 
<< m1 >>
rect 372 166 373 167 
<< m1 >>
rect 383 166 384 167 
<< m1 >>
rect 402 166 403 167 
<< m1 >>
rect 406 166 407 167 
<< m2 >>
rect 411 166 412 167 
<< m1 >>
rect 412 166 413 167 
<< m1 >>
rect 415 166 416 167 
<< m1 >>
rect 417 166 418 167 
<< m1 >>
rect 423 166 424 167 
<< m1 >>
rect 425 166 426 167 
<< m1 >>
rect 433 166 434 167 
<< m1 >>
rect 434 166 435 167 
<< m1 >>
rect 435 166 436 167 
<< m1 >>
rect 436 166 437 167 
<< m1 >>
rect 437 166 438 167 
<< m1 >>
rect 438 166 439 167 
<< m1 >>
rect 439 166 440 167 
<< m1 >>
rect 440 166 441 167 
<< m1 >>
rect 441 166 442 167 
<< m1 >>
rect 442 166 443 167 
<< m1 >>
rect 443 166 444 167 
<< m1 >>
rect 444 166 445 167 
<< m2 >>
rect 444 166 445 167 
<< m1 >>
rect 445 166 446 167 
<< m1 >>
rect 446 166 447 167 
<< m1 >>
rect 447 166 448 167 
<< m1 >>
rect 448 166 449 167 
<< m2 >>
rect 456 166 457 167 
<< m1 >>
rect 478 166 479 167 
<< m1 >>
rect 34 167 35 168 
<< m1 >>
rect 64 167 65 168 
<< m2 >>
rect 97 167 98 168 
<< m1 >>
rect 98 167 99 168 
<< m1 >>
rect 100 167 101 168 
<< m1 >>
rect 114 167 115 168 
<< m2 >>
rect 114 167 115 168 
<< m2c >>
rect 114 167 115 168 
<< m1 >>
rect 114 167 115 168 
<< m2 >>
rect 114 167 115 168 
<< m2 >>
rect 117 167 118 168 
<< m1 >>
rect 118 167 119 168 
<< m1 >>
rect 127 167 128 168 
<< m1 >>
rect 129 167 130 168 
<< m1 >>
rect 160 167 161 168 
<< m2 >>
rect 160 167 161 168 
<< m2c >>
rect 160 167 161 168 
<< m1 >>
rect 160 167 161 168 
<< m2 >>
rect 160 167 161 168 
<< m1 >>
rect 175 167 176 168 
<< m2 >>
rect 192 167 193 168 
<< m1 >>
rect 193 167 194 168 
<< m2 >>
rect 193 167 194 168 
<< m2 >>
rect 194 167 195 168 
<< m1 >>
rect 195 167 196 168 
<< m2 >>
rect 195 167 196 168 
<< m2c >>
rect 195 167 196 168 
<< m1 >>
rect 195 167 196 168 
<< m2 >>
rect 195 167 196 168 
<< m1 >>
rect 196 167 197 168 
<< m1 >>
rect 197 167 198 168 
<< m1 >>
rect 198 167 199 168 
<< m1 >>
rect 199 167 200 168 
<< m2 >>
rect 199 167 200 168 
<< m1 >>
rect 221 167 222 168 
<< m2 >>
rect 221 167 222 168 
<< m2c >>
rect 221 167 222 168 
<< m1 >>
rect 221 167 222 168 
<< m2 >>
rect 221 167 222 168 
<< m1 >>
rect 226 167 227 168 
<< m2 >>
rect 226 167 227 168 
<< m2c >>
rect 226 167 227 168 
<< m1 >>
rect 226 167 227 168 
<< m2 >>
rect 226 167 227 168 
<< m1 >>
rect 235 167 236 168 
<< m1 >>
rect 244 167 245 168 
<< m1 >>
rect 253 167 254 168 
<< m1 >>
rect 278 167 279 168 
<< m1 >>
rect 280 167 281 168 
<< m2 >>
rect 280 167 281 168 
<< m1 >>
rect 288 167 289 168 
<< m2 >>
rect 288 167 289 168 
<< m2c >>
rect 288 167 289 168 
<< m1 >>
rect 288 167 289 168 
<< m2 >>
rect 288 167 289 168 
<< m1 >>
rect 319 167 320 168 
<< m1 >>
rect 320 167 321 168 
<< m2 >>
rect 320 167 321 168 
<< m2c >>
rect 320 167 321 168 
<< m1 >>
rect 320 167 321 168 
<< m2 >>
rect 320 167 321 168 
<< m2 >>
rect 321 167 322 168 
<< m1 >>
rect 322 167 323 168 
<< m2 >>
rect 322 167 323 168 
<< m2 >>
rect 323 167 324 168 
<< m1 >>
rect 324 167 325 168 
<< m2 >>
rect 324 167 325 168 
<< m2c >>
rect 324 167 325 168 
<< m1 >>
rect 324 167 325 168 
<< m2 >>
rect 324 167 325 168 
<< m1 >>
rect 325 167 326 168 
<< m1 >>
rect 326 167 327 168 
<< m1 >>
rect 327 167 328 168 
<< m1 >>
rect 328 167 329 168 
<< m1 >>
rect 329 167 330 168 
<< m1 >>
rect 330 167 331 168 
<< m1 >>
rect 331 167 332 168 
<< m1 >>
rect 332 167 333 168 
<< m1 >>
rect 333 167 334 168 
<< m1 >>
rect 334 167 335 168 
<< m2 >>
rect 334 167 335 168 
<< m2c >>
rect 334 167 335 168 
<< m1 >>
rect 334 167 335 168 
<< m2 >>
rect 334 167 335 168 
<< m2 >>
rect 335 167 336 168 
<< m1 >>
rect 336 167 337 168 
<< m2 >>
rect 336 167 337 168 
<< m2 >>
rect 337 167 338 168 
<< m1 >>
rect 338 167 339 168 
<< m2 >>
rect 338 167 339 168 
<< m2c >>
rect 338 167 339 168 
<< m1 >>
rect 338 167 339 168 
<< m2 >>
rect 338 167 339 168 
<< m1 >>
rect 339 167 340 168 
<< m1 >>
rect 340 167 341 168 
<< m1 >>
rect 341 167 342 168 
<< m2 >>
rect 341 167 342 168 
<< m2c >>
rect 341 167 342 168 
<< m1 >>
rect 341 167 342 168 
<< m2 >>
rect 341 167 342 168 
<< m2 >>
rect 342 167 343 168 
<< m1 >>
rect 343 167 344 168 
<< m2 >>
rect 343 167 344 168 
<< m2 >>
rect 344 167 345 168 
<< m1 >>
rect 345 167 346 168 
<< m2 >>
rect 345 167 346 168 
<< m2 >>
rect 346 167 347 168 
<< m1 >>
rect 347 167 348 168 
<< m2 >>
rect 347 167 348 168 
<< m2c >>
rect 347 167 348 168 
<< m1 >>
rect 347 167 348 168 
<< m2 >>
rect 347 167 348 168 
<< m1 >>
rect 348 167 349 168 
<< m1 >>
rect 354 167 355 168 
<< m2 >>
rect 366 167 367 168 
<< m1 >>
rect 372 167 373 168 
<< m1 >>
rect 373 167 374 168 
<< m1 >>
rect 374 167 375 168 
<< m1 >>
rect 375 167 376 168 
<< m1 >>
rect 376 167 377 168 
<< m1 >>
rect 377 167 378 168 
<< m1 >>
rect 378 167 379 168 
<< m1 >>
rect 379 167 380 168 
<< m1 >>
rect 380 167 381 168 
<< m1 >>
rect 381 167 382 168 
<< m2 >>
rect 381 167 382 168 
<< m2c >>
rect 381 167 382 168 
<< m1 >>
rect 381 167 382 168 
<< m2 >>
rect 381 167 382 168 
<< m2 >>
rect 382 167 383 168 
<< m1 >>
rect 383 167 384 168 
<< m2 >>
rect 383 167 384 168 
<< m2 >>
rect 384 167 385 168 
<< m1 >>
rect 385 167 386 168 
<< m2 >>
rect 385 167 386 168 
<< m2c >>
rect 385 167 386 168 
<< m1 >>
rect 385 167 386 168 
<< m2 >>
rect 385 167 386 168 
<< m1 >>
rect 386 167 387 168 
<< m1 >>
rect 387 167 388 168 
<< m1 >>
rect 388 167 389 168 
<< m1 >>
rect 389 167 390 168 
<< m1 >>
rect 390 167 391 168 
<< m1 >>
rect 391 167 392 168 
<< m1 >>
rect 392 167 393 168 
<< m1 >>
rect 393 167 394 168 
<< m1 >>
rect 394 167 395 168 
<< m1 >>
rect 395 167 396 168 
<< m1 >>
rect 396 167 397 168 
<< m1 >>
rect 397 167 398 168 
<< m1 >>
rect 398 167 399 168 
<< m1 >>
rect 399 167 400 168 
<< m1 >>
rect 400 167 401 168 
<< m2 >>
rect 400 167 401 168 
<< m2c >>
rect 400 167 401 168 
<< m1 >>
rect 400 167 401 168 
<< m2 >>
rect 400 167 401 168 
<< m2 >>
rect 401 167 402 168 
<< m1 >>
rect 402 167 403 168 
<< m2 >>
rect 402 167 403 168 
<< m2 >>
rect 403 167 404 168 
<< m1 >>
rect 404 167 405 168 
<< m2 >>
rect 404 167 405 168 
<< m2c >>
rect 404 167 405 168 
<< m1 >>
rect 404 167 405 168 
<< m2 >>
rect 404 167 405 168 
<< m2 >>
rect 405 167 406 168 
<< m1 >>
rect 406 167 407 168 
<< m2 >>
rect 406 167 407 168 
<< m2 >>
rect 407 167 408 168 
<< m1 >>
rect 408 167 409 168 
<< m2 >>
rect 408 167 409 168 
<< m2c >>
rect 408 167 409 168 
<< m1 >>
rect 408 167 409 168 
<< m2 >>
rect 408 167 409 168 
<< m1 >>
rect 409 167 410 168 
<< m1 >>
rect 410 167 411 168 
<< m2 >>
rect 410 167 411 168 
<< m2c >>
rect 410 167 411 168 
<< m1 >>
rect 410 167 411 168 
<< m2 >>
rect 410 167 411 168 
<< m2 >>
rect 411 167 412 168 
<< m1 >>
rect 412 167 413 168 
<< m1 >>
rect 413 167 414 168 
<< m2 >>
rect 413 167 414 168 
<< m2c >>
rect 413 167 414 168 
<< m1 >>
rect 413 167 414 168 
<< m2 >>
rect 413 167 414 168 
<< m2 >>
rect 414 167 415 168 
<< m1 >>
rect 415 167 416 168 
<< m2 >>
rect 415 167 416 168 
<< m2 >>
rect 416 167 417 168 
<< m1 >>
rect 417 167 418 168 
<< m2 >>
rect 417 167 418 168 
<< m2 >>
rect 418 167 419 168 
<< m1 >>
rect 423 167 424 168 
<< m1 >>
rect 425 167 426 168 
<< m2 >>
rect 444 167 445 168 
<< m2 >>
rect 445 167 446 168 
<< m2 >>
rect 446 167 447 168 
<< m2 >>
rect 447 167 448 168 
<< m2 >>
rect 448 167 449 168 
<< m2 >>
rect 449 167 450 168 
<< m1 >>
rect 450 167 451 168 
<< m2 >>
rect 450 167 451 168 
<< m2c >>
rect 450 167 451 168 
<< m1 >>
rect 450 167 451 168 
<< m2 >>
rect 450 167 451 168 
<< m1 >>
rect 451 167 452 168 
<< m1 >>
rect 452 167 453 168 
<< m1 >>
rect 453 167 454 168 
<< m1 >>
rect 454 167 455 168 
<< m1 >>
rect 455 167 456 168 
<< m1 >>
rect 456 167 457 168 
<< m2 >>
rect 456 167 457 168 
<< m1 >>
rect 457 167 458 168 
<< m1 >>
rect 458 167 459 168 
<< m1 >>
rect 459 167 460 168 
<< m1 >>
rect 460 167 461 168 
<< m1 >>
rect 461 167 462 168 
<< m1 >>
rect 462 167 463 168 
<< m1 >>
rect 463 167 464 168 
<< m1 >>
rect 478 167 479 168 
<< m1 >>
rect 34 168 35 169 
<< m1 >>
rect 64 168 65 169 
<< m2 >>
rect 97 168 98 169 
<< m1 >>
rect 98 168 99 169 
<< m1 >>
rect 100 168 101 169 
<< m1 >>
rect 114 168 115 169 
<< m2 >>
rect 117 168 118 169 
<< m1 >>
rect 118 168 119 169 
<< m1 >>
rect 127 168 128 169 
<< m1 >>
rect 129 168 130 169 
<< m2 >>
rect 160 168 161 169 
<< m2 >>
rect 161 168 162 169 
<< m2 >>
rect 162 168 163 169 
<< m2 >>
rect 163 168 164 169 
<< m1 >>
rect 175 168 176 169 
<< m2 >>
rect 192 168 193 169 
<< m1 >>
rect 193 168 194 169 
<< m2 >>
rect 199 168 200 169 
<< m2 >>
rect 221 168 222 169 
<< m2 >>
rect 226 168 227 169 
<< m2 >>
rect 231 168 232 169 
<< m2 >>
rect 232 168 233 169 
<< m2 >>
rect 233 168 234 169 
<< m2 >>
rect 234 168 235 169 
<< m1 >>
rect 235 168 236 169 
<< m2 >>
rect 235 168 236 169 
<< m2 >>
rect 236 168 237 169 
<< m1 >>
rect 237 168 238 169 
<< m2 >>
rect 237 168 238 169 
<< m2c >>
rect 237 168 238 169 
<< m1 >>
rect 237 168 238 169 
<< m2 >>
rect 237 168 238 169 
<< m1 >>
rect 238 168 239 169 
<< m1 >>
rect 239 168 240 169 
<< m1 >>
rect 240 168 241 169 
<< m1 >>
rect 241 168 242 169 
<< m1 >>
rect 242 168 243 169 
<< m2 >>
rect 242 168 243 169 
<< m2c >>
rect 242 168 243 169 
<< m1 >>
rect 242 168 243 169 
<< m2 >>
rect 242 168 243 169 
<< m2 >>
rect 243 168 244 169 
<< m1 >>
rect 244 168 245 169 
<< m2 >>
rect 244 168 245 169 
<< m2 >>
rect 245 168 246 169 
<< m1 >>
rect 246 168 247 169 
<< m2 >>
rect 246 168 247 169 
<< m2c >>
rect 246 168 247 169 
<< m1 >>
rect 246 168 247 169 
<< m2 >>
rect 246 168 247 169 
<< m1 >>
rect 247 168 248 169 
<< m1 >>
rect 248 168 249 169 
<< m1 >>
rect 249 168 250 169 
<< m1 >>
rect 250 168 251 169 
<< m1 >>
rect 251 168 252 169 
<< m1 >>
rect 253 168 254 169 
<< m1 >>
rect 278 168 279 169 
<< m1 >>
rect 280 168 281 169 
<< m2 >>
rect 280 168 281 169 
<< m2 >>
rect 288 168 289 169 
<< m2 >>
rect 289 168 290 169 
<< m2 >>
rect 290 168 291 169 
<< m2 >>
rect 291 168 292 169 
<< m2 >>
rect 292 168 293 169 
<< m2 >>
rect 293 168 294 169 
<< m2 >>
rect 294 168 295 169 
<< m2 >>
rect 295 168 296 169 
<< m2 >>
rect 296 168 297 169 
<< m2 >>
rect 297 168 298 169 
<< m2 >>
rect 298 168 299 169 
<< m2 >>
rect 299 168 300 169 
<< m2 >>
rect 300 168 301 169 
<< m2 >>
rect 301 168 302 169 
<< m2 >>
rect 302 168 303 169 
<< m1 >>
rect 322 168 323 169 
<< m1 >>
rect 336 168 337 169 
<< m1 >>
rect 343 168 344 169 
<< m1 >>
rect 345 168 346 169 
<< m1 >>
rect 348 168 349 169 
<< m1 >>
rect 354 168 355 169 
<< m1 >>
rect 366 168 367 169 
<< m2 >>
rect 366 168 367 169 
<< m2c >>
rect 366 168 367 169 
<< m1 >>
rect 366 168 367 169 
<< m2 >>
rect 366 168 367 169 
<< m1 >>
rect 383 168 384 169 
<< m1 >>
rect 402 168 403 169 
<< m1 >>
rect 406 168 407 169 
<< m1 >>
rect 415 168 416 169 
<< m1 >>
rect 417 168 418 169 
<< m2 >>
rect 418 168 419 169 
<< m1 >>
rect 423 168 424 169 
<< m1 >>
rect 425 168 426 169 
<< m1 >>
rect 426 168 427 169 
<< m1 >>
rect 427 168 428 169 
<< m1 >>
rect 428 168 429 169 
<< m1 >>
rect 429 168 430 169 
<< m1 >>
rect 430 168 431 169 
<< m1 >>
rect 431 168 432 169 
<< m1 >>
rect 432 168 433 169 
<< m1 >>
rect 433 168 434 169 
<< m2 >>
rect 456 168 457 169 
<< m1 >>
rect 463 168 464 169 
<< m1 >>
rect 478 168 479 169 
<< m1 >>
rect 34 169 35 170 
<< m1 >>
rect 64 169 65 170 
<< m2 >>
rect 97 169 98 170 
<< m1 >>
rect 98 169 99 170 
<< m1 >>
rect 100 169 101 170 
<< m1 >>
rect 114 169 115 170 
<< m2 >>
rect 117 169 118 170 
<< m1 >>
rect 118 169 119 170 
<< m1 >>
rect 127 169 128 170 
<< m1 >>
rect 129 169 130 170 
<< m1 >>
rect 131 169 132 170 
<< m1 >>
rect 132 169 133 170 
<< m1 >>
rect 133 169 134 170 
<< m1 >>
rect 134 169 135 170 
<< m1 >>
rect 135 169 136 170 
<< m1 >>
rect 136 169 137 170 
<< m1 >>
rect 137 169 138 170 
<< m1 >>
rect 138 169 139 170 
<< m1 >>
rect 139 169 140 170 
<< m1 >>
rect 140 169 141 170 
<< m1 >>
rect 141 169 142 170 
<< m1 >>
rect 142 169 143 170 
<< m1 >>
rect 143 169 144 170 
<< m1 >>
rect 144 169 145 170 
<< m1 >>
rect 145 169 146 170 
<< m1 >>
rect 146 169 147 170 
<< m1 >>
rect 147 169 148 170 
<< m1 >>
rect 148 169 149 170 
<< m1 >>
rect 149 169 150 170 
<< m1 >>
rect 150 169 151 170 
<< m1 >>
rect 151 169 152 170 
<< m1 >>
rect 152 169 153 170 
<< m1 >>
rect 153 169 154 170 
<< m1 >>
rect 154 169 155 170 
<< m1 >>
rect 155 169 156 170 
<< m1 >>
rect 156 169 157 170 
<< m1 >>
rect 157 169 158 170 
<< m1 >>
rect 158 169 159 170 
<< m1 >>
rect 159 169 160 170 
<< m1 >>
rect 160 169 161 170 
<< m1 >>
rect 161 169 162 170 
<< m1 >>
rect 162 169 163 170 
<< m1 >>
rect 163 169 164 170 
<< m2 >>
rect 163 169 164 170 
<< m1 >>
rect 164 169 165 170 
<< m1 >>
rect 165 169 166 170 
<< m1 >>
rect 166 169 167 170 
<< m1 >>
rect 167 169 168 170 
<< m1 >>
rect 168 169 169 170 
<< m1 >>
rect 169 169 170 170 
<< m1 >>
rect 170 169 171 170 
<< m1 >>
rect 171 169 172 170 
<< m1 >>
rect 172 169 173 170 
<< m1 >>
rect 173 169 174 170 
<< m2 >>
rect 173 169 174 170 
<< m2c >>
rect 173 169 174 170 
<< m1 >>
rect 173 169 174 170 
<< m2 >>
rect 173 169 174 170 
<< m2 >>
rect 174 169 175 170 
<< m1 >>
rect 175 169 176 170 
<< m2 >>
rect 175 169 176 170 
<< m1 >>
rect 176 169 177 170 
<< m2 >>
rect 176 169 177 170 
<< m1 >>
rect 177 169 178 170 
<< m2 >>
rect 177 169 178 170 
<< m1 >>
rect 178 169 179 170 
<< m2 >>
rect 178 169 179 170 
<< m1 >>
rect 179 169 180 170 
<< m2 >>
rect 179 169 180 170 
<< m1 >>
rect 180 169 181 170 
<< m2 >>
rect 180 169 181 170 
<< m1 >>
rect 181 169 182 170 
<< m2 >>
rect 181 169 182 170 
<< m1 >>
rect 182 169 183 170 
<< m2 >>
rect 182 169 183 170 
<< m1 >>
rect 183 169 184 170 
<< m2 >>
rect 183 169 184 170 
<< m1 >>
rect 184 169 185 170 
<< m2 >>
rect 184 169 185 170 
<< m1 >>
rect 185 169 186 170 
<< m1 >>
rect 186 169 187 170 
<< m1 >>
rect 187 169 188 170 
<< m1 >>
rect 188 169 189 170 
<< m1 >>
rect 189 169 190 170 
<< m1 >>
rect 190 169 191 170 
<< m2 >>
rect 192 169 193 170 
<< m1 >>
rect 193 169 194 170 
<< m1 >>
rect 194 169 195 170 
<< m1 >>
rect 195 169 196 170 
<< m1 >>
rect 196 169 197 170 
<< m1 >>
rect 197 169 198 170 
<< m1 >>
rect 198 169 199 170 
<< m1 >>
rect 199 169 200 170 
<< m2 >>
rect 199 169 200 170 
<< m1 >>
rect 200 169 201 170 
<< m1 >>
rect 201 169 202 170 
<< m1 >>
rect 202 169 203 170 
<< m1 >>
rect 203 169 204 170 
<< m1 >>
rect 204 169 205 170 
<< m1 >>
rect 205 169 206 170 
<< m1 >>
rect 206 169 207 170 
<< m1 >>
rect 207 169 208 170 
<< m1 >>
rect 208 169 209 170 
<< m1 >>
rect 209 169 210 170 
<< m1 >>
rect 210 169 211 170 
<< m1 >>
rect 211 169 212 170 
<< m1 >>
rect 212 169 213 170 
<< m1 >>
rect 213 169 214 170 
<< m1 >>
rect 214 169 215 170 
<< m1 >>
rect 215 169 216 170 
<< m1 >>
rect 216 169 217 170 
<< m1 >>
rect 217 169 218 170 
<< m1 >>
rect 218 169 219 170 
<< m1 >>
rect 219 169 220 170 
<< m1 >>
rect 220 169 221 170 
<< m1 >>
rect 221 169 222 170 
<< m2 >>
rect 221 169 222 170 
<< m1 >>
rect 222 169 223 170 
<< m1 >>
rect 223 169 224 170 
<< m1 >>
rect 224 169 225 170 
<< m1 >>
rect 225 169 226 170 
<< m1 >>
rect 226 169 227 170 
<< m2 >>
rect 226 169 227 170 
<< m1 >>
rect 227 169 228 170 
<< m1 >>
rect 228 169 229 170 
<< m1 >>
rect 229 169 230 170 
<< m1 >>
rect 230 169 231 170 
<< m1 >>
rect 231 169 232 170 
<< m2 >>
rect 231 169 232 170 
<< m1 >>
rect 232 169 233 170 
<< m1 >>
rect 233 169 234 170 
<< m1 >>
rect 235 169 236 170 
<< m1 >>
rect 244 169 245 170 
<< m1 >>
rect 251 169 252 170 
<< m1 >>
rect 253 169 254 170 
<< m1 >>
rect 278 169 279 170 
<< m1 >>
rect 280 169 281 170 
<< m2 >>
rect 280 169 281 170 
<< m1 >>
rect 286 169 287 170 
<< m2 >>
rect 286 169 287 170 
<< m2c >>
rect 286 169 287 170 
<< m1 >>
rect 286 169 287 170 
<< m2 >>
rect 286 169 287 170 
<< m1 >>
rect 287 169 288 170 
<< m1 >>
rect 288 169 289 170 
<< m1 >>
rect 289 169 290 170 
<< m1 >>
rect 290 169 291 170 
<< m1 >>
rect 291 169 292 170 
<< m1 >>
rect 292 169 293 170 
<< m1 >>
rect 293 169 294 170 
<< m1 >>
rect 294 169 295 170 
<< m1 >>
rect 295 169 296 170 
<< m1 >>
rect 296 169 297 170 
<< m1 >>
rect 297 169 298 170 
<< m1 >>
rect 298 169 299 170 
<< m1 >>
rect 299 169 300 170 
<< m1 >>
rect 300 169 301 170 
<< m1 >>
rect 301 169 302 170 
<< m1 >>
rect 302 169 303 170 
<< m2 >>
rect 302 169 303 170 
<< m1 >>
rect 303 169 304 170 
<< m1 >>
rect 304 169 305 170 
<< m1 >>
rect 305 169 306 170 
<< m1 >>
rect 306 169 307 170 
<< m1 >>
rect 307 169 308 170 
<< m1 >>
rect 308 169 309 170 
<< m1 >>
rect 309 169 310 170 
<< m1 >>
rect 310 169 311 170 
<< m1 >>
rect 311 169 312 170 
<< m1 >>
rect 312 169 313 170 
<< m1 >>
rect 313 169 314 170 
<< m1 >>
rect 314 169 315 170 
<< m1 >>
rect 315 169 316 170 
<< m1 >>
rect 316 169 317 170 
<< m1 >>
rect 317 169 318 170 
<< m1 >>
rect 318 169 319 170 
<< m1 >>
rect 319 169 320 170 
<< m1 >>
rect 320 169 321 170 
<< m2 >>
rect 320 169 321 170 
<< m2c >>
rect 320 169 321 170 
<< m1 >>
rect 320 169 321 170 
<< m2 >>
rect 320 169 321 170 
<< m2 >>
rect 321 169 322 170 
<< m1 >>
rect 322 169 323 170 
<< m2 >>
rect 322 169 323 170 
<< m2 >>
rect 323 169 324 170 
<< m1 >>
rect 324 169 325 170 
<< m2 >>
rect 324 169 325 170 
<< m2c >>
rect 324 169 325 170 
<< m1 >>
rect 324 169 325 170 
<< m2 >>
rect 324 169 325 170 
<< m1 >>
rect 325 169 326 170 
<< m1 >>
rect 326 169 327 170 
<< m1 >>
rect 327 169 328 170 
<< m1 >>
rect 328 169 329 170 
<< m1 >>
rect 329 169 330 170 
<< m1 >>
rect 330 169 331 170 
<< m1 >>
rect 331 169 332 170 
<< m1 >>
rect 332 169 333 170 
<< m1 >>
rect 333 169 334 170 
<< m1 >>
rect 334 169 335 170 
<< m2 >>
rect 334 169 335 170 
<< m2c >>
rect 334 169 335 170 
<< m1 >>
rect 334 169 335 170 
<< m2 >>
rect 334 169 335 170 
<< m2 >>
rect 335 169 336 170 
<< m1 >>
rect 336 169 337 170 
<< m2 >>
rect 336 169 337 170 
<< m2 >>
rect 337 169 338 170 
<< m1 >>
rect 338 169 339 170 
<< m2 >>
rect 338 169 339 170 
<< m2c >>
rect 338 169 339 170 
<< m1 >>
rect 338 169 339 170 
<< m2 >>
rect 338 169 339 170 
<< m1 >>
rect 339 169 340 170 
<< m1 >>
rect 340 169 341 170 
<< m1 >>
rect 341 169 342 170 
<< m2 >>
rect 341 169 342 170 
<< m2c >>
rect 341 169 342 170 
<< m1 >>
rect 341 169 342 170 
<< m2 >>
rect 341 169 342 170 
<< m2 >>
rect 342 169 343 170 
<< m1 >>
rect 343 169 344 170 
<< m2 >>
rect 343 169 344 170 
<< m2 >>
rect 344 169 345 170 
<< m1 >>
rect 345 169 346 170 
<< m2 >>
rect 345 169 346 170 
<< m2c >>
rect 345 169 346 170 
<< m1 >>
rect 345 169 346 170 
<< m2 >>
rect 345 169 346 170 
<< m1 >>
rect 348 169 349 170 
<< m1 >>
rect 354 169 355 170 
<< m1 >>
rect 366 169 367 170 
<< m1 >>
rect 383 169 384 170 
<< m1 >>
rect 402 169 403 170 
<< m1 >>
rect 406 169 407 170 
<< m1 >>
rect 408 169 409 170 
<< m1 >>
rect 409 169 410 170 
<< m1 >>
rect 410 169 411 170 
<< m1 >>
rect 411 169 412 170 
<< m1 >>
rect 412 169 413 170 
<< m1 >>
rect 413 169 414 170 
<< m2 >>
rect 413 169 414 170 
<< m2c >>
rect 413 169 414 170 
<< m1 >>
rect 413 169 414 170 
<< m2 >>
rect 413 169 414 170 
<< m2 >>
rect 414 169 415 170 
<< m1 >>
rect 415 169 416 170 
<< m2 >>
rect 415 169 416 170 
<< m1 >>
rect 417 169 418 170 
<< m2 >>
rect 418 169 419 170 
<< m1 >>
rect 423 169 424 170 
<< m1 >>
rect 433 169 434 170 
<< m1 >>
rect 456 169 457 170 
<< m2 >>
rect 456 169 457 170 
<< m2c >>
rect 456 169 457 170 
<< m1 >>
rect 456 169 457 170 
<< m2 >>
rect 456 169 457 170 
<< m1 >>
rect 463 169 464 170 
<< m1 >>
rect 478 169 479 170 
<< m1 >>
rect 34 170 35 171 
<< m1 >>
rect 64 170 65 171 
<< m2 >>
rect 97 170 98 171 
<< m1 >>
rect 98 170 99 171 
<< m1 >>
rect 100 170 101 171 
<< m1 >>
rect 114 170 115 171 
<< m2 >>
rect 117 170 118 171 
<< m1 >>
rect 118 170 119 171 
<< m1 >>
rect 127 170 128 171 
<< m1 >>
rect 129 170 130 171 
<< m1 >>
rect 131 170 132 171 
<< m2 >>
rect 163 170 164 171 
<< m2 >>
rect 184 170 185 171 
<< m1 >>
rect 190 170 191 171 
<< m2 >>
rect 190 170 191 171 
<< m2c >>
rect 190 170 191 171 
<< m1 >>
rect 190 170 191 171 
<< m2 >>
rect 190 170 191 171 
<< m2 >>
rect 192 170 193 171 
<< m2 >>
rect 199 170 200 171 
<< m2 >>
rect 221 170 222 171 
<< m2 >>
rect 226 170 227 171 
<< m2 >>
rect 231 170 232 171 
<< m1 >>
rect 233 170 234 171 
<< m1 >>
rect 235 170 236 171 
<< m1 >>
rect 244 170 245 171 
<< m2 >>
rect 244 170 245 171 
<< m2c >>
rect 244 170 245 171 
<< m1 >>
rect 244 170 245 171 
<< m2 >>
rect 244 170 245 171 
<< m1 >>
rect 251 170 252 171 
<< m1 >>
rect 253 170 254 171 
<< m1 >>
rect 278 170 279 171 
<< m1 >>
rect 280 170 281 171 
<< m2 >>
rect 280 170 281 171 
<< m2 >>
rect 286 170 287 171 
<< m2 >>
rect 302 170 303 171 
<< m1 >>
rect 322 170 323 171 
<< m1 >>
rect 336 170 337 171 
<< m1 >>
rect 343 170 344 171 
<< m1 >>
rect 348 170 349 171 
<< m1 >>
rect 354 170 355 171 
<< m1 >>
rect 366 170 367 171 
<< m1 >>
rect 383 170 384 171 
<< m2 >>
rect 383 170 384 171 
<< m2c >>
rect 383 170 384 171 
<< m1 >>
rect 383 170 384 171 
<< m2 >>
rect 383 170 384 171 
<< m1 >>
rect 402 170 403 171 
<< m1 >>
rect 406 170 407 171 
<< m1 >>
rect 408 170 409 171 
<< m1 >>
rect 415 170 416 171 
<< m2 >>
rect 415 170 416 171 
<< m1 >>
rect 417 170 418 171 
<< m2 >>
rect 418 170 419 171 
<< m1 >>
rect 423 170 424 171 
<< m1 >>
rect 433 170 434 171 
<< m1 >>
rect 456 170 457 171 
<< m1 >>
rect 463 170 464 171 
<< m1 >>
rect 478 170 479 171 
<< m2 >>
rect 478 170 479 171 
<< m2c >>
rect 478 170 479 171 
<< m1 >>
rect 478 170 479 171 
<< m2 >>
rect 478 170 479 171 
<< m1 >>
rect 34 171 35 172 
<< m1 >>
rect 64 171 65 172 
<< m2 >>
rect 97 171 98 172 
<< m1 >>
rect 98 171 99 172 
<< m1 >>
rect 100 171 101 172 
<< m1 >>
rect 114 171 115 172 
<< m2 >>
rect 117 171 118 172 
<< m1 >>
rect 118 171 119 172 
<< m1 >>
rect 127 171 128 172 
<< m1 >>
rect 129 171 130 172 
<< m1 >>
rect 131 171 132 172 
<< m2 >>
rect 163 171 164 172 
<< m2 >>
rect 184 171 185 172 
<< m2 >>
rect 190 171 191 172 
<< m1 >>
rect 192 171 193 172 
<< m2 >>
rect 192 171 193 172 
<< m2c >>
rect 192 171 193 172 
<< m1 >>
rect 192 171 193 172 
<< m2 >>
rect 192 171 193 172 
<< m2 >>
rect 199 171 200 172 
<< m1 >>
rect 211 171 212 172 
<< m1 >>
rect 212 171 213 172 
<< m1 >>
rect 213 171 214 172 
<< m1 >>
rect 214 171 215 172 
<< m1 >>
rect 215 171 216 172 
<< m1 >>
rect 216 171 217 172 
<< m1 >>
rect 217 171 218 172 
<< m1 >>
rect 221 171 222 172 
<< m2 >>
rect 221 171 222 172 
<< m2c >>
rect 221 171 222 172 
<< m1 >>
rect 221 171 222 172 
<< m2 >>
rect 221 171 222 172 
<< m1 >>
rect 226 171 227 172 
<< m2 >>
rect 226 171 227 172 
<< m2c >>
rect 226 171 227 172 
<< m1 >>
rect 226 171 227 172 
<< m2 >>
rect 226 171 227 172 
<< m1 >>
rect 229 171 230 172 
<< m1 >>
rect 230 171 231 172 
<< m1 >>
rect 231 171 232 172 
<< m2 >>
rect 231 171 232 172 
<< m2c >>
rect 231 171 232 172 
<< m1 >>
rect 231 171 232 172 
<< m2 >>
rect 231 171 232 172 
<< m1 >>
rect 233 171 234 172 
<< m1 >>
rect 235 171 236 172 
<< m2 >>
rect 244 171 245 172 
<< m1 >>
rect 251 171 252 172 
<< m1 >>
rect 253 171 254 172 
<< m1 >>
rect 278 171 279 172 
<< m1 >>
rect 280 171 281 172 
<< m2 >>
rect 280 171 281 172 
<< m1 >>
rect 283 171 284 172 
<< m1 >>
rect 284 171 285 172 
<< m1 >>
rect 285 171 286 172 
<< m1 >>
rect 286 171 287 172 
<< m2 >>
rect 286 171 287 172 
<< m1 >>
rect 287 171 288 172 
<< m1 >>
rect 288 171 289 172 
<< m1 >>
rect 289 171 290 172 
<< m1 >>
rect 302 171 303 172 
<< m2 >>
rect 302 171 303 172 
<< m2c >>
rect 302 171 303 172 
<< m1 >>
rect 302 171 303 172 
<< m2 >>
rect 302 171 303 172 
<< m1 >>
rect 303 171 304 172 
<< m1 >>
rect 304 171 305 172 
<< m1 >>
rect 305 171 306 172 
<< m1 >>
rect 306 171 307 172 
<< m1 >>
rect 307 171 308 172 
<< m2 >>
rect 321 171 322 172 
<< m1 >>
rect 322 171 323 172 
<< m2 >>
rect 322 171 323 172 
<< m2 >>
rect 323 171 324 172 
<< m2 >>
rect 324 171 325 172 
<< m2 >>
rect 325 171 326 172 
<< m1 >>
rect 336 171 337 172 
<< m1 >>
rect 343 171 344 172 
<< m1 >>
rect 348 171 349 172 
<< m1 >>
rect 354 171 355 172 
<< m1 >>
rect 366 171 367 172 
<< m2 >>
rect 383 171 384 172 
<< m1 >>
rect 402 171 403 172 
<< m1 >>
rect 406 171 407 172 
<< m1 >>
rect 408 171 409 172 
<< m1 >>
rect 415 171 416 172 
<< m2 >>
rect 415 171 416 172 
<< m1 >>
rect 417 171 418 172 
<< m2 >>
rect 418 171 419 172 
<< m1 >>
rect 423 171 424 172 
<< m1 >>
rect 433 171 434 172 
<< m1 >>
rect 456 171 457 172 
<< m1 >>
rect 463 171 464 172 
<< m2 >>
rect 478 171 479 172 
<< m1 >>
rect 28 172 29 173 
<< m1 >>
rect 29 172 30 173 
<< m1 >>
rect 30 172 31 173 
<< m1 >>
rect 31 172 32 173 
<< m1 >>
rect 34 172 35 173 
<< m1 >>
rect 64 172 65 173 
<< m2 >>
rect 97 172 98 173 
<< m1 >>
rect 98 172 99 173 
<< m1 >>
rect 100 172 101 173 
<< m1 >>
rect 114 172 115 173 
<< m2 >>
rect 117 172 118 173 
<< m1 >>
rect 118 172 119 173 
<< m1 >>
rect 127 172 128 173 
<< m1 >>
rect 129 172 130 173 
<< m1 >>
rect 131 172 132 173 
<< m1 >>
rect 160 172 161 173 
<< m1 >>
rect 161 172 162 173 
<< m1 >>
rect 162 172 163 173 
<< m1 >>
rect 163 172 164 173 
<< m2 >>
rect 163 172 164 173 
<< m2 >>
rect 184 172 185 173 
<< m1 >>
rect 185 172 186 173 
<< m1 >>
rect 186 172 187 173 
<< m1 >>
rect 187 172 188 173 
<< m1 >>
rect 188 172 189 173 
<< m1 >>
rect 189 172 190 173 
<< m1 >>
rect 190 172 191 173 
<< m2 >>
rect 190 172 191 173 
<< m1 >>
rect 191 172 192 173 
<< m1 >>
rect 192 172 193 173 
<< m1 >>
rect 196 172 197 173 
<< m1 >>
rect 197 172 198 173 
<< m1 >>
rect 198 172 199 173 
<< m1 >>
rect 199 172 200 173 
<< m2 >>
rect 199 172 200 173 
<< m1 >>
rect 211 172 212 173 
<< m1 >>
rect 217 172 218 173 
<< m1 >>
rect 221 172 222 173 
<< m1 >>
rect 226 172 227 173 
<< m1 >>
rect 229 172 230 173 
<< m1 >>
rect 233 172 234 173 
<< m2 >>
rect 233 172 234 173 
<< m2c >>
rect 233 172 234 173 
<< m1 >>
rect 233 172 234 173 
<< m2 >>
rect 233 172 234 173 
<< m2 >>
rect 234 172 235 173 
<< m1 >>
rect 235 172 236 173 
<< m2 >>
rect 235 172 236 173 
<< m2 >>
rect 236 172 237 173 
<< m1 >>
rect 244 172 245 173 
<< m2 >>
rect 244 172 245 173 
<< m1 >>
rect 245 172 246 173 
<< m1 >>
rect 246 172 247 173 
<< m1 >>
rect 247 172 248 173 
<< m1 >>
rect 251 172 252 173 
<< m2 >>
rect 251 172 252 173 
<< m2c >>
rect 251 172 252 173 
<< m1 >>
rect 251 172 252 173 
<< m2 >>
rect 251 172 252 173 
<< m2 >>
rect 252 172 253 173 
<< m1 >>
rect 253 172 254 173 
<< m2 >>
rect 253 172 254 173 
<< m1 >>
rect 278 172 279 173 
<< m1 >>
rect 280 172 281 173 
<< m2 >>
rect 280 172 281 173 
<< m1 >>
rect 283 172 284 173 
<< m2 >>
rect 286 172 287 173 
<< m1 >>
rect 289 172 290 173 
<< m1 >>
rect 307 172 308 173 
<< m1 >>
rect 319 172 320 173 
<< m1 >>
rect 320 172 321 173 
<< m2 >>
rect 320 172 321 173 
<< m2c >>
rect 320 172 321 173 
<< m1 >>
rect 320 172 321 173 
<< m2 >>
rect 320 172 321 173 
<< m2 >>
rect 321 172 322 173 
<< m1 >>
rect 322 172 323 173 
<< m1 >>
rect 325 172 326 173 
<< m2 >>
rect 325 172 326 173 
<< m1 >>
rect 326 172 327 173 
<< m1 >>
rect 327 172 328 173 
<< m1 >>
rect 328 172 329 173 
<< m1 >>
rect 329 172 330 173 
<< m1 >>
rect 330 172 331 173 
<< m1 >>
rect 331 172 332 173 
<< m1 >>
rect 332 172 333 173 
<< m1 >>
rect 333 172 334 173 
<< m1 >>
rect 334 172 335 173 
<< m1 >>
rect 335 172 336 173 
<< m1 >>
rect 336 172 337 173 
<< m1 >>
rect 343 172 344 173 
<< m1 >>
rect 348 172 349 173 
<< m1 >>
rect 354 172 355 173 
<< m1 >>
rect 366 172 367 173 
<< m1 >>
rect 376 172 377 173 
<< m1 >>
rect 377 172 378 173 
<< m1 >>
rect 378 172 379 173 
<< m1 >>
rect 379 172 380 173 
<< m2 >>
rect 380 172 381 173 
<< m1 >>
rect 381 172 382 173 
<< m2 >>
rect 381 172 382 173 
<< m2c >>
rect 381 172 382 173 
<< m1 >>
rect 381 172 382 173 
<< m2 >>
rect 381 172 382 173 
<< m1 >>
rect 382 172 383 173 
<< m1 >>
rect 383 172 384 173 
<< m2 >>
rect 383 172 384 173 
<< m1 >>
rect 384 172 385 173 
<< m1 >>
rect 385 172 386 173 
<< m1 >>
rect 386 172 387 173 
<< m1 >>
rect 387 172 388 173 
<< m1 >>
rect 388 172 389 173 
<< m1 >>
rect 389 172 390 173 
<< m1 >>
rect 390 172 391 173 
<< m1 >>
rect 391 172 392 173 
<< m1 >>
rect 402 172 403 173 
<< m2 >>
rect 405 172 406 173 
<< m1 >>
rect 406 172 407 173 
<< m2 >>
rect 406 172 407 173 
<< m2 >>
rect 407 172 408 173 
<< m1 >>
rect 408 172 409 173 
<< m2 >>
rect 408 172 409 173 
<< m2c >>
rect 408 172 409 173 
<< m1 >>
rect 408 172 409 173 
<< m2 >>
rect 408 172 409 173 
<< m1 >>
rect 415 172 416 173 
<< m2 >>
rect 415 172 416 173 
<< m1 >>
rect 417 172 418 173 
<< m2 >>
rect 418 172 419 173 
<< m1 >>
rect 423 172 424 173 
<< m1 >>
rect 433 172 434 173 
<< m1 >>
rect 456 172 457 173 
<< m1 >>
rect 463 172 464 173 
<< m1 >>
rect 478 172 479 173 
<< m2 >>
rect 478 172 479 173 
<< m1 >>
rect 479 172 480 173 
<< m1 >>
rect 480 172 481 173 
<< m1 >>
rect 481 172 482 173 
<< m1 >>
rect 28 173 29 174 
<< m1 >>
rect 31 173 32 174 
<< m1 >>
rect 34 173 35 174 
<< m1 >>
rect 64 173 65 174 
<< m2 >>
rect 97 173 98 174 
<< m1 >>
rect 98 173 99 174 
<< m1 >>
rect 100 173 101 174 
<< m1 >>
rect 114 173 115 174 
<< m2 >>
rect 117 173 118 174 
<< m1 >>
rect 118 173 119 174 
<< m1 >>
rect 127 173 128 174 
<< m1 >>
rect 129 173 130 174 
<< m1 >>
rect 131 173 132 174 
<< m1 >>
rect 160 173 161 174 
<< m1 >>
rect 163 173 164 174 
<< m2 >>
rect 163 173 164 174 
<< m2 >>
rect 184 173 185 174 
<< m1 >>
rect 185 173 186 174 
<< m2 >>
rect 190 173 191 174 
<< m1 >>
rect 196 173 197 174 
<< m1 >>
rect 199 173 200 174 
<< m2 >>
rect 199 173 200 174 
<< m1 >>
rect 211 173 212 174 
<< m1 >>
rect 217 173 218 174 
<< m1 >>
rect 221 173 222 174 
<< m1 >>
rect 226 173 227 174 
<< m1 >>
rect 229 173 230 174 
<< m1 >>
rect 235 173 236 174 
<< m2 >>
rect 236 173 237 174 
<< m1 >>
rect 244 173 245 174 
<< m2 >>
rect 244 173 245 174 
<< m1 >>
rect 247 173 248 174 
<< m1 >>
rect 253 173 254 174 
<< m2 >>
rect 253 173 254 174 
<< m1 >>
rect 278 173 279 174 
<< m1 >>
rect 280 173 281 174 
<< m2 >>
rect 280 173 281 174 
<< m1 >>
rect 283 173 284 174 
<< m1 >>
rect 286 173 287 174 
<< m2 >>
rect 286 173 287 174 
<< m1 >>
rect 289 173 290 174 
<< m1 >>
rect 307 173 308 174 
<< m1 >>
rect 319 173 320 174 
<< m1 >>
rect 322 173 323 174 
<< m1 >>
rect 325 173 326 174 
<< m2 >>
rect 325 173 326 174 
<< m1 >>
rect 343 173 344 174 
<< m1 >>
rect 348 173 349 174 
<< m1 >>
rect 354 173 355 174 
<< m1 >>
rect 366 173 367 174 
<< m1 >>
rect 376 173 377 174 
<< m1 >>
rect 379 173 380 174 
<< m2 >>
rect 380 173 381 174 
<< m2 >>
rect 383 173 384 174 
<< m1 >>
rect 391 173 392 174 
<< m1 >>
rect 402 173 403 174 
<< m2 >>
rect 405 173 406 174 
<< m1 >>
rect 406 173 407 174 
<< m1 >>
rect 415 173 416 174 
<< m2 >>
rect 415 173 416 174 
<< m1 >>
rect 417 173 418 174 
<< m2 >>
rect 418 173 419 174 
<< m1 >>
rect 423 173 424 174 
<< m1 >>
rect 433 173 434 174 
<< m1 >>
rect 456 173 457 174 
<< m1 >>
rect 463 173 464 174 
<< m1 >>
rect 478 173 479 174 
<< m2 >>
rect 478 173 479 174 
<< m1 >>
rect 481 173 482 174 
<< pdiffusion >>
rect 12 174 13 175 
<< pdiffusion >>
rect 13 174 14 175 
<< pdiffusion >>
rect 14 174 15 175 
<< pdiffusion >>
rect 15 174 16 175 
<< pdiffusion >>
rect 16 174 17 175 
<< pdiffusion >>
rect 17 174 18 175 
<< m1 >>
rect 28 174 29 175 
<< pdiffusion >>
rect 30 174 31 175 
<< m1 >>
rect 31 174 32 175 
<< pdiffusion >>
rect 31 174 32 175 
<< pdiffusion >>
rect 32 174 33 175 
<< pdiffusion >>
rect 33 174 34 175 
<< m1 >>
rect 34 174 35 175 
<< pdiffusion >>
rect 34 174 35 175 
<< pdiffusion >>
rect 35 174 36 175 
<< pdiffusion >>
rect 48 174 49 175 
<< pdiffusion >>
rect 49 174 50 175 
<< pdiffusion >>
rect 50 174 51 175 
<< pdiffusion >>
rect 51 174 52 175 
<< pdiffusion >>
rect 52 174 53 175 
<< pdiffusion >>
rect 53 174 54 175 
<< m1 >>
rect 64 174 65 175 
<< pdiffusion >>
rect 66 174 67 175 
<< pdiffusion >>
rect 67 174 68 175 
<< pdiffusion >>
rect 68 174 69 175 
<< pdiffusion >>
rect 69 174 70 175 
<< pdiffusion >>
rect 70 174 71 175 
<< pdiffusion >>
rect 71 174 72 175 
<< pdiffusion >>
rect 84 174 85 175 
<< pdiffusion >>
rect 85 174 86 175 
<< pdiffusion >>
rect 86 174 87 175 
<< pdiffusion >>
rect 87 174 88 175 
<< pdiffusion >>
rect 88 174 89 175 
<< pdiffusion >>
rect 89 174 90 175 
<< m2 >>
rect 97 174 98 175 
<< m1 >>
rect 98 174 99 175 
<< m1 >>
rect 100 174 101 175 
<< pdiffusion >>
rect 102 174 103 175 
<< pdiffusion >>
rect 103 174 104 175 
<< pdiffusion >>
rect 104 174 105 175 
<< pdiffusion >>
rect 105 174 106 175 
<< pdiffusion >>
rect 106 174 107 175 
<< pdiffusion >>
rect 107 174 108 175 
<< m1 >>
rect 114 174 115 175 
<< m2 >>
rect 117 174 118 175 
<< m1 >>
rect 118 174 119 175 
<< pdiffusion >>
rect 120 174 121 175 
<< pdiffusion >>
rect 121 174 122 175 
<< pdiffusion >>
rect 122 174 123 175 
<< pdiffusion >>
rect 123 174 124 175 
<< pdiffusion >>
rect 124 174 125 175 
<< pdiffusion >>
rect 125 174 126 175 
<< m1 >>
rect 127 174 128 175 
<< m1 >>
rect 129 174 130 175 
<< m1 >>
rect 131 174 132 175 
<< pdiffusion >>
rect 138 174 139 175 
<< pdiffusion >>
rect 139 174 140 175 
<< pdiffusion >>
rect 140 174 141 175 
<< pdiffusion >>
rect 141 174 142 175 
<< pdiffusion >>
rect 142 174 143 175 
<< pdiffusion >>
rect 143 174 144 175 
<< pdiffusion >>
rect 156 174 157 175 
<< pdiffusion >>
rect 157 174 158 175 
<< pdiffusion >>
rect 158 174 159 175 
<< pdiffusion >>
rect 159 174 160 175 
<< m1 >>
rect 160 174 161 175 
<< pdiffusion >>
rect 160 174 161 175 
<< pdiffusion >>
rect 161 174 162 175 
<< m1 >>
rect 163 174 164 175 
<< m2 >>
rect 163 174 164 175 
<< pdiffusion >>
rect 174 174 175 175 
<< pdiffusion >>
rect 175 174 176 175 
<< pdiffusion >>
rect 176 174 177 175 
<< pdiffusion >>
rect 177 174 178 175 
<< pdiffusion >>
rect 178 174 179 175 
<< pdiffusion >>
rect 179 174 180 175 
<< m2 >>
rect 184 174 185 175 
<< m1 >>
rect 185 174 186 175 
<< m2 >>
rect 185 174 186 175 
<< m2 >>
rect 186 174 187 175 
<< m1 >>
rect 187 174 188 175 
<< m2 >>
rect 187 174 188 175 
<< m2c >>
rect 187 174 188 175 
<< m1 >>
rect 187 174 188 175 
<< m2 >>
rect 187 174 188 175 
<< m1 >>
rect 190 174 191 175 
<< m2 >>
rect 190 174 191 175 
<< m2c >>
rect 190 174 191 175 
<< m1 >>
rect 190 174 191 175 
<< m2 >>
rect 190 174 191 175 
<< pdiffusion >>
rect 192 174 193 175 
<< pdiffusion >>
rect 193 174 194 175 
<< pdiffusion >>
rect 194 174 195 175 
<< pdiffusion >>
rect 195 174 196 175 
<< m1 >>
rect 196 174 197 175 
<< pdiffusion >>
rect 196 174 197 175 
<< pdiffusion >>
rect 197 174 198 175 
<< m1 >>
rect 199 174 200 175 
<< m2 >>
rect 199 174 200 175 
<< pdiffusion >>
rect 210 174 211 175 
<< m1 >>
rect 211 174 212 175 
<< pdiffusion >>
rect 211 174 212 175 
<< pdiffusion >>
rect 212 174 213 175 
<< pdiffusion >>
rect 213 174 214 175 
<< pdiffusion >>
rect 214 174 215 175 
<< pdiffusion >>
rect 215 174 216 175 
<< m1 >>
rect 217 174 218 175 
<< m1 >>
rect 221 174 222 175 
<< m1 >>
rect 226 174 227 175 
<< pdiffusion >>
rect 228 174 229 175 
<< m1 >>
rect 229 174 230 175 
<< pdiffusion >>
rect 229 174 230 175 
<< pdiffusion >>
rect 230 174 231 175 
<< pdiffusion >>
rect 231 174 232 175 
<< pdiffusion >>
rect 232 174 233 175 
<< pdiffusion >>
rect 233 174 234 175 
<< m1 >>
rect 235 174 236 175 
<< m2 >>
rect 236 174 237 175 
<< m1 >>
rect 244 174 245 175 
<< m2 >>
rect 244 174 245 175 
<< pdiffusion >>
rect 246 174 247 175 
<< m1 >>
rect 247 174 248 175 
<< pdiffusion >>
rect 247 174 248 175 
<< pdiffusion >>
rect 248 174 249 175 
<< pdiffusion >>
rect 249 174 250 175 
<< pdiffusion >>
rect 250 174 251 175 
<< pdiffusion >>
rect 251 174 252 175 
<< m1 >>
rect 253 174 254 175 
<< m2 >>
rect 253 174 254 175 
<< pdiffusion >>
rect 264 174 265 175 
<< pdiffusion >>
rect 265 174 266 175 
<< pdiffusion >>
rect 266 174 267 175 
<< pdiffusion >>
rect 267 174 268 175 
<< pdiffusion >>
rect 268 174 269 175 
<< pdiffusion >>
rect 269 174 270 175 
<< m1 >>
rect 278 174 279 175 
<< m1 >>
rect 280 174 281 175 
<< m2 >>
rect 280 174 281 175 
<< pdiffusion >>
rect 282 174 283 175 
<< m1 >>
rect 283 174 284 175 
<< pdiffusion >>
rect 283 174 284 175 
<< pdiffusion >>
rect 284 174 285 175 
<< m1 >>
rect 285 174 286 175 
<< m2 >>
rect 285 174 286 175 
<< m2c >>
rect 285 174 286 175 
<< m1 >>
rect 285 174 286 175 
<< m2 >>
rect 285 174 286 175 
<< pdiffusion >>
rect 285 174 286 175 
<< m1 >>
rect 286 174 287 175 
<< pdiffusion >>
rect 286 174 287 175 
<< pdiffusion >>
rect 287 174 288 175 
<< m1 >>
rect 289 174 290 175 
<< pdiffusion >>
rect 300 174 301 175 
<< pdiffusion >>
rect 301 174 302 175 
<< pdiffusion >>
rect 302 174 303 175 
<< pdiffusion >>
rect 303 174 304 175 
<< pdiffusion >>
rect 304 174 305 175 
<< pdiffusion >>
rect 305 174 306 175 
<< m1 >>
rect 307 174 308 175 
<< pdiffusion >>
rect 318 174 319 175 
<< m1 >>
rect 319 174 320 175 
<< pdiffusion >>
rect 319 174 320 175 
<< pdiffusion >>
rect 320 174 321 175 
<< pdiffusion >>
rect 321 174 322 175 
<< m1 >>
rect 322 174 323 175 
<< pdiffusion >>
rect 322 174 323 175 
<< pdiffusion >>
rect 323 174 324 175 
<< m1 >>
rect 325 174 326 175 
<< m2 >>
rect 325 174 326 175 
<< m2 >>
rect 326 174 327 175 
<< m1 >>
rect 327 174 328 175 
<< m2 >>
rect 327 174 328 175 
<< m2c >>
rect 327 174 328 175 
<< m1 >>
rect 327 174 328 175 
<< m2 >>
rect 327 174 328 175 
<< m1 >>
rect 328 174 329 175 
<< m1 >>
rect 329 174 330 175 
<< pdiffusion >>
rect 336 174 337 175 
<< pdiffusion >>
rect 337 174 338 175 
<< pdiffusion >>
rect 338 174 339 175 
<< pdiffusion >>
rect 339 174 340 175 
<< pdiffusion >>
rect 340 174 341 175 
<< pdiffusion >>
rect 341 174 342 175 
<< m1 >>
rect 343 174 344 175 
<< m1 >>
rect 348 174 349 175 
<< m1 >>
rect 354 174 355 175 
<< m1 >>
rect 366 174 367 175 
<< pdiffusion >>
rect 372 174 373 175 
<< pdiffusion >>
rect 373 174 374 175 
<< pdiffusion >>
rect 374 174 375 175 
<< pdiffusion >>
rect 375 174 376 175 
<< m1 >>
rect 376 174 377 175 
<< pdiffusion >>
rect 376 174 377 175 
<< pdiffusion >>
rect 377 174 378 175 
<< m1 >>
rect 379 174 380 175 
<< m2 >>
rect 380 174 381 175 
<< m1 >>
rect 383 174 384 175 
<< m2 >>
rect 383 174 384 175 
<< m2c >>
rect 383 174 384 175 
<< m1 >>
rect 383 174 384 175 
<< m2 >>
rect 383 174 384 175 
<< pdiffusion >>
rect 390 174 391 175 
<< m1 >>
rect 391 174 392 175 
<< pdiffusion >>
rect 391 174 392 175 
<< pdiffusion >>
rect 392 174 393 175 
<< pdiffusion >>
rect 393 174 394 175 
<< pdiffusion >>
rect 394 174 395 175 
<< pdiffusion >>
rect 395 174 396 175 
<< m1 >>
rect 402 174 403 175 
<< m2 >>
rect 405 174 406 175 
<< m1 >>
rect 406 174 407 175 
<< pdiffusion >>
rect 408 174 409 175 
<< pdiffusion >>
rect 409 174 410 175 
<< pdiffusion >>
rect 410 174 411 175 
<< pdiffusion >>
rect 411 174 412 175 
<< pdiffusion >>
rect 412 174 413 175 
<< pdiffusion >>
rect 413 174 414 175 
<< m1 >>
rect 415 174 416 175 
<< m2 >>
rect 415 174 416 175 
<< m1 >>
rect 417 174 418 175 
<< m2 >>
rect 418 174 419 175 
<< m1 >>
rect 423 174 424 175 
<< pdiffusion >>
rect 426 174 427 175 
<< pdiffusion >>
rect 427 174 428 175 
<< pdiffusion >>
rect 428 174 429 175 
<< pdiffusion >>
rect 429 174 430 175 
<< pdiffusion >>
rect 430 174 431 175 
<< pdiffusion >>
rect 431 174 432 175 
<< m1 >>
rect 433 174 434 175 
<< m1 >>
rect 456 174 457 175 
<< pdiffusion >>
rect 462 174 463 175 
<< m1 >>
rect 463 174 464 175 
<< pdiffusion >>
rect 463 174 464 175 
<< pdiffusion >>
rect 464 174 465 175 
<< pdiffusion >>
rect 465 174 466 175 
<< pdiffusion >>
rect 466 174 467 175 
<< pdiffusion >>
rect 467 174 468 175 
<< m1 >>
rect 478 174 479 175 
<< m2 >>
rect 478 174 479 175 
<< pdiffusion >>
rect 480 174 481 175 
<< m1 >>
rect 481 174 482 175 
<< pdiffusion >>
rect 481 174 482 175 
<< pdiffusion >>
rect 482 174 483 175 
<< pdiffusion >>
rect 483 174 484 175 
<< pdiffusion >>
rect 484 174 485 175 
<< pdiffusion >>
rect 485 174 486 175 
<< pdiffusion >>
rect 498 174 499 175 
<< pdiffusion >>
rect 499 174 500 175 
<< pdiffusion >>
rect 500 174 501 175 
<< pdiffusion >>
rect 501 174 502 175 
<< pdiffusion >>
rect 502 174 503 175 
<< pdiffusion >>
rect 503 174 504 175 
<< pdiffusion >>
rect 12 175 13 176 
<< pdiffusion >>
rect 13 175 14 176 
<< pdiffusion >>
rect 14 175 15 176 
<< pdiffusion >>
rect 15 175 16 176 
<< pdiffusion >>
rect 16 175 17 176 
<< pdiffusion >>
rect 17 175 18 176 
<< m1 >>
rect 28 175 29 176 
<< pdiffusion >>
rect 30 175 31 176 
<< pdiffusion >>
rect 31 175 32 176 
<< pdiffusion >>
rect 32 175 33 176 
<< pdiffusion >>
rect 33 175 34 176 
<< pdiffusion >>
rect 34 175 35 176 
<< pdiffusion >>
rect 35 175 36 176 
<< pdiffusion >>
rect 48 175 49 176 
<< pdiffusion >>
rect 49 175 50 176 
<< pdiffusion >>
rect 50 175 51 176 
<< pdiffusion >>
rect 51 175 52 176 
<< pdiffusion >>
rect 52 175 53 176 
<< pdiffusion >>
rect 53 175 54 176 
<< m1 >>
rect 64 175 65 176 
<< pdiffusion >>
rect 66 175 67 176 
<< pdiffusion >>
rect 67 175 68 176 
<< pdiffusion >>
rect 68 175 69 176 
<< pdiffusion >>
rect 69 175 70 176 
<< pdiffusion >>
rect 70 175 71 176 
<< pdiffusion >>
rect 71 175 72 176 
<< pdiffusion >>
rect 84 175 85 176 
<< pdiffusion >>
rect 85 175 86 176 
<< pdiffusion >>
rect 86 175 87 176 
<< pdiffusion >>
rect 87 175 88 176 
<< pdiffusion >>
rect 88 175 89 176 
<< pdiffusion >>
rect 89 175 90 176 
<< m2 >>
rect 97 175 98 176 
<< m1 >>
rect 98 175 99 176 
<< m1 >>
rect 100 175 101 176 
<< pdiffusion >>
rect 102 175 103 176 
<< pdiffusion >>
rect 103 175 104 176 
<< pdiffusion >>
rect 104 175 105 176 
<< pdiffusion >>
rect 105 175 106 176 
<< pdiffusion >>
rect 106 175 107 176 
<< pdiffusion >>
rect 107 175 108 176 
<< m1 >>
rect 114 175 115 176 
<< m2 >>
rect 117 175 118 176 
<< m1 >>
rect 118 175 119 176 
<< pdiffusion >>
rect 120 175 121 176 
<< pdiffusion >>
rect 121 175 122 176 
<< pdiffusion >>
rect 122 175 123 176 
<< pdiffusion >>
rect 123 175 124 176 
<< pdiffusion >>
rect 124 175 125 176 
<< pdiffusion >>
rect 125 175 126 176 
<< m1 >>
rect 127 175 128 176 
<< m1 >>
rect 129 175 130 176 
<< m1 >>
rect 131 175 132 176 
<< pdiffusion >>
rect 138 175 139 176 
<< pdiffusion >>
rect 139 175 140 176 
<< pdiffusion >>
rect 140 175 141 176 
<< pdiffusion >>
rect 141 175 142 176 
<< pdiffusion >>
rect 142 175 143 176 
<< pdiffusion >>
rect 143 175 144 176 
<< pdiffusion >>
rect 156 175 157 176 
<< pdiffusion >>
rect 157 175 158 176 
<< pdiffusion >>
rect 158 175 159 176 
<< pdiffusion >>
rect 159 175 160 176 
<< pdiffusion >>
rect 160 175 161 176 
<< pdiffusion >>
rect 161 175 162 176 
<< m1 >>
rect 163 175 164 176 
<< m2 >>
rect 163 175 164 176 
<< pdiffusion >>
rect 174 175 175 176 
<< pdiffusion >>
rect 175 175 176 176 
<< pdiffusion >>
rect 176 175 177 176 
<< pdiffusion >>
rect 177 175 178 176 
<< pdiffusion >>
rect 178 175 179 176 
<< pdiffusion >>
rect 179 175 180 176 
<< m1 >>
rect 185 175 186 176 
<< m1 >>
rect 187 175 188 176 
<< m1 >>
rect 190 175 191 176 
<< pdiffusion >>
rect 192 175 193 176 
<< pdiffusion >>
rect 193 175 194 176 
<< pdiffusion >>
rect 194 175 195 176 
<< pdiffusion >>
rect 195 175 196 176 
<< pdiffusion >>
rect 196 175 197 176 
<< pdiffusion >>
rect 197 175 198 176 
<< m1 >>
rect 199 175 200 176 
<< m2 >>
rect 199 175 200 176 
<< pdiffusion >>
rect 210 175 211 176 
<< pdiffusion >>
rect 211 175 212 176 
<< pdiffusion >>
rect 212 175 213 176 
<< pdiffusion >>
rect 213 175 214 176 
<< pdiffusion >>
rect 214 175 215 176 
<< pdiffusion >>
rect 215 175 216 176 
<< m1 >>
rect 217 175 218 176 
<< m1 >>
rect 221 175 222 176 
<< m1 >>
rect 226 175 227 176 
<< pdiffusion >>
rect 228 175 229 176 
<< pdiffusion >>
rect 229 175 230 176 
<< pdiffusion >>
rect 230 175 231 176 
<< pdiffusion >>
rect 231 175 232 176 
<< pdiffusion >>
rect 232 175 233 176 
<< pdiffusion >>
rect 233 175 234 176 
<< m1 >>
rect 235 175 236 176 
<< m2 >>
rect 236 175 237 176 
<< m1 >>
rect 244 175 245 176 
<< m2 >>
rect 244 175 245 176 
<< pdiffusion >>
rect 246 175 247 176 
<< pdiffusion >>
rect 247 175 248 176 
<< pdiffusion >>
rect 248 175 249 176 
<< pdiffusion >>
rect 249 175 250 176 
<< pdiffusion >>
rect 250 175 251 176 
<< pdiffusion >>
rect 251 175 252 176 
<< m1 >>
rect 253 175 254 176 
<< m2 >>
rect 253 175 254 176 
<< pdiffusion >>
rect 264 175 265 176 
<< pdiffusion >>
rect 265 175 266 176 
<< pdiffusion >>
rect 266 175 267 176 
<< pdiffusion >>
rect 267 175 268 176 
<< pdiffusion >>
rect 268 175 269 176 
<< pdiffusion >>
rect 269 175 270 176 
<< m1 >>
rect 278 175 279 176 
<< m1 >>
rect 280 175 281 176 
<< m2 >>
rect 280 175 281 176 
<< pdiffusion >>
rect 282 175 283 176 
<< pdiffusion >>
rect 283 175 284 176 
<< pdiffusion >>
rect 284 175 285 176 
<< pdiffusion >>
rect 285 175 286 176 
<< pdiffusion >>
rect 286 175 287 176 
<< pdiffusion >>
rect 287 175 288 176 
<< m1 >>
rect 289 175 290 176 
<< pdiffusion >>
rect 300 175 301 176 
<< pdiffusion >>
rect 301 175 302 176 
<< pdiffusion >>
rect 302 175 303 176 
<< pdiffusion >>
rect 303 175 304 176 
<< pdiffusion >>
rect 304 175 305 176 
<< pdiffusion >>
rect 305 175 306 176 
<< m1 >>
rect 307 175 308 176 
<< pdiffusion >>
rect 318 175 319 176 
<< pdiffusion >>
rect 319 175 320 176 
<< pdiffusion >>
rect 320 175 321 176 
<< pdiffusion >>
rect 321 175 322 176 
<< pdiffusion >>
rect 322 175 323 176 
<< pdiffusion >>
rect 323 175 324 176 
<< m1 >>
rect 325 175 326 176 
<< m1 >>
rect 329 175 330 176 
<< pdiffusion >>
rect 336 175 337 176 
<< pdiffusion >>
rect 337 175 338 176 
<< pdiffusion >>
rect 338 175 339 176 
<< pdiffusion >>
rect 339 175 340 176 
<< pdiffusion >>
rect 340 175 341 176 
<< pdiffusion >>
rect 341 175 342 176 
<< m1 >>
rect 343 175 344 176 
<< m1 >>
rect 348 175 349 176 
<< m1 >>
rect 354 175 355 176 
<< m1 >>
rect 366 175 367 176 
<< pdiffusion >>
rect 372 175 373 176 
<< pdiffusion >>
rect 373 175 374 176 
<< pdiffusion >>
rect 374 175 375 176 
<< pdiffusion >>
rect 375 175 376 176 
<< pdiffusion >>
rect 376 175 377 176 
<< pdiffusion >>
rect 377 175 378 176 
<< m1 >>
rect 379 175 380 176 
<< m2 >>
rect 380 175 381 176 
<< m1 >>
rect 383 175 384 176 
<< pdiffusion >>
rect 390 175 391 176 
<< pdiffusion >>
rect 391 175 392 176 
<< pdiffusion >>
rect 392 175 393 176 
<< pdiffusion >>
rect 393 175 394 176 
<< pdiffusion >>
rect 394 175 395 176 
<< pdiffusion >>
rect 395 175 396 176 
<< m1 >>
rect 402 175 403 176 
<< m2 >>
rect 405 175 406 176 
<< m1 >>
rect 406 175 407 176 
<< pdiffusion >>
rect 408 175 409 176 
<< pdiffusion >>
rect 409 175 410 176 
<< pdiffusion >>
rect 410 175 411 176 
<< pdiffusion >>
rect 411 175 412 176 
<< pdiffusion >>
rect 412 175 413 176 
<< pdiffusion >>
rect 413 175 414 176 
<< m1 >>
rect 415 175 416 176 
<< m2 >>
rect 415 175 416 176 
<< m1 >>
rect 417 175 418 176 
<< m2 >>
rect 418 175 419 176 
<< m1 >>
rect 423 175 424 176 
<< pdiffusion >>
rect 426 175 427 176 
<< pdiffusion >>
rect 427 175 428 176 
<< pdiffusion >>
rect 428 175 429 176 
<< pdiffusion >>
rect 429 175 430 176 
<< pdiffusion >>
rect 430 175 431 176 
<< pdiffusion >>
rect 431 175 432 176 
<< m1 >>
rect 433 175 434 176 
<< m1 >>
rect 456 175 457 176 
<< pdiffusion >>
rect 462 175 463 176 
<< pdiffusion >>
rect 463 175 464 176 
<< pdiffusion >>
rect 464 175 465 176 
<< pdiffusion >>
rect 465 175 466 176 
<< pdiffusion >>
rect 466 175 467 176 
<< pdiffusion >>
rect 467 175 468 176 
<< m1 >>
rect 478 175 479 176 
<< m2 >>
rect 478 175 479 176 
<< pdiffusion >>
rect 480 175 481 176 
<< pdiffusion >>
rect 481 175 482 176 
<< pdiffusion >>
rect 482 175 483 176 
<< pdiffusion >>
rect 483 175 484 176 
<< pdiffusion >>
rect 484 175 485 176 
<< pdiffusion >>
rect 485 175 486 176 
<< pdiffusion >>
rect 498 175 499 176 
<< pdiffusion >>
rect 499 175 500 176 
<< pdiffusion >>
rect 500 175 501 176 
<< pdiffusion >>
rect 501 175 502 176 
<< pdiffusion >>
rect 502 175 503 176 
<< pdiffusion >>
rect 503 175 504 176 
<< pdiffusion >>
rect 12 176 13 177 
<< pdiffusion >>
rect 13 176 14 177 
<< pdiffusion >>
rect 14 176 15 177 
<< pdiffusion >>
rect 15 176 16 177 
<< pdiffusion >>
rect 16 176 17 177 
<< pdiffusion >>
rect 17 176 18 177 
<< m1 >>
rect 28 176 29 177 
<< pdiffusion >>
rect 30 176 31 177 
<< pdiffusion >>
rect 31 176 32 177 
<< pdiffusion >>
rect 32 176 33 177 
<< pdiffusion >>
rect 33 176 34 177 
<< pdiffusion >>
rect 34 176 35 177 
<< pdiffusion >>
rect 35 176 36 177 
<< pdiffusion >>
rect 48 176 49 177 
<< pdiffusion >>
rect 49 176 50 177 
<< pdiffusion >>
rect 50 176 51 177 
<< pdiffusion >>
rect 51 176 52 177 
<< pdiffusion >>
rect 52 176 53 177 
<< pdiffusion >>
rect 53 176 54 177 
<< m1 >>
rect 64 176 65 177 
<< pdiffusion >>
rect 66 176 67 177 
<< pdiffusion >>
rect 67 176 68 177 
<< pdiffusion >>
rect 68 176 69 177 
<< pdiffusion >>
rect 69 176 70 177 
<< pdiffusion >>
rect 70 176 71 177 
<< pdiffusion >>
rect 71 176 72 177 
<< pdiffusion >>
rect 84 176 85 177 
<< pdiffusion >>
rect 85 176 86 177 
<< pdiffusion >>
rect 86 176 87 177 
<< pdiffusion >>
rect 87 176 88 177 
<< pdiffusion >>
rect 88 176 89 177 
<< pdiffusion >>
rect 89 176 90 177 
<< m2 >>
rect 97 176 98 177 
<< m1 >>
rect 98 176 99 177 
<< m1 >>
rect 100 176 101 177 
<< pdiffusion >>
rect 102 176 103 177 
<< pdiffusion >>
rect 103 176 104 177 
<< pdiffusion >>
rect 104 176 105 177 
<< pdiffusion >>
rect 105 176 106 177 
<< pdiffusion >>
rect 106 176 107 177 
<< pdiffusion >>
rect 107 176 108 177 
<< m1 >>
rect 114 176 115 177 
<< m2 >>
rect 117 176 118 177 
<< m1 >>
rect 118 176 119 177 
<< pdiffusion >>
rect 120 176 121 177 
<< pdiffusion >>
rect 121 176 122 177 
<< pdiffusion >>
rect 122 176 123 177 
<< pdiffusion >>
rect 123 176 124 177 
<< pdiffusion >>
rect 124 176 125 177 
<< pdiffusion >>
rect 125 176 126 177 
<< m1 >>
rect 127 176 128 177 
<< m1 >>
rect 129 176 130 177 
<< m1 >>
rect 131 176 132 177 
<< pdiffusion >>
rect 138 176 139 177 
<< pdiffusion >>
rect 139 176 140 177 
<< pdiffusion >>
rect 140 176 141 177 
<< pdiffusion >>
rect 141 176 142 177 
<< pdiffusion >>
rect 142 176 143 177 
<< pdiffusion >>
rect 143 176 144 177 
<< pdiffusion >>
rect 156 176 157 177 
<< pdiffusion >>
rect 157 176 158 177 
<< pdiffusion >>
rect 158 176 159 177 
<< pdiffusion >>
rect 159 176 160 177 
<< pdiffusion >>
rect 160 176 161 177 
<< pdiffusion >>
rect 161 176 162 177 
<< m1 >>
rect 163 176 164 177 
<< m2 >>
rect 163 176 164 177 
<< pdiffusion >>
rect 174 176 175 177 
<< pdiffusion >>
rect 175 176 176 177 
<< pdiffusion >>
rect 176 176 177 177 
<< pdiffusion >>
rect 177 176 178 177 
<< pdiffusion >>
rect 178 176 179 177 
<< pdiffusion >>
rect 179 176 180 177 
<< m1 >>
rect 185 176 186 177 
<< m1 >>
rect 187 176 188 177 
<< m1 >>
rect 188 176 189 177 
<< m2 >>
rect 188 176 189 177 
<< m2c >>
rect 188 176 189 177 
<< m1 >>
rect 188 176 189 177 
<< m2 >>
rect 188 176 189 177 
<< m2 >>
rect 189 176 190 177 
<< m1 >>
rect 190 176 191 177 
<< pdiffusion >>
rect 192 176 193 177 
<< pdiffusion >>
rect 193 176 194 177 
<< pdiffusion >>
rect 194 176 195 177 
<< pdiffusion >>
rect 195 176 196 177 
<< pdiffusion >>
rect 196 176 197 177 
<< pdiffusion >>
rect 197 176 198 177 
<< m1 >>
rect 199 176 200 177 
<< m2 >>
rect 199 176 200 177 
<< pdiffusion >>
rect 210 176 211 177 
<< pdiffusion >>
rect 211 176 212 177 
<< pdiffusion >>
rect 212 176 213 177 
<< pdiffusion >>
rect 213 176 214 177 
<< pdiffusion >>
rect 214 176 215 177 
<< pdiffusion >>
rect 215 176 216 177 
<< m1 >>
rect 217 176 218 177 
<< m1 >>
rect 221 176 222 177 
<< m1 >>
rect 226 176 227 177 
<< pdiffusion >>
rect 228 176 229 177 
<< pdiffusion >>
rect 229 176 230 177 
<< pdiffusion >>
rect 230 176 231 177 
<< pdiffusion >>
rect 231 176 232 177 
<< pdiffusion >>
rect 232 176 233 177 
<< pdiffusion >>
rect 233 176 234 177 
<< m1 >>
rect 235 176 236 177 
<< m2 >>
rect 236 176 237 177 
<< m1 >>
rect 244 176 245 177 
<< m2 >>
rect 244 176 245 177 
<< pdiffusion >>
rect 246 176 247 177 
<< pdiffusion >>
rect 247 176 248 177 
<< pdiffusion >>
rect 248 176 249 177 
<< pdiffusion >>
rect 249 176 250 177 
<< pdiffusion >>
rect 250 176 251 177 
<< pdiffusion >>
rect 251 176 252 177 
<< m1 >>
rect 253 176 254 177 
<< m2 >>
rect 253 176 254 177 
<< pdiffusion >>
rect 264 176 265 177 
<< pdiffusion >>
rect 265 176 266 177 
<< pdiffusion >>
rect 266 176 267 177 
<< pdiffusion >>
rect 267 176 268 177 
<< pdiffusion >>
rect 268 176 269 177 
<< pdiffusion >>
rect 269 176 270 177 
<< m1 >>
rect 278 176 279 177 
<< m1 >>
rect 280 176 281 177 
<< m2 >>
rect 280 176 281 177 
<< pdiffusion >>
rect 282 176 283 177 
<< pdiffusion >>
rect 283 176 284 177 
<< pdiffusion >>
rect 284 176 285 177 
<< pdiffusion >>
rect 285 176 286 177 
<< pdiffusion >>
rect 286 176 287 177 
<< pdiffusion >>
rect 287 176 288 177 
<< m1 >>
rect 289 176 290 177 
<< pdiffusion >>
rect 300 176 301 177 
<< pdiffusion >>
rect 301 176 302 177 
<< pdiffusion >>
rect 302 176 303 177 
<< pdiffusion >>
rect 303 176 304 177 
<< pdiffusion >>
rect 304 176 305 177 
<< pdiffusion >>
rect 305 176 306 177 
<< m1 >>
rect 307 176 308 177 
<< pdiffusion >>
rect 318 176 319 177 
<< pdiffusion >>
rect 319 176 320 177 
<< pdiffusion >>
rect 320 176 321 177 
<< pdiffusion >>
rect 321 176 322 177 
<< pdiffusion >>
rect 322 176 323 177 
<< pdiffusion >>
rect 323 176 324 177 
<< m1 >>
rect 325 176 326 177 
<< m1 >>
rect 329 176 330 177 
<< pdiffusion >>
rect 336 176 337 177 
<< pdiffusion >>
rect 337 176 338 177 
<< pdiffusion >>
rect 338 176 339 177 
<< pdiffusion >>
rect 339 176 340 177 
<< pdiffusion >>
rect 340 176 341 177 
<< pdiffusion >>
rect 341 176 342 177 
<< m1 >>
rect 343 176 344 177 
<< m1 >>
rect 348 176 349 177 
<< m1 >>
rect 354 176 355 177 
<< m1 >>
rect 366 176 367 177 
<< pdiffusion >>
rect 372 176 373 177 
<< pdiffusion >>
rect 373 176 374 177 
<< pdiffusion >>
rect 374 176 375 177 
<< pdiffusion >>
rect 375 176 376 177 
<< pdiffusion >>
rect 376 176 377 177 
<< pdiffusion >>
rect 377 176 378 177 
<< m1 >>
rect 379 176 380 177 
<< m2 >>
rect 380 176 381 177 
<< m1 >>
rect 383 176 384 177 
<< pdiffusion >>
rect 390 176 391 177 
<< pdiffusion >>
rect 391 176 392 177 
<< pdiffusion >>
rect 392 176 393 177 
<< pdiffusion >>
rect 393 176 394 177 
<< pdiffusion >>
rect 394 176 395 177 
<< pdiffusion >>
rect 395 176 396 177 
<< m1 >>
rect 402 176 403 177 
<< m2 >>
rect 405 176 406 177 
<< m1 >>
rect 406 176 407 177 
<< pdiffusion >>
rect 408 176 409 177 
<< pdiffusion >>
rect 409 176 410 177 
<< pdiffusion >>
rect 410 176 411 177 
<< pdiffusion >>
rect 411 176 412 177 
<< pdiffusion >>
rect 412 176 413 177 
<< pdiffusion >>
rect 413 176 414 177 
<< m1 >>
rect 415 176 416 177 
<< m2 >>
rect 415 176 416 177 
<< m1 >>
rect 417 176 418 177 
<< m2 >>
rect 418 176 419 177 
<< m1 >>
rect 423 176 424 177 
<< pdiffusion >>
rect 426 176 427 177 
<< pdiffusion >>
rect 427 176 428 177 
<< pdiffusion >>
rect 428 176 429 177 
<< pdiffusion >>
rect 429 176 430 177 
<< pdiffusion >>
rect 430 176 431 177 
<< pdiffusion >>
rect 431 176 432 177 
<< m1 >>
rect 433 176 434 177 
<< m1 >>
rect 456 176 457 177 
<< pdiffusion >>
rect 462 176 463 177 
<< pdiffusion >>
rect 463 176 464 177 
<< pdiffusion >>
rect 464 176 465 177 
<< pdiffusion >>
rect 465 176 466 177 
<< pdiffusion >>
rect 466 176 467 177 
<< pdiffusion >>
rect 467 176 468 177 
<< m1 >>
rect 478 176 479 177 
<< m2 >>
rect 478 176 479 177 
<< pdiffusion >>
rect 480 176 481 177 
<< pdiffusion >>
rect 481 176 482 177 
<< pdiffusion >>
rect 482 176 483 177 
<< pdiffusion >>
rect 483 176 484 177 
<< pdiffusion >>
rect 484 176 485 177 
<< pdiffusion >>
rect 485 176 486 177 
<< pdiffusion >>
rect 498 176 499 177 
<< pdiffusion >>
rect 499 176 500 177 
<< pdiffusion >>
rect 500 176 501 177 
<< pdiffusion >>
rect 501 176 502 177 
<< pdiffusion >>
rect 502 176 503 177 
<< pdiffusion >>
rect 503 176 504 177 
<< pdiffusion >>
rect 12 177 13 178 
<< pdiffusion >>
rect 13 177 14 178 
<< pdiffusion >>
rect 14 177 15 178 
<< pdiffusion >>
rect 15 177 16 178 
<< pdiffusion >>
rect 16 177 17 178 
<< pdiffusion >>
rect 17 177 18 178 
<< m1 >>
rect 28 177 29 178 
<< pdiffusion >>
rect 30 177 31 178 
<< pdiffusion >>
rect 31 177 32 178 
<< pdiffusion >>
rect 32 177 33 178 
<< pdiffusion >>
rect 33 177 34 178 
<< pdiffusion >>
rect 34 177 35 178 
<< pdiffusion >>
rect 35 177 36 178 
<< pdiffusion >>
rect 48 177 49 178 
<< pdiffusion >>
rect 49 177 50 178 
<< pdiffusion >>
rect 50 177 51 178 
<< pdiffusion >>
rect 51 177 52 178 
<< pdiffusion >>
rect 52 177 53 178 
<< pdiffusion >>
rect 53 177 54 178 
<< m1 >>
rect 64 177 65 178 
<< pdiffusion >>
rect 66 177 67 178 
<< pdiffusion >>
rect 67 177 68 178 
<< pdiffusion >>
rect 68 177 69 178 
<< pdiffusion >>
rect 69 177 70 178 
<< pdiffusion >>
rect 70 177 71 178 
<< pdiffusion >>
rect 71 177 72 178 
<< pdiffusion >>
rect 84 177 85 178 
<< pdiffusion >>
rect 85 177 86 178 
<< pdiffusion >>
rect 86 177 87 178 
<< pdiffusion >>
rect 87 177 88 178 
<< pdiffusion >>
rect 88 177 89 178 
<< pdiffusion >>
rect 89 177 90 178 
<< m2 >>
rect 97 177 98 178 
<< m1 >>
rect 98 177 99 178 
<< m1 >>
rect 100 177 101 178 
<< pdiffusion >>
rect 102 177 103 178 
<< pdiffusion >>
rect 103 177 104 178 
<< pdiffusion >>
rect 104 177 105 178 
<< pdiffusion >>
rect 105 177 106 178 
<< pdiffusion >>
rect 106 177 107 178 
<< pdiffusion >>
rect 107 177 108 178 
<< m1 >>
rect 114 177 115 178 
<< m2 >>
rect 117 177 118 178 
<< m1 >>
rect 118 177 119 178 
<< pdiffusion >>
rect 120 177 121 178 
<< pdiffusion >>
rect 121 177 122 178 
<< pdiffusion >>
rect 122 177 123 178 
<< pdiffusion >>
rect 123 177 124 178 
<< pdiffusion >>
rect 124 177 125 178 
<< pdiffusion >>
rect 125 177 126 178 
<< m1 >>
rect 127 177 128 178 
<< m1 >>
rect 129 177 130 178 
<< m1 >>
rect 131 177 132 178 
<< pdiffusion >>
rect 138 177 139 178 
<< pdiffusion >>
rect 139 177 140 178 
<< pdiffusion >>
rect 140 177 141 178 
<< pdiffusion >>
rect 141 177 142 178 
<< pdiffusion >>
rect 142 177 143 178 
<< pdiffusion >>
rect 143 177 144 178 
<< pdiffusion >>
rect 156 177 157 178 
<< pdiffusion >>
rect 157 177 158 178 
<< pdiffusion >>
rect 158 177 159 178 
<< pdiffusion >>
rect 159 177 160 178 
<< pdiffusion >>
rect 160 177 161 178 
<< pdiffusion >>
rect 161 177 162 178 
<< m1 >>
rect 163 177 164 178 
<< m2 >>
rect 163 177 164 178 
<< pdiffusion >>
rect 174 177 175 178 
<< pdiffusion >>
rect 175 177 176 178 
<< pdiffusion >>
rect 176 177 177 178 
<< pdiffusion >>
rect 177 177 178 178 
<< pdiffusion >>
rect 178 177 179 178 
<< pdiffusion >>
rect 179 177 180 178 
<< m1 >>
rect 185 177 186 178 
<< m2 >>
rect 189 177 190 178 
<< m1 >>
rect 190 177 191 178 
<< pdiffusion >>
rect 192 177 193 178 
<< pdiffusion >>
rect 193 177 194 178 
<< pdiffusion >>
rect 194 177 195 178 
<< pdiffusion >>
rect 195 177 196 178 
<< pdiffusion >>
rect 196 177 197 178 
<< pdiffusion >>
rect 197 177 198 178 
<< m1 >>
rect 199 177 200 178 
<< m2 >>
rect 199 177 200 178 
<< pdiffusion >>
rect 210 177 211 178 
<< pdiffusion >>
rect 211 177 212 178 
<< pdiffusion >>
rect 212 177 213 178 
<< pdiffusion >>
rect 213 177 214 178 
<< pdiffusion >>
rect 214 177 215 178 
<< pdiffusion >>
rect 215 177 216 178 
<< m1 >>
rect 217 177 218 178 
<< m1 >>
rect 221 177 222 178 
<< m1 >>
rect 226 177 227 178 
<< pdiffusion >>
rect 228 177 229 178 
<< pdiffusion >>
rect 229 177 230 178 
<< pdiffusion >>
rect 230 177 231 178 
<< pdiffusion >>
rect 231 177 232 178 
<< pdiffusion >>
rect 232 177 233 178 
<< pdiffusion >>
rect 233 177 234 178 
<< m1 >>
rect 235 177 236 178 
<< m2 >>
rect 236 177 237 178 
<< m1 >>
rect 244 177 245 178 
<< m2 >>
rect 244 177 245 178 
<< pdiffusion >>
rect 246 177 247 178 
<< pdiffusion >>
rect 247 177 248 178 
<< pdiffusion >>
rect 248 177 249 178 
<< pdiffusion >>
rect 249 177 250 178 
<< pdiffusion >>
rect 250 177 251 178 
<< pdiffusion >>
rect 251 177 252 178 
<< m1 >>
rect 253 177 254 178 
<< m2 >>
rect 253 177 254 178 
<< pdiffusion >>
rect 264 177 265 178 
<< pdiffusion >>
rect 265 177 266 178 
<< pdiffusion >>
rect 266 177 267 178 
<< pdiffusion >>
rect 267 177 268 178 
<< pdiffusion >>
rect 268 177 269 178 
<< pdiffusion >>
rect 269 177 270 178 
<< m1 >>
rect 278 177 279 178 
<< m1 >>
rect 280 177 281 178 
<< m2 >>
rect 280 177 281 178 
<< pdiffusion >>
rect 282 177 283 178 
<< pdiffusion >>
rect 283 177 284 178 
<< pdiffusion >>
rect 284 177 285 178 
<< pdiffusion >>
rect 285 177 286 178 
<< pdiffusion >>
rect 286 177 287 178 
<< pdiffusion >>
rect 287 177 288 178 
<< m1 >>
rect 289 177 290 178 
<< pdiffusion >>
rect 300 177 301 178 
<< pdiffusion >>
rect 301 177 302 178 
<< pdiffusion >>
rect 302 177 303 178 
<< pdiffusion >>
rect 303 177 304 178 
<< pdiffusion >>
rect 304 177 305 178 
<< pdiffusion >>
rect 305 177 306 178 
<< m1 >>
rect 307 177 308 178 
<< pdiffusion >>
rect 318 177 319 178 
<< pdiffusion >>
rect 319 177 320 178 
<< pdiffusion >>
rect 320 177 321 178 
<< pdiffusion >>
rect 321 177 322 178 
<< pdiffusion >>
rect 322 177 323 178 
<< pdiffusion >>
rect 323 177 324 178 
<< m1 >>
rect 325 177 326 178 
<< m1 >>
rect 329 177 330 178 
<< pdiffusion >>
rect 336 177 337 178 
<< pdiffusion >>
rect 337 177 338 178 
<< pdiffusion >>
rect 338 177 339 178 
<< pdiffusion >>
rect 339 177 340 178 
<< pdiffusion >>
rect 340 177 341 178 
<< pdiffusion >>
rect 341 177 342 178 
<< m1 >>
rect 343 177 344 178 
<< m1 >>
rect 348 177 349 178 
<< m1 >>
rect 354 177 355 178 
<< m1 >>
rect 366 177 367 178 
<< pdiffusion >>
rect 372 177 373 178 
<< pdiffusion >>
rect 373 177 374 178 
<< pdiffusion >>
rect 374 177 375 178 
<< pdiffusion >>
rect 375 177 376 178 
<< pdiffusion >>
rect 376 177 377 178 
<< pdiffusion >>
rect 377 177 378 178 
<< m1 >>
rect 379 177 380 178 
<< m2 >>
rect 380 177 381 178 
<< m1 >>
rect 383 177 384 178 
<< pdiffusion >>
rect 390 177 391 178 
<< pdiffusion >>
rect 391 177 392 178 
<< pdiffusion >>
rect 392 177 393 178 
<< pdiffusion >>
rect 393 177 394 178 
<< pdiffusion >>
rect 394 177 395 178 
<< pdiffusion >>
rect 395 177 396 178 
<< m1 >>
rect 402 177 403 178 
<< m2 >>
rect 405 177 406 178 
<< m1 >>
rect 406 177 407 178 
<< pdiffusion >>
rect 408 177 409 178 
<< pdiffusion >>
rect 409 177 410 178 
<< pdiffusion >>
rect 410 177 411 178 
<< pdiffusion >>
rect 411 177 412 178 
<< pdiffusion >>
rect 412 177 413 178 
<< pdiffusion >>
rect 413 177 414 178 
<< m1 >>
rect 415 177 416 178 
<< m2 >>
rect 415 177 416 178 
<< m1 >>
rect 417 177 418 178 
<< m2 >>
rect 418 177 419 178 
<< m1 >>
rect 423 177 424 178 
<< pdiffusion >>
rect 426 177 427 178 
<< pdiffusion >>
rect 427 177 428 178 
<< pdiffusion >>
rect 428 177 429 178 
<< pdiffusion >>
rect 429 177 430 178 
<< pdiffusion >>
rect 430 177 431 178 
<< pdiffusion >>
rect 431 177 432 178 
<< m1 >>
rect 433 177 434 178 
<< m1 >>
rect 456 177 457 178 
<< pdiffusion >>
rect 462 177 463 178 
<< pdiffusion >>
rect 463 177 464 178 
<< pdiffusion >>
rect 464 177 465 178 
<< pdiffusion >>
rect 465 177 466 178 
<< pdiffusion >>
rect 466 177 467 178 
<< pdiffusion >>
rect 467 177 468 178 
<< m1 >>
rect 478 177 479 178 
<< m2 >>
rect 478 177 479 178 
<< pdiffusion >>
rect 480 177 481 178 
<< pdiffusion >>
rect 481 177 482 178 
<< pdiffusion >>
rect 482 177 483 178 
<< pdiffusion >>
rect 483 177 484 178 
<< pdiffusion >>
rect 484 177 485 178 
<< pdiffusion >>
rect 485 177 486 178 
<< pdiffusion >>
rect 498 177 499 178 
<< pdiffusion >>
rect 499 177 500 178 
<< pdiffusion >>
rect 500 177 501 178 
<< pdiffusion >>
rect 501 177 502 178 
<< pdiffusion >>
rect 502 177 503 178 
<< pdiffusion >>
rect 503 177 504 178 
<< pdiffusion >>
rect 12 178 13 179 
<< pdiffusion >>
rect 13 178 14 179 
<< pdiffusion >>
rect 14 178 15 179 
<< pdiffusion >>
rect 15 178 16 179 
<< pdiffusion >>
rect 16 178 17 179 
<< pdiffusion >>
rect 17 178 18 179 
<< m1 >>
rect 28 178 29 179 
<< pdiffusion >>
rect 30 178 31 179 
<< pdiffusion >>
rect 31 178 32 179 
<< pdiffusion >>
rect 32 178 33 179 
<< pdiffusion >>
rect 33 178 34 179 
<< pdiffusion >>
rect 34 178 35 179 
<< pdiffusion >>
rect 35 178 36 179 
<< pdiffusion >>
rect 48 178 49 179 
<< pdiffusion >>
rect 49 178 50 179 
<< pdiffusion >>
rect 50 178 51 179 
<< pdiffusion >>
rect 51 178 52 179 
<< pdiffusion >>
rect 52 178 53 179 
<< pdiffusion >>
rect 53 178 54 179 
<< m1 >>
rect 64 178 65 179 
<< pdiffusion >>
rect 66 178 67 179 
<< pdiffusion >>
rect 67 178 68 179 
<< pdiffusion >>
rect 68 178 69 179 
<< pdiffusion >>
rect 69 178 70 179 
<< pdiffusion >>
rect 70 178 71 179 
<< pdiffusion >>
rect 71 178 72 179 
<< pdiffusion >>
rect 84 178 85 179 
<< pdiffusion >>
rect 85 178 86 179 
<< pdiffusion >>
rect 86 178 87 179 
<< pdiffusion >>
rect 87 178 88 179 
<< pdiffusion >>
rect 88 178 89 179 
<< pdiffusion >>
rect 89 178 90 179 
<< m2 >>
rect 97 178 98 179 
<< m1 >>
rect 98 178 99 179 
<< m1 >>
rect 100 178 101 179 
<< pdiffusion >>
rect 102 178 103 179 
<< pdiffusion >>
rect 103 178 104 179 
<< pdiffusion >>
rect 104 178 105 179 
<< pdiffusion >>
rect 105 178 106 179 
<< pdiffusion >>
rect 106 178 107 179 
<< pdiffusion >>
rect 107 178 108 179 
<< m1 >>
rect 114 178 115 179 
<< m2 >>
rect 117 178 118 179 
<< m1 >>
rect 118 178 119 179 
<< pdiffusion >>
rect 120 178 121 179 
<< pdiffusion >>
rect 121 178 122 179 
<< pdiffusion >>
rect 122 178 123 179 
<< pdiffusion >>
rect 123 178 124 179 
<< pdiffusion >>
rect 124 178 125 179 
<< pdiffusion >>
rect 125 178 126 179 
<< m1 >>
rect 127 178 128 179 
<< m1 >>
rect 129 178 130 179 
<< m1 >>
rect 131 178 132 179 
<< pdiffusion >>
rect 138 178 139 179 
<< pdiffusion >>
rect 139 178 140 179 
<< pdiffusion >>
rect 140 178 141 179 
<< pdiffusion >>
rect 141 178 142 179 
<< pdiffusion >>
rect 142 178 143 179 
<< pdiffusion >>
rect 143 178 144 179 
<< pdiffusion >>
rect 156 178 157 179 
<< pdiffusion >>
rect 157 178 158 179 
<< pdiffusion >>
rect 158 178 159 179 
<< pdiffusion >>
rect 159 178 160 179 
<< pdiffusion >>
rect 160 178 161 179 
<< pdiffusion >>
rect 161 178 162 179 
<< m1 >>
rect 163 178 164 179 
<< m2 >>
rect 163 178 164 179 
<< pdiffusion >>
rect 174 178 175 179 
<< pdiffusion >>
rect 175 178 176 179 
<< pdiffusion >>
rect 176 178 177 179 
<< pdiffusion >>
rect 177 178 178 179 
<< pdiffusion >>
rect 178 178 179 179 
<< pdiffusion >>
rect 179 178 180 179 
<< m1 >>
rect 185 178 186 179 
<< m2 >>
rect 189 178 190 179 
<< m1 >>
rect 190 178 191 179 
<< pdiffusion >>
rect 192 178 193 179 
<< pdiffusion >>
rect 193 178 194 179 
<< pdiffusion >>
rect 194 178 195 179 
<< pdiffusion >>
rect 195 178 196 179 
<< pdiffusion >>
rect 196 178 197 179 
<< pdiffusion >>
rect 197 178 198 179 
<< m1 >>
rect 199 178 200 179 
<< m2 >>
rect 199 178 200 179 
<< pdiffusion >>
rect 210 178 211 179 
<< pdiffusion >>
rect 211 178 212 179 
<< pdiffusion >>
rect 212 178 213 179 
<< pdiffusion >>
rect 213 178 214 179 
<< pdiffusion >>
rect 214 178 215 179 
<< pdiffusion >>
rect 215 178 216 179 
<< m1 >>
rect 217 178 218 179 
<< m1 >>
rect 221 178 222 179 
<< m1 >>
rect 226 178 227 179 
<< pdiffusion >>
rect 228 178 229 179 
<< pdiffusion >>
rect 229 178 230 179 
<< pdiffusion >>
rect 230 178 231 179 
<< pdiffusion >>
rect 231 178 232 179 
<< pdiffusion >>
rect 232 178 233 179 
<< pdiffusion >>
rect 233 178 234 179 
<< m1 >>
rect 235 178 236 179 
<< m2 >>
rect 236 178 237 179 
<< m1 >>
rect 244 178 245 179 
<< m2 >>
rect 244 178 245 179 
<< pdiffusion >>
rect 246 178 247 179 
<< pdiffusion >>
rect 247 178 248 179 
<< pdiffusion >>
rect 248 178 249 179 
<< pdiffusion >>
rect 249 178 250 179 
<< pdiffusion >>
rect 250 178 251 179 
<< pdiffusion >>
rect 251 178 252 179 
<< m1 >>
rect 253 178 254 179 
<< m2 >>
rect 253 178 254 179 
<< pdiffusion >>
rect 264 178 265 179 
<< pdiffusion >>
rect 265 178 266 179 
<< pdiffusion >>
rect 266 178 267 179 
<< pdiffusion >>
rect 267 178 268 179 
<< pdiffusion >>
rect 268 178 269 179 
<< pdiffusion >>
rect 269 178 270 179 
<< m1 >>
rect 278 178 279 179 
<< m1 >>
rect 280 178 281 179 
<< m2 >>
rect 280 178 281 179 
<< pdiffusion >>
rect 282 178 283 179 
<< pdiffusion >>
rect 283 178 284 179 
<< pdiffusion >>
rect 284 178 285 179 
<< pdiffusion >>
rect 285 178 286 179 
<< pdiffusion >>
rect 286 178 287 179 
<< pdiffusion >>
rect 287 178 288 179 
<< m1 >>
rect 289 178 290 179 
<< pdiffusion >>
rect 300 178 301 179 
<< pdiffusion >>
rect 301 178 302 179 
<< pdiffusion >>
rect 302 178 303 179 
<< pdiffusion >>
rect 303 178 304 179 
<< pdiffusion >>
rect 304 178 305 179 
<< pdiffusion >>
rect 305 178 306 179 
<< m1 >>
rect 307 178 308 179 
<< pdiffusion >>
rect 318 178 319 179 
<< pdiffusion >>
rect 319 178 320 179 
<< pdiffusion >>
rect 320 178 321 179 
<< pdiffusion >>
rect 321 178 322 179 
<< pdiffusion >>
rect 322 178 323 179 
<< pdiffusion >>
rect 323 178 324 179 
<< m1 >>
rect 325 178 326 179 
<< m1 >>
rect 329 178 330 179 
<< pdiffusion >>
rect 336 178 337 179 
<< pdiffusion >>
rect 337 178 338 179 
<< pdiffusion >>
rect 338 178 339 179 
<< pdiffusion >>
rect 339 178 340 179 
<< pdiffusion >>
rect 340 178 341 179 
<< pdiffusion >>
rect 341 178 342 179 
<< m1 >>
rect 343 178 344 179 
<< m1 >>
rect 348 178 349 179 
<< m1 >>
rect 354 178 355 179 
<< m1 >>
rect 366 178 367 179 
<< pdiffusion >>
rect 372 178 373 179 
<< pdiffusion >>
rect 373 178 374 179 
<< pdiffusion >>
rect 374 178 375 179 
<< pdiffusion >>
rect 375 178 376 179 
<< pdiffusion >>
rect 376 178 377 179 
<< pdiffusion >>
rect 377 178 378 179 
<< m1 >>
rect 379 178 380 179 
<< m2 >>
rect 380 178 381 179 
<< m1 >>
rect 383 178 384 179 
<< pdiffusion >>
rect 390 178 391 179 
<< pdiffusion >>
rect 391 178 392 179 
<< pdiffusion >>
rect 392 178 393 179 
<< pdiffusion >>
rect 393 178 394 179 
<< pdiffusion >>
rect 394 178 395 179 
<< pdiffusion >>
rect 395 178 396 179 
<< m1 >>
rect 402 178 403 179 
<< m2 >>
rect 405 178 406 179 
<< m1 >>
rect 406 178 407 179 
<< pdiffusion >>
rect 408 178 409 179 
<< pdiffusion >>
rect 409 178 410 179 
<< pdiffusion >>
rect 410 178 411 179 
<< pdiffusion >>
rect 411 178 412 179 
<< pdiffusion >>
rect 412 178 413 179 
<< pdiffusion >>
rect 413 178 414 179 
<< m1 >>
rect 415 178 416 179 
<< m2 >>
rect 415 178 416 179 
<< m1 >>
rect 417 178 418 179 
<< m2 >>
rect 418 178 419 179 
<< m1 >>
rect 419 178 420 179 
<< m2 >>
rect 419 178 420 179 
<< m2c >>
rect 419 178 420 179 
<< m1 >>
rect 419 178 420 179 
<< m2 >>
rect 419 178 420 179 
<< m1 >>
rect 420 178 421 179 
<< m1 >>
rect 421 178 422 179 
<< m1 >>
rect 423 178 424 179 
<< pdiffusion >>
rect 426 178 427 179 
<< pdiffusion >>
rect 427 178 428 179 
<< pdiffusion >>
rect 428 178 429 179 
<< pdiffusion >>
rect 429 178 430 179 
<< pdiffusion >>
rect 430 178 431 179 
<< pdiffusion >>
rect 431 178 432 179 
<< m1 >>
rect 433 178 434 179 
<< m1 >>
rect 456 178 457 179 
<< pdiffusion >>
rect 462 178 463 179 
<< pdiffusion >>
rect 463 178 464 179 
<< pdiffusion >>
rect 464 178 465 179 
<< pdiffusion >>
rect 465 178 466 179 
<< pdiffusion >>
rect 466 178 467 179 
<< pdiffusion >>
rect 467 178 468 179 
<< m1 >>
rect 478 178 479 179 
<< m2 >>
rect 478 178 479 179 
<< pdiffusion >>
rect 480 178 481 179 
<< pdiffusion >>
rect 481 178 482 179 
<< pdiffusion >>
rect 482 178 483 179 
<< pdiffusion >>
rect 483 178 484 179 
<< pdiffusion >>
rect 484 178 485 179 
<< pdiffusion >>
rect 485 178 486 179 
<< pdiffusion >>
rect 498 178 499 179 
<< pdiffusion >>
rect 499 178 500 179 
<< pdiffusion >>
rect 500 178 501 179 
<< pdiffusion >>
rect 501 178 502 179 
<< pdiffusion >>
rect 502 178 503 179 
<< pdiffusion >>
rect 503 178 504 179 
<< pdiffusion >>
rect 12 179 13 180 
<< pdiffusion >>
rect 13 179 14 180 
<< pdiffusion >>
rect 14 179 15 180 
<< pdiffusion >>
rect 15 179 16 180 
<< pdiffusion >>
rect 16 179 17 180 
<< pdiffusion >>
rect 17 179 18 180 
<< m1 >>
rect 28 179 29 180 
<< pdiffusion >>
rect 30 179 31 180 
<< pdiffusion >>
rect 31 179 32 180 
<< pdiffusion >>
rect 32 179 33 180 
<< pdiffusion >>
rect 33 179 34 180 
<< pdiffusion >>
rect 34 179 35 180 
<< pdiffusion >>
rect 35 179 36 180 
<< pdiffusion >>
rect 48 179 49 180 
<< pdiffusion >>
rect 49 179 50 180 
<< pdiffusion >>
rect 50 179 51 180 
<< pdiffusion >>
rect 51 179 52 180 
<< pdiffusion >>
rect 52 179 53 180 
<< pdiffusion >>
rect 53 179 54 180 
<< m1 >>
rect 64 179 65 180 
<< pdiffusion >>
rect 66 179 67 180 
<< pdiffusion >>
rect 67 179 68 180 
<< pdiffusion >>
rect 68 179 69 180 
<< pdiffusion >>
rect 69 179 70 180 
<< pdiffusion >>
rect 70 179 71 180 
<< pdiffusion >>
rect 71 179 72 180 
<< pdiffusion >>
rect 84 179 85 180 
<< pdiffusion >>
rect 85 179 86 180 
<< pdiffusion >>
rect 86 179 87 180 
<< pdiffusion >>
rect 87 179 88 180 
<< pdiffusion >>
rect 88 179 89 180 
<< pdiffusion >>
rect 89 179 90 180 
<< m2 >>
rect 97 179 98 180 
<< m1 >>
rect 98 179 99 180 
<< m1 >>
rect 100 179 101 180 
<< pdiffusion >>
rect 102 179 103 180 
<< pdiffusion >>
rect 103 179 104 180 
<< pdiffusion >>
rect 104 179 105 180 
<< pdiffusion >>
rect 105 179 106 180 
<< pdiffusion >>
rect 106 179 107 180 
<< pdiffusion >>
rect 107 179 108 180 
<< m1 >>
rect 114 179 115 180 
<< m2 >>
rect 117 179 118 180 
<< m1 >>
rect 118 179 119 180 
<< pdiffusion >>
rect 120 179 121 180 
<< pdiffusion >>
rect 121 179 122 180 
<< pdiffusion >>
rect 122 179 123 180 
<< pdiffusion >>
rect 123 179 124 180 
<< pdiffusion >>
rect 124 179 125 180 
<< pdiffusion >>
rect 125 179 126 180 
<< m1 >>
rect 127 179 128 180 
<< m1 >>
rect 129 179 130 180 
<< m1 >>
rect 131 179 132 180 
<< pdiffusion >>
rect 138 179 139 180 
<< pdiffusion >>
rect 139 179 140 180 
<< pdiffusion >>
rect 140 179 141 180 
<< pdiffusion >>
rect 141 179 142 180 
<< pdiffusion >>
rect 142 179 143 180 
<< pdiffusion >>
rect 143 179 144 180 
<< pdiffusion >>
rect 156 179 157 180 
<< pdiffusion >>
rect 157 179 158 180 
<< pdiffusion >>
rect 158 179 159 180 
<< pdiffusion >>
rect 159 179 160 180 
<< pdiffusion >>
rect 160 179 161 180 
<< pdiffusion >>
rect 161 179 162 180 
<< m1 >>
rect 163 179 164 180 
<< m2 >>
rect 163 179 164 180 
<< pdiffusion >>
rect 174 179 175 180 
<< m1 >>
rect 175 179 176 180 
<< pdiffusion >>
rect 175 179 176 180 
<< pdiffusion >>
rect 176 179 177 180 
<< pdiffusion >>
rect 177 179 178 180 
<< pdiffusion >>
rect 178 179 179 180 
<< pdiffusion >>
rect 179 179 180 180 
<< m1 >>
rect 185 179 186 180 
<< m2 >>
rect 189 179 190 180 
<< m1 >>
rect 190 179 191 180 
<< pdiffusion >>
rect 192 179 193 180 
<< pdiffusion >>
rect 193 179 194 180 
<< pdiffusion >>
rect 194 179 195 180 
<< pdiffusion >>
rect 195 179 196 180 
<< m1 >>
rect 196 179 197 180 
<< pdiffusion >>
rect 196 179 197 180 
<< pdiffusion >>
rect 197 179 198 180 
<< m1 >>
rect 199 179 200 180 
<< m2 >>
rect 199 179 200 180 
<< pdiffusion >>
rect 210 179 211 180 
<< pdiffusion >>
rect 211 179 212 180 
<< pdiffusion >>
rect 212 179 213 180 
<< pdiffusion >>
rect 213 179 214 180 
<< m1 >>
rect 214 179 215 180 
<< pdiffusion >>
rect 214 179 215 180 
<< pdiffusion >>
rect 215 179 216 180 
<< m1 >>
rect 217 179 218 180 
<< m1 >>
rect 221 179 222 180 
<< m1 >>
rect 226 179 227 180 
<< pdiffusion >>
rect 228 179 229 180 
<< pdiffusion >>
rect 229 179 230 180 
<< pdiffusion >>
rect 230 179 231 180 
<< pdiffusion >>
rect 231 179 232 180 
<< m1 >>
rect 232 179 233 180 
<< pdiffusion >>
rect 232 179 233 180 
<< pdiffusion >>
rect 233 179 234 180 
<< m1 >>
rect 235 179 236 180 
<< m2 >>
rect 236 179 237 180 
<< m1 >>
rect 244 179 245 180 
<< m2 >>
rect 244 179 245 180 
<< pdiffusion >>
rect 246 179 247 180 
<< pdiffusion >>
rect 247 179 248 180 
<< pdiffusion >>
rect 248 179 249 180 
<< pdiffusion >>
rect 249 179 250 180 
<< pdiffusion >>
rect 250 179 251 180 
<< pdiffusion >>
rect 251 179 252 180 
<< m1 >>
rect 253 179 254 180 
<< m2 >>
rect 253 179 254 180 
<< pdiffusion >>
rect 264 179 265 180 
<< pdiffusion >>
rect 265 179 266 180 
<< pdiffusion >>
rect 266 179 267 180 
<< pdiffusion >>
rect 267 179 268 180 
<< pdiffusion >>
rect 268 179 269 180 
<< pdiffusion >>
rect 269 179 270 180 
<< m1 >>
rect 278 179 279 180 
<< m1 >>
rect 280 179 281 180 
<< m2 >>
rect 280 179 281 180 
<< pdiffusion >>
rect 282 179 283 180 
<< pdiffusion >>
rect 283 179 284 180 
<< pdiffusion >>
rect 284 179 285 180 
<< pdiffusion >>
rect 285 179 286 180 
<< pdiffusion >>
rect 286 179 287 180 
<< pdiffusion >>
rect 287 179 288 180 
<< m1 >>
rect 289 179 290 180 
<< pdiffusion >>
rect 300 179 301 180 
<< pdiffusion >>
rect 301 179 302 180 
<< pdiffusion >>
rect 302 179 303 180 
<< pdiffusion >>
rect 303 179 304 180 
<< m1 >>
rect 304 179 305 180 
<< pdiffusion >>
rect 304 179 305 180 
<< pdiffusion >>
rect 305 179 306 180 
<< m1 >>
rect 307 179 308 180 
<< pdiffusion >>
rect 318 179 319 180 
<< pdiffusion >>
rect 319 179 320 180 
<< pdiffusion >>
rect 320 179 321 180 
<< pdiffusion >>
rect 321 179 322 180 
<< m1 >>
rect 322 179 323 180 
<< pdiffusion >>
rect 322 179 323 180 
<< pdiffusion >>
rect 323 179 324 180 
<< m1 >>
rect 325 179 326 180 
<< m1 >>
rect 329 179 330 180 
<< pdiffusion >>
rect 336 179 337 180 
<< pdiffusion >>
rect 337 179 338 180 
<< pdiffusion >>
rect 338 179 339 180 
<< pdiffusion >>
rect 339 179 340 180 
<< pdiffusion >>
rect 340 179 341 180 
<< pdiffusion >>
rect 341 179 342 180 
<< m1 >>
rect 343 179 344 180 
<< m1 >>
rect 348 179 349 180 
<< m1 >>
rect 354 179 355 180 
<< m1 >>
rect 366 179 367 180 
<< pdiffusion >>
rect 372 179 373 180 
<< m1 >>
rect 373 179 374 180 
<< pdiffusion >>
rect 373 179 374 180 
<< pdiffusion >>
rect 374 179 375 180 
<< pdiffusion >>
rect 375 179 376 180 
<< pdiffusion >>
rect 376 179 377 180 
<< pdiffusion >>
rect 377 179 378 180 
<< m1 >>
rect 379 179 380 180 
<< m2 >>
rect 380 179 381 180 
<< m1 >>
rect 383 179 384 180 
<< pdiffusion >>
rect 390 179 391 180 
<< m1 >>
rect 391 179 392 180 
<< pdiffusion >>
rect 391 179 392 180 
<< pdiffusion >>
rect 392 179 393 180 
<< pdiffusion >>
rect 393 179 394 180 
<< pdiffusion >>
rect 394 179 395 180 
<< pdiffusion >>
rect 395 179 396 180 
<< m1 >>
rect 402 179 403 180 
<< m2 >>
rect 405 179 406 180 
<< m1 >>
rect 406 179 407 180 
<< pdiffusion >>
rect 408 179 409 180 
<< m1 >>
rect 409 179 410 180 
<< pdiffusion >>
rect 409 179 410 180 
<< pdiffusion >>
rect 410 179 411 180 
<< pdiffusion >>
rect 411 179 412 180 
<< pdiffusion >>
rect 412 179 413 180 
<< pdiffusion >>
rect 413 179 414 180 
<< m1 >>
rect 415 179 416 180 
<< m2 >>
rect 415 179 416 180 
<< m1 >>
rect 417 179 418 180 
<< m1 >>
rect 421 179 422 180 
<< m2 >>
rect 421 179 422 180 
<< m2c >>
rect 421 179 422 180 
<< m1 >>
rect 421 179 422 180 
<< m2 >>
rect 421 179 422 180 
<< m1 >>
rect 423 179 424 180 
<< m2 >>
rect 423 179 424 180 
<< m2c >>
rect 423 179 424 180 
<< m1 >>
rect 423 179 424 180 
<< m2 >>
rect 423 179 424 180 
<< pdiffusion >>
rect 426 179 427 180 
<< pdiffusion >>
rect 427 179 428 180 
<< pdiffusion >>
rect 428 179 429 180 
<< pdiffusion >>
rect 429 179 430 180 
<< pdiffusion >>
rect 430 179 431 180 
<< pdiffusion >>
rect 431 179 432 180 
<< m1 >>
rect 433 179 434 180 
<< m1 >>
rect 456 179 457 180 
<< pdiffusion >>
rect 462 179 463 180 
<< pdiffusion >>
rect 463 179 464 180 
<< pdiffusion >>
rect 464 179 465 180 
<< pdiffusion >>
rect 465 179 466 180 
<< pdiffusion >>
rect 466 179 467 180 
<< pdiffusion >>
rect 467 179 468 180 
<< m1 >>
rect 478 179 479 180 
<< m2 >>
rect 478 179 479 180 
<< pdiffusion >>
rect 480 179 481 180 
<< pdiffusion >>
rect 481 179 482 180 
<< pdiffusion >>
rect 482 179 483 180 
<< pdiffusion >>
rect 483 179 484 180 
<< pdiffusion >>
rect 484 179 485 180 
<< pdiffusion >>
rect 485 179 486 180 
<< pdiffusion >>
rect 498 179 499 180 
<< pdiffusion >>
rect 499 179 500 180 
<< pdiffusion >>
rect 500 179 501 180 
<< pdiffusion >>
rect 501 179 502 180 
<< pdiffusion >>
rect 502 179 503 180 
<< pdiffusion >>
rect 503 179 504 180 
<< m1 >>
rect 28 180 29 181 
<< m1 >>
rect 64 180 65 181 
<< m2 >>
rect 97 180 98 181 
<< m1 >>
rect 98 180 99 181 
<< m1 >>
rect 100 180 101 181 
<< m1 >>
rect 114 180 115 181 
<< m2 >>
rect 117 180 118 181 
<< m1 >>
rect 118 180 119 181 
<< m1 >>
rect 127 180 128 181 
<< m1 >>
rect 129 180 130 181 
<< m1 >>
rect 131 180 132 181 
<< m1 >>
rect 163 180 164 181 
<< m2 >>
rect 163 180 164 181 
<< m1 >>
rect 175 180 176 181 
<< m1 >>
rect 185 180 186 181 
<< m2 >>
rect 189 180 190 181 
<< m1 >>
rect 190 180 191 181 
<< m1 >>
rect 196 180 197 181 
<< m1 >>
rect 199 180 200 181 
<< m2 >>
rect 199 180 200 181 
<< m1 >>
rect 214 180 215 181 
<< m1 >>
rect 217 180 218 181 
<< m1 >>
rect 221 180 222 181 
<< m1 >>
rect 226 180 227 181 
<< m1 >>
rect 232 180 233 181 
<< m1 >>
rect 235 180 236 181 
<< m2 >>
rect 236 180 237 181 
<< m1 >>
rect 244 180 245 181 
<< m2 >>
rect 244 180 245 181 
<< m1 >>
rect 253 180 254 181 
<< m2 >>
rect 253 180 254 181 
<< m1 >>
rect 278 180 279 181 
<< m1 >>
rect 280 180 281 181 
<< m2 >>
rect 280 180 281 181 
<< m1 >>
rect 289 180 290 181 
<< m1 >>
rect 304 180 305 181 
<< m1 >>
rect 307 180 308 181 
<< m1 >>
rect 322 180 323 181 
<< m1 >>
rect 325 180 326 181 
<< m1 >>
rect 329 180 330 181 
<< m1 >>
rect 343 180 344 181 
<< m1 >>
rect 348 180 349 181 
<< m1 >>
rect 354 180 355 181 
<< m1 >>
rect 366 180 367 181 
<< m1 >>
rect 373 180 374 181 
<< m1 >>
rect 379 180 380 181 
<< m2 >>
rect 380 180 381 181 
<< m1 >>
rect 383 180 384 181 
<< m1 >>
rect 391 180 392 181 
<< m1 >>
rect 402 180 403 181 
<< m2 >>
rect 405 180 406 181 
<< m1 >>
rect 406 180 407 181 
<< m1 >>
rect 409 180 410 181 
<< m1 >>
rect 415 180 416 181 
<< m2 >>
rect 415 180 416 181 
<< m2 >>
rect 416 180 417 181 
<< m1 >>
rect 417 180 418 181 
<< m2 >>
rect 417 180 418 181 
<< m2 >>
rect 418 180 419 181 
<< m2 >>
rect 419 180 420 181 
<< m2 >>
rect 421 180 422 181 
<< m2 >>
rect 423 180 424 181 
<< m1 >>
rect 433 180 434 181 
<< m1 >>
rect 456 180 457 181 
<< m1 >>
rect 478 180 479 181 
<< m2 >>
rect 478 180 479 181 
<< m1 >>
rect 28 181 29 182 
<< m1 >>
rect 64 181 65 182 
<< m2 >>
rect 97 181 98 182 
<< m1 >>
rect 98 181 99 182 
<< m1 >>
rect 100 181 101 182 
<< m1 >>
rect 114 181 115 182 
<< m2 >>
rect 117 181 118 182 
<< m1 >>
rect 118 181 119 182 
<< m2 >>
rect 118 181 119 182 
<< m2 >>
rect 119 181 120 182 
<< m1 >>
rect 120 181 121 182 
<< m2 >>
rect 120 181 121 182 
<< m2c >>
rect 120 181 121 182 
<< m1 >>
rect 120 181 121 182 
<< m2 >>
rect 120 181 121 182 
<< m1 >>
rect 127 181 128 182 
<< m1 >>
rect 129 181 130 182 
<< m1 >>
rect 131 181 132 182 
<< m1 >>
rect 163 181 164 182 
<< m2 >>
rect 163 181 164 182 
<< m1 >>
rect 164 181 165 182 
<< m1 >>
rect 165 181 166 182 
<< m1 >>
rect 166 181 167 182 
<< m1 >>
rect 167 181 168 182 
<< m1 >>
rect 168 181 169 182 
<< m1 >>
rect 169 181 170 182 
<< m1 >>
rect 170 181 171 182 
<< m1 >>
rect 171 181 172 182 
<< m1 >>
rect 172 181 173 182 
<< m1 >>
rect 173 181 174 182 
<< m1 >>
rect 174 181 175 182 
<< m1 >>
rect 175 181 176 182 
<< m1 >>
rect 185 181 186 182 
<< m2 >>
rect 189 181 190 182 
<< m1 >>
rect 190 181 191 182 
<< m1 >>
rect 196 181 197 182 
<< m1 >>
rect 197 181 198 182 
<< m1 >>
rect 198 181 199 182 
<< m1 >>
rect 199 181 200 182 
<< m2 >>
rect 199 181 200 182 
<< m1 >>
rect 214 181 215 182 
<< m1 >>
rect 217 181 218 182 
<< m1 >>
rect 221 181 222 182 
<< m1 >>
rect 226 181 227 182 
<< m1 >>
rect 231 181 232 182 
<< m1 >>
rect 232 181 233 182 
<< m1 >>
rect 235 181 236 182 
<< m2 >>
rect 236 181 237 182 
<< m1 >>
rect 244 181 245 182 
<< m2 >>
rect 244 181 245 182 
<< m1 >>
rect 253 181 254 182 
<< m2 >>
rect 253 181 254 182 
<< m1 >>
rect 278 181 279 182 
<< m1 >>
rect 280 181 281 182 
<< m2 >>
rect 280 181 281 182 
<< m1 >>
rect 289 181 290 182 
<< m1 >>
rect 304 181 305 182 
<< m1 >>
rect 305 181 306 182 
<< m1 >>
rect 306 181 307 182 
<< m1 >>
rect 307 181 308 182 
<< m1 >>
rect 321 181 322 182 
<< m1 >>
rect 322 181 323 182 
<< m1 >>
rect 325 181 326 182 
<< m1 >>
rect 329 181 330 182 
<< m1 >>
rect 343 181 344 182 
<< m1 >>
rect 348 181 349 182 
<< m1 >>
rect 354 181 355 182 
<< m1 >>
rect 366 181 367 182 
<< m1 >>
rect 367 181 368 182 
<< m1 >>
rect 368 181 369 182 
<< m1 >>
rect 369 181 370 182 
<< m1 >>
rect 370 181 371 182 
<< m1 >>
rect 371 181 372 182 
<< m1 >>
rect 372 181 373 182 
<< m1 >>
rect 373 181 374 182 
<< m1 >>
rect 377 181 378 182 
<< m2 >>
rect 377 181 378 182 
<< m2c >>
rect 377 181 378 182 
<< m1 >>
rect 377 181 378 182 
<< m2 >>
rect 377 181 378 182 
<< m2 >>
rect 378 181 379 182 
<< m1 >>
rect 379 181 380 182 
<< m2 >>
rect 379 181 380 182 
<< m2 >>
rect 380 181 381 182 
<< m1 >>
rect 383 181 384 182 
<< m1 >>
rect 391 181 392 182 
<< m1 >>
rect 402 181 403 182 
<< m2 >>
rect 405 181 406 182 
<< m1 >>
rect 406 181 407 182 
<< m1 >>
rect 409 181 410 182 
<< m1 >>
rect 410 181 411 182 
<< m1 >>
rect 415 181 416 182 
<< m1 >>
rect 417 181 418 182 
<< m1 >>
rect 418 181 419 182 
<< m1 >>
rect 419 181 420 182 
<< m2 >>
rect 419 181 420 182 
<< m1 >>
rect 420 181 421 182 
<< m1 >>
rect 421 181 422 182 
<< m2 >>
rect 421 181 422 182 
<< m1 >>
rect 422 181 423 182 
<< m1 >>
rect 423 181 424 182 
<< m2 >>
rect 423 181 424 182 
<< m1 >>
rect 424 181 425 182 
<< m1 >>
rect 425 181 426 182 
<< m1 >>
rect 426 181 427 182 
<< m1 >>
rect 433 181 434 182 
<< m1 >>
rect 456 181 457 182 
<< m1 >>
rect 478 181 479 182 
<< m2 >>
rect 478 181 479 182 
<< m1 >>
rect 28 182 29 183 
<< m1 >>
rect 64 182 65 183 
<< m2 >>
rect 97 182 98 183 
<< m1 >>
rect 98 182 99 183 
<< m1 >>
rect 100 182 101 183 
<< m1 >>
rect 114 182 115 183 
<< m1 >>
rect 118 182 119 183 
<< m1 >>
rect 120 182 121 183 
<< m1 >>
rect 122 182 123 183 
<< m2 >>
rect 122 182 123 183 
<< m2c >>
rect 122 182 123 183 
<< m1 >>
rect 122 182 123 183 
<< m2 >>
rect 122 182 123 183 
<< m1 >>
rect 123 182 124 183 
<< m1 >>
rect 124 182 125 183 
<< m1 >>
rect 125 182 126 183 
<< m2 >>
rect 125 182 126 183 
<< m2c >>
rect 125 182 126 183 
<< m1 >>
rect 125 182 126 183 
<< m2 >>
rect 125 182 126 183 
<< m2 >>
rect 126 182 127 183 
<< m1 >>
rect 127 182 128 183 
<< m2 >>
rect 127 182 128 183 
<< m2 >>
rect 128 182 129 183 
<< m1 >>
rect 129 182 130 183 
<< m2 >>
rect 129 182 130 183 
<< m2 >>
rect 130 182 131 183 
<< m1 >>
rect 131 182 132 183 
<< m2 >>
rect 131 182 132 183 
<< m2c >>
rect 131 182 132 183 
<< m1 >>
rect 131 182 132 183 
<< m2 >>
rect 131 182 132 183 
<< m2 >>
rect 163 182 164 183 
<< m1 >>
rect 185 182 186 183 
<< m2 >>
rect 189 182 190 183 
<< m1 >>
rect 190 182 191 183 
<< m1 >>
rect 191 182 192 183 
<< m1 >>
rect 192 182 193 183 
<< m2 >>
rect 192 182 193 183 
<< m2c >>
rect 192 182 193 183 
<< m1 >>
rect 192 182 193 183 
<< m2 >>
rect 192 182 193 183 
<< m2 >>
rect 199 182 200 183 
<< m1 >>
rect 214 182 215 183 
<< m1 >>
rect 217 182 218 183 
<< m1 >>
rect 221 182 222 183 
<< m2 >>
rect 221 182 222 183 
<< m2c >>
rect 221 182 222 183 
<< m1 >>
rect 221 182 222 183 
<< m2 >>
rect 221 182 222 183 
<< m1 >>
rect 226 182 227 183 
<< m2 >>
rect 226 182 227 183 
<< m2c >>
rect 226 182 227 183 
<< m1 >>
rect 226 182 227 183 
<< m2 >>
rect 226 182 227 183 
<< m1 >>
rect 231 182 232 183 
<< m2 >>
rect 231 182 232 183 
<< m2c >>
rect 231 182 232 183 
<< m1 >>
rect 231 182 232 183 
<< m2 >>
rect 231 182 232 183 
<< m1 >>
rect 235 182 236 183 
<< m2 >>
rect 236 182 237 183 
<< m1 >>
rect 237 182 238 183 
<< m2 >>
rect 237 182 238 183 
<< m2c >>
rect 237 182 238 183 
<< m1 >>
rect 237 182 238 183 
<< m2 >>
rect 237 182 238 183 
<< m1 >>
rect 238 182 239 183 
<< m1 >>
rect 239 182 240 183 
<< m1 >>
rect 240 182 241 183 
<< m1 >>
rect 241 182 242 183 
<< m1 >>
rect 242 182 243 183 
<< m1 >>
rect 244 182 245 183 
<< m2 >>
rect 244 182 245 183 
<< m1 >>
rect 253 182 254 183 
<< m2 >>
rect 253 182 254 183 
<< m1 >>
rect 278 182 279 183 
<< m1 >>
rect 280 182 281 183 
<< m2 >>
rect 280 182 281 183 
<< m1 >>
rect 289 182 290 183 
<< m1 >>
rect 321 182 322 183 
<< m2 >>
rect 321 182 322 183 
<< m2c >>
rect 321 182 322 183 
<< m1 >>
rect 321 182 322 183 
<< m2 >>
rect 321 182 322 183 
<< m1 >>
rect 325 182 326 183 
<< m1 >>
rect 329 182 330 183 
<< m2 >>
rect 329 182 330 183 
<< m2c >>
rect 329 182 330 183 
<< m1 >>
rect 329 182 330 183 
<< m2 >>
rect 329 182 330 183 
<< m1 >>
rect 343 182 344 183 
<< m1 >>
rect 348 182 349 183 
<< m2 >>
rect 348 182 349 183 
<< m2c >>
rect 348 182 349 183 
<< m1 >>
rect 348 182 349 183 
<< m2 >>
rect 348 182 349 183 
<< m1 >>
rect 354 182 355 183 
<< m2 >>
rect 354 182 355 183 
<< m2c >>
rect 354 182 355 183 
<< m1 >>
rect 354 182 355 183 
<< m2 >>
rect 354 182 355 183 
<< m1 >>
rect 377 182 378 183 
<< m1 >>
rect 379 182 380 183 
<< m1 >>
rect 383 182 384 183 
<< m2 >>
rect 383 182 384 183 
<< m2c >>
rect 383 182 384 183 
<< m1 >>
rect 383 182 384 183 
<< m2 >>
rect 383 182 384 183 
<< m1 >>
rect 391 182 392 183 
<< m1 >>
rect 392 182 393 183 
<< m1 >>
rect 393 182 394 183 
<< m1 >>
rect 394 182 395 183 
<< m1 >>
rect 395 182 396 183 
<< m1 >>
rect 396 182 397 183 
<< m1 >>
rect 397 182 398 183 
<< m1 >>
rect 398 182 399 183 
<< m1 >>
rect 399 182 400 183 
<< m1 >>
rect 400 182 401 183 
<< m2 >>
rect 400 182 401 183 
<< m2c >>
rect 400 182 401 183 
<< m1 >>
rect 400 182 401 183 
<< m2 >>
rect 400 182 401 183 
<< m2 >>
rect 401 182 402 183 
<< m1 >>
rect 402 182 403 183 
<< m2 >>
rect 402 182 403 183 
<< m2 >>
rect 403 182 404 183 
<< m1 >>
rect 404 182 405 183 
<< m2 >>
rect 404 182 405 183 
<< m2c >>
rect 404 182 405 183 
<< m1 >>
rect 404 182 405 183 
<< m2 >>
rect 404 182 405 183 
<< m2 >>
rect 405 182 406 183 
<< m1 >>
rect 406 182 407 183 
<< m1 >>
rect 410 182 411 183 
<< m2 >>
rect 410 182 411 183 
<< m2c >>
rect 410 182 411 183 
<< m1 >>
rect 410 182 411 183 
<< m2 >>
rect 410 182 411 183 
<< m1 >>
rect 415 182 416 183 
<< m2 >>
rect 419 182 420 183 
<< m2 >>
rect 421 182 422 183 
<< m2 >>
rect 423 182 424 183 
<< m1 >>
rect 426 182 427 183 
<< m2 >>
rect 426 182 427 183 
<< m2c >>
rect 426 182 427 183 
<< m1 >>
rect 426 182 427 183 
<< m2 >>
rect 426 182 427 183 
<< m1 >>
rect 433 182 434 183 
<< m2 >>
rect 433 182 434 183 
<< m2c >>
rect 433 182 434 183 
<< m1 >>
rect 433 182 434 183 
<< m2 >>
rect 433 182 434 183 
<< m1 >>
rect 456 182 457 183 
<< m2 >>
rect 456 182 457 183 
<< m2c >>
rect 456 182 457 183 
<< m1 >>
rect 456 182 457 183 
<< m2 >>
rect 456 182 457 183 
<< m1 >>
rect 478 182 479 183 
<< m2 >>
rect 478 182 479 183 
<< m1 >>
rect 28 183 29 184 
<< m1 >>
rect 64 183 65 184 
<< m2 >>
rect 97 183 98 184 
<< m1 >>
rect 98 183 99 184 
<< m1 >>
rect 100 183 101 184 
<< m1 >>
rect 114 183 115 184 
<< m1 >>
rect 115 183 116 184 
<< m1 >>
rect 116 183 117 184 
<< m2 >>
rect 116 183 117 184 
<< m2c >>
rect 116 183 117 184 
<< m1 >>
rect 116 183 117 184 
<< m2 >>
rect 116 183 117 184 
<< m2 >>
rect 117 183 118 184 
<< m1 >>
rect 118 183 119 184 
<< m2 >>
rect 118 183 119 184 
<< m2 >>
rect 119 183 120 184 
<< m1 >>
rect 120 183 121 184 
<< m2 >>
rect 120 183 121 184 
<< m2 >>
rect 122 183 123 184 
<< m1 >>
rect 127 183 128 184 
<< m1 >>
rect 129 183 130 184 
<< m2 >>
rect 163 183 164 184 
<< m1 >>
rect 185 183 186 184 
<< m2 >>
rect 189 183 190 184 
<< m2 >>
rect 192 183 193 184 
<< m1 >>
rect 199 183 200 184 
<< m2 >>
rect 199 183 200 184 
<< m2c >>
rect 199 183 200 184 
<< m1 >>
rect 199 183 200 184 
<< m2 >>
rect 199 183 200 184 
<< m1 >>
rect 214 183 215 184 
<< m1 >>
rect 217 183 218 184 
<< m2 >>
rect 221 183 222 184 
<< m2 >>
rect 226 183 227 184 
<< m2 >>
rect 231 183 232 184 
<< m1 >>
rect 235 183 236 184 
<< m1 >>
rect 242 183 243 184 
<< m1 >>
rect 244 183 245 184 
<< m2 >>
rect 244 183 245 184 
<< m1 >>
rect 253 183 254 184 
<< m2 >>
rect 253 183 254 184 
<< m1 >>
rect 278 183 279 184 
<< m1 >>
rect 280 183 281 184 
<< m2 >>
rect 280 183 281 184 
<< m1 >>
rect 289 183 290 184 
<< m2 >>
rect 321 183 322 184 
<< m1 >>
rect 325 183 326 184 
<< m2 >>
rect 329 183 330 184 
<< m1 >>
rect 343 183 344 184 
<< m2 >>
rect 348 183 349 184 
<< m2 >>
rect 354 183 355 184 
<< m1 >>
rect 377 183 378 184 
<< m1 >>
rect 379 183 380 184 
<< m2 >>
rect 383 183 384 184 
<< m1 >>
rect 402 183 403 184 
<< m1 >>
rect 406 183 407 184 
<< m2 >>
rect 410 183 411 184 
<< m1 >>
rect 415 183 416 184 
<< m1 >>
rect 419 183 420 184 
<< m2 >>
rect 419 183 420 184 
<< m2c >>
rect 419 183 420 184 
<< m1 >>
rect 419 183 420 184 
<< m2 >>
rect 419 183 420 184 
<< m1 >>
rect 421 183 422 184 
<< m2 >>
rect 421 183 422 184 
<< m2c >>
rect 421 183 422 184 
<< m1 >>
rect 421 183 422 184 
<< m2 >>
rect 421 183 422 184 
<< m1 >>
rect 423 183 424 184 
<< m2 >>
rect 423 183 424 184 
<< m2c >>
rect 423 183 424 184 
<< m1 >>
rect 423 183 424 184 
<< m2 >>
rect 423 183 424 184 
<< m2 >>
rect 426 183 427 184 
<< m2 >>
rect 433 183 434 184 
<< m2 >>
rect 456 183 457 184 
<< m1 >>
rect 478 183 479 184 
<< m2 >>
rect 478 183 479 184 
<< m1 >>
rect 28 184 29 185 
<< m1 >>
rect 64 184 65 185 
<< m2 >>
rect 97 184 98 185 
<< m1 >>
rect 98 184 99 185 
<< m1 >>
rect 100 184 101 185 
<< m1 >>
rect 118 184 119 185 
<< m1 >>
rect 120 184 121 185 
<< m2 >>
rect 120 184 121 185 
<< m1 >>
rect 121 184 122 185 
<< m2 >>
rect 121 184 122 185 
<< m1 >>
rect 122 184 123 185 
<< m2 >>
rect 122 184 123 185 
<< m1 >>
rect 123 184 124 185 
<< m1 >>
rect 124 184 125 185 
<< m1 >>
rect 125 184 126 185 
<< m2 >>
rect 125 184 126 185 
<< m2c >>
rect 125 184 126 185 
<< m1 >>
rect 125 184 126 185 
<< m2 >>
rect 125 184 126 185 
<< m2 >>
rect 126 184 127 185 
<< m1 >>
rect 127 184 128 185 
<< m2 >>
rect 127 184 128 185 
<< m2 >>
rect 128 184 129 185 
<< m1 >>
rect 129 184 130 185 
<< m2 >>
rect 129 184 130 185 
<< m1 >>
rect 130 184 131 185 
<< m2 >>
rect 130 184 131 185 
<< m1 >>
rect 131 184 132 185 
<< m2 >>
rect 131 184 132 185 
<< m1 >>
rect 132 184 133 185 
<< m2 >>
rect 132 184 133 185 
<< m1 >>
rect 133 184 134 185 
<< m2 >>
rect 133 184 134 185 
<< m1 >>
rect 134 184 135 185 
<< m2 >>
rect 134 184 135 185 
<< m1 >>
rect 135 184 136 185 
<< m2 >>
rect 135 184 136 185 
<< m1 >>
rect 136 184 137 185 
<< m2 >>
rect 136 184 137 185 
<< m1 >>
rect 137 184 138 185 
<< m2 >>
rect 137 184 138 185 
<< m1 >>
rect 138 184 139 185 
<< m2 >>
rect 138 184 139 185 
<< m1 >>
rect 139 184 140 185 
<< m2 >>
rect 139 184 140 185 
<< m1 >>
rect 140 184 141 185 
<< m2 >>
rect 140 184 141 185 
<< m1 >>
rect 141 184 142 185 
<< m1 >>
rect 142 184 143 185 
<< m1 >>
rect 143 184 144 185 
<< m1 >>
rect 144 184 145 185 
<< m1 >>
rect 145 184 146 185 
<< m1 >>
rect 146 184 147 185 
<< m1 >>
rect 147 184 148 185 
<< m1 >>
rect 148 184 149 185 
<< m1 >>
rect 149 184 150 185 
<< m1 >>
rect 150 184 151 185 
<< m1 >>
rect 151 184 152 185 
<< m1 >>
rect 152 184 153 185 
<< m1 >>
rect 153 184 154 185 
<< m1 >>
rect 154 184 155 185 
<< m1 >>
rect 155 184 156 185 
<< m1 >>
rect 156 184 157 185 
<< m1 >>
rect 157 184 158 185 
<< m1 >>
rect 158 184 159 185 
<< m1 >>
rect 159 184 160 185 
<< m1 >>
rect 160 184 161 185 
<< m1 >>
rect 161 184 162 185 
<< m1 >>
rect 162 184 163 185 
<< m1 >>
rect 163 184 164 185 
<< m2 >>
rect 163 184 164 185 
<< m1 >>
rect 164 184 165 185 
<< m1 >>
rect 165 184 166 185 
<< m1 >>
rect 166 184 167 185 
<< m1 >>
rect 167 184 168 185 
<< m1 >>
rect 168 184 169 185 
<< m1 >>
rect 169 184 170 185 
<< m1 >>
rect 170 184 171 185 
<< m1 >>
rect 171 184 172 185 
<< m1 >>
rect 172 184 173 185 
<< m1 >>
rect 173 184 174 185 
<< m1 >>
rect 174 184 175 185 
<< m1 >>
rect 175 184 176 185 
<< m1 >>
rect 176 184 177 185 
<< m2 >>
rect 176 184 177 185 
<< m2c >>
rect 176 184 177 185 
<< m1 >>
rect 176 184 177 185 
<< m2 >>
rect 176 184 177 185 
<< m2 >>
rect 177 184 178 185 
<< m1 >>
rect 178 184 179 185 
<< m1 >>
rect 179 184 180 185 
<< m1 >>
rect 180 184 181 185 
<< m1 >>
rect 181 184 182 185 
<< m1 >>
rect 182 184 183 185 
<< m1 >>
rect 183 184 184 185 
<< m2 >>
rect 183 184 184 185 
<< m2c >>
rect 183 184 184 185 
<< m1 >>
rect 183 184 184 185 
<< m2 >>
rect 183 184 184 185 
<< m2 >>
rect 184 184 185 185 
<< m1 >>
rect 185 184 186 185 
<< m2 >>
rect 185 184 186 185 
<< m2 >>
rect 186 184 187 185 
<< m1 >>
rect 187 184 188 185 
<< m2 >>
rect 187 184 188 185 
<< m2c >>
rect 187 184 188 185 
<< m1 >>
rect 187 184 188 185 
<< m2 >>
rect 187 184 188 185 
<< m1 >>
rect 188 184 189 185 
<< m1 >>
rect 189 184 190 185 
<< m2 >>
rect 189 184 190 185 
<< m1 >>
rect 190 184 191 185 
<< m1 >>
rect 191 184 192 185 
<< m1 >>
rect 192 184 193 185 
<< m2 >>
rect 192 184 193 185 
<< m1 >>
rect 193 184 194 185 
<< m1 >>
rect 194 184 195 185 
<< m1 >>
rect 195 184 196 185 
<< m1 >>
rect 196 184 197 185 
<< m1 >>
rect 197 184 198 185 
<< m1 >>
rect 198 184 199 185 
<< m1 >>
rect 199 184 200 185 
<< m1 >>
rect 214 184 215 185 
<< m1 >>
rect 217 184 218 185 
<< m1 >>
rect 218 184 219 185 
<< m1 >>
rect 219 184 220 185 
<< m1 >>
rect 220 184 221 185 
<< m1 >>
rect 221 184 222 185 
<< m2 >>
rect 221 184 222 185 
<< m1 >>
rect 222 184 223 185 
<< m1 >>
rect 223 184 224 185 
<< m1 >>
rect 224 184 225 185 
<< m1 >>
rect 225 184 226 185 
<< m1 >>
rect 226 184 227 185 
<< m2 >>
rect 226 184 227 185 
<< m1 >>
rect 227 184 228 185 
<< m1 >>
rect 228 184 229 185 
<< m1 >>
rect 229 184 230 185 
<< m1 >>
rect 230 184 231 185 
<< m1 >>
rect 231 184 232 185 
<< m2 >>
rect 231 184 232 185 
<< m1 >>
rect 232 184 233 185 
<< m1 >>
rect 233 184 234 185 
<< m2 >>
rect 233 184 234 185 
<< m2c >>
rect 233 184 234 185 
<< m1 >>
rect 233 184 234 185 
<< m2 >>
rect 233 184 234 185 
<< m2 >>
rect 234 184 235 185 
<< m1 >>
rect 235 184 236 185 
<< m2 >>
rect 235 184 236 185 
<< m2 >>
rect 236 184 237 185 
<< m1 >>
rect 237 184 238 185 
<< m2 >>
rect 237 184 238 185 
<< m2c >>
rect 237 184 238 185 
<< m1 >>
rect 237 184 238 185 
<< m2 >>
rect 237 184 238 185 
<< m1 >>
rect 240 184 241 185 
<< m2 >>
rect 240 184 241 185 
<< m2c >>
rect 240 184 241 185 
<< m1 >>
rect 240 184 241 185 
<< m2 >>
rect 240 184 241 185 
<< m2 >>
rect 241 184 242 185 
<< m1 >>
rect 242 184 243 185 
<< m2 >>
rect 242 184 243 185 
<< m2 >>
rect 243 184 244 185 
<< m1 >>
rect 244 184 245 185 
<< m2 >>
rect 244 184 245 185 
<< m1 >>
rect 253 184 254 185 
<< m2 >>
rect 253 184 254 185 
<< m1 >>
rect 278 184 279 185 
<< m1 >>
rect 280 184 281 185 
<< m2 >>
rect 280 184 281 185 
<< m1 >>
rect 289 184 290 185 
<< m1 >>
rect 290 184 291 185 
<< m1 >>
rect 291 184 292 185 
<< m1 >>
rect 292 184 293 185 
<< m1 >>
rect 293 184 294 185 
<< m1 >>
rect 294 184 295 185 
<< m1 >>
rect 295 184 296 185 
<< m1 >>
rect 296 184 297 185 
<< m1 >>
rect 297 184 298 185 
<< m1 >>
rect 298 184 299 185 
<< m1 >>
rect 299 184 300 185 
<< m1 >>
rect 300 184 301 185 
<< m2 >>
rect 300 184 301 185 
<< m1 >>
rect 301 184 302 185 
<< m2 >>
rect 301 184 302 185 
<< m1 >>
rect 302 184 303 185 
<< m2 >>
rect 302 184 303 185 
<< m1 >>
rect 303 184 304 185 
<< m2 >>
rect 303 184 304 185 
<< m1 >>
rect 304 184 305 185 
<< m2 >>
rect 304 184 305 185 
<< m1 >>
rect 305 184 306 185 
<< m2 >>
rect 305 184 306 185 
<< m1 >>
rect 306 184 307 185 
<< m2 >>
rect 306 184 307 185 
<< m1 >>
rect 307 184 308 185 
<< m2 >>
rect 307 184 308 185 
<< m1 >>
rect 308 184 309 185 
<< m2 >>
rect 308 184 309 185 
<< m1 >>
rect 309 184 310 185 
<< m2 >>
rect 309 184 310 185 
<< m1 >>
rect 310 184 311 185 
<< m2 >>
rect 310 184 311 185 
<< m1 >>
rect 311 184 312 185 
<< m2 >>
rect 311 184 312 185 
<< m1 >>
rect 312 184 313 185 
<< m2 >>
rect 312 184 313 185 
<< m1 >>
rect 313 184 314 185 
<< m2 >>
rect 313 184 314 185 
<< m1 >>
rect 314 184 315 185 
<< m2 >>
rect 314 184 315 185 
<< m1 >>
rect 315 184 316 185 
<< m2 >>
rect 315 184 316 185 
<< m1 >>
rect 316 184 317 185 
<< m2 >>
rect 316 184 317 185 
<< m1 >>
rect 317 184 318 185 
<< m2 >>
rect 317 184 318 185 
<< m1 >>
rect 318 184 319 185 
<< m2 >>
rect 318 184 319 185 
<< m1 >>
rect 319 184 320 185 
<< m2 >>
rect 319 184 320 185 
<< m1 >>
rect 320 184 321 185 
<< m2 >>
rect 320 184 321 185 
<< m1 >>
rect 321 184 322 185 
<< m2 >>
rect 321 184 322 185 
<< m1 >>
rect 322 184 323 185 
<< m1 >>
rect 323 184 324 185 
<< m2 >>
rect 323 184 324 185 
<< m2c >>
rect 323 184 324 185 
<< m1 >>
rect 323 184 324 185 
<< m2 >>
rect 323 184 324 185 
<< m2 >>
rect 324 184 325 185 
<< m1 >>
rect 325 184 326 185 
<< m2 >>
rect 325 184 326 185 
<< m2 >>
rect 326 184 327 185 
<< m1 >>
rect 327 184 328 185 
<< m2 >>
rect 327 184 328 185 
<< m2c >>
rect 327 184 328 185 
<< m1 >>
rect 327 184 328 185 
<< m2 >>
rect 327 184 328 185 
<< m1 >>
rect 328 184 329 185 
<< m1 >>
rect 329 184 330 185 
<< m2 >>
rect 329 184 330 185 
<< m1 >>
rect 330 184 331 185 
<< m2 >>
rect 330 184 331 185 
<< m1 >>
rect 331 184 332 185 
<< m2 >>
rect 331 184 332 185 
<< m1 >>
rect 332 184 333 185 
<< m2 >>
rect 332 184 333 185 
<< m1 >>
rect 333 184 334 185 
<< m2 >>
rect 333 184 334 185 
<< m1 >>
rect 334 184 335 185 
<< m2 >>
rect 334 184 335 185 
<< m1 >>
rect 335 184 336 185 
<< m2 >>
rect 335 184 336 185 
<< m1 >>
rect 336 184 337 185 
<< m2 >>
rect 336 184 337 185 
<< m1 >>
rect 337 184 338 185 
<< m2 >>
rect 337 184 338 185 
<< m1 >>
rect 338 184 339 185 
<< m2 >>
rect 338 184 339 185 
<< m1 >>
rect 339 184 340 185 
<< m2 >>
rect 339 184 340 185 
<< m1 >>
rect 340 184 341 185 
<< m2 >>
rect 340 184 341 185 
<< m2 >>
rect 341 184 342 185 
<< m2 >>
rect 342 184 343 185 
<< m1 >>
rect 343 184 344 185 
<< m2 >>
rect 343 184 344 185 
<< m2 >>
rect 344 184 345 185 
<< m1 >>
rect 345 184 346 185 
<< m2 >>
rect 345 184 346 185 
<< m2c >>
rect 345 184 346 185 
<< m1 >>
rect 345 184 346 185 
<< m2 >>
rect 345 184 346 185 
<< m1 >>
rect 346 184 347 185 
<< m1 >>
rect 347 184 348 185 
<< m1 >>
rect 348 184 349 185 
<< m2 >>
rect 348 184 349 185 
<< m1 >>
rect 349 184 350 185 
<< m1 >>
rect 350 184 351 185 
<< m1 >>
rect 351 184 352 185 
<< m1 >>
rect 352 184 353 185 
<< m1 >>
rect 353 184 354 185 
<< m1 >>
rect 354 184 355 185 
<< m2 >>
rect 354 184 355 185 
<< m1 >>
rect 355 184 356 185 
<< m1 >>
rect 356 184 357 185 
<< m2 >>
rect 356 184 357 185 
<< m2c >>
rect 356 184 357 185 
<< m1 >>
rect 356 184 357 185 
<< m2 >>
rect 356 184 357 185 
<< m2 >>
rect 357 184 358 185 
<< m1 >>
rect 358 184 359 185 
<< m2 >>
rect 358 184 359 185 
<< m1 >>
rect 359 184 360 185 
<< m2 >>
rect 359 184 360 185 
<< m1 >>
rect 360 184 361 185 
<< m2 >>
rect 360 184 361 185 
<< m1 >>
rect 361 184 362 185 
<< m2 >>
rect 361 184 362 185 
<< m1 >>
rect 362 184 363 185 
<< m2 >>
rect 362 184 363 185 
<< m1 >>
rect 363 184 364 185 
<< m2 >>
rect 363 184 364 185 
<< m1 >>
rect 364 184 365 185 
<< m2 >>
rect 364 184 365 185 
<< m1 >>
rect 365 184 366 185 
<< m2 >>
rect 365 184 366 185 
<< m1 >>
rect 366 184 367 185 
<< m2 >>
rect 366 184 367 185 
<< m1 >>
rect 367 184 368 185 
<< m2 >>
rect 367 184 368 185 
<< m1 >>
rect 368 184 369 185 
<< m2 >>
rect 368 184 369 185 
<< m1 >>
rect 369 184 370 185 
<< m2 >>
rect 369 184 370 185 
<< m1 >>
rect 370 184 371 185 
<< m2 >>
rect 370 184 371 185 
<< m1 >>
rect 371 184 372 185 
<< m2 >>
rect 371 184 372 185 
<< m1 >>
rect 372 184 373 185 
<< m2 >>
rect 372 184 373 185 
<< m1 >>
rect 373 184 374 185 
<< m2 >>
rect 373 184 374 185 
<< m1 >>
rect 374 184 375 185 
<< m2 >>
rect 374 184 375 185 
<< m1 >>
rect 375 184 376 185 
<< m2 >>
rect 375 184 376 185 
<< m1 >>
rect 376 184 377 185 
<< m2 >>
rect 376 184 377 185 
<< m1 >>
rect 377 184 378 185 
<< m2 >>
rect 377 184 378 185 
<< m2 >>
rect 378 184 379 185 
<< m1 >>
rect 379 184 380 185 
<< m2 >>
rect 379 184 380 185 
<< m2 >>
rect 380 184 381 185 
<< m1 >>
rect 381 184 382 185 
<< m2 >>
rect 381 184 382 185 
<< m2c >>
rect 381 184 382 185 
<< m1 >>
rect 381 184 382 185 
<< m2 >>
rect 381 184 382 185 
<< m1 >>
rect 382 184 383 185 
<< m1 >>
rect 383 184 384 185 
<< m2 >>
rect 383 184 384 185 
<< m1 >>
rect 384 184 385 185 
<< m2 >>
rect 384 184 385 185 
<< m1 >>
rect 385 184 386 185 
<< m2 >>
rect 385 184 386 185 
<< m1 >>
rect 386 184 387 185 
<< m2 >>
rect 386 184 387 185 
<< m1 >>
rect 387 184 388 185 
<< m2 >>
rect 387 184 388 185 
<< m1 >>
rect 388 184 389 185 
<< m2 >>
rect 388 184 389 185 
<< m1 >>
rect 389 184 390 185 
<< m2 >>
rect 389 184 390 185 
<< m1 >>
rect 390 184 391 185 
<< m2 >>
rect 390 184 391 185 
<< m1 >>
rect 391 184 392 185 
<< m2 >>
rect 391 184 392 185 
<< m1 >>
rect 392 184 393 185 
<< m2 >>
rect 392 184 393 185 
<< m1 >>
rect 393 184 394 185 
<< m2 >>
rect 393 184 394 185 
<< m1 >>
rect 394 184 395 185 
<< m2 >>
rect 394 184 395 185 
<< m1 >>
rect 395 184 396 185 
<< m2 >>
rect 395 184 396 185 
<< m1 >>
rect 396 184 397 185 
<< m2 >>
rect 396 184 397 185 
<< m1 >>
rect 397 184 398 185 
<< m1 >>
rect 398 184 399 185 
<< m1 >>
rect 399 184 400 185 
<< m1 >>
rect 400 184 401 185 
<< m2 >>
rect 400 184 401 185 
<< m2c >>
rect 400 184 401 185 
<< m1 >>
rect 400 184 401 185 
<< m2 >>
rect 400 184 401 185 
<< m2 >>
rect 401 184 402 185 
<< m1 >>
rect 402 184 403 185 
<< m2 >>
rect 402 184 403 185 
<< m2 >>
rect 403 184 404 185 
<< m1 >>
rect 404 184 405 185 
<< m2 >>
rect 404 184 405 185 
<< m2c >>
rect 404 184 405 185 
<< m1 >>
rect 404 184 405 185 
<< m2 >>
rect 404 184 405 185 
<< m2 >>
rect 405 184 406 185 
<< m1 >>
rect 406 184 407 185 
<< m2 >>
rect 406 184 407 185 
<< m2 >>
rect 407 184 408 185 
<< m1 >>
rect 408 184 409 185 
<< m2 >>
rect 408 184 409 185 
<< m2c >>
rect 408 184 409 185 
<< m1 >>
rect 408 184 409 185 
<< m2 >>
rect 408 184 409 185 
<< m1 >>
rect 409 184 410 185 
<< m1 >>
rect 410 184 411 185 
<< m2 >>
rect 410 184 411 185 
<< m1 >>
rect 411 184 412 185 
<< m1 >>
rect 412 184 413 185 
<< m1 >>
rect 413 184 414 185 
<< m2 >>
rect 413 184 414 185 
<< m2c >>
rect 413 184 414 185 
<< m1 >>
rect 413 184 414 185 
<< m2 >>
rect 413 184 414 185 
<< m2 >>
rect 414 184 415 185 
<< m1 >>
rect 415 184 416 185 
<< m2 >>
rect 415 184 416 185 
<< m2 >>
rect 416 184 417 185 
<< m1 >>
rect 417 184 418 185 
<< m2 >>
rect 417 184 418 185 
<< m2c >>
rect 417 184 418 185 
<< m1 >>
rect 417 184 418 185 
<< m2 >>
rect 417 184 418 185 
<< m1 >>
rect 419 184 420 185 
<< m1 >>
rect 421 184 422 185 
<< m1 >>
rect 423 184 424 185 
<< m2 >>
rect 426 184 427 185 
<< m1 >>
rect 427 184 428 185 
<< m1 >>
rect 428 184 429 185 
<< m1 >>
rect 429 184 430 185 
<< m1 >>
rect 430 184 431 185 
<< m1 >>
rect 431 184 432 185 
<< m1 >>
rect 432 184 433 185 
<< m1 >>
rect 433 184 434 185 
<< m2 >>
rect 433 184 434 185 
<< m1 >>
rect 434 184 435 185 
<< m1 >>
rect 435 184 436 185 
<< m1 >>
rect 436 184 437 185 
<< m1 >>
rect 437 184 438 185 
<< m1 >>
rect 438 184 439 185 
<< m1 >>
rect 439 184 440 185 
<< m1 >>
rect 440 184 441 185 
<< m1 >>
rect 441 184 442 185 
<< m1 >>
rect 442 184 443 185 
<< m1 >>
rect 443 184 444 185 
<< m1 >>
rect 444 184 445 185 
<< m1 >>
rect 445 184 446 185 
<< m1 >>
rect 446 184 447 185 
<< m1 >>
rect 447 184 448 185 
<< m1 >>
rect 448 184 449 185 
<< m1 >>
rect 449 184 450 185 
<< m1 >>
rect 450 184 451 185 
<< m1 >>
rect 451 184 452 185 
<< m1 >>
rect 452 184 453 185 
<< m1 >>
rect 453 184 454 185 
<< m1 >>
rect 454 184 455 185 
<< m1 >>
rect 455 184 456 185 
<< m1 >>
rect 456 184 457 185 
<< m2 >>
rect 456 184 457 185 
<< m1 >>
rect 457 184 458 185 
<< m1 >>
rect 458 184 459 185 
<< m1 >>
rect 459 184 460 185 
<< m1 >>
rect 460 184 461 185 
<< m1 >>
rect 461 184 462 185 
<< m1 >>
rect 462 184 463 185 
<< m1 >>
rect 463 184 464 185 
<< m1 >>
rect 464 184 465 185 
<< m1 >>
rect 465 184 466 185 
<< m1 >>
rect 466 184 467 185 
<< m1 >>
rect 467 184 468 185 
<< m1 >>
rect 468 184 469 185 
<< m1 >>
rect 469 184 470 185 
<< m1 >>
rect 470 184 471 185 
<< m1 >>
rect 471 184 472 185 
<< m1 >>
rect 472 184 473 185 
<< m1 >>
rect 473 184 474 185 
<< m1 >>
rect 474 184 475 185 
<< m1 >>
rect 475 184 476 185 
<< m1 >>
rect 476 184 477 185 
<< m1 >>
rect 477 184 478 185 
<< m1 >>
rect 478 184 479 185 
<< m2 >>
rect 478 184 479 185 
<< m1 >>
rect 28 185 29 186 
<< m1 >>
rect 64 185 65 186 
<< m2 >>
rect 97 185 98 186 
<< m1 >>
rect 98 185 99 186 
<< m1 >>
rect 100 185 101 186 
<< m1 >>
rect 118 185 119 186 
<< m2 >>
rect 118 185 119 186 
<< m2c >>
rect 118 185 119 186 
<< m1 >>
rect 118 185 119 186 
<< m2 >>
rect 118 185 119 186 
<< m1 >>
rect 127 185 128 186 
<< m2 >>
rect 140 185 141 186 
<< m2 >>
rect 163 185 164 186 
<< m2 >>
rect 177 185 178 186 
<< m1 >>
rect 178 185 179 186 
<< m1 >>
rect 185 185 186 186 
<< m2 >>
rect 189 185 190 186 
<< m2 >>
rect 192 185 193 186 
<< m2 >>
rect 193 185 194 186 
<< m2 >>
rect 194 185 195 186 
<< m2 >>
rect 195 185 196 186 
<< m2 >>
rect 196 185 197 186 
<< m2 >>
rect 197 185 198 186 
<< m2 >>
rect 198 185 199 186 
<< m2 >>
rect 199 185 200 186 
<< m2 >>
rect 200 185 201 186 
<< m1 >>
rect 201 185 202 186 
<< m2 >>
rect 201 185 202 186 
<< m2c >>
rect 201 185 202 186 
<< m1 >>
rect 201 185 202 186 
<< m2 >>
rect 201 185 202 186 
<< m1 >>
rect 202 185 203 186 
<< m1 >>
rect 203 185 204 186 
<< m1 >>
rect 204 185 205 186 
<< m1 >>
rect 205 185 206 186 
<< m1 >>
rect 206 185 207 186 
<< m1 >>
rect 207 185 208 186 
<< m1 >>
rect 208 185 209 186 
<< m1 >>
rect 209 185 210 186 
<< m1 >>
rect 210 185 211 186 
<< m1 >>
rect 211 185 212 186 
<< m1 >>
rect 212 185 213 186 
<< m1 >>
rect 213 185 214 186 
<< m1 >>
rect 214 185 215 186 
<< m2 >>
rect 221 185 222 186 
<< m2 >>
rect 226 185 227 186 
<< m2 >>
rect 231 185 232 186 
<< m1 >>
rect 235 185 236 186 
<< m1 >>
rect 237 185 238 186 
<< m1 >>
rect 240 185 241 186 
<< m1 >>
rect 242 185 243 186 
<< m1 >>
rect 244 185 245 186 
<< m1 >>
rect 246 185 247 186 
<< m2 >>
rect 246 185 247 186 
<< m2c >>
rect 246 185 247 186 
<< m1 >>
rect 246 185 247 186 
<< m2 >>
rect 246 185 247 186 
<< m1 >>
rect 247 185 248 186 
<< m1 >>
rect 248 185 249 186 
<< m1 >>
rect 249 185 250 186 
<< m1 >>
rect 250 185 251 186 
<< m1 >>
rect 251 185 252 186 
<< m1 >>
rect 252 185 253 186 
<< m1 >>
rect 253 185 254 186 
<< m2 >>
rect 253 185 254 186 
<< m1 >>
rect 278 185 279 186 
<< m2 >>
rect 278 185 279 186 
<< m2c >>
rect 278 185 279 186 
<< m1 >>
rect 278 185 279 186 
<< m2 >>
rect 278 185 279 186 
<< m1 >>
rect 280 185 281 186 
<< m2 >>
rect 280 185 281 186 
<< m1 >>
rect 281 185 282 186 
<< m1 >>
rect 282 185 283 186 
<< m1 >>
rect 283 185 284 186 
<< m1 >>
rect 284 185 285 186 
<< m1 >>
rect 285 185 286 186 
<< m1 >>
rect 286 185 287 186 
<< m1 >>
rect 287 185 288 186 
<< m2 >>
rect 287 185 288 186 
<< m2c >>
rect 287 185 288 186 
<< m1 >>
rect 287 185 288 186 
<< m2 >>
rect 287 185 288 186 
<< m2 >>
rect 288 185 289 186 
<< m2 >>
rect 289 185 290 186 
<< m2 >>
rect 290 185 291 186 
<< m2 >>
rect 291 185 292 186 
<< m2 >>
rect 292 185 293 186 
<< m2 >>
rect 293 185 294 186 
<< m2 >>
rect 294 185 295 186 
<< m2 >>
rect 295 185 296 186 
<< m2 >>
rect 296 185 297 186 
<< m2 >>
rect 297 185 298 186 
<< m2 >>
rect 298 185 299 186 
<< m2 >>
rect 300 185 301 186 
<< m1 >>
rect 325 185 326 186 
<< m1 >>
rect 340 185 341 186 
<< m1 >>
rect 343 185 344 186 
<< m2 >>
rect 348 185 349 186 
<< m2 >>
rect 354 185 355 186 
<< m1 >>
rect 358 185 359 186 
<< m1 >>
rect 379 185 380 186 
<< m2 >>
rect 396 185 397 186 
<< m1 >>
rect 402 185 403 186 
<< m1 >>
rect 406 185 407 186 
<< m2 >>
rect 410 185 411 186 
<< m1 >>
rect 415 185 416 186 
<< m1 >>
rect 417 185 418 186 
<< m1 >>
rect 419 185 420 186 
<< m1 >>
rect 421 185 422 186 
<< m1 >>
rect 423 185 424 186 
<< m2 >>
rect 426 185 427 186 
<< m1 >>
rect 427 185 428 186 
<< m2 >>
rect 433 185 434 186 
<< m2 >>
rect 456 185 457 186 
<< m2 >>
rect 478 185 479 186 
<< m1 >>
rect 28 186 29 187 
<< m1 >>
rect 64 186 65 187 
<< m2 >>
rect 97 186 98 187 
<< m1 >>
rect 98 186 99 187 
<< m1 >>
rect 100 186 101 187 
<< m2 >>
rect 118 186 119 187 
<< m1 >>
rect 127 186 128 187 
<< m2 >>
rect 140 186 141 187 
<< m1 >>
rect 163 186 164 187 
<< m2 >>
rect 163 186 164 187 
<< m2c >>
rect 163 186 164 187 
<< m1 >>
rect 163 186 164 187 
<< m2 >>
rect 163 186 164 187 
<< m2 >>
rect 177 186 178 187 
<< m1 >>
rect 178 186 179 187 
<< m2 >>
rect 178 186 179 187 
<< m2 >>
rect 179 186 180 187 
<< m1 >>
rect 180 186 181 187 
<< m2 >>
rect 180 186 181 187 
<< m2c >>
rect 180 186 181 187 
<< m1 >>
rect 180 186 181 187 
<< m2 >>
rect 180 186 181 187 
<< m1 >>
rect 181 186 182 187 
<< m1 >>
rect 182 186 183 187 
<< m1 >>
rect 183 186 184 187 
<< m2 >>
rect 183 186 184 187 
<< m2c >>
rect 183 186 184 187 
<< m1 >>
rect 183 186 184 187 
<< m2 >>
rect 183 186 184 187 
<< m2 >>
rect 184 186 185 187 
<< m1 >>
rect 185 186 186 187 
<< m2 >>
rect 185 186 186 187 
<< m2 >>
rect 186 186 187 187 
<< m1 >>
rect 187 186 188 187 
<< m2 >>
rect 187 186 188 187 
<< m2c >>
rect 187 186 188 187 
<< m1 >>
rect 187 186 188 187 
<< m2 >>
rect 187 186 188 187 
<< m1 >>
rect 189 186 190 187 
<< m2 >>
rect 189 186 190 187 
<< m2c >>
rect 189 186 190 187 
<< m1 >>
rect 189 186 190 187 
<< m2 >>
rect 189 186 190 187 
<< m1 >>
rect 221 186 222 187 
<< m2 >>
rect 221 186 222 187 
<< m2c >>
rect 221 186 222 187 
<< m1 >>
rect 221 186 222 187 
<< m2 >>
rect 221 186 222 187 
<< m1 >>
rect 226 186 227 187 
<< m2 >>
rect 226 186 227 187 
<< m2c >>
rect 226 186 227 187 
<< m1 >>
rect 226 186 227 187 
<< m2 >>
rect 226 186 227 187 
<< m1 >>
rect 231 186 232 187 
<< m2 >>
rect 231 186 232 187 
<< m2c >>
rect 231 186 232 187 
<< m1 >>
rect 231 186 232 187 
<< m2 >>
rect 231 186 232 187 
<< m1 >>
rect 233 186 234 187 
<< m2 >>
rect 233 186 234 187 
<< m2c >>
rect 233 186 234 187 
<< m1 >>
rect 233 186 234 187 
<< m2 >>
rect 233 186 234 187 
<< m2 >>
rect 234 186 235 187 
<< m1 >>
rect 235 186 236 187 
<< m2 >>
rect 235 186 236 187 
<< m2 >>
rect 236 186 237 187 
<< m1 >>
rect 237 186 238 187 
<< m2 >>
rect 237 186 238 187 
<< m2 >>
rect 238 186 239 187 
<< m1 >>
rect 239 186 240 187 
<< m2 >>
rect 239 186 240 187 
<< m2c >>
rect 239 186 240 187 
<< m1 >>
rect 239 186 240 187 
<< m2 >>
rect 239 186 240 187 
<< m1 >>
rect 240 186 241 187 
<< m1 >>
rect 242 186 243 187 
<< m1 >>
rect 244 186 245 187 
<< m2 >>
rect 246 186 247 187 
<< m2 >>
rect 253 186 254 187 
<< m2 >>
rect 278 186 279 187 
<< m2 >>
rect 280 186 281 187 
<< m2 >>
rect 298 186 299 187 
<< m2 >>
rect 300 186 301 187 
<< m1 >>
rect 325 186 326 187 
<< m1 >>
rect 334 186 335 187 
<< m1 >>
rect 335 186 336 187 
<< m1 >>
rect 336 186 337 187 
<< m1 >>
rect 337 186 338 187 
<< m1 >>
rect 338 186 339 187 
<< m2 >>
rect 338 186 339 187 
<< m2c >>
rect 338 186 339 187 
<< m1 >>
rect 338 186 339 187 
<< m2 >>
rect 338 186 339 187 
<< m2 >>
rect 339 186 340 187 
<< m1 >>
rect 340 186 341 187 
<< m2 >>
rect 340 186 341 187 
<< m2 >>
rect 341 186 342 187 
<< m2 >>
rect 342 186 343 187 
<< m1 >>
rect 343 186 344 187 
<< m2 >>
rect 343 186 344 187 
<< m2 >>
rect 344 186 345 187 
<< m1 >>
rect 345 186 346 187 
<< m2 >>
rect 345 186 346 187 
<< m2c >>
rect 345 186 346 187 
<< m1 >>
rect 345 186 346 187 
<< m2 >>
rect 345 186 346 187 
<< m1 >>
rect 346 186 347 187 
<< m1 >>
rect 347 186 348 187 
<< m1 >>
rect 348 186 349 187 
<< m2 >>
rect 348 186 349 187 
<< m1 >>
rect 349 186 350 187 
<< m1 >>
rect 350 186 351 187 
<< m2 >>
rect 350 186 351 187 
<< m2c >>
rect 350 186 351 187 
<< m1 >>
rect 350 186 351 187 
<< m2 >>
rect 350 186 351 187 
<< m2 >>
rect 351 186 352 187 
<< m2 >>
rect 352 186 353 187 
<< m2 >>
rect 353 186 354 187 
<< m2 >>
rect 354 186 355 187 
<< m1 >>
rect 358 186 359 187 
<< m1 >>
rect 379 186 380 187 
<< m1 >>
rect 396 186 397 187 
<< m2 >>
rect 396 186 397 187 
<< m2c >>
rect 396 186 397 187 
<< m1 >>
rect 396 186 397 187 
<< m2 >>
rect 396 186 397 187 
<< m1 >>
rect 402 186 403 187 
<< m1 >>
rect 406 186 407 187 
<< m1 >>
rect 410 186 411 187 
<< m2 >>
rect 410 186 411 187 
<< m2c >>
rect 410 186 411 187 
<< m1 >>
rect 410 186 411 187 
<< m2 >>
rect 410 186 411 187 
<< m1 >>
rect 411 186 412 187 
<< m1 >>
rect 412 186 413 187 
<< m1 >>
rect 413 186 414 187 
<< m2 >>
rect 413 186 414 187 
<< m2c >>
rect 413 186 414 187 
<< m1 >>
rect 413 186 414 187 
<< m2 >>
rect 413 186 414 187 
<< m2 >>
rect 414 186 415 187 
<< m1 >>
rect 415 186 416 187 
<< m2 >>
rect 415 186 416 187 
<< m2 >>
rect 416 186 417 187 
<< m1 >>
rect 417 186 418 187 
<< m2 >>
rect 417 186 418 187 
<< m2 >>
rect 418 186 419 187 
<< m1 >>
rect 419 186 420 187 
<< m2 >>
rect 419 186 420 187 
<< m2 >>
rect 420 186 421 187 
<< m1 >>
rect 421 186 422 187 
<< m2 >>
rect 421 186 422 187 
<< m2c >>
rect 421 186 422 187 
<< m1 >>
rect 421 186 422 187 
<< m2 >>
rect 421 186 422 187 
<< m1 >>
rect 423 186 424 187 
<< m2 >>
rect 426 186 427 187 
<< m1 >>
rect 427 186 428 187 
<< m2 >>
rect 427 186 428 187 
<< m2 >>
rect 428 186 429 187 
<< m1 >>
rect 429 186 430 187 
<< m2 >>
rect 429 186 430 187 
<< m2c >>
rect 429 186 430 187 
<< m1 >>
rect 429 186 430 187 
<< m2 >>
rect 429 186 430 187 
<< m1 >>
rect 430 186 431 187 
<< m1 >>
rect 431 186 432 187 
<< m1 >>
rect 432 186 433 187 
<< m1 >>
rect 433 186 434 187 
<< m2 >>
rect 433 186 434 187 
<< m1 >>
rect 456 186 457 187 
<< m2 >>
rect 456 186 457 187 
<< m2c >>
rect 456 186 457 187 
<< m1 >>
rect 456 186 457 187 
<< m2 >>
rect 456 186 457 187 
<< m1 >>
rect 478 186 479 187 
<< m2 >>
rect 478 186 479 187 
<< m2c >>
rect 478 186 479 187 
<< m1 >>
rect 478 186 479 187 
<< m2 >>
rect 478 186 479 187 
<< m1 >>
rect 28 187 29 188 
<< m1 >>
rect 64 187 65 188 
<< m2 >>
rect 97 187 98 188 
<< m1 >>
rect 98 187 99 188 
<< m1 >>
rect 100 187 101 188 
<< m1 >>
rect 101 187 102 188 
<< m1 >>
rect 102 187 103 188 
<< m1 >>
rect 103 187 104 188 
<< m1 >>
rect 104 187 105 188 
<< m1 >>
rect 105 187 106 188 
<< m1 >>
rect 106 187 107 188 
<< m1 >>
rect 107 187 108 188 
<< m1 >>
rect 108 187 109 188 
<< m1 >>
rect 109 187 110 188 
<< m1 >>
rect 110 187 111 188 
<< m1 >>
rect 111 187 112 188 
<< m1 >>
rect 112 187 113 188 
<< m1 >>
rect 113 187 114 188 
<< m1 >>
rect 114 187 115 188 
<< m1 >>
rect 115 187 116 188 
<< m1 >>
rect 116 187 117 188 
<< m1 >>
rect 117 187 118 188 
<< m1 >>
rect 118 187 119 188 
<< m2 >>
rect 118 187 119 188 
<< m1 >>
rect 119 187 120 188 
<< m1 >>
rect 120 187 121 188 
<< m1 >>
rect 121 187 122 188 
<< m1 >>
rect 122 187 123 188 
<< m1 >>
rect 123 187 124 188 
<< m1 >>
rect 124 187 125 188 
<< m1 >>
rect 125 187 126 188 
<< m2 >>
rect 125 187 126 188 
<< m2c >>
rect 125 187 126 188 
<< m1 >>
rect 125 187 126 188 
<< m2 >>
rect 125 187 126 188 
<< m2 >>
rect 126 187 127 188 
<< m1 >>
rect 127 187 128 188 
<< m2 >>
rect 127 187 128 188 
<< m2 >>
rect 128 187 129 188 
<< m1 >>
rect 129 187 130 188 
<< m2 >>
rect 129 187 130 188 
<< m2c >>
rect 129 187 130 188 
<< m1 >>
rect 129 187 130 188 
<< m2 >>
rect 129 187 130 188 
<< m1 >>
rect 130 187 131 188 
<< m1 >>
rect 131 187 132 188 
<< m1 >>
rect 132 187 133 188 
<< m1 >>
rect 133 187 134 188 
<< m1 >>
rect 134 187 135 188 
<< m1 >>
rect 135 187 136 188 
<< m1 >>
rect 136 187 137 188 
<< m1 >>
rect 137 187 138 188 
<< m1 >>
rect 138 187 139 188 
<< m1 >>
rect 139 187 140 188 
<< m1 >>
rect 140 187 141 188 
<< m2 >>
rect 140 187 141 188 
<< m1 >>
rect 141 187 142 188 
<< m1 >>
rect 142 187 143 188 
<< m1 >>
rect 143 187 144 188 
<< m1 >>
rect 144 187 145 188 
<< m1 >>
rect 145 187 146 188 
<< m1 >>
rect 146 187 147 188 
<< m1 >>
rect 147 187 148 188 
<< m1 >>
rect 148 187 149 188 
<< m1 >>
rect 149 187 150 188 
<< m1 >>
rect 150 187 151 188 
<< m1 >>
rect 151 187 152 188 
<< m1 >>
rect 152 187 153 188 
<< m1 >>
rect 153 187 154 188 
<< m1 >>
rect 154 187 155 188 
<< m1 >>
rect 163 187 164 188 
<< m1 >>
rect 178 187 179 188 
<< m1 >>
rect 185 187 186 188 
<< m1 >>
rect 187 187 188 188 
<< m1 >>
rect 189 187 190 188 
<< m1 >>
rect 190 187 191 188 
<< m1 >>
rect 191 187 192 188 
<< m1 >>
rect 192 187 193 188 
<< m1 >>
rect 193 187 194 188 
<< m1 >>
rect 194 187 195 188 
<< m1 >>
rect 195 187 196 188 
<< m1 >>
rect 196 187 197 188 
<< m1 >>
rect 197 187 198 188 
<< m1 >>
rect 198 187 199 188 
<< m1 >>
rect 199 187 200 188 
<< m1 >>
rect 200 187 201 188 
<< m1 >>
rect 201 187 202 188 
<< m1 >>
rect 202 187 203 188 
<< m1 >>
rect 203 187 204 188 
<< m1 >>
rect 204 187 205 188 
<< m1 >>
rect 205 187 206 188 
<< m1 >>
rect 206 187 207 188 
<< m1 >>
rect 207 187 208 188 
<< m1 >>
rect 208 187 209 188 
<< m1 >>
rect 209 187 210 188 
<< m1 >>
rect 210 187 211 188 
<< m1 >>
rect 211 187 212 188 
<< m1 >>
rect 212 187 213 188 
<< m1 >>
rect 213 187 214 188 
<< m1 >>
rect 214 187 215 188 
<< m1 >>
rect 221 187 222 188 
<< m1 >>
rect 226 187 227 188 
<< m2 >>
rect 231 187 232 188 
<< m1 >>
rect 233 187 234 188 
<< m1 >>
rect 235 187 236 188 
<< m1 >>
rect 237 187 238 188 
<< m1 >>
rect 242 187 243 188 
<< m1 >>
rect 244 187 245 188 
<< m2 >>
rect 246 187 247 188 
<< m1 >>
rect 247 187 248 188 
<< m1 >>
rect 248 187 249 188 
<< m1 >>
rect 249 187 250 188 
<< m1 >>
rect 250 187 251 188 
<< m1 >>
rect 251 187 252 188 
<< m1 >>
rect 252 187 253 188 
<< m1 >>
rect 253 187 254 188 
<< m2 >>
rect 253 187 254 188 
<< m1 >>
rect 254 187 255 188 
<< m1 >>
rect 255 187 256 188 
<< m1 >>
rect 256 187 257 188 
<< m1 >>
rect 257 187 258 188 
<< m1 >>
rect 258 187 259 188 
<< m1 >>
rect 259 187 260 188 
<< m1 >>
rect 260 187 261 188 
<< m1 >>
rect 261 187 262 188 
<< m1 >>
rect 262 187 263 188 
<< m1 >>
rect 263 187 264 188 
<< m1 >>
rect 264 187 265 188 
<< m1 >>
rect 265 187 266 188 
<< m1 >>
rect 266 187 267 188 
<< m1 >>
rect 267 187 268 188 
<< m1 >>
rect 268 187 269 188 
<< m1 >>
rect 269 187 270 188 
<< m1 >>
rect 270 187 271 188 
<< m1 >>
rect 271 187 272 188 
<< m1 >>
rect 272 187 273 188 
<< m1 >>
rect 273 187 274 188 
<< m1 >>
rect 274 187 275 188 
<< m1 >>
rect 275 187 276 188 
<< m1 >>
rect 276 187 277 188 
<< m1 >>
rect 277 187 278 188 
<< m1 >>
rect 278 187 279 188 
<< m2 >>
rect 278 187 279 188 
<< m1 >>
rect 279 187 280 188 
<< m1 >>
rect 280 187 281 188 
<< m2 >>
rect 280 187 281 188 
<< m1 >>
rect 281 187 282 188 
<< m2 >>
rect 281 187 282 188 
<< m1 >>
rect 282 187 283 188 
<< m2 >>
rect 282 187 283 188 
<< m1 >>
rect 283 187 284 188 
<< m2 >>
rect 283 187 284 188 
<< m1 >>
rect 284 187 285 188 
<< m2 >>
rect 284 187 285 188 
<< m1 >>
rect 285 187 286 188 
<< m2 >>
rect 285 187 286 188 
<< m1 >>
rect 286 187 287 188 
<< m2 >>
rect 286 187 287 188 
<< m1 >>
rect 287 187 288 188 
<< m2 >>
rect 287 187 288 188 
<< m1 >>
rect 288 187 289 188 
<< m2 >>
rect 288 187 289 188 
<< m1 >>
rect 289 187 290 188 
<< m2 >>
rect 289 187 290 188 
<< m1 >>
rect 290 187 291 188 
<< m2 >>
rect 290 187 291 188 
<< m1 >>
rect 291 187 292 188 
<< m2 >>
rect 291 187 292 188 
<< m1 >>
rect 292 187 293 188 
<< m2 >>
rect 292 187 293 188 
<< m1 >>
rect 293 187 294 188 
<< m2 >>
rect 293 187 294 188 
<< m1 >>
rect 294 187 295 188 
<< m2 >>
rect 294 187 295 188 
<< m1 >>
rect 295 187 296 188 
<< m2 >>
rect 295 187 296 188 
<< m1 >>
rect 296 187 297 188 
<< m1 >>
rect 297 187 298 188 
<< m1 >>
rect 298 187 299 188 
<< m2 >>
rect 298 187 299 188 
<< m1 >>
rect 299 187 300 188 
<< m1 >>
rect 300 187 301 188 
<< m2 >>
rect 300 187 301 188 
<< m1 >>
rect 301 187 302 188 
<< m1 >>
rect 302 187 303 188 
<< m1 >>
rect 303 187 304 188 
<< m1 >>
rect 304 187 305 188 
<< m1 >>
rect 305 187 306 188 
<< m1 >>
rect 306 187 307 188 
<< m1 >>
rect 307 187 308 188 
<< m1 >>
rect 308 187 309 188 
<< m1 >>
rect 309 187 310 188 
<< m1 >>
rect 310 187 311 188 
<< m1 >>
rect 311 187 312 188 
<< m1 >>
rect 312 187 313 188 
<< m1 >>
rect 313 187 314 188 
<< m1 >>
rect 314 187 315 188 
<< m1 >>
rect 315 187 316 188 
<< m1 >>
rect 316 187 317 188 
<< m1 >>
rect 317 187 318 188 
<< m1 >>
rect 318 187 319 188 
<< m1 >>
rect 319 187 320 188 
<< m1 >>
rect 320 187 321 188 
<< m1 >>
rect 321 187 322 188 
<< m1 >>
rect 322 187 323 188 
<< m1 >>
rect 323 187 324 188 
<< m1 >>
rect 324 187 325 188 
<< m1 >>
rect 325 187 326 188 
<< m1 >>
rect 334 187 335 188 
<< m1 >>
rect 340 187 341 188 
<< m1 >>
rect 343 187 344 188 
<< m2 >>
rect 348 187 349 188 
<< m1 >>
rect 352 187 353 188 
<< m1 >>
rect 353 187 354 188 
<< m1 >>
rect 354 187 355 188 
<< m1 >>
rect 355 187 356 188 
<< m1 >>
rect 356 187 357 188 
<< m2 >>
rect 356 187 357 188 
<< m2c >>
rect 356 187 357 188 
<< m1 >>
rect 356 187 357 188 
<< m2 >>
rect 356 187 357 188 
<< m2 >>
rect 357 187 358 188 
<< m1 >>
rect 358 187 359 188 
<< m2 >>
rect 358 187 359 188 
<< m2 >>
rect 359 187 360 188 
<< m1 >>
rect 360 187 361 188 
<< m2 >>
rect 360 187 361 188 
<< m2c >>
rect 360 187 361 188 
<< m1 >>
rect 360 187 361 188 
<< m2 >>
rect 360 187 361 188 
<< m1 >>
rect 361 187 362 188 
<< m1 >>
rect 362 187 363 188 
<< m1 >>
rect 363 187 364 188 
<< m1 >>
rect 364 187 365 188 
<< m1 >>
rect 365 187 366 188 
<< m1 >>
rect 366 187 367 188 
<< m1 >>
rect 367 187 368 188 
<< m1 >>
rect 368 187 369 188 
<< m1 >>
rect 369 187 370 188 
<< m1 >>
rect 370 187 371 188 
<< m1 >>
rect 371 187 372 188 
<< m1 >>
rect 372 187 373 188 
<< m1 >>
rect 373 187 374 188 
<< m1 >>
rect 374 187 375 188 
<< m1 >>
rect 375 187 376 188 
<< m1 >>
rect 376 187 377 188 
<< m1 >>
rect 377 187 378 188 
<< m2 >>
rect 377 187 378 188 
<< m2c >>
rect 377 187 378 188 
<< m1 >>
rect 377 187 378 188 
<< m2 >>
rect 377 187 378 188 
<< m2 >>
rect 378 187 379 188 
<< m1 >>
rect 379 187 380 188 
<< m2 >>
rect 379 187 380 188 
<< m2 >>
rect 380 187 381 188 
<< m1 >>
rect 381 187 382 188 
<< m2 >>
rect 381 187 382 188 
<< m2c >>
rect 381 187 382 188 
<< m1 >>
rect 381 187 382 188 
<< m2 >>
rect 381 187 382 188 
<< m1 >>
rect 382 187 383 188 
<< m1 >>
rect 383 187 384 188 
<< m1 >>
rect 384 187 385 188 
<< m1 >>
rect 385 187 386 188 
<< m1 >>
rect 386 187 387 188 
<< m1 >>
rect 387 187 388 188 
<< m1 >>
rect 388 187 389 188 
<< m1 >>
rect 389 187 390 188 
<< m1 >>
rect 390 187 391 188 
<< m1 >>
rect 391 187 392 188 
<< m1 >>
rect 392 187 393 188 
<< m1 >>
rect 393 187 394 188 
<< m1 >>
rect 394 187 395 188 
<< m2 >>
rect 394 187 395 188 
<< m2c >>
rect 394 187 395 188 
<< m1 >>
rect 394 187 395 188 
<< m2 >>
rect 394 187 395 188 
<< m1 >>
rect 396 187 397 188 
<< m2 >>
rect 396 187 397 188 
<< m1 >>
rect 402 187 403 188 
<< m2 >>
rect 402 187 403 188 
<< m2c >>
rect 402 187 403 188 
<< m1 >>
rect 402 187 403 188 
<< m2 >>
rect 402 187 403 188 
<< m1 >>
rect 406 187 407 188 
<< m1 >>
rect 415 187 416 188 
<< m1 >>
rect 417 187 418 188 
<< m1 >>
rect 419 187 420 188 
<< m1 >>
rect 423 187 424 188 
<< m1 >>
rect 427 187 428 188 
<< m1 >>
rect 433 187 434 188 
<< m2 >>
rect 433 187 434 188 
<< m1 >>
rect 456 187 457 188 
<< m1 >>
rect 478 187 479 188 
<< m1 >>
rect 28 188 29 189 
<< m1 >>
rect 64 188 65 189 
<< m2 >>
rect 97 188 98 189 
<< m1 >>
rect 98 188 99 189 
<< m2 >>
rect 118 188 119 189 
<< m1 >>
rect 127 188 128 189 
<< m2 >>
rect 140 188 141 189 
<< m1 >>
rect 154 188 155 189 
<< m1 >>
rect 163 188 164 189 
<< m1 >>
rect 178 188 179 189 
<< m1 >>
rect 185 188 186 189 
<< m1 >>
rect 187 188 188 189 
<< m1 >>
rect 214 188 215 189 
<< m1 >>
rect 221 188 222 189 
<< m1 >>
rect 224 188 225 189 
<< m2 >>
rect 224 188 225 189 
<< m2c >>
rect 224 188 225 189 
<< m1 >>
rect 224 188 225 189 
<< m2 >>
rect 224 188 225 189 
<< m2 >>
rect 225 188 226 189 
<< m1 >>
rect 226 188 227 189 
<< m2 >>
rect 226 188 227 189 
<< m2 >>
rect 227 188 228 189 
<< m1 >>
rect 228 188 229 189 
<< m2 >>
rect 228 188 229 189 
<< m2c >>
rect 228 188 229 189 
<< m1 >>
rect 228 188 229 189 
<< m2 >>
rect 228 188 229 189 
<< m1 >>
rect 229 188 230 189 
<< m1 >>
rect 230 188 231 189 
<< m1 >>
rect 231 188 232 189 
<< m2 >>
rect 231 188 232 189 
<< m1 >>
rect 232 188 233 189 
<< m1 >>
rect 233 188 234 189 
<< m1 >>
rect 235 188 236 189 
<< m1 >>
rect 237 188 238 189 
<< m1 >>
rect 242 188 243 189 
<< m1 >>
rect 244 188 245 189 
<< m2 >>
rect 246 188 247 189 
<< m1 >>
rect 247 188 248 189 
<< m2 >>
rect 253 188 254 189 
<< m2 >>
rect 278 188 279 189 
<< m2 >>
rect 295 188 296 189 
<< m2 >>
rect 298 188 299 189 
<< m2 >>
rect 300 188 301 189 
<< m1 >>
rect 334 188 335 189 
<< m1 >>
rect 340 188 341 189 
<< m1 >>
rect 343 188 344 189 
<< m1 >>
rect 348 188 349 189 
<< m2 >>
rect 348 188 349 189 
<< m2c >>
rect 348 188 349 189 
<< m1 >>
rect 348 188 349 189 
<< m2 >>
rect 348 188 349 189 
<< m1 >>
rect 352 188 353 189 
<< m1 >>
rect 358 188 359 189 
<< m1 >>
rect 379 188 380 189 
<< m2 >>
rect 394 188 395 189 
<< m2 >>
rect 396 188 397 189 
<< m2 >>
rect 397 188 398 189 
<< m2 >>
rect 402 188 403 189 
<< m1 >>
rect 406 188 407 189 
<< m1 >>
rect 415 188 416 189 
<< m1 >>
rect 417 188 418 189 
<< m1 >>
rect 419 188 420 189 
<< m1 >>
rect 423 188 424 189 
<< m1 >>
rect 427 188 428 189 
<< m1 >>
rect 433 188 434 189 
<< m2 >>
rect 433 188 434 189 
<< m1 >>
rect 456 188 457 189 
<< m1 >>
rect 478 188 479 189 
<< m1 >>
rect 28 189 29 190 
<< m1 >>
rect 64 189 65 190 
<< m2 >>
rect 97 189 98 190 
<< m1 >>
rect 98 189 99 190 
<< m2 >>
rect 98 189 99 190 
<< m2 >>
rect 99 189 100 190 
<< m1 >>
rect 100 189 101 190 
<< m2 >>
rect 100 189 101 190 
<< m2c >>
rect 100 189 101 190 
<< m1 >>
rect 100 189 101 190 
<< m2 >>
rect 100 189 101 190 
<< m1 >>
rect 101 189 102 190 
<< m1 >>
rect 102 189 103 190 
<< m1 >>
rect 103 189 104 190 
<< m1 >>
rect 106 189 107 190 
<< m1 >>
rect 107 189 108 190 
<< m1 >>
rect 108 189 109 190 
<< m1 >>
rect 109 189 110 190 
<< m1 >>
rect 110 189 111 190 
<< m1 >>
rect 111 189 112 190 
<< m1 >>
rect 112 189 113 190 
<< m1 >>
rect 113 189 114 190 
<< m1 >>
rect 114 189 115 190 
<< m1 >>
rect 115 189 116 190 
<< m1 >>
rect 116 189 117 190 
<< m1 >>
rect 117 189 118 190 
<< m1 >>
rect 118 189 119 190 
<< m2 >>
rect 118 189 119 190 
<< m2c >>
rect 118 189 119 190 
<< m1 >>
rect 118 189 119 190 
<< m2 >>
rect 118 189 119 190 
<< m1 >>
rect 127 189 128 190 
<< m1 >>
rect 140 189 141 190 
<< m2 >>
rect 140 189 141 190 
<< m2c >>
rect 140 189 141 190 
<< m1 >>
rect 140 189 141 190 
<< m2 >>
rect 140 189 141 190 
<< m1 >>
rect 141 189 142 190 
<< m1 >>
rect 142 189 143 190 
<< m1 >>
rect 143 189 144 190 
<< m1 >>
rect 144 189 145 190 
<< m1 >>
rect 145 189 146 190 
<< m1 >>
rect 146 189 147 190 
<< m1 >>
rect 147 189 148 190 
<< m1 >>
rect 154 189 155 190 
<< m1 >>
rect 163 189 164 190 
<< m1 >>
rect 178 189 179 190 
<< m1 >>
rect 185 189 186 190 
<< m1 >>
rect 187 189 188 190 
<< m1 >>
rect 214 189 215 190 
<< m1 >>
rect 221 189 222 190 
<< m1 >>
rect 224 189 225 190 
<< m1 >>
rect 226 189 227 190 
<< m2 >>
rect 231 189 232 190 
<< m1 >>
rect 235 189 236 190 
<< m1 >>
rect 237 189 238 190 
<< m1 >>
rect 242 189 243 190 
<< m1 >>
rect 244 189 245 190 
<< m2 >>
rect 246 189 247 190 
<< m1 >>
rect 247 189 248 190 
<< m1 >>
rect 253 189 254 190 
<< m2 >>
rect 253 189 254 190 
<< m2c >>
rect 253 189 254 190 
<< m1 >>
rect 253 189 254 190 
<< m2 >>
rect 253 189 254 190 
<< m1 >>
rect 278 189 279 190 
<< m2 >>
rect 278 189 279 190 
<< m2c >>
rect 278 189 279 190 
<< m1 >>
rect 278 189 279 190 
<< m2 >>
rect 278 189 279 190 
<< m2 >>
rect 295 189 296 190 
<< m1 >>
rect 296 189 297 190 
<< m1 >>
rect 297 189 298 190 
<< m1 >>
rect 298 189 299 190 
<< m2 >>
rect 298 189 299 190 
<< m1 >>
rect 299 189 300 190 
<< m1 >>
rect 300 189 301 190 
<< m2 >>
rect 300 189 301 190 
<< m2c >>
rect 300 189 301 190 
<< m1 >>
rect 300 189 301 190 
<< m2 >>
rect 300 189 301 190 
<< m1 >>
rect 334 189 335 190 
<< m1 >>
rect 340 189 341 190 
<< m1 >>
rect 343 189 344 190 
<< m1 >>
rect 348 189 349 190 
<< m1 >>
rect 352 189 353 190 
<< m1 >>
rect 358 189 359 190 
<< m1 >>
rect 379 189 380 190 
<< m1 >>
rect 391 189 392 190 
<< m1 >>
rect 392 189 393 190 
<< m1 >>
rect 393 189 394 190 
<< m1 >>
rect 394 189 395 190 
<< m2 >>
rect 394 189 395 190 
<< m1 >>
rect 395 189 396 190 
<< m1 >>
rect 396 189 397 190 
<< m1 >>
rect 397 189 398 190 
<< m2 >>
rect 397 189 398 190 
<< m1 >>
rect 398 189 399 190 
<< m1 >>
rect 399 189 400 190 
<< m1 >>
rect 400 189 401 190 
<< m1 >>
rect 401 189 402 190 
<< m1 >>
rect 402 189 403 190 
<< m2 >>
rect 402 189 403 190 
<< m1 >>
rect 403 189 404 190 
<< m1 >>
rect 404 189 405 190 
<< m2 >>
rect 404 189 405 190 
<< m2c >>
rect 404 189 405 190 
<< m1 >>
rect 404 189 405 190 
<< m2 >>
rect 404 189 405 190 
<< m2 >>
rect 405 189 406 190 
<< m1 >>
rect 406 189 407 190 
<< m1 >>
rect 415 189 416 190 
<< m1 >>
rect 417 189 418 190 
<< m1 >>
rect 419 189 420 190 
<< m1 >>
rect 423 189 424 190 
<< m1 >>
rect 427 189 428 190 
<< m1 >>
rect 433 189 434 190 
<< m2 >>
rect 433 189 434 190 
<< m1 >>
rect 456 189 457 190 
<< m1 >>
rect 478 189 479 190 
<< m1 >>
rect 28 190 29 191 
<< m1 >>
rect 64 190 65 191 
<< m1 >>
rect 98 190 99 191 
<< m1 >>
rect 103 190 104 191 
<< m1 >>
rect 106 190 107 191 
<< m1 >>
rect 127 190 128 191 
<< m1 >>
rect 147 190 148 191 
<< m1 >>
rect 154 190 155 191 
<< m1 >>
rect 163 190 164 191 
<< m1 >>
rect 178 190 179 191 
<< m1 >>
rect 185 190 186 191 
<< m1 >>
rect 187 190 188 191 
<< m1 >>
rect 208 190 209 191 
<< m1 >>
rect 209 190 210 191 
<< m1 >>
rect 210 190 211 191 
<< m1 >>
rect 211 190 212 191 
<< m1 >>
rect 214 190 215 191 
<< m1 >>
rect 219 190 220 191 
<< m2 >>
rect 219 190 220 191 
<< m2c >>
rect 219 190 220 191 
<< m1 >>
rect 219 190 220 191 
<< m2 >>
rect 219 190 220 191 
<< m2 >>
rect 220 190 221 191 
<< m1 >>
rect 221 190 222 191 
<< m2 >>
rect 221 190 222 191 
<< m2 >>
rect 222 190 223 191 
<< m2 >>
rect 223 190 224 191 
<< m1 >>
rect 224 190 225 191 
<< m2 >>
rect 224 190 225 191 
<< m2 >>
rect 225 190 226 191 
<< m1 >>
rect 226 190 227 191 
<< m2 >>
rect 226 190 227 191 
<< m2 >>
rect 227 190 228 191 
<< m1 >>
rect 228 190 229 191 
<< m2 >>
rect 228 190 229 191 
<< m2c >>
rect 228 190 229 191 
<< m1 >>
rect 228 190 229 191 
<< m2 >>
rect 228 190 229 191 
<< m1 >>
rect 229 190 230 191 
<< m1 >>
rect 230 190 231 191 
<< m1 >>
rect 231 190 232 191 
<< m2 >>
rect 231 190 232 191 
<< m2c >>
rect 231 190 232 191 
<< m1 >>
rect 231 190 232 191 
<< m2 >>
rect 231 190 232 191 
<< m1 >>
rect 235 190 236 191 
<< m1 >>
rect 237 190 238 191 
<< m2 >>
rect 241 190 242 191 
<< m1 >>
rect 242 190 243 191 
<< m2 >>
rect 242 190 243 191 
<< m2 >>
rect 243 190 244 191 
<< m1 >>
rect 244 190 245 191 
<< m2 >>
rect 244 190 245 191 
<< m2 >>
rect 245 190 246 191 
<< m2 >>
rect 246 190 247 191 
<< m1 >>
rect 247 190 248 191 
<< m1 >>
rect 253 190 254 191 
<< m1 >>
rect 262 190 263 191 
<< m1 >>
rect 263 190 264 191 
<< m1 >>
rect 264 190 265 191 
<< m1 >>
rect 265 190 266 191 
<< m1 >>
rect 278 190 279 191 
<< m2 >>
rect 295 190 296 191 
<< m1 >>
rect 296 190 297 191 
<< m2 >>
rect 298 190 299 191 
<< m1 >>
rect 304 190 305 191 
<< m1 >>
rect 305 190 306 191 
<< m1 >>
rect 306 190 307 191 
<< m1 >>
rect 307 190 308 191 
<< m1 >>
rect 308 190 309 191 
<< m1 >>
rect 334 190 335 191 
<< m1 >>
rect 340 190 341 191 
<< m1 >>
rect 343 190 344 191 
<< m1 >>
rect 348 190 349 191 
<< m1 >>
rect 349 190 350 191 
<< m1 >>
rect 350 190 351 191 
<< m2 >>
rect 350 190 351 191 
<< m2c >>
rect 350 190 351 191 
<< m1 >>
rect 350 190 351 191 
<< m2 >>
rect 350 190 351 191 
<< m2 >>
rect 351 190 352 191 
<< m1 >>
rect 352 190 353 191 
<< m2 >>
rect 352 190 353 191 
<< m2 >>
rect 353 190 354 191 
<< m1 >>
rect 354 190 355 191 
<< m2 >>
rect 354 190 355 191 
<< m2c >>
rect 354 190 355 191 
<< m1 >>
rect 354 190 355 191 
<< m2 >>
rect 354 190 355 191 
<< m1 >>
rect 355 190 356 191 
<< m1 >>
rect 358 190 359 191 
<< m1 >>
rect 379 190 380 191 
<< m1 >>
rect 391 190 392 191 
<< m2 >>
rect 394 190 395 191 
<< m2 >>
rect 397 190 398 191 
<< m2 >>
rect 402 190 403 191 
<< m2 >>
rect 405 190 406 191 
<< m1 >>
rect 406 190 407 191 
<< m1 >>
rect 415 190 416 191 
<< m1 >>
rect 417 190 418 191 
<< m1 >>
rect 419 190 420 191 
<< m1 >>
rect 423 190 424 191 
<< m1 >>
rect 427 190 428 191 
<< m1 >>
rect 433 190 434 191 
<< m2 >>
rect 433 190 434 191 
<< m1 >>
rect 456 190 457 191 
<< m1 >>
rect 478 190 479 191 
<< m1 >>
rect 28 191 29 192 
<< m1 >>
rect 64 191 65 192 
<< m1 >>
rect 98 191 99 192 
<< m1 >>
rect 103 191 104 192 
<< m1 >>
rect 106 191 107 192 
<< m1 >>
rect 127 191 128 192 
<< m1 >>
rect 147 191 148 192 
<< m1 >>
rect 154 191 155 192 
<< m1 >>
rect 163 191 164 192 
<< m1 >>
rect 178 191 179 192 
<< m1 >>
rect 185 191 186 192 
<< m1 >>
rect 187 191 188 192 
<< m1 >>
rect 208 191 209 192 
<< m1 >>
rect 211 191 212 192 
<< m1 >>
rect 214 191 215 192 
<< m1 >>
rect 219 191 220 192 
<< m1 >>
rect 221 191 222 192 
<< m1 >>
rect 224 191 225 192 
<< m1 >>
rect 226 191 227 192 
<< m1 >>
rect 235 191 236 192 
<< m1 >>
rect 237 191 238 192 
<< m2 >>
rect 241 191 242 192 
<< m1 >>
rect 242 191 243 192 
<< m1 >>
rect 244 191 245 192 
<< m1 >>
rect 247 191 248 192 
<< m1 >>
rect 253 191 254 192 
<< m1 >>
rect 262 191 263 192 
<< m1 >>
rect 265 191 266 192 
<< m1 >>
rect 278 191 279 192 
<< m2 >>
rect 295 191 296 192 
<< m1 >>
rect 296 191 297 192 
<< m1 >>
rect 298 191 299 192 
<< m2 >>
rect 298 191 299 192 
<< m2c >>
rect 298 191 299 192 
<< m1 >>
rect 298 191 299 192 
<< m2 >>
rect 298 191 299 192 
<< m1 >>
rect 304 191 305 192 
<< m1 >>
rect 308 191 309 192 
<< m1 >>
rect 334 191 335 192 
<< m1 >>
rect 340 191 341 192 
<< m1 >>
rect 343 191 344 192 
<< m1 >>
rect 352 191 353 192 
<< m1 >>
rect 355 191 356 192 
<< m1 >>
rect 358 191 359 192 
<< m1 >>
rect 379 191 380 192 
<< m1 >>
rect 391 191 392 192 
<< m1 >>
rect 394 191 395 192 
<< m2 >>
rect 394 191 395 192 
<< m1 >>
rect 397 191 398 192 
<< m2 >>
rect 397 191 398 192 
<< m2c >>
rect 397 191 398 192 
<< m1 >>
rect 397 191 398 192 
<< m2 >>
rect 397 191 398 192 
<< m1 >>
rect 402 191 403 192 
<< m2 >>
rect 402 191 403 192 
<< m2c >>
rect 402 191 403 192 
<< m1 >>
rect 402 191 403 192 
<< m2 >>
rect 402 191 403 192 
<< m2 >>
rect 405 191 406 192 
<< m1 >>
rect 406 191 407 192 
<< m1 >>
rect 415 191 416 192 
<< m1 >>
rect 417 191 418 192 
<< m1 >>
rect 419 191 420 192 
<< m1 >>
rect 423 191 424 192 
<< m1 >>
rect 427 191 428 192 
<< m1 >>
rect 433 191 434 192 
<< m2 >>
rect 433 191 434 192 
<< m1 >>
rect 456 191 457 192 
<< m1 >>
rect 478 191 479 192 
<< m1 >>
rect 28 192 29 193 
<< pdiffusion >>
rect 30 192 31 193 
<< pdiffusion >>
rect 31 192 32 193 
<< pdiffusion >>
rect 32 192 33 193 
<< pdiffusion >>
rect 33 192 34 193 
<< pdiffusion >>
rect 34 192 35 193 
<< pdiffusion >>
rect 35 192 36 193 
<< pdiffusion >>
rect 48 192 49 193 
<< pdiffusion >>
rect 49 192 50 193 
<< pdiffusion >>
rect 50 192 51 193 
<< pdiffusion >>
rect 51 192 52 193 
<< pdiffusion >>
rect 52 192 53 193 
<< pdiffusion >>
rect 53 192 54 193 
<< m1 >>
rect 64 192 65 193 
<< pdiffusion >>
rect 66 192 67 193 
<< pdiffusion >>
rect 67 192 68 193 
<< pdiffusion >>
rect 68 192 69 193 
<< pdiffusion >>
rect 69 192 70 193 
<< pdiffusion >>
rect 70 192 71 193 
<< pdiffusion >>
rect 71 192 72 193 
<< pdiffusion >>
rect 84 192 85 193 
<< pdiffusion >>
rect 85 192 86 193 
<< pdiffusion >>
rect 86 192 87 193 
<< pdiffusion >>
rect 87 192 88 193 
<< pdiffusion >>
rect 88 192 89 193 
<< pdiffusion >>
rect 89 192 90 193 
<< m1 >>
rect 98 192 99 193 
<< pdiffusion >>
rect 102 192 103 193 
<< m1 >>
rect 103 192 104 193 
<< pdiffusion >>
rect 103 192 104 193 
<< pdiffusion >>
rect 104 192 105 193 
<< pdiffusion >>
rect 105 192 106 193 
<< m1 >>
rect 106 192 107 193 
<< pdiffusion >>
rect 106 192 107 193 
<< pdiffusion >>
rect 107 192 108 193 
<< pdiffusion >>
rect 120 192 121 193 
<< pdiffusion >>
rect 121 192 122 193 
<< pdiffusion >>
rect 122 192 123 193 
<< pdiffusion >>
rect 123 192 124 193 
<< pdiffusion >>
rect 124 192 125 193 
<< pdiffusion >>
rect 125 192 126 193 
<< m1 >>
rect 127 192 128 193 
<< pdiffusion >>
rect 138 192 139 193 
<< pdiffusion >>
rect 139 192 140 193 
<< pdiffusion >>
rect 140 192 141 193 
<< pdiffusion >>
rect 141 192 142 193 
<< pdiffusion >>
rect 142 192 143 193 
<< pdiffusion >>
rect 143 192 144 193 
<< m1 >>
rect 147 192 148 193 
<< m1 >>
rect 154 192 155 193 
<< pdiffusion >>
rect 156 192 157 193 
<< pdiffusion >>
rect 157 192 158 193 
<< pdiffusion >>
rect 158 192 159 193 
<< pdiffusion >>
rect 159 192 160 193 
<< pdiffusion >>
rect 160 192 161 193 
<< pdiffusion >>
rect 161 192 162 193 
<< m1 >>
rect 163 192 164 193 
<< pdiffusion >>
rect 174 192 175 193 
<< pdiffusion >>
rect 175 192 176 193 
<< pdiffusion >>
rect 176 192 177 193 
<< pdiffusion >>
rect 177 192 178 193 
<< m1 >>
rect 178 192 179 193 
<< pdiffusion >>
rect 178 192 179 193 
<< pdiffusion >>
rect 179 192 180 193 
<< m1 >>
rect 185 192 186 193 
<< m1 >>
rect 187 192 188 193 
<< pdiffusion >>
rect 192 192 193 193 
<< pdiffusion >>
rect 193 192 194 193 
<< pdiffusion >>
rect 194 192 195 193 
<< pdiffusion >>
rect 195 192 196 193 
<< pdiffusion >>
rect 196 192 197 193 
<< pdiffusion >>
rect 197 192 198 193 
<< m1 >>
rect 208 192 209 193 
<< pdiffusion >>
rect 210 192 211 193 
<< m1 >>
rect 211 192 212 193 
<< pdiffusion >>
rect 211 192 212 193 
<< pdiffusion >>
rect 212 192 213 193 
<< pdiffusion >>
rect 213 192 214 193 
<< m1 >>
rect 214 192 215 193 
<< pdiffusion >>
rect 214 192 215 193 
<< pdiffusion >>
rect 215 192 216 193 
<< m1 >>
rect 219 192 220 193 
<< m1 >>
rect 221 192 222 193 
<< m1 >>
rect 224 192 225 193 
<< m1 >>
rect 226 192 227 193 
<< m1 >>
rect 235 192 236 193 
<< m1 >>
rect 237 192 238 193 
<< m2 >>
rect 241 192 242 193 
<< m1 >>
rect 242 192 243 193 
<< m1 >>
rect 244 192 245 193 
<< pdiffusion >>
rect 246 192 247 193 
<< m1 >>
rect 247 192 248 193 
<< pdiffusion >>
rect 247 192 248 193 
<< pdiffusion >>
rect 248 192 249 193 
<< pdiffusion >>
rect 249 192 250 193 
<< pdiffusion >>
rect 250 192 251 193 
<< pdiffusion >>
rect 251 192 252 193 
<< m1 >>
rect 253 192 254 193 
<< m1 >>
rect 262 192 263 193 
<< pdiffusion >>
rect 264 192 265 193 
<< m1 >>
rect 265 192 266 193 
<< pdiffusion >>
rect 265 192 266 193 
<< pdiffusion >>
rect 266 192 267 193 
<< pdiffusion >>
rect 267 192 268 193 
<< pdiffusion >>
rect 268 192 269 193 
<< pdiffusion >>
rect 269 192 270 193 
<< m1 >>
rect 278 192 279 193 
<< pdiffusion >>
rect 282 192 283 193 
<< pdiffusion >>
rect 283 192 284 193 
<< pdiffusion >>
rect 284 192 285 193 
<< pdiffusion >>
rect 285 192 286 193 
<< pdiffusion >>
rect 286 192 287 193 
<< pdiffusion >>
rect 287 192 288 193 
<< m2 >>
rect 295 192 296 193 
<< m1 >>
rect 296 192 297 193 
<< m1 >>
rect 298 192 299 193 
<< pdiffusion >>
rect 300 192 301 193 
<< pdiffusion >>
rect 301 192 302 193 
<< pdiffusion >>
rect 302 192 303 193 
<< pdiffusion >>
rect 303 192 304 193 
<< m1 >>
rect 304 192 305 193 
<< pdiffusion >>
rect 304 192 305 193 
<< pdiffusion >>
rect 305 192 306 193 
<< m1 >>
rect 308 192 309 193 
<< pdiffusion >>
rect 318 192 319 193 
<< pdiffusion >>
rect 319 192 320 193 
<< pdiffusion >>
rect 320 192 321 193 
<< pdiffusion >>
rect 321 192 322 193 
<< pdiffusion >>
rect 322 192 323 193 
<< pdiffusion >>
rect 323 192 324 193 
<< m1 >>
rect 334 192 335 193 
<< pdiffusion >>
rect 336 192 337 193 
<< pdiffusion >>
rect 337 192 338 193 
<< pdiffusion >>
rect 338 192 339 193 
<< pdiffusion >>
rect 339 192 340 193 
<< m1 >>
rect 340 192 341 193 
<< pdiffusion >>
rect 340 192 341 193 
<< pdiffusion >>
rect 341 192 342 193 
<< m1 >>
rect 343 192 344 193 
<< m1 >>
rect 352 192 353 193 
<< pdiffusion >>
rect 354 192 355 193 
<< m1 >>
rect 355 192 356 193 
<< pdiffusion >>
rect 355 192 356 193 
<< pdiffusion >>
rect 356 192 357 193 
<< pdiffusion >>
rect 357 192 358 193 
<< m1 >>
rect 358 192 359 193 
<< pdiffusion >>
rect 358 192 359 193 
<< pdiffusion >>
rect 359 192 360 193 
<< pdiffusion >>
rect 372 192 373 193 
<< pdiffusion >>
rect 373 192 374 193 
<< pdiffusion >>
rect 374 192 375 193 
<< pdiffusion >>
rect 375 192 376 193 
<< pdiffusion >>
rect 376 192 377 193 
<< pdiffusion >>
rect 377 192 378 193 
<< m1 >>
rect 379 192 380 193 
<< pdiffusion >>
rect 390 192 391 193 
<< m1 >>
rect 391 192 392 193 
<< pdiffusion >>
rect 391 192 392 193 
<< pdiffusion >>
rect 392 192 393 193 
<< m1 >>
rect 393 192 394 193 
<< m2 >>
rect 393 192 394 193 
<< m2c >>
rect 393 192 394 193 
<< m1 >>
rect 393 192 394 193 
<< m2 >>
rect 393 192 394 193 
<< pdiffusion >>
rect 393 192 394 193 
<< m1 >>
rect 394 192 395 193 
<< pdiffusion >>
rect 394 192 395 193 
<< pdiffusion >>
rect 395 192 396 193 
<< m1 >>
rect 397 192 398 193 
<< m1 >>
rect 402 192 403 193 
<< m2 >>
rect 405 192 406 193 
<< m1 >>
rect 406 192 407 193 
<< pdiffusion >>
rect 408 192 409 193 
<< pdiffusion >>
rect 409 192 410 193 
<< pdiffusion >>
rect 410 192 411 193 
<< pdiffusion >>
rect 411 192 412 193 
<< pdiffusion >>
rect 412 192 413 193 
<< pdiffusion >>
rect 413 192 414 193 
<< m1 >>
rect 415 192 416 193 
<< m1 >>
rect 417 192 418 193 
<< m1 >>
rect 419 192 420 193 
<< m1 >>
rect 423 192 424 193 
<< pdiffusion >>
rect 426 192 427 193 
<< m1 >>
rect 427 192 428 193 
<< pdiffusion >>
rect 427 192 428 193 
<< pdiffusion >>
rect 428 192 429 193 
<< pdiffusion >>
rect 429 192 430 193 
<< pdiffusion >>
rect 430 192 431 193 
<< pdiffusion >>
rect 431 192 432 193 
<< m1 >>
rect 433 192 434 193 
<< m2 >>
rect 433 192 434 193 
<< pdiffusion >>
rect 444 192 445 193 
<< pdiffusion >>
rect 445 192 446 193 
<< pdiffusion >>
rect 446 192 447 193 
<< pdiffusion >>
rect 447 192 448 193 
<< pdiffusion >>
rect 448 192 449 193 
<< pdiffusion >>
rect 449 192 450 193 
<< m1 >>
rect 456 192 457 193 
<< pdiffusion >>
rect 462 192 463 193 
<< pdiffusion >>
rect 463 192 464 193 
<< pdiffusion >>
rect 464 192 465 193 
<< pdiffusion >>
rect 465 192 466 193 
<< pdiffusion >>
rect 466 192 467 193 
<< pdiffusion >>
rect 467 192 468 193 
<< m1 >>
rect 478 192 479 193 
<< pdiffusion >>
rect 480 192 481 193 
<< pdiffusion >>
rect 481 192 482 193 
<< pdiffusion >>
rect 482 192 483 193 
<< pdiffusion >>
rect 483 192 484 193 
<< pdiffusion >>
rect 484 192 485 193 
<< pdiffusion >>
rect 485 192 486 193 
<< pdiffusion >>
rect 498 192 499 193 
<< pdiffusion >>
rect 499 192 500 193 
<< pdiffusion >>
rect 500 192 501 193 
<< pdiffusion >>
rect 501 192 502 193 
<< pdiffusion >>
rect 502 192 503 193 
<< pdiffusion >>
rect 503 192 504 193 
<< pdiffusion >>
rect 516 192 517 193 
<< pdiffusion >>
rect 517 192 518 193 
<< pdiffusion >>
rect 518 192 519 193 
<< pdiffusion >>
rect 519 192 520 193 
<< pdiffusion >>
rect 520 192 521 193 
<< pdiffusion >>
rect 521 192 522 193 
<< m1 >>
rect 28 193 29 194 
<< pdiffusion >>
rect 30 193 31 194 
<< pdiffusion >>
rect 31 193 32 194 
<< pdiffusion >>
rect 32 193 33 194 
<< pdiffusion >>
rect 33 193 34 194 
<< pdiffusion >>
rect 34 193 35 194 
<< pdiffusion >>
rect 35 193 36 194 
<< pdiffusion >>
rect 48 193 49 194 
<< pdiffusion >>
rect 49 193 50 194 
<< pdiffusion >>
rect 50 193 51 194 
<< pdiffusion >>
rect 51 193 52 194 
<< pdiffusion >>
rect 52 193 53 194 
<< pdiffusion >>
rect 53 193 54 194 
<< m1 >>
rect 64 193 65 194 
<< pdiffusion >>
rect 66 193 67 194 
<< pdiffusion >>
rect 67 193 68 194 
<< pdiffusion >>
rect 68 193 69 194 
<< pdiffusion >>
rect 69 193 70 194 
<< pdiffusion >>
rect 70 193 71 194 
<< pdiffusion >>
rect 71 193 72 194 
<< pdiffusion >>
rect 84 193 85 194 
<< pdiffusion >>
rect 85 193 86 194 
<< pdiffusion >>
rect 86 193 87 194 
<< pdiffusion >>
rect 87 193 88 194 
<< pdiffusion >>
rect 88 193 89 194 
<< pdiffusion >>
rect 89 193 90 194 
<< m1 >>
rect 98 193 99 194 
<< pdiffusion >>
rect 102 193 103 194 
<< pdiffusion >>
rect 103 193 104 194 
<< pdiffusion >>
rect 104 193 105 194 
<< pdiffusion >>
rect 105 193 106 194 
<< pdiffusion >>
rect 106 193 107 194 
<< pdiffusion >>
rect 107 193 108 194 
<< pdiffusion >>
rect 120 193 121 194 
<< pdiffusion >>
rect 121 193 122 194 
<< pdiffusion >>
rect 122 193 123 194 
<< pdiffusion >>
rect 123 193 124 194 
<< pdiffusion >>
rect 124 193 125 194 
<< pdiffusion >>
rect 125 193 126 194 
<< m1 >>
rect 127 193 128 194 
<< pdiffusion >>
rect 138 193 139 194 
<< pdiffusion >>
rect 139 193 140 194 
<< pdiffusion >>
rect 140 193 141 194 
<< pdiffusion >>
rect 141 193 142 194 
<< pdiffusion >>
rect 142 193 143 194 
<< pdiffusion >>
rect 143 193 144 194 
<< m1 >>
rect 147 193 148 194 
<< m1 >>
rect 154 193 155 194 
<< pdiffusion >>
rect 156 193 157 194 
<< pdiffusion >>
rect 157 193 158 194 
<< pdiffusion >>
rect 158 193 159 194 
<< pdiffusion >>
rect 159 193 160 194 
<< pdiffusion >>
rect 160 193 161 194 
<< pdiffusion >>
rect 161 193 162 194 
<< m1 >>
rect 163 193 164 194 
<< pdiffusion >>
rect 174 193 175 194 
<< pdiffusion >>
rect 175 193 176 194 
<< pdiffusion >>
rect 176 193 177 194 
<< pdiffusion >>
rect 177 193 178 194 
<< pdiffusion >>
rect 178 193 179 194 
<< pdiffusion >>
rect 179 193 180 194 
<< m1 >>
rect 185 193 186 194 
<< m1 >>
rect 187 193 188 194 
<< pdiffusion >>
rect 192 193 193 194 
<< pdiffusion >>
rect 193 193 194 194 
<< pdiffusion >>
rect 194 193 195 194 
<< pdiffusion >>
rect 195 193 196 194 
<< pdiffusion >>
rect 196 193 197 194 
<< pdiffusion >>
rect 197 193 198 194 
<< m1 >>
rect 208 193 209 194 
<< pdiffusion >>
rect 210 193 211 194 
<< pdiffusion >>
rect 211 193 212 194 
<< pdiffusion >>
rect 212 193 213 194 
<< pdiffusion >>
rect 213 193 214 194 
<< pdiffusion >>
rect 214 193 215 194 
<< pdiffusion >>
rect 215 193 216 194 
<< m1 >>
rect 219 193 220 194 
<< m1 >>
rect 221 193 222 194 
<< m1 >>
rect 224 193 225 194 
<< m1 >>
rect 226 193 227 194 
<< m1 >>
rect 235 193 236 194 
<< m1 >>
rect 237 193 238 194 
<< m2 >>
rect 241 193 242 194 
<< m1 >>
rect 242 193 243 194 
<< m1 >>
rect 244 193 245 194 
<< pdiffusion >>
rect 246 193 247 194 
<< pdiffusion >>
rect 247 193 248 194 
<< pdiffusion >>
rect 248 193 249 194 
<< pdiffusion >>
rect 249 193 250 194 
<< pdiffusion >>
rect 250 193 251 194 
<< pdiffusion >>
rect 251 193 252 194 
<< m1 >>
rect 253 193 254 194 
<< m1 >>
rect 262 193 263 194 
<< pdiffusion >>
rect 264 193 265 194 
<< pdiffusion >>
rect 265 193 266 194 
<< pdiffusion >>
rect 266 193 267 194 
<< pdiffusion >>
rect 267 193 268 194 
<< pdiffusion >>
rect 268 193 269 194 
<< pdiffusion >>
rect 269 193 270 194 
<< m1 >>
rect 278 193 279 194 
<< pdiffusion >>
rect 282 193 283 194 
<< pdiffusion >>
rect 283 193 284 194 
<< pdiffusion >>
rect 284 193 285 194 
<< pdiffusion >>
rect 285 193 286 194 
<< pdiffusion >>
rect 286 193 287 194 
<< pdiffusion >>
rect 287 193 288 194 
<< m2 >>
rect 295 193 296 194 
<< m1 >>
rect 296 193 297 194 
<< m1 >>
rect 298 193 299 194 
<< pdiffusion >>
rect 300 193 301 194 
<< pdiffusion >>
rect 301 193 302 194 
<< pdiffusion >>
rect 302 193 303 194 
<< pdiffusion >>
rect 303 193 304 194 
<< pdiffusion >>
rect 304 193 305 194 
<< pdiffusion >>
rect 305 193 306 194 
<< m1 >>
rect 308 193 309 194 
<< pdiffusion >>
rect 318 193 319 194 
<< pdiffusion >>
rect 319 193 320 194 
<< pdiffusion >>
rect 320 193 321 194 
<< pdiffusion >>
rect 321 193 322 194 
<< pdiffusion >>
rect 322 193 323 194 
<< pdiffusion >>
rect 323 193 324 194 
<< m1 >>
rect 334 193 335 194 
<< pdiffusion >>
rect 336 193 337 194 
<< pdiffusion >>
rect 337 193 338 194 
<< pdiffusion >>
rect 338 193 339 194 
<< pdiffusion >>
rect 339 193 340 194 
<< pdiffusion >>
rect 340 193 341 194 
<< pdiffusion >>
rect 341 193 342 194 
<< m1 >>
rect 343 193 344 194 
<< m1 >>
rect 352 193 353 194 
<< pdiffusion >>
rect 354 193 355 194 
<< pdiffusion >>
rect 355 193 356 194 
<< pdiffusion >>
rect 356 193 357 194 
<< pdiffusion >>
rect 357 193 358 194 
<< pdiffusion >>
rect 358 193 359 194 
<< pdiffusion >>
rect 359 193 360 194 
<< pdiffusion >>
rect 372 193 373 194 
<< pdiffusion >>
rect 373 193 374 194 
<< pdiffusion >>
rect 374 193 375 194 
<< pdiffusion >>
rect 375 193 376 194 
<< pdiffusion >>
rect 376 193 377 194 
<< pdiffusion >>
rect 377 193 378 194 
<< m1 >>
rect 379 193 380 194 
<< pdiffusion >>
rect 390 193 391 194 
<< pdiffusion >>
rect 391 193 392 194 
<< pdiffusion >>
rect 392 193 393 194 
<< pdiffusion >>
rect 393 193 394 194 
<< pdiffusion >>
rect 394 193 395 194 
<< pdiffusion >>
rect 395 193 396 194 
<< m1 >>
rect 397 193 398 194 
<< m1 >>
rect 398 193 399 194 
<< m1 >>
rect 399 193 400 194 
<< m1 >>
rect 400 193 401 194 
<< m2 >>
rect 400 193 401 194 
<< m2c >>
rect 400 193 401 194 
<< m1 >>
rect 400 193 401 194 
<< m2 >>
rect 400 193 401 194 
<< m2 >>
rect 401 193 402 194 
<< m1 >>
rect 402 193 403 194 
<< m2 >>
rect 402 193 403 194 
<< m2 >>
rect 403 193 404 194 
<< m1 >>
rect 404 193 405 194 
<< m2 >>
rect 404 193 405 194 
<< m2c >>
rect 404 193 405 194 
<< m1 >>
rect 404 193 405 194 
<< m2 >>
rect 404 193 405 194 
<< m2 >>
rect 405 193 406 194 
<< m1 >>
rect 406 193 407 194 
<< pdiffusion >>
rect 408 193 409 194 
<< pdiffusion >>
rect 409 193 410 194 
<< pdiffusion >>
rect 410 193 411 194 
<< pdiffusion >>
rect 411 193 412 194 
<< pdiffusion >>
rect 412 193 413 194 
<< pdiffusion >>
rect 413 193 414 194 
<< m1 >>
rect 415 193 416 194 
<< m1 >>
rect 417 193 418 194 
<< m1 >>
rect 419 193 420 194 
<< m1 >>
rect 423 193 424 194 
<< pdiffusion >>
rect 426 193 427 194 
<< pdiffusion >>
rect 427 193 428 194 
<< pdiffusion >>
rect 428 193 429 194 
<< pdiffusion >>
rect 429 193 430 194 
<< pdiffusion >>
rect 430 193 431 194 
<< pdiffusion >>
rect 431 193 432 194 
<< m1 >>
rect 433 193 434 194 
<< m2 >>
rect 433 193 434 194 
<< pdiffusion >>
rect 444 193 445 194 
<< pdiffusion >>
rect 445 193 446 194 
<< pdiffusion >>
rect 446 193 447 194 
<< pdiffusion >>
rect 447 193 448 194 
<< pdiffusion >>
rect 448 193 449 194 
<< pdiffusion >>
rect 449 193 450 194 
<< m1 >>
rect 456 193 457 194 
<< pdiffusion >>
rect 462 193 463 194 
<< pdiffusion >>
rect 463 193 464 194 
<< pdiffusion >>
rect 464 193 465 194 
<< pdiffusion >>
rect 465 193 466 194 
<< pdiffusion >>
rect 466 193 467 194 
<< pdiffusion >>
rect 467 193 468 194 
<< m1 >>
rect 478 193 479 194 
<< pdiffusion >>
rect 480 193 481 194 
<< pdiffusion >>
rect 481 193 482 194 
<< pdiffusion >>
rect 482 193 483 194 
<< pdiffusion >>
rect 483 193 484 194 
<< pdiffusion >>
rect 484 193 485 194 
<< pdiffusion >>
rect 485 193 486 194 
<< pdiffusion >>
rect 498 193 499 194 
<< pdiffusion >>
rect 499 193 500 194 
<< pdiffusion >>
rect 500 193 501 194 
<< pdiffusion >>
rect 501 193 502 194 
<< pdiffusion >>
rect 502 193 503 194 
<< pdiffusion >>
rect 503 193 504 194 
<< pdiffusion >>
rect 516 193 517 194 
<< pdiffusion >>
rect 517 193 518 194 
<< pdiffusion >>
rect 518 193 519 194 
<< pdiffusion >>
rect 519 193 520 194 
<< pdiffusion >>
rect 520 193 521 194 
<< pdiffusion >>
rect 521 193 522 194 
<< m1 >>
rect 28 194 29 195 
<< pdiffusion >>
rect 30 194 31 195 
<< pdiffusion >>
rect 31 194 32 195 
<< pdiffusion >>
rect 32 194 33 195 
<< pdiffusion >>
rect 33 194 34 195 
<< pdiffusion >>
rect 34 194 35 195 
<< pdiffusion >>
rect 35 194 36 195 
<< pdiffusion >>
rect 48 194 49 195 
<< pdiffusion >>
rect 49 194 50 195 
<< pdiffusion >>
rect 50 194 51 195 
<< pdiffusion >>
rect 51 194 52 195 
<< pdiffusion >>
rect 52 194 53 195 
<< pdiffusion >>
rect 53 194 54 195 
<< m1 >>
rect 64 194 65 195 
<< pdiffusion >>
rect 66 194 67 195 
<< pdiffusion >>
rect 67 194 68 195 
<< pdiffusion >>
rect 68 194 69 195 
<< pdiffusion >>
rect 69 194 70 195 
<< pdiffusion >>
rect 70 194 71 195 
<< pdiffusion >>
rect 71 194 72 195 
<< pdiffusion >>
rect 84 194 85 195 
<< pdiffusion >>
rect 85 194 86 195 
<< pdiffusion >>
rect 86 194 87 195 
<< pdiffusion >>
rect 87 194 88 195 
<< pdiffusion >>
rect 88 194 89 195 
<< pdiffusion >>
rect 89 194 90 195 
<< m1 >>
rect 98 194 99 195 
<< pdiffusion >>
rect 102 194 103 195 
<< pdiffusion >>
rect 103 194 104 195 
<< pdiffusion >>
rect 104 194 105 195 
<< pdiffusion >>
rect 105 194 106 195 
<< pdiffusion >>
rect 106 194 107 195 
<< pdiffusion >>
rect 107 194 108 195 
<< pdiffusion >>
rect 120 194 121 195 
<< pdiffusion >>
rect 121 194 122 195 
<< pdiffusion >>
rect 122 194 123 195 
<< pdiffusion >>
rect 123 194 124 195 
<< pdiffusion >>
rect 124 194 125 195 
<< pdiffusion >>
rect 125 194 126 195 
<< m1 >>
rect 127 194 128 195 
<< pdiffusion >>
rect 138 194 139 195 
<< pdiffusion >>
rect 139 194 140 195 
<< pdiffusion >>
rect 140 194 141 195 
<< pdiffusion >>
rect 141 194 142 195 
<< pdiffusion >>
rect 142 194 143 195 
<< pdiffusion >>
rect 143 194 144 195 
<< m1 >>
rect 147 194 148 195 
<< m1 >>
rect 154 194 155 195 
<< pdiffusion >>
rect 156 194 157 195 
<< pdiffusion >>
rect 157 194 158 195 
<< pdiffusion >>
rect 158 194 159 195 
<< pdiffusion >>
rect 159 194 160 195 
<< pdiffusion >>
rect 160 194 161 195 
<< pdiffusion >>
rect 161 194 162 195 
<< m1 >>
rect 163 194 164 195 
<< pdiffusion >>
rect 174 194 175 195 
<< pdiffusion >>
rect 175 194 176 195 
<< pdiffusion >>
rect 176 194 177 195 
<< pdiffusion >>
rect 177 194 178 195 
<< pdiffusion >>
rect 178 194 179 195 
<< pdiffusion >>
rect 179 194 180 195 
<< m1 >>
rect 185 194 186 195 
<< m1 >>
rect 187 194 188 195 
<< pdiffusion >>
rect 192 194 193 195 
<< pdiffusion >>
rect 193 194 194 195 
<< pdiffusion >>
rect 194 194 195 195 
<< pdiffusion >>
rect 195 194 196 195 
<< pdiffusion >>
rect 196 194 197 195 
<< pdiffusion >>
rect 197 194 198 195 
<< m1 >>
rect 208 194 209 195 
<< pdiffusion >>
rect 210 194 211 195 
<< pdiffusion >>
rect 211 194 212 195 
<< pdiffusion >>
rect 212 194 213 195 
<< pdiffusion >>
rect 213 194 214 195 
<< pdiffusion >>
rect 214 194 215 195 
<< pdiffusion >>
rect 215 194 216 195 
<< m1 >>
rect 219 194 220 195 
<< m1 >>
rect 221 194 222 195 
<< m1 >>
rect 224 194 225 195 
<< m1 >>
rect 226 194 227 195 
<< m1 >>
rect 235 194 236 195 
<< m1 >>
rect 237 194 238 195 
<< m2 >>
rect 241 194 242 195 
<< m1 >>
rect 242 194 243 195 
<< m1 >>
rect 244 194 245 195 
<< pdiffusion >>
rect 246 194 247 195 
<< pdiffusion >>
rect 247 194 248 195 
<< pdiffusion >>
rect 248 194 249 195 
<< pdiffusion >>
rect 249 194 250 195 
<< pdiffusion >>
rect 250 194 251 195 
<< pdiffusion >>
rect 251 194 252 195 
<< m1 >>
rect 253 194 254 195 
<< m1 >>
rect 262 194 263 195 
<< pdiffusion >>
rect 264 194 265 195 
<< pdiffusion >>
rect 265 194 266 195 
<< pdiffusion >>
rect 266 194 267 195 
<< pdiffusion >>
rect 267 194 268 195 
<< pdiffusion >>
rect 268 194 269 195 
<< pdiffusion >>
rect 269 194 270 195 
<< m1 >>
rect 278 194 279 195 
<< pdiffusion >>
rect 282 194 283 195 
<< pdiffusion >>
rect 283 194 284 195 
<< pdiffusion >>
rect 284 194 285 195 
<< pdiffusion >>
rect 285 194 286 195 
<< pdiffusion >>
rect 286 194 287 195 
<< pdiffusion >>
rect 287 194 288 195 
<< m2 >>
rect 295 194 296 195 
<< m1 >>
rect 296 194 297 195 
<< m1 >>
rect 298 194 299 195 
<< pdiffusion >>
rect 300 194 301 195 
<< pdiffusion >>
rect 301 194 302 195 
<< pdiffusion >>
rect 302 194 303 195 
<< pdiffusion >>
rect 303 194 304 195 
<< pdiffusion >>
rect 304 194 305 195 
<< pdiffusion >>
rect 305 194 306 195 
<< m1 >>
rect 308 194 309 195 
<< pdiffusion >>
rect 318 194 319 195 
<< pdiffusion >>
rect 319 194 320 195 
<< pdiffusion >>
rect 320 194 321 195 
<< pdiffusion >>
rect 321 194 322 195 
<< pdiffusion >>
rect 322 194 323 195 
<< pdiffusion >>
rect 323 194 324 195 
<< m1 >>
rect 334 194 335 195 
<< pdiffusion >>
rect 336 194 337 195 
<< pdiffusion >>
rect 337 194 338 195 
<< pdiffusion >>
rect 338 194 339 195 
<< pdiffusion >>
rect 339 194 340 195 
<< pdiffusion >>
rect 340 194 341 195 
<< pdiffusion >>
rect 341 194 342 195 
<< m1 >>
rect 343 194 344 195 
<< m1 >>
rect 352 194 353 195 
<< pdiffusion >>
rect 354 194 355 195 
<< pdiffusion >>
rect 355 194 356 195 
<< pdiffusion >>
rect 356 194 357 195 
<< pdiffusion >>
rect 357 194 358 195 
<< pdiffusion >>
rect 358 194 359 195 
<< pdiffusion >>
rect 359 194 360 195 
<< pdiffusion >>
rect 372 194 373 195 
<< pdiffusion >>
rect 373 194 374 195 
<< pdiffusion >>
rect 374 194 375 195 
<< pdiffusion >>
rect 375 194 376 195 
<< pdiffusion >>
rect 376 194 377 195 
<< pdiffusion >>
rect 377 194 378 195 
<< m1 >>
rect 379 194 380 195 
<< pdiffusion >>
rect 390 194 391 195 
<< pdiffusion >>
rect 391 194 392 195 
<< pdiffusion >>
rect 392 194 393 195 
<< pdiffusion >>
rect 393 194 394 195 
<< pdiffusion >>
rect 394 194 395 195 
<< pdiffusion >>
rect 395 194 396 195 
<< m1 >>
rect 402 194 403 195 
<< m1 >>
rect 404 194 405 195 
<< m2 >>
rect 405 194 406 195 
<< m1 >>
rect 406 194 407 195 
<< pdiffusion >>
rect 408 194 409 195 
<< pdiffusion >>
rect 409 194 410 195 
<< pdiffusion >>
rect 410 194 411 195 
<< pdiffusion >>
rect 411 194 412 195 
<< pdiffusion >>
rect 412 194 413 195 
<< pdiffusion >>
rect 413 194 414 195 
<< m1 >>
rect 415 194 416 195 
<< m1 >>
rect 417 194 418 195 
<< m1 >>
rect 419 194 420 195 
<< m1 >>
rect 423 194 424 195 
<< pdiffusion >>
rect 426 194 427 195 
<< pdiffusion >>
rect 427 194 428 195 
<< pdiffusion >>
rect 428 194 429 195 
<< pdiffusion >>
rect 429 194 430 195 
<< pdiffusion >>
rect 430 194 431 195 
<< pdiffusion >>
rect 431 194 432 195 
<< m1 >>
rect 433 194 434 195 
<< m2 >>
rect 433 194 434 195 
<< pdiffusion >>
rect 444 194 445 195 
<< pdiffusion >>
rect 445 194 446 195 
<< pdiffusion >>
rect 446 194 447 195 
<< pdiffusion >>
rect 447 194 448 195 
<< pdiffusion >>
rect 448 194 449 195 
<< pdiffusion >>
rect 449 194 450 195 
<< m1 >>
rect 456 194 457 195 
<< pdiffusion >>
rect 462 194 463 195 
<< pdiffusion >>
rect 463 194 464 195 
<< pdiffusion >>
rect 464 194 465 195 
<< pdiffusion >>
rect 465 194 466 195 
<< pdiffusion >>
rect 466 194 467 195 
<< pdiffusion >>
rect 467 194 468 195 
<< m1 >>
rect 478 194 479 195 
<< pdiffusion >>
rect 480 194 481 195 
<< pdiffusion >>
rect 481 194 482 195 
<< pdiffusion >>
rect 482 194 483 195 
<< pdiffusion >>
rect 483 194 484 195 
<< pdiffusion >>
rect 484 194 485 195 
<< pdiffusion >>
rect 485 194 486 195 
<< pdiffusion >>
rect 498 194 499 195 
<< pdiffusion >>
rect 499 194 500 195 
<< pdiffusion >>
rect 500 194 501 195 
<< pdiffusion >>
rect 501 194 502 195 
<< pdiffusion >>
rect 502 194 503 195 
<< pdiffusion >>
rect 503 194 504 195 
<< pdiffusion >>
rect 516 194 517 195 
<< pdiffusion >>
rect 517 194 518 195 
<< pdiffusion >>
rect 518 194 519 195 
<< pdiffusion >>
rect 519 194 520 195 
<< pdiffusion >>
rect 520 194 521 195 
<< pdiffusion >>
rect 521 194 522 195 
<< m1 >>
rect 28 195 29 196 
<< pdiffusion >>
rect 30 195 31 196 
<< pdiffusion >>
rect 31 195 32 196 
<< pdiffusion >>
rect 32 195 33 196 
<< pdiffusion >>
rect 33 195 34 196 
<< pdiffusion >>
rect 34 195 35 196 
<< pdiffusion >>
rect 35 195 36 196 
<< pdiffusion >>
rect 48 195 49 196 
<< pdiffusion >>
rect 49 195 50 196 
<< pdiffusion >>
rect 50 195 51 196 
<< pdiffusion >>
rect 51 195 52 196 
<< pdiffusion >>
rect 52 195 53 196 
<< pdiffusion >>
rect 53 195 54 196 
<< m1 >>
rect 64 195 65 196 
<< pdiffusion >>
rect 66 195 67 196 
<< pdiffusion >>
rect 67 195 68 196 
<< pdiffusion >>
rect 68 195 69 196 
<< pdiffusion >>
rect 69 195 70 196 
<< pdiffusion >>
rect 70 195 71 196 
<< pdiffusion >>
rect 71 195 72 196 
<< pdiffusion >>
rect 84 195 85 196 
<< pdiffusion >>
rect 85 195 86 196 
<< pdiffusion >>
rect 86 195 87 196 
<< pdiffusion >>
rect 87 195 88 196 
<< pdiffusion >>
rect 88 195 89 196 
<< pdiffusion >>
rect 89 195 90 196 
<< m1 >>
rect 98 195 99 196 
<< pdiffusion >>
rect 102 195 103 196 
<< pdiffusion >>
rect 103 195 104 196 
<< pdiffusion >>
rect 104 195 105 196 
<< pdiffusion >>
rect 105 195 106 196 
<< pdiffusion >>
rect 106 195 107 196 
<< pdiffusion >>
rect 107 195 108 196 
<< pdiffusion >>
rect 120 195 121 196 
<< pdiffusion >>
rect 121 195 122 196 
<< pdiffusion >>
rect 122 195 123 196 
<< pdiffusion >>
rect 123 195 124 196 
<< pdiffusion >>
rect 124 195 125 196 
<< pdiffusion >>
rect 125 195 126 196 
<< m1 >>
rect 127 195 128 196 
<< pdiffusion >>
rect 138 195 139 196 
<< pdiffusion >>
rect 139 195 140 196 
<< pdiffusion >>
rect 140 195 141 196 
<< pdiffusion >>
rect 141 195 142 196 
<< pdiffusion >>
rect 142 195 143 196 
<< pdiffusion >>
rect 143 195 144 196 
<< m1 >>
rect 147 195 148 196 
<< m1 >>
rect 154 195 155 196 
<< pdiffusion >>
rect 156 195 157 196 
<< pdiffusion >>
rect 157 195 158 196 
<< pdiffusion >>
rect 158 195 159 196 
<< pdiffusion >>
rect 159 195 160 196 
<< pdiffusion >>
rect 160 195 161 196 
<< pdiffusion >>
rect 161 195 162 196 
<< m1 >>
rect 163 195 164 196 
<< pdiffusion >>
rect 174 195 175 196 
<< pdiffusion >>
rect 175 195 176 196 
<< pdiffusion >>
rect 176 195 177 196 
<< pdiffusion >>
rect 177 195 178 196 
<< pdiffusion >>
rect 178 195 179 196 
<< pdiffusion >>
rect 179 195 180 196 
<< m1 >>
rect 185 195 186 196 
<< m1 >>
rect 187 195 188 196 
<< pdiffusion >>
rect 192 195 193 196 
<< pdiffusion >>
rect 193 195 194 196 
<< pdiffusion >>
rect 194 195 195 196 
<< pdiffusion >>
rect 195 195 196 196 
<< pdiffusion >>
rect 196 195 197 196 
<< pdiffusion >>
rect 197 195 198 196 
<< m1 >>
rect 208 195 209 196 
<< pdiffusion >>
rect 210 195 211 196 
<< pdiffusion >>
rect 211 195 212 196 
<< pdiffusion >>
rect 212 195 213 196 
<< pdiffusion >>
rect 213 195 214 196 
<< pdiffusion >>
rect 214 195 215 196 
<< pdiffusion >>
rect 215 195 216 196 
<< m1 >>
rect 219 195 220 196 
<< m1 >>
rect 221 195 222 196 
<< m1 >>
rect 224 195 225 196 
<< m1 >>
rect 226 195 227 196 
<< m1 >>
rect 235 195 236 196 
<< m1 >>
rect 237 195 238 196 
<< m2 >>
rect 241 195 242 196 
<< m1 >>
rect 242 195 243 196 
<< m1 >>
rect 244 195 245 196 
<< pdiffusion >>
rect 246 195 247 196 
<< pdiffusion >>
rect 247 195 248 196 
<< pdiffusion >>
rect 248 195 249 196 
<< pdiffusion >>
rect 249 195 250 196 
<< pdiffusion >>
rect 250 195 251 196 
<< pdiffusion >>
rect 251 195 252 196 
<< m1 >>
rect 253 195 254 196 
<< m1 >>
rect 262 195 263 196 
<< pdiffusion >>
rect 264 195 265 196 
<< pdiffusion >>
rect 265 195 266 196 
<< pdiffusion >>
rect 266 195 267 196 
<< pdiffusion >>
rect 267 195 268 196 
<< pdiffusion >>
rect 268 195 269 196 
<< pdiffusion >>
rect 269 195 270 196 
<< m1 >>
rect 278 195 279 196 
<< pdiffusion >>
rect 282 195 283 196 
<< pdiffusion >>
rect 283 195 284 196 
<< pdiffusion >>
rect 284 195 285 196 
<< pdiffusion >>
rect 285 195 286 196 
<< pdiffusion >>
rect 286 195 287 196 
<< pdiffusion >>
rect 287 195 288 196 
<< m2 >>
rect 295 195 296 196 
<< m1 >>
rect 296 195 297 196 
<< m1 >>
rect 298 195 299 196 
<< pdiffusion >>
rect 300 195 301 196 
<< pdiffusion >>
rect 301 195 302 196 
<< pdiffusion >>
rect 302 195 303 196 
<< pdiffusion >>
rect 303 195 304 196 
<< pdiffusion >>
rect 304 195 305 196 
<< pdiffusion >>
rect 305 195 306 196 
<< m1 >>
rect 308 195 309 196 
<< pdiffusion >>
rect 318 195 319 196 
<< pdiffusion >>
rect 319 195 320 196 
<< pdiffusion >>
rect 320 195 321 196 
<< pdiffusion >>
rect 321 195 322 196 
<< pdiffusion >>
rect 322 195 323 196 
<< pdiffusion >>
rect 323 195 324 196 
<< m1 >>
rect 334 195 335 196 
<< pdiffusion >>
rect 336 195 337 196 
<< pdiffusion >>
rect 337 195 338 196 
<< pdiffusion >>
rect 338 195 339 196 
<< pdiffusion >>
rect 339 195 340 196 
<< pdiffusion >>
rect 340 195 341 196 
<< pdiffusion >>
rect 341 195 342 196 
<< m1 >>
rect 343 195 344 196 
<< m1 >>
rect 352 195 353 196 
<< pdiffusion >>
rect 354 195 355 196 
<< pdiffusion >>
rect 355 195 356 196 
<< pdiffusion >>
rect 356 195 357 196 
<< pdiffusion >>
rect 357 195 358 196 
<< pdiffusion >>
rect 358 195 359 196 
<< pdiffusion >>
rect 359 195 360 196 
<< pdiffusion >>
rect 372 195 373 196 
<< pdiffusion >>
rect 373 195 374 196 
<< pdiffusion >>
rect 374 195 375 196 
<< pdiffusion >>
rect 375 195 376 196 
<< pdiffusion >>
rect 376 195 377 196 
<< pdiffusion >>
rect 377 195 378 196 
<< m1 >>
rect 379 195 380 196 
<< pdiffusion >>
rect 390 195 391 196 
<< pdiffusion >>
rect 391 195 392 196 
<< pdiffusion >>
rect 392 195 393 196 
<< pdiffusion >>
rect 393 195 394 196 
<< pdiffusion >>
rect 394 195 395 196 
<< pdiffusion >>
rect 395 195 396 196 
<< m1 >>
rect 402 195 403 196 
<< m1 >>
rect 404 195 405 196 
<< m2 >>
rect 405 195 406 196 
<< m1 >>
rect 406 195 407 196 
<< pdiffusion >>
rect 408 195 409 196 
<< pdiffusion >>
rect 409 195 410 196 
<< pdiffusion >>
rect 410 195 411 196 
<< pdiffusion >>
rect 411 195 412 196 
<< pdiffusion >>
rect 412 195 413 196 
<< pdiffusion >>
rect 413 195 414 196 
<< m1 >>
rect 415 195 416 196 
<< m1 >>
rect 417 195 418 196 
<< m1 >>
rect 419 195 420 196 
<< m1 >>
rect 423 195 424 196 
<< pdiffusion >>
rect 426 195 427 196 
<< pdiffusion >>
rect 427 195 428 196 
<< pdiffusion >>
rect 428 195 429 196 
<< pdiffusion >>
rect 429 195 430 196 
<< pdiffusion >>
rect 430 195 431 196 
<< pdiffusion >>
rect 431 195 432 196 
<< m1 >>
rect 433 195 434 196 
<< m2 >>
rect 433 195 434 196 
<< pdiffusion >>
rect 444 195 445 196 
<< pdiffusion >>
rect 445 195 446 196 
<< pdiffusion >>
rect 446 195 447 196 
<< pdiffusion >>
rect 447 195 448 196 
<< pdiffusion >>
rect 448 195 449 196 
<< pdiffusion >>
rect 449 195 450 196 
<< m1 >>
rect 456 195 457 196 
<< pdiffusion >>
rect 462 195 463 196 
<< pdiffusion >>
rect 463 195 464 196 
<< pdiffusion >>
rect 464 195 465 196 
<< pdiffusion >>
rect 465 195 466 196 
<< pdiffusion >>
rect 466 195 467 196 
<< pdiffusion >>
rect 467 195 468 196 
<< m1 >>
rect 478 195 479 196 
<< pdiffusion >>
rect 480 195 481 196 
<< pdiffusion >>
rect 481 195 482 196 
<< pdiffusion >>
rect 482 195 483 196 
<< pdiffusion >>
rect 483 195 484 196 
<< pdiffusion >>
rect 484 195 485 196 
<< pdiffusion >>
rect 485 195 486 196 
<< pdiffusion >>
rect 498 195 499 196 
<< pdiffusion >>
rect 499 195 500 196 
<< pdiffusion >>
rect 500 195 501 196 
<< pdiffusion >>
rect 501 195 502 196 
<< pdiffusion >>
rect 502 195 503 196 
<< pdiffusion >>
rect 503 195 504 196 
<< pdiffusion >>
rect 516 195 517 196 
<< pdiffusion >>
rect 517 195 518 196 
<< pdiffusion >>
rect 518 195 519 196 
<< pdiffusion >>
rect 519 195 520 196 
<< pdiffusion >>
rect 520 195 521 196 
<< pdiffusion >>
rect 521 195 522 196 
<< m1 >>
rect 28 196 29 197 
<< pdiffusion >>
rect 30 196 31 197 
<< pdiffusion >>
rect 31 196 32 197 
<< pdiffusion >>
rect 32 196 33 197 
<< pdiffusion >>
rect 33 196 34 197 
<< pdiffusion >>
rect 34 196 35 197 
<< pdiffusion >>
rect 35 196 36 197 
<< pdiffusion >>
rect 48 196 49 197 
<< pdiffusion >>
rect 49 196 50 197 
<< pdiffusion >>
rect 50 196 51 197 
<< pdiffusion >>
rect 51 196 52 197 
<< pdiffusion >>
rect 52 196 53 197 
<< pdiffusion >>
rect 53 196 54 197 
<< m1 >>
rect 64 196 65 197 
<< pdiffusion >>
rect 66 196 67 197 
<< pdiffusion >>
rect 67 196 68 197 
<< pdiffusion >>
rect 68 196 69 197 
<< pdiffusion >>
rect 69 196 70 197 
<< pdiffusion >>
rect 70 196 71 197 
<< pdiffusion >>
rect 71 196 72 197 
<< pdiffusion >>
rect 84 196 85 197 
<< pdiffusion >>
rect 85 196 86 197 
<< pdiffusion >>
rect 86 196 87 197 
<< pdiffusion >>
rect 87 196 88 197 
<< pdiffusion >>
rect 88 196 89 197 
<< pdiffusion >>
rect 89 196 90 197 
<< m1 >>
rect 98 196 99 197 
<< pdiffusion >>
rect 102 196 103 197 
<< pdiffusion >>
rect 103 196 104 197 
<< pdiffusion >>
rect 104 196 105 197 
<< pdiffusion >>
rect 105 196 106 197 
<< pdiffusion >>
rect 106 196 107 197 
<< pdiffusion >>
rect 107 196 108 197 
<< pdiffusion >>
rect 120 196 121 197 
<< pdiffusion >>
rect 121 196 122 197 
<< pdiffusion >>
rect 122 196 123 197 
<< pdiffusion >>
rect 123 196 124 197 
<< pdiffusion >>
rect 124 196 125 197 
<< pdiffusion >>
rect 125 196 126 197 
<< m1 >>
rect 127 196 128 197 
<< pdiffusion >>
rect 138 196 139 197 
<< pdiffusion >>
rect 139 196 140 197 
<< pdiffusion >>
rect 140 196 141 197 
<< pdiffusion >>
rect 141 196 142 197 
<< pdiffusion >>
rect 142 196 143 197 
<< pdiffusion >>
rect 143 196 144 197 
<< m1 >>
rect 147 196 148 197 
<< m1 >>
rect 154 196 155 197 
<< pdiffusion >>
rect 156 196 157 197 
<< pdiffusion >>
rect 157 196 158 197 
<< pdiffusion >>
rect 158 196 159 197 
<< pdiffusion >>
rect 159 196 160 197 
<< pdiffusion >>
rect 160 196 161 197 
<< pdiffusion >>
rect 161 196 162 197 
<< m1 >>
rect 163 196 164 197 
<< pdiffusion >>
rect 174 196 175 197 
<< pdiffusion >>
rect 175 196 176 197 
<< pdiffusion >>
rect 176 196 177 197 
<< pdiffusion >>
rect 177 196 178 197 
<< pdiffusion >>
rect 178 196 179 197 
<< pdiffusion >>
rect 179 196 180 197 
<< m1 >>
rect 185 196 186 197 
<< m1 >>
rect 187 196 188 197 
<< pdiffusion >>
rect 192 196 193 197 
<< pdiffusion >>
rect 193 196 194 197 
<< pdiffusion >>
rect 194 196 195 197 
<< pdiffusion >>
rect 195 196 196 197 
<< pdiffusion >>
rect 196 196 197 197 
<< pdiffusion >>
rect 197 196 198 197 
<< m1 >>
rect 208 196 209 197 
<< pdiffusion >>
rect 210 196 211 197 
<< pdiffusion >>
rect 211 196 212 197 
<< pdiffusion >>
rect 212 196 213 197 
<< pdiffusion >>
rect 213 196 214 197 
<< pdiffusion >>
rect 214 196 215 197 
<< pdiffusion >>
rect 215 196 216 197 
<< m1 >>
rect 219 196 220 197 
<< m1 >>
rect 221 196 222 197 
<< m1 >>
rect 224 196 225 197 
<< m1 >>
rect 226 196 227 197 
<< m1 >>
rect 235 196 236 197 
<< m1 >>
rect 237 196 238 197 
<< m2 >>
rect 241 196 242 197 
<< m1 >>
rect 242 196 243 197 
<< m1 >>
rect 244 196 245 197 
<< pdiffusion >>
rect 246 196 247 197 
<< pdiffusion >>
rect 247 196 248 197 
<< pdiffusion >>
rect 248 196 249 197 
<< pdiffusion >>
rect 249 196 250 197 
<< pdiffusion >>
rect 250 196 251 197 
<< pdiffusion >>
rect 251 196 252 197 
<< m1 >>
rect 253 196 254 197 
<< m1 >>
rect 262 196 263 197 
<< pdiffusion >>
rect 264 196 265 197 
<< pdiffusion >>
rect 265 196 266 197 
<< pdiffusion >>
rect 266 196 267 197 
<< pdiffusion >>
rect 267 196 268 197 
<< pdiffusion >>
rect 268 196 269 197 
<< pdiffusion >>
rect 269 196 270 197 
<< m1 >>
rect 278 196 279 197 
<< pdiffusion >>
rect 282 196 283 197 
<< pdiffusion >>
rect 283 196 284 197 
<< pdiffusion >>
rect 284 196 285 197 
<< pdiffusion >>
rect 285 196 286 197 
<< pdiffusion >>
rect 286 196 287 197 
<< pdiffusion >>
rect 287 196 288 197 
<< m2 >>
rect 295 196 296 197 
<< m1 >>
rect 296 196 297 197 
<< m1 >>
rect 298 196 299 197 
<< pdiffusion >>
rect 300 196 301 197 
<< pdiffusion >>
rect 301 196 302 197 
<< pdiffusion >>
rect 302 196 303 197 
<< pdiffusion >>
rect 303 196 304 197 
<< pdiffusion >>
rect 304 196 305 197 
<< pdiffusion >>
rect 305 196 306 197 
<< m1 >>
rect 308 196 309 197 
<< pdiffusion >>
rect 318 196 319 197 
<< pdiffusion >>
rect 319 196 320 197 
<< pdiffusion >>
rect 320 196 321 197 
<< pdiffusion >>
rect 321 196 322 197 
<< pdiffusion >>
rect 322 196 323 197 
<< pdiffusion >>
rect 323 196 324 197 
<< m1 >>
rect 334 196 335 197 
<< pdiffusion >>
rect 336 196 337 197 
<< pdiffusion >>
rect 337 196 338 197 
<< pdiffusion >>
rect 338 196 339 197 
<< pdiffusion >>
rect 339 196 340 197 
<< pdiffusion >>
rect 340 196 341 197 
<< pdiffusion >>
rect 341 196 342 197 
<< m1 >>
rect 343 196 344 197 
<< m1 >>
rect 352 196 353 197 
<< pdiffusion >>
rect 354 196 355 197 
<< pdiffusion >>
rect 355 196 356 197 
<< pdiffusion >>
rect 356 196 357 197 
<< pdiffusion >>
rect 357 196 358 197 
<< pdiffusion >>
rect 358 196 359 197 
<< pdiffusion >>
rect 359 196 360 197 
<< pdiffusion >>
rect 372 196 373 197 
<< pdiffusion >>
rect 373 196 374 197 
<< pdiffusion >>
rect 374 196 375 197 
<< pdiffusion >>
rect 375 196 376 197 
<< pdiffusion >>
rect 376 196 377 197 
<< pdiffusion >>
rect 377 196 378 197 
<< m1 >>
rect 379 196 380 197 
<< pdiffusion >>
rect 390 196 391 197 
<< pdiffusion >>
rect 391 196 392 197 
<< pdiffusion >>
rect 392 196 393 197 
<< pdiffusion >>
rect 393 196 394 197 
<< pdiffusion >>
rect 394 196 395 197 
<< pdiffusion >>
rect 395 196 396 197 
<< m1 >>
rect 402 196 403 197 
<< m1 >>
rect 404 196 405 197 
<< m2 >>
rect 405 196 406 197 
<< m1 >>
rect 406 196 407 197 
<< pdiffusion >>
rect 408 196 409 197 
<< pdiffusion >>
rect 409 196 410 197 
<< pdiffusion >>
rect 410 196 411 197 
<< pdiffusion >>
rect 411 196 412 197 
<< pdiffusion >>
rect 412 196 413 197 
<< pdiffusion >>
rect 413 196 414 197 
<< m1 >>
rect 415 196 416 197 
<< m1 >>
rect 417 196 418 197 
<< m1 >>
rect 419 196 420 197 
<< m1 >>
rect 423 196 424 197 
<< pdiffusion >>
rect 426 196 427 197 
<< pdiffusion >>
rect 427 196 428 197 
<< pdiffusion >>
rect 428 196 429 197 
<< pdiffusion >>
rect 429 196 430 197 
<< pdiffusion >>
rect 430 196 431 197 
<< pdiffusion >>
rect 431 196 432 197 
<< m1 >>
rect 433 196 434 197 
<< m2 >>
rect 433 196 434 197 
<< pdiffusion >>
rect 444 196 445 197 
<< pdiffusion >>
rect 445 196 446 197 
<< pdiffusion >>
rect 446 196 447 197 
<< pdiffusion >>
rect 447 196 448 197 
<< pdiffusion >>
rect 448 196 449 197 
<< pdiffusion >>
rect 449 196 450 197 
<< m1 >>
rect 456 196 457 197 
<< pdiffusion >>
rect 462 196 463 197 
<< pdiffusion >>
rect 463 196 464 197 
<< pdiffusion >>
rect 464 196 465 197 
<< pdiffusion >>
rect 465 196 466 197 
<< pdiffusion >>
rect 466 196 467 197 
<< pdiffusion >>
rect 467 196 468 197 
<< m1 >>
rect 478 196 479 197 
<< pdiffusion >>
rect 480 196 481 197 
<< pdiffusion >>
rect 481 196 482 197 
<< pdiffusion >>
rect 482 196 483 197 
<< pdiffusion >>
rect 483 196 484 197 
<< pdiffusion >>
rect 484 196 485 197 
<< pdiffusion >>
rect 485 196 486 197 
<< pdiffusion >>
rect 498 196 499 197 
<< pdiffusion >>
rect 499 196 500 197 
<< pdiffusion >>
rect 500 196 501 197 
<< pdiffusion >>
rect 501 196 502 197 
<< pdiffusion >>
rect 502 196 503 197 
<< pdiffusion >>
rect 503 196 504 197 
<< pdiffusion >>
rect 516 196 517 197 
<< pdiffusion >>
rect 517 196 518 197 
<< pdiffusion >>
rect 518 196 519 197 
<< pdiffusion >>
rect 519 196 520 197 
<< pdiffusion >>
rect 520 196 521 197 
<< pdiffusion >>
rect 521 196 522 197 
<< m1 >>
rect 28 197 29 198 
<< pdiffusion >>
rect 30 197 31 198 
<< pdiffusion >>
rect 31 197 32 198 
<< pdiffusion >>
rect 32 197 33 198 
<< pdiffusion >>
rect 33 197 34 198 
<< pdiffusion >>
rect 34 197 35 198 
<< pdiffusion >>
rect 35 197 36 198 
<< pdiffusion >>
rect 48 197 49 198 
<< pdiffusion >>
rect 49 197 50 198 
<< pdiffusion >>
rect 50 197 51 198 
<< pdiffusion >>
rect 51 197 52 198 
<< pdiffusion >>
rect 52 197 53 198 
<< pdiffusion >>
rect 53 197 54 198 
<< m1 >>
rect 64 197 65 198 
<< pdiffusion >>
rect 66 197 67 198 
<< pdiffusion >>
rect 67 197 68 198 
<< pdiffusion >>
rect 68 197 69 198 
<< pdiffusion >>
rect 69 197 70 198 
<< pdiffusion >>
rect 70 197 71 198 
<< pdiffusion >>
rect 71 197 72 198 
<< pdiffusion >>
rect 84 197 85 198 
<< pdiffusion >>
rect 85 197 86 198 
<< pdiffusion >>
rect 86 197 87 198 
<< pdiffusion >>
rect 87 197 88 198 
<< pdiffusion >>
rect 88 197 89 198 
<< pdiffusion >>
rect 89 197 90 198 
<< m1 >>
rect 98 197 99 198 
<< pdiffusion >>
rect 102 197 103 198 
<< pdiffusion >>
rect 103 197 104 198 
<< pdiffusion >>
rect 104 197 105 198 
<< pdiffusion >>
rect 105 197 106 198 
<< m1 >>
rect 106 197 107 198 
<< pdiffusion >>
rect 106 197 107 198 
<< pdiffusion >>
rect 107 197 108 198 
<< pdiffusion >>
rect 120 197 121 198 
<< m1 >>
rect 121 197 122 198 
<< pdiffusion >>
rect 121 197 122 198 
<< pdiffusion >>
rect 122 197 123 198 
<< pdiffusion >>
rect 123 197 124 198 
<< pdiffusion >>
rect 124 197 125 198 
<< pdiffusion >>
rect 125 197 126 198 
<< m1 >>
rect 127 197 128 198 
<< pdiffusion >>
rect 138 197 139 198 
<< pdiffusion >>
rect 139 197 140 198 
<< pdiffusion >>
rect 140 197 141 198 
<< pdiffusion >>
rect 141 197 142 198 
<< pdiffusion >>
rect 142 197 143 198 
<< pdiffusion >>
rect 143 197 144 198 
<< m1 >>
rect 147 197 148 198 
<< m1 >>
rect 154 197 155 198 
<< pdiffusion >>
rect 156 197 157 198 
<< m1 >>
rect 157 197 158 198 
<< pdiffusion >>
rect 157 197 158 198 
<< pdiffusion >>
rect 158 197 159 198 
<< pdiffusion >>
rect 159 197 160 198 
<< pdiffusion >>
rect 160 197 161 198 
<< pdiffusion >>
rect 161 197 162 198 
<< m1 >>
rect 163 197 164 198 
<< pdiffusion >>
rect 174 197 175 198 
<< pdiffusion >>
rect 175 197 176 198 
<< pdiffusion >>
rect 176 197 177 198 
<< pdiffusion >>
rect 177 197 178 198 
<< m1 >>
rect 178 197 179 198 
<< pdiffusion >>
rect 178 197 179 198 
<< pdiffusion >>
rect 179 197 180 198 
<< m1 >>
rect 185 197 186 198 
<< m1 >>
rect 187 197 188 198 
<< pdiffusion >>
rect 192 197 193 198 
<< pdiffusion >>
rect 193 197 194 198 
<< pdiffusion >>
rect 194 197 195 198 
<< pdiffusion >>
rect 195 197 196 198 
<< pdiffusion >>
rect 196 197 197 198 
<< pdiffusion >>
rect 197 197 198 198 
<< m1 >>
rect 208 197 209 198 
<< pdiffusion >>
rect 210 197 211 198 
<< pdiffusion >>
rect 211 197 212 198 
<< pdiffusion >>
rect 212 197 213 198 
<< pdiffusion >>
rect 213 197 214 198 
<< m1 >>
rect 214 197 215 198 
<< pdiffusion >>
rect 214 197 215 198 
<< pdiffusion >>
rect 215 197 216 198 
<< m1 >>
rect 219 197 220 198 
<< m2 >>
rect 219 197 220 198 
<< m2c >>
rect 219 197 220 198 
<< m1 >>
rect 219 197 220 198 
<< m2 >>
rect 219 197 220 198 
<< m1 >>
rect 221 197 222 198 
<< m2 >>
rect 221 197 222 198 
<< m2c >>
rect 221 197 222 198 
<< m1 >>
rect 221 197 222 198 
<< m2 >>
rect 221 197 222 198 
<< m1 >>
rect 224 197 225 198 
<< m1 >>
rect 226 197 227 198 
<< m1 >>
rect 235 197 236 198 
<< m1 >>
rect 237 197 238 198 
<< m2 >>
rect 241 197 242 198 
<< m1 >>
rect 242 197 243 198 
<< m1 >>
rect 244 197 245 198 
<< pdiffusion >>
rect 246 197 247 198 
<< pdiffusion >>
rect 247 197 248 198 
<< pdiffusion >>
rect 248 197 249 198 
<< pdiffusion >>
rect 249 197 250 198 
<< pdiffusion >>
rect 250 197 251 198 
<< pdiffusion >>
rect 251 197 252 198 
<< m1 >>
rect 253 197 254 198 
<< m1 >>
rect 262 197 263 198 
<< pdiffusion >>
rect 264 197 265 198 
<< pdiffusion >>
rect 265 197 266 198 
<< pdiffusion >>
rect 266 197 267 198 
<< pdiffusion >>
rect 267 197 268 198 
<< pdiffusion >>
rect 268 197 269 198 
<< pdiffusion >>
rect 269 197 270 198 
<< m1 >>
rect 278 197 279 198 
<< pdiffusion >>
rect 282 197 283 198 
<< m1 >>
rect 283 197 284 198 
<< pdiffusion >>
rect 283 197 284 198 
<< pdiffusion >>
rect 284 197 285 198 
<< pdiffusion >>
rect 285 197 286 198 
<< pdiffusion >>
rect 286 197 287 198 
<< pdiffusion >>
rect 287 197 288 198 
<< m2 >>
rect 295 197 296 198 
<< m1 >>
rect 296 197 297 198 
<< m1 >>
rect 298 197 299 198 
<< pdiffusion >>
rect 300 197 301 198 
<< pdiffusion >>
rect 301 197 302 198 
<< pdiffusion >>
rect 302 197 303 198 
<< pdiffusion >>
rect 303 197 304 198 
<< m1 >>
rect 304 197 305 198 
<< pdiffusion >>
rect 304 197 305 198 
<< pdiffusion >>
rect 305 197 306 198 
<< m1 >>
rect 308 197 309 198 
<< pdiffusion >>
rect 318 197 319 198 
<< m1 >>
rect 319 197 320 198 
<< pdiffusion >>
rect 319 197 320 198 
<< pdiffusion >>
rect 320 197 321 198 
<< pdiffusion >>
rect 321 197 322 198 
<< m1 >>
rect 322 197 323 198 
<< pdiffusion >>
rect 322 197 323 198 
<< pdiffusion >>
rect 323 197 324 198 
<< m1 >>
rect 334 197 335 198 
<< pdiffusion >>
rect 336 197 337 198 
<< m1 >>
rect 337 197 338 198 
<< pdiffusion >>
rect 337 197 338 198 
<< pdiffusion >>
rect 338 197 339 198 
<< pdiffusion >>
rect 339 197 340 198 
<< pdiffusion >>
rect 340 197 341 198 
<< pdiffusion >>
rect 341 197 342 198 
<< m1 >>
rect 343 197 344 198 
<< m1 >>
rect 352 197 353 198 
<< m2 >>
rect 352 197 353 198 
<< m2c >>
rect 352 197 353 198 
<< m1 >>
rect 352 197 353 198 
<< m2 >>
rect 352 197 353 198 
<< pdiffusion >>
rect 354 197 355 198 
<< m1 >>
rect 355 197 356 198 
<< pdiffusion >>
rect 355 197 356 198 
<< pdiffusion >>
rect 356 197 357 198 
<< pdiffusion >>
rect 357 197 358 198 
<< pdiffusion >>
rect 358 197 359 198 
<< pdiffusion >>
rect 359 197 360 198 
<< pdiffusion >>
rect 372 197 373 198 
<< pdiffusion >>
rect 373 197 374 198 
<< pdiffusion >>
rect 374 197 375 198 
<< pdiffusion >>
rect 375 197 376 198 
<< pdiffusion >>
rect 376 197 377 198 
<< pdiffusion >>
rect 377 197 378 198 
<< m1 >>
rect 379 197 380 198 
<< pdiffusion >>
rect 390 197 391 198 
<< pdiffusion >>
rect 391 197 392 198 
<< pdiffusion >>
rect 392 197 393 198 
<< pdiffusion >>
rect 393 197 394 198 
<< m1 >>
rect 394 197 395 198 
<< pdiffusion >>
rect 394 197 395 198 
<< pdiffusion >>
rect 395 197 396 198 
<< m1 >>
rect 402 197 403 198 
<< m1 >>
rect 404 197 405 198 
<< m2 >>
rect 405 197 406 198 
<< m1 >>
rect 406 197 407 198 
<< pdiffusion >>
rect 408 197 409 198 
<< pdiffusion >>
rect 409 197 410 198 
<< pdiffusion >>
rect 410 197 411 198 
<< pdiffusion >>
rect 411 197 412 198 
<< pdiffusion >>
rect 412 197 413 198 
<< pdiffusion >>
rect 413 197 414 198 
<< m1 >>
rect 415 197 416 198 
<< m1 >>
rect 417 197 418 198 
<< m1 >>
rect 419 197 420 198 
<< m1 >>
rect 423 197 424 198 
<< pdiffusion >>
rect 426 197 427 198 
<< pdiffusion >>
rect 427 197 428 198 
<< pdiffusion >>
rect 428 197 429 198 
<< pdiffusion >>
rect 429 197 430 198 
<< m1 >>
rect 430 197 431 198 
<< pdiffusion >>
rect 430 197 431 198 
<< pdiffusion >>
rect 431 197 432 198 
<< m1 >>
rect 433 197 434 198 
<< m2 >>
rect 433 197 434 198 
<< pdiffusion >>
rect 444 197 445 198 
<< m1 >>
rect 445 197 446 198 
<< pdiffusion >>
rect 445 197 446 198 
<< pdiffusion >>
rect 446 197 447 198 
<< pdiffusion >>
rect 447 197 448 198 
<< m1 >>
rect 448 197 449 198 
<< pdiffusion >>
rect 448 197 449 198 
<< pdiffusion >>
rect 449 197 450 198 
<< m1 >>
rect 456 197 457 198 
<< pdiffusion >>
rect 462 197 463 198 
<< pdiffusion >>
rect 463 197 464 198 
<< pdiffusion >>
rect 464 197 465 198 
<< pdiffusion >>
rect 465 197 466 198 
<< pdiffusion >>
rect 466 197 467 198 
<< pdiffusion >>
rect 467 197 468 198 
<< m1 >>
rect 478 197 479 198 
<< pdiffusion >>
rect 480 197 481 198 
<< pdiffusion >>
rect 481 197 482 198 
<< pdiffusion >>
rect 482 197 483 198 
<< pdiffusion >>
rect 483 197 484 198 
<< pdiffusion >>
rect 484 197 485 198 
<< pdiffusion >>
rect 485 197 486 198 
<< pdiffusion >>
rect 498 197 499 198 
<< pdiffusion >>
rect 499 197 500 198 
<< pdiffusion >>
rect 500 197 501 198 
<< pdiffusion >>
rect 501 197 502 198 
<< pdiffusion >>
rect 502 197 503 198 
<< pdiffusion >>
rect 503 197 504 198 
<< pdiffusion >>
rect 516 197 517 198 
<< pdiffusion >>
rect 517 197 518 198 
<< pdiffusion >>
rect 518 197 519 198 
<< pdiffusion >>
rect 519 197 520 198 
<< pdiffusion >>
rect 520 197 521 198 
<< pdiffusion >>
rect 521 197 522 198 
<< m1 >>
rect 28 198 29 199 
<< m1 >>
rect 64 198 65 199 
<< m1 >>
rect 98 198 99 199 
<< m1 >>
rect 106 198 107 199 
<< m1 >>
rect 121 198 122 199 
<< m1 >>
rect 127 198 128 199 
<< m1 >>
rect 147 198 148 199 
<< m1 >>
rect 154 198 155 199 
<< m1 >>
rect 157 198 158 199 
<< m1 >>
rect 163 198 164 199 
<< m1 >>
rect 178 198 179 199 
<< m1 >>
rect 185 198 186 199 
<< m1 >>
rect 187 198 188 199 
<< m1 >>
rect 208 198 209 199 
<< m1 >>
rect 214 198 215 199 
<< m2 >>
rect 219 198 220 199 
<< m2 >>
rect 221 198 222 199 
<< m1 >>
rect 224 198 225 199 
<< m1 >>
rect 226 198 227 199 
<< m1 >>
rect 235 198 236 199 
<< m1 >>
rect 237 198 238 199 
<< m1 >>
rect 239 198 240 199 
<< m1 >>
rect 240 198 241 199 
<< m2 >>
rect 240 198 241 199 
<< m2c >>
rect 240 198 241 199 
<< m1 >>
rect 240 198 241 199 
<< m2 >>
rect 240 198 241 199 
<< m2 >>
rect 241 198 242 199 
<< m1 >>
rect 242 198 243 199 
<< m1 >>
rect 244 198 245 199 
<< m1 >>
rect 253 198 254 199 
<< m1 >>
rect 262 198 263 199 
<< m1 >>
rect 278 198 279 199 
<< m1 >>
rect 283 198 284 199 
<< m2 >>
rect 295 198 296 199 
<< m1 >>
rect 296 198 297 199 
<< m1 >>
rect 298 198 299 199 
<< m1 >>
rect 304 198 305 199 
<< m1 >>
rect 308 198 309 199 
<< m1 >>
rect 319 198 320 199 
<< m1 >>
rect 322 198 323 199 
<< m1 >>
rect 334 198 335 199 
<< m1 >>
rect 337 198 338 199 
<< m1 >>
rect 343 198 344 199 
<< m2 >>
rect 352 198 353 199 
<< m1 >>
rect 355 198 356 199 
<< m1 >>
rect 379 198 380 199 
<< m1 >>
rect 394 198 395 199 
<< m1 >>
rect 402 198 403 199 
<< m1 >>
rect 404 198 405 199 
<< m2 >>
rect 405 198 406 199 
<< m1 >>
rect 406 198 407 199 
<< m1 >>
rect 415 198 416 199 
<< m1 >>
rect 417 198 418 199 
<< m1 >>
rect 419 198 420 199 
<< m1 >>
rect 423 198 424 199 
<< m1 >>
rect 430 198 431 199 
<< m1 >>
rect 433 198 434 199 
<< m2 >>
rect 433 198 434 199 
<< m1 >>
rect 445 198 446 199 
<< m1 >>
rect 448 198 449 199 
<< m1 >>
rect 456 198 457 199 
<< m1 >>
rect 478 198 479 199 
<< m1 >>
rect 28 199 29 200 
<< m1 >>
rect 64 199 65 200 
<< m1 >>
rect 98 199 99 200 
<< m1 >>
rect 106 199 107 200 
<< m2 >>
rect 107 199 108 200 
<< m1 >>
rect 108 199 109 200 
<< m2 >>
rect 108 199 109 200 
<< m2c >>
rect 108 199 109 200 
<< m1 >>
rect 108 199 109 200 
<< m2 >>
rect 108 199 109 200 
<< m1 >>
rect 109 199 110 200 
<< m1 >>
rect 110 199 111 200 
<< m1 >>
rect 111 199 112 200 
<< m1 >>
rect 112 199 113 200 
<< m1 >>
rect 113 199 114 200 
<< m1 >>
rect 114 199 115 200 
<< m1 >>
rect 115 199 116 200 
<< m1 >>
rect 116 199 117 200 
<< m1 >>
rect 117 199 118 200 
<< m1 >>
rect 118 199 119 200 
<< m1 >>
rect 119 199 120 200 
<< m1 >>
rect 120 199 121 200 
<< m1 >>
rect 121 199 122 200 
<< m1 >>
rect 127 199 128 200 
<< m1 >>
rect 147 199 148 200 
<< m1 >>
rect 154 199 155 200 
<< m1 >>
rect 155 199 156 200 
<< m1 >>
rect 156 199 157 200 
<< m1 >>
rect 157 199 158 200 
<< m1 >>
rect 163 199 164 200 
<< m1 >>
rect 178 199 179 200 
<< m1 >>
rect 179 199 180 200 
<< m1 >>
rect 180 199 181 200 
<< m1 >>
rect 181 199 182 200 
<< m1 >>
rect 185 199 186 200 
<< m1 >>
rect 187 199 188 200 
<< m1 >>
rect 208 199 209 200 
<< m1 >>
rect 214 199 215 200 
<< m2 >>
rect 215 199 216 200 
<< m1 >>
rect 216 199 217 200 
<< m2 >>
rect 216 199 217 200 
<< m2c >>
rect 216 199 217 200 
<< m1 >>
rect 216 199 217 200 
<< m2 >>
rect 216 199 217 200 
<< m1 >>
rect 217 199 218 200 
<< m1 >>
rect 218 199 219 200 
<< m1 >>
rect 219 199 220 200 
<< m2 >>
rect 219 199 220 200 
<< m1 >>
rect 220 199 221 200 
<< m1 >>
rect 221 199 222 200 
<< m2 >>
rect 221 199 222 200 
<< m1 >>
rect 222 199 223 200 
<< m1 >>
rect 223 199 224 200 
<< m1 >>
rect 224 199 225 200 
<< m1 >>
rect 226 199 227 200 
<< m1 >>
rect 235 199 236 200 
<< m1 >>
rect 237 199 238 200 
<< m1 >>
rect 239 199 240 200 
<< m1 >>
rect 242 199 243 200 
<< m1 >>
rect 244 199 245 200 
<< m1 >>
rect 253 199 254 200 
<< m1 >>
rect 262 199 263 200 
<< m1 >>
rect 278 199 279 200 
<< m1 >>
rect 279 199 280 200 
<< m1 >>
rect 280 199 281 200 
<< m1 >>
rect 281 199 282 200 
<< m1 >>
rect 282 199 283 200 
<< m1 >>
rect 283 199 284 200 
<< m2 >>
rect 295 199 296 200 
<< m1 >>
rect 296 199 297 200 
<< m1 >>
rect 298 199 299 200 
<< m1 >>
rect 304 199 305 200 
<< m1 >>
rect 308 199 309 200 
<< m1 >>
rect 316 199 317 200 
<< m1 >>
rect 317 199 318 200 
<< m1 >>
rect 318 199 319 200 
<< m1 >>
rect 319 199 320 200 
<< m1 >>
rect 322 199 323 200 
<< m1 >>
rect 334 199 335 200 
<< m1 >>
rect 337 199 338 200 
<< m1 >>
rect 341 199 342 200 
<< m2 >>
rect 341 199 342 200 
<< m2c >>
rect 341 199 342 200 
<< m1 >>
rect 341 199 342 200 
<< m2 >>
rect 341 199 342 200 
<< m2 >>
rect 342 199 343 200 
<< m1 >>
rect 343 199 344 200 
<< m2 >>
rect 343 199 344 200 
<< m1 >>
rect 344 199 345 200 
<< m2 >>
rect 344 199 345 200 
<< m1 >>
rect 345 199 346 200 
<< m2 >>
rect 345 199 346 200 
<< m1 >>
rect 346 199 347 200 
<< m2 >>
rect 346 199 347 200 
<< m1 >>
rect 347 199 348 200 
<< m2 >>
rect 347 199 348 200 
<< m1 >>
rect 348 199 349 200 
<< m2 >>
rect 348 199 349 200 
<< m1 >>
rect 349 199 350 200 
<< m2 >>
rect 349 199 350 200 
<< m1 >>
rect 350 199 351 200 
<< m2 >>
rect 350 199 351 200 
<< m1 >>
rect 351 199 352 200 
<< m2 >>
rect 351 199 352 200 
<< m1 >>
rect 352 199 353 200 
<< m2 >>
rect 352 199 353 200 
<< m1 >>
rect 353 199 354 200 
<< m1 >>
rect 354 199 355 200 
<< m1 >>
rect 355 199 356 200 
<< m1 >>
rect 379 199 380 200 
<< m1 >>
rect 394 199 395 200 
<< m1 >>
rect 402 199 403 200 
<< m1 >>
rect 404 199 405 200 
<< m2 >>
rect 405 199 406 200 
<< m1 >>
rect 406 199 407 200 
<< m1 >>
rect 415 199 416 200 
<< m1 >>
rect 417 199 418 200 
<< m1 >>
rect 419 199 420 200 
<< m1 >>
rect 423 199 424 200 
<< m1 >>
rect 430 199 431 200 
<< m1 >>
rect 433 199 434 200 
<< m2 >>
rect 433 199 434 200 
<< m1 >>
rect 434 199 435 200 
<< m1 >>
rect 435 199 436 200 
<< m1 >>
rect 436 199 437 200 
<< m1 >>
rect 437 199 438 200 
<< m1 >>
rect 438 199 439 200 
<< m1 >>
rect 439 199 440 200 
<< m1 >>
rect 440 199 441 200 
<< m1 >>
rect 441 199 442 200 
<< m1 >>
rect 442 199 443 200 
<< m1 >>
rect 443 199 444 200 
<< m1 >>
rect 444 199 445 200 
<< m1 >>
rect 445 199 446 200 
<< m1 >>
rect 448 199 449 200 
<< m1 >>
rect 456 199 457 200 
<< m1 >>
rect 478 199 479 200 
<< m1 >>
rect 28 200 29 201 
<< m1 >>
rect 64 200 65 201 
<< m1 >>
rect 98 200 99 201 
<< m1 >>
rect 106 200 107 201 
<< m2 >>
rect 107 200 108 201 
<< m1 >>
rect 127 200 128 201 
<< m1 >>
rect 147 200 148 201 
<< m2 >>
rect 147 200 148 201 
<< m2c >>
rect 147 200 148 201 
<< m1 >>
rect 147 200 148 201 
<< m2 >>
rect 147 200 148 201 
<< m1 >>
rect 163 200 164 201 
<< m2 >>
rect 163 200 164 201 
<< m2c >>
rect 163 200 164 201 
<< m1 >>
rect 163 200 164 201 
<< m2 >>
rect 163 200 164 201 
<< m1 >>
rect 181 200 182 201 
<< m1 >>
rect 185 200 186 201 
<< m2 >>
rect 185 200 186 201 
<< m2c >>
rect 185 200 186 201 
<< m1 >>
rect 185 200 186 201 
<< m2 >>
rect 185 200 186 201 
<< m1 >>
rect 187 200 188 201 
<< m2 >>
rect 187 200 188 201 
<< m2c >>
rect 187 200 188 201 
<< m1 >>
rect 187 200 188 201 
<< m2 >>
rect 187 200 188 201 
<< m1 >>
rect 208 200 209 201 
<< m1 >>
rect 212 200 213 201 
<< m2 >>
rect 212 200 213 201 
<< m2c >>
rect 212 200 213 201 
<< m1 >>
rect 212 200 213 201 
<< m2 >>
rect 212 200 213 201 
<< m2 >>
rect 213 200 214 201 
<< m1 >>
rect 214 200 215 201 
<< m2 >>
rect 214 200 215 201 
<< m2 >>
rect 215 200 216 201 
<< m2 >>
rect 219 200 220 201 
<< m2 >>
rect 221 200 222 201 
<< m1 >>
rect 226 200 227 201 
<< m2 >>
rect 234 200 235 201 
<< m1 >>
rect 235 200 236 201 
<< m2 >>
rect 235 200 236 201 
<< m2 >>
rect 236 200 237 201 
<< m1 >>
rect 237 200 238 201 
<< m2 >>
rect 237 200 238 201 
<< m2 >>
rect 238 200 239 201 
<< m1 >>
rect 239 200 240 201 
<< m2 >>
rect 239 200 240 201 
<< m2c >>
rect 239 200 240 201 
<< m1 >>
rect 239 200 240 201 
<< m2 >>
rect 239 200 240 201 
<< m1 >>
rect 242 200 243 201 
<< m2 >>
rect 242 200 243 201 
<< m2c >>
rect 242 200 243 201 
<< m1 >>
rect 242 200 243 201 
<< m2 >>
rect 242 200 243 201 
<< m1 >>
rect 244 200 245 201 
<< m2 >>
rect 244 200 245 201 
<< m2c >>
rect 244 200 245 201 
<< m1 >>
rect 244 200 245 201 
<< m2 >>
rect 244 200 245 201 
<< m1 >>
rect 253 200 254 201 
<< m2 >>
rect 253 200 254 201 
<< m2c >>
rect 253 200 254 201 
<< m1 >>
rect 253 200 254 201 
<< m2 >>
rect 253 200 254 201 
<< m1 >>
rect 262 200 263 201 
<< m2 >>
rect 262 200 263 201 
<< m2c >>
rect 262 200 263 201 
<< m1 >>
rect 262 200 263 201 
<< m2 >>
rect 262 200 263 201 
<< m2 >>
rect 295 200 296 201 
<< m1 >>
rect 296 200 297 201 
<< m1 >>
rect 298 200 299 201 
<< m1 >>
rect 304 200 305 201 
<< m1 >>
rect 308 200 309 201 
<< m2 >>
rect 308 200 309 201 
<< m2c >>
rect 308 200 309 201 
<< m1 >>
rect 308 200 309 201 
<< m2 >>
rect 308 200 309 201 
<< m1 >>
rect 316 200 317 201 
<< m1 >>
rect 322 200 323 201 
<< m1 >>
rect 323 200 324 201 
<< m1 >>
rect 324 200 325 201 
<< m1 >>
rect 325 200 326 201 
<< m1 >>
rect 326 200 327 201 
<< m1 >>
rect 327 200 328 201 
<< m1 >>
rect 328 200 329 201 
<< m1 >>
rect 329 200 330 201 
<< m1 >>
rect 330 200 331 201 
<< m2 >>
rect 330 200 331 201 
<< m2c >>
rect 330 200 331 201 
<< m1 >>
rect 330 200 331 201 
<< m2 >>
rect 330 200 331 201 
<< m1 >>
rect 334 200 335 201 
<< m1 >>
rect 337 200 338 201 
<< m1 >>
rect 338 200 339 201 
<< m1 >>
rect 339 200 340 201 
<< m1 >>
rect 340 200 341 201 
<< m1 >>
rect 341 200 342 201 
<< m1 >>
rect 379 200 380 201 
<< m1 >>
rect 394 200 395 201 
<< m1 >>
rect 402 200 403 201 
<< m1 >>
rect 404 200 405 201 
<< m2 >>
rect 405 200 406 201 
<< m1 >>
rect 406 200 407 201 
<< m1 >>
rect 415 200 416 201 
<< m1 >>
rect 417 200 418 201 
<< m1 >>
rect 419 200 420 201 
<< m1 >>
rect 423 200 424 201 
<< m2 >>
rect 423 200 424 201 
<< m2c >>
rect 423 200 424 201 
<< m1 >>
rect 423 200 424 201 
<< m2 >>
rect 423 200 424 201 
<< m1 >>
rect 430 200 431 201 
<< m2 >>
rect 433 200 434 201 
<< m1 >>
rect 448 200 449 201 
<< m1 >>
rect 456 200 457 201 
<< m1 >>
rect 478 200 479 201 
<< m1 >>
rect 28 201 29 202 
<< m1 >>
rect 64 201 65 202 
<< m1 >>
rect 98 201 99 202 
<< m1 >>
rect 106 201 107 202 
<< m2 >>
rect 107 201 108 202 
<< m1 >>
rect 127 201 128 202 
<< m2 >>
rect 147 201 148 202 
<< m2 >>
rect 163 201 164 202 
<< m1 >>
rect 181 201 182 202 
<< m2 >>
rect 185 201 186 202 
<< m2 >>
rect 187 201 188 202 
<< m1 >>
rect 208 201 209 202 
<< m1 >>
rect 212 201 213 202 
<< m1 >>
rect 214 201 215 202 
<< m1 >>
rect 219 201 220 202 
<< m2 >>
rect 219 201 220 202 
<< m2c >>
rect 219 201 220 202 
<< m1 >>
rect 219 201 220 202 
<< m2 >>
rect 219 201 220 202 
<< m1 >>
rect 221 201 222 202 
<< m2 >>
rect 221 201 222 202 
<< m2c >>
rect 221 201 222 202 
<< m1 >>
rect 221 201 222 202 
<< m2 >>
rect 221 201 222 202 
<< m1 >>
rect 226 201 227 202 
<< m2 >>
rect 234 201 235 202 
<< m1 >>
rect 235 201 236 202 
<< m1 >>
rect 237 201 238 202 
<< m2 >>
rect 242 201 243 202 
<< m2 >>
rect 244 201 245 202 
<< m2 >>
rect 253 201 254 202 
<< m2 >>
rect 262 201 263 202 
<< m2 >>
rect 295 201 296 202 
<< m1 >>
rect 296 201 297 202 
<< m1 >>
rect 298 201 299 202 
<< m1 >>
rect 304 201 305 202 
<< m2 >>
rect 308 201 309 202 
<< m1 >>
rect 316 201 317 202 
<< m2 >>
rect 330 201 331 202 
<< m1 >>
rect 334 201 335 202 
<< m1 >>
rect 379 201 380 202 
<< m1 >>
rect 394 201 395 202 
<< m1 >>
rect 402 201 403 202 
<< m1 >>
rect 404 201 405 202 
<< m2 >>
rect 405 201 406 202 
<< m1 >>
rect 406 201 407 202 
<< m1 >>
rect 415 201 416 202 
<< m1 >>
rect 417 201 418 202 
<< m1 >>
rect 419 201 420 202 
<< m2 >>
rect 423 201 424 202 
<< m1 >>
rect 430 201 431 202 
<< m1 >>
rect 433 201 434 202 
<< m2 >>
rect 433 201 434 202 
<< m2c >>
rect 433 201 434 202 
<< m1 >>
rect 433 201 434 202 
<< m2 >>
rect 433 201 434 202 
<< m1 >>
rect 448 201 449 202 
<< m1 >>
rect 456 201 457 202 
<< m2 >>
rect 456 201 457 202 
<< m2c >>
rect 456 201 457 202 
<< m1 >>
rect 456 201 457 202 
<< m2 >>
rect 456 201 457 202 
<< m1 >>
rect 478 201 479 202 
<< m1 >>
rect 28 202 29 203 
<< m1 >>
rect 64 202 65 203 
<< m1 >>
rect 98 202 99 203 
<< m1 >>
rect 106 202 107 203 
<< m2 >>
rect 107 202 108 203 
<< m1 >>
rect 127 202 128 203 
<< m2 >>
rect 147 202 148 203 
<< m1 >>
rect 148 202 149 203 
<< m1 >>
rect 149 202 150 203 
<< m1 >>
rect 150 202 151 203 
<< m1 >>
rect 151 202 152 203 
<< m1 >>
rect 152 202 153 203 
<< m1 >>
rect 153 202 154 203 
<< m1 >>
rect 154 202 155 203 
<< m1 >>
rect 155 202 156 203 
<< m1 >>
rect 156 202 157 203 
<< m1 >>
rect 157 202 158 203 
<< m1 >>
rect 158 202 159 203 
<< m1 >>
rect 159 202 160 203 
<< m1 >>
rect 160 202 161 203 
<< m1 >>
rect 161 202 162 203 
<< m1 >>
rect 162 202 163 203 
<< m1 >>
rect 163 202 164 203 
<< m2 >>
rect 163 202 164 203 
<< m1 >>
rect 164 202 165 203 
<< m1 >>
rect 165 202 166 203 
<< m1 >>
rect 166 202 167 203 
<< m1 >>
rect 167 202 168 203 
<< m1 >>
rect 168 202 169 203 
<< m1 >>
rect 169 202 170 203 
<< m1 >>
rect 170 202 171 203 
<< m1 >>
rect 171 202 172 203 
<< m1 >>
rect 172 202 173 203 
<< m1 >>
rect 173 202 174 203 
<< m1 >>
rect 174 202 175 203 
<< m1 >>
rect 175 202 176 203 
<< m1 >>
rect 176 202 177 203 
<< m1 >>
rect 177 202 178 203 
<< m1 >>
rect 178 202 179 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m2c >>
rect 179 202 180 203 
<< m1 >>
rect 179 202 180 203 
<< m2 >>
rect 179 202 180 203 
<< m2 >>
rect 180 202 181 203 
<< m1 >>
rect 181 202 182 203 
<< m2 >>
rect 181 202 182 203 
<< m2 >>
rect 182 202 183 203 
<< m1 >>
rect 183 202 184 203 
<< m2 >>
rect 183 202 184 203 
<< m2c >>
rect 183 202 184 203 
<< m1 >>
rect 183 202 184 203 
<< m2 >>
rect 183 202 184 203 
<< m1 >>
rect 184 202 185 203 
<< m1 >>
rect 185 202 186 203 
<< m2 >>
rect 185 202 186 203 
<< m1 >>
rect 186 202 187 203 
<< m1 >>
rect 187 202 188 203 
<< m2 >>
rect 187 202 188 203 
<< m1 >>
rect 188 202 189 203 
<< m1 >>
rect 189 202 190 203 
<< m1 >>
rect 190 202 191 203 
<< m1 >>
rect 191 202 192 203 
<< m1 >>
rect 192 202 193 203 
<< m2 >>
rect 192 202 193 203 
<< m1 >>
rect 193 202 194 203 
<< m2 >>
rect 193 202 194 203 
<< m1 >>
rect 194 202 195 203 
<< m2 >>
rect 194 202 195 203 
<< m1 >>
rect 195 202 196 203 
<< m2 >>
rect 195 202 196 203 
<< m1 >>
rect 196 202 197 203 
<< m2 >>
rect 196 202 197 203 
<< m1 >>
rect 197 202 198 203 
<< m2 >>
rect 197 202 198 203 
<< m1 >>
rect 198 202 199 203 
<< m2 >>
rect 198 202 199 203 
<< m1 >>
rect 199 202 200 203 
<< m2 >>
rect 199 202 200 203 
<< m1 >>
rect 200 202 201 203 
<< m2 >>
rect 200 202 201 203 
<< m1 >>
rect 201 202 202 203 
<< m2 >>
rect 201 202 202 203 
<< m1 >>
rect 202 202 203 203 
<< m2 >>
rect 202 202 203 203 
<< m1 >>
rect 203 202 204 203 
<< m2 >>
rect 203 202 204 203 
<< m1 >>
rect 204 202 205 203 
<< m2 >>
rect 204 202 205 203 
<< m1 >>
rect 205 202 206 203 
<< m2 >>
rect 205 202 206 203 
<< m1 >>
rect 206 202 207 203 
<< m2 >>
rect 206 202 207 203 
<< m1 >>
rect 207 202 208 203 
<< m2 >>
rect 207 202 208 203 
<< m1 >>
rect 208 202 209 203 
<< m2 >>
rect 208 202 209 203 
<< m2 >>
rect 209 202 210 203 
<< m1 >>
rect 210 202 211 203 
<< m2 >>
rect 210 202 211 203 
<< m2c >>
rect 210 202 211 203 
<< m1 >>
rect 210 202 211 203 
<< m2 >>
rect 210 202 211 203 
<< m1 >>
rect 211 202 212 203 
<< m1 >>
rect 212 202 213 203 
<< m1 >>
rect 214 202 215 203 
<< m2 >>
rect 215 202 216 203 
<< m1 >>
rect 216 202 217 203 
<< m2 >>
rect 216 202 217 203 
<< m2c >>
rect 216 202 217 203 
<< m1 >>
rect 216 202 217 203 
<< m2 >>
rect 216 202 217 203 
<< m1 >>
rect 217 202 218 203 
<< m1 >>
rect 218 202 219 203 
<< m1 >>
rect 219 202 220 203 
<< m1 >>
rect 221 202 222 203 
<< m1 >>
rect 226 202 227 203 
<< m2 >>
rect 234 202 235 203 
<< m1 >>
rect 235 202 236 203 
<< m1 >>
rect 237 202 238 203 
<< m1 >>
rect 238 202 239 203 
<< m1 >>
rect 239 202 240 203 
<< m1 >>
rect 240 202 241 203 
<< m1 >>
rect 241 202 242 203 
<< m1 >>
rect 242 202 243 203 
<< m2 >>
rect 242 202 243 203 
<< m1 >>
rect 243 202 244 203 
<< m1 >>
rect 244 202 245 203 
<< m2 >>
rect 244 202 245 203 
<< m1 >>
rect 245 202 246 203 
<< m1 >>
rect 246 202 247 203 
<< m1 >>
rect 247 202 248 203 
<< m1 >>
rect 248 202 249 203 
<< m1 >>
rect 249 202 250 203 
<< m1 >>
rect 250 202 251 203 
<< m1 >>
rect 251 202 252 203 
<< m1 >>
rect 252 202 253 203 
<< m1 >>
rect 253 202 254 203 
<< m2 >>
rect 253 202 254 203 
<< m1 >>
rect 254 202 255 203 
<< m1 >>
rect 255 202 256 203 
<< m1 >>
rect 256 202 257 203 
<< m1 >>
rect 257 202 258 203 
<< m1 >>
rect 258 202 259 203 
<< m1 >>
rect 259 202 260 203 
<< m1 >>
rect 260 202 261 203 
<< m1 >>
rect 261 202 262 203 
<< m1 >>
rect 262 202 263 203 
<< m2 >>
rect 262 202 263 203 
<< m1 >>
rect 263 202 264 203 
<< m1 >>
rect 264 202 265 203 
<< m1 >>
rect 265 202 266 203 
<< m1 >>
rect 266 202 267 203 
<< m1 >>
rect 267 202 268 203 
<< m1 >>
rect 268 202 269 203 
<< m1 >>
rect 269 202 270 203 
<< m1 >>
rect 270 202 271 203 
<< m1 >>
rect 271 202 272 203 
<< m1 >>
rect 272 202 273 203 
<< m1 >>
rect 273 202 274 203 
<< m1 >>
rect 274 202 275 203 
<< m1 >>
rect 275 202 276 203 
<< m1 >>
rect 276 202 277 203 
<< m1 >>
rect 277 202 278 203 
<< m1 >>
rect 278 202 279 203 
<< m1 >>
rect 279 202 280 203 
<< m1 >>
rect 280 202 281 203 
<< m1 >>
rect 281 202 282 203 
<< m1 >>
rect 282 202 283 203 
<< m1 >>
rect 283 202 284 203 
<< m2 >>
rect 295 202 296 203 
<< m1 >>
rect 296 202 297 203 
<< m1 >>
rect 298 202 299 203 
<< m1 >>
rect 299 202 300 203 
<< m1 >>
rect 300 202 301 203 
<< m1 >>
rect 301 202 302 203 
<< m1 >>
rect 302 202 303 203 
<< m2 >>
rect 302 202 303 203 
<< m2c >>
rect 302 202 303 203 
<< m1 >>
rect 302 202 303 203 
<< m2 >>
rect 302 202 303 203 
<< m2 >>
rect 303 202 304 203 
<< m1 >>
rect 304 202 305 203 
<< m2 >>
rect 304 202 305 203 
<< m2 >>
rect 305 202 306 203 
<< m1 >>
rect 306 202 307 203 
<< m2 >>
rect 306 202 307 203 
<< m2c >>
rect 306 202 307 203 
<< m1 >>
rect 306 202 307 203 
<< m2 >>
rect 306 202 307 203 
<< m1 >>
rect 307 202 308 203 
<< m1 >>
rect 308 202 309 203 
<< m2 >>
rect 308 202 309 203 
<< m1 >>
rect 309 202 310 203 
<< m1 >>
rect 310 202 311 203 
<< m1 >>
rect 311 202 312 203 
<< m1 >>
rect 312 202 313 203 
<< m1 >>
rect 313 202 314 203 
<< m1 >>
rect 314 202 315 203 
<< m2 >>
rect 314 202 315 203 
<< m2c >>
rect 314 202 315 203 
<< m1 >>
rect 314 202 315 203 
<< m2 >>
rect 314 202 315 203 
<< m2 >>
rect 315 202 316 203 
<< m1 >>
rect 316 202 317 203 
<< m2 >>
rect 316 202 317 203 
<< m2 >>
rect 317 202 318 203 
<< m1 >>
rect 318 202 319 203 
<< m2 >>
rect 318 202 319 203 
<< m2c >>
rect 318 202 319 203 
<< m1 >>
rect 318 202 319 203 
<< m2 >>
rect 318 202 319 203 
<< m1 >>
rect 319 202 320 203 
<< m1 >>
rect 320 202 321 203 
<< m1 >>
rect 321 202 322 203 
<< m1 >>
rect 322 202 323 203 
<< m1 >>
rect 323 202 324 203 
<< m1 >>
rect 324 202 325 203 
<< m1 >>
rect 325 202 326 203 
<< m1 >>
rect 326 202 327 203 
<< m1 >>
rect 327 202 328 203 
<< m1 >>
rect 328 202 329 203 
<< m1 >>
rect 329 202 330 203 
<< m1 >>
rect 330 202 331 203 
<< m2 >>
rect 330 202 331 203 
<< m1 >>
rect 331 202 332 203 
<< m1 >>
rect 332 202 333 203 
<< m2 >>
rect 332 202 333 203 
<< m2c >>
rect 332 202 333 203 
<< m1 >>
rect 332 202 333 203 
<< m2 >>
rect 332 202 333 203 
<< m2 >>
rect 333 202 334 203 
<< m1 >>
rect 334 202 335 203 
<< m2 >>
rect 334 202 335 203 
<< m2 >>
rect 335 202 336 203 
<< m1 >>
rect 336 202 337 203 
<< m2 >>
rect 336 202 337 203 
<< m2c >>
rect 336 202 337 203 
<< m1 >>
rect 336 202 337 203 
<< m2 >>
rect 336 202 337 203 
<< m1 >>
rect 337 202 338 203 
<< m1 >>
rect 338 202 339 203 
<< m1 >>
rect 339 202 340 203 
<< m1 >>
rect 340 202 341 203 
<< m1 >>
rect 341 202 342 203 
<< m1 >>
rect 342 202 343 203 
<< m1 >>
rect 343 202 344 203 
<< m1 >>
rect 344 202 345 203 
<< m1 >>
rect 345 202 346 203 
<< m1 >>
rect 346 202 347 203 
<< m1 >>
rect 347 202 348 203 
<< m1 >>
rect 348 202 349 203 
<< m1 >>
rect 349 202 350 203 
<< m1 >>
rect 350 202 351 203 
<< m1 >>
rect 351 202 352 203 
<< m1 >>
rect 352 202 353 203 
<< m1 >>
rect 353 202 354 203 
<< m1 >>
rect 354 202 355 203 
<< m1 >>
rect 355 202 356 203 
<< m1 >>
rect 356 202 357 203 
<< m1 >>
rect 357 202 358 203 
<< m1 >>
rect 358 202 359 203 
<< m1 >>
rect 359 202 360 203 
<< m1 >>
rect 360 202 361 203 
<< m1 >>
rect 361 202 362 203 
<< m1 >>
rect 362 202 363 203 
<< m1 >>
rect 363 202 364 203 
<< m1 >>
rect 364 202 365 203 
<< m1 >>
rect 365 202 366 203 
<< m1 >>
rect 366 202 367 203 
<< m1 >>
rect 367 202 368 203 
<< m1 >>
rect 368 202 369 203 
<< m1 >>
rect 369 202 370 203 
<< m1 >>
rect 370 202 371 203 
<< m1 >>
rect 371 202 372 203 
<< m1 >>
rect 372 202 373 203 
<< m1 >>
rect 373 202 374 203 
<< m1 >>
rect 374 202 375 203 
<< m1 >>
rect 375 202 376 203 
<< m1 >>
rect 376 202 377 203 
<< m1 >>
rect 377 202 378 203 
<< m2 >>
rect 377 202 378 203 
<< m2c >>
rect 377 202 378 203 
<< m1 >>
rect 377 202 378 203 
<< m2 >>
rect 377 202 378 203 
<< m2 >>
rect 378 202 379 203 
<< m1 >>
rect 379 202 380 203 
<< m2 >>
rect 379 202 380 203 
<< m2 >>
rect 380 202 381 203 
<< m1 >>
rect 381 202 382 203 
<< m2 >>
rect 381 202 382 203 
<< m2c >>
rect 381 202 382 203 
<< m1 >>
rect 381 202 382 203 
<< m2 >>
rect 381 202 382 203 
<< m1 >>
rect 382 202 383 203 
<< m1 >>
rect 383 202 384 203 
<< m1 >>
rect 384 202 385 203 
<< m1 >>
rect 385 202 386 203 
<< m1 >>
rect 386 202 387 203 
<< m1 >>
rect 387 202 388 203 
<< m1 >>
rect 388 202 389 203 
<< m1 >>
rect 389 202 390 203 
<< m1 >>
rect 390 202 391 203 
<< m1 >>
rect 391 202 392 203 
<< m1 >>
rect 392 202 393 203 
<< m1 >>
rect 393 202 394 203 
<< m1 >>
rect 394 202 395 203 
<< m1 >>
rect 402 202 403 203 
<< m1 >>
rect 404 202 405 203 
<< m2 >>
rect 405 202 406 203 
<< m1 >>
rect 406 202 407 203 
<< m1 >>
rect 415 202 416 203 
<< m1 >>
rect 417 202 418 203 
<< m1 >>
rect 419 202 420 203 
<< m1 >>
rect 420 202 421 203 
<< m1 >>
rect 421 202 422 203 
<< m1 >>
rect 422 202 423 203 
<< m1 >>
rect 423 202 424 203 
<< m2 >>
rect 423 202 424 203 
<< m1 >>
rect 424 202 425 203 
<< m1 >>
rect 425 202 426 203 
<< m1 >>
rect 426 202 427 203 
<< m1 >>
rect 427 202 428 203 
<< m1 >>
rect 428 202 429 203 
<< m1 >>
rect 429 202 430 203 
<< m1 >>
rect 430 202 431 203 
<< m1 >>
rect 433 202 434 203 
<< m1 >>
rect 448 202 449 203 
<< m2 >>
rect 456 202 457 203 
<< m1 >>
rect 478 202 479 203 
<< m1 >>
rect 28 203 29 204 
<< m1 >>
rect 64 203 65 204 
<< m2 >>
rect 64 203 65 204 
<< m2c >>
rect 64 203 65 204 
<< m1 >>
rect 64 203 65 204 
<< m2 >>
rect 64 203 65 204 
<< m1 >>
rect 98 203 99 204 
<< m1 >>
rect 99 203 100 204 
<< m1 >>
rect 100 203 101 204 
<< m2 >>
rect 100 203 101 204 
<< m2c >>
rect 100 203 101 204 
<< m1 >>
rect 100 203 101 204 
<< m2 >>
rect 100 203 101 204 
<< m1 >>
rect 106 203 107 204 
<< m2 >>
rect 107 203 108 204 
<< m1 >>
rect 127 203 128 204 
<< m2 >>
rect 147 203 148 204 
<< m1 >>
rect 148 203 149 204 
<< m2 >>
rect 163 203 164 204 
<< m1 >>
rect 181 203 182 204 
<< m2 >>
rect 185 203 186 204 
<< m2 >>
rect 187 203 188 204 
<< m2 >>
rect 192 203 193 204 
<< m1 >>
rect 214 203 215 204 
<< m2 >>
rect 215 203 216 204 
<< m1 >>
rect 221 203 222 204 
<< m1 >>
rect 226 203 227 204 
<< m2 >>
rect 234 203 235 204 
<< m1 >>
rect 235 203 236 204 
<< m2 >>
rect 242 203 243 204 
<< m2 >>
rect 244 203 245 204 
<< m2 >>
rect 253 203 254 204 
<< m2 >>
rect 262 203 263 204 
<< m1 >>
rect 283 203 284 204 
<< m2 >>
rect 295 203 296 204 
<< m1 >>
rect 296 203 297 204 
<< m1 >>
rect 304 203 305 204 
<< m2 >>
rect 308 203 309 204 
<< m1 >>
rect 316 203 317 204 
<< m2 >>
rect 330 203 331 204 
<< m1 >>
rect 334 203 335 204 
<< m1 >>
rect 379 203 380 204 
<< m1 >>
rect 402 203 403 204 
<< m1 >>
rect 404 203 405 204 
<< m2 >>
rect 405 203 406 204 
<< m1 >>
rect 406 203 407 204 
<< m1 >>
rect 415 203 416 204 
<< m2 >>
rect 415 203 416 204 
<< m2c >>
rect 415 203 416 204 
<< m1 >>
rect 415 203 416 204 
<< m2 >>
rect 415 203 416 204 
<< m1 >>
rect 417 203 418 204 
<< m2 >>
rect 417 203 418 204 
<< m2c >>
rect 417 203 418 204 
<< m1 >>
rect 417 203 418 204 
<< m2 >>
rect 417 203 418 204 
<< m2 >>
rect 423 203 424 204 
<< m1 >>
rect 433 203 434 204 
<< m2 >>
rect 433 203 434 204 
<< m2c >>
rect 433 203 434 204 
<< m1 >>
rect 433 203 434 204 
<< m2 >>
rect 433 203 434 204 
<< m1 >>
rect 448 203 449 204 
<< m1 >>
rect 449 203 450 204 
<< m1 >>
rect 450 203 451 204 
<< m1 >>
rect 451 203 452 204 
<< m1 >>
rect 452 203 453 204 
<< m1 >>
rect 453 203 454 204 
<< m1 >>
rect 454 203 455 204 
<< m1 >>
rect 455 203 456 204 
<< m1 >>
rect 456 203 457 204 
<< m2 >>
rect 456 203 457 204 
<< m1 >>
rect 457 203 458 204 
<< m1 >>
rect 458 203 459 204 
<< m2 >>
rect 458 203 459 204 
<< m2c >>
rect 458 203 459 204 
<< m1 >>
rect 458 203 459 204 
<< m2 >>
rect 458 203 459 204 
<< m1 >>
rect 478 203 479 204 
<< m1 >>
rect 28 204 29 205 
<< m2 >>
rect 64 204 65 205 
<< m2 >>
rect 100 204 101 205 
<< m2 >>
rect 102 204 103 205 
<< m2 >>
rect 103 204 104 205 
<< m2 >>
rect 104 204 105 205 
<< m2 >>
rect 105 204 106 205 
<< m1 >>
rect 106 204 107 205 
<< m2 >>
rect 106 204 107 205 
<< m2 >>
rect 107 204 108 205 
<< m1 >>
rect 127 204 128 205 
<< m2 >>
rect 147 204 148 205 
<< m1 >>
rect 148 204 149 205 
<< m2 >>
rect 148 204 149 205 
<< m2 >>
rect 149 204 150 205 
<< m1 >>
rect 150 204 151 205 
<< m2 >>
rect 150 204 151 205 
<< m2c >>
rect 150 204 151 205 
<< m1 >>
rect 150 204 151 205 
<< m2 >>
rect 150 204 151 205 
<< m1 >>
rect 163 204 164 205 
<< m2 >>
rect 163 204 164 205 
<< m2c >>
rect 163 204 164 205 
<< m1 >>
rect 163 204 164 205 
<< m2 >>
rect 163 204 164 205 
<< m1 >>
rect 181 204 182 205 
<< m1 >>
rect 185 204 186 205 
<< m2 >>
rect 185 204 186 205 
<< m2c >>
rect 185 204 186 205 
<< m1 >>
rect 185 204 186 205 
<< m2 >>
rect 185 204 186 205 
<< m1 >>
rect 187 204 188 205 
<< m2 >>
rect 187 204 188 205 
<< m2c >>
rect 187 204 188 205 
<< m1 >>
rect 187 204 188 205 
<< m2 >>
rect 187 204 188 205 
<< m1 >>
rect 188 204 189 205 
<< m1 >>
rect 189 204 190 205 
<< m1 >>
rect 190 204 191 205 
<< m1 >>
rect 191 204 192 205 
<< m1 >>
rect 192 204 193 205 
<< m2 >>
rect 192 204 193 205 
<< m1 >>
rect 193 204 194 205 
<< m1 >>
rect 205 204 206 205 
<< m2 >>
rect 205 204 206 205 
<< m2c >>
rect 205 204 206 205 
<< m1 >>
rect 205 204 206 205 
<< m2 >>
rect 205 204 206 205 
<< m2 >>
rect 206 204 207 205 
<< m1 >>
rect 207 204 208 205 
<< m2 >>
rect 207 204 208 205 
<< m1 >>
rect 208 204 209 205 
<< m2 >>
rect 208 204 209 205 
<< m1 >>
rect 209 204 210 205 
<< m2 >>
rect 209 204 210 205 
<< m1 >>
rect 210 204 211 205 
<< m2 >>
rect 210 204 211 205 
<< m1 >>
rect 211 204 212 205 
<< m2 >>
rect 211 204 212 205 
<< m1 >>
rect 212 204 213 205 
<< m2 >>
rect 212 204 213 205 
<< m1 >>
rect 213 204 214 205 
<< m2 >>
rect 213 204 214 205 
<< m1 >>
rect 214 204 215 205 
<< m2 >>
rect 214 204 215 205 
<< m2 >>
rect 215 204 216 205 
<< m1 >>
rect 221 204 222 205 
<< m2 >>
rect 221 204 222 205 
<< m2c >>
rect 221 204 222 205 
<< m1 >>
rect 221 204 222 205 
<< m2 >>
rect 221 204 222 205 
<< m1 >>
rect 226 204 227 205 
<< m2 >>
rect 234 204 235 205 
<< m1 >>
rect 235 204 236 205 
<< m1 >>
rect 242 204 243 205 
<< m2 >>
rect 242 204 243 205 
<< m2c >>
rect 242 204 243 205 
<< m1 >>
rect 242 204 243 205 
<< m2 >>
rect 242 204 243 205 
<< m1 >>
rect 244 204 245 205 
<< m2 >>
rect 244 204 245 205 
<< m2c >>
rect 244 204 245 205 
<< m1 >>
rect 244 204 245 205 
<< m2 >>
rect 244 204 245 205 
<< m1 >>
rect 253 204 254 205 
<< m2 >>
rect 253 204 254 205 
<< m2c >>
rect 253 204 254 205 
<< m1 >>
rect 253 204 254 205 
<< m2 >>
rect 253 204 254 205 
<< m1 >>
rect 262 204 263 205 
<< m2 >>
rect 262 204 263 205 
<< m2c >>
rect 262 204 263 205 
<< m1 >>
rect 262 204 263 205 
<< m2 >>
rect 262 204 263 205 
<< m1 >>
rect 283 204 284 205 
<< m2 >>
rect 295 204 296 205 
<< m1 >>
rect 296 204 297 205 
<< m2 >>
rect 296 204 297 205 
<< m2 >>
rect 297 204 298 205 
<< m2 >>
rect 298 204 299 205 
<< m2 >>
rect 299 204 300 205 
<< m2 >>
rect 300 204 301 205 
<< m2 >>
rect 301 204 302 205 
<< m2 >>
rect 302 204 303 205 
<< m2 >>
rect 303 204 304 205 
<< m1 >>
rect 304 204 305 205 
<< m2 >>
rect 304 204 305 205 
<< m2 >>
rect 305 204 306 205 
<< m1 >>
rect 306 204 307 205 
<< m2 >>
rect 306 204 307 205 
<< m2c >>
rect 306 204 307 205 
<< m1 >>
rect 306 204 307 205 
<< m2 >>
rect 306 204 307 205 
<< m1 >>
rect 307 204 308 205 
<< m1 >>
rect 308 204 309 205 
<< m2 >>
rect 308 204 309 205 
<< m2c >>
rect 308 204 309 205 
<< m1 >>
rect 308 204 309 205 
<< m2 >>
rect 308 204 309 205 
<< m1 >>
rect 316 204 317 205 
<< m1 >>
rect 330 204 331 205 
<< m2 >>
rect 330 204 331 205 
<< m2c >>
rect 330 204 331 205 
<< m1 >>
rect 330 204 331 205 
<< m2 >>
rect 330 204 331 205 
<< m1 >>
rect 334 204 335 205 
<< m1 >>
rect 379 204 380 205 
<< m1 >>
rect 402 204 403 205 
<< m1 >>
rect 404 204 405 205 
<< m2 >>
rect 405 204 406 205 
<< m1 >>
rect 406 204 407 205 
<< m2 >>
rect 406 204 407 205 
<< m2 >>
rect 407 204 408 205 
<< m2 >>
rect 408 204 409 205 
<< m2 >>
rect 409 204 410 205 
<< m2 >>
rect 410 204 411 205 
<< m2 >>
rect 415 204 416 205 
<< m2 >>
rect 417 204 418 205 
<< m2 >>
rect 418 204 419 205 
<< m2 >>
rect 419 204 420 205 
<< m2 >>
rect 420 204 421 205 
<< m2 >>
rect 423 204 424 205 
<< m2 >>
rect 433 204 434 205 
<< m2 >>
rect 456 204 457 205 
<< m2 >>
rect 458 204 459 205 
<< m2 >>
rect 460 204 461 205 
<< m2 >>
rect 461 204 462 205 
<< m1 >>
rect 462 204 463 205 
<< m2 >>
rect 462 204 463 205 
<< m2c >>
rect 462 204 463 205 
<< m1 >>
rect 462 204 463 205 
<< m2 >>
rect 462 204 463 205 
<< m1 >>
rect 463 204 464 205 
<< m1 >>
rect 464 204 465 205 
<< m1 >>
rect 465 204 466 205 
<< m1 >>
rect 466 204 467 205 
<< m1 >>
rect 467 204 468 205 
<< m1 >>
rect 468 204 469 205 
<< m1 >>
rect 469 204 470 205 
<< m1 >>
rect 470 204 471 205 
<< m1 >>
rect 471 204 472 205 
<< m1 >>
rect 472 204 473 205 
<< m1 >>
rect 473 204 474 205 
<< m1 >>
rect 474 204 475 205 
<< m1 >>
rect 475 204 476 205 
<< m1 >>
rect 476 204 477 205 
<< m1 >>
rect 477 204 478 205 
<< m1 >>
rect 478 204 479 205 
<< m1 >>
rect 28 205 29 206 
<< m1 >>
rect 30 205 31 206 
<< m1 >>
rect 31 205 32 206 
<< m1 >>
rect 32 205 33 206 
<< m1 >>
rect 33 205 34 206 
<< m1 >>
rect 34 205 35 206 
<< m1 >>
rect 35 205 36 206 
<< m1 >>
rect 36 205 37 206 
<< m1 >>
rect 37 205 38 206 
<< m1 >>
rect 38 205 39 206 
<< m1 >>
rect 39 205 40 206 
<< m1 >>
rect 40 205 41 206 
<< m1 >>
rect 41 205 42 206 
<< m1 >>
rect 42 205 43 206 
<< m1 >>
rect 43 205 44 206 
<< m1 >>
rect 44 205 45 206 
<< m1 >>
rect 45 205 46 206 
<< m1 >>
rect 46 205 47 206 
<< m1 >>
rect 47 205 48 206 
<< m1 >>
rect 48 205 49 206 
<< m1 >>
rect 49 205 50 206 
<< m1 >>
rect 50 205 51 206 
<< m1 >>
rect 51 205 52 206 
<< m1 >>
rect 52 205 53 206 
<< m1 >>
rect 53 205 54 206 
<< m1 >>
rect 54 205 55 206 
<< m1 >>
rect 55 205 56 206 
<< m1 >>
rect 56 205 57 206 
<< m1 >>
rect 57 205 58 206 
<< m1 >>
rect 58 205 59 206 
<< m1 >>
rect 59 205 60 206 
<< m1 >>
rect 60 205 61 206 
<< m1 >>
rect 61 205 62 206 
<< m1 >>
rect 62 205 63 206 
<< m1 >>
rect 63 205 64 206 
<< m1 >>
rect 64 205 65 206 
<< m2 >>
rect 64 205 65 206 
<< m1 >>
rect 65 205 66 206 
<< m1 >>
rect 66 205 67 206 
<< m1 >>
rect 67 205 68 206 
<< m1 >>
rect 68 205 69 206 
<< m1 >>
rect 69 205 70 206 
<< m1 >>
rect 70 205 71 206 
<< m1 >>
rect 71 205 72 206 
<< m1 >>
rect 72 205 73 206 
<< m1 >>
rect 73 205 74 206 
<< m1 >>
rect 74 205 75 206 
<< m1 >>
rect 75 205 76 206 
<< m1 >>
rect 76 205 77 206 
<< m1 >>
rect 77 205 78 206 
<< m1 >>
rect 78 205 79 206 
<< m1 >>
rect 79 205 80 206 
<< m1 >>
rect 80 205 81 206 
<< m1 >>
rect 81 205 82 206 
<< m1 >>
rect 82 205 83 206 
<< m1 >>
rect 83 205 84 206 
<< m1 >>
rect 84 205 85 206 
<< m1 >>
rect 85 205 86 206 
<< m1 >>
rect 86 205 87 206 
<< m1 >>
rect 87 205 88 206 
<< m1 >>
rect 88 205 89 206 
<< m1 >>
rect 89 205 90 206 
<< m1 >>
rect 90 205 91 206 
<< m1 >>
rect 91 205 92 206 
<< m1 >>
rect 92 205 93 206 
<< m1 >>
rect 93 205 94 206 
<< m1 >>
rect 94 205 95 206 
<< m1 >>
rect 95 205 96 206 
<< m1 >>
rect 96 205 97 206 
<< m1 >>
rect 97 205 98 206 
<< m1 >>
rect 98 205 99 206 
<< m1 >>
rect 99 205 100 206 
<< m1 >>
rect 100 205 101 206 
<< m2 >>
rect 100 205 101 206 
<< m1 >>
rect 101 205 102 206 
<< m1 >>
rect 102 205 103 206 
<< m2 >>
rect 102 205 103 206 
<< m1 >>
rect 103 205 104 206 
<< m1 >>
rect 104 205 105 206 
<< m1 >>
rect 105 205 106 206 
<< m1 >>
rect 106 205 107 206 
<< m1 >>
rect 127 205 128 206 
<< m1 >>
rect 148 205 149 206 
<< m1 >>
rect 150 205 151 206 
<< m1 >>
rect 163 205 164 206 
<< m1 >>
rect 181 205 182 206 
<< m1 >>
rect 185 205 186 206 
<< m2 >>
rect 192 205 193 206 
<< m1 >>
rect 193 205 194 206 
<< m1 >>
rect 205 205 206 206 
<< m1 >>
rect 207 205 208 206 
<< m2 >>
rect 221 205 222 206 
<< m2 >>
rect 225 205 226 206 
<< m1 >>
rect 226 205 227 206 
<< m2 >>
rect 226 205 227 206 
<< m2 >>
rect 227 205 228 206 
<< m1 >>
rect 228 205 229 206 
<< m2 >>
rect 228 205 229 206 
<< m1 >>
rect 229 205 230 206 
<< m2 >>
rect 229 205 230 206 
<< m1 >>
rect 230 205 231 206 
<< m2 >>
rect 230 205 231 206 
<< m1 >>
rect 231 205 232 206 
<< m1 >>
rect 232 205 233 206 
<< m1 >>
rect 233 205 234 206 
<< m2 >>
rect 233 205 234 206 
<< m2c >>
rect 233 205 234 206 
<< m1 >>
rect 233 205 234 206 
<< m2 >>
rect 233 205 234 206 
<< m2 >>
rect 234 205 235 206 
<< m1 >>
rect 235 205 236 206 
<< m1 >>
rect 242 205 243 206 
<< m1 >>
rect 244 205 245 206 
<< m1 >>
rect 246 205 247 206 
<< m1 >>
rect 247 205 248 206 
<< m1 >>
rect 248 205 249 206 
<< m1 >>
rect 249 205 250 206 
<< m1 >>
rect 250 205 251 206 
<< m1 >>
rect 253 205 254 206 
<< m1 >>
rect 262 205 263 206 
<< m1 >>
rect 283 205 284 206 
<< m1 >>
rect 296 205 297 206 
<< m1 >>
rect 298 205 299 206 
<< m1 >>
rect 299 205 300 206 
<< m1 >>
rect 300 205 301 206 
<< m1 >>
rect 301 205 302 206 
<< m1 >>
rect 302 205 303 206 
<< m1 >>
rect 303 205 304 206 
<< m1 >>
rect 304 205 305 206 
<< m1 >>
rect 316 205 317 206 
<< m1 >>
rect 330 205 331 206 
<< m1 >>
rect 334 205 335 206 
<< m1 >>
rect 379 205 380 206 
<< m1 >>
rect 402 205 403 206 
<< m1 >>
rect 404 205 405 206 
<< m1 >>
rect 406 205 407 206 
<< m1 >>
rect 407 205 408 206 
<< m1 >>
rect 408 205 409 206 
<< m1 >>
rect 409 205 410 206 
<< m1 >>
rect 410 205 411 206 
<< m2 >>
rect 410 205 411 206 
<< m1 >>
rect 411 205 412 206 
<< m1 >>
rect 412 205 413 206 
<< m1 >>
rect 413 205 414 206 
<< m1 >>
rect 414 205 415 206 
<< m1 >>
rect 415 205 416 206 
<< m2 >>
rect 415 205 416 206 
<< m1 >>
rect 416 205 417 206 
<< m1 >>
rect 417 205 418 206 
<< m1 >>
rect 418 205 419 206 
<< m1 >>
rect 419 205 420 206 
<< m1 >>
rect 420 205 421 206 
<< m2 >>
rect 420 205 421 206 
<< m1 >>
rect 421 205 422 206 
<< m1 >>
rect 422 205 423 206 
<< m1 >>
rect 423 205 424 206 
<< m2 >>
rect 423 205 424 206 
<< m1 >>
rect 424 205 425 206 
<< m1 >>
rect 425 205 426 206 
<< m1 >>
rect 426 205 427 206 
<< m1 >>
rect 427 205 428 206 
<< m1 >>
rect 428 205 429 206 
<< m1 >>
rect 429 205 430 206 
<< m1 >>
rect 430 205 431 206 
<< m1 >>
rect 431 205 432 206 
<< m1 >>
rect 432 205 433 206 
<< m1 >>
rect 433 205 434 206 
<< m2 >>
rect 433 205 434 206 
<< m1 >>
rect 434 205 435 206 
<< m1 >>
rect 435 205 436 206 
<< m1 >>
rect 436 205 437 206 
<< m1 >>
rect 437 205 438 206 
<< m1 >>
rect 438 205 439 206 
<< m1 >>
rect 439 205 440 206 
<< m1 >>
rect 440 205 441 206 
<< m1 >>
rect 441 205 442 206 
<< m1 >>
rect 442 205 443 206 
<< m1 >>
rect 443 205 444 206 
<< m1 >>
rect 444 205 445 206 
<< m1 >>
rect 445 205 446 206 
<< m1 >>
rect 446 205 447 206 
<< m1 >>
rect 447 205 448 206 
<< m1 >>
rect 448 205 449 206 
<< m1 >>
rect 449 205 450 206 
<< m1 >>
rect 450 205 451 206 
<< m1 >>
rect 451 205 452 206 
<< m1 >>
rect 452 205 453 206 
<< m1 >>
rect 453 205 454 206 
<< m1 >>
rect 454 205 455 206 
<< m1 >>
rect 455 205 456 206 
<< m1 >>
rect 456 205 457 206 
<< m2 >>
rect 456 205 457 206 
<< m1 >>
rect 457 205 458 206 
<< m1 >>
rect 458 205 459 206 
<< m2 >>
rect 458 205 459 206 
<< m1 >>
rect 459 205 460 206 
<< m1 >>
rect 460 205 461 206 
<< m2 >>
rect 460 205 461 206 
<< m1 >>
rect 28 206 29 207 
<< m1 >>
rect 30 206 31 207 
<< m2 >>
rect 64 206 65 207 
<< m2 >>
rect 100 206 101 207 
<< m2 >>
rect 102 206 103 207 
<< m1 >>
rect 127 206 128 207 
<< m1 >>
rect 148 206 149 207 
<< m1 >>
rect 150 206 151 207 
<< m1 >>
rect 163 206 164 207 
<< m2 >>
rect 163 206 164 207 
<< m2c >>
rect 163 206 164 207 
<< m1 >>
rect 163 206 164 207 
<< m2 >>
rect 163 206 164 207 
<< m1 >>
rect 181 206 182 207 
<< m1 >>
rect 185 206 186 207 
<< m1 >>
rect 190 206 191 207 
<< m1 >>
rect 191 206 192 207 
<< m2 >>
rect 191 206 192 207 
<< m2c >>
rect 191 206 192 207 
<< m1 >>
rect 191 206 192 207 
<< m2 >>
rect 191 206 192 207 
<< m2 >>
rect 192 206 193 207 
<< m1 >>
rect 193 206 194 207 
<< m1 >>
rect 205 206 206 207 
<< m1 >>
rect 207 206 208 207 
<< m1 >>
rect 217 206 218 207 
<< m1 >>
rect 218 206 219 207 
<< m1 >>
rect 219 206 220 207 
<< m1 >>
rect 220 206 221 207 
<< m1 >>
rect 221 206 222 207 
<< m2 >>
rect 221 206 222 207 
<< m1 >>
rect 222 206 223 207 
<< m1 >>
rect 223 206 224 207 
<< m1 >>
rect 224 206 225 207 
<< m2 >>
rect 224 206 225 207 
<< m2c >>
rect 224 206 225 207 
<< m1 >>
rect 224 206 225 207 
<< m2 >>
rect 224 206 225 207 
<< m2 >>
rect 225 206 226 207 
<< m1 >>
rect 226 206 227 207 
<< m1 >>
rect 228 206 229 207 
<< m2 >>
rect 230 206 231 207 
<< m1 >>
rect 235 206 236 207 
<< m1 >>
rect 242 206 243 207 
<< m2 >>
rect 242 206 243 207 
<< m2c >>
rect 242 206 243 207 
<< m1 >>
rect 242 206 243 207 
<< m2 >>
rect 242 206 243 207 
<< m2 >>
rect 243 206 244 207 
<< m1 >>
rect 244 206 245 207 
<< m2 >>
rect 244 206 245 207 
<< m2 >>
rect 245 206 246 207 
<< m1 >>
rect 246 206 247 207 
<< m2 >>
rect 246 206 247 207 
<< m2c >>
rect 246 206 247 207 
<< m1 >>
rect 246 206 247 207 
<< m2 >>
rect 246 206 247 207 
<< m1 >>
rect 250 206 251 207 
<< m1 >>
rect 253 206 254 207 
<< m2 >>
rect 254 206 255 207 
<< m1 >>
rect 255 206 256 207 
<< m2 >>
rect 255 206 256 207 
<< m2c >>
rect 255 206 256 207 
<< m1 >>
rect 255 206 256 207 
<< m2 >>
rect 255 206 256 207 
<< m1 >>
rect 256 206 257 207 
<< m1 >>
rect 257 206 258 207 
<< m1 >>
rect 258 206 259 207 
<< m1 >>
rect 259 206 260 207 
<< m1 >>
rect 260 206 261 207 
<< m1 >>
rect 261 206 262 207 
<< m1 >>
rect 262 206 263 207 
<< m1 >>
rect 283 206 284 207 
<< m1 >>
rect 296 206 297 207 
<< m1 >>
rect 298 206 299 207 
<< m1 >>
rect 316 206 317 207 
<< m1 >>
rect 330 206 331 207 
<< m1 >>
rect 334 206 335 207 
<< m1 >>
rect 379 206 380 207 
<< m1 >>
rect 402 206 403 207 
<< m1 >>
rect 404 206 405 207 
<< m2 >>
rect 410 206 411 207 
<< m2 >>
rect 415 206 416 207 
<< m2 >>
rect 420 206 421 207 
<< m2 >>
rect 423 206 424 207 
<< m2 >>
rect 433 206 434 207 
<< m2 >>
rect 456 206 457 207 
<< m2 >>
rect 458 206 459 207 
<< m1 >>
rect 460 206 461 207 
<< m2 >>
rect 460 206 461 207 
<< m1 >>
rect 28 207 29 208 
<< m1 >>
rect 30 207 31 208 
<< m1 >>
rect 64 207 65 208 
<< m2 >>
rect 64 207 65 208 
<< m2c >>
rect 64 207 65 208 
<< m1 >>
rect 64 207 65 208 
<< m2 >>
rect 64 207 65 208 
<< m1 >>
rect 100 207 101 208 
<< m2 >>
rect 100 207 101 208 
<< m1 >>
rect 101 207 102 208 
<< m1 >>
rect 102 207 103 208 
<< m2 >>
rect 102 207 103 208 
<< m2c >>
rect 102 207 103 208 
<< m1 >>
rect 102 207 103 208 
<< m2 >>
rect 102 207 103 208 
<< m1 >>
rect 127 207 128 208 
<< m1 >>
rect 148 207 149 208 
<< m1 >>
rect 150 207 151 208 
<< m2 >>
rect 163 207 164 208 
<< m1 >>
rect 181 207 182 208 
<< m1 >>
rect 185 207 186 208 
<< m1 >>
rect 190 207 191 208 
<< m1 >>
rect 193 207 194 208 
<< m1 >>
rect 205 207 206 208 
<< m1 >>
rect 207 207 208 208 
<< m1 >>
rect 217 207 218 208 
<< m2 >>
rect 221 207 222 208 
<< m1 >>
rect 226 207 227 208 
<< m1 >>
rect 228 207 229 208 
<< m1 >>
rect 230 207 231 208 
<< m2 >>
rect 230 207 231 208 
<< m2c >>
rect 230 207 231 208 
<< m1 >>
rect 230 207 231 208 
<< m2 >>
rect 230 207 231 208 
<< m1 >>
rect 231 207 232 208 
<< m1 >>
rect 232 207 233 208 
<< m1 >>
rect 233 207 234 208 
<< m2 >>
rect 233 207 234 208 
<< m2c >>
rect 233 207 234 208 
<< m1 >>
rect 233 207 234 208 
<< m2 >>
rect 233 207 234 208 
<< m2 >>
rect 234 207 235 208 
<< m1 >>
rect 235 207 236 208 
<< m2 >>
rect 235 207 236 208 
<< m2 >>
rect 236 207 237 208 
<< m1 >>
rect 237 207 238 208 
<< m2 >>
rect 237 207 238 208 
<< m2c >>
rect 237 207 238 208 
<< m1 >>
rect 237 207 238 208 
<< m2 >>
rect 237 207 238 208 
<< m1 >>
rect 244 207 245 208 
<< m1 >>
rect 248 207 249 208 
<< m2 >>
rect 248 207 249 208 
<< m2c >>
rect 248 207 249 208 
<< m1 >>
rect 248 207 249 208 
<< m2 >>
rect 248 207 249 208 
<< m2 >>
rect 249 207 250 208 
<< m1 >>
rect 250 207 251 208 
<< m2 >>
rect 250 207 251 208 
<< m2 >>
rect 251 207 252 208 
<< m2 >>
rect 252 207 253 208 
<< m1 >>
rect 253 207 254 208 
<< m2 >>
rect 253 207 254 208 
<< m2 >>
rect 254 207 255 208 
<< m1 >>
rect 283 207 284 208 
<< m1 >>
rect 296 207 297 208 
<< m1 >>
rect 298 207 299 208 
<< m1 >>
rect 316 207 317 208 
<< m1 >>
rect 330 207 331 208 
<< m1 >>
rect 334 207 335 208 
<< m1 >>
rect 379 207 380 208 
<< m1 >>
rect 402 207 403 208 
<< m1 >>
rect 404 207 405 208 
<< m1 >>
rect 410 207 411 208 
<< m2 >>
rect 410 207 411 208 
<< m2c >>
rect 410 207 411 208 
<< m1 >>
rect 410 207 411 208 
<< m2 >>
rect 410 207 411 208 
<< m1 >>
rect 411 207 412 208 
<< m1 >>
rect 412 207 413 208 
<< m1 >>
rect 413 207 414 208 
<< m1 >>
rect 414 207 415 208 
<< m1 >>
rect 415 207 416 208 
<< m2 >>
rect 415 207 416 208 
<< m1 >>
rect 416 207 417 208 
<< m2 >>
rect 416 207 417 208 
<< m2 >>
rect 417 207 418 208 
<< m1 >>
rect 418 207 419 208 
<< m2 >>
rect 418 207 419 208 
<< m2c >>
rect 418 207 419 208 
<< m1 >>
rect 418 207 419 208 
<< m2 >>
rect 418 207 419 208 
<< m1 >>
rect 420 207 421 208 
<< m2 >>
rect 420 207 421 208 
<< m2c >>
rect 420 207 421 208 
<< m1 >>
rect 420 207 421 208 
<< m2 >>
rect 420 207 421 208 
<< m1 >>
rect 423 207 424 208 
<< m2 >>
rect 423 207 424 208 
<< m2c >>
rect 423 207 424 208 
<< m1 >>
rect 423 207 424 208 
<< m2 >>
rect 423 207 424 208 
<< m1 >>
rect 433 207 434 208 
<< m2 >>
rect 433 207 434 208 
<< m2c >>
rect 433 207 434 208 
<< m1 >>
rect 433 207 434 208 
<< m2 >>
rect 433 207 434 208 
<< m1 >>
rect 456 207 457 208 
<< m2 >>
rect 456 207 457 208 
<< m2c >>
rect 456 207 457 208 
<< m1 >>
rect 456 207 457 208 
<< m2 >>
rect 456 207 457 208 
<< m1 >>
rect 458 207 459 208 
<< m2 >>
rect 458 207 459 208 
<< m2c >>
rect 458 207 459 208 
<< m1 >>
rect 458 207 459 208 
<< m2 >>
rect 458 207 459 208 
<< m1 >>
rect 460 207 461 208 
<< m2 >>
rect 460 207 461 208 
<< m2 >>
rect 27 208 28 209 
<< m1 >>
rect 28 208 29 209 
<< m2 >>
rect 28 208 29 209 
<< m2 >>
rect 29 208 30 209 
<< m1 >>
rect 30 208 31 209 
<< m2 >>
rect 30 208 31 209 
<< m2c >>
rect 30 208 31 209 
<< m1 >>
rect 30 208 31 209 
<< m2 >>
rect 30 208 31 209 
<< m1 >>
rect 64 208 65 209 
<< m1 >>
rect 73 208 74 209 
<< m1 >>
rect 74 208 75 209 
<< m1 >>
rect 75 208 76 209 
<< m1 >>
rect 76 208 77 209 
<< m1 >>
rect 77 208 78 209 
<< m1 >>
rect 78 208 79 209 
<< m1 >>
rect 79 208 80 209 
<< m1 >>
rect 80 208 81 209 
<< m1 >>
rect 81 208 82 209 
<< m1 >>
rect 82 208 83 209 
<< m1 >>
rect 83 208 84 209 
<< m1 >>
rect 84 208 85 209 
<< m1 >>
rect 85 208 86 209 
<< m1 >>
rect 100 208 101 209 
<< m2 >>
rect 100 208 101 209 
<< m1 >>
rect 127 208 128 209 
<< m1 >>
rect 142 208 143 209 
<< m1 >>
rect 143 208 144 209 
<< m1 >>
rect 144 208 145 209 
<< m1 >>
rect 145 208 146 209 
<< m1 >>
rect 148 208 149 209 
<< m1 >>
rect 150 208 151 209 
<< m1 >>
rect 160 208 161 209 
<< m1 >>
rect 161 208 162 209 
<< m1 >>
rect 162 208 163 209 
<< m1 >>
rect 163 208 164 209 
<< m2 >>
rect 163 208 164 209 
<< m1 >>
rect 164 208 165 209 
<< m1 >>
rect 165 208 166 209 
<< m1 >>
rect 166 208 167 209 
<< m1 >>
rect 167 208 168 209 
<< m1 >>
rect 168 208 169 209 
<< m1 >>
rect 169 208 170 209 
<< m1 >>
rect 170 208 171 209 
<< m1 >>
rect 171 208 172 209 
<< m1 >>
rect 172 208 173 209 
<< m1 >>
rect 181 208 182 209 
<< m1 >>
rect 185 208 186 209 
<< m1 >>
rect 190 208 191 209 
<< m1 >>
rect 193 208 194 209 
<< m1 >>
rect 205 208 206 209 
<< m1 >>
rect 207 208 208 209 
<< m1 >>
rect 217 208 218 209 
<< m1 >>
rect 221 208 222 209 
<< m2 >>
rect 221 208 222 209 
<< m2c >>
rect 221 208 222 209 
<< m1 >>
rect 221 208 222 209 
<< m2 >>
rect 221 208 222 209 
<< m2 >>
rect 225 208 226 209 
<< m1 >>
rect 226 208 227 209 
<< m2 >>
rect 226 208 227 209 
<< m2 >>
rect 227 208 228 209 
<< m1 >>
rect 228 208 229 209 
<< m2 >>
rect 228 208 229 209 
<< m2c >>
rect 228 208 229 209 
<< m1 >>
rect 228 208 229 209 
<< m2 >>
rect 228 208 229 209 
<< m1 >>
rect 235 208 236 209 
<< m1 >>
rect 237 208 238 209 
<< m1 >>
rect 238 208 239 209 
<< m1 >>
rect 239 208 240 209 
<< m1 >>
rect 240 208 241 209 
<< m1 >>
rect 241 208 242 209 
<< m1 >>
rect 242 208 243 209 
<< m2 >>
rect 242 208 243 209 
<< m2c >>
rect 242 208 243 209 
<< m1 >>
rect 242 208 243 209 
<< m2 >>
rect 242 208 243 209 
<< m2 >>
rect 243 208 244 209 
<< m1 >>
rect 244 208 245 209 
<< m1 >>
rect 247 208 248 209 
<< m1 >>
rect 248 208 249 209 
<< m1 >>
rect 250 208 251 209 
<< m1 >>
rect 253 208 254 209 
<< m1 >>
rect 283 208 284 209 
<< m1 >>
rect 296 208 297 209 
<< m1 >>
rect 298 208 299 209 
<< m1 >>
rect 316 208 317 209 
<< m1 >>
rect 330 208 331 209 
<< m1 >>
rect 334 208 335 209 
<< m1 >>
rect 340 208 341 209 
<< m1 >>
rect 341 208 342 209 
<< m1 >>
rect 342 208 343 209 
<< m1 >>
rect 343 208 344 209 
<< m1 >>
rect 358 208 359 209 
<< m1 >>
rect 359 208 360 209 
<< m1 >>
rect 360 208 361 209 
<< m1 >>
rect 361 208 362 209 
<< m1 >>
rect 379 208 380 209 
<< m1 >>
rect 402 208 403 209 
<< m1 >>
rect 404 208 405 209 
<< m1 >>
rect 416 208 417 209 
<< m1 >>
rect 418 208 419 209 
<< m1 >>
rect 420 208 421 209 
<< m1 >>
rect 423 208 424 209 
<< m1 >>
rect 433 208 434 209 
<< m1 >>
rect 456 208 457 209 
<< m1 >>
rect 458 208 459 209 
<< m1 >>
rect 460 208 461 209 
<< m2 >>
rect 460 208 461 209 
<< m1 >>
rect 520 208 521 209 
<< m1 >>
rect 521 208 522 209 
<< m1 >>
rect 522 208 523 209 
<< m1 >>
rect 523 208 524 209 
<< m2 >>
rect 27 209 28 210 
<< m1 >>
rect 28 209 29 210 
<< m1 >>
rect 64 209 65 210 
<< m1 >>
rect 73 209 74 210 
<< m1 >>
rect 85 209 86 210 
<< m1 >>
rect 100 209 101 210 
<< m2 >>
rect 100 209 101 210 
<< m1 >>
rect 127 209 128 210 
<< m1 >>
rect 142 209 143 210 
<< m1 >>
rect 145 209 146 210 
<< m1 >>
rect 148 209 149 210 
<< m1 >>
rect 150 209 151 210 
<< m1 >>
rect 160 209 161 210 
<< m2 >>
rect 163 209 164 210 
<< m1 >>
rect 172 209 173 210 
<< m1 >>
rect 181 209 182 210 
<< m1 >>
rect 185 209 186 210 
<< m1 >>
rect 190 209 191 210 
<< m1 >>
rect 193 209 194 210 
<< m1 >>
rect 205 209 206 210 
<< m1 >>
rect 207 209 208 210 
<< m1 >>
rect 217 209 218 210 
<< m1 >>
rect 221 209 222 210 
<< m2 >>
rect 225 209 226 210 
<< m1 >>
rect 226 209 227 210 
<< m1 >>
rect 235 209 236 210 
<< m2 >>
rect 243 209 244 210 
<< m1 >>
rect 244 209 245 210 
<< m1 >>
rect 247 209 248 210 
<< m1 >>
rect 250 209 251 210 
<< m1 >>
rect 253 209 254 210 
<< m1 >>
rect 283 209 284 210 
<< m1 >>
rect 296 209 297 210 
<< m1 >>
rect 298 209 299 210 
<< m1 >>
rect 316 209 317 210 
<< m1 >>
rect 330 209 331 210 
<< m1 >>
rect 334 209 335 210 
<< m1 >>
rect 340 209 341 210 
<< m1 >>
rect 343 209 344 210 
<< m1 >>
rect 358 209 359 210 
<< m1 >>
rect 361 209 362 210 
<< m1 >>
rect 379 209 380 210 
<< m1 >>
rect 402 209 403 210 
<< m1 >>
rect 404 209 405 210 
<< m1 >>
rect 416 209 417 210 
<< m1 >>
rect 418 209 419 210 
<< m1 >>
rect 420 209 421 210 
<< m1 >>
rect 423 209 424 210 
<< m1 >>
rect 433 209 434 210 
<< m1 >>
rect 456 209 457 210 
<< m1 >>
rect 458 209 459 210 
<< m1 >>
rect 460 209 461 210 
<< m2 >>
rect 460 209 461 210 
<< m1 >>
rect 520 209 521 210 
<< m1 >>
rect 523 209 524 210 
<< pdiffusion >>
rect 12 210 13 211 
<< pdiffusion >>
rect 13 210 14 211 
<< pdiffusion >>
rect 14 210 15 211 
<< pdiffusion >>
rect 15 210 16 211 
<< pdiffusion >>
rect 16 210 17 211 
<< pdiffusion >>
rect 17 210 18 211 
<< m2 >>
rect 27 210 28 211 
<< m1 >>
rect 28 210 29 211 
<< pdiffusion >>
rect 30 210 31 211 
<< pdiffusion >>
rect 31 210 32 211 
<< pdiffusion >>
rect 32 210 33 211 
<< pdiffusion >>
rect 33 210 34 211 
<< pdiffusion >>
rect 34 210 35 211 
<< pdiffusion >>
rect 35 210 36 211 
<< pdiffusion >>
rect 48 210 49 211 
<< pdiffusion >>
rect 49 210 50 211 
<< pdiffusion >>
rect 50 210 51 211 
<< pdiffusion >>
rect 51 210 52 211 
<< pdiffusion >>
rect 52 210 53 211 
<< pdiffusion >>
rect 53 210 54 211 
<< m1 >>
rect 64 210 65 211 
<< pdiffusion >>
rect 66 210 67 211 
<< pdiffusion >>
rect 67 210 68 211 
<< pdiffusion >>
rect 68 210 69 211 
<< pdiffusion >>
rect 69 210 70 211 
<< pdiffusion >>
rect 70 210 71 211 
<< pdiffusion >>
rect 71 210 72 211 
<< m1 >>
rect 73 210 74 211 
<< pdiffusion >>
rect 84 210 85 211 
<< m1 >>
rect 85 210 86 211 
<< pdiffusion >>
rect 85 210 86 211 
<< pdiffusion >>
rect 86 210 87 211 
<< pdiffusion >>
rect 87 210 88 211 
<< pdiffusion >>
rect 88 210 89 211 
<< pdiffusion >>
rect 89 210 90 211 
<< m1 >>
rect 100 210 101 211 
<< m2 >>
rect 100 210 101 211 
<< pdiffusion >>
rect 102 210 103 211 
<< pdiffusion >>
rect 103 210 104 211 
<< pdiffusion >>
rect 104 210 105 211 
<< pdiffusion >>
rect 105 210 106 211 
<< pdiffusion >>
rect 106 210 107 211 
<< pdiffusion >>
rect 107 210 108 211 
<< m1 >>
rect 127 210 128 211 
<< pdiffusion >>
rect 138 210 139 211 
<< pdiffusion >>
rect 139 210 140 211 
<< pdiffusion >>
rect 140 210 141 211 
<< pdiffusion >>
rect 141 210 142 211 
<< m1 >>
rect 142 210 143 211 
<< pdiffusion >>
rect 142 210 143 211 
<< pdiffusion >>
rect 143 210 144 211 
<< m1 >>
rect 145 210 146 211 
<< m1 >>
rect 148 210 149 211 
<< m1 >>
rect 150 210 151 211 
<< pdiffusion >>
rect 156 210 157 211 
<< pdiffusion >>
rect 157 210 158 211 
<< pdiffusion >>
rect 158 210 159 211 
<< pdiffusion >>
rect 159 210 160 211 
<< m1 >>
rect 160 210 161 211 
<< pdiffusion >>
rect 160 210 161 211 
<< pdiffusion >>
rect 161 210 162 211 
<< m1 >>
rect 163 210 164 211 
<< m2 >>
rect 163 210 164 211 
<< m2c >>
rect 163 210 164 211 
<< m1 >>
rect 163 210 164 211 
<< m2 >>
rect 163 210 164 211 
<< m1 >>
rect 172 210 173 211 
<< pdiffusion >>
rect 174 210 175 211 
<< pdiffusion >>
rect 175 210 176 211 
<< pdiffusion >>
rect 176 210 177 211 
<< pdiffusion >>
rect 177 210 178 211 
<< pdiffusion >>
rect 178 210 179 211 
<< pdiffusion >>
rect 179 210 180 211 
<< m1 >>
rect 181 210 182 211 
<< m1 >>
rect 185 210 186 211 
<< m1 >>
rect 190 210 191 211 
<< pdiffusion >>
rect 192 210 193 211 
<< m1 >>
rect 193 210 194 211 
<< pdiffusion >>
rect 193 210 194 211 
<< pdiffusion >>
rect 194 210 195 211 
<< pdiffusion >>
rect 195 210 196 211 
<< pdiffusion >>
rect 196 210 197 211 
<< pdiffusion >>
rect 197 210 198 211 
<< m1 >>
rect 205 210 206 211 
<< m1 >>
rect 207 210 208 211 
<< pdiffusion >>
rect 210 210 211 211 
<< pdiffusion >>
rect 211 210 212 211 
<< pdiffusion >>
rect 212 210 213 211 
<< pdiffusion >>
rect 213 210 214 211 
<< pdiffusion >>
rect 214 210 215 211 
<< pdiffusion >>
rect 215 210 216 211 
<< m1 >>
rect 217 210 218 211 
<< m1 >>
rect 221 210 222 211 
<< m2 >>
rect 225 210 226 211 
<< m1 >>
rect 226 210 227 211 
<< pdiffusion >>
rect 228 210 229 211 
<< pdiffusion >>
rect 229 210 230 211 
<< pdiffusion >>
rect 230 210 231 211 
<< pdiffusion >>
rect 231 210 232 211 
<< pdiffusion >>
rect 232 210 233 211 
<< pdiffusion >>
rect 233 210 234 211 
<< m1 >>
rect 235 210 236 211 
<< m2 >>
rect 243 210 244 211 
<< m1 >>
rect 244 210 245 211 
<< pdiffusion >>
rect 246 210 247 211 
<< m1 >>
rect 247 210 248 211 
<< pdiffusion >>
rect 247 210 248 211 
<< pdiffusion >>
rect 248 210 249 211 
<< pdiffusion >>
rect 249 210 250 211 
<< m1 >>
rect 250 210 251 211 
<< pdiffusion >>
rect 250 210 251 211 
<< pdiffusion >>
rect 251 210 252 211 
<< m1 >>
rect 253 210 254 211 
<< pdiffusion >>
rect 264 210 265 211 
<< pdiffusion >>
rect 265 210 266 211 
<< pdiffusion >>
rect 266 210 267 211 
<< pdiffusion >>
rect 267 210 268 211 
<< pdiffusion >>
rect 268 210 269 211 
<< pdiffusion >>
rect 269 210 270 211 
<< pdiffusion >>
rect 282 210 283 211 
<< m1 >>
rect 283 210 284 211 
<< pdiffusion >>
rect 283 210 284 211 
<< pdiffusion >>
rect 284 210 285 211 
<< pdiffusion >>
rect 285 210 286 211 
<< pdiffusion >>
rect 286 210 287 211 
<< pdiffusion >>
rect 287 210 288 211 
<< m1 >>
rect 296 210 297 211 
<< m1 >>
rect 298 210 299 211 
<< pdiffusion >>
rect 300 210 301 211 
<< pdiffusion >>
rect 301 210 302 211 
<< pdiffusion >>
rect 302 210 303 211 
<< pdiffusion >>
rect 303 210 304 211 
<< pdiffusion >>
rect 304 210 305 211 
<< pdiffusion >>
rect 305 210 306 211 
<< m1 >>
rect 316 210 317 211 
<< pdiffusion >>
rect 318 210 319 211 
<< pdiffusion >>
rect 319 210 320 211 
<< pdiffusion >>
rect 320 210 321 211 
<< pdiffusion >>
rect 321 210 322 211 
<< pdiffusion >>
rect 322 210 323 211 
<< pdiffusion >>
rect 323 210 324 211 
<< m1 >>
rect 330 210 331 211 
<< m1 >>
rect 334 210 335 211 
<< pdiffusion >>
rect 336 210 337 211 
<< pdiffusion >>
rect 337 210 338 211 
<< pdiffusion >>
rect 338 210 339 211 
<< pdiffusion >>
rect 339 210 340 211 
<< m1 >>
rect 340 210 341 211 
<< pdiffusion >>
rect 340 210 341 211 
<< pdiffusion >>
rect 341 210 342 211 
<< m1 >>
rect 343 210 344 211 
<< pdiffusion >>
rect 354 210 355 211 
<< pdiffusion >>
rect 355 210 356 211 
<< pdiffusion >>
rect 356 210 357 211 
<< pdiffusion >>
rect 357 210 358 211 
<< m1 >>
rect 358 210 359 211 
<< pdiffusion >>
rect 358 210 359 211 
<< pdiffusion >>
rect 359 210 360 211 
<< m1 >>
rect 361 210 362 211 
<< pdiffusion >>
rect 372 210 373 211 
<< pdiffusion >>
rect 373 210 374 211 
<< pdiffusion >>
rect 374 210 375 211 
<< pdiffusion >>
rect 375 210 376 211 
<< pdiffusion >>
rect 376 210 377 211 
<< pdiffusion >>
rect 377 210 378 211 
<< m1 >>
rect 379 210 380 211 
<< pdiffusion >>
rect 390 210 391 211 
<< pdiffusion >>
rect 391 210 392 211 
<< pdiffusion >>
rect 392 210 393 211 
<< pdiffusion >>
rect 393 210 394 211 
<< pdiffusion >>
rect 394 210 395 211 
<< pdiffusion >>
rect 395 210 396 211 
<< m1 >>
rect 402 210 403 211 
<< m1 >>
rect 404 210 405 211 
<< pdiffusion >>
rect 408 210 409 211 
<< pdiffusion >>
rect 409 210 410 211 
<< pdiffusion >>
rect 410 210 411 211 
<< pdiffusion >>
rect 411 210 412 211 
<< pdiffusion >>
rect 412 210 413 211 
<< pdiffusion >>
rect 413 210 414 211 
<< m1 >>
rect 416 210 417 211 
<< m1 >>
rect 418 210 419 211 
<< m1 >>
rect 420 210 421 211 
<< m1 >>
rect 423 210 424 211 
<< pdiffusion >>
rect 426 210 427 211 
<< pdiffusion >>
rect 427 210 428 211 
<< pdiffusion >>
rect 428 210 429 211 
<< pdiffusion >>
rect 429 210 430 211 
<< pdiffusion >>
rect 430 210 431 211 
<< pdiffusion >>
rect 431 210 432 211 
<< m1 >>
rect 433 210 434 211 
<< pdiffusion >>
rect 444 210 445 211 
<< pdiffusion >>
rect 445 210 446 211 
<< pdiffusion >>
rect 446 210 447 211 
<< pdiffusion >>
rect 447 210 448 211 
<< pdiffusion >>
rect 448 210 449 211 
<< pdiffusion >>
rect 449 210 450 211 
<< m1 >>
rect 456 210 457 211 
<< m1 >>
rect 458 210 459 211 
<< m1 >>
rect 460 210 461 211 
<< m2 >>
rect 460 210 461 211 
<< pdiffusion >>
rect 462 210 463 211 
<< pdiffusion >>
rect 463 210 464 211 
<< pdiffusion >>
rect 464 210 465 211 
<< pdiffusion >>
rect 465 210 466 211 
<< pdiffusion >>
rect 466 210 467 211 
<< pdiffusion >>
rect 467 210 468 211 
<< pdiffusion >>
rect 480 210 481 211 
<< pdiffusion >>
rect 481 210 482 211 
<< pdiffusion >>
rect 482 210 483 211 
<< pdiffusion >>
rect 483 210 484 211 
<< pdiffusion >>
rect 484 210 485 211 
<< pdiffusion >>
rect 485 210 486 211 
<< pdiffusion >>
rect 498 210 499 211 
<< pdiffusion >>
rect 499 210 500 211 
<< pdiffusion >>
rect 500 210 501 211 
<< pdiffusion >>
rect 501 210 502 211 
<< pdiffusion >>
rect 502 210 503 211 
<< pdiffusion >>
rect 503 210 504 211 
<< pdiffusion >>
rect 516 210 517 211 
<< pdiffusion >>
rect 517 210 518 211 
<< pdiffusion >>
rect 518 210 519 211 
<< pdiffusion >>
rect 519 210 520 211 
<< m1 >>
rect 520 210 521 211 
<< pdiffusion >>
rect 520 210 521 211 
<< pdiffusion >>
rect 521 210 522 211 
<< m1 >>
rect 523 210 524 211 
<< pdiffusion >>
rect 12 211 13 212 
<< pdiffusion >>
rect 13 211 14 212 
<< pdiffusion >>
rect 14 211 15 212 
<< pdiffusion >>
rect 15 211 16 212 
<< pdiffusion >>
rect 16 211 17 212 
<< pdiffusion >>
rect 17 211 18 212 
<< m2 >>
rect 27 211 28 212 
<< m1 >>
rect 28 211 29 212 
<< pdiffusion >>
rect 30 211 31 212 
<< pdiffusion >>
rect 31 211 32 212 
<< pdiffusion >>
rect 32 211 33 212 
<< pdiffusion >>
rect 33 211 34 212 
<< pdiffusion >>
rect 34 211 35 212 
<< pdiffusion >>
rect 35 211 36 212 
<< pdiffusion >>
rect 48 211 49 212 
<< pdiffusion >>
rect 49 211 50 212 
<< pdiffusion >>
rect 50 211 51 212 
<< pdiffusion >>
rect 51 211 52 212 
<< pdiffusion >>
rect 52 211 53 212 
<< pdiffusion >>
rect 53 211 54 212 
<< m1 >>
rect 64 211 65 212 
<< pdiffusion >>
rect 66 211 67 212 
<< pdiffusion >>
rect 67 211 68 212 
<< pdiffusion >>
rect 68 211 69 212 
<< pdiffusion >>
rect 69 211 70 212 
<< pdiffusion >>
rect 70 211 71 212 
<< pdiffusion >>
rect 71 211 72 212 
<< m1 >>
rect 73 211 74 212 
<< pdiffusion >>
rect 84 211 85 212 
<< pdiffusion >>
rect 85 211 86 212 
<< pdiffusion >>
rect 86 211 87 212 
<< pdiffusion >>
rect 87 211 88 212 
<< pdiffusion >>
rect 88 211 89 212 
<< pdiffusion >>
rect 89 211 90 212 
<< m1 >>
rect 100 211 101 212 
<< m2 >>
rect 100 211 101 212 
<< pdiffusion >>
rect 102 211 103 212 
<< pdiffusion >>
rect 103 211 104 212 
<< pdiffusion >>
rect 104 211 105 212 
<< pdiffusion >>
rect 105 211 106 212 
<< pdiffusion >>
rect 106 211 107 212 
<< pdiffusion >>
rect 107 211 108 212 
<< m1 >>
rect 127 211 128 212 
<< pdiffusion >>
rect 138 211 139 212 
<< pdiffusion >>
rect 139 211 140 212 
<< pdiffusion >>
rect 140 211 141 212 
<< pdiffusion >>
rect 141 211 142 212 
<< pdiffusion >>
rect 142 211 143 212 
<< pdiffusion >>
rect 143 211 144 212 
<< m1 >>
rect 145 211 146 212 
<< m1 >>
rect 148 211 149 212 
<< m1 >>
rect 150 211 151 212 
<< pdiffusion >>
rect 156 211 157 212 
<< pdiffusion >>
rect 157 211 158 212 
<< pdiffusion >>
rect 158 211 159 212 
<< pdiffusion >>
rect 159 211 160 212 
<< pdiffusion >>
rect 160 211 161 212 
<< pdiffusion >>
rect 161 211 162 212 
<< m1 >>
rect 163 211 164 212 
<< m1 >>
rect 172 211 173 212 
<< pdiffusion >>
rect 174 211 175 212 
<< pdiffusion >>
rect 175 211 176 212 
<< pdiffusion >>
rect 176 211 177 212 
<< pdiffusion >>
rect 177 211 178 212 
<< pdiffusion >>
rect 178 211 179 212 
<< pdiffusion >>
rect 179 211 180 212 
<< m1 >>
rect 181 211 182 212 
<< m1 >>
rect 185 211 186 212 
<< m1 >>
rect 190 211 191 212 
<< pdiffusion >>
rect 192 211 193 212 
<< pdiffusion >>
rect 193 211 194 212 
<< pdiffusion >>
rect 194 211 195 212 
<< pdiffusion >>
rect 195 211 196 212 
<< pdiffusion >>
rect 196 211 197 212 
<< pdiffusion >>
rect 197 211 198 212 
<< m1 >>
rect 205 211 206 212 
<< m1 >>
rect 207 211 208 212 
<< pdiffusion >>
rect 210 211 211 212 
<< pdiffusion >>
rect 211 211 212 212 
<< pdiffusion >>
rect 212 211 213 212 
<< pdiffusion >>
rect 213 211 214 212 
<< pdiffusion >>
rect 214 211 215 212 
<< pdiffusion >>
rect 215 211 216 212 
<< m1 >>
rect 217 211 218 212 
<< m1 >>
rect 221 211 222 212 
<< m2 >>
rect 225 211 226 212 
<< m1 >>
rect 226 211 227 212 
<< pdiffusion >>
rect 228 211 229 212 
<< pdiffusion >>
rect 229 211 230 212 
<< pdiffusion >>
rect 230 211 231 212 
<< pdiffusion >>
rect 231 211 232 212 
<< pdiffusion >>
rect 232 211 233 212 
<< pdiffusion >>
rect 233 211 234 212 
<< m1 >>
rect 235 211 236 212 
<< m2 >>
rect 243 211 244 212 
<< m1 >>
rect 244 211 245 212 
<< pdiffusion >>
rect 246 211 247 212 
<< pdiffusion >>
rect 247 211 248 212 
<< pdiffusion >>
rect 248 211 249 212 
<< pdiffusion >>
rect 249 211 250 212 
<< pdiffusion >>
rect 250 211 251 212 
<< pdiffusion >>
rect 251 211 252 212 
<< m1 >>
rect 253 211 254 212 
<< pdiffusion >>
rect 264 211 265 212 
<< pdiffusion >>
rect 265 211 266 212 
<< pdiffusion >>
rect 266 211 267 212 
<< pdiffusion >>
rect 267 211 268 212 
<< pdiffusion >>
rect 268 211 269 212 
<< pdiffusion >>
rect 269 211 270 212 
<< pdiffusion >>
rect 282 211 283 212 
<< pdiffusion >>
rect 283 211 284 212 
<< pdiffusion >>
rect 284 211 285 212 
<< pdiffusion >>
rect 285 211 286 212 
<< pdiffusion >>
rect 286 211 287 212 
<< pdiffusion >>
rect 287 211 288 212 
<< m1 >>
rect 296 211 297 212 
<< m1 >>
rect 298 211 299 212 
<< pdiffusion >>
rect 300 211 301 212 
<< pdiffusion >>
rect 301 211 302 212 
<< pdiffusion >>
rect 302 211 303 212 
<< pdiffusion >>
rect 303 211 304 212 
<< pdiffusion >>
rect 304 211 305 212 
<< pdiffusion >>
rect 305 211 306 212 
<< m1 >>
rect 316 211 317 212 
<< pdiffusion >>
rect 318 211 319 212 
<< pdiffusion >>
rect 319 211 320 212 
<< pdiffusion >>
rect 320 211 321 212 
<< pdiffusion >>
rect 321 211 322 212 
<< pdiffusion >>
rect 322 211 323 212 
<< pdiffusion >>
rect 323 211 324 212 
<< m1 >>
rect 330 211 331 212 
<< m1 >>
rect 334 211 335 212 
<< pdiffusion >>
rect 336 211 337 212 
<< pdiffusion >>
rect 337 211 338 212 
<< pdiffusion >>
rect 338 211 339 212 
<< pdiffusion >>
rect 339 211 340 212 
<< pdiffusion >>
rect 340 211 341 212 
<< pdiffusion >>
rect 341 211 342 212 
<< m1 >>
rect 343 211 344 212 
<< pdiffusion >>
rect 354 211 355 212 
<< pdiffusion >>
rect 355 211 356 212 
<< pdiffusion >>
rect 356 211 357 212 
<< pdiffusion >>
rect 357 211 358 212 
<< pdiffusion >>
rect 358 211 359 212 
<< pdiffusion >>
rect 359 211 360 212 
<< m1 >>
rect 361 211 362 212 
<< pdiffusion >>
rect 372 211 373 212 
<< pdiffusion >>
rect 373 211 374 212 
<< pdiffusion >>
rect 374 211 375 212 
<< pdiffusion >>
rect 375 211 376 212 
<< pdiffusion >>
rect 376 211 377 212 
<< pdiffusion >>
rect 377 211 378 212 
<< m1 >>
rect 379 211 380 212 
<< pdiffusion >>
rect 390 211 391 212 
<< pdiffusion >>
rect 391 211 392 212 
<< pdiffusion >>
rect 392 211 393 212 
<< pdiffusion >>
rect 393 211 394 212 
<< pdiffusion >>
rect 394 211 395 212 
<< pdiffusion >>
rect 395 211 396 212 
<< m1 >>
rect 402 211 403 212 
<< m1 >>
rect 404 211 405 212 
<< pdiffusion >>
rect 408 211 409 212 
<< pdiffusion >>
rect 409 211 410 212 
<< pdiffusion >>
rect 410 211 411 212 
<< pdiffusion >>
rect 411 211 412 212 
<< pdiffusion >>
rect 412 211 413 212 
<< pdiffusion >>
rect 413 211 414 212 
<< m1 >>
rect 416 211 417 212 
<< m1 >>
rect 418 211 419 212 
<< m1 >>
rect 420 211 421 212 
<< m1 >>
rect 423 211 424 212 
<< pdiffusion >>
rect 426 211 427 212 
<< pdiffusion >>
rect 427 211 428 212 
<< pdiffusion >>
rect 428 211 429 212 
<< pdiffusion >>
rect 429 211 430 212 
<< pdiffusion >>
rect 430 211 431 212 
<< pdiffusion >>
rect 431 211 432 212 
<< m1 >>
rect 433 211 434 212 
<< pdiffusion >>
rect 444 211 445 212 
<< pdiffusion >>
rect 445 211 446 212 
<< pdiffusion >>
rect 446 211 447 212 
<< pdiffusion >>
rect 447 211 448 212 
<< pdiffusion >>
rect 448 211 449 212 
<< pdiffusion >>
rect 449 211 450 212 
<< m1 >>
rect 456 211 457 212 
<< m1 >>
rect 458 211 459 212 
<< m1 >>
rect 460 211 461 212 
<< m2 >>
rect 460 211 461 212 
<< pdiffusion >>
rect 462 211 463 212 
<< pdiffusion >>
rect 463 211 464 212 
<< pdiffusion >>
rect 464 211 465 212 
<< pdiffusion >>
rect 465 211 466 212 
<< pdiffusion >>
rect 466 211 467 212 
<< pdiffusion >>
rect 467 211 468 212 
<< pdiffusion >>
rect 480 211 481 212 
<< pdiffusion >>
rect 481 211 482 212 
<< pdiffusion >>
rect 482 211 483 212 
<< pdiffusion >>
rect 483 211 484 212 
<< pdiffusion >>
rect 484 211 485 212 
<< pdiffusion >>
rect 485 211 486 212 
<< pdiffusion >>
rect 498 211 499 212 
<< pdiffusion >>
rect 499 211 500 212 
<< pdiffusion >>
rect 500 211 501 212 
<< pdiffusion >>
rect 501 211 502 212 
<< pdiffusion >>
rect 502 211 503 212 
<< pdiffusion >>
rect 503 211 504 212 
<< pdiffusion >>
rect 516 211 517 212 
<< pdiffusion >>
rect 517 211 518 212 
<< pdiffusion >>
rect 518 211 519 212 
<< pdiffusion >>
rect 519 211 520 212 
<< pdiffusion >>
rect 520 211 521 212 
<< pdiffusion >>
rect 521 211 522 212 
<< m1 >>
rect 523 211 524 212 
<< pdiffusion >>
rect 12 212 13 213 
<< pdiffusion >>
rect 13 212 14 213 
<< pdiffusion >>
rect 14 212 15 213 
<< pdiffusion >>
rect 15 212 16 213 
<< pdiffusion >>
rect 16 212 17 213 
<< pdiffusion >>
rect 17 212 18 213 
<< m2 >>
rect 27 212 28 213 
<< m1 >>
rect 28 212 29 213 
<< pdiffusion >>
rect 30 212 31 213 
<< pdiffusion >>
rect 31 212 32 213 
<< pdiffusion >>
rect 32 212 33 213 
<< pdiffusion >>
rect 33 212 34 213 
<< pdiffusion >>
rect 34 212 35 213 
<< pdiffusion >>
rect 35 212 36 213 
<< pdiffusion >>
rect 48 212 49 213 
<< pdiffusion >>
rect 49 212 50 213 
<< pdiffusion >>
rect 50 212 51 213 
<< pdiffusion >>
rect 51 212 52 213 
<< pdiffusion >>
rect 52 212 53 213 
<< pdiffusion >>
rect 53 212 54 213 
<< m1 >>
rect 64 212 65 213 
<< pdiffusion >>
rect 66 212 67 213 
<< pdiffusion >>
rect 67 212 68 213 
<< pdiffusion >>
rect 68 212 69 213 
<< pdiffusion >>
rect 69 212 70 213 
<< pdiffusion >>
rect 70 212 71 213 
<< pdiffusion >>
rect 71 212 72 213 
<< m1 >>
rect 73 212 74 213 
<< pdiffusion >>
rect 84 212 85 213 
<< pdiffusion >>
rect 85 212 86 213 
<< pdiffusion >>
rect 86 212 87 213 
<< pdiffusion >>
rect 87 212 88 213 
<< pdiffusion >>
rect 88 212 89 213 
<< pdiffusion >>
rect 89 212 90 213 
<< m1 >>
rect 100 212 101 213 
<< m2 >>
rect 100 212 101 213 
<< pdiffusion >>
rect 102 212 103 213 
<< pdiffusion >>
rect 103 212 104 213 
<< pdiffusion >>
rect 104 212 105 213 
<< pdiffusion >>
rect 105 212 106 213 
<< pdiffusion >>
rect 106 212 107 213 
<< pdiffusion >>
rect 107 212 108 213 
<< m1 >>
rect 127 212 128 213 
<< pdiffusion >>
rect 138 212 139 213 
<< pdiffusion >>
rect 139 212 140 213 
<< pdiffusion >>
rect 140 212 141 213 
<< pdiffusion >>
rect 141 212 142 213 
<< pdiffusion >>
rect 142 212 143 213 
<< pdiffusion >>
rect 143 212 144 213 
<< m1 >>
rect 145 212 146 213 
<< m1 >>
rect 148 212 149 213 
<< m1 >>
rect 150 212 151 213 
<< pdiffusion >>
rect 156 212 157 213 
<< pdiffusion >>
rect 157 212 158 213 
<< pdiffusion >>
rect 158 212 159 213 
<< pdiffusion >>
rect 159 212 160 213 
<< pdiffusion >>
rect 160 212 161 213 
<< pdiffusion >>
rect 161 212 162 213 
<< m1 >>
rect 163 212 164 213 
<< m1 >>
rect 172 212 173 213 
<< pdiffusion >>
rect 174 212 175 213 
<< pdiffusion >>
rect 175 212 176 213 
<< pdiffusion >>
rect 176 212 177 213 
<< pdiffusion >>
rect 177 212 178 213 
<< pdiffusion >>
rect 178 212 179 213 
<< pdiffusion >>
rect 179 212 180 213 
<< m1 >>
rect 181 212 182 213 
<< m1 >>
rect 185 212 186 213 
<< m1 >>
rect 190 212 191 213 
<< pdiffusion >>
rect 192 212 193 213 
<< pdiffusion >>
rect 193 212 194 213 
<< pdiffusion >>
rect 194 212 195 213 
<< pdiffusion >>
rect 195 212 196 213 
<< pdiffusion >>
rect 196 212 197 213 
<< pdiffusion >>
rect 197 212 198 213 
<< m1 >>
rect 205 212 206 213 
<< m1 >>
rect 207 212 208 213 
<< pdiffusion >>
rect 210 212 211 213 
<< pdiffusion >>
rect 211 212 212 213 
<< pdiffusion >>
rect 212 212 213 213 
<< pdiffusion >>
rect 213 212 214 213 
<< pdiffusion >>
rect 214 212 215 213 
<< pdiffusion >>
rect 215 212 216 213 
<< m1 >>
rect 217 212 218 213 
<< m1 >>
rect 221 212 222 213 
<< m2 >>
rect 225 212 226 213 
<< m1 >>
rect 226 212 227 213 
<< pdiffusion >>
rect 228 212 229 213 
<< pdiffusion >>
rect 229 212 230 213 
<< pdiffusion >>
rect 230 212 231 213 
<< pdiffusion >>
rect 231 212 232 213 
<< pdiffusion >>
rect 232 212 233 213 
<< pdiffusion >>
rect 233 212 234 213 
<< m1 >>
rect 235 212 236 213 
<< m2 >>
rect 243 212 244 213 
<< m1 >>
rect 244 212 245 213 
<< pdiffusion >>
rect 246 212 247 213 
<< pdiffusion >>
rect 247 212 248 213 
<< pdiffusion >>
rect 248 212 249 213 
<< pdiffusion >>
rect 249 212 250 213 
<< pdiffusion >>
rect 250 212 251 213 
<< pdiffusion >>
rect 251 212 252 213 
<< m1 >>
rect 253 212 254 213 
<< pdiffusion >>
rect 264 212 265 213 
<< pdiffusion >>
rect 265 212 266 213 
<< pdiffusion >>
rect 266 212 267 213 
<< pdiffusion >>
rect 267 212 268 213 
<< pdiffusion >>
rect 268 212 269 213 
<< pdiffusion >>
rect 269 212 270 213 
<< pdiffusion >>
rect 282 212 283 213 
<< pdiffusion >>
rect 283 212 284 213 
<< pdiffusion >>
rect 284 212 285 213 
<< pdiffusion >>
rect 285 212 286 213 
<< pdiffusion >>
rect 286 212 287 213 
<< pdiffusion >>
rect 287 212 288 213 
<< m1 >>
rect 296 212 297 213 
<< m1 >>
rect 298 212 299 213 
<< pdiffusion >>
rect 300 212 301 213 
<< pdiffusion >>
rect 301 212 302 213 
<< pdiffusion >>
rect 302 212 303 213 
<< pdiffusion >>
rect 303 212 304 213 
<< pdiffusion >>
rect 304 212 305 213 
<< pdiffusion >>
rect 305 212 306 213 
<< m1 >>
rect 316 212 317 213 
<< pdiffusion >>
rect 318 212 319 213 
<< pdiffusion >>
rect 319 212 320 213 
<< pdiffusion >>
rect 320 212 321 213 
<< pdiffusion >>
rect 321 212 322 213 
<< pdiffusion >>
rect 322 212 323 213 
<< pdiffusion >>
rect 323 212 324 213 
<< m1 >>
rect 330 212 331 213 
<< m1 >>
rect 334 212 335 213 
<< pdiffusion >>
rect 336 212 337 213 
<< pdiffusion >>
rect 337 212 338 213 
<< pdiffusion >>
rect 338 212 339 213 
<< pdiffusion >>
rect 339 212 340 213 
<< pdiffusion >>
rect 340 212 341 213 
<< pdiffusion >>
rect 341 212 342 213 
<< m1 >>
rect 343 212 344 213 
<< pdiffusion >>
rect 354 212 355 213 
<< pdiffusion >>
rect 355 212 356 213 
<< pdiffusion >>
rect 356 212 357 213 
<< pdiffusion >>
rect 357 212 358 213 
<< pdiffusion >>
rect 358 212 359 213 
<< pdiffusion >>
rect 359 212 360 213 
<< m1 >>
rect 361 212 362 213 
<< pdiffusion >>
rect 372 212 373 213 
<< pdiffusion >>
rect 373 212 374 213 
<< pdiffusion >>
rect 374 212 375 213 
<< pdiffusion >>
rect 375 212 376 213 
<< pdiffusion >>
rect 376 212 377 213 
<< pdiffusion >>
rect 377 212 378 213 
<< m1 >>
rect 379 212 380 213 
<< pdiffusion >>
rect 390 212 391 213 
<< pdiffusion >>
rect 391 212 392 213 
<< pdiffusion >>
rect 392 212 393 213 
<< pdiffusion >>
rect 393 212 394 213 
<< pdiffusion >>
rect 394 212 395 213 
<< pdiffusion >>
rect 395 212 396 213 
<< m1 >>
rect 402 212 403 213 
<< m1 >>
rect 404 212 405 213 
<< pdiffusion >>
rect 408 212 409 213 
<< pdiffusion >>
rect 409 212 410 213 
<< pdiffusion >>
rect 410 212 411 213 
<< pdiffusion >>
rect 411 212 412 213 
<< pdiffusion >>
rect 412 212 413 213 
<< pdiffusion >>
rect 413 212 414 213 
<< m1 >>
rect 416 212 417 213 
<< m1 >>
rect 418 212 419 213 
<< m1 >>
rect 420 212 421 213 
<< m1 >>
rect 423 212 424 213 
<< pdiffusion >>
rect 426 212 427 213 
<< pdiffusion >>
rect 427 212 428 213 
<< pdiffusion >>
rect 428 212 429 213 
<< pdiffusion >>
rect 429 212 430 213 
<< pdiffusion >>
rect 430 212 431 213 
<< pdiffusion >>
rect 431 212 432 213 
<< m1 >>
rect 433 212 434 213 
<< pdiffusion >>
rect 444 212 445 213 
<< pdiffusion >>
rect 445 212 446 213 
<< pdiffusion >>
rect 446 212 447 213 
<< pdiffusion >>
rect 447 212 448 213 
<< pdiffusion >>
rect 448 212 449 213 
<< pdiffusion >>
rect 449 212 450 213 
<< m1 >>
rect 456 212 457 213 
<< m1 >>
rect 458 212 459 213 
<< m1 >>
rect 460 212 461 213 
<< m2 >>
rect 460 212 461 213 
<< pdiffusion >>
rect 462 212 463 213 
<< pdiffusion >>
rect 463 212 464 213 
<< pdiffusion >>
rect 464 212 465 213 
<< pdiffusion >>
rect 465 212 466 213 
<< pdiffusion >>
rect 466 212 467 213 
<< pdiffusion >>
rect 467 212 468 213 
<< pdiffusion >>
rect 480 212 481 213 
<< pdiffusion >>
rect 481 212 482 213 
<< pdiffusion >>
rect 482 212 483 213 
<< pdiffusion >>
rect 483 212 484 213 
<< pdiffusion >>
rect 484 212 485 213 
<< pdiffusion >>
rect 485 212 486 213 
<< pdiffusion >>
rect 498 212 499 213 
<< pdiffusion >>
rect 499 212 500 213 
<< pdiffusion >>
rect 500 212 501 213 
<< pdiffusion >>
rect 501 212 502 213 
<< pdiffusion >>
rect 502 212 503 213 
<< pdiffusion >>
rect 503 212 504 213 
<< pdiffusion >>
rect 516 212 517 213 
<< pdiffusion >>
rect 517 212 518 213 
<< pdiffusion >>
rect 518 212 519 213 
<< pdiffusion >>
rect 519 212 520 213 
<< pdiffusion >>
rect 520 212 521 213 
<< pdiffusion >>
rect 521 212 522 213 
<< m1 >>
rect 523 212 524 213 
<< pdiffusion >>
rect 12 213 13 214 
<< pdiffusion >>
rect 13 213 14 214 
<< pdiffusion >>
rect 14 213 15 214 
<< pdiffusion >>
rect 15 213 16 214 
<< pdiffusion >>
rect 16 213 17 214 
<< pdiffusion >>
rect 17 213 18 214 
<< m2 >>
rect 27 213 28 214 
<< m1 >>
rect 28 213 29 214 
<< pdiffusion >>
rect 30 213 31 214 
<< pdiffusion >>
rect 31 213 32 214 
<< pdiffusion >>
rect 32 213 33 214 
<< pdiffusion >>
rect 33 213 34 214 
<< pdiffusion >>
rect 34 213 35 214 
<< pdiffusion >>
rect 35 213 36 214 
<< pdiffusion >>
rect 48 213 49 214 
<< pdiffusion >>
rect 49 213 50 214 
<< pdiffusion >>
rect 50 213 51 214 
<< pdiffusion >>
rect 51 213 52 214 
<< pdiffusion >>
rect 52 213 53 214 
<< pdiffusion >>
rect 53 213 54 214 
<< m1 >>
rect 64 213 65 214 
<< pdiffusion >>
rect 66 213 67 214 
<< pdiffusion >>
rect 67 213 68 214 
<< pdiffusion >>
rect 68 213 69 214 
<< pdiffusion >>
rect 69 213 70 214 
<< pdiffusion >>
rect 70 213 71 214 
<< pdiffusion >>
rect 71 213 72 214 
<< m1 >>
rect 73 213 74 214 
<< pdiffusion >>
rect 84 213 85 214 
<< pdiffusion >>
rect 85 213 86 214 
<< pdiffusion >>
rect 86 213 87 214 
<< pdiffusion >>
rect 87 213 88 214 
<< pdiffusion >>
rect 88 213 89 214 
<< pdiffusion >>
rect 89 213 90 214 
<< m1 >>
rect 100 213 101 214 
<< m2 >>
rect 100 213 101 214 
<< pdiffusion >>
rect 102 213 103 214 
<< pdiffusion >>
rect 103 213 104 214 
<< pdiffusion >>
rect 104 213 105 214 
<< pdiffusion >>
rect 105 213 106 214 
<< pdiffusion >>
rect 106 213 107 214 
<< pdiffusion >>
rect 107 213 108 214 
<< m1 >>
rect 127 213 128 214 
<< pdiffusion >>
rect 138 213 139 214 
<< pdiffusion >>
rect 139 213 140 214 
<< pdiffusion >>
rect 140 213 141 214 
<< pdiffusion >>
rect 141 213 142 214 
<< pdiffusion >>
rect 142 213 143 214 
<< pdiffusion >>
rect 143 213 144 214 
<< m1 >>
rect 145 213 146 214 
<< m1 >>
rect 148 213 149 214 
<< m1 >>
rect 150 213 151 214 
<< pdiffusion >>
rect 156 213 157 214 
<< pdiffusion >>
rect 157 213 158 214 
<< pdiffusion >>
rect 158 213 159 214 
<< pdiffusion >>
rect 159 213 160 214 
<< pdiffusion >>
rect 160 213 161 214 
<< pdiffusion >>
rect 161 213 162 214 
<< m1 >>
rect 163 213 164 214 
<< m1 >>
rect 172 213 173 214 
<< pdiffusion >>
rect 174 213 175 214 
<< pdiffusion >>
rect 175 213 176 214 
<< pdiffusion >>
rect 176 213 177 214 
<< pdiffusion >>
rect 177 213 178 214 
<< pdiffusion >>
rect 178 213 179 214 
<< pdiffusion >>
rect 179 213 180 214 
<< m1 >>
rect 181 213 182 214 
<< m1 >>
rect 185 213 186 214 
<< m1 >>
rect 190 213 191 214 
<< pdiffusion >>
rect 192 213 193 214 
<< pdiffusion >>
rect 193 213 194 214 
<< pdiffusion >>
rect 194 213 195 214 
<< pdiffusion >>
rect 195 213 196 214 
<< pdiffusion >>
rect 196 213 197 214 
<< pdiffusion >>
rect 197 213 198 214 
<< m1 >>
rect 205 213 206 214 
<< m1 >>
rect 207 213 208 214 
<< pdiffusion >>
rect 210 213 211 214 
<< pdiffusion >>
rect 211 213 212 214 
<< pdiffusion >>
rect 212 213 213 214 
<< pdiffusion >>
rect 213 213 214 214 
<< pdiffusion >>
rect 214 213 215 214 
<< pdiffusion >>
rect 215 213 216 214 
<< m1 >>
rect 217 213 218 214 
<< m1 >>
rect 221 213 222 214 
<< m2 >>
rect 225 213 226 214 
<< m1 >>
rect 226 213 227 214 
<< pdiffusion >>
rect 228 213 229 214 
<< pdiffusion >>
rect 229 213 230 214 
<< pdiffusion >>
rect 230 213 231 214 
<< pdiffusion >>
rect 231 213 232 214 
<< pdiffusion >>
rect 232 213 233 214 
<< pdiffusion >>
rect 233 213 234 214 
<< m1 >>
rect 235 213 236 214 
<< m2 >>
rect 243 213 244 214 
<< m1 >>
rect 244 213 245 214 
<< pdiffusion >>
rect 246 213 247 214 
<< pdiffusion >>
rect 247 213 248 214 
<< pdiffusion >>
rect 248 213 249 214 
<< pdiffusion >>
rect 249 213 250 214 
<< pdiffusion >>
rect 250 213 251 214 
<< pdiffusion >>
rect 251 213 252 214 
<< m1 >>
rect 253 213 254 214 
<< pdiffusion >>
rect 264 213 265 214 
<< pdiffusion >>
rect 265 213 266 214 
<< pdiffusion >>
rect 266 213 267 214 
<< pdiffusion >>
rect 267 213 268 214 
<< pdiffusion >>
rect 268 213 269 214 
<< pdiffusion >>
rect 269 213 270 214 
<< pdiffusion >>
rect 282 213 283 214 
<< pdiffusion >>
rect 283 213 284 214 
<< pdiffusion >>
rect 284 213 285 214 
<< pdiffusion >>
rect 285 213 286 214 
<< pdiffusion >>
rect 286 213 287 214 
<< pdiffusion >>
rect 287 213 288 214 
<< m1 >>
rect 296 213 297 214 
<< m1 >>
rect 298 213 299 214 
<< pdiffusion >>
rect 300 213 301 214 
<< pdiffusion >>
rect 301 213 302 214 
<< pdiffusion >>
rect 302 213 303 214 
<< pdiffusion >>
rect 303 213 304 214 
<< pdiffusion >>
rect 304 213 305 214 
<< pdiffusion >>
rect 305 213 306 214 
<< m1 >>
rect 316 213 317 214 
<< pdiffusion >>
rect 318 213 319 214 
<< pdiffusion >>
rect 319 213 320 214 
<< pdiffusion >>
rect 320 213 321 214 
<< pdiffusion >>
rect 321 213 322 214 
<< pdiffusion >>
rect 322 213 323 214 
<< pdiffusion >>
rect 323 213 324 214 
<< m1 >>
rect 330 213 331 214 
<< m1 >>
rect 334 213 335 214 
<< pdiffusion >>
rect 336 213 337 214 
<< pdiffusion >>
rect 337 213 338 214 
<< pdiffusion >>
rect 338 213 339 214 
<< pdiffusion >>
rect 339 213 340 214 
<< pdiffusion >>
rect 340 213 341 214 
<< pdiffusion >>
rect 341 213 342 214 
<< m1 >>
rect 343 213 344 214 
<< pdiffusion >>
rect 354 213 355 214 
<< pdiffusion >>
rect 355 213 356 214 
<< pdiffusion >>
rect 356 213 357 214 
<< pdiffusion >>
rect 357 213 358 214 
<< pdiffusion >>
rect 358 213 359 214 
<< pdiffusion >>
rect 359 213 360 214 
<< m1 >>
rect 361 213 362 214 
<< pdiffusion >>
rect 372 213 373 214 
<< pdiffusion >>
rect 373 213 374 214 
<< pdiffusion >>
rect 374 213 375 214 
<< pdiffusion >>
rect 375 213 376 214 
<< pdiffusion >>
rect 376 213 377 214 
<< pdiffusion >>
rect 377 213 378 214 
<< m1 >>
rect 379 213 380 214 
<< pdiffusion >>
rect 390 213 391 214 
<< pdiffusion >>
rect 391 213 392 214 
<< pdiffusion >>
rect 392 213 393 214 
<< pdiffusion >>
rect 393 213 394 214 
<< pdiffusion >>
rect 394 213 395 214 
<< pdiffusion >>
rect 395 213 396 214 
<< m1 >>
rect 402 213 403 214 
<< m1 >>
rect 404 213 405 214 
<< pdiffusion >>
rect 408 213 409 214 
<< pdiffusion >>
rect 409 213 410 214 
<< pdiffusion >>
rect 410 213 411 214 
<< pdiffusion >>
rect 411 213 412 214 
<< pdiffusion >>
rect 412 213 413 214 
<< pdiffusion >>
rect 413 213 414 214 
<< m1 >>
rect 416 213 417 214 
<< m1 >>
rect 418 213 419 214 
<< m1 >>
rect 420 213 421 214 
<< m1 >>
rect 423 213 424 214 
<< pdiffusion >>
rect 426 213 427 214 
<< pdiffusion >>
rect 427 213 428 214 
<< pdiffusion >>
rect 428 213 429 214 
<< pdiffusion >>
rect 429 213 430 214 
<< pdiffusion >>
rect 430 213 431 214 
<< pdiffusion >>
rect 431 213 432 214 
<< m1 >>
rect 433 213 434 214 
<< pdiffusion >>
rect 444 213 445 214 
<< pdiffusion >>
rect 445 213 446 214 
<< pdiffusion >>
rect 446 213 447 214 
<< pdiffusion >>
rect 447 213 448 214 
<< pdiffusion >>
rect 448 213 449 214 
<< pdiffusion >>
rect 449 213 450 214 
<< m1 >>
rect 456 213 457 214 
<< m1 >>
rect 458 213 459 214 
<< m1 >>
rect 460 213 461 214 
<< m2 >>
rect 460 213 461 214 
<< pdiffusion >>
rect 462 213 463 214 
<< pdiffusion >>
rect 463 213 464 214 
<< pdiffusion >>
rect 464 213 465 214 
<< pdiffusion >>
rect 465 213 466 214 
<< pdiffusion >>
rect 466 213 467 214 
<< pdiffusion >>
rect 467 213 468 214 
<< pdiffusion >>
rect 480 213 481 214 
<< pdiffusion >>
rect 481 213 482 214 
<< pdiffusion >>
rect 482 213 483 214 
<< pdiffusion >>
rect 483 213 484 214 
<< pdiffusion >>
rect 484 213 485 214 
<< pdiffusion >>
rect 485 213 486 214 
<< pdiffusion >>
rect 498 213 499 214 
<< pdiffusion >>
rect 499 213 500 214 
<< pdiffusion >>
rect 500 213 501 214 
<< pdiffusion >>
rect 501 213 502 214 
<< pdiffusion >>
rect 502 213 503 214 
<< pdiffusion >>
rect 503 213 504 214 
<< pdiffusion >>
rect 516 213 517 214 
<< pdiffusion >>
rect 517 213 518 214 
<< pdiffusion >>
rect 518 213 519 214 
<< pdiffusion >>
rect 519 213 520 214 
<< pdiffusion >>
rect 520 213 521 214 
<< pdiffusion >>
rect 521 213 522 214 
<< m1 >>
rect 523 213 524 214 
<< pdiffusion >>
rect 12 214 13 215 
<< pdiffusion >>
rect 13 214 14 215 
<< pdiffusion >>
rect 14 214 15 215 
<< pdiffusion >>
rect 15 214 16 215 
<< pdiffusion >>
rect 16 214 17 215 
<< pdiffusion >>
rect 17 214 18 215 
<< m2 >>
rect 27 214 28 215 
<< m1 >>
rect 28 214 29 215 
<< pdiffusion >>
rect 30 214 31 215 
<< pdiffusion >>
rect 31 214 32 215 
<< pdiffusion >>
rect 32 214 33 215 
<< pdiffusion >>
rect 33 214 34 215 
<< pdiffusion >>
rect 34 214 35 215 
<< pdiffusion >>
rect 35 214 36 215 
<< pdiffusion >>
rect 48 214 49 215 
<< pdiffusion >>
rect 49 214 50 215 
<< pdiffusion >>
rect 50 214 51 215 
<< pdiffusion >>
rect 51 214 52 215 
<< pdiffusion >>
rect 52 214 53 215 
<< pdiffusion >>
rect 53 214 54 215 
<< m1 >>
rect 64 214 65 215 
<< pdiffusion >>
rect 66 214 67 215 
<< pdiffusion >>
rect 67 214 68 215 
<< pdiffusion >>
rect 68 214 69 215 
<< pdiffusion >>
rect 69 214 70 215 
<< pdiffusion >>
rect 70 214 71 215 
<< pdiffusion >>
rect 71 214 72 215 
<< m1 >>
rect 73 214 74 215 
<< pdiffusion >>
rect 84 214 85 215 
<< pdiffusion >>
rect 85 214 86 215 
<< pdiffusion >>
rect 86 214 87 215 
<< pdiffusion >>
rect 87 214 88 215 
<< pdiffusion >>
rect 88 214 89 215 
<< pdiffusion >>
rect 89 214 90 215 
<< m1 >>
rect 100 214 101 215 
<< m2 >>
rect 100 214 101 215 
<< pdiffusion >>
rect 102 214 103 215 
<< pdiffusion >>
rect 103 214 104 215 
<< pdiffusion >>
rect 104 214 105 215 
<< pdiffusion >>
rect 105 214 106 215 
<< pdiffusion >>
rect 106 214 107 215 
<< pdiffusion >>
rect 107 214 108 215 
<< m1 >>
rect 127 214 128 215 
<< pdiffusion >>
rect 138 214 139 215 
<< pdiffusion >>
rect 139 214 140 215 
<< pdiffusion >>
rect 140 214 141 215 
<< pdiffusion >>
rect 141 214 142 215 
<< pdiffusion >>
rect 142 214 143 215 
<< pdiffusion >>
rect 143 214 144 215 
<< m1 >>
rect 145 214 146 215 
<< m1 >>
rect 148 214 149 215 
<< m1 >>
rect 150 214 151 215 
<< pdiffusion >>
rect 156 214 157 215 
<< pdiffusion >>
rect 157 214 158 215 
<< pdiffusion >>
rect 158 214 159 215 
<< pdiffusion >>
rect 159 214 160 215 
<< pdiffusion >>
rect 160 214 161 215 
<< pdiffusion >>
rect 161 214 162 215 
<< m1 >>
rect 163 214 164 215 
<< m1 >>
rect 172 214 173 215 
<< pdiffusion >>
rect 174 214 175 215 
<< pdiffusion >>
rect 175 214 176 215 
<< pdiffusion >>
rect 176 214 177 215 
<< pdiffusion >>
rect 177 214 178 215 
<< pdiffusion >>
rect 178 214 179 215 
<< pdiffusion >>
rect 179 214 180 215 
<< m1 >>
rect 181 214 182 215 
<< m1 >>
rect 185 214 186 215 
<< m1 >>
rect 190 214 191 215 
<< pdiffusion >>
rect 192 214 193 215 
<< pdiffusion >>
rect 193 214 194 215 
<< pdiffusion >>
rect 194 214 195 215 
<< pdiffusion >>
rect 195 214 196 215 
<< pdiffusion >>
rect 196 214 197 215 
<< pdiffusion >>
rect 197 214 198 215 
<< m1 >>
rect 205 214 206 215 
<< m1 >>
rect 207 214 208 215 
<< pdiffusion >>
rect 210 214 211 215 
<< pdiffusion >>
rect 211 214 212 215 
<< pdiffusion >>
rect 212 214 213 215 
<< pdiffusion >>
rect 213 214 214 215 
<< pdiffusion >>
rect 214 214 215 215 
<< pdiffusion >>
rect 215 214 216 215 
<< m1 >>
rect 217 214 218 215 
<< m1 >>
rect 221 214 222 215 
<< m2 >>
rect 225 214 226 215 
<< m1 >>
rect 226 214 227 215 
<< pdiffusion >>
rect 228 214 229 215 
<< pdiffusion >>
rect 229 214 230 215 
<< pdiffusion >>
rect 230 214 231 215 
<< pdiffusion >>
rect 231 214 232 215 
<< pdiffusion >>
rect 232 214 233 215 
<< pdiffusion >>
rect 233 214 234 215 
<< m1 >>
rect 235 214 236 215 
<< m2 >>
rect 243 214 244 215 
<< m1 >>
rect 244 214 245 215 
<< pdiffusion >>
rect 246 214 247 215 
<< pdiffusion >>
rect 247 214 248 215 
<< pdiffusion >>
rect 248 214 249 215 
<< pdiffusion >>
rect 249 214 250 215 
<< pdiffusion >>
rect 250 214 251 215 
<< pdiffusion >>
rect 251 214 252 215 
<< m1 >>
rect 253 214 254 215 
<< pdiffusion >>
rect 264 214 265 215 
<< pdiffusion >>
rect 265 214 266 215 
<< pdiffusion >>
rect 266 214 267 215 
<< pdiffusion >>
rect 267 214 268 215 
<< pdiffusion >>
rect 268 214 269 215 
<< pdiffusion >>
rect 269 214 270 215 
<< pdiffusion >>
rect 282 214 283 215 
<< pdiffusion >>
rect 283 214 284 215 
<< pdiffusion >>
rect 284 214 285 215 
<< pdiffusion >>
rect 285 214 286 215 
<< pdiffusion >>
rect 286 214 287 215 
<< pdiffusion >>
rect 287 214 288 215 
<< m1 >>
rect 296 214 297 215 
<< m1 >>
rect 298 214 299 215 
<< pdiffusion >>
rect 300 214 301 215 
<< pdiffusion >>
rect 301 214 302 215 
<< pdiffusion >>
rect 302 214 303 215 
<< pdiffusion >>
rect 303 214 304 215 
<< pdiffusion >>
rect 304 214 305 215 
<< pdiffusion >>
rect 305 214 306 215 
<< m1 >>
rect 316 214 317 215 
<< pdiffusion >>
rect 318 214 319 215 
<< pdiffusion >>
rect 319 214 320 215 
<< pdiffusion >>
rect 320 214 321 215 
<< pdiffusion >>
rect 321 214 322 215 
<< pdiffusion >>
rect 322 214 323 215 
<< pdiffusion >>
rect 323 214 324 215 
<< m1 >>
rect 330 214 331 215 
<< m1 >>
rect 334 214 335 215 
<< pdiffusion >>
rect 336 214 337 215 
<< pdiffusion >>
rect 337 214 338 215 
<< pdiffusion >>
rect 338 214 339 215 
<< pdiffusion >>
rect 339 214 340 215 
<< pdiffusion >>
rect 340 214 341 215 
<< pdiffusion >>
rect 341 214 342 215 
<< m1 >>
rect 343 214 344 215 
<< pdiffusion >>
rect 354 214 355 215 
<< pdiffusion >>
rect 355 214 356 215 
<< pdiffusion >>
rect 356 214 357 215 
<< pdiffusion >>
rect 357 214 358 215 
<< pdiffusion >>
rect 358 214 359 215 
<< pdiffusion >>
rect 359 214 360 215 
<< m1 >>
rect 361 214 362 215 
<< pdiffusion >>
rect 372 214 373 215 
<< pdiffusion >>
rect 373 214 374 215 
<< pdiffusion >>
rect 374 214 375 215 
<< pdiffusion >>
rect 375 214 376 215 
<< pdiffusion >>
rect 376 214 377 215 
<< pdiffusion >>
rect 377 214 378 215 
<< m1 >>
rect 379 214 380 215 
<< pdiffusion >>
rect 390 214 391 215 
<< pdiffusion >>
rect 391 214 392 215 
<< pdiffusion >>
rect 392 214 393 215 
<< pdiffusion >>
rect 393 214 394 215 
<< pdiffusion >>
rect 394 214 395 215 
<< pdiffusion >>
rect 395 214 396 215 
<< m1 >>
rect 402 214 403 215 
<< m1 >>
rect 404 214 405 215 
<< pdiffusion >>
rect 408 214 409 215 
<< pdiffusion >>
rect 409 214 410 215 
<< pdiffusion >>
rect 410 214 411 215 
<< pdiffusion >>
rect 411 214 412 215 
<< pdiffusion >>
rect 412 214 413 215 
<< pdiffusion >>
rect 413 214 414 215 
<< m1 >>
rect 416 214 417 215 
<< m1 >>
rect 418 214 419 215 
<< m1 >>
rect 420 214 421 215 
<< m1 >>
rect 423 214 424 215 
<< pdiffusion >>
rect 426 214 427 215 
<< pdiffusion >>
rect 427 214 428 215 
<< pdiffusion >>
rect 428 214 429 215 
<< pdiffusion >>
rect 429 214 430 215 
<< pdiffusion >>
rect 430 214 431 215 
<< pdiffusion >>
rect 431 214 432 215 
<< m1 >>
rect 433 214 434 215 
<< pdiffusion >>
rect 444 214 445 215 
<< pdiffusion >>
rect 445 214 446 215 
<< pdiffusion >>
rect 446 214 447 215 
<< pdiffusion >>
rect 447 214 448 215 
<< pdiffusion >>
rect 448 214 449 215 
<< pdiffusion >>
rect 449 214 450 215 
<< m1 >>
rect 456 214 457 215 
<< m1 >>
rect 458 214 459 215 
<< m1 >>
rect 460 214 461 215 
<< m2 >>
rect 460 214 461 215 
<< pdiffusion >>
rect 462 214 463 215 
<< pdiffusion >>
rect 463 214 464 215 
<< pdiffusion >>
rect 464 214 465 215 
<< pdiffusion >>
rect 465 214 466 215 
<< pdiffusion >>
rect 466 214 467 215 
<< pdiffusion >>
rect 467 214 468 215 
<< pdiffusion >>
rect 480 214 481 215 
<< pdiffusion >>
rect 481 214 482 215 
<< pdiffusion >>
rect 482 214 483 215 
<< pdiffusion >>
rect 483 214 484 215 
<< pdiffusion >>
rect 484 214 485 215 
<< pdiffusion >>
rect 485 214 486 215 
<< pdiffusion >>
rect 498 214 499 215 
<< pdiffusion >>
rect 499 214 500 215 
<< pdiffusion >>
rect 500 214 501 215 
<< pdiffusion >>
rect 501 214 502 215 
<< pdiffusion >>
rect 502 214 503 215 
<< pdiffusion >>
rect 503 214 504 215 
<< pdiffusion >>
rect 516 214 517 215 
<< pdiffusion >>
rect 517 214 518 215 
<< pdiffusion >>
rect 518 214 519 215 
<< pdiffusion >>
rect 519 214 520 215 
<< pdiffusion >>
rect 520 214 521 215 
<< pdiffusion >>
rect 521 214 522 215 
<< m1 >>
rect 523 214 524 215 
<< pdiffusion >>
rect 12 215 13 216 
<< m1 >>
rect 13 215 14 216 
<< pdiffusion >>
rect 13 215 14 216 
<< pdiffusion >>
rect 14 215 15 216 
<< pdiffusion >>
rect 15 215 16 216 
<< pdiffusion >>
rect 16 215 17 216 
<< pdiffusion >>
rect 17 215 18 216 
<< m2 >>
rect 27 215 28 216 
<< m1 >>
rect 28 215 29 216 
<< pdiffusion >>
rect 30 215 31 216 
<< pdiffusion >>
rect 31 215 32 216 
<< pdiffusion >>
rect 32 215 33 216 
<< pdiffusion >>
rect 33 215 34 216 
<< pdiffusion >>
rect 34 215 35 216 
<< pdiffusion >>
rect 35 215 36 216 
<< pdiffusion >>
rect 48 215 49 216 
<< pdiffusion >>
rect 49 215 50 216 
<< pdiffusion >>
rect 50 215 51 216 
<< pdiffusion >>
rect 51 215 52 216 
<< pdiffusion >>
rect 52 215 53 216 
<< pdiffusion >>
rect 53 215 54 216 
<< m1 >>
rect 64 215 65 216 
<< pdiffusion >>
rect 66 215 67 216 
<< pdiffusion >>
rect 67 215 68 216 
<< pdiffusion >>
rect 68 215 69 216 
<< pdiffusion >>
rect 69 215 70 216 
<< pdiffusion >>
rect 70 215 71 216 
<< pdiffusion >>
rect 71 215 72 216 
<< m1 >>
rect 73 215 74 216 
<< pdiffusion >>
rect 84 215 85 216 
<< m1 >>
rect 85 215 86 216 
<< pdiffusion >>
rect 85 215 86 216 
<< pdiffusion >>
rect 86 215 87 216 
<< pdiffusion >>
rect 87 215 88 216 
<< pdiffusion >>
rect 88 215 89 216 
<< pdiffusion >>
rect 89 215 90 216 
<< m1 >>
rect 100 215 101 216 
<< m2 >>
rect 100 215 101 216 
<< pdiffusion >>
rect 102 215 103 216 
<< pdiffusion >>
rect 103 215 104 216 
<< pdiffusion >>
rect 104 215 105 216 
<< pdiffusion >>
rect 105 215 106 216 
<< pdiffusion >>
rect 106 215 107 216 
<< pdiffusion >>
rect 107 215 108 216 
<< m1 >>
rect 127 215 128 216 
<< pdiffusion >>
rect 138 215 139 216 
<< pdiffusion >>
rect 139 215 140 216 
<< pdiffusion >>
rect 140 215 141 216 
<< pdiffusion >>
rect 141 215 142 216 
<< pdiffusion >>
rect 142 215 143 216 
<< pdiffusion >>
rect 143 215 144 216 
<< m1 >>
rect 145 215 146 216 
<< m1 >>
rect 148 215 149 216 
<< m1 >>
rect 150 215 151 216 
<< pdiffusion >>
rect 156 215 157 216 
<< pdiffusion >>
rect 157 215 158 216 
<< pdiffusion >>
rect 158 215 159 216 
<< pdiffusion >>
rect 159 215 160 216 
<< pdiffusion >>
rect 160 215 161 216 
<< pdiffusion >>
rect 161 215 162 216 
<< m1 >>
rect 163 215 164 216 
<< m1 >>
rect 172 215 173 216 
<< pdiffusion >>
rect 174 215 175 216 
<< pdiffusion >>
rect 175 215 176 216 
<< pdiffusion >>
rect 176 215 177 216 
<< pdiffusion >>
rect 177 215 178 216 
<< pdiffusion >>
rect 178 215 179 216 
<< pdiffusion >>
rect 179 215 180 216 
<< m1 >>
rect 181 215 182 216 
<< m1 >>
rect 185 215 186 216 
<< m1 >>
rect 190 215 191 216 
<< pdiffusion >>
rect 192 215 193 216 
<< pdiffusion >>
rect 193 215 194 216 
<< pdiffusion >>
rect 194 215 195 216 
<< pdiffusion >>
rect 195 215 196 216 
<< pdiffusion >>
rect 196 215 197 216 
<< pdiffusion >>
rect 197 215 198 216 
<< m1 >>
rect 205 215 206 216 
<< m1 >>
rect 207 215 208 216 
<< pdiffusion >>
rect 210 215 211 216 
<< pdiffusion >>
rect 211 215 212 216 
<< pdiffusion >>
rect 212 215 213 216 
<< pdiffusion >>
rect 213 215 214 216 
<< pdiffusion >>
rect 214 215 215 216 
<< pdiffusion >>
rect 215 215 216 216 
<< m1 >>
rect 217 215 218 216 
<< m1 >>
rect 221 215 222 216 
<< m2 >>
rect 225 215 226 216 
<< m1 >>
rect 226 215 227 216 
<< pdiffusion >>
rect 228 215 229 216 
<< pdiffusion >>
rect 229 215 230 216 
<< pdiffusion >>
rect 230 215 231 216 
<< pdiffusion >>
rect 231 215 232 216 
<< m1 >>
rect 232 215 233 216 
<< pdiffusion >>
rect 232 215 233 216 
<< pdiffusion >>
rect 233 215 234 216 
<< m1 >>
rect 235 215 236 216 
<< m2 >>
rect 243 215 244 216 
<< m1 >>
rect 244 215 245 216 
<< pdiffusion >>
rect 246 215 247 216 
<< pdiffusion >>
rect 247 215 248 216 
<< pdiffusion >>
rect 248 215 249 216 
<< pdiffusion >>
rect 249 215 250 216 
<< pdiffusion >>
rect 250 215 251 216 
<< pdiffusion >>
rect 251 215 252 216 
<< m1 >>
rect 253 215 254 216 
<< pdiffusion >>
rect 264 215 265 216 
<< pdiffusion >>
rect 265 215 266 216 
<< pdiffusion >>
rect 266 215 267 216 
<< pdiffusion >>
rect 267 215 268 216 
<< pdiffusion >>
rect 268 215 269 216 
<< pdiffusion >>
rect 269 215 270 216 
<< pdiffusion >>
rect 282 215 283 216 
<< m1 >>
rect 283 215 284 216 
<< pdiffusion >>
rect 283 215 284 216 
<< pdiffusion >>
rect 284 215 285 216 
<< pdiffusion >>
rect 285 215 286 216 
<< pdiffusion >>
rect 286 215 287 216 
<< pdiffusion >>
rect 287 215 288 216 
<< m1 >>
rect 296 215 297 216 
<< m1 >>
rect 298 215 299 216 
<< pdiffusion >>
rect 300 215 301 216 
<< pdiffusion >>
rect 301 215 302 216 
<< pdiffusion >>
rect 302 215 303 216 
<< pdiffusion >>
rect 303 215 304 216 
<< m1 >>
rect 304 215 305 216 
<< pdiffusion >>
rect 304 215 305 216 
<< pdiffusion >>
rect 305 215 306 216 
<< m1 >>
rect 316 215 317 216 
<< pdiffusion >>
rect 318 215 319 216 
<< m1 >>
rect 319 215 320 216 
<< pdiffusion >>
rect 319 215 320 216 
<< pdiffusion >>
rect 320 215 321 216 
<< pdiffusion >>
rect 321 215 322 216 
<< pdiffusion >>
rect 322 215 323 216 
<< pdiffusion >>
rect 323 215 324 216 
<< m1 >>
rect 330 215 331 216 
<< m1 >>
rect 334 215 335 216 
<< pdiffusion >>
rect 336 215 337 216 
<< pdiffusion >>
rect 337 215 338 216 
<< pdiffusion >>
rect 338 215 339 216 
<< pdiffusion >>
rect 339 215 340 216 
<< m1 >>
rect 340 215 341 216 
<< pdiffusion >>
rect 340 215 341 216 
<< pdiffusion >>
rect 341 215 342 216 
<< m1 >>
rect 343 215 344 216 
<< pdiffusion >>
rect 354 215 355 216 
<< pdiffusion >>
rect 355 215 356 216 
<< pdiffusion >>
rect 356 215 357 216 
<< pdiffusion >>
rect 357 215 358 216 
<< pdiffusion >>
rect 358 215 359 216 
<< pdiffusion >>
rect 359 215 360 216 
<< m1 >>
rect 361 215 362 216 
<< pdiffusion >>
rect 372 215 373 216 
<< pdiffusion >>
rect 373 215 374 216 
<< pdiffusion >>
rect 374 215 375 216 
<< pdiffusion >>
rect 375 215 376 216 
<< pdiffusion >>
rect 376 215 377 216 
<< pdiffusion >>
rect 377 215 378 216 
<< m1 >>
rect 379 215 380 216 
<< pdiffusion >>
rect 390 215 391 216 
<< pdiffusion >>
rect 391 215 392 216 
<< pdiffusion >>
rect 392 215 393 216 
<< pdiffusion >>
rect 393 215 394 216 
<< pdiffusion >>
rect 394 215 395 216 
<< pdiffusion >>
rect 395 215 396 216 
<< m1 >>
rect 402 215 403 216 
<< m1 >>
rect 404 215 405 216 
<< pdiffusion >>
rect 408 215 409 216 
<< pdiffusion >>
rect 409 215 410 216 
<< pdiffusion >>
rect 410 215 411 216 
<< pdiffusion >>
rect 411 215 412 216 
<< pdiffusion >>
rect 412 215 413 216 
<< pdiffusion >>
rect 413 215 414 216 
<< m1 >>
rect 416 215 417 216 
<< m1 >>
rect 418 215 419 216 
<< m1 >>
rect 420 215 421 216 
<< m2 >>
rect 420 215 421 216 
<< m2c >>
rect 420 215 421 216 
<< m1 >>
rect 420 215 421 216 
<< m2 >>
rect 420 215 421 216 
<< m1 >>
rect 423 215 424 216 
<< m2 >>
rect 423 215 424 216 
<< m2c >>
rect 423 215 424 216 
<< m1 >>
rect 423 215 424 216 
<< m2 >>
rect 423 215 424 216 
<< pdiffusion >>
rect 426 215 427 216 
<< m1 >>
rect 427 215 428 216 
<< pdiffusion >>
rect 427 215 428 216 
<< pdiffusion >>
rect 428 215 429 216 
<< pdiffusion >>
rect 429 215 430 216 
<< pdiffusion >>
rect 430 215 431 216 
<< pdiffusion >>
rect 431 215 432 216 
<< m1 >>
rect 433 215 434 216 
<< pdiffusion >>
rect 444 215 445 216 
<< pdiffusion >>
rect 445 215 446 216 
<< pdiffusion >>
rect 446 215 447 216 
<< pdiffusion >>
rect 447 215 448 216 
<< pdiffusion >>
rect 448 215 449 216 
<< pdiffusion >>
rect 449 215 450 216 
<< m1 >>
rect 456 215 457 216 
<< m1 >>
rect 458 215 459 216 
<< m1 >>
rect 460 215 461 216 
<< m2 >>
rect 460 215 461 216 
<< pdiffusion >>
rect 462 215 463 216 
<< m1 >>
rect 463 215 464 216 
<< pdiffusion >>
rect 463 215 464 216 
<< pdiffusion >>
rect 464 215 465 216 
<< pdiffusion >>
rect 465 215 466 216 
<< pdiffusion >>
rect 466 215 467 216 
<< pdiffusion >>
rect 467 215 468 216 
<< pdiffusion >>
rect 480 215 481 216 
<< pdiffusion >>
rect 481 215 482 216 
<< pdiffusion >>
rect 482 215 483 216 
<< pdiffusion >>
rect 483 215 484 216 
<< m1 >>
rect 484 215 485 216 
<< pdiffusion >>
rect 484 215 485 216 
<< pdiffusion >>
rect 485 215 486 216 
<< pdiffusion >>
rect 498 215 499 216 
<< pdiffusion >>
rect 499 215 500 216 
<< pdiffusion >>
rect 500 215 501 216 
<< pdiffusion >>
rect 501 215 502 216 
<< pdiffusion >>
rect 502 215 503 216 
<< pdiffusion >>
rect 503 215 504 216 
<< pdiffusion >>
rect 516 215 517 216 
<< pdiffusion >>
rect 517 215 518 216 
<< pdiffusion >>
rect 518 215 519 216 
<< pdiffusion >>
rect 519 215 520 216 
<< pdiffusion >>
rect 520 215 521 216 
<< pdiffusion >>
rect 521 215 522 216 
<< m1 >>
rect 523 215 524 216 
<< m1 >>
rect 13 216 14 217 
<< m2 >>
rect 27 216 28 217 
<< m1 >>
rect 28 216 29 217 
<< m1 >>
rect 64 216 65 217 
<< m1 >>
rect 73 216 74 217 
<< m1 >>
rect 85 216 86 217 
<< m1 >>
rect 100 216 101 217 
<< m2 >>
rect 100 216 101 217 
<< m1 >>
rect 127 216 128 217 
<< m1 >>
rect 145 216 146 217 
<< m1 >>
rect 148 216 149 217 
<< m1 >>
rect 150 216 151 217 
<< m1 >>
rect 163 216 164 217 
<< m1 >>
rect 172 216 173 217 
<< m1 >>
rect 181 216 182 217 
<< m1 >>
rect 185 216 186 217 
<< m1 >>
rect 190 216 191 217 
<< m1 >>
rect 205 216 206 217 
<< m1 >>
rect 207 216 208 217 
<< m1 >>
rect 217 216 218 217 
<< m1 >>
rect 221 216 222 217 
<< m2 >>
rect 225 216 226 217 
<< m1 >>
rect 226 216 227 217 
<< m1 >>
rect 232 216 233 217 
<< m1 >>
rect 235 216 236 217 
<< m2 >>
rect 243 216 244 217 
<< m1 >>
rect 244 216 245 217 
<< m1 >>
rect 253 216 254 217 
<< m1 >>
rect 283 216 284 217 
<< m1 >>
rect 296 216 297 217 
<< m1 >>
rect 298 216 299 217 
<< m1 >>
rect 304 216 305 217 
<< m1 >>
rect 316 216 317 217 
<< m1 >>
rect 319 216 320 217 
<< m1 >>
rect 330 216 331 217 
<< m1 >>
rect 331 216 332 217 
<< m1 >>
rect 332 216 333 217 
<< m2 >>
rect 332 216 333 217 
<< m2c >>
rect 332 216 333 217 
<< m1 >>
rect 332 216 333 217 
<< m2 >>
rect 332 216 333 217 
<< m2 >>
rect 333 216 334 217 
<< m1 >>
rect 334 216 335 217 
<< m2 >>
rect 334 216 335 217 
<< m1 >>
rect 340 216 341 217 
<< m1 >>
rect 343 216 344 217 
<< m1 >>
rect 361 216 362 217 
<< m1 >>
rect 379 216 380 217 
<< m1 >>
rect 402 216 403 217 
<< m1 >>
rect 404 216 405 217 
<< m1 >>
rect 416 216 417 217 
<< m1 >>
rect 418 216 419 217 
<< m2 >>
rect 420 216 421 217 
<< m2 >>
rect 423 216 424 217 
<< m1 >>
rect 427 216 428 217 
<< m1 >>
rect 433 216 434 217 
<< m1 >>
rect 456 216 457 217 
<< m1 >>
rect 458 216 459 217 
<< m1 >>
rect 460 216 461 217 
<< m2 >>
rect 460 216 461 217 
<< m1 >>
rect 463 216 464 217 
<< m1 >>
rect 484 216 485 217 
<< m1 >>
rect 523 216 524 217 
<< m1 >>
rect 13 217 14 218 
<< m2 >>
rect 27 217 28 218 
<< m1 >>
rect 28 217 29 218 
<< m1 >>
rect 64 217 65 218 
<< m1 >>
rect 73 217 74 218 
<< m1 >>
rect 85 217 86 218 
<< m1 >>
rect 100 217 101 218 
<< m2 >>
rect 100 217 101 218 
<< m1 >>
rect 127 217 128 218 
<< m1 >>
rect 145 217 146 218 
<< m1 >>
rect 148 217 149 218 
<< m1 >>
rect 150 217 151 218 
<< m1 >>
rect 163 217 164 218 
<< m1 >>
rect 172 217 173 218 
<< m1 >>
rect 181 217 182 218 
<< m1 >>
rect 185 217 186 218 
<< m1 >>
rect 190 217 191 218 
<< m1 >>
rect 205 217 206 218 
<< m1 >>
rect 207 217 208 218 
<< m1 >>
rect 215 217 216 218 
<< m2 >>
rect 215 217 216 218 
<< m2c >>
rect 215 217 216 218 
<< m1 >>
rect 215 217 216 218 
<< m2 >>
rect 215 217 216 218 
<< m1 >>
rect 216 217 217 218 
<< m1 >>
rect 217 217 218 218 
<< m1 >>
rect 221 217 222 218 
<< m2 >>
rect 221 217 222 218 
<< m2c >>
rect 221 217 222 218 
<< m1 >>
rect 221 217 222 218 
<< m2 >>
rect 221 217 222 218 
<< m2 >>
rect 225 217 226 218 
<< m1 >>
rect 226 217 227 218 
<< m1 >>
rect 232 217 233 218 
<< m1 >>
rect 235 217 236 218 
<< m2 >>
rect 243 217 244 218 
<< m1 >>
rect 244 217 245 218 
<< m2 >>
rect 244 217 245 218 
<< m2 >>
rect 245 217 246 218 
<< m1 >>
rect 246 217 247 218 
<< m2 >>
rect 246 217 247 218 
<< m2c >>
rect 246 217 247 218 
<< m1 >>
rect 246 217 247 218 
<< m2 >>
rect 246 217 247 218 
<< m1 >>
rect 253 217 254 218 
<< m1 >>
rect 283 217 284 218 
<< m1 >>
rect 287 217 288 218 
<< m1 >>
rect 288 217 289 218 
<< m2 >>
rect 288 217 289 218 
<< m2c >>
rect 288 217 289 218 
<< m1 >>
rect 288 217 289 218 
<< m2 >>
rect 288 217 289 218 
<< m2 >>
rect 289 217 290 218 
<< m1 >>
rect 290 217 291 218 
<< m2 >>
rect 290 217 291 218 
<< m1 >>
rect 291 217 292 218 
<< m2 >>
rect 291 217 292 218 
<< m1 >>
rect 292 217 293 218 
<< m2 >>
rect 292 217 293 218 
<< m1 >>
rect 293 217 294 218 
<< m1 >>
rect 294 217 295 218 
<< m2 >>
rect 294 217 295 218 
<< m2c >>
rect 294 217 295 218 
<< m1 >>
rect 294 217 295 218 
<< m2 >>
rect 294 217 295 218 
<< m2 >>
rect 295 217 296 218 
<< m1 >>
rect 296 217 297 218 
<< m2 >>
rect 296 217 297 218 
<< m2 >>
rect 297 217 298 218 
<< m1 >>
rect 298 217 299 218 
<< m2 >>
rect 298 217 299 218 
<< m2c >>
rect 298 217 299 218 
<< m1 >>
rect 298 217 299 218 
<< m2 >>
rect 298 217 299 218 
<< m1 >>
rect 304 217 305 218 
<< m1 >>
rect 316 217 317 218 
<< m1 >>
rect 319 217 320 218 
<< m1 >>
rect 334 217 335 218 
<< m2 >>
rect 334 217 335 218 
<< m1 >>
rect 340 217 341 218 
<< m1 >>
rect 341 217 342 218 
<< m2 >>
rect 341 217 342 218 
<< m2c >>
rect 341 217 342 218 
<< m1 >>
rect 341 217 342 218 
<< m2 >>
rect 341 217 342 218 
<< m2 >>
rect 342 217 343 218 
<< m1 >>
rect 343 217 344 218 
<< m2 >>
rect 343 217 344 218 
<< m2 >>
rect 344 217 345 218 
<< m1 >>
rect 345 217 346 218 
<< m2 >>
rect 345 217 346 218 
<< m2c >>
rect 345 217 346 218 
<< m1 >>
rect 345 217 346 218 
<< m2 >>
rect 345 217 346 218 
<< m1 >>
rect 361 217 362 218 
<< m1 >>
rect 379 217 380 218 
<< m1 >>
rect 402 217 403 218 
<< m1 >>
rect 404 217 405 218 
<< m1 >>
rect 416 217 417 218 
<< m1 >>
rect 418 217 419 218 
<< m1 >>
rect 419 217 420 218 
<< m1 >>
rect 420 217 421 218 
<< m2 >>
rect 420 217 421 218 
<< m1 >>
rect 421 217 422 218 
<< m1 >>
rect 422 217 423 218 
<< m1 >>
rect 423 217 424 218 
<< m2 >>
rect 423 217 424 218 
<< m1 >>
rect 424 217 425 218 
<< m1 >>
rect 425 217 426 218 
<< m1 >>
rect 426 217 427 218 
<< m1 >>
rect 427 217 428 218 
<< m1 >>
rect 433 217 434 218 
<< m1 >>
rect 456 217 457 218 
<< m2 >>
rect 456 217 457 218 
<< m2c >>
rect 456 217 457 218 
<< m1 >>
rect 456 217 457 218 
<< m2 >>
rect 456 217 457 218 
<< m1 >>
rect 458 217 459 218 
<< m2 >>
rect 458 217 459 218 
<< m2c >>
rect 458 217 459 218 
<< m1 >>
rect 458 217 459 218 
<< m2 >>
rect 458 217 459 218 
<< m1 >>
rect 460 217 461 218 
<< m2 >>
rect 460 217 461 218 
<< m1 >>
rect 461 217 462 218 
<< m1 >>
rect 462 217 463 218 
<< m1 >>
rect 463 217 464 218 
<< m1 >>
rect 484 217 485 218 
<< m1 >>
rect 523 217 524 218 
<< m1 >>
rect 13 218 14 219 
<< m1 >>
rect 14 218 15 219 
<< m1 >>
rect 15 218 16 219 
<< m1 >>
rect 16 218 17 219 
<< m1 >>
rect 17 218 18 219 
<< m1 >>
rect 18 218 19 219 
<< m1 >>
rect 19 218 20 219 
<< m1 >>
rect 20 218 21 219 
<< m1 >>
rect 21 218 22 219 
<< m1 >>
rect 22 218 23 219 
<< m1 >>
rect 23 218 24 219 
<< m1 >>
rect 24 218 25 219 
<< m1 >>
rect 25 218 26 219 
<< m1 >>
rect 26 218 27 219 
<< m1 >>
rect 27 218 28 219 
<< m2 >>
rect 27 218 28 219 
<< m1 >>
rect 28 218 29 219 
<< m1 >>
rect 64 218 65 219 
<< m1 >>
rect 73 218 74 219 
<< m1 >>
rect 85 218 86 219 
<< m1 >>
rect 86 218 87 219 
<< m1 >>
rect 87 218 88 219 
<< m1 >>
rect 88 218 89 219 
<< m1 >>
rect 89 218 90 219 
<< m1 >>
rect 90 218 91 219 
<< m1 >>
rect 91 218 92 219 
<< m1 >>
rect 92 218 93 219 
<< m1 >>
rect 93 218 94 219 
<< m1 >>
rect 94 218 95 219 
<< m1 >>
rect 95 218 96 219 
<< m1 >>
rect 96 218 97 219 
<< m1 >>
rect 97 218 98 219 
<< m1 >>
rect 98 218 99 219 
<< m1 >>
rect 99 218 100 219 
<< m1 >>
rect 100 218 101 219 
<< m2 >>
rect 100 218 101 219 
<< m1 >>
rect 127 218 128 219 
<< m1 >>
rect 145 218 146 219 
<< m1 >>
rect 148 218 149 219 
<< m1 >>
rect 150 218 151 219 
<< m1 >>
rect 163 218 164 219 
<< m1 >>
rect 172 218 173 219 
<< m1 >>
rect 181 218 182 219 
<< m1 >>
rect 185 218 186 219 
<< m1 >>
rect 190 218 191 219 
<< m1 >>
rect 205 218 206 219 
<< m1 >>
rect 207 218 208 219 
<< m2 >>
rect 215 218 216 219 
<< m2 >>
rect 221 218 222 219 
<< m2 >>
rect 225 218 226 219 
<< m1 >>
rect 226 218 227 219 
<< m1 >>
rect 232 218 233 219 
<< m1 >>
rect 235 218 236 219 
<< m1 >>
rect 244 218 245 219 
<< m1 >>
rect 246 218 247 219 
<< m1 >>
rect 253 218 254 219 
<< m1 >>
rect 283 218 284 219 
<< m1 >>
rect 287 218 288 219 
<< m1 >>
rect 290 218 291 219 
<< m2 >>
rect 292 218 293 219 
<< m1 >>
rect 296 218 297 219 
<< m1 >>
rect 304 218 305 219 
<< m1 >>
rect 316 218 317 219 
<< m1 >>
rect 319 218 320 219 
<< m2 >>
rect 320 218 321 219 
<< m1 >>
rect 321 218 322 219 
<< m2 >>
rect 321 218 322 219 
<< m2c >>
rect 321 218 322 219 
<< m1 >>
rect 321 218 322 219 
<< m2 >>
rect 321 218 322 219 
<< m1 >>
rect 322 218 323 219 
<< m1 >>
rect 323 218 324 219 
<< m1 >>
rect 324 218 325 219 
<< m1 >>
rect 325 218 326 219 
<< m1 >>
rect 326 218 327 219 
<< m1 >>
rect 327 218 328 219 
<< m1 >>
rect 328 218 329 219 
<< m1 >>
rect 329 218 330 219 
<< m1 >>
rect 330 218 331 219 
<< m1 >>
rect 331 218 332 219 
<< m1 >>
rect 332 218 333 219 
<< m1 >>
rect 333 218 334 219 
<< m1 >>
rect 334 218 335 219 
<< m2 >>
rect 334 218 335 219 
<< m1 >>
rect 343 218 344 219 
<< m1 >>
rect 345 218 346 219 
<< m1 >>
rect 361 218 362 219 
<< m1 >>
rect 374 218 375 219 
<< m2 >>
rect 374 218 375 219 
<< m2c >>
rect 374 218 375 219 
<< m1 >>
rect 374 218 375 219 
<< m2 >>
rect 374 218 375 219 
<< m1 >>
rect 375 218 376 219 
<< m1 >>
rect 376 218 377 219 
<< m1 >>
rect 377 218 378 219 
<< m2 >>
rect 377 218 378 219 
<< m2c >>
rect 377 218 378 219 
<< m1 >>
rect 377 218 378 219 
<< m2 >>
rect 377 218 378 219 
<< m2 >>
rect 378 218 379 219 
<< m1 >>
rect 379 218 380 219 
<< m2 >>
rect 379 218 380 219 
<< m2 >>
rect 380 218 381 219 
<< m1 >>
rect 381 218 382 219 
<< m2 >>
rect 381 218 382 219 
<< m2c >>
rect 381 218 382 219 
<< m1 >>
rect 381 218 382 219 
<< m2 >>
rect 381 218 382 219 
<< m1 >>
rect 382 218 383 219 
<< m1 >>
rect 383 218 384 219 
<< m2 >>
rect 383 218 384 219 
<< m2c >>
rect 383 218 384 219 
<< m1 >>
rect 383 218 384 219 
<< m2 >>
rect 383 218 384 219 
<< m1 >>
rect 402 218 403 219 
<< m2 >>
rect 402 218 403 219 
<< m2c >>
rect 402 218 403 219 
<< m1 >>
rect 402 218 403 219 
<< m2 >>
rect 402 218 403 219 
<< m1 >>
rect 404 218 405 219 
<< m2 >>
rect 404 218 405 219 
<< m2c >>
rect 404 218 405 219 
<< m1 >>
rect 404 218 405 219 
<< m2 >>
rect 404 218 405 219 
<< m1 >>
rect 416 218 417 219 
<< m2 >>
rect 420 218 421 219 
<< m2 >>
rect 423 218 424 219 
<< m1 >>
rect 433 218 434 219 
<< m2 >>
rect 433 218 434 219 
<< m2c >>
rect 433 218 434 219 
<< m1 >>
rect 433 218 434 219 
<< m2 >>
rect 433 218 434 219 
<< m2 >>
rect 456 218 457 219 
<< m2 >>
rect 458 218 459 219 
<< m2 >>
rect 460 218 461 219 
<< m1 >>
rect 484 218 485 219 
<< m1 >>
rect 523 218 524 219 
<< m2 >>
rect 19 219 20 220 
<< m2 >>
rect 20 219 21 220 
<< m2 >>
rect 21 219 22 220 
<< m2 >>
rect 22 219 23 220 
<< m2 >>
rect 23 219 24 220 
<< m2 >>
rect 24 219 25 220 
<< m2 >>
rect 25 219 26 220 
<< m2 >>
rect 26 219 27 220 
<< m2 >>
rect 27 219 28 220 
<< m1 >>
rect 64 219 65 220 
<< m1 >>
rect 73 219 74 220 
<< m2 >>
rect 100 219 101 220 
<< m1 >>
rect 127 219 128 220 
<< m1 >>
rect 145 219 146 220 
<< m1 >>
rect 148 219 149 220 
<< m1 >>
rect 150 219 151 220 
<< m1 >>
rect 163 219 164 220 
<< m1 >>
rect 172 219 173 220 
<< m1 >>
rect 181 219 182 220 
<< m1 >>
rect 185 219 186 220 
<< m1 >>
rect 190 219 191 220 
<< m1 >>
rect 205 219 206 220 
<< m1 >>
rect 207 219 208 220 
<< m1 >>
rect 212 219 213 220 
<< m1 >>
rect 213 219 214 220 
<< m1 >>
rect 214 219 215 220 
<< m1 >>
rect 215 219 216 220 
<< m2 >>
rect 215 219 216 220 
<< m1 >>
rect 216 219 217 220 
<< m1 >>
rect 217 219 218 220 
<< m1 >>
rect 218 219 219 220 
<< m1 >>
rect 219 219 220 220 
<< m1 >>
rect 220 219 221 220 
<< m1 >>
rect 221 219 222 220 
<< m2 >>
rect 221 219 222 220 
<< m1 >>
rect 222 219 223 220 
<< m1 >>
rect 223 219 224 220 
<< m1 >>
rect 224 219 225 220 
<< m2 >>
rect 224 219 225 220 
<< m2c >>
rect 224 219 225 220 
<< m1 >>
rect 224 219 225 220 
<< m2 >>
rect 224 219 225 220 
<< m2 >>
rect 225 219 226 220 
<< m1 >>
rect 226 219 227 220 
<< m1 >>
rect 232 219 233 220 
<< m1 >>
rect 235 219 236 220 
<< m1 >>
rect 244 219 245 220 
<< m1 >>
rect 246 219 247 220 
<< m1 >>
rect 253 219 254 220 
<< m1 >>
rect 283 219 284 220 
<< m2 >>
rect 284 219 285 220 
<< m1 >>
rect 285 219 286 220 
<< m2 >>
rect 285 219 286 220 
<< m2c >>
rect 285 219 286 220 
<< m1 >>
rect 285 219 286 220 
<< m2 >>
rect 285 219 286 220 
<< m1 >>
rect 286 219 287 220 
<< m1 >>
rect 287 219 288 220 
<< m1 >>
rect 290 219 291 220 
<< m2 >>
rect 290 219 291 220 
<< m2c >>
rect 290 219 291 220 
<< m1 >>
rect 290 219 291 220 
<< m2 >>
rect 290 219 291 220 
<< m1 >>
rect 292 219 293 220 
<< m2 >>
rect 292 219 293 220 
<< m2c >>
rect 292 219 293 220 
<< m1 >>
rect 292 219 293 220 
<< m2 >>
rect 292 219 293 220 
<< m1 >>
rect 296 219 297 220 
<< m2 >>
rect 296 219 297 220 
<< m2c >>
rect 296 219 297 220 
<< m1 >>
rect 296 219 297 220 
<< m2 >>
rect 296 219 297 220 
<< m1 >>
rect 304 219 305 220 
<< m1 >>
rect 316 219 317 220 
<< m1 >>
rect 319 219 320 220 
<< m2 >>
rect 320 219 321 220 
<< m2 >>
rect 334 219 335 220 
<< m2 >>
rect 335 219 336 220 
<< m2 >>
rect 336 219 337 220 
<< m1 >>
rect 343 219 344 220 
<< m1 >>
rect 345 219 346 220 
<< m1 >>
rect 361 219 362 220 
<< m2 >>
rect 374 219 375 220 
<< m1 >>
rect 379 219 380 220 
<< m2 >>
rect 383 219 384 220 
<< m2 >>
rect 402 219 403 220 
<< m2 >>
rect 404 219 405 220 
<< m1 >>
rect 416 219 417 220 
<< m2 >>
rect 420 219 421 220 
<< m1 >>
rect 421 219 422 220 
<< m2 >>
rect 421 219 422 220 
<< m2c >>
rect 421 219 422 220 
<< m1 >>
rect 421 219 422 220 
<< m2 >>
rect 421 219 422 220 
<< m2 >>
rect 423 219 424 220 
<< m2 >>
rect 433 219 434 220 
<< m2 >>
rect 449 219 450 220 
<< m1 >>
rect 450 219 451 220 
<< m2 >>
rect 450 219 451 220 
<< m2c >>
rect 450 219 451 220 
<< m1 >>
rect 450 219 451 220 
<< m2 >>
rect 450 219 451 220 
<< m1 >>
rect 451 219 452 220 
<< m1 >>
rect 452 219 453 220 
<< m1 >>
rect 453 219 454 220 
<< m1 >>
rect 454 219 455 220 
<< m1 >>
rect 455 219 456 220 
<< m1 >>
rect 456 219 457 220 
<< m2 >>
rect 456 219 457 220 
<< m1 >>
rect 457 219 458 220 
<< m1 >>
rect 458 219 459 220 
<< m2 >>
rect 458 219 459 220 
<< m1 >>
rect 459 219 460 220 
<< m1 >>
rect 460 219 461 220 
<< m2 >>
rect 460 219 461 220 
<< m2c >>
rect 460 219 461 220 
<< m1 >>
rect 460 219 461 220 
<< m2 >>
rect 460 219 461 220 
<< m1 >>
rect 484 219 485 220 
<< m1 >>
rect 523 219 524 220 
<< m1 >>
rect 19 220 20 221 
<< m2 >>
rect 19 220 20 221 
<< m2c >>
rect 19 220 20 221 
<< m1 >>
rect 19 220 20 221 
<< m2 >>
rect 19 220 20 221 
<< m1 >>
rect 64 220 65 221 
<< m1 >>
rect 73 220 74 221 
<< m1 >>
rect 100 220 101 221 
<< m2 >>
rect 100 220 101 221 
<< m2c >>
rect 100 220 101 221 
<< m1 >>
rect 100 220 101 221 
<< m2 >>
rect 100 220 101 221 
<< m1 >>
rect 127 220 128 221 
<< m1 >>
rect 145 220 146 221 
<< m1 >>
rect 148 220 149 221 
<< m1 >>
rect 150 220 151 221 
<< m1 >>
rect 151 220 152 221 
<< m1 >>
rect 152 220 153 221 
<< m1 >>
rect 153 220 154 221 
<< m1 >>
rect 154 220 155 221 
<< m1 >>
rect 155 220 156 221 
<< m1 >>
rect 156 220 157 221 
<< m1 >>
rect 157 220 158 221 
<< m1 >>
rect 158 220 159 221 
<< m1 >>
rect 159 220 160 221 
<< m1 >>
rect 160 220 161 221 
<< m1 >>
rect 163 220 164 221 
<< m1 >>
rect 172 220 173 221 
<< m1 >>
rect 181 220 182 221 
<< m1 >>
rect 185 220 186 221 
<< m2 >>
rect 186 220 187 221 
<< m1 >>
rect 187 220 188 221 
<< m2 >>
rect 187 220 188 221 
<< m1 >>
rect 188 220 189 221 
<< m2 >>
rect 188 220 189 221 
<< m2c >>
rect 188 220 189 221 
<< m1 >>
rect 188 220 189 221 
<< m2 >>
rect 188 220 189 221 
<< m2 >>
rect 189 220 190 221 
<< m1 >>
rect 190 220 191 221 
<< m2 >>
rect 190 220 191 221 
<< m2 >>
rect 191 220 192 221 
<< m1 >>
rect 192 220 193 221 
<< m2 >>
rect 192 220 193 221 
<< m2c >>
rect 192 220 193 221 
<< m1 >>
rect 192 220 193 221 
<< m2 >>
rect 192 220 193 221 
<< m1 >>
rect 193 220 194 221 
<< m1 >>
rect 194 220 195 221 
<< m1 >>
rect 195 220 196 221 
<< m1 >>
rect 196 220 197 221 
<< m1 >>
rect 197 220 198 221 
<< m1 >>
rect 198 220 199 221 
<< m1 >>
rect 199 220 200 221 
<< m1 >>
rect 200 220 201 221 
<< m1 >>
rect 201 220 202 221 
<< m1 >>
rect 202 220 203 221 
<< m1 >>
rect 203 220 204 221 
<< m1 >>
rect 204 220 205 221 
<< m1 >>
rect 205 220 206 221 
<< m1 >>
rect 207 220 208 221 
<< m2 >>
rect 211 220 212 221 
<< m1 >>
rect 212 220 213 221 
<< m2 >>
rect 212 220 213 221 
<< m2 >>
rect 213 220 214 221 
<< m2 >>
rect 214 220 215 221 
<< m2 >>
rect 215 220 216 221 
<< m2 >>
rect 221 220 222 221 
<< m1 >>
rect 226 220 227 221 
<< m1 >>
rect 232 220 233 221 
<< m1 >>
rect 235 220 236 221 
<< m1 >>
rect 244 220 245 221 
<< m1 >>
rect 246 220 247 221 
<< m1 >>
rect 247 220 248 221 
<< m1 >>
rect 248 220 249 221 
<< m1 >>
rect 249 220 250 221 
<< m1 >>
rect 250 220 251 221 
<< m1 >>
rect 251 220 252 221 
<< m1 >>
rect 252 220 253 221 
<< m1 >>
rect 253 220 254 221 
<< m1 >>
rect 283 220 284 221 
<< m2 >>
rect 284 220 285 221 
<< m2 >>
rect 290 220 291 221 
<< m2 >>
rect 292 220 293 221 
<< m2 >>
rect 296 220 297 221 
<< m1 >>
rect 304 220 305 221 
<< m1 >>
rect 316 220 317 221 
<< m2 >>
rect 318 220 319 221 
<< m1 >>
rect 319 220 320 221 
<< m2 >>
rect 319 220 320 221 
<< m2 >>
rect 320 220 321 221 
<< m2 >>
rect 336 220 337 221 
<< m1 >>
rect 337 220 338 221 
<< m1 >>
rect 338 220 339 221 
<< m1 >>
rect 339 220 340 221 
<< m1 >>
rect 340 220 341 221 
<< m1 >>
rect 341 220 342 221 
<< m1 >>
rect 342 220 343 221 
<< m1 >>
rect 343 220 344 221 
<< m1 >>
rect 345 220 346 221 
<< m1 >>
rect 346 220 347 221 
<< m1 >>
rect 347 220 348 221 
<< m1 >>
rect 348 220 349 221 
<< m1 >>
rect 349 220 350 221 
<< m1 >>
rect 350 220 351 221 
<< m1 >>
rect 351 220 352 221 
<< m1 >>
rect 352 220 353 221 
<< m1 >>
rect 353 220 354 221 
<< m1 >>
rect 354 220 355 221 
<< m1 >>
rect 355 220 356 221 
<< m1 >>
rect 356 220 357 221 
<< m1 >>
rect 357 220 358 221 
<< m1 >>
rect 358 220 359 221 
<< m1 >>
rect 359 220 360 221 
<< m2 >>
rect 359 220 360 221 
<< m2c >>
rect 359 220 360 221 
<< m1 >>
rect 359 220 360 221 
<< m2 >>
rect 359 220 360 221 
<< m2 >>
rect 360 220 361 221 
<< m1 >>
rect 361 220 362 221 
<< m2 >>
rect 361 220 362 221 
<< m1 >>
rect 362 220 363 221 
<< m2 >>
rect 362 220 363 221 
<< m1 >>
rect 363 220 364 221 
<< m2 >>
rect 363 220 364 221 
<< m1 >>
rect 364 220 365 221 
<< m2 >>
rect 364 220 365 221 
<< m1 >>
rect 365 220 366 221 
<< m2 >>
rect 365 220 366 221 
<< m1 >>
rect 366 220 367 221 
<< m2 >>
rect 366 220 367 221 
<< m1 >>
rect 367 220 368 221 
<< m2 >>
rect 367 220 368 221 
<< m1 >>
rect 368 220 369 221 
<< m2 >>
rect 368 220 369 221 
<< m1 >>
rect 369 220 370 221 
<< m2 >>
rect 369 220 370 221 
<< m1 >>
rect 370 220 371 221 
<< m2 >>
rect 370 220 371 221 
<< m1 >>
rect 371 220 372 221 
<< m2 >>
rect 371 220 372 221 
<< m1 >>
rect 372 220 373 221 
<< m2 >>
rect 372 220 373 221 
<< m1 >>
rect 373 220 374 221 
<< m2 >>
rect 373 220 374 221 
<< m1 >>
rect 374 220 375 221 
<< m2 >>
rect 374 220 375 221 
<< m1 >>
rect 375 220 376 221 
<< m1 >>
rect 376 220 377 221 
<< m1 >>
rect 377 220 378 221 
<< m2 >>
rect 377 220 378 221 
<< m2c >>
rect 377 220 378 221 
<< m1 >>
rect 377 220 378 221 
<< m2 >>
rect 377 220 378 221 
<< m2 >>
rect 378 220 379 221 
<< m1 >>
rect 379 220 380 221 
<< m2 >>
rect 379 220 380 221 
<< m2 >>
rect 380 220 381 221 
<< m1 >>
rect 381 220 382 221 
<< m2 >>
rect 381 220 382 221 
<< m2c >>
rect 381 220 382 221 
<< m1 >>
rect 381 220 382 221 
<< m2 >>
rect 381 220 382 221 
<< m1 >>
rect 382 220 383 221 
<< m1 >>
rect 383 220 384 221 
<< m2 >>
rect 383 220 384 221 
<< m1 >>
rect 384 220 385 221 
<< m1 >>
rect 385 220 386 221 
<< m1 >>
rect 386 220 387 221 
<< m1 >>
rect 387 220 388 221 
<< m1 >>
rect 388 220 389 221 
<< m1 >>
rect 389 220 390 221 
<< m1 >>
rect 390 220 391 221 
<< m1 >>
rect 391 220 392 221 
<< m1 >>
rect 392 220 393 221 
<< m1 >>
rect 393 220 394 221 
<< m1 >>
rect 394 220 395 221 
<< m1 >>
rect 395 220 396 221 
<< m1 >>
rect 396 220 397 221 
<< m1 >>
rect 397 220 398 221 
<< m1 >>
rect 398 220 399 221 
<< m1 >>
rect 399 220 400 221 
<< m1 >>
rect 400 220 401 221 
<< m1 >>
rect 401 220 402 221 
<< m1 >>
rect 402 220 403 221 
<< m2 >>
rect 402 220 403 221 
<< m1 >>
rect 403 220 404 221 
<< m1 >>
rect 404 220 405 221 
<< m2 >>
rect 404 220 405 221 
<< m1 >>
rect 405 220 406 221 
<< m1 >>
rect 406 220 407 221 
<< m1 >>
rect 407 220 408 221 
<< m1 >>
rect 408 220 409 221 
<< m1 >>
rect 409 220 410 221 
<< m1 >>
rect 410 220 411 221 
<< m1 >>
rect 411 220 412 221 
<< m1 >>
rect 412 220 413 221 
<< m1 >>
rect 413 220 414 221 
<< m1 >>
rect 414 220 415 221 
<< m2 >>
rect 414 220 415 221 
<< m2c >>
rect 414 220 415 221 
<< m1 >>
rect 414 220 415 221 
<< m2 >>
rect 414 220 415 221 
<< m2 >>
rect 415 220 416 221 
<< m1 >>
rect 416 220 417 221 
<< m2 >>
rect 416 220 417 221 
<< m2 >>
rect 417 220 418 221 
<< m1 >>
rect 418 220 419 221 
<< m2 >>
rect 418 220 419 221 
<< m2c >>
rect 418 220 419 221 
<< m1 >>
rect 418 220 419 221 
<< m2 >>
rect 418 220 419 221 
<< m1 >>
rect 419 220 420 221 
<< m1 >>
rect 421 220 422 221 
<< m1 >>
rect 422 220 423 221 
<< m1 >>
rect 423 220 424 221 
<< m2 >>
rect 423 220 424 221 
<< m1 >>
rect 424 220 425 221 
<< m1 >>
rect 425 220 426 221 
<< m1 >>
rect 426 220 427 221 
<< m1 >>
rect 427 220 428 221 
<< m1 >>
rect 428 220 429 221 
<< m1 >>
rect 429 220 430 221 
<< m1 >>
rect 430 220 431 221 
<< m1 >>
rect 431 220 432 221 
<< m1 >>
rect 432 220 433 221 
<< m1 >>
rect 433 220 434 221 
<< m2 >>
rect 433 220 434 221 
<< m1 >>
rect 434 220 435 221 
<< m1 >>
rect 435 220 436 221 
<< m1 >>
rect 436 220 437 221 
<< m1 >>
rect 437 220 438 221 
<< m1 >>
rect 438 220 439 221 
<< m1 >>
rect 439 220 440 221 
<< m1 >>
rect 440 220 441 221 
<< m1 >>
rect 441 220 442 221 
<< m1 >>
rect 442 220 443 221 
<< m1 >>
rect 443 220 444 221 
<< m1 >>
rect 444 220 445 221 
<< m1 >>
rect 445 220 446 221 
<< m1 >>
rect 446 220 447 221 
<< m1 >>
rect 447 220 448 221 
<< m1 >>
rect 448 220 449 221 
<< m2 >>
rect 449 220 450 221 
<< m2 >>
rect 456 220 457 221 
<< m2 >>
rect 458 220 459 221 
<< m1 >>
rect 484 220 485 221 
<< m1 >>
rect 523 220 524 221 
<< m1 >>
rect 19 221 20 222 
<< m1 >>
rect 64 221 65 222 
<< m2 >>
rect 64 221 65 222 
<< m2c >>
rect 64 221 65 222 
<< m1 >>
rect 64 221 65 222 
<< m2 >>
rect 64 221 65 222 
<< m1 >>
rect 73 221 74 222 
<< m1 >>
rect 100 221 101 222 
<< m1 >>
rect 127 221 128 222 
<< m1 >>
rect 145 221 146 222 
<< m1 >>
rect 148 221 149 222 
<< m1 >>
rect 160 221 161 222 
<< m1 >>
rect 163 221 164 222 
<< m1 >>
rect 172 221 173 222 
<< m1 >>
rect 181 221 182 222 
<< m1 >>
rect 185 221 186 222 
<< m2 >>
rect 186 221 187 222 
<< m1 >>
rect 190 221 191 222 
<< m1 >>
rect 207 221 208 222 
<< m2 >>
rect 211 221 212 222 
<< m1 >>
rect 212 221 213 222 
<< m1 >>
rect 221 221 222 222 
<< m2 >>
rect 221 221 222 222 
<< m2c >>
rect 221 221 222 222 
<< m1 >>
rect 221 221 222 222 
<< m2 >>
rect 221 221 222 222 
<< m1 >>
rect 226 221 227 222 
<< m2 >>
rect 226 221 227 222 
<< m2c >>
rect 226 221 227 222 
<< m1 >>
rect 226 221 227 222 
<< m2 >>
rect 226 221 227 222 
<< m1 >>
rect 232 221 233 222 
<< m1 >>
rect 235 221 236 222 
<< m1 >>
rect 244 221 245 222 
<< m2 >>
rect 244 221 245 222 
<< m2c >>
rect 244 221 245 222 
<< m1 >>
rect 244 221 245 222 
<< m2 >>
rect 244 221 245 222 
<< m2 >>
rect 246 221 247 222 
<< m2 >>
rect 247 221 248 222 
<< m2 >>
rect 248 221 249 222 
<< m2 >>
rect 249 221 250 222 
<< m2 >>
rect 250 221 251 222 
<< m2 >>
rect 251 221 252 222 
<< m2 >>
rect 252 221 253 222 
<< m2 >>
rect 253 221 254 222 
<< m2 >>
rect 254 221 255 222 
<< m1 >>
rect 255 221 256 222 
<< m2 >>
rect 255 221 256 222 
<< m2c >>
rect 255 221 256 222 
<< m1 >>
rect 255 221 256 222 
<< m2 >>
rect 255 221 256 222 
<< m1 >>
rect 256 221 257 222 
<< m1 >>
rect 257 221 258 222 
<< m1 >>
rect 258 221 259 222 
<< m1 >>
rect 259 221 260 222 
<< m1 >>
rect 260 221 261 222 
<< m1 >>
rect 261 221 262 222 
<< m1 >>
rect 262 221 263 222 
<< m1 >>
rect 263 221 264 222 
<< m1 >>
rect 264 221 265 222 
<< m1 >>
rect 265 221 266 222 
<< m1 >>
rect 266 221 267 222 
<< m1 >>
rect 267 221 268 222 
<< m1 >>
rect 268 221 269 222 
<< m1 >>
rect 269 221 270 222 
<< m1 >>
rect 270 221 271 222 
<< m1 >>
rect 271 221 272 222 
<< m1 >>
rect 272 221 273 222 
<< m1 >>
rect 273 221 274 222 
<< m1 >>
rect 274 221 275 222 
<< m1 >>
rect 275 221 276 222 
<< m1 >>
rect 276 221 277 222 
<< m1 >>
rect 277 221 278 222 
<< m1 >>
rect 278 221 279 222 
<< m1 >>
rect 279 221 280 222 
<< m1 >>
rect 280 221 281 222 
<< m1 >>
rect 281 221 282 222 
<< m2 >>
rect 281 221 282 222 
<< m2c >>
rect 281 221 282 222 
<< m1 >>
rect 281 221 282 222 
<< m2 >>
rect 281 221 282 222 
<< m2 >>
rect 282 221 283 222 
<< m1 >>
rect 283 221 284 222 
<< m2 >>
rect 283 221 284 222 
<< m1 >>
rect 284 221 285 222 
<< m2 >>
rect 284 221 285 222 
<< m1 >>
rect 285 221 286 222 
<< m1 >>
rect 286 221 287 222 
<< m1 >>
rect 287 221 288 222 
<< m1 >>
rect 288 221 289 222 
<< m1 >>
rect 289 221 290 222 
<< m1 >>
rect 290 221 291 222 
<< m2 >>
rect 290 221 291 222 
<< m1 >>
rect 291 221 292 222 
<< m1 >>
rect 292 221 293 222 
<< m2 >>
rect 292 221 293 222 
<< m1 >>
rect 293 221 294 222 
<< m1 >>
rect 294 221 295 222 
<< m1 >>
rect 295 221 296 222 
<< m1 >>
rect 296 221 297 222 
<< m2 >>
rect 296 221 297 222 
<< m1 >>
rect 297 221 298 222 
<< m1 >>
rect 298 221 299 222 
<< m2 >>
rect 298 221 299 222 
<< m2c >>
rect 298 221 299 222 
<< m1 >>
rect 298 221 299 222 
<< m2 >>
rect 298 221 299 222 
<< m1 >>
rect 304 221 305 222 
<< m1 >>
rect 316 221 317 222 
<< m2 >>
rect 316 221 317 222 
<< m2c >>
rect 316 221 317 222 
<< m1 >>
rect 316 221 317 222 
<< m2 >>
rect 316 221 317 222 
<< m2 >>
rect 318 221 319 222 
<< m1 >>
rect 319 221 320 222 
<< m2 >>
rect 336 221 337 222 
<< m1 >>
rect 337 221 338 222 
<< m1 >>
rect 379 221 380 222 
<< m2 >>
rect 383 221 384 222 
<< m2 >>
rect 402 221 403 222 
<< m2 >>
rect 404 221 405 222 
<< m1 >>
rect 416 221 417 222 
<< m1 >>
rect 419 221 420 222 
<< m2 >>
rect 423 221 424 222 
<< m2 >>
rect 433 221 434 222 
<< m1 >>
rect 448 221 449 222 
<< m2 >>
rect 449 221 450 222 
<< m1 >>
rect 456 221 457 222 
<< m2 >>
rect 456 221 457 222 
<< m2c >>
rect 456 221 457 222 
<< m1 >>
rect 456 221 457 222 
<< m2 >>
rect 456 221 457 222 
<< m1 >>
rect 458 221 459 222 
<< m2 >>
rect 458 221 459 222 
<< m2c >>
rect 458 221 459 222 
<< m1 >>
rect 458 221 459 222 
<< m2 >>
rect 458 221 459 222 
<< m1 >>
rect 484 221 485 222 
<< m1 >>
rect 523 221 524 222 
<< m1 >>
rect 19 222 20 223 
<< m2 >>
rect 64 222 65 223 
<< m1 >>
rect 73 222 74 223 
<< m1 >>
rect 100 222 101 223 
<< m1 >>
rect 127 222 128 223 
<< m1 >>
rect 145 222 146 223 
<< m1 >>
rect 148 222 149 223 
<< m1 >>
rect 160 222 161 223 
<< m1 >>
rect 163 222 164 223 
<< m1 >>
rect 172 222 173 223 
<< m1 >>
rect 181 222 182 223 
<< m1 >>
rect 185 222 186 223 
<< m2 >>
rect 186 222 187 223 
<< m1 >>
rect 190 222 191 223 
<< m1 >>
rect 207 222 208 223 
<< m2 >>
rect 211 222 212 223 
<< m1 >>
rect 212 222 213 223 
<< m2 >>
rect 221 222 222 223 
<< m2 >>
rect 226 222 227 223 
<< m1 >>
rect 232 222 233 223 
<< m1 >>
rect 235 222 236 223 
<< m2 >>
rect 238 222 239 223 
<< m2 >>
rect 239 222 240 223 
<< m2 >>
rect 240 222 241 223 
<< m2 >>
rect 241 222 242 223 
<< m2 >>
rect 242 222 243 223 
<< m2 >>
rect 243 222 244 223 
<< m2 >>
rect 244 222 245 223 
<< m2 >>
rect 246 222 247 223 
<< m2 >>
rect 290 222 291 223 
<< m2 >>
rect 292 222 293 223 
<< m2 >>
rect 296 222 297 223 
<< m2 >>
rect 298 222 299 223 
<< m1 >>
rect 304 222 305 223 
<< m2 >>
rect 308 222 309 223 
<< m2 >>
rect 309 222 310 223 
<< m2 >>
rect 310 222 311 223 
<< m2 >>
rect 311 222 312 223 
<< m2 >>
rect 312 222 313 223 
<< m2 >>
rect 313 222 314 223 
<< m2 >>
rect 314 222 315 223 
<< m2 >>
rect 315 222 316 223 
<< m2 >>
rect 316 222 317 223 
<< m2 >>
rect 318 222 319 223 
<< m1 >>
rect 319 222 320 223 
<< m2 >>
rect 336 222 337 223 
<< m1 >>
rect 337 222 338 223 
<< m1 >>
rect 379 222 380 223 
<< m2 >>
rect 380 222 381 223 
<< m1 >>
rect 381 222 382 223 
<< m2 >>
rect 381 222 382 223 
<< m2c >>
rect 381 222 382 223 
<< m1 >>
rect 381 222 382 223 
<< m2 >>
rect 381 222 382 223 
<< m1 >>
rect 382 222 383 223 
<< m1 >>
rect 383 222 384 223 
<< m2 >>
rect 383 222 384 223 
<< m1 >>
rect 384 222 385 223 
<< m1 >>
rect 385 222 386 223 
<< m1 >>
rect 386 222 387 223 
<< m1 >>
rect 387 222 388 223 
<< m1 >>
rect 388 222 389 223 
<< m1 >>
rect 389 222 390 223 
<< m1 >>
rect 390 222 391 223 
<< m1 >>
rect 391 222 392 223 
<< m1 >>
rect 392 222 393 223 
<< m1 >>
rect 393 222 394 223 
<< m1 >>
rect 394 222 395 223 
<< m1 >>
rect 395 222 396 223 
<< m1 >>
rect 396 222 397 223 
<< m1 >>
rect 397 222 398 223 
<< m1 >>
rect 398 222 399 223 
<< m1 >>
rect 399 222 400 223 
<< m1 >>
rect 400 222 401 223 
<< m1 >>
rect 401 222 402 223 
<< m1 >>
rect 402 222 403 223 
<< m2 >>
rect 402 222 403 223 
<< m2c >>
rect 402 222 403 223 
<< m1 >>
rect 402 222 403 223 
<< m2 >>
rect 402 222 403 223 
<< m1 >>
rect 404 222 405 223 
<< m2 >>
rect 404 222 405 223 
<< m2c >>
rect 404 222 405 223 
<< m1 >>
rect 404 222 405 223 
<< m2 >>
rect 404 222 405 223 
<< m1 >>
rect 405 222 406 223 
<< m1 >>
rect 406 222 407 223 
<< m1 >>
rect 407 222 408 223 
<< m1 >>
rect 408 222 409 223 
<< m1 >>
rect 409 222 410 223 
<< m1 >>
rect 410 222 411 223 
<< m1 >>
rect 411 222 412 223 
<< m1 >>
rect 412 222 413 223 
<< m1 >>
rect 413 222 414 223 
<< m1 >>
rect 414 222 415 223 
<< m2 >>
rect 414 222 415 223 
<< m2c >>
rect 414 222 415 223 
<< m1 >>
rect 414 222 415 223 
<< m2 >>
rect 414 222 415 223 
<< m2 >>
rect 415 222 416 223 
<< m1 >>
rect 416 222 417 223 
<< m2 >>
rect 416 222 417 223 
<< m2 >>
rect 417 222 418 223 
<< m2 >>
rect 418 222 419 223 
<< m1 >>
rect 419 222 420 223 
<< m2 >>
rect 419 222 420 223 
<< m2 >>
rect 420 222 421 223 
<< m1 >>
rect 421 222 422 223 
<< m2 >>
rect 421 222 422 223 
<< m2c >>
rect 421 222 422 223 
<< m1 >>
rect 421 222 422 223 
<< m2 >>
rect 421 222 422 223 
<< m1 >>
rect 423 222 424 223 
<< m2 >>
rect 423 222 424 223 
<< m2c >>
rect 423 222 424 223 
<< m1 >>
rect 423 222 424 223 
<< m2 >>
rect 423 222 424 223 
<< m1 >>
rect 433 222 434 223 
<< m2 >>
rect 433 222 434 223 
<< m2c >>
rect 433 222 434 223 
<< m1 >>
rect 433 222 434 223 
<< m2 >>
rect 433 222 434 223 
<< m1 >>
rect 434 222 435 223 
<< m1 >>
rect 442 222 443 223 
<< m1 >>
rect 443 222 444 223 
<< m1 >>
rect 444 222 445 223 
<< m1 >>
rect 445 222 446 223 
<< m1 >>
rect 446 222 447 223 
<< m2 >>
rect 446 222 447 223 
<< m2c >>
rect 446 222 447 223 
<< m1 >>
rect 446 222 447 223 
<< m2 >>
rect 446 222 447 223 
<< m2 >>
rect 447 222 448 223 
<< m1 >>
rect 448 222 449 223 
<< m2 >>
rect 448 222 449 223 
<< m2 >>
rect 449 222 450 223 
<< m1 >>
rect 456 222 457 223 
<< m1 >>
rect 458 222 459 223 
<< m2 >>
rect 480 222 481 223 
<< m2 >>
rect 481 222 482 223 
<< m2 >>
rect 482 222 483 223 
<< m1 >>
rect 483 222 484 223 
<< m2 >>
rect 483 222 484 223 
<< m2c >>
rect 483 222 484 223 
<< m1 >>
rect 483 222 484 223 
<< m2 >>
rect 483 222 484 223 
<< m1 >>
rect 484 222 485 223 
<< m1 >>
rect 523 222 524 223 
<< m1 >>
rect 19 223 20 224 
<< m1 >>
rect 37 223 38 224 
<< m1 >>
rect 38 223 39 224 
<< m1 >>
rect 39 223 40 224 
<< m1 >>
rect 40 223 41 224 
<< m1 >>
rect 41 223 42 224 
<< m1 >>
rect 42 223 43 224 
<< m1 >>
rect 43 223 44 224 
<< m1 >>
rect 44 223 45 224 
<< m1 >>
rect 45 223 46 224 
<< m1 >>
rect 46 223 47 224 
<< m1 >>
rect 47 223 48 224 
<< m1 >>
rect 48 223 49 224 
<< m1 >>
rect 49 223 50 224 
<< m1 >>
rect 50 223 51 224 
<< m1 >>
rect 51 223 52 224 
<< m1 >>
rect 52 223 53 224 
<< m1 >>
rect 53 223 54 224 
<< m1 >>
rect 54 223 55 224 
<< m1 >>
rect 55 223 56 224 
<< m1 >>
rect 56 223 57 224 
<< m1 >>
rect 57 223 58 224 
<< m1 >>
rect 58 223 59 224 
<< m1 >>
rect 59 223 60 224 
<< m1 >>
rect 60 223 61 224 
<< m1 >>
rect 61 223 62 224 
<< m1 >>
rect 62 223 63 224 
<< m1 >>
rect 63 223 64 224 
<< m1 >>
rect 64 223 65 224 
<< m2 >>
rect 64 223 65 224 
<< m1 >>
rect 65 223 66 224 
<< m1 >>
rect 66 223 67 224 
<< m1 >>
rect 67 223 68 224 
<< m1 >>
rect 68 223 69 224 
<< m1 >>
rect 69 223 70 224 
<< m1 >>
rect 70 223 71 224 
<< m1 >>
rect 71 223 72 224 
<< m1 >>
rect 72 223 73 224 
<< m1 >>
rect 73 223 74 224 
<< m1 >>
rect 100 223 101 224 
<< m1 >>
rect 127 223 128 224 
<< m1 >>
rect 145 223 146 224 
<< m1 >>
rect 148 223 149 224 
<< m1 >>
rect 160 223 161 224 
<< m1 >>
rect 163 223 164 224 
<< m1 >>
rect 172 223 173 224 
<< m1 >>
rect 181 223 182 224 
<< m1 >>
rect 185 223 186 224 
<< m2 >>
rect 186 223 187 224 
<< m1 >>
rect 190 223 191 224 
<< m2 >>
rect 206 223 207 224 
<< m1 >>
rect 207 223 208 224 
<< m2 >>
rect 207 223 208 224 
<< m2 >>
rect 208 223 209 224 
<< m1 >>
rect 209 223 210 224 
<< m2 >>
rect 209 223 210 224 
<< m1 >>
rect 210 223 211 224 
<< m2 >>
rect 210 223 211 224 
<< m1 >>
rect 211 223 212 224 
<< m2 >>
rect 211 223 212 224 
<< m1 >>
rect 212 223 213 224 
<< m1 >>
rect 217 223 218 224 
<< m1 >>
rect 218 223 219 224 
<< m1 >>
rect 219 223 220 224 
<< m1 >>
rect 220 223 221 224 
<< m1 >>
rect 221 223 222 224 
<< m2 >>
rect 221 223 222 224 
<< m1 >>
rect 222 223 223 224 
<< m1 >>
rect 223 223 224 224 
<< m1 >>
rect 224 223 225 224 
<< m1 >>
rect 225 223 226 224 
<< m1 >>
rect 226 223 227 224 
<< m2 >>
rect 226 223 227 224 
<< m1 >>
rect 227 223 228 224 
<< m1 >>
rect 228 223 229 224 
<< m1 >>
rect 229 223 230 224 
<< m1 >>
rect 230 223 231 224 
<< m1 >>
rect 231 223 232 224 
<< m1 >>
rect 232 223 233 224 
<< m1 >>
rect 235 223 236 224 
<< m1 >>
rect 237 223 238 224 
<< m1 >>
rect 238 223 239 224 
<< m2 >>
rect 238 223 239 224 
<< m1 >>
rect 239 223 240 224 
<< m1 >>
rect 240 223 241 224 
<< m1 >>
rect 241 223 242 224 
<< m1 >>
rect 242 223 243 224 
<< m1 >>
rect 243 223 244 224 
<< m1 >>
rect 244 223 245 224 
<< m1 >>
rect 245 223 246 224 
<< m1 >>
rect 246 223 247 224 
<< m2 >>
rect 246 223 247 224 
<< m1 >>
rect 247 223 248 224 
<< m1 >>
rect 248 223 249 224 
<< m1 >>
rect 249 223 250 224 
<< m1 >>
rect 250 223 251 224 
<< m1 >>
rect 251 223 252 224 
<< m1 >>
rect 252 223 253 224 
<< m1 >>
rect 253 223 254 224 
<< m2 >>
rect 253 223 254 224 
<< m1 >>
rect 254 223 255 224 
<< m2 >>
rect 254 223 255 224 
<< m1 >>
rect 255 223 256 224 
<< m2 >>
rect 255 223 256 224 
<< m1 >>
rect 256 223 257 224 
<< m2 >>
rect 256 223 257 224 
<< m1 >>
rect 257 223 258 224 
<< m2 >>
rect 257 223 258 224 
<< m1 >>
rect 258 223 259 224 
<< m2 >>
rect 258 223 259 224 
<< m1 >>
rect 259 223 260 224 
<< m2 >>
rect 259 223 260 224 
<< m1 >>
rect 260 223 261 224 
<< m2 >>
rect 260 223 261 224 
<< m1 >>
rect 261 223 262 224 
<< m2 >>
rect 261 223 262 224 
<< m1 >>
rect 262 223 263 224 
<< m2 >>
rect 262 223 263 224 
<< m1 >>
rect 263 223 264 224 
<< m2 >>
rect 263 223 264 224 
<< m1 >>
rect 264 223 265 224 
<< m2 >>
rect 264 223 265 224 
<< m1 >>
rect 265 223 266 224 
<< m2 >>
rect 265 223 266 224 
<< m1 >>
rect 266 223 267 224 
<< m2 >>
rect 266 223 267 224 
<< m1 >>
rect 267 223 268 224 
<< m2 >>
rect 267 223 268 224 
<< m1 >>
rect 268 223 269 224 
<< m2 >>
rect 268 223 269 224 
<< m1 >>
rect 269 223 270 224 
<< m2 >>
rect 269 223 270 224 
<< m1 >>
rect 270 223 271 224 
<< m2 >>
rect 270 223 271 224 
<< m1 >>
rect 271 223 272 224 
<< m2 >>
rect 271 223 272 224 
<< m1 >>
rect 272 223 273 224 
<< m2 >>
rect 272 223 273 224 
<< m1 >>
rect 273 223 274 224 
<< m2 >>
rect 273 223 274 224 
<< m1 >>
rect 274 223 275 224 
<< m2 >>
rect 274 223 275 224 
<< m1 >>
rect 275 223 276 224 
<< m2 >>
rect 275 223 276 224 
<< m1 >>
rect 276 223 277 224 
<< m2 >>
rect 276 223 277 224 
<< m1 >>
rect 277 223 278 224 
<< m2 >>
rect 277 223 278 224 
<< m1 >>
rect 278 223 279 224 
<< m2 >>
rect 278 223 279 224 
<< m1 >>
rect 279 223 280 224 
<< m2 >>
rect 279 223 280 224 
<< m1 >>
rect 280 223 281 224 
<< m2 >>
rect 280 223 281 224 
<< m1 >>
rect 281 223 282 224 
<< m2 >>
rect 281 223 282 224 
<< m1 >>
rect 282 223 283 224 
<< m2 >>
rect 282 223 283 224 
<< m1 >>
rect 283 223 284 224 
<< m2 >>
rect 283 223 284 224 
<< m1 >>
rect 284 223 285 224 
<< m2 >>
rect 284 223 285 224 
<< m1 >>
rect 285 223 286 224 
<< m2 >>
rect 285 223 286 224 
<< m1 >>
rect 286 223 287 224 
<< m2 >>
rect 286 223 287 224 
<< m2 >>
rect 287 223 288 224 
<< m1 >>
rect 288 223 289 224 
<< m2 >>
rect 288 223 289 224 
<< m2c >>
rect 288 223 289 224 
<< m1 >>
rect 288 223 289 224 
<< m2 >>
rect 288 223 289 224 
<< m1 >>
rect 289 223 290 224 
<< m1 >>
rect 290 223 291 224 
<< m2 >>
rect 290 223 291 224 
<< m1 >>
rect 291 223 292 224 
<< m1 >>
rect 292 223 293 224 
<< m2 >>
rect 292 223 293 224 
<< m1 >>
rect 293 223 294 224 
<< m1 >>
rect 294 223 295 224 
<< m1 >>
rect 295 223 296 224 
<< m1 >>
rect 296 223 297 224 
<< m2 >>
rect 296 223 297 224 
<< m1 >>
rect 297 223 298 224 
<< m1 >>
rect 298 223 299 224 
<< m2 >>
rect 298 223 299 224 
<< m1 >>
rect 299 223 300 224 
<< m1 >>
rect 300 223 301 224 
<< m1 >>
rect 301 223 302 224 
<< m1 >>
rect 302 223 303 224 
<< m1 >>
rect 303 223 304 224 
<< m1 >>
rect 304 223 305 224 
<< m1 >>
rect 307 223 308 224 
<< m1 >>
rect 308 223 309 224 
<< m2 >>
rect 308 223 309 224 
<< m1 >>
rect 309 223 310 224 
<< m1 >>
rect 310 223 311 224 
<< m1 >>
rect 311 223 312 224 
<< m1 >>
rect 312 223 313 224 
<< m1 >>
rect 313 223 314 224 
<< m1 >>
rect 314 223 315 224 
<< m1 >>
rect 315 223 316 224 
<< m1 >>
rect 316 223 317 224 
<< m1 >>
rect 317 223 318 224 
<< m1 >>
rect 318 223 319 224 
<< m2 >>
rect 318 223 319 224 
<< m1 >>
rect 319 223 320 224 
<< m2 >>
rect 336 223 337 224 
<< m1 >>
rect 337 223 338 224 
<< m2 >>
rect 337 223 338 224 
<< m2 >>
rect 338 223 339 224 
<< m1 >>
rect 379 223 380 224 
<< m2 >>
rect 380 223 381 224 
<< m2 >>
rect 383 223 384 224 
<< m1 >>
rect 416 223 417 224 
<< m1 >>
rect 419 223 420 224 
<< m1 >>
rect 421 223 422 224 
<< m1 >>
rect 423 223 424 224 
<< m1 >>
rect 434 223 435 224 
<< m1 >>
rect 442 223 443 224 
<< m1 >>
rect 448 223 449 224 
<< m1 >>
rect 456 223 457 224 
<< m1 >>
rect 458 223 459 224 
<< m1 >>
rect 459 223 460 224 
<< m1 >>
rect 460 223 461 224 
<< m1 >>
rect 461 223 462 224 
<< m1 >>
rect 462 223 463 224 
<< m1 >>
rect 463 223 464 224 
<< m1 >>
rect 464 223 465 224 
<< m1 >>
rect 465 223 466 224 
<< m1 >>
rect 466 223 467 224 
<< m1 >>
rect 467 223 468 224 
<< m1 >>
rect 468 223 469 224 
<< m1 >>
rect 469 223 470 224 
<< m1 >>
rect 470 223 471 224 
<< m1 >>
rect 471 223 472 224 
<< m1 >>
rect 472 223 473 224 
<< m1 >>
rect 473 223 474 224 
<< m1 >>
rect 474 223 475 224 
<< m1 >>
rect 475 223 476 224 
<< m1 >>
rect 476 223 477 224 
<< m1 >>
rect 477 223 478 224 
<< m1 >>
rect 478 223 479 224 
<< m1 >>
rect 479 223 480 224 
<< m1 >>
rect 480 223 481 224 
<< m2 >>
rect 480 223 481 224 
<< m1 >>
rect 481 223 482 224 
<< m1 >>
rect 523 223 524 224 
<< m1 >>
rect 19 224 20 225 
<< m1 >>
rect 37 224 38 225 
<< m2 >>
rect 64 224 65 225 
<< m1 >>
rect 100 224 101 225 
<< m1 >>
rect 127 224 128 225 
<< m1 >>
rect 145 224 146 225 
<< m1 >>
rect 148 224 149 225 
<< m1 >>
rect 160 224 161 225 
<< m1 >>
rect 163 224 164 225 
<< m1 >>
rect 172 224 173 225 
<< m1 >>
rect 181 224 182 225 
<< m1 >>
rect 185 224 186 225 
<< m2 >>
rect 186 224 187 225 
<< m1 >>
rect 190 224 191 225 
<< m1 >>
rect 196 224 197 225 
<< m1 >>
rect 197 224 198 225 
<< m1 >>
rect 198 224 199 225 
<< m1 >>
rect 199 224 200 225 
<< m1 >>
rect 200 224 201 225 
<< m1 >>
rect 201 224 202 225 
<< m1 >>
rect 202 224 203 225 
<< m1 >>
rect 203 224 204 225 
<< m1 >>
rect 204 224 205 225 
<< m1 >>
rect 205 224 206 225 
<< m2 >>
rect 205 224 206 225 
<< m2c >>
rect 205 224 206 225 
<< m1 >>
rect 205 224 206 225 
<< m2 >>
rect 205 224 206 225 
<< m2 >>
rect 206 224 207 225 
<< m1 >>
rect 207 224 208 225 
<< m1 >>
rect 209 224 210 225 
<< m1 >>
rect 217 224 218 225 
<< m2 >>
rect 221 224 222 225 
<< m2 >>
rect 226 224 227 225 
<< m1 >>
rect 235 224 236 225 
<< m1 >>
rect 237 224 238 225 
<< m2 >>
rect 238 224 239 225 
<< m2 >>
rect 240 224 241 225 
<< m2 >>
rect 241 224 242 225 
<< m2 >>
rect 242 224 243 225 
<< m2 >>
rect 243 224 244 225 
<< m2 >>
rect 244 224 245 225 
<< m2 >>
rect 245 224 246 225 
<< m2 >>
rect 246 224 247 225 
<< m2 >>
rect 253 224 254 225 
<< m1 >>
rect 286 224 287 225 
<< m2 >>
rect 290 224 291 225 
<< m2 >>
rect 292 224 293 225 
<< m2 >>
rect 296 224 297 225 
<< m2 >>
rect 298 224 299 225 
<< m1 >>
rect 307 224 308 225 
<< m2 >>
rect 308 224 309 225 
<< m2 >>
rect 318 224 319 225 
<< m1 >>
rect 337 224 338 225 
<< m2 >>
rect 338 224 339 225 
<< m1 >>
rect 379 224 380 225 
<< m2 >>
rect 380 224 381 225 
<< m1 >>
rect 383 224 384 225 
<< m2 >>
rect 383 224 384 225 
<< m2c >>
rect 383 224 384 225 
<< m1 >>
rect 383 224 384 225 
<< m2 >>
rect 383 224 384 225 
<< m1 >>
rect 416 224 417 225 
<< m1 >>
rect 419 224 420 225 
<< m1 >>
rect 421 224 422 225 
<< m2 >>
rect 422 224 423 225 
<< m1 >>
rect 423 224 424 225 
<< m2 >>
rect 423 224 424 225 
<< m2c >>
rect 423 224 424 225 
<< m1 >>
rect 423 224 424 225 
<< m2 >>
rect 423 224 424 225 
<< m1 >>
rect 434 224 435 225 
<< m1 >>
rect 442 224 443 225 
<< m1 >>
rect 448 224 449 225 
<< m1 >>
rect 456 224 457 225 
<< m2 >>
rect 480 224 481 225 
<< m1 >>
rect 481 224 482 225 
<< m1 >>
rect 523 224 524 225 
<< m1 >>
rect 19 225 20 226 
<< m1 >>
rect 37 225 38 226 
<< m1 >>
rect 64 225 65 226 
<< m2 >>
rect 64 225 65 226 
<< m2c >>
rect 64 225 65 226 
<< m1 >>
rect 64 225 65 226 
<< m2 >>
rect 64 225 65 226 
<< m1 >>
rect 100 225 101 226 
<< m1 >>
rect 127 225 128 226 
<< m1 >>
rect 145 225 146 226 
<< m1 >>
rect 148 225 149 226 
<< m1 >>
rect 160 225 161 226 
<< m1 >>
rect 163 225 164 226 
<< m1 >>
rect 172 225 173 226 
<< m1 >>
rect 181 225 182 226 
<< m1 >>
rect 185 225 186 226 
<< m2 >>
rect 186 225 187 226 
<< m1 >>
rect 190 225 191 226 
<< m1 >>
rect 196 225 197 226 
<< m1 >>
rect 207 225 208 226 
<< m1 >>
rect 209 225 210 226 
<< m1 >>
rect 217 225 218 226 
<< m1 >>
rect 221 225 222 226 
<< m2 >>
rect 221 225 222 226 
<< m2c >>
rect 221 225 222 226 
<< m1 >>
rect 221 225 222 226 
<< m2 >>
rect 221 225 222 226 
<< m1 >>
rect 226 225 227 226 
<< m2 >>
rect 226 225 227 226 
<< m2c >>
rect 226 225 227 226 
<< m1 >>
rect 226 225 227 226 
<< m2 >>
rect 226 225 227 226 
<< m1 >>
rect 235 225 236 226 
<< m1 >>
rect 237 225 238 226 
<< m2 >>
rect 238 225 239 226 
<< m1 >>
rect 240 225 241 226 
<< m2 >>
rect 240 225 241 226 
<< m2c >>
rect 240 225 241 226 
<< m1 >>
rect 240 225 241 226 
<< m2 >>
rect 240 225 241 226 
<< m1 >>
rect 253 225 254 226 
<< m2 >>
rect 253 225 254 226 
<< m2c >>
rect 253 225 254 226 
<< m1 >>
rect 253 225 254 226 
<< m2 >>
rect 253 225 254 226 
<< m1 >>
rect 286 225 287 226 
<< m1 >>
rect 290 225 291 226 
<< m2 >>
rect 290 225 291 226 
<< m2c >>
rect 290 225 291 226 
<< m1 >>
rect 290 225 291 226 
<< m2 >>
rect 290 225 291 226 
<< m1 >>
rect 292 225 293 226 
<< m2 >>
rect 292 225 293 226 
<< m2c >>
rect 292 225 293 226 
<< m1 >>
rect 292 225 293 226 
<< m2 >>
rect 292 225 293 226 
<< m1 >>
rect 296 225 297 226 
<< m2 >>
rect 296 225 297 226 
<< m2c >>
rect 296 225 297 226 
<< m1 >>
rect 296 225 297 226 
<< m2 >>
rect 296 225 297 226 
<< m1 >>
rect 298 225 299 226 
<< m2 >>
rect 298 225 299 226 
<< m2c >>
rect 298 225 299 226 
<< m1 >>
rect 298 225 299 226 
<< m2 >>
rect 298 225 299 226 
<< m1 >>
rect 307 225 308 226 
<< m2 >>
rect 308 225 309 226 
<< m1 >>
rect 316 225 317 226 
<< m1 >>
rect 317 225 318 226 
<< m1 >>
rect 318 225 319 226 
<< m2 >>
rect 318 225 319 226 
<< m2c >>
rect 318 225 319 226 
<< m1 >>
rect 318 225 319 226 
<< m2 >>
rect 318 225 319 226 
<< m1 >>
rect 337 225 338 226 
<< m2 >>
rect 338 225 339 226 
<< m1 >>
rect 339 225 340 226 
<< m2 >>
rect 339 225 340 226 
<< m2c >>
rect 339 225 340 226 
<< m1 >>
rect 339 225 340 226 
<< m2 >>
rect 339 225 340 226 
<< m1 >>
rect 340 225 341 226 
<< m1 >>
rect 341 225 342 226 
<< m1 >>
rect 342 225 343 226 
<< m1 >>
rect 343 225 344 226 
<< m1 >>
rect 344 225 345 226 
<< m1 >>
rect 345 225 346 226 
<< m1 >>
rect 346 225 347 226 
<< m1 >>
rect 347 225 348 226 
<< m1 >>
rect 348 225 349 226 
<< m1 >>
rect 349 225 350 226 
<< m1 >>
rect 350 225 351 226 
<< m1 >>
rect 351 225 352 226 
<< m1 >>
rect 352 225 353 226 
<< m1 >>
rect 379 225 380 226 
<< m2 >>
rect 380 225 381 226 
<< m1 >>
rect 383 225 384 226 
<< m1 >>
rect 416 225 417 226 
<< m1 >>
rect 419 225 420 226 
<< m1 >>
rect 421 225 422 226 
<< m2 >>
rect 422 225 423 226 
<< m1 >>
rect 434 225 435 226 
<< m1 >>
rect 442 225 443 226 
<< m1 >>
rect 448 225 449 226 
<< m1 >>
rect 456 225 457 226 
<< m1 >>
rect 478 225 479 226 
<< m1 >>
rect 479 225 480 226 
<< m2 >>
rect 479 225 480 226 
<< m2c >>
rect 479 225 480 226 
<< m1 >>
rect 479 225 480 226 
<< m2 >>
rect 479 225 480 226 
<< m2 >>
rect 480 225 481 226 
<< m1 >>
rect 481 225 482 226 
<< m1 >>
rect 523 225 524 226 
<< m1 >>
rect 19 226 20 227 
<< m1 >>
rect 37 226 38 227 
<< m1 >>
rect 64 226 65 227 
<< m1 >>
rect 100 226 101 227 
<< m1 >>
rect 118 226 119 227 
<< m1 >>
rect 119 226 120 227 
<< m1 >>
rect 120 226 121 227 
<< m1 >>
rect 121 226 122 227 
<< m1 >>
rect 127 226 128 227 
<< m1 >>
rect 145 226 146 227 
<< m1 >>
rect 148 226 149 227 
<< m1 >>
rect 160 226 161 227 
<< m1 >>
rect 163 226 164 227 
<< m1 >>
rect 172 226 173 227 
<< m1 >>
rect 181 226 182 227 
<< m1 >>
rect 185 226 186 227 
<< m2 >>
rect 186 226 187 227 
<< m1 >>
rect 190 226 191 227 
<< m1 >>
rect 196 226 197 227 
<< m2 >>
rect 206 226 207 227 
<< m1 >>
rect 207 226 208 227 
<< m2 >>
rect 207 226 208 227 
<< m2 >>
rect 208 226 209 227 
<< m1 >>
rect 209 226 210 227 
<< m2 >>
rect 209 226 210 227 
<< m2c >>
rect 209 226 210 227 
<< m1 >>
rect 209 226 210 227 
<< m2 >>
rect 209 226 210 227 
<< m1 >>
rect 214 226 215 227 
<< m1 >>
rect 215 226 216 227 
<< m2 >>
rect 215 226 216 227 
<< m2c >>
rect 215 226 216 227 
<< m1 >>
rect 215 226 216 227 
<< m2 >>
rect 215 226 216 227 
<< m2 >>
rect 216 226 217 227 
<< m1 >>
rect 217 226 218 227 
<< m2 >>
rect 217 226 218 227 
<< m1 >>
rect 221 226 222 227 
<< m1 >>
rect 226 226 227 227 
<< m1 >>
rect 235 226 236 227 
<< m1 >>
rect 237 226 238 227 
<< m2 >>
rect 238 226 239 227 
<< m1 >>
rect 240 226 241 227 
<< m1 >>
rect 253 226 254 227 
<< m1 >>
rect 272 226 273 227 
<< m1 >>
rect 273 226 274 227 
<< m1 >>
rect 274 226 275 227 
<< m1 >>
rect 275 226 276 227 
<< m1 >>
rect 276 226 277 227 
<< m1 >>
rect 277 226 278 227 
<< m1 >>
rect 278 226 279 227 
<< m1 >>
rect 279 226 280 227 
<< m1 >>
rect 280 226 281 227 
<< m1 >>
rect 281 226 282 227 
<< m1 >>
rect 282 226 283 227 
<< m1 >>
rect 283 226 284 227 
<< m1 >>
rect 286 226 287 227 
<< m1 >>
rect 290 226 291 227 
<< m1 >>
rect 292 226 293 227 
<< m1 >>
rect 296 226 297 227 
<< m1 >>
rect 298 226 299 227 
<< m1 >>
rect 307 226 308 227 
<< m2 >>
rect 308 226 309 227 
<< m1 >>
rect 316 226 317 227 
<< m1 >>
rect 337 226 338 227 
<< m1 >>
rect 352 226 353 227 
<< m1 >>
rect 379 226 380 227 
<< m2 >>
rect 380 226 381 227 
<< m1 >>
rect 383 226 384 227 
<< m1 >>
rect 416 226 417 227 
<< m1 >>
rect 419 226 420 227 
<< m1 >>
rect 421 226 422 227 
<< m2 >>
rect 422 226 423 227 
<< m1 >>
rect 434 226 435 227 
<< m1 >>
rect 442 226 443 227 
<< m1 >>
rect 448 226 449 227 
<< m1 >>
rect 456 226 457 227 
<< m1 >>
rect 457 226 458 227 
<< m1 >>
rect 458 226 459 227 
<< m1 >>
rect 459 226 460 227 
<< m1 >>
rect 460 226 461 227 
<< m1 >>
rect 461 226 462 227 
<< m1 >>
rect 462 226 463 227 
<< m1 >>
rect 463 226 464 227 
<< m1 >>
rect 478 226 479 227 
<< m1 >>
rect 481 226 482 227 
<< m1 >>
rect 487 226 488 227 
<< m1 >>
rect 488 226 489 227 
<< m1 >>
rect 489 226 490 227 
<< m1 >>
rect 490 226 491 227 
<< m1 >>
rect 491 226 492 227 
<< m1 >>
rect 492 226 493 227 
<< m1 >>
rect 493 226 494 227 
<< m1 >>
rect 494 226 495 227 
<< m1 >>
rect 495 226 496 227 
<< m1 >>
rect 496 226 497 227 
<< m1 >>
rect 497 226 498 227 
<< m1 >>
rect 498 226 499 227 
<< m1 >>
rect 499 226 500 227 
<< m1 >>
rect 523 226 524 227 
<< m1 >>
rect 19 227 20 228 
<< m1 >>
rect 37 227 38 228 
<< m1 >>
rect 64 227 65 228 
<< m1 >>
rect 100 227 101 228 
<< m1 >>
rect 118 227 119 228 
<< m1 >>
rect 121 227 122 228 
<< m1 >>
rect 127 227 128 228 
<< m1 >>
rect 145 227 146 228 
<< m1 >>
rect 148 227 149 228 
<< m1 >>
rect 160 227 161 228 
<< m1 >>
rect 163 227 164 228 
<< m1 >>
rect 172 227 173 228 
<< m1 >>
rect 181 227 182 228 
<< m1 >>
rect 185 227 186 228 
<< m2 >>
rect 186 227 187 228 
<< m1 >>
rect 190 227 191 228 
<< m1 >>
rect 196 227 197 228 
<< m2 >>
rect 206 227 207 228 
<< m1 >>
rect 207 227 208 228 
<< m1 >>
rect 214 227 215 228 
<< m1 >>
rect 217 227 218 228 
<< m2 >>
rect 217 227 218 228 
<< m1 >>
rect 221 227 222 228 
<< m1 >>
rect 226 227 227 228 
<< m1 >>
rect 235 227 236 228 
<< m1 >>
rect 237 227 238 228 
<< m2 >>
rect 238 227 239 228 
<< m1 >>
rect 240 227 241 228 
<< m1 >>
rect 253 227 254 228 
<< m1 >>
rect 272 227 273 228 
<< m1 >>
rect 283 227 284 228 
<< m1 >>
rect 286 227 287 228 
<< m1 >>
rect 290 227 291 228 
<< m1 >>
rect 292 227 293 228 
<< m1 >>
rect 296 227 297 228 
<< m1 >>
rect 298 227 299 228 
<< m1 >>
rect 307 227 308 228 
<< m2 >>
rect 308 227 309 228 
<< m1 >>
rect 316 227 317 228 
<< m1 >>
rect 337 227 338 228 
<< m1 >>
rect 352 227 353 228 
<< m1 >>
rect 379 227 380 228 
<< m2 >>
rect 380 227 381 228 
<< m1 >>
rect 383 227 384 228 
<< m1 >>
rect 416 227 417 228 
<< m1 >>
rect 419 227 420 228 
<< m1 >>
rect 421 227 422 228 
<< m2 >>
rect 422 227 423 228 
<< m1 >>
rect 434 227 435 228 
<< m1 >>
rect 442 227 443 228 
<< m1 >>
rect 448 227 449 228 
<< m1 >>
rect 463 227 464 228 
<< m1 >>
rect 478 227 479 228 
<< m1 >>
rect 481 227 482 228 
<< m1 >>
rect 487 227 488 228 
<< m1 >>
rect 499 227 500 228 
<< m1 >>
rect 523 227 524 228 
<< pdiffusion >>
rect 12 228 13 229 
<< pdiffusion >>
rect 13 228 14 229 
<< pdiffusion >>
rect 14 228 15 229 
<< pdiffusion >>
rect 15 228 16 229 
<< pdiffusion >>
rect 16 228 17 229 
<< pdiffusion >>
rect 17 228 18 229 
<< m1 >>
rect 19 228 20 229 
<< pdiffusion >>
rect 30 228 31 229 
<< pdiffusion >>
rect 31 228 32 229 
<< pdiffusion >>
rect 32 228 33 229 
<< pdiffusion >>
rect 33 228 34 229 
<< pdiffusion >>
rect 34 228 35 229 
<< pdiffusion >>
rect 35 228 36 229 
<< m1 >>
rect 37 228 38 229 
<< pdiffusion >>
rect 48 228 49 229 
<< pdiffusion >>
rect 49 228 50 229 
<< pdiffusion >>
rect 50 228 51 229 
<< pdiffusion >>
rect 51 228 52 229 
<< pdiffusion >>
rect 52 228 53 229 
<< pdiffusion >>
rect 53 228 54 229 
<< m1 >>
rect 64 228 65 229 
<< pdiffusion >>
rect 66 228 67 229 
<< pdiffusion >>
rect 67 228 68 229 
<< pdiffusion >>
rect 68 228 69 229 
<< pdiffusion >>
rect 69 228 70 229 
<< pdiffusion >>
rect 70 228 71 229 
<< pdiffusion >>
rect 71 228 72 229 
<< pdiffusion >>
rect 84 228 85 229 
<< pdiffusion >>
rect 85 228 86 229 
<< pdiffusion >>
rect 86 228 87 229 
<< pdiffusion >>
rect 87 228 88 229 
<< pdiffusion >>
rect 88 228 89 229 
<< pdiffusion >>
rect 89 228 90 229 
<< m1 >>
rect 100 228 101 229 
<< pdiffusion >>
rect 102 228 103 229 
<< pdiffusion >>
rect 103 228 104 229 
<< pdiffusion >>
rect 104 228 105 229 
<< pdiffusion >>
rect 105 228 106 229 
<< pdiffusion >>
rect 106 228 107 229 
<< pdiffusion >>
rect 107 228 108 229 
<< m1 >>
rect 118 228 119 229 
<< pdiffusion >>
rect 120 228 121 229 
<< m1 >>
rect 121 228 122 229 
<< pdiffusion >>
rect 121 228 122 229 
<< pdiffusion >>
rect 122 228 123 229 
<< pdiffusion >>
rect 123 228 124 229 
<< pdiffusion >>
rect 124 228 125 229 
<< pdiffusion >>
rect 125 228 126 229 
<< m1 >>
rect 127 228 128 229 
<< pdiffusion >>
rect 138 228 139 229 
<< pdiffusion >>
rect 139 228 140 229 
<< pdiffusion >>
rect 140 228 141 229 
<< pdiffusion >>
rect 141 228 142 229 
<< pdiffusion >>
rect 142 228 143 229 
<< pdiffusion >>
rect 143 228 144 229 
<< m1 >>
rect 145 228 146 229 
<< m1 >>
rect 148 228 149 229 
<< pdiffusion >>
rect 156 228 157 229 
<< pdiffusion >>
rect 157 228 158 229 
<< pdiffusion >>
rect 158 228 159 229 
<< pdiffusion >>
rect 159 228 160 229 
<< m1 >>
rect 160 228 161 229 
<< pdiffusion >>
rect 160 228 161 229 
<< pdiffusion >>
rect 161 228 162 229 
<< m1 >>
rect 163 228 164 229 
<< m1 >>
rect 172 228 173 229 
<< pdiffusion >>
rect 174 228 175 229 
<< pdiffusion >>
rect 175 228 176 229 
<< pdiffusion >>
rect 176 228 177 229 
<< pdiffusion >>
rect 177 228 178 229 
<< pdiffusion >>
rect 178 228 179 229 
<< pdiffusion >>
rect 179 228 180 229 
<< m1 >>
rect 181 228 182 229 
<< m1 >>
rect 185 228 186 229 
<< m2 >>
rect 186 228 187 229 
<< m1 >>
rect 190 228 191 229 
<< pdiffusion >>
rect 192 228 193 229 
<< pdiffusion >>
rect 193 228 194 229 
<< pdiffusion >>
rect 194 228 195 229 
<< pdiffusion >>
rect 195 228 196 229 
<< m1 >>
rect 196 228 197 229 
<< pdiffusion >>
rect 196 228 197 229 
<< pdiffusion >>
rect 197 228 198 229 
<< m2 >>
rect 206 228 207 229 
<< m1 >>
rect 207 228 208 229 
<< pdiffusion >>
rect 210 228 211 229 
<< pdiffusion >>
rect 211 228 212 229 
<< pdiffusion >>
rect 212 228 213 229 
<< pdiffusion >>
rect 213 228 214 229 
<< m1 >>
rect 214 228 215 229 
<< pdiffusion >>
rect 214 228 215 229 
<< pdiffusion >>
rect 215 228 216 229 
<< m1 >>
rect 217 228 218 229 
<< m2 >>
rect 217 228 218 229 
<< m1 >>
rect 221 228 222 229 
<< m1 >>
rect 226 228 227 229 
<< pdiffusion >>
rect 228 228 229 229 
<< pdiffusion >>
rect 229 228 230 229 
<< pdiffusion >>
rect 230 228 231 229 
<< pdiffusion >>
rect 231 228 232 229 
<< pdiffusion >>
rect 232 228 233 229 
<< pdiffusion >>
rect 233 228 234 229 
<< m1 >>
rect 235 228 236 229 
<< m1 >>
rect 237 228 238 229 
<< m2 >>
rect 238 228 239 229 
<< m1 >>
rect 240 228 241 229 
<< pdiffusion >>
rect 246 228 247 229 
<< pdiffusion >>
rect 247 228 248 229 
<< pdiffusion >>
rect 248 228 249 229 
<< pdiffusion >>
rect 249 228 250 229 
<< pdiffusion >>
rect 250 228 251 229 
<< pdiffusion >>
rect 251 228 252 229 
<< m1 >>
rect 253 228 254 229 
<< pdiffusion >>
rect 264 228 265 229 
<< pdiffusion >>
rect 265 228 266 229 
<< pdiffusion >>
rect 266 228 267 229 
<< pdiffusion >>
rect 267 228 268 229 
<< pdiffusion >>
rect 268 228 269 229 
<< pdiffusion >>
rect 269 228 270 229 
<< m1 >>
rect 272 228 273 229 
<< pdiffusion >>
rect 282 228 283 229 
<< m1 >>
rect 283 228 284 229 
<< pdiffusion >>
rect 283 228 284 229 
<< pdiffusion >>
rect 284 228 285 229 
<< pdiffusion >>
rect 285 228 286 229 
<< m1 >>
rect 286 228 287 229 
<< pdiffusion >>
rect 286 228 287 229 
<< pdiffusion >>
rect 287 228 288 229 
<< m1 >>
rect 290 228 291 229 
<< m1 >>
rect 292 228 293 229 
<< m1 >>
rect 296 228 297 229 
<< m1 >>
rect 298 228 299 229 
<< pdiffusion >>
rect 300 228 301 229 
<< pdiffusion >>
rect 301 228 302 229 
<< pdiffusion >>
rect 302 228 303 229 
<< pdiffusion >>
rect 303 228 304 229 
<< pdiffusion >>
rect 304 228 305 229 
<< pdiffusion >>
rect 305 228 306 229 
<< m1 >>
rect 307 228 308 229 
<< m2 >>
rect 308 228 309 229 
<< m1 >>
rect 316 228 317 229 
<< pdiffusion >>
rect 318 228 319 229 
<< pdiffusion >>
rect 319 228 320 229 
<< pdiffusion >>
rect 320 228 321 229 
<< pdiffusion >>
rect 321 228 322 229 
<< pdiffusion >>
rect 322 228 323 229 
<< pdiffusion >>
rect 323 228 324 229 
<< pdiffusion >>
rect 336 228 337 229 
<< m1 >>
rect 337 228 338 229 
<< pdiffusion >>
rect 337 228 338 229 
<< pdiffusion >>
rect 338 228 339 229 
<< pdiffusion >>
rect 339 228 340 229 
<< pdiffusion >>
rect 340 228 341 229 
<< pdiffusion >>
rect 341 228 342 229 
<< m1 >>
rect 352 228 353 229 
<< pdiffusion >>
rect 354 228 355 229 
<< pdiffusion >>
rect 355 228 356 229 
<< pdiffusion >>
rect 356 228 357 229 
<< pdiffusion >>
rect 357 228 358 229 
<< pdiffusion >>
rect 358 228 359 229 
<< pdiffusion >>
rect 359 228 360 229 
<< pdiffusion >>
rect 372 228 373 229 
<< pdiffusion >>
rect 373 228 374 229 
<< pdiffusion >>
rect 374 228 375 229 
<< pdiffusion >>
rect 375 228 376 229 
<< pdiffusion >>
rect 376 228 377 229 
<< pdiffusion >>
rect 377 228 378 229 
<< m1 >>
rect 379 228 380 229 
<< m2 >>
rect 380 228 381 229 
<< m1 >>
rect 383 228 384 229 
<< pdiffusion >>
rect 390 228 391 229 
<< pdiffusion >>
rect 391 228 392 229 
<< pdiffusion >>
rect 392 228 393 229 
<< pdiffusion >>
rect 393 228 394 229 
<< pdiffusion >>
rect 394 228 395 229 
<< pdiffusion >>
rect 395 228 396 229 
<< pdiffusion >>
rect 408 228 409 229 
<< pdiffusion >>
rect 409 228 410 229 
<< pdiffusion >>
rect 410 228 411 229 
<< pdiffusion >>
rect 411 228 412 229 
<< pdiffusion >>
rect 412 228 413 229 
<< pdiffusion >>
rect 413 228 414 229 
<< m1 >>
rect 416 228 417 229 
<< m1 >>
rect 419 228 420 229 
<< m1 >>
rect 421 228 422 229 
<< m2 >>
rect 422 228 423 229 
<< pdiffusion >>
rect 426 228 427 229 
<< pdiffusion >>
rect 427 228 428 229 
<< pdiffusion >>
rect 428 228 429 229 
<< pdiffusion >>
rect 429 228 430 229 
<< pdiffusion >>
rect 430 228 431 229 
<< pdiffusion >>
rect 431 228 432 229 
<< m1 >>
rect 434 228 435 229 
<< m1 >>
rect 442 228 443 229 
<< pdiffusion >>
rect 444 228 445 229 
<< pdiffusion >>
rect 445 228 446 229 
<< pdiffusion >>
rect 446 228 447 229 
<< pdiffusion >>
rect 447 228 448 229 
<< m1 >>
rect 448 228 449 229 
<< pdiffusion >>
rect 448 228 449 229 
<< pdiffusion >>
rect 449 228 450 229 
<< pdiffusion >>
rect 462 228 463 229 
<< m1 >>
rect 463 228 464 229 
<< pdiffusion >>
rect 463 228 464 229 
<< pdiffusion >>
rect 464 228 465 229 
<< pdiffusion >>
rect 465 228 466 229 
<< pdiffusion >>
rect 466 228 467 229 
<< pdiffusion >>
rect 467 228 468 229 
<< m1 >>
rect 478 228 479 229 
<< pdiffusion >>
rect 480 228 481 229 
<< m1 >>
rect 481 228 482 229 
<< pdiffusion >>
rect 481 228 482 229 
<< pdiffusion >>
rect 482 228 483 229 
<< pdiffusion >>
rect 483 228 484 229 
<< pdiffusion >>
rect 484 228 485 229 
<< pdiffusion >>
rect 485 228 486 229 
<< m1 >>
rect 487 228 488 229 
<< pdiffusion >>
rect 498 228 499 229 
<< m1 >>
rect 499 228 500 229 
<< pdiffusion >>
rect 499 228 500 229 
<< pdiffusion >>
rect 500 228 501 229 
<< pdiffusion >>
rect 501 228 502 229 
<< pdiffusion >>
rect 502 228 503 229 
<< pdiffusion >>
rect 503 228 504 229 
<< m1 >>
rect 523 228 524 229 
<< pdiffusion >>
rect 12 229 13 230 
<< pdiffusion >>
rect 13 229 14 230 
<< pdiffusion >>
rect 14 229 15 230 
<< pdiffusion >>
rect 15 229 16 230 
<< pdiffusion >>
rect 16 229 17 230 
<< pdiffusion >>
rect 17 229 18 230 
<< m1 >>
rect 19 229 20 230 
<< pdiffusion >>
rect 30 229 31 230 
<< pdiffusion >>
rect 31 229 32 230 
<< pdiffusion >>
rect 32 229 33 230 
<< pdiffusion >>
rect 33 229 34 230 
<< pdiffusion >>
rect 34 229 35 230 
<< pdiffusion >>
rect 35 229 36 230 
<< m1 >>
rect 37 229 38 230 
<< pdiffusion >>
rect 48 229 49 230 
<< pdiffusion >>
rect 49 229 50 230 
<< pdiffusion >>
rect 50 229 51 230 
<< pdiffusion >>
rect 51 229 52 230 
<< pdiffusion >>
rect 52 229 53 230 
<< pdiffusion >>
rect 53 229 54 230 
<< m1 >>
rect 64 229 65 230 
<< pdiffusion >>
rect 66 229 67 230 
<< pdiffusion >>
rect 67 229 68 230 
<< pdiffusion >>
rect 68 229 69 230 
<< pdiffusion >>
rect 69 229 70 230 
<< pdiffusion >>
rect 70 229 71 230 
<< pdiffusion >>
rect 71 229 72 230 
<< pdiffusion >>
rect 84 229 85 230 
<< pdiffusion >>
rect 85 229 86 230 
<< pdiffusion >>
rect 86 229 87 230 
<< pdiffusion >>
rect 87 229 88 230 
<< pdiffusion >>
rect 88 229 89 230 
<< pdiffusion >>
rect 89 229 90 230 
<< m1 >>
rect 100 229 101 230 
<< pdiffusion >>
rect 102 229 103 230 
<< pdiffusion >>
rect 103 229 104 230 
<< pdiffusion >>
rect 104 229 105 230 
<< pdiffusion >>
rect 105 229 106 230 
<< pdiffusion >>
rect 106 229 107 230 
<< pdiffusion >>
rect 107 229 108 230 
<< m1 >>
rect 118 229 119 230 
<< pdiffusion >>
rect 120 229 121 230 
<< pdiffusion >>
rect 121 229 122 230 
<< pdiffusion >>
rect 122 229 123 230 
<< pdiffusion >>
rect 123 229 124 230 
<< pdiffusion >>
rect 124 229 125 230 
<< pdiffusion >>
rect 125 229 126 230 
<< m1 >>
rect 127 229 128 230 
<< pdiffusion >>
rect 138 229 139 230 
<< pdiffusion >>
rect 139 229 140 230 
<< pdiffusion >>
rect 140 229 141 230 
<< pdiffusion >>
rect 141 229 142 230 
<< pdiffusion >>
rect 142 229 143 230 
<< pdiffusion >>
rect 143 229 144 230 
<< m1 >>
rect 145 229 146 230 
<< m1 >>
rect 148 229 149 230 
<< pdiffusion >>
rect 156 229 157 230 
<< pdiffusion >>
rect 157 229 158 230 
<< pdiffusion >>
rect 158 229 159 230 
<< pdiffusion >>
rect 159 229 160 230 
<< pdiffusion >>
rect 160 229 161 230 
<< pdiffusion >>
rect 161 229 162 230 
<< m1 >>
rect 163 229 164 230 
<< m1 >>
rect 172 229 173 230 
<< pdiffusion >>
rect 174 229 175 230 
<< pdiffusion >>
rect 175 229 176 230 
<< pdiffusion >>
rect 176 229 177 230 
<< pdiffusion >>
rect 177 229 178 230 
<< pdiffusion >>
rect 178 229 179 230 
<< pdiffusion >>
rect 179 229 180 230 
<< m1 >>
rect 181 229 182 230 
<< m1 >>
rect 185 229 186 230 
<< m2 >>
rect 186 229 187 230 
<< m1 >>
rect 190 229 191 230 
<< pdiffusion >>
rect 192 229 193 230 
<< pdiffusion >>
rect 193 229 194 230 
<< pdiffusion >>
rect 194 229 195 230 
<< pdiffusion >>
rect 195 229 196 230 
<< pdiffusion >>
rect 196 229 197 230 
<< pdiffusion >>
rect 197 229 198 230 
<< m2 >>
rect 206 229 207 230 
<< m1 >>
rect 207 229 208 230 
<< pdiffusion >>
rect 210 229 211 230 
<< pdiffusion >>
rect 211 229 212 230 
<< pdiffusion >>
rect 212 229 213 230 
<< pdiffusion >>
rect 213 229 214 230 
<< pdiffusion >>
rect 214 229 215 230 
<< pdiffusion >>
rect 215 229 216 230 
<< m1 >>
rect 217 229 218 230 
<< m2 >>
rect 217 229 218 230 
<< m1 >>
rect 221 229 222 230 
<< m1 >>
rect 226 229 227 230 
<< pdiffusion >>
rect 228 229 229 230 
<< pdiffusion >>
rect 229 229 230 230 
<< pdiffusion >>
rect 230 229 231 230 
<< pdiffusion >>
rect 231 229 232 230 
<< pdiffusion >>
rect 232 229 233 230 
<< pdiffusion >>
rect 233 229 234 230 
<< m1 >>
rect 235 229 236 230 
<< m1 >>
rect 237 229 238 230 
<< m2 >>
rect 238 229 239 230 
<< m1 >>
rect 240 229 241 230 
<< pdiffusion >>
rect 246 229 247 230 
<< pdiffusion >>
rect 247 229 248 230 
<< pdiffusion >>
rect 248 229 249 230 
<< pdiffusion >>
rect 249 229 250 230 
<< pdiffusion >>
rect 250 229 251 230 
<< pdiffusion >>
rect 251 229 252 230 
<< m1 >>
rect 253 229 254 230 
<< pdiffusion >>
rect 264 229 265 230 
<< pdiffusion >>
rect 265 229 266 230 
<< pdiffusion >>
rect 266 229 267 230 
<< pdiffusion >>
rect 267 229 268 230 
<< pdiffusion >>
rect 268 229 269 230 
<< pdiffusion >>
rect 269 229 270 230 
<< m1 >>
rect 272 229 273 230 
<< pdiffusion >>
rect 282 229 283 230 
<< pdiffusion >>
rect 283 229 284 230 
<< pdiffusion >>
rect 284 229 285 230 
<< pdiffusion >>
rect 285 229 286 230 
<< pdiffusion >>
rect 286 229 287 230 
<< pdiffusion >>
rect 287 229 288 230 
<< m1 >>
rect 290 229 291 230 
<< m1 >>
rect 292 229 293 230 
<< m1 >>
rect 296 229 297 230 
<< m1 >>
rect 298 229 299 230 
<< pdiffusion >>
rect 300 229 301 230 
<< pdiffusion >>
rect 301 229 302 230 
<< pdiffusion >>
rect 302 229 303 230 
<< pdiffusion >>
rect 303 229 304 230 
<< pdiffusion >>
rect 304 229 305 230 
<< pdiffusion >>
rect 305 229 306 230 
<< m1 >>
rect 307 229 308 230 
<< m2 >>
rect 308 229 309 230 
<< m1 >>
rect 316 229 317 230 
<< pdiffusion >>
rect 318 229 319 230 
<< pdiffusion >>
rect 319 229 320 230 
<< pdiffusion >>
rect 320 229 321 230 
<< pdiffusion >>
rect 321 229 322 230 
<< pdiffusion >>
rect 322 229 323 230 
<< pdiffusion >>
rect 323 229 324 230 
<< pdiffusion >>
rect 336 229 337 230 
<< pdiffusion >>
rect 337 229 338 230 
<< pdiffusion >>
rect 338 229 339 230 
<< pdiffusion >>
rect 339 229 340 230 
<< pdiffusion >>
rect 340 229 341 230 
<< pdiffusion >>
rect 341 229 342 230 
<< m1 >>
rect 352 229 353 230 
<< pdiffusion >>
rect 354 229 355 230 
<< pdiffusion >>
rect 355 229 356 230 
<< pdiffusion >>
rect 356 229 357 230 
<< pdiffusion >>
rect 357 229 358 230 
<< pdiffusion >>
rect 358 229 359 230 
<< pdiffusion >>
rect 359 229 360 230 
<< pdiffusion >>
rect 372 229 373 230 
<< pdiffusion >>
rect 373 229 374 230 
<< pdiffusion >>
rect 374 229 375 230 
<< pdiffusion >>
rect 375 229 376 230 
<< pdiffusion >>
rect 376 229 377 230 
<< pdiffusion >>
rect 377 229 378 230 
<< m1 >>
rect 379 229 380 230 
<< m2 >>
rect 380 229 381 230 
<< m1 >>
rect 383 229 384 230 
<< pdiffusion >>
rect 390 229 391 230 
<< pdiffusion >>
rect 391 229 392 230 
<< pdiffusion >>
rect 392 229 393 230 
<< pdiffusion >>
rect 393 229 394 230 
<< pdiffusion >>
rect 394 229 395 230 
<< pdiffusion >>
rect 395 229 396 230 
<< pdiffusion >>
rect 408 229 409 230 
<< pdiffusion >>
rect 409 229 410 230 
<< pdiffusion >>
rect 410 229 411 230 
<< pdiffusion >>
rect 411 229 412 230 
<< pdiffusion >>
rect 412 229 413 230 
<< pdiffusion >>
rect 413 229 414 230 
<< m1 >>
rect 416 229 417 230 
<< m1 >>
rect 419 229 420 230 
<< m1 >>
rect 421 229 422 230 
<< m2 >>
rect 422 229 423 230 
<< pdiffusion >>
rect 426 229 427 230 
<< pdiffusion >>
rect 427 229 428 230 
<< pdiffusion >>
rect 428 229 429 230 
<< pdiffusion >>
rect 429 229 430 230 
<< pdiffusion >>
rect 430 229 431 230 
<< pdiffusion >>
rect 431 229 432 230 
<< m1 >>
rect 434 229 435 230 
<< m1 >>
rect 442 229 443 230 
<< pdiffusion >>
rect 444 229 445 230 
<< pdiffusion >>
rect 445 229 446 230 
<< pdiffusion >>
rect 446 229 447 230 
<< pdiffusion >>
rect 447 229 448 230 
<< pdiffusion >>
rect 448 229 449 230 
<< pdiffusion >>
rect 449 229 450 230 
<< pdiffusion >>
rect 462 229 463 230 
<< pdiffusion >>
rect 463 229 464 230 
<< pdiffusion >>
rect 464 229 465 230 
<< pdiffusion >>
rect 465 229 466 230 
<< pdiffusion >>
rect 466 229 467 230 
<< pdiffusion >>
rect 467 229 468 230 
<< m1 >>
rect 478 229 479 230 
<< pdiffusion >>
rect 480 229 481 230 
<< pdiffusion >>
rect 481 229 482 230 
<< pdiffusion >>
rect 482 229 483 230 
<< pdiffusion >>
rect 483 229 484 230 
<< pdiffusion >>
rect 484 229 485 230 
<< pdiffusion >>
rect 485 229 486 230 
<< m1 >>
rect 487 229 488 230 
<< pdiffusion >>
rect 498 229 499 230 
<< pdiffusion >>
rect 499 229 500 230 
<< pdiffusion >>
rect 500 229 501 230 
<< pdiffusion >>
rect 501 229 502 230 
<< pdiffusion >>
rect 502 229 503 230 
<< pdiffusion >>
rect 503 229 504 230 
<< m1 >>
rect 523 229 524 230 
<< pdiffusion >>
rect 12 230 13 231 
<< pdiffusion >>
rect 13 230 14 231 
<< pdiffusion >>
rect 14 230 15 231 
<< pdiffusion >>
rect 15 230 16 231 
<< pdiffusion >>
rect 16 230 17 231 
<< pdiffusion >>
rect 17 230 18 231 
<< m1 >>
rect 19 230 20 231 
<< pdiffusion >>
rect 30 230 31 231 
<< pdiffusion >>
rect 31 230 32 231 
<< pdiffusion >>
rect 32 230 33 231 
<< pdiffusion >>
rect 33 230 34 231 
<< pdiffusion >>
rect 34 230 35 231 
<< pdiffusion >>
rect 35 230 36 231 
<< m1 >>
rect 37 230 38 231 
<< pdiffusion >>
rect 48 230 49 231 
<< pdiffusion >>
rect 49 230 50 231 
<< pdiffusion >>
rect 50 230 51 231 
<< pdiffusion >>
rect 51 230 52 231 
<< pdiffusion >>
rect 52 230 53 231 
<< pdiffusion >>
rect 53 230 54 231 
<< m1 >>
rect 64 230 65 231 
<< pdiffusion >>
rect 66 230 67 231 
<< pdiffusion >>
rect 67 230 68 231 
<< pdiffusion >>
rect 68 230 69 231 
<< pdiffusion >>
rect 69 230 70 231 
<< pdiffusion >>
rect 70 230 71 231 
<< pdiffusion >>
rect 71 230 72 231 
<< pdiffusion >>
rect 84 230 85 231 
<< pdiffusion >>
rect 85 230 86 231 
<< pdiffusion >>
rect 86 230 87 231 
<< pdiffusion >>
rect 87 230 88 231 
<< pdiffusion >>
rect 88 230 89 231 
<< pdiffusion >>
rect 89 230 90 231 
<< m1 >>
rect 100 230 101 231 
<< pdiffusion >>
rect 102 230 103 231 
<< pdiffusion >>
rect 103 230 104 231 
<< pdiffusion >>
rect 104 230 105 231 
<< pdiffusion >>
rect 105 230 106 231 
<< pdiffusion >>
rect 106 230 107 231 
<< pdiffusion >>
rect 107 230 108 231 
<< m1 >>
rect 118 230 119 231 
<< pdiffusion >>
rect 120 230 121 231 
<< pdiffusion >>
rect 121 230 122 231 
<< pdiffusion >>
rect 122 230 123 231 
<< pdiffusion >>
rect 123 230 124 231 
<< pdiffusion >>
rect 124 230 125 231 
<< pdiffusion >>
rect 125 230 126 231 
<< m1 >>
rect 127 230 128 231 
<< pdiffusion >>
rect 138 230 139 231 
<< pdiffusion >>
rect 139 230 140 231 
<< pdiffusion >>
rect 140 230 141 231 
<< pdiffusion >>
rect 141 230 142 231 
<< pdiffusion >>
rect 142 230 143 231 
<< pdiffusion >>
rect 143 230 144 231 
<< m1 >>
rect 145 230 146 231 
<< m1 >>
rect 148 230 149 231 
<< pdiffusion >>
rect 156 230 157 231 
<< pdiffusion >>
rect 157 230 158 231 
<< pdiffusion >>
rect 158 230 159 231 
<< pdiffusion >>
rect 159 230 160 231 
<< pdiffusion >>
rect 160 230 161 231 
<< pdiffusion >>
rect 161 230 162 231 
<< m1 >>
rect 163 230 164 231 
<< m1 >>
rect 172 230 173 231 
<< pdiffusion >>
rect 174 230 175 231 
<< pdiffusion >>
rect 175 230 176 231 
<< pdiffusion >>
rect 176 230 177 231 
<< pdiffusion >>
rect 177 230 178 231 
<< pdiffusion >>
rect 178 230 179 231 
<< pdiffusion >>
rect 179 230 180 231 
<< m1 >>
rect 181 230 182 231 
<< m1 >>
rect 185 230 186 231 
<< m2 >>
rect 186 230 187 231 
<< m1 >>
rect 190 230 191 231 
<< pdiffusion >>
rect 192 230 193 231 
<< pdiffusion >>
rect 193 230 194 231 
<< pdiffusion >>
rect 194 230 195 231 
<< pdiffusion >>
rect 195 230 196 231 
<< pdiffusion >>
rect 196 230 197 231 
<< pdiffusion >>
rect 197 230 198 231 
<< m2 >>
rect 206 230 207 231 
<< m1 >>
rect 207 230 208 231 
<< pdiffusion >>
rect 210 230 211 231 
<< pdiffusion >>
rect 211 230 212 231 
<< pdiffusion >>
rect 212 230 213 231 
<< pdiffusion >>
rect 213 230 214 231 
<< pdiffusion >>
rect 214 230 215 231 
<< pdiffusion >>
rect 215 230 216 231 
<< m1 >>
rect 217 230 218 231 
<< m2 >>
rect 217 230 218 231 
<< m1 >>
rect 221 230 222 231 
<< m1 >>
rect 226 230 227 231 
<< pdiffusion >>
rect 228 230 229 231 
<< pdiffusion >>
rect 229 230 230 231 
<< pdiffusion >>
rect 230 230 231 231 
<< pdiffusion >>
rect 231 230 232 231 
<< pdiffusion >>
rect 232 230 233 231 
<< pdiffusion >>
rect 233 230 234 231 
<< m1 >>
rect 235 230 236 231 
<< m1 >>
rect 237 230 238 231 
<< m2 >>
rect 238 230 239 231 
<< m1 >>
rect 240 230 241 231 
<< pdiffusion >>
rect 246 230 247 231 
<< pdiffusion >>
rect 247 230 248 231 
<< pdiffusion >>
rect 248 230 249 231 
<< pdiffusion >>
rect 249 230 250 231 
<< pdiffusion >>
rect 250 230 251 231 
<< pdiffusion >>
rect 251 230 252 231 
<< m1 >>
rect 253 230 254 231 
<< pdiffusion >>
rect 264 230 265 231 
<< pdiffusion >>
rect 265 230 266 231 
<< pdiffusion >>
rect 266 230 267 231 
<< pdiffusion >>
rect 267 230 268 231 
<< pdiffusion >>
rect 268 230 269 231 
<< pdiffusion >>
rect 269 230 270 231 
<< m1 >>
rect 272 230 273 231 
<< pdiffusion >>
rect 282 230 283 231 
<< pdiffusion >>
rect 283 230 284 231 
<< pdiffusion >>
rect 284 230 285 231 
<< pdiffusion >>
rect 285 230 286 231 
<< pdiffusion >>
rect 286 230 287 231 
<< pdiffusion >>
rect 287 230 288 231 
<< m1 >>
rect 290 230 291 231 
<< m1 >>
rect 292 230 293 231 
<< m1 >>
rect 296 230 297 231 
<< m1 >>
rect 298 230 299 231 
<< pdiffusion >>
rect 300 230 301 231 
<< pdiffusion >>
rect 301 230 302 231 
<< pdiffusion >>
rect 302 230 303 231 
<< pdiffusion >>
rect 303 230 304 231 
<< pdiffusion >>
rect 304 230 305 231 
<< pdiffusion >>
rect 305 230 306 231 
<< m1 >>
rect 307 230 308 231 
<< m2 >>
rect 308 230 309 231 
<< m1 >>
rect 316 230 317 231 
<< pdiffusion >>
rect 318 230 319 231 
<< pdiffusion >>
rect 319 230 320 231 
<< pdiffusion >>
rect 320 230 321 231 
<< pdiffusion >>
rect 321 230 322 231 
<< pdiffusion >>
rect 322 230 323 231 
<< pdiffusion >>
rect 323 230 324 231 
<< pdiffusion >>
rect 336 230 337 231 
<< pdiffusion >>
rect 337 230 338 231 
<< pdiffusion >>
rect 338 230 339 231 
<< pdiffusion >>
rect 339 230 340 231 
<< pdiffusion >>
rect 340 230 341 231 
<< pdiffusion >>
rect 341 230 342 231 
<< m1 >>
rect 352 230 353 231 
<< pdiffusion >>
rect 354 230 355 231 
<< pdiffusion >>
rect 355 230 356 231 
<< pdiffusion >>
rect 356 230 357 231 
<< pdiffusion >>
rect 357 230 358 231 
<< pdiffusion >>
rect 358 230 359 231 
<< pdiffusion >>
rect 359 230 360 231 
<< pdiffusion >>
rect 372 230 373 231 
<< pdiffusion >>
rect 373 230 374 231 
<< pdiffusion >>
rect 374 230 375 231 
<< pdiffusion >>
rect 375 230 376 231 
<< pdiffusion >>
rect 376 230 377 231 
<< pdiffusion >>
rect 377 230 378 231 
<< m1 >>
rect 379 230 380 231 
<< m2 >>
rect 380 230 381 231 
<< m1 >>
rect 383 230 384 231 
<< pdiffusion >>
rect 390 230 391 231 
<< pdiffusion >>
rect 391 230 392 231 
<< pdiffusion >>
rect 392 230 393 231 
<< pdiffusion >>
rect 393 230 394 231 
<< pdiffusion >>
rect 394 230 395 231 
<< pdiffusion >>
rect 395 230 396 231 
<< pdiffusion >>
rect 408 230 409 231 
<< pdiffusion >>
rect 409 230 410 231 
<< pdiffusion >>
rect 410 230 411 231 
<< pdiffusion >>
rect 411 230 412 231 
<< pdiffusion >>
rect 412 230 413 231 
<< pdiffusion >>
rect 413 230 414 231 
<< m1 >>
rect 416 230 417 231 
<< m1 >>
rect 419 230 420 231 
<< m1 >>
rect 421 230 422 231 
<< m2 >>
rect 422 230 423 231 
<< pdiffusion >>
rect 426 230 427 231 
<< pdiffusion >>
rect 427 230 428 231 
<< pdiffusion >>
rect 428 230 429 231 
<< pdiffusion >>
rect 429 230 430 231 
<< pdiffusion >>
rect 430 230 431 231 
<< pdiffusion >>
rect 431 230 432 231 
<< m1 >>
rect 434 230 435 231 
<< m1 >>
rect 442 230 443 231 
<< pdiffusion >>
rect 444 230 445 231 
<< pdiffusion >>
rect 445 230 446 231 
<< pdiffusion >>
rect 446 230 447 231 
<< pdiffusion >>
rect 447 230 448 231 
<< pdiffusion >>
rect 448 230 449 231 
<< pdiffusion >>
rect 449 230 450 231 
<< pdiffusion >>
rect 462 230 463 231 
<< pdiffusion >>
rect 463 230 464 231 
<< pdiffusion >>
rect 464 230 465 231 
<< pdiffusion >>
rect 465 230 466 231 
<< pdiffusion >>
rect 466 230 467 231 
<< pdiffusion >>
rect 467 230 468 231 
<< m1 >>
rect 478 230 479 231 
<< pdiffusion >>
rect 480 230 481 231 
<< pdiffusion >>
rect 481 230 482 231 
<< pdiffusion >>
rect 482 230 483 231 
<< pdiffusion >>
rect 483 230 484 231 
<< pdiffusion >>
rect 484 230 485 231 
<< pdiffusion >>
rect 485 230 486 231 
<< m1 >>
rect 487 230 488 231 
<< pdiffusion >>
rect 498 230 499 231 
<< pdiffusion >>
rect 499 230 500 231 
<< pdiffusion >>
rect 500 230 501 231 
<< pdiffusion >>
rect 501 230 502 231 
<< pdiffusion >>
rect 502 230 503 231 
<< pdiffusion >>
rect 503 230 504 231 
<< m1 >>
rect 523 230 524 231 
<< pdiffusion >>
rect 12 231 13 232 
<< pdiffusion >>
rect 13 231 14 232 
<< pdiffusion >>
rect 14 231 15 232 
<< pdiffusion >>
rect 15 231 16 232 
<< pdiffusion >>
rect 16 231 17 232 
<< pdiffusion >>
rect 17 231 18 232 
<< m1 >>
rect 19 231 20 232 
<< pdiffusion >>
rect 30 231 31 232 
<< pdiffusion >>
rect 31 231 32 232 
<< pdiffusion >>
rect 32 231 33 232 
<< pdiffusion >>
rect 33 231 34 232 
<< pdiffusion >>
rect 34 231 35 232 
<< pdiffusion >>
rect 35 231 36 232 
<< m1 >>
rect 37 231 38 232 
<< pdiffusion >>
rect 48 231 49 232 
<< pdiffusion >>
rect 49 231 50 232 
<< pdiffusion >>
rect 50 231 51 232 
<< pdiffusion >>
rect 51 231 52 232 
<< pdiffusion >>
rect 52 231 53 232 
<< pdiffusion >>
rect 53 231 54 232 
<< m1 >>
rect 64 231 65 232 
<< pdiffusion >>
rect 66 231 67 232 
<< pdiffusion >>
rect 67 231 68 232 
<< pdiffusion >>
rect 68 231 69 232 
<< pdiffusion >>
rect 69 231 70 232 
<< pdiffusion >>
rect 70 231 71 232 
<< pdiffusion >>
rect 71 231 72 232 
<< pdiffusion >>
rect 84 231 85 232 
<< pdiffusion >>
rect 85 231 86 232 
<< pdiffusion >>
rect 86 231 87 232 
<< pdiffusion >>
rect 87 231 88 232 
<< pdiffusion >>
rect 88 231 89 232 
<< pdiffusion >>
rect 89 231 90 232 
<< m1 >>
rect 100 231 101 232 
<< pdiffusion >>
rect 102 231 103 232 
<< pdiffusion >>
rect 103 231 104 232 
<< pdiffusion >>
rect 104 231 105 232 
<< pdiffusion >>
rect 105 231 106 232 
<< pdiffusion >>
rect 106 231 107 232 
<< pdiffusion >>
rect 107 231 108 232 
<< m1 >>
rect 118 231 119 232 
<< pdiffusion >>
rect 120 231 121 232 
<< pdiffusion >>
rect 121 231 122 232 
<< pdiffusion >>
rect 122 231 123 232 
<< pdiffusion >>
rect 123 231 124 232 
<< pdiffusion >>
rect 124 231 125 232 
<< pdiffusion >>
rect 125 231 126 232 
<< m1 >>
rect 127 231 128 232 
<< pdiffusion >>
rect 138 231 139 232 
<< pdiffusion >>
rect 139 231 140 232 
<< pdiffusion >>
rect 140 231 141 232 
<< pdiffusion >>
rect 141 231 142 232 
<< pdiffusion >>
rect 142 231 143 232 
<< pdiffusion >>
rect 143 231 144 232 
<< m1 >>
rect 145 231 146 232 
<< m1 >>
rect 148 231 149 232 
<< pdiffusion >>
rect 156 231 157 232 
<< pdiffusion >>
rect 157 231 158 232 
<< pdiffusion >>
rect 158 231 159 232 
<< pdiffusion >>
rect 159 231 160 232 
<< pdiffusion >>
rect 160 231 161 232 
<< pdiffusion >>
rect 161 231 162 232 
<< m1 >>
rect 163 231 164 232 
<< m1 >>
rect 172 231 173 232 
<< pdiffusion >>
rect 174 231 175 232 
<< pdiffusion >>
rect 175 231 176 232 
<< pdiffusion >>
rect 176 231 177 232 
<< pdiffusion >>
rect 177 231 178 232 
<< pdiffusion >>
rect 178 231 179 232 
<< pdiffusion >>
rect 179 231 180 232 
<< m1 >>
rect 181 231 182 232 
<< m1 >>
rect 185 231 186 232 
<< m2 >>
rect 186 231 187 232 
<< m1 >>
rect 190 231 191 232 
<< pdiffusion >>
rect 192 231 193 232 
<< pdiffusion >>
rect 193 231 194 232 
<< pdiffusion >>
rect 194 231 195 232 
<< pdiffusion >>
rect 195 231 196 232 
<< pdiffusion >>
rect 196 231 197 232 
<< pdiffusion >>
rect 197 231 198 232 
<< m2 >>
rect 206 231 207 232 
<< m1 >>
rect 207 231 208 232 
<< pdiffusion >>
rect 210 231 211 232 
<< pdiffusion >>
rect 211 231 212 232 
<< pdiffusion >>
rect 212 231 213 232 
<< pdiffusion >>
rect 213 231 214 232 
<< pdiffusion >>
rect 214 231 215 232 
<< pdiffusion >>
rect 215 231 216 232 
<< m1 >>
rect 217 231 218 232 
<< m2 >>
rect 217 231 218 232 
<< m1 >>
rect 221 231 222 232 
<< m1 >>
rect 226 231 227 232 
<< pdiffusion >>
rect 228 231 229 232 
<< pdiffusion >>
rect 229 231 230 232 
<< pdiffusion >>
rect 230 231 231 232 
<< pdiffusion >>
rect 231 231 232 232 
<< pdiffusion >>
rect 232 231 233 232 
<< pdiffusion >>
rect 233 231 234 232 
<< m1 >>
rect 235 231 236 232 
<< m1 >>
rect 237 231 238 232 
<< m2 >>
rect 238 231 239 232 
<< m1 >>
rect 240 231 241 232 
<< pdiffusion >>
rect 246 231 247 232 
<< pdiffusion >>
rect 247 231 248 232 
<< pdiffusion >>
rect 248 231 249 232 
<< pdiffusion >>
rect 249 231 250 232 
<< pdiffusion >>
rect 250 231 251 232 
<< pdiffusion >>
rect 251 231 252 232 
<< m1 >>
rect 253 231 254 232 
<< pdiffusion >>
rect 264 231 265 232 
<< pdiffusion >>
rect 265 231 266 232 
<< pdiffusion >>
rect 266 231 267 232 
<< pdiffusion >>
rect 267 231 268 232 
<< pdiffusion >>
rect 268 231 269 232 
<< pdiffusion >>
rect 269 231 270 232 
<< m1 >>
rect 272 231 273 232 
<< pdiffusion >>
rect 282 231 283 232 
<< pdiffusion >>
rect 283 231 284 232 
<< pdiffusion >>
rect 284 231 285 232 
<< pdiffusion >>
rect 285 231 286 232 
<< pdiffusion >>
rect 286 231 287 232 
<< pdiffusion >>
rect 287 231 288 232 
<< m1 >>
rect 290 231 291 232 
<< m1 >>
rect 292 231 293 232 
<< m1 >>
rect 296 231 297 232 
<< m1 >>
rect 298 231 299 232 
<< pdiffusion >>
rect 300 231 301 232 
<< pdiffusion >>
rect 301 231 302 232 
<< pdiffusion >>
rect 302 231 303 232 
<< pdiffusion >>
rect 303 231 304 232 
<< pdiffusion >>
rect 304 231 305 232 
<< pdiffusion >>
rect 305 231 306 232 
<< m1 >>
rect 307 231 308 232 
<< m2 >>
rect 308 231 309 232 
<< m1 >>
rect 316 231 317 232 
<< pdiffusion >>
rect 318 231 319 232 
<< pdiffusion >>
rect 319 231 320 232 
<< pdiffusion >>
rect 320 231 321 232 
<< pdiffusion >>
rect 321 231 322 232 
<< pdiffusion >>
rect 322 231 323 232 
<< pdiffusion >>
rect 323 231 324 232 
<< pdiffusion >>
rect 336 231 337 232 
<< pdiffusion >>
rect 337 231 338 232 
<< pdiffusion >>
rect 338 231 339 232 
<< pdiffusion >>
rect 339 231 340 232 
<< pdiffusion >>
rect 340 231 341 232 
<< pdiffusion >>
rect 341 231 342 232 
<< m1 >>
rect 352 231 353 232 
<< pdiffusion >>
rect 354 231 355 232 
<< pdiffusion >>
rect 355 231 356 232 
<< pdiffusion >>
rect 356 231 357 232 
<< pdiffusion >>
rect 357 231 358 232 
<< pdiffusion >>
rect 358 231 359 232 
<< pdiffusion >>
rect 359 231 360 232 
<< pdiffusion >>
rect 372 231 373 232 
<< pdiffusion >>
rect 373 231 374 232 
<< pdiffusion >>
rect 374 231 375 232 
<< pdiffusion >>
rect 375 231 376 232 
<< pdiffusion >>
rect 376 231 377 232 
<< pdiffusion >>
rect 377 231 378 232 
<< m1 >>
rect 379 231 380 232 
<< m2 >>
rect 380 231 381 232 
<< m1 >>
rect 383 231 384 232 
<< pdiffusion >>
rect 390 231 391 232 
<< pdiffusion >>
rect 391 231 392 232 
<< pdiffusion >>
rect 392 231 393 232 
<< pdiffusion >>
rect 393 231 394 232 
<< pdiffusion >>
rect 394 231 395 232 
<< pdiffusion >>
rect 395 231 396 232 
<< pdiffusion >>
rect 408 231 409 232 
<< pdiffusion >>
rect 409 231 410 232 
<< pdiffusion >>
rect 410 231 411 232 
<< pdiffusion >>
rect 411 231 412 232 
<< pdiffusion >>
rect 412 231 413 232 
<< pdiffusion >>
rect 413 231 414 232 
<< m1 >>
rect 416 231 417 232 
<< m1 >>
rect 419 231 420 232 
<< m1 >>
rect 421 231 422 232 
<< m2 >>
rect 422 231 423 232 
<< pdiffusion >>
rect 426 231 427 232 
<< pdiffusion >>
rect 427 231 428 232 
<< pdiffusion >>
rect 428 231 429 232 
<< pdiffusion >>
rect 429 231 430 232 
<< pdiffusion >>
rect 430 231 431 232 
<< pdiffusion >>
rect 431 231 432 232 
<< m1 >>
rect 434 231 435 232 
<< m1 >>
rect 442 231 443 232 
<< pdiffusion >>
rect 444 231 445 232 
<< pdiffusion >>
rect 445 231 446 232 
<< pdiffusion >>
rect 446 231 447 232 
<< pdiffusion >>
rect 447 231 448 232 
<< pdiffusion >>
rect 448 231 449 232 
<< pdiffusion >>
rect 449 231 450 232 
<< pdiffusion >>
rect 462 231 463 232 
<< pdiffusion >>
rect 463 231 464 232 
<< pdiffusion >>
rect 464 231 465 232 
<< pdiffusion >>
rect 465 231 466 232 
<< pdiffusion >>
rect 466 231 467 232 
<< pdiffusion >>
rect 467 231 468 232 
<< m1 >>
rect 478 231 479 232 
<< pdiffusion >>
rect 480 231 481 232 
<< pdiffusion >>
rect 481 231 482 232 
<< pdiffusion >>
rect 482 231 483 232 
<< pdiffusion >>
rect 483 231 484 232 
<< pdiffusion >>
rect 484 231 485 232 
<< pdiffusion >>
rect 485 231 486 232 
<< m1 >>
rect 487 231 488 232 
<< pdiffusion >>
rect 498 231 499 232 
<< pdiffusion >>
rect 499 231 500 232 
<< pdiffusion >>
rect 500 231 501 232 
<< pdiffusion >>
rect 501 231 502 232 
<< pdiffusion >>
rect 502 231 503 232 
<< pdiffusion >>
rect 503 231 504 232 
<< m1 >>
rect 523 231 524 232 
<< pdiffusion >>
rect 12 232 13 233 
<< pdiffusion >>
rect 13 232 14 233 
<< pdiffusion >>
rect 14 232 15 233 
<< pdiffusion >>
rect 15 232 16 233 
<< pdiffusion >>
rect 16 232 17 233 
<< pdiffusion >>
rect 17 232 18 233 
<< m1 >>
rect 19 232 20 233 
<< pdiffusion >>
rect 30 232 31 233 
<< pdiffusion >>
rect 31 232 32 233 
<< pdiffusion >>
rect 32 232 33 233 
<< pdiffusion >>
rect 33 232 34 233 
<< pdiffusion >>
rect 34 232 35 233 
<< pdiffusion >>
rect 35 232 36 233 
<< m1 >>
rect 37 232 38 233 
<< pdiffusion >>
rect 48 232 49 233 
<< pdiffusion >>
rect 49 232 50 233 
<< pdiffusion >>
rect 50 232 51 233 
<< pdiffusion >>
rect 51 232 52 233 
<< pdiffusion >>
rect 52 232 53 233 
<< pdiffusion >>
rect 53 232 54 233 
<< m1 >>
rect 64 232 65 233 
<< pdiffusion >>
rect 66 232 67 233 
<< pdiffusion >>
rect 67 232 68 233 
<< pdiffusion >>
rect 68 232 69 233 
<< pdiffusion >>
rect 69 232 70 233 
<< pdiffusion >>
rect 70 232 71 233 
<< pdiffusion >>
rect 71 232 72 233 
<< pdiffusion >>
rect 84 232 85 233 
<< pdiffusion >>
rect 85 232 86 233 
<< pdiffusion >>
rect 86 232 87 233 
<< pdiffusion >>
rect 87 232 88 233 
<< pdiffusion >>
rect 88 232 89 233 
<< pdiffusion >>
rect 89 232 90 233 
<< m1 >>
rect 100 232 101 233 
<< pdiffusion >>
rect 102 232 103 233 
<< pdiffusion >>
rect 103 232 104 233 
<< pdiffusion >>
rect 104 232 105 233 
<< pdiffusion >>
rect 105 232 106 233 
<< pdiffusion >>
rect 106 232 107 233 
<< pdiffusion >>
rect 107 232 108 233 
<< m1 >>
rect 118 232 119 233 
<< pdiffusion >>
rect 120 232 121 233 
<< pdiffusion >>
rect 121 232 122 233 
<< pdiffusion >>
rect 122 232 123 233 
<< pdiffusion >>
rect 123 232 124 233 
<< pdiffusion >>
rect 124 232 125 233 
<< pdiffusion >>
rect 125 232 126 233 
<< m1 >>
rect 127 232 128 233 
<< pdiffusion >>
rect 138 232 139 233 
<< pdiffusion >>
rect 139 232 140 233 
<< pdiffusion >>
rect 140 232 141 233 
<< pdiffusion >>
rect 141 232 142 233 
<< pdiffusion >>
rect 142 232 143 233 
<< pdiffusion >>
rect 143 232 144 233 
<< m1 >>
rect 145 232 146 233 
<< m1 >>
rect 148 232 149 233 
<< pdiffusion >>
rect 156 232 157 233 
<< pdiffusion >>
rect 157 232 158 233 
<< pdiffusion >>
rect 158 232 159 233 
<< pdiffusion >>
rect 159 232 160 233 
<< pdiffusion >>
rect 160 232 161 233 
<< pdiffusion >>
rect 161 232 162 233 
<< m1 >>
rect 163 232 164 233 
<< m1 >>
rect 172 232 173 233 
<< pdiffusion >>
rect 174 232 175 233 
<< pdiffusion >>
rect 175 232 176 233 
<< pdiffusion >>
rect 176 232 177 233 
<< pdiffusion >>
rect 177 232 178 233 
<< pdiffusion >>
rect 178 232 179 233 
<< pdiffusion >>
rect 179 232 180 233 
<< m1 >>
rect 181 232 182 233 
<< m1 >>
rect 185 232 186 233 
<< m2 >>
rect 186 232 187 233 
<< m1 >>
rect 190 232 191 233 
<< pdiffusion >>
rect 192 232 193 233 
<< pdiffusion >>
rect 193 232 194 233 
<< pdiffusion >>
rect 194 232 195 233 
<< pdiffusion >>
rect 195 232 196 233 
<< pdiffusion >>
rect 196 232 197 233 
<< pdiffusion >>
rect 197 232 198 233 
<< m2 >>
rect 206 232 207 233 
<< m1 >>
rect 207 232 208 233 
<< pdiffusion >>
rect 210 232 211 233 
<< pdiffusion >>
rect 211 232 212 233 
<< pdiffusion >>
rect 212 232 213 233 
<< pdiffusion >>
rect 213 232 214 233 
<< pdiffusion >>
rect 214 232 215 233 
<< pdiffusion >>
rect 215 232 216 233 
<< m1 >>
rect 217 232 218 233 
<< m2 >>
rect 217 232 218 233 
<< m1 >>
rect 221 232 222 233 
<< m1 >>
rect 226 232 227 233 
<< pdiffusion >>
rect 228 232 229 233 
<< pdiffusion >>
rect 229 232 230 233 
<< pdiffusion >>
rect 230 232 231 233 
<< pdiffusion >>
rect 231 232 232 233 
<< pdiffusion >>
rect 232 232 233 233 
<< pdiffusion >>
rect 233 232 234 233 
<< m1 >>
rect 235 232 236 233 
<< m1 >>
rect 237 232 238 233 
<< m2 >>
rect 238 232 239 233 
<< m1 >>
rect 240 232 241 233 
<< pdiffusion >>
rect 246 232 247 233 
<< pdiffusion >>
rect 247 232 248 233 
<< pdiffusion >>
rect 248 232 249 233 
<< pdiffusion >>
rect 249 232 250 233 
<< pdiffusion >>
rect 250 232 251 233 
<< pdiffusion >>
rect 251 232 252 233 
<< m1 >>
rect 253 232 254 233 
<< pdiffusion >>
rect 264 232 265 233 
<< pdiffusion >>
rect 265 232 266 233 
<< pdiffusion >>
rect 266 232 267 233 
<< pdiffusion >>
rect 267 232 268 233 
<< pdiffusion >>
rect 268 232 269 233 
<< pdiffusion >>
rect 269 232 270 233 
<< m1 >>
rect 272 232 273 233 
<< pdiffusion >>
rect 282 232 283 233 
<< pdiffusion >>
rect 283 232 284 233 
<< pdiffusion >>
rect 284 232 285 233 
<< pdiffusion >>
rect 285 232 286 233 
<< pdiffusion >>
rect 286 232 287 233 
<< pdiffusion >>
rect 287 232 288 233 
<< m1 >>
rect 290 232 291 233 
<< m1 >>
rect 292 232 293 233 
<< m1 >>
rect 296 232 297 233 
<< m1 >>
rect 298 232 299 233 
<< pdiffusion >>
rect 300 232 301 233 
<< pdiffusion >>
rect 301 232 302 233 
<< pdiffusion >>
rect 302 232 303 233 
<< pdiffusion >>
rect 303 232 304 233 
<< pdiffusion >>
rect 304 232 305 233 
<< pdiffusion >>
rect 305 232 306 233 
<< m1 >>
rect 307 232 308 233 
<< m2 >>
rect 308 232 309 233 
<< m1 >>
rect 316 232 317 233 
<< pdiffusion >>
rect 318 232 319 233 
<< pdiffusion >>
rect 319 232 320 233 
<< pdiffusion >>
rect 320 232 321 233 
<< pdiffusion >>
rect 321 232 322 233 
<< pdiffusion >>
rect 322 232 323 233 
<< pdiffusion >>
rect 323 232 324 233 
<< pdiffusion >>
rect 336 232 337 233 
<< pdiffusion >>
rect 337 232 338 233 
<< pdiffusion >>
rect 338 232 339 233 
<< pdiffusion >>
rect 339 232 340 233 
<< pdiffusion >>
rect 340 232 341 233 
<< pdiffusion >>
rect 341 232 342 233 
<< m1 >>
rect 352 232 353 233 
<< pdiffusion >>
rect 354 232 355 233 
<< pdiffusion >>
rect 355 232 356 233 
<< pdiffusion >>
rect 356 232 357 233 
<< pdiffusion >>
rect 357 232 358 233 
<< pdiffusion >>
rect 358 232 359 233 
<< pdiffusion >>
rect 359 232 360 233 
<< pdiffusion >>
rect 372 232 373 233 
<< pdiffusion >>
rect 373 232 374 233 
<< pdiffusion >>
rect 374 232 375 233 
<< pdiffusion >>
rect 375 232 376 233 
<< pdiffusion >>
rect 376 232 377 233 
<< pdiffusion >>
rect 377 232 378 233 
<< m1 >>
rect 379 232 380 233 
<< m2 >>
rect 380 232 381 233 
<< m1 >>
rect 383 232 384 233 
<< pdiffusion >>
rect 390 232 391 233 
<< pdiffusion >>
rect 391 232 392 233 
<< pdiffusion >>
rect 392 232 393 233 
<< pdiffusion >>
rect 393 232 394 233 
<< pdiffusion >>
rect 394 232 395 233 
<< pdiffusion >>
rect 395 232 396 233 
<< pdiffusion >>
rect 408 232 409 233 
<< pdiffusion >>
rect 409 232 410 233 
<< pdiffusion >>
rect 410 232 411 233 
<< pdiffusion >>
rect 411 232 412 233 
<< pdiffusion >>
rect 412 232 413 233 
<< pdiffusion >>
rect 413 232 414 233 
<< m1 >>
rect 416 232 417 233 
<< m1 >>
rect 419 232 420 233 
<< m1 >>
rect 421 232 422 233 
<< m2 >>
rect 422 232 423 233 
<< pdiffusion >>
rect 426 232 427 233 
<< pdiffusion >>
rect 427 232 428 233 
<< pdiffusion >>
rect 428 232 429 233 
<< pdiffusion >>
rect 429 232 430 233 
<< pdiffusion >>
rect 430 232 431 233 
<< pdiffusion >>
rect 431 232 432 233 
<< m1 >>
rect 434 232 435 233 
<< m1 >>
rect 442 232 443 233 
<< pdiffusion >>
rect 444 232 445 233 
<< pdiffusion >>
rect 445 232 446 233 
<< pdiffusion >>
rect 446 232 447 233 
<< pdiffusion >>
rect 447 232 448 233 
<< pdiffusion >>
rect 448 232 449 233 
<< pdiffusion >>
rect 449 232 450 233 
<< pdiffusion >>
rect 462 232 463 233 
<< pdiffusion >>
rect 463 232 464 233 
<< pdiffusion >>
rect 464 232 465 233 
<< pdiffusion >>
rect 465 232 466 233 
<< pdiffusion >>
rect 466 232 467 233 
<< pdiffusion >>
rect 467 232 468 233 
<< m1 >>
rect 478 232 479 233 
<< pdiffusion >>
rect 480 232 481 233 
<< pdiffusion >>
rect 481 232 482 233 
<< pdiffusion >>
rect 482 232 483 233 
<< pdiffusion >>
rect 483 232 484 233 
<< pdiffusion >>
rect 484 232 485 233 
<< pdiffusion >>
rect 485 232 486 233 
<< m1 >>
rect 487 232 488 233 
<< pdiffusion >>
rect 498 232 499 233 
<< pdiffusion >>
rect 499 232 500 233 
<< pdiffusion >>
rect 500 232 501 233 
<< pdiffusion >>
rect 501 232 502 233 
<< pdiffusion >>
rect 502 232 503 233 
<< pdiffusion >>
rect 503 232 504 233 
<< m1 >>
rect 523 232 524 233 
<< pdiffusion >>
rect 12 233 13 234 
<< pdiffusion >>
rect 13 233 14 234 
<< pdiffusion >>
rect 14 233 15 234 
<< pdiffusion >>
rect 15 233 16 234 
<< m1 >>
rect 16 233 17 234 
<< pdiffusion >>
rect 16 233 17 234 
<< pdiffusion >>
rect 17 233 18 234 
<< m1 >>
rect 19 233 20 234 
<< pdiffusion >>
rect 30 233 31 234 
<< pdiffusion >>
rect 31 233 32 234 
<< pdiffusion >>
rect 32 233 33 234 
<< pdiffusion >>
rect 33 233 34 234 
<< m1 >>
rect 34 233 35 234 
<< pdiffusion >>
rect 34 233 35 234 
<< pdiffusion >>
rect 35 233 36 234 
<< m1 >>
rect 37 233 38 234 
<< pdiffusion >>
rect 48 233 49 234 
<< pdiffusion >>
rect 49 233 50 234 
<< pdiffusion >>
rect 50 233 51 234 
<< pdiffusion >>
rect 51 233 52 234 
<< m1 >>
rect 52 233 53 234 
<< pdiffusion >>
rect 52 233 53 234 
<< pdiffusion >>
rect 53 233 54 234 
<< m1 >>
rect 64 233 65 234 
<< pdiffusion >>
rect 66 233 67 234 
<< pdiffusion >>
rect 67 233 68 234 
<< pdiffusion >>
rect 68 233 69 234 
<< pdiffusion >>
rect 69 233 70 234 
<< pdiffusion >>
rect 70 233 71 234 
<< pdiffusion >>
rect 71 233 72 234 
<< pdiffusion >>
rect 84 233 85 234 
<< m1 >>
rect 85 233 86 234 
<< pdiffusion >>
rect 85 233 86 234 
<< pdiffusion >>
rect 86 233 87 234 
<< pdiffusion >>
rect 87 233 88 234 
<< pdiffusion >>
rect 88 233 89 234 
<< pdiffusion >>
rect 89 233 90 234 
<< m1 >>
rect 100 233 101 234 
<< pdiffusion >>
rect 102 233 103 234 
<< pdiffusion >>
rect 103 233 104 234 
<< pdiffusion >>
rect 104 233 105 234 
<< pdiffusion >>
rect 105 233 106 234 
<< pdiffusion >>
rect 106 233 107 234 
<< pdiffusion >>
rect 107 233 108 234 
<< m1 >>
rect 118 233 119 234 
<< pdiffusion >>
rect 120 233 121 234 
<< pdiffusion >>
rect 121 233 122 234 
<< pdiffusion >>
rect 122 233 123 234 
<< pdiffusion >>
rect 123 233 124 234 
<< pdiffusion >>
rect 124 233 125 234 
<< pdiffusion >>
rect 125 233 126 234 
<< m1 >>
rect 127 233 128 234 
<< pdiffusion >>
rect 138 233 139 234 
<< pdiffusion >>
rect 139 233 140 234 
<< pdiffusion >>
rect 140 233 141 234 
<< pdiffusion >>
rect 141 233 142 234 
<< m1 >>
rect 142 233 143 234 
<< pdiffusion >>
rect 142 233 143 234 
<< pdiffusion >>
rect 143 233 144 234 
<< m1 >>
rect 145 233 146 234 
<< m1 >>
rect 148 233 149 234 
<< pdiffusion >>
rect 156 233 157 234 
<< pdiffusion >>
rect 157 233 158 234 
<< pdiffusion >>
rect 158 233 159 234 
<< pdiffusion >>
rect 159 233 160 234 
<< pdiffusion >>
rect 160 233 161 234 
<< pdiffusion >>
rect 161 233 162 234 
<< m1 >>
rect 163 233 164 234 
<< m1 >>
rect 172 233 173 234 
<< pdiffusion >>
rect 174 233 175 234 
<< m1 >>
rect 175 233 176 234 
<< pdiffusion >>
rect 175 233 176 234 
<< pdiffusion >>
rect 176 233 177 234 
<< pdiffusion >>
rect 177 233 178 234 
<< pdiffusion >>
rect 178 233 179 234 
<< pdiffusion >>
rect 179 233 180 234 
<< m1 >>
rect 181 233 182 234 
<< m1 >>
rect 185 233 186 234 
<< m2 >>
rect 186 233 187 234 
<< m1 >>
rect 190 233 191 234 
<< pdiffusion >>
rect 192 233 193 234 
<< pdiffusion >>
rect 193 233 194 234 
<< pdiffusion >>
rect 194 233 195 234 
<< pdiffusion >>
rect 195 233 196 234 
<< pdiffusion >>
rect 196 233 197 234 
<< pdiffusion >>
rect 197 233 198 234 
<< m2 >>
rect 206 233 207 234 
<< m1 >>
rect 207 233 208 234 
<< pdiffusion >>
rect 210 233 211 234 
<< pdiffusion >>
rect 211 233 212 234 
<< pdiffusion >>
rect 212 233 213 234 
<< pdiffusion >>
rect 213 233 214 234 
<< m1 >>
rect 214 233 215 234 
<< pdiffusion >>
rect 214 233 215 234 
<< pdiffusion >>
rect 215 233 216 234 
<< m1 >>
rect 217 233 218 234 
<< m2 >>
rect 217 233 218 234 
<< m1 >>
rect 221 233 222 234 
<< m1 >>
rect 226 233 227 234 
<< pdiffusion >>
rect 228 233 229 234 
<< m1 >>
rect 229 233 230 234 
<< pdiffusion >>
rect 229 233 230 234 
<< pdiffusion >>
rect 230 233 231 234 
<< pdiffusion >>
rect 231 233 232 234 
<< pdiffusion >>
rect 232 233 233 234 
<< pdiffusion >>
rect 233 233 234 234 
<< m1 >>
rect 235 233 236 234 
<< m1 >>
rect 237 233 238 234 
<< m2 >>
rect 238 233 239 234 
<< m1 >>
rect 240 233 241 234 
<< pdiffusion >>
rect 246 233 247 234 
<< pdiffusion >>
rect 247 233 248 234 
<< pdiffusion >>
rect 248 233 249 234 
<< pdiffusion >>
rect 249 233 250 234 
<< m1 >>
rect 250 233 251 234 
<< pdiffusion >>
rect 250 233 251 234 
<< pdiffusion >>
rect 251 233 252 234 
<< m1 >>
rect 253 233 254 234 
<< pdiffusion >>
rect 264 233 265 234 
<< pdiffusion >>
rect 265 233 266 234 
<< pdiffusion >>
rect 266 233 267 234 
<< pdiffusion >>
rect 267 233 268 234 
<< pdiffusion >>
rect 268 233 269 234 
<< pdiffusion >>
rect 269 233 270 234 
<< m1 >>
rect 272 233 273 234 
<< pdiffusion >>
rect 282 233 283 234 
<< pdiffusion >>
rect 283 233 284 234 
<< pdiffusion >>
rect 284 233 285 234 
<< pdiffusion >>
rect 285 233 286 234 
<< pdiffusion >>
rect 286 233 287 234 
<< pdiffusion >>
rect 287 233 288 234 
<< m1 >>
rect 290 233 291 234 
<< m1 >>
rect 292 233 293 234 
<< m1 >>
rect 296 233 297 234 
<< m1 >>
rect 298 233 299 234 
<< pdiffusion >>
rect 300 233 301 234 
<< m1 >>
rect 301 233 302 234 
<< pdiffusion >>
rect 301 233 302 234 
<< pdiffusion >>
rect 302 233 303 234 
<< pdiffusion >>
rect 303 233 304 234 
<< pdiffusion >>
rect 304 233 305 234 
<< pdiffusion >>
rect 305 233 306 234 
<< m1 >>
rect 307 233 308 234 
<< m2 >>
rect 308 233 309 234 
<< m1 >>
rect 316 233 317 234 
<< pdiffusion >>
rect 318 233 319 234 
<< pdiffusion >>
rect 319 233 320 234 
<< pdiffusion >>
rect 320 233 321 234 
<< pdiffusion >>
rect 321 233 322 234 
<< pdiffusion >>
rect 322 233 323 234 
<< pdiffusion >>
rect 323 233 324 234 
<< pdiffusion >>
rect 336 233 337 234 
<< m1 >>
rect 337 233 338 234 
<< pdiffusion >>
rect 337 233 338 234 
<< pdiffusion >>
rect 338 233 339 234 
<< pdiffusion >>
rect 339 233 340 234 
<< pdiffusion >>
rect 340 233 341 234 
<< pdiffusion >>
rect 341 233 342 234 
<< m1 >>
rect 352 233 353 234 
<< pdiffusion >>
rect 354 233 355 234 
<< pdiffusion >>
rect 355 233 356 234 
<< pdiffusion >>
rect 356 233 357 234 
<< pdiffusion >>
rect 357 233 358 234 
<< pdiffusion >>
rect 358 233 359 234 
<< pdiffusion >>
rect 359 233 360 234 
<< pdiffusion >>
rect 372 233 373 234 
<< pdiffusion >>
rect 373 233 374 234 
<< pdiffusion >>
rect 374 233 375 234 
<< pdiffusion >>
rect 375 233 376 234 
<< pdiffusion >>
rect 376 233 377 234 
<< pdiffusion >>
rect 377 233 378 234 
<< m1 >>
rect 379 233 380 234 
<< m2 >>
rect 380 233 381 234 
<< m1 >>
rect 383 233 384 234 
<< pdiffusion >>
rect 390 233 391 234 
<< pdiffusion >>
rect 391 233 392 234 
<< pdiffusion >>
rect 392 233 393 234 
<< pdiffusion >>
rect 393 233 394 234 
<< m1 >>
rect 394 233 395 234 
<< pdiffusion >>
rect 394 233 395 234 
<< pdiffusion >>
rect 395 233 396 234 
<< pdiffusion >>
rect 408 233 409 234 
<< pdiffusion >>
rect 409 233 410 234 
<< pdiffusion >>
rect 410 233 411 234 
<< pdiffusion >>
rect 411 233 412 234 
<< pdiffusion >>
rect 412 233 413 234 
<< pdiffusion >>
rect 413 233 414 234 
<< m1 >>
rect 416 233 417 234 
<< m1 >>
rect 419 233 420 234 
<< m1 >>
rect 421 233 422 234 
<< m2 >>
rect 422 233 423 234 
<< pdiffusion >>
rect 426 233 427 234 
<< pdiffusion >>
rect 427 233 428 234 
<< pdiffusion >>
rect 428 233 429 234 
<< pdiffusion >>
rect 429 233 430 234 
<< pdiffusion >>
rect 430 233 431 234 
<< pdiffusion >>
rect 431 233 432 234 
<< m1 >>
rect 434 233 435 234 
<< m1 >>
rect 442 233 443 234 
<< pdiffusion >>
rect 444 233 445 234 
<< pdiffusion >>
rect 445 233 446 234 
<< pdiffusion >>
rect 446 233 447 234 
<< pdiffusion >>
rect 447 233 448 234 
<< pdiffusion >>
rect 448 233 449 234 
<< pdiffusion >>
rect 449 233 450 234 
<< pdiffusion >>
rect 462 233 463 234 
<< pdiffusion >>
rect 463 233 464 234 
<< pdiffusion >>
rect 464 233 465 234 
<< pdiffusion >>
rect 465 233 466 234 
<< pdiffusion >>
rect 466 233 467 234 
<< pdiffusion >>
rect 467 233 468 234 
<< m1 >>
rect 478 233 479 234 
<< pdiffusion >>
rect 480 233 481 234 
<< pdiffusion >>
rect 481 233 482 234 
<< pdiffusion >>
rect 482 233 483 234 
<< pdiffusion >>
rect 483 233 484 234 
<< pdiffusion >>
rect 484 233 485 234 
<< pdiffusion >>
rect 485 233 486 234 
<< m1 >>
rect 487 233 488 234 
<< pdiffusion >>
rect 498 233 499 234 
<< pdiffusion >>
rect 499 233 500 234 
<< pdiffusion >>
rect 500 233 501 234 
<< pdiffusion >>
rect 501 233 502 234 
<< pdiffusion >>
rect 502 233 503 234 
<< pdiffusion >>
rect 503 233 504 234 
<< m1 >>
rect 523 233 524 234 
<< m1 >>
rect 16 234 17 235 
<< m1 >>
rect 19 234 20 235 
<< m1 >>
rect 34 234 35 235 
<< m1 >>
rect 37 234 38 235 
<< m1 >>
rect 52 234 53 235 
<< m2 >>
rect 56 234 57 235 
<< m1 >>
rect 57 234 58 235 
<< m2 >>
rect 57 234 58 235 
<< m2c >>
rect 57 234 58 235 
<< m1 >>
rect 57 234 58 235 
<< m2 >>
rect 57 234 58 235 
<< m1 >>
rect 58 234 59 235 
<< m1 >>
rect 59 234 60 235 
<< m1 >>
rect 60 234 61 235 
<< m1 >>
rect 61 234 62 235 
<< m1 >>
rect 62 234 63 235 
<< m1 >>
rect 63 234 64 235 
<< m1 >>
rect 64 234 65 235 
<< m1 >>
rect 85 234 86 235 
<< m1 >>
rect 100 234 101 235 
<< m1 >>
rect 118 234 119 235 
<< m1 >>
rect 127 234 128 235 
<< m1 >>
rect 142 234 143 235 
<< m1 >>
rect 145 234 146 235 
<< m1 >>
rect 148 234 149 235 
<< m1 >>
rect 163 234 164 235 
<< m1 >>
rect 172 234 173 235 
<< m1 >>
rect 175 234 176 235 
<< m1 >>
rect 181 234 182 235 
<< m1 >>
rect 185 234 186 235 
<< m2 >>
rect 186 234 187 235 
<< m1 >>
rect 190 234 191 235 
<< m1 >>
rect 199 234 200 235 
<< m1 >>
rect 200 234 201 235 
<< m1 >>
rect 201 234 202 235 
<< m1 >>
rect 202 234 203 235 
<< m1 >>
rect 203 234 204 235 
<< m1 >>
rect 204 234 205 235 
<< m1 >>
rect 205 234 206 235 
<< m2 >>
rect 205 234 206 235 
<< m2c >>
rect 205 234 206 235 
<< m1 >>
rect 205 234 206 235 
<< m2 >>
rect 205 234 206 235 
<< m2 >>
rect 206 234 207 235 
<< m1 >>
rect 207 234 208 235 
<< m1 >>
rect 214 234 215 235 
<< m1 >>
rect 217 234 218 235 
<< m2 >>
rect 217 234 218 235 
<< m1 >>
rect 221 234 222 235 
<< m1 >>
rect 226 234 227 235 
<< m1 >>
rect 229 234 230 235 
<< m1 >>
rect 235 234 236 235 
<< m1 >>
rect 237 234 238 235 
<< m2 >>
rect 238 234 239 235 
<< m1 >>
rect 240 234 241 235 
<< m1 >>
rect 250 234 251 235 
<< m1 >>
rect 253 234 254 235 
<< m1 >>
rect 272 234 273 235 
<< m1 >>
rect 290 234 291 235 
<< m1 >>
rect 292 234 293 235 
<< m1 >>
rect 296 234 297 235 
<< m1 >>
rect 298 234 299 235 
<< m1 >>
rect 301 234 302 235 
<< m1 >>
rect 307 234 308 235 
<< m2 >>
rect 308 234 309 235 
<< m1 >>
rect 316 234 317 235 
<< m1 >>
rect 337 234 338 235 
<< m1 >>
rect 352 234 353 235 
<< m1 >>
rect 379 234 380 235 
<< m2 >>
rect 380 234 381 235 
<< m1 >>
rect 383 234 384 235 
<< m1 >>
rect 394 234 395 235 
<< m1 >>
rect 416 234 417 235 
<< m1 >>
rect 419 234 420 235 
<< m1 >>
rect 421 234 422 235 
<< m2 >>
rect 422 234 423 235 
<< m1 >>
rect 434 234 435 235 
<< m1 >>
rect 442 234 443 235 
<< m1 >>
rect 478 234 479 235 
<< m1 >>
rect 487 234 488 235 
<< m1 >>
rect 523 234 524 235 
<< m1 >>
rect 16 235 17 236 
<< m1 >>
rect 17 235 18 236 
<< m2 >>
rect 17 235 18 236 
<< m2c >>
rect 17 235 18 236 
<< m1 >>
rect 17 235 18 236 
<< m2 >>
rect 17 235 18 236 
<< m2 >>
rect 18 235 19 236 
<< m1 >>
rect 19 235 20 236 
<< m2 >>
rect 19 235 20 236 
<< m2 >>
rect 20 235 21 236 
<< m1 >>
rect 21 235 22 236 
<< m2 >>
rect 21 235 22 236 
<< m2c >>
rect 21 235 22 236 
<< m1 >>
rect 21 235 22 236 
<< m2 >>
rect 21 235 22 236 
<< m1 >>
rect 22 235 23 236 
<< m1 >>
rect 34 235 35 236 
<< m1 >>
rect 35 235 36 236 
<< m1 >>
rect 36 235 37 236 
<< m1 >>
rect 37 235 38 236 
<< m1 >>
rect 52 235 53 236 
<< m1 >>
rect 53 235 54 236 
<< m1 >>
rect 54 235 55 236 
<< m1 >>
rect 55 235 56 236 
<< m2 >>
rect 56 235 57 236 
<< m1 >>
rect 85 235 86 236 
<< m1 >>
rect 100 235 101 236 
<< m1 >>
rect 118 235 119 236 
<< m1 >>
rect 127 235 128 236 
<< m1 >>
rect 142 235 143 236 
<< m1 >>
rect 143 235 144 236 
<< m1 >>
rect 144 235 145 236 
<< m1 >>
rect 145 235 146 236 
<< m1 >>
rect 148 235 149 236 
<< m1 >>
rect 163 235 164 236 
<< m1 >>
rect 172 235 173 236 
<< m1 >>
rect 175 235 176 236 
<< m1 >>
rect 181 235 182 236 
<< m1 >>
rect 185 235 186 236 
<< m2 >>
rect 186 235 187 236 
<< m1 >>
rect 190 235 191 236 
<< m1 >>
rect 199 235 200 236 
<< m1 >>
rect 207 235 208 236 
<< m1 >>
rect 214 235 215 236 
<< m1 >>
rect 215 235 216 236 
<< m1 >>
rect 216 235 217 236 
<< m1 >>
rect 217 235 218 236 
<< m2 >>
rect 217 235 218 236 
<< m1 >>
rect 221 235 222 236 
<< m1 >>
rect 226 235 227 236 
<< m1 >>
rect 229 235 230 236 
<< m1 >>
rect 233 235 234 236 
<< m2 >>
rect 233 235 234 236 
<< m2c >>
rect 233 235 234 236 
<< m1 >>
rect 233 235 234 236 
<< m2 >>
rect 233 235 234 236 
<< m2 >>
rect 234 235 235 236 
<< m1 >>
rect 235 235 236 236 
<< m2 >>
rect 235 235 236 236 
<< m2 >>
rect 236 235 237 236 
<< m1 >>
rect 237 235 238 236 
<< m2 >>
rect 237 235 238 236 
<< m2 >>
rect 238 235 239 236 
<< m1 >>
rect 240 235 241 236 
<< m1 >>
rect 250 235 251 236 
<< m1 >>
rect 251 235 252 236 
<< m1 >>
rect 252 235 253 236 
<< m1 >>
rect 253 235 254 236 
<< m1 >>
rect 272 235 273 236 
<< m1 >>
rect 290 235 291 236 
<< m1 >>
rect 292 235 293 236 
<< m1 >>
rect 296 235 297 236 
<< m1 >>
rect 298 235 299 236 
<< m1 >>
rect 301 235 302 236 
<< m1 >>
rect 305 235 306 236 
<< m2 >>
rect 305 235 306 236 
<< m2c >>
rect 305 235 306 236 
<< m1 >>
rect 305 235 306 236 
<< m2 >>
rect 305 235 306 236 
<< m2 >>
rect 306 235 307 236 
<< m1 >>
rect 307 235 308 236 
<< m2 >>
rect 307 235 308 236 
<< m2 >>
rect 308 235 309 236 
<< m1 >>
rect 316 235 317 236 
<< m1 >>
rect 337 235 338 236 
<< m1 >>
rect 352 235 353 236 
<< m1 >>
rect 379 235 380 236 
<< m2 >>
rect 380 235 381 236 
<< m1 >>
rect 383 235 384 236 
<< m1 >>
rect 394 235 395 236 
<< m1 >>
rect 416 235 417 236 
<< m1 >>
rect 419 235 420 236 
<< m1 >>
rect 421 235 422 236 
<< m2 >>
rect 422 235 423 236 
<< m1 >>
rect 434 235 435 236 
<< m1 >>
rect 442 235 443 236 
<< m1 >>
rect 478 235 479 236 
<< m1 >>
rect 487 235 488 236 
<< m1 >>
rect 523 235 524 236 
<< m1 >>
rect 19 236 20 237 
<< m1 >>
rect 22 236 23 237 
<< m1 >>
rect 55 236 56 237 
<< m2 >>
rect 56 236 57 237 
<< m1 >>
rect 85 236 86 237 
<< m1 >>
rect 100 236 101 237 
<< m1 >>
rect 118 236 119 237 
<< m1 >>
rect 127 236 128 237 
<< m1 >>
rect 148 236 149 237 
<< m1 >>
rect 163 236 164 237 
<< m1 >>
rect 172 236 173 237 
<< m1 >>
rect 175 236 176 237 
<< m1 >>
rect 176 236 177 237 
<< m1 >>
rect 177 236 178 237 
<< m1 >>
rect 178 236 179 237 
<< m1 >>
rect 179 236 180 237 
<< m2 >>
rect 179 236 180 237 
<< m2c >>
rect 179 236 180 237 
<< m1 >>
rect 179 236 180 237 
<< m2 >>
rect 179 236 180 237 
<< m2 >>
rect 180 236 181 237 
<< m1 >>
rect 181 236 182 237 
<< m2 >>
rect 181 236 182 237 
<< m2 >>
rect 182 236 183 237 
<< m1 >>
rect 183 236 184 237 
<< m2 >>
rect 183 236 184 237 
<< m2c >>
rect 183 236 184 237 
<< m1 >>
rect 183 236 184 237 
<< m2 >>
rect 183 236 184 237 
<< m1 >>
rect 184 236 185 237 
<< m1 >>
rect 185 236 186 237 
<< m2 >>
rect 186 236 187 237 
<< m1 >>
rect 190 236 191 237 
<< m1 >>
rect 194 236 195 237 
<< m2 >>
rect 194 236 195 237 
<< m2c >>
rect 194 236 195 237 
<< m1 >>
rect 194 236 195 237 
<< m2 >>
rect 194 236 195 237 
<< m1 >>
rect 195 236 196 237 
<< m1 >>
rect 196 236 197 237 
<< m1 >>
rect 197 236 198 237 
<< m1 >>
rect 198 236 199 237 
<< m1 >>
rect 199 236 200 237 
<< m1 >>
rect 207 236 208 237 
<< m2 >>
rect 207 236 208 237 
<< m2c >>
rect 207 236 208 237 
<< m1 >>
rect 207 236 208 237 
<< m2 >>
rect 207 236 208 237 
<< m2 >>
rect 217 236 218 237 
<< m1 >>
rect 221 236 222 237 
<< m2 >>
rect 221 236 222 237 
<< m2c >>
rect 221 236 222 237 
<< m1 >>
rect 221 236 222 237 
<< m2 >>
rect 221 236 222 237 
<< m1 >>
rect 226 236 227 237 
<< m2 >>
rect 226 236 227 237 
<< m2c >>
rect 226 236 227 237 
<< m1 >>
rect 226 236 227 237 
<< m2 >>
rect 226 236 227 237 
<< m1 >>
rect 229 236 230 237 
<< m2 >>
rect 229 236 230 237 
<< m2c >>
rect 229 236 230 237 
<< m1 >>
rect 229 236 230 237 
<< m2 >>
rect 229 236 230 237 
<< m1 >>
rect 233 236 234 237 
<< m1 >>
rect 235 236 236 237 
<< m1 >>
rect 237 236 238 237 
<< m1 >>
rect 240 236 241 237 
<< m1 >>
rect 272 236 273 237 
<< m1 >>
rect 284 236 285 237 
<< m2 >>
rect 284 236 285 237 
<< m2c >>
rect 284 236 285 237 
<< m1 >>
rect 284 236 285 237 
<< m2 >>
rect 284 236 285 237 
<< m1 >>
rect 285 236 286 237 
<< m1 >>
rect 286 236 287 237 
<< m1 >>
rect 287 236 288 237 
<< m1 >>
rect 288 236 289 237 
<< m1 >>
rect 289 236 290 237 
<< m1 >>
rect 290 236 291 237 
<< m1 >>
rect 292 236 293 237 
<< m2 >>
rect 292 236 293 237 
<< m2c >>
rect 292 236 293 237 
<< m1 >>
rect 292 236 293 237 
<< m2 >>
rect 292 236 293 237 
<< m1 >>
rect 296 236 297 237 
<< m1 >>
rect 298 236 299 237 
<< m1 >>
rect 301 236 302 237 
<< m1 >>
rect 302 236 303 237 
<< m1 >>
rect 303 236 304 237 
<< m1 >>
rect 304 236 305 237 
<< m1 >>
rect 305 236 306 237 
<< m1 >>
rect 307 236 308 237 
<< m1 >>
rect 316 236 317 237 
<< m1 >>
rect 337 236 338 237 
<< m1 >>
rect 352 236 353 237 
<< m1 >>
rect 379 236 380 237 
<< m2 >>
rect 380 236 381 237 
<< m1 >>
rect 383 236 384 237 
<< m1 >>
rect 394 236 395 237 
<< m1 >>
rect 416 236 417 237 
<< m1 >>
rect 419 236 420 237 
<< m1 >>
rect 421 236 422 237 
<< m2 >>
rect 422 236 423 237 
<< m1 >>
rect 434 236 435 237 
<< m1 >>
rect 442 236 443 237 
<< m1 >>
rect 478 236 479 237 
<< m1 >>
rect 487 236 488 237 
<< m1 >>
rect 523 236 524 237 
<< m1 >>
rect 19 237 20 238 
<< m1 >>
rect 22 237 23 238 
<< m1 >>
rect 55 237 56 238 
<< m2 >>
rect 56 237 57 238 
<< m1 >>
rect 85 237 86 238 
<< m1 >>
rect 100 237 101 238 
<< m1 >>
rect 118 237 119 238 
<< m1 >>
rect 127 237 128 238 
<< m1 >>
rect 148 237 149 238 
<< m1 >>
rect 163 237 164 238 
<< m1 >>
rect 172 237 173 238 
<< m1 >>
rect 181 237 182 238 
<< m2 >>
rect 186 237 187 238 
<< m1 >>
rect 190 237 191 238 
<< m2 >>
rect 194 237 195 238 
<< m2 >>
rect 207 237 208 238 
<< m2 >>
rect 217 237 218 238 
<< m2 >>
rect 221 237 222 238 
<< m2 >>
rect 226 237 227 238 
<< m2 >>
rect 229 237 230 238 
<< m2 >>
rect 230 237 231 238 
<< m2 >>
rect 231 237 232 238 
<< m2 >>
rect 232 237 233 238 
<< m1 >>
rect 233 237 234 238 
<< m2 >>
rect 233 237 234 238 
<< m2 >>
rect 234 237 235 238 
<< m1 >>
rect 235 237 236 238 
<< m2 >>
rect 235 237 236 238 
<< m2 >>
rect 236 237 237 238 
<< m1 >>
rect 237 237 238 238 
<< m2 >>
rect 237 237 238 238 
<< m2 >>
rect 238 237 239 238 
<< m1 >>
rect 239 237 240 238 
<< m2 >>
rect 239 237 240 238 
<< m2c >>
rect 239 237 240 238 
<< m1 >>
rect 239 237 240 238 
<< m2 >>
rect 239 237 240 238 
<< m1 >>
rect 240 237 241 238 
<< m1 >>
rect 272 237 273 238 
<< m2 >>
rect 284 237 285 238 
<< m2 >>
rect 292 237 293 238 
<< m1 >>
rect 296 237 297 238 
<< m1 >>
rect 298 237 299 238 
<< m1 >>
rect 307 237 308 238 
<< m2 >>
rect 308 237 309 238 
<< m1 >>
rect 309 237 310 238 
<< m2 >>
rect 309 237 310 238 
<< m2c >>
rect 309 237 310 238 
<< m1 >>
rect 309 237 310 238 
<< m2 >>
rect 309 237 310 238 
<< m1 >>
rect 310 237 311 238 
<< m1 >>
rect 311 237 312 238 
<< m1 >>
rect 312 237 313 238 
<< m1 >>
rect 313 237 314 238 
<< m1 >>
rect 314 237 315 238 
<< m1 >>
rect 315 237 316 238 
<< m1 >>
rect 316 237 317 238 
<< m1 >>
rect 337 237 338 238 
<< m1 >>
rect 352 237 353 238 
<< m1 >>
rect 379 237 380 238 
<< m2 >>
rect 380 237 381 238 
<< m1 >>
rect 383 237 384 238 
<< m1 >>
rect 394 237 395 238 
<< m1 >>
rect 416 237 417 238 
<< m1 >>
rect 419 237 420 238 
<< m1 >>
rect 421 237 422 238 
<< m2 >>
rect 422 237 423 238 
<< m1 >>
rect 434 237 435 238 
<< m1 >>
rect 442 237 443 238 
<< m1 >>
rect 478 237 479 238 
<< m1 >>
rect 487 237 488 238 
<< m1 >>
rect 523 237 524 238 
<< m1 >>
rect 19 238 20 239 
<< m1 >>
rect 22 238 23 239 
<< m1 >>
rect 55 238 56 239 
<< m2 >>
rect 56 238 57 239 
<< m1 >>
rect 64 238 65 239 
<< m1 >>
rect 65 238 66 239 
<< m1 >>
rect 66 238 67 239 
<< m1 >>
rect 67 238 68 239 
<< m1 >>
rect 68 238 69 239 
<< m1 >>
rect 69 238 70 239 
<< m1 >>
rect 70 238 71 239 
<< m1 >>
rect 71 238 72 239 
<< m1 >>
rect 72 238 73 239 
<< m1 >>
rect 73 238 74 239 
<< m1 >>
rect 74 238 75 239 
<< m1 >>
rect 75 238 76 239 
<< m1 >>
rect 76 238 77 239 
<< m1 >>
rect 77 238 78 239 
<< m1 >>
rect 78 238 79 239 
<< m1 >>
rect 79 238 80 239 
<< m1 >>
rect 80 238 81 239 
<< m1 >>
rect 81 238 82 239 
<< m1 >>
rect 82 238 83 239 
<< m1 >>
rect 83 238 84 239 
<< m1 >>
rect 84 238 85 239 
<< m1 >>
rect 85 238 86 239 
<< m1 >>
rect 100 238 101 239 
<< m1 >>
rect 118 238 119 239 
<< m1 >>
rect 127 238 128 239 
<< m1 >>
rect 148 238 149 239 
<< m1 >>
rect 163 238 164 239 
<< m1 >>
rect 172 238 173 239 
<< m1 >>
rect 181 238 182 239 
<< m2 >>
rect 186 238 187 239 
<< m1 >>
rect 190 238 191 239 
<< m1 >>
rect 193 238 194 239 
<< m1 >>
rect 194 238 195 239 
<< m2 >>
rect 194 238 195 239 
<< m1 >>
rect 195 238 196 239 
<< m1 >>
rect 196 238 197 239 
<< m1 >>
rect 197 238 198 239 
<< m1 >>
rect 198 238 199 239 
<< m1 >>
rect 199 238 200 239 
<< m1 >>
rect 200 238 201 239 
<< m1 >>
rect 201 238 202 239 
<< m1 >>
rect 202 238 203 239 
<< m1 >>
rect 203 238 204 239 
<< m1 >>
rect 204 238 205 239 
<< m1 >>
rect 205 238 206 239 
<< m1 >>
rect 206 238 207 239 
<< m1 >>
rect 207 238 208 239 
<< m2 >>
rect 207 238 208 239 
<< m1 >>
rect 208 238 209 239 
<< m1 >>
rect 209 238 210 239 
<< m2 >>
rect 209 238 210 239 
<< m2c >>
rect 209 238 210 239 
<< m1 >>
rect 209 238 210 239 
<< m2 >>
rect 209 238 210 239 
<< m2 >>
rect 210 238 211 239 
<< m1 >>
rect 211 238 212 239 
<< m2 >>
rect 211 238 212 239 
<< m1 >>
rect 212 238 213 239 
<< m2 >>
rect 212 238 213 239 
<< m1 >>
rect 213 238 214 239 
<< m2 >>
rect 213 238 214 239 
<< m1 >>
rect 214 238 215 239 
<< m2 >>
rect 214 238 215 239 
<< m1 >>
rect 215 238 216 239 
<< m2 >>
rect 215 238 216 239 
<< m1 >>
rect 216 238 217 239 
<< m2 >>
rect 216 238 217 239 
<< m1 >>
rect 217 238 218 239 
<< m2 >>
rect 217 238 218 239 
<< m1 >>
rect 218 238 219 239 
<< m1 >>
rect 219 238 220 239 
<< m1 >>
rect 220 238 221 239 
<< m1 >>
rect 221 238 222 239 
<< m2 >>
rect 221 238 222 239 
<< m1 >>
rect 222 238 223 239 
<< m1 >>
rect 223 238 224 239 
<< m1 >>
rect 224 238 225 239 
<< m1 >>
rect 225 238 226 239 
<< m1 >>
rect 226 238 227 239 
<< m2 >>
rect 226 238 227 239 
<< m1 >>
rect 227 238 228 239 
<< m1 >>
rect 228 238 229 239 
<< m1 >>
rect 229 238 230 239 
<< m1 >>
rect 230 238 231 239 
<< m1 >>
rect 231 238 232 239 
<< m1 >>
rect 232 238 233 239 
<< m1 >>
rect 233 238 234 239 
<< m1 >>
rect 235 238 236 239 
<< m1 >>
rect 237 238 238 239 
<< m1 >>
rect 272 238 273 239 
<< m1 >>
rect 276 238 277 239 
<< m1 >>
rect 277 238 278 239 
<< m1 >>
rect 278 238 279 239 
<< m1 >>
rect 279 238 280 239 
<< m1 >>
rect 280 238 281 239 
<< m1 >>
rect 281 238 282 239 
<< m1 >>
rect 282 238 283 239 
<< m1 >>
rect 283 238 284 239 
<< m1 >>
rect 284 238 285 239 
<< m2 >>
rect 284 238 285 239 
<< m1 >>
rect 285 238 286 239 
<< m1 >>
rect 286 238 287 239 
<< m1 >>
rect 287 238 288 239 
<< m1 >>
rect 288 238 289 239 
<< m1 >>
rect 289 238 290 239 
<< m1 >>
rect 290 238 291 239 
<< m1 >>
rect 291 238 292 239 
<< m1 >>
rect 292 238 293 239 
<< m2 >>
rect 292 238 293 239 
<< m1 >>
rect 293 238 294 239 
<< m1 >>
rect 294 238 295 239 
<< m1 >>
rect 295 238 296 239 
<< m1 >>
rect 296 238 297 239 
<< m1 >>
rect 298 238 299 239 
<< m1 >>
rect 307 238 308 239 
<< m2 >>
rect 308 238 309 239 
<< m1 >>
rect 337 238 338 239 
<< m1 >>
rect 352 238 353 239 
<< m1 >>
rect 379 238 380 239 
<< m2 >>
rect 380 238 381 239 
<< m1 >>
rect 383 238 384 239 
<< m1 >>
rect 384 238 385 239 
<< m1 >>
rect 385 238 386 239 
<< m1 >>
rect 386 238 387 239 
<< m1 >>
rect 387 238 388 239 
<< m1 >>
rect 388 238 389 239 
<< m1 >>
rect 389 238 390 239 
<< m1 >>
rect 390 238 391 239 
<< m1 >>
rect 391 238 392 239 
<< m1 >>
rect 392 238 393 239 
<< m1 >>
rect 393 238 394 239 
<< m1 >>
rect 394 238 395 239 
<< m1 >>
rect 416 238 417 239 
<< m1 >>
rect 419 238 420 239 
<< m1 >>
rect 421 238 422 239 
<< m2 >>
rect 422 238 423 239 
<< m1 >>
rect 434 238 435 239 
<< m1 >>
rect 442 238 443 239 
<< m2 >>
rect 442 238 443 239 
<< m2 >>
rect 443 238 444 239 
<< m1 >>
rect 444 238 445 239 
<< m2 >>
rect 444 238 445 239 
<< m2c >>
rect 444 238 445 239 
<< m1 >>
rect 444 238 445 239 
<< m2 >>
rect 444 238 445 239 
<< m1 >>
rect 445 238 446 239 
<< m1 >>
rect 446 238 447 239 
<< m1 >>
rect 447 238 448 239 
<< m1 >>
rect 448 238 449 239 
<< m1 >>
rect 449 238 450 239 
<< m1 >>
rect 450 238 451 239 
<< m1 >>
rect 451 238 452 239 
<< m1 >>
rect 452 238 453 239 
<< m1 >>
rect 453 238 454 239 
<< m1 >>
rect 454 238 455 239 
<< m1 >>
rect 455 238 456 239 
<< m1 >>
rect 456 238 457 239 
<< m1 >>
rect 457 238 458 239 
<< m1 >>
rect 458 238 459 239 
<< m1 >>
rect 459 238 460 239 
<< m1 >>
rect 460 238 461 239 
<< m1 >>
rect 461 238 462 239 
<< m1 >>
rect 462 238 463 239 
<< m1 >>
rect 463 238 464 239 
<< m1 >>
rect 464 238 465 239 
<< m1 >>
rect 465 238 466 239 
<< m1 >>
rect 466 238 467 239 
<< m1 >>
rect 467 238 468 239 
<< m1 >>
rect 468 238 469 239 
<< m1 >>
rect 469 238 470 239 
<< m1 >>
rect 470 238 471 239 
<< m1 >>
rect 471 238 472 239 
<< m1 >>
rect 472 238 473 239 
<< m1 >>
rect 473 238 474 239 
<< m1 >>
rect 474 238 475 239 
<< m1 >>
rect 475 238 476 239 
<< m1 >>
rect 476 238 477 239 
<< m1 >>
rect 477 238 478 239 
<< m1 >>
rect 478 238 479 239 
<< m1 >>
rect 487 238 488 239 
<< m1 >>
rect 523 238 524 239 
<< m1 >>
rect 19 239 20 240 
<< m1 >>
rect 22 239 23 240 
<< m1 >>
rect 55 239 56 240 
<< m2 >>
rect 56 239 57 240 
<< m1 >>
rect 64 239 65 240 
<< m1 >>
rect 100 239 101 240 
<< m1 >>
rect 118 239 119 240 
<< m1 >>
rect 127 239 128 240 
<< m1 >>
rect 148 239 149 240 
<< m1 >>
rect 163 239 164 240 
<< m1 >>
rect 172 239 173 240 
<< m2 >>
rect 180 239 181 240 
<< m1 >>
rect 181 239 182 240 
<< m2 >>
rect 181 239 182 240 
<< m2 >>
rect 182 239 183 240 
<< m1 >>
rect 183 239 184 240 
<< m2 >>
rect 183 239 184 240 
<< m2c >>
rect 183 239 184 240 
<< m1 >>
rect 183 239 184 240 
<< m2 >>
rect 183 239 184 240 
<< m1 >>
rect 184 239 185 240 
<< m1 >>
rect 185 239 186 240 
<< m1 >>
rect 186 239 187 240 
<< m2 >>
rect 186 239 187 240 
<< m1 >>
rect 187 239 188 240 
<< m1 >>
rect 188 239 189 240 
<< m2 >>
rect 188 239 189 240 
<< m2c >>
rect 188 239 189 240 
<< m1 >>
rect 188 239 189 240 
<< m2 >>
rect 188 239 189 240 
<< m2 >>
rect 189 239 190 240 
<< m1 >>
rect 190 239 191 240 
<< m2 >>
rect 190 239 191 240 
<< m2 >>
rect 191 239 192 240 
<< m2 >>
rect 192 239 193 240 
<< m1 >>
rect 193 239 194 240 
<< m2 >>
rect 193 239 194 240 
<< m2 >>
rect 194 239 195 240 
<< m2 >>
rect 207 239 208 240 
<< m1 >>
rect 211 239 212 240 
<< m2 >>
rect 221 239 222 240 
<< m2 >>
rect 226 239 227 240 
<< m1 >>
rect 235 239 236 240 
<< m1 >>
rect 237 239 238 240 
<< m1 >>
rect 272 239 273 240 
<< m2 >>
rect 272 239 273 240 
<< m2c >>
rect 272 239 273 240 
<< m1 >>
rect 272 239 273 240 
<< m2 >>
rect 272 239 273 240 
<< m2 >>
rect 275 239 276 240 
<< m1 >>
rect 276 239 277 240 
<< m2 >>
rect 276 239 277 240 
<< m2 >>
rect 277 239 278 240 
<< m2 >>
rect 278 239 279 240 
<< m2 >>
rect 279 239 280 240 
<< m2 >>
rect 280 239 281 240 
<< m2 >>
rect 281 239 282 240 
<< m2 >>
rect 282 239 283 240 
<< m2 >>
rect 283 239 284 240 
<< m2 >>
rect 284 239 285 240 
<< m2 >>
rect 292 239 293 240 
<< m1 >>
rect 298 239 299 240 
<< m1 >>
rect 307 239 308 240 
<< m2 >>
rect 308 239 309 240 
<< m1 >>
rect 337 239 338 240 
<< m1 >>
rect 352 239 353 240 
<< m1 >>
rect 379 239 380 240 
<< m2 >>
rect 380 239 381 240 
<< m1 >>
rect 416 239 417 240 
<< m1 >>
rect 419 239 420 240 
<< m1 >>
rect 421 239 422 240 
<< m2 >>
rect 422 239 423 240 
<< m1 >>
rect 434 239 435 240 
<< m1 >>
rect 442 239 443 240 
<< m2 >>
rect 442 239 443 240 
<< m1 >>
rect 487 239 488 240 
<< m1 >>
rect 523 239 524 240 
<< m1 >>
rect 19 240 20 241 
<< m1 >>
rect 22 240 23 241 
<< m1 >>
rect 55 240 56 241 
<< m2 >>
rect 56 240 57 241 
<< m1 >>
rect 64 240 65 241 
<< m1 >>
rect 100 240 101 241 
<< m1 >>
rect 118 240 119 241 
<< m1 >>
rect 127 240 128 241 
<< m1 >>
rect 148 240 149 241 
<< m1 >>
rect 163 240 164 241 
<< m1 >>
rect 172 240 173 241 
<< m2 >>
rect 180 240 181 241 
<< m1 >>
rect 181 240 182 241 
<< m2 >>
rect 186 240 187 241 
<< m1 >>
rect 190 240 191 241 
<< m1 >>
rect 193 240 194 241 
<< m1 >>
rect 207 240 208 241 
<< m2 >>
rect 207 240 208 241 
<< m2c >>
rect 207 240 208 241 
<< m1 >>
rect 207 240 208 241 
<< m2 >>
rect 207 240 208 241 
<< m1 >>
rect 211 240 212 241 
<< m1 >>
rect 221 240 222 241 
<< m2 >>
rect 221 240 222 241 
<< m2c >>
rect 221 240 222 241 
<< m1 >>
rect 221 240 222 241 
<< m2 >>
rect 221 240 222 241 
<< m1 >>
rect 226 240 227 241 
<< m2 >>
rect 226 240 227 241 
<< m2c >>
rect 226 240 227 241 
<< m1 >>
rect 226 240 227 241 
<< m2 >>
rect 226 240 227 241 
<< m1 >>
rect 235 240 236 241 
<< m1 >>
rect 237 240 238 241 
<< m2 >>
rect 272 240 273 241 
<< m2 >>
rect 275 240 276 241 
<< m1 >>
rect 276 240 277 241 
<< m2 >>
rect 292 240 293 241 
<< m1 >>
rect 296 240 297 241 
<< m2 >>
rect 296 240 297 241 
<< m2c >>
rect 296 240 297 241 
<< m1 >>
rect 296 240 297 241 
<< m2 >>
rect 296 240 297 241 
<< m2 >>
rect 297 240 298 241 
<< m1 >>
rect 298 240 299 241 
<< m2 >>
rect 298 240 299 241 
<< m2 >>
rect 299 240 300 241 
<< m2 >>
rect 300 240 301 241 
<< m2 >>
rect 301 240 302 241 
<< m2 >>
rect 302 240 303 241 
<< m2 >>
rect 303 240 304 241 
<< m2 >>
rect 304 240 305 241 
<< m2 >>
rect 305 240 306 241 
<< m2 >>
rect 306 240 307 241 
<< m1 >>
rect 307 240 308 241 
<< m2 >>
rect 307 240 308 241 
<< m2 >>
rect 308 240 309 241 
<< m1 >>
rect 337 240 338 241 
<< m1 >>
rect 352 240 353 241 
<< m1 >>
rect 379 240 380 241 
<< m2 >>
rect 380 240 381 241 
<< m1 >>
rect 416 240 417 241 
<< m1 >>
rect 419 240 420 241 
<< m1 >>
rect 421 240 422 241 
<< m2 >>
rect 422 240 423 241 
<< m1 >>
rect 434 240 435 241 
<< m1 >>
rect 442 240 443 241 
<< m2 >>
rect 442 240 443 241 
<< m1 >>
rect 487 240 488 241 
<< m1 >>
rect 523 240 524 241 
<< m1 >>
rect 19 241 20 242 
<< m1 >>
rect 22 241 23 242 
<< m1 >>
rect 44 241 45 242 
<< m1 >>
rect 45 241 46 242 
<< m1 >>
rect 46 241 47 242 
<< m1 >>
rect 47 241 48 242 
<< m1 >>
rect 48 241 49 242 
<< m1 >>
rect 49 241 50 242 
<< m1 >>
rect 50 241 51 242 
<< m1 >>
rect 51 241 52 242 
<< m1 >>
rect 52 241 53 242 
<< m1 >>
rect 55 241 56 242 
<< m2 >>
rect 56 241 57 242 
<< m1 >>
rect 64 241 65 242 
<< m1 >>
rect 100 241 101 242 
<< m1 >>
rect 101 241 102 242 
<< m1 >>
rect 102 241 103 242 
<< m1 >>
rect 103 241 104 242 
<< m1 >>
rect 104 241 105 242 
<< m1 >>
rect 105 241 106 242 
<< m1 >>
rect 106 241 107 242 
<< m1 >>
rect 118 241 119 242 
<< m1 >>
rect 127 241 128 242 
<< m1 >>
rect 148 241 149 242 
<< m1 >>
rect 163 241 164 242 
<< m1 >>
rect 172 241 173 242 
<< m1 >>
rect 174 241 175 242 
<< m1 >>
rect 175 241 176 242 
<< m1 >>
rect 176 241 177 242 
<< m1 >>
rect 177 241 178 242 
<< m1 >>
rect 178 241 179 242 
<< m1 >>
rect 179 241 180 242 
<< m2 >>
rect 179 241 180 242 
<< m2c >>
rect 179 241 180 242 
<< m1 >>
rect 179 241 180 242 
<< m2 >>
rect 179 241 180 242 
<< m2 >>
rect 180 241 181 242 
<< m1 >>
rect 181 241 182 242 
<< m2 >>
rect 182 241 183 242 
<< m1 >>
rect 183 241 184 242 
<< m2 >>
rect 183 241 184 242 
<< m2c >>
rect 183 241 184 242 
<< m1 >>
rect 183 241 184 242 
<< m2 >>
rect 183 241 184 242 
<< m1 >>
rect 184 241 185 242 
<< m1 >>
rect 185 241 186 242 
<< m1 >>
rect 186 241 187 242 
<< m2 >>
rect 186 241 187 242 
<< m1 >>
rect 187 241 188 242 
<< m1 >>
rect 188 241 189 242 
<< m2 >>
rect 188 241 189 242 
<< m2c >>
rect 188 241 189 242 
<< m1 >>
rect 188 241 189 242 
<< m2 >>
rect 188 241 189 242 
<< m2 >>
rect 189 241 190 242 
<< m1 >>
rect 190 241 191 242 
<< m2 >>
rect 190 241 191 242 
<< m2 >>
rect 191 241 192 242 
<< m2 >>
rect 192 241 193 242 
<< m1 >>
rect 193 241 194 242 
<< m2 >>
rect 193 241 194 242 
<< m2 >>
rect 194 241 195 242 
<< m1 >>
rect 207 241 208 242 
<< m1 >>
rect 209 241 210 242 
<< m2 >>
rect 209 241 210 242 
<< m2c >>
rect 209 241 210 242 
<< m1 >>
rect 209 241 210 242 
<< m2 >>
rect 209 241 210 242 
<< m2 >>
rect 210 241 211 242 
<< m1 >>
rect 211 241 212 242 
<< m2 >>
rect 211 241 212 242 
<< m2 >>
rect 212 241 213 242 
<< m1 >>
rect 221 241 222 242 
<< m2 >>
rect 221 241 222 242 
<< m1 >>
rect 226 241 227 242 
<< m1 >>
rect 228 241 229 242 
<< m1 >>
rect 229 241 230 242 
<< m1 >>
rect 230 241 231 242 
<< m1 >>
rect 231 241 232 242 
<< m1 >>
rect 232 241 233 242 
<< m1 >>
rect 233 241 234 242 
<< m2 >>
rect 233 241 234 242 
<< m2c >>
rect 233 241 234 242 
<< m1 >>
rect 233 241 234 242 
<< m2 >>
rect 233 241 234 242 
<< m2 >>
rect 234 241 235 242 
<< m1 >>
rect 235 241 236 242 
<< m2 >>
rect 235 241 236 242 
<< m2 >>
rect 236 241 237 242 
<< m1 >>
rect 237 241 238 242 
<< m2 >>
rect 237 241 238 242 
<< m2 >>
rect 238 241 239 242 
<< m1 >>
rect 239 241 240 242 
<< m2 >>
rect 239 241 240 242 
<< m2c >>
rect 239 241 240 242 
<< m1 >>
rect 239 241 240 242 
<< m2 >>
rect 239 241 240 242 
<< m1 >>
rect 240 241 241 242 
<< m1 >>
rect 241 241 242 242 
<< m1 >>
rect 242 241 243 242 
<< m1 >>
rect 243 241 244 242 
<< m1 >>
rect 244 241 245 242 
<< m1 >>
rect 245 241 246 242 
<< m1 >>
rect 246 241 247 242 
<< m1 >>
rect 247 241 248 242 
<< m1 >>
rect 248 241 249 242 
<< m1 >>
rect 249 241 250 242 
<< m1 >>
rect 262 241 263 242 
<< m1 >>
rect 263 241 264 242 
<< m1 >>
rect 264 241 265 242 
<< m1 >>
rect 265 241 266 242 
<< m1 >>
rect 266 241 267 242 
<< m1 >>
rect 267 241 268 242 
<< m1 >>
rect 268 241 269 242 
<< m1 >>
rect 269 241 270 242 
<< m1 >>
rect 270 241 271 242 
<< m1 >>
rect 271 241 272 242 
<< m1 >>
rect 272 241 273 242 
<< m2 >>
rect 272 241 273 242 
<< m1 >>
rect 273 241 274 242 
<< m1 >>
rect 274 241 275 242 
<< m2 >>
rect 274 241 275 242 
<< m2c >>
rect 274 241 275 242 
<< m1 >>
rect 274 241 275 242 
<< m2 >>
rect 274 241 275 242 
<< m2 >>
rect 275 241 276 242 
<< m1 >>
rect 276 241 277 242 
<< m2 >>
rect 277 241 278 242 
<< m1 >>
rect 278 241 279 242 
<< m2 >>
rect 278 241 279 242 
<< m2c >>
rect 278 241 279 242 
<< m1 >>
rect 278 241 279 242 
<< m2 >>
rect 278 241 279 242 
<< m1 >>
rect 279 241 280 242 
<< m1 >>
rect 280 241 281 242 
<< m1 >>
rect 281 241 282 242 
<< m1 >>
rect 282 241 283 242 
<< m1 >>
rect 283 241 284 242 
<< m1 >>
rect 284 241 285 242 
<< m1 >>
rect 285 241 286 242 
<< m1 >>
rect 286 241 287 242 
<< m1 >>
rect 287 241 288 242 
<< m1 >>
rect 288 241 289 242 
<< m1 >>
rect 289 241 290 242 
<< m1 >>
rect 290 241 291 242 
<< m1 >>
rect 291 241 292 242 
<< m1 >>
rect 292 241 293 242 
<< m2 >>
rect 292 241 293 242 
<< m1 >>
rect 293 241 294 242 
<< m1 >>
rect 294 241 295 242 
<< m1 >>
rect 295 241 296 242 
<< m1 >>
rect 296 241 297 242 
<< m1 >>
rect 298 241 299 242 
<< m1 >>
rect 299 241 300 242 
<< m1 >>
rect 300 241 301 242 
<< m1 >>
rect 301 241 302 242 
<< m1 >>
rect 302 241 303 242 
<< m1 >>
rect 303 241 304 242 
<< m1 >>
rect 304 241 305 242 
<< m1 >>
rect 305 241 306 242 
<< m1 >>
rect 307 241 308 242 
<< m1 >>
rect 337 241 338 242 
<< m1 >>
rect 338 241 339 242 
<< m1 >>
rect 339 241 340 242 
<< m1 >>
rect 340 241 341 242 
<< m1 >>
rect 341 241 342 242 
<< m1 >>
rect 342 241 343 242 
<< m1 >>
rect 343 241 344 242 
<< m1 >>
rect 344 241 345 242 
<< m1 >>
rect 345 241 346 242 
<< m1 >>
rect 346 241 347 242 
<< m1 >>
rect 352 241 353 242 
<< m1 >>
rect 379 241 380 242 
<< m2 >>
rect 380 241 381 242 
<< m1 >>
rect 416 241 417 242 
<< m1 >>
rect 419 241 420 242 
<< m1 >>
rect 421 241 422 242 
<< m2 >>
rect 422 241 423 242 
<< m1 >>
rect 434 241 435 242 
<< m1 >>
rect 442 241 443 242 
<< m2 >>
rect 442 241 443 242 
<< m1 >>
rect 487 241 488 242 
<< m1 >>
rect 523 241 524 242 
<< m1 >>
rect 19 242 20 243 
<< m1 >>
rect 22 242 23 243 
<< m1 >>
rect 44 242 45 243 
<< m1 >>
rect 52 242 53 243 
<< m1 >>
rect 55 242 56 243 
<< m2 >>
rect 56 242 57 243 
<< m1 >>
rect 64 242 65 243 
<< m1 >>
rect 106 242 107 243 
<< m1 >>
rect 118 242 119 243 
<< m1 >>
rect 127 242 128 243 
<< m1 >>
rect 148 242 149 243 
<< m1 >>
rect 163 242 164 243 
<< m1 >>
rect 172 242 173 243 
<< m1 >>
rect 174 242 175 243 
<< m1 >>
rect 181 242 182 243 
<< m2 >>
rect 182 242 183 243 
<< m2 >>
rect 186 242 187 243 
<< m1 >>
rect 190 242 191 243 
<< m1 >>
rect 193 242 194 243 
<< m2 >>
rect 194 242 195 243 
<< m1 >>
rect 195 242 196 243 
<< m2 >>
rect 195 242 196 243 
<< m2c >>
rect 195 242 196 243 
<< m1 >>
rect 195 242 196 243 
<< m2 >>
rect 195 242 196 243 
<< m1 >>
rect 196 242 197 243 
<< m1 >>
rect 197 242 198 243 
<< m1 >>
rect 198 242 199 243 
<< m1 >>
rect 199 242 200 243 
<< m1 >>
rect 200 242 201 243 
<< m1 >>
rect 201 242 202 243 
<< m1 >>
rect 202 242 203 243 
<< m1 >>
rect 203 242 204 243 
<< m1 >>
rect 204 242 205 243 
<< m1 >>
rect 205 242 206 243 
<< m2 >>
rect 205 242 206 243 
<< m2c >>
rect 205 242 206 243 
<< m1 >>
rect 205 242 206 243 
<< m2 >>
rect 205 242 206 243 
<< m2 >>
rect 206 242 207 243 
<< m1 >>
rect 207 242 208 243 
<< m2 >>
rect 207 242 208 243 
<< m2 >>
rect 208 242 209 243 
<< m1 >>
rect 209 242 210 243 
<< m2 >>
rect 209 242 210 243 
<< m1 >>
rect 211 242 212 243 
<< m2 >>
rect 212 242 213 243 
<< m2 >>
rect 221 242 222 243 
<< m2 >>
rect 222 242 223 243 
<< m2 >>
rect 223 242 224 243 
<< m2 >>
rect 224 242 225 243 
<< m2 >>
rect 225 242 226 243 
<< m1 >>
rect 226 242 227 243 
<< m2 >>
rect 226 242 227 243 
<< m2 >>
rect 227 242 228 243 
<< m1 >>
rect 228 242 229 243 
<< m2 >>
rect 228 242 229 243 
<< m2c >>
rect 228 242 229 243 
<< m1 >>
rect 228 242 229 243 
<< m2 >>
rect 228 242 229 243 
<< m1 >>
rect 235 242 236 243 
<< m1 >>
rect 237 242 238 243 
<< m1 >>
rect 249 242 250 243 
<< m2 >>
rect 249 242 250 243 
<< m2c >>
rect 249 242 250 243 
<< m1 >>
rect 249 242 250 243 
<< m2 >>
rect 249 242 250 243 
<< m1 >>
rect 262 242 263 243 
<< m2 >>
rect 262 242 263 243 
<< m2c >>
rect 262 242 263 243 
<< m1 >>
rect 262 242 263 243 
<< m2 >>
rect 262 242 263 243 
<< m2 >>
rect 272 242 273 243 
<< m1 >>
rect 276 242 277 243 
<< m2 >>
rect 277 242 278 243 
<< m2 >>
rect 292 242 293 243 
<< m1 >>
rect 305 242 306 243 
<< m1 >>
rect 307 242 308 243 
<< m1 >>
rect 346 242 347 243 
<< m1 >>
rect 352 242 353 243 
<< m1 >>
rect 379 242 380 243 
<< m2 >>
rect 380 242 381 243 
<< m1 >>
rect 416 242 417 243 
<< m1 >>
rect 419 242 420 243 
<< m1 >>
rect 421 242 422 243 
<< m2 >>
rect 422 242 423 243 
<< m1 >>
rect 434 242 435 243 
<< m1 >>
rect 442 242 443 243 
<< m2 >>
rect 442 242 443 243 
<< m1 >>
rect 487 242 488 243 
<< m1 >>
rect 523 242 524 243 
<< m1 >>
rect 19 243 20 244 
<< m1 >>
rect 22 243 23 244 
<< m1 >>
rect 44 243 45 244 
<< m1 >>
rect 52 243 53 244 
<< m1 >>
rect 55 243 56 244 
<< m2 >>
rect 56 243 57 244 
<< m1 >>
rect 64 243 65 244 
<< m1 >>
rect 106 243 107 244 
<< m1 >>
rect 118 243 119 244 
<< m1 >>
rect 127 243 128 244 
<< m1 >>
rect 148 243 149 244 
<< m1 >>
rect 163 243 164 244 
<< m1 >>
rect 172 243 173 244 
<< m1 >>
rect 174 243 175 244 
<< m1 >>
rect 181 243 182 244 
<< m2 >>
rect 182 243 183 244 
<< m1 >>
rect 186 243 187 244 
<< m2 >>
rect 186 243 187 244 
<< m2c >>
rect 186 243 187 244 
<< m1 >>
rect 186 243 187 244 
<< m2 >>
rect 186 243 187 244 
<< m1 >>
rect 190 243 191 244 
<< m1 >>
rect 193 243 194 244 
<< m1 >>
rect 207 243 208 244 
<< m1 >>
rect 211 243 212 244 
<< m2 >>
rect 212 243 213 244 
<< m1 >>
rect 213 243 214 244 
<< m2 >>
rect 213 243 214 244 
<< m2c >>
rect 213 243 214 244 
<< m1 >>
rect 213 243 214 244 
<< m2 >>
rect 213 243 214 244 
<< m1 >>
rect 214 243 215 244 
<< m1 >>
rect 215 243 216 244 
<< m1 >>
rect 216 243 217 244 
<< m1 >>
rect 217 243 218 244 
<< m1 >>
rect 218 243 219 244 
<< m1 >>
rect 219 243 220 244 
<< m1 >>
rect 220 243 221 244 
<< m1 >>
rect 221 243 222 244 
<< m1 >>
rect 222 243 223 244 
<< m1 >>
rect 223 243 224 244 
<< m1 >>
rect 224 243 225 244 
<< m1 >>
rect 226 243 227 244 
<< m1 >>
rect 235 243 236 244 
<< m1 >>
rect 237 243 238 244 
<< m2 >>
rect 249 243 250 244 
<< m2 >>
rect 250 243 251 244 
<< m2 >>
rect 251 243 252 244 
<< m2 >>
rect 252 243 253 244 
<< m2 >>
rect 253 243 254 244 
<< m2 >>
rect 262 243 263 244 
<< m1 >>
rect 272 243 273 244 
<< m2 >>
rect 272 243 273 244 
<< m2c >>
rect 272 243 273 244 
<< m1 >>
rect 272 243 273 244 
<< m2 >>
rect 272 243 273 244 
<< m1 >>
rect 273 243 274 244 
<< m1 >>
rect 274 243 275 244 
<< m2 >>
rect 274 243 275 244 
<< m2c >>
rect 274 243 275 244 
<< m1 >>
rect 274 243 275 244 
<< m2 >>
rect 274 243 275 244 
<< m2 >>
rect 275 243 276 244 
<< m1 >>
rect 276 243 277 244 
<< m2 >>
rect 276 243 277 244 
<< m2 >>
rect 277 243 278 244 
<< m1 >>
rect 292 243 293 244 
<< m2 >>
rect 292 243 293 244 
<< m2c >>
rect 292 243 293 244 
<< m1 >>
rect 292 243 293 244 
<< m2 >>
rect 292 243 293 244 
<< m1 >>
rect 305 243 306 244 
<< m1 >>
rect 307 243 308 244 
<< m1 >>
rect 346 243 347 244 
<< m1 >>
rect 352 243 353 244 
<< m1 >>
rect 379 243 380 244 
<< m2 >>
rect 380 243 381 244 
<< m1 >>
rect 416 243 417 244 
<< m1 >>
rect 419 243 420 244 
<< m1 >>
rect 421 243 422 244 
<< m2 >>
rect 422 243 423 244 
<< m1 >>
rect 434 243 435 244 
<< m1 >>
rect 442 243 443 244 
<< m2 >>
rect 442 243 443 244 
<< m1 >>
rect 481 243 482 244 
<< m1 >>
rect 482 243 483 244 
<< m1 >>
rect 483 243 484 244 
<< m1 >>
rect 484 243 485 244 
<< m1 >>
rect 485 243 486 244 
<< m1 >>
rect 486 243 487 244 
<< m1 >>
rect 487 243 488 244 
<< m1 >>
rect 523 243 524 244 
<< m1 >>
rect 19 244 20 245 
<< m1 >>
rect 22 244 23 245 
<< m1 >>
rect 44 244 45 245 
<< m1 >>
rect 52 244 53 245 
<< m1 >>
rect 55 244 56 245 
<< m2 >>
rect 56 244 57 245 
<< m1 >>
rect 64 244 65 245 
<< m1 >>
rect 106 244 107 245 
<< m1 >>
rect 118 244 119 245 
<< m1 >>
rect 127 244 128 245 
<< m1 >>
rect 148 244 149 245 
<< m1 >>
rect 163 244 164 245 
<< m2 >>
rect 171 244 172 245 
<< m1 >>
rect 172 244 173 245 
<< m2 >>
rect 172 244 173 245 
<< m2 >>
rect 173 244 174 245 
<< m1 >>
rect 174 244 175 245 
<< m2 >>
rect 174 244 175 245 
<< m2c >>
rect 174 244 175 245 
<< m1 >>
rect 174 244 175 245 
<< m2 >>
rect 174 244 175 245 
<< m1 >>
rect 181 244 182 245 
<< m2 >>
rect 182 244 183 245 
<< m1 >>
rect 186 244 187 245 
<< m1 >>
rect 190 244 191 245 
<< m1 >>
rect 193 244 194 245 
<< m1 >>
rect 207 244 208 245 
<< m1 >>
rect 211 244 212 245 
<< m1 >>
rect 224 244 225 245 
<< m1 >>
rect 226 244 227 245 
<< m1 >>
rect 235 244 236 245 
<< m1 >>
rect 237 244 238 245 
<< m1 >>
rect 250 244 251 245 
<< m1 >>
rect 251 244 252 245 
<< m1 >>
rect 252 244 253 245 
<< m1 >>
rect 253 244 254 245 
<< m2 >>
rect 253 244 254 245 
<< m1 >>
rect 254 244 255 245 
<< m1 >>
rect 255 244 256 245 
<< m1 >>
rect 256 244 257 245 
<< m1 >>
rect 257 244 258 245 
<< m1 >>
rect 258 244 259 245 
<< m1 >>
rect 259 244 260 245 
<< m1 >>
rect 260 244 261 245 
<< m1 >>
rect 261 244 262 245 
<< m1 >>
rect 262 244 263 245 
<< m2 >>
rect 262 244 263 245 
<< m1 >>
rect 276 244 277 245 
<< m1 >>
rect 292 244 293 245 
<< m1 >>
rect 305 244 306 245 
<< m2 >>
rect 305 244 306 245 
<< m2c >>
rect 305 244 306 245 
<< m1 >>
rect 305 244 306 245 
<< m2 >>
rect 305 244 306 245 
<< m2 >>
rect 306 244 307 245 
<< m1 >>
rect 307 244 308 245 
<< m2 >>
rect 307 244 308 245 
<< m2 >>
rect 308 244 309 245 
<< m1 >>
rect 334 244 335 245 
<< m1 >>
rect 335 244 336 245 
<< m1 >>
rect 336 244 337 245 
<< m1 >>
rect 337 244 338 245 
<< m1 >>
rect 346 244 347 245 
<< m1 >>
rect 352 244 353 245 
<< m1 >>
rect 379 244 380 245 
<< m2 >>
rect 380 244 381 245 
<< m1 >>
rect 416 244 417 245 
<< m1 >>
rect 419 244 420 245 
<< m1 >>
rect 421 244 422 245 
<< m2 >>
rect 422 244 423 245 
<< m1 >>
rect 434 244 435 245 
<< m1 >>
rect 442 244 443 245 
<< m2 >>
rect 442 244 443 245 
<< m1 >>
rect 481 244 482 245 
<< m1 >>
rect 496 244 497 245 
<< m1 >>
rect 497 244 498 245 
<< m1 >>
rect 498 244 499 245 
<< m1 >>
rect 499 244 500 245 
<< m1 >>
rect 523 244 524 245 
<< m1 >>
rect 19 245 20 246 
<< m1 >>
rect 22 245 23 246 
<< m1 >>
rect 44 245 45 246 
<< m1 >>
rect 52 245 53 246 
<< m1 >>
rect 55 245 56 246 
<< m2 >>
rect 56 245 57 246 
<< m1 >>
rect 64 245 65 246 
<< m1 >>
rect 106 245 107 246 
<< m1 >>
rect 118 245 119 246 
<< m1 >>
rect 127 245 128 246 
<< m1 >>
rect 148 245 149 246 
<< m1 >>
rect 163 245 164 246 
<< m2 >>
rect 171 245 172 246 
<< m1 >>
rect 172 245 173 246 
<< m1 >>
rect 181 245 182 246 
<< m2 >>
rect 182 245 183 246 
<< m1 >>
rect 186 245 187 246 
<< m1 >>
rect 190 245 191 246 
<< m1 >>
rect 193 245 194 246 
<< m1 >>
rect 207 245 208 246 
<< m1 >>
rect 211 245 212 246 
<< m1 >>
rect 224 245 225 246 
<< m1 >>
rect 226 245 227 246 
<< m1 >>
rect 235 245 236 246 
<< m1 >>
rect 237 245 238 246 
<< m1 >>
rect 250 245 251 246 
<< m2 >>
rect 253 245 254 246 
<< m1 >>
rect 262 245 263 246 
<< m2 >>
rect 262 245 263 246 
<< m1 >>
rect 274 245 275 246 
<< m2 >>
rect 274 245 275 246 
<< m2c >>
rect 274 245 275 246 
<< m1 >>
rect 274 245 275 246 
<< m2 >>
rect 274 245 275 246 
<< m2 >>
rect 275 245 276 246 
<< m1 >>
rect 276 245 277 246 
<< m2 >>
rect 276 245 277 246 
<< m2 >>
rect 277 245 278 246 
<< m1 >>
rect 278 245 279 246 
<< m2 >>
rect 278 245 279 246 
<< m2c >>
rect 278 245 279 246 
<< m1 >>
rect 278 245 279 246 
<< m2 >>
rect 278 245 279 246 
<< m1 >>
rect 279 245 280 246 
<< m1 >>
rect 280 245 281 246 
<< m1 >>
rect 281 245 282 246 
<< m1 >>
rect 282 245 283 246 
<< m1 >>
rect 283 245 284 246 
<< m1 >>
rect 284 245 285 246 
<< m1 >>
rect 285 245 286 246 
<< m1 >>
rect 286 245 287 246 
<< m1 >>
rect 287 245 288 246 
<< m1 >>
rect 288 245 289 246 
<< m1 >>
rect 289 245 290 246 
<< m1 >>
rect 290 245 291 246 
<< m1 >>
rect 291 245 292 246 
<< m1 >>
rect 292 245 293 246 
<< m1 >>
rect 307 245 308 246 
<< m2 >>
rect 308 245 309 246 
<< m1 >>
rect 334 245 335 246 
<< m1 >>
rect 337 245 338 246 
<< m1 >>
rect 346 245 347 246 
<< m1 >>
rect 352 245 353 246 
<< m1 >>
rect 379 245 380 246 
<< m2 >>
rect 380 245 381 246 
<< m1 >>
rect 416 245 417 246 
<< m1 >>
rect 419 245 420 246 
<< m1 >>
rect 421 245 422 246 
<< m2 >>
rect 422 245 423 246 
<< m1 >>
rect 434 245 435 246 
<< m1 >>
rect 442 245 443 246 
<< m2 >>
rect 442 245 443 246 
<< m1 >>
rect 481 245 482 246 
<< m1 >>
rect 496 245 497 246 
<< m1 >>
rect 499 245 500 246 
<< m1 >>
rect 523 245 524 246 
<< pdiffusion >>
rect 12 246 13 247 
<< pdiffusion >>
rect 13 246 14 247 
<< pdiffusion >>
rect 14 246 15 247 
<< pdiffusion >>
rect 15 246 16 247 
<< pdiffusion >>
rect 16 246 17 247 
<< pdiffusion >>
rect 17 246 18 247 
<< m1 >>
rect 19 246 20 247 
<< m1 >>
rect 22 246 23 247 
<< pdiffusion >>
rect 30 246 31 247 
<< pdiffusion >>
rect 31 246 32 247 
<< pdiffusion >>
rect 32 246 33 247 
<< pdiffusion >>
rect 33 246 34 247 
<< pdiffusion >>
rect 34 246 35 247 
<< pdiffusion >>
rect 35 246 36 247 
<< m1 >>
rect 44 246 45 247 
<< pdiffusion >>
rect 48 246 49 247 
<< pdiffusion >>
rect 49 246 50 247 
<< pdiffusion >>
rect 50 246 51 247 
<< pdiffusion >>
rect 51 246 52 247 
<< m1 >>
rect 52 246 53 247 
<< pdiffusion >>
rect 52 246 53 247 
<< pdiffusion >>
rect 53 246 54 247 
<< m1 >>
rect 55 246 56 247 
<< m2 >>
rect 56 246 57 247 
<< m1 >>
rect 64 246 65 247 
<< pdiffusion >>
rect 66 246 67 247 
<< pdiffusion >>
rect 67 246 68 247 
<< pdiffusion >>
rect 68 246 69 247 
<< pdiffusion >>
rect 69 246 70 247 
<< pdiffusion >>
rect 70 246 71 247 
<< pdiffusion >>
rect 71 246 72 247 
<< pdiffusion >>
rect 84 246 85 247 
<< pdiffusion >>
rect 85 246 86 247 
<< pdiffusion >>
rect 86 246 87 247 
<< pdiffusion >>
rect 87 246 88 247 
<< pdiffusion >>
rect 88 246 89 247 
<< pdiffusion >>
rect 89 246 90 247 
<< pdiffusion >>
rect 102 246 103 247 
<< pdiffusion >>
rect 103 246 104 247 
<< pdiffusion >>
rect 104 246 105 247 
<< pdiffusion >>
rect 105 246 106 247 
<< m1 >>
rect 106 246 107 247 
<< pdiffusion >>
rect 106 246 107 247 
<< pdiffusion >>
rect 107 246 108 247 
<< m1 >>
rect 118 246 119 247 
<< pdiffusion >>
rect 120 246 121 247 
<< pdiffusion >>
rect 121 246 122 247 
<< pdiffusion >>
rect 122 246 123 247 
<< pdiffusion >>
rect 123 246 124 247 
<< pdiffusion >>
rect 124 246 125 247 
<< pdiffusion >>
rect 125 246 126 247 
<< m1 >>
rect 127 246 128 247 
<< pdiffusion >>
rect 138 246 139 247 
<< pdiffusion >>
rect 139 246 140 247 
<< pdiffusion >>
rect 140 246 141 247 
<< pdiffusion >>
rect 141 246 142 247 
<< pdiffusion >>
rect 142 246 143 247 
<< pdiffusion >>
rect 143 246 144 247 
<< m1 >>
rect 148 246 149 247 
<< pdiffusion >>
rect 156 246 157 247 
<< pdiffusion >>
rect 157 246 158 247 
<< pdiffusion >>
rect 158 246 159 247 
<< pdiffusion >>
rect 159 246 160 247 
<< pdiffusion >>
rect 160 246 161 247 
<< pdiffusion >>
rect 161 246 162 247 
<< m1 >>
rect 163 246 164 247 
<< m2 >>
rect 171 246 172 247 
<< m1 >>
rect 172 246 173 247 
<< pdiffusion >>
rect 174 246 175 247 
<< pdiffusion >>
rect 175 246 176 247 
<< pdiffusion >>
rect 176 246 177 247 
<< pdiffusion >>
rect 177 246 178 247 
<< pdiffusion >>
rect 178 246 179 247 
<< pdiffusion >>
rect 179 246 180 247 
<< m1 >>
rect 181 246 182 247 
<< m2 >>
rect 182 246 183 247 
<< m1 >>
rect 186 246 187 247 
<< m1 >>
rect 190 246 191 247 
<< pdiffusion >>
rect 192 246 193 247 
<< m1 >>
rect 193 246 194 247 
<< pdiffusion >>
rect 193 246 194 247 
<< pdiffusion >>
rect 194 246 195 247 
<< pdiffusion >>
rect 195 246 196 247 
<< pdiffusion >>
rect 196 246 197 247 
<< pdiffusion >>
rect 197 246 198 247 
<< m1 >>
rect 207 246 208 247 
<< pdiffusion >>
rect 210 246 211 247 
<< m1 >>
rect 211 246 212 247 
<< pdiffusion >>
rect 211 246 212 247 
<< pdiffusion >>
rect 212 246 213 247 
<< pdiffusion >>
rect 213 246 214 247 
<< pdiffusion >>
rect 214 246 215 247 
<< pdiffusion >>
rect 215 246 216 247 
<< m1 >>
rect 224 246 225 247 
<< m1 >>
rect 226 246 227 247 
<< pdiffusion >>
rect 228 246 229 247 
<< pdiffusion >>
rect 229 246 230 247 
<< pdiffusion >>
rect 230 246 231 247 
<< pdiffusion >>
rect 231 246 232 247 
<< pdiffusion >>
rect 232 246 233 247 
<< pdiffusion >>
rect 233 246 234 247 
<< m1 >>
rect 235 246 236 247 
<< m1 >>
rect 237 246 238 247 
<< pdiffusion >>
rect 246 246 247 247 
<< pdiffusion >>
rect 247 246 248 247 
<< pdiffusion >>
rect 248 246 249 247 
<< pdiffusion >>
rect 249 246 250 247 
<< m1 >>
rect 250 246 251 247 
<< pdiffusion >>
rect 250 246 251 247 
<< pdiffusion >>
rect 251 246 252 247 
<< m1 >>
rect 253 246 254 247 
<< m2 >>
rect 253 246 254 247 
<< m2c >>
rect 253 246 254 247 
<< m1 >>
rect 253 246 254 247 
<< m2 >>
rect 253 246 254 247 
<< m1 >>
rect 254 246 255 247 
<< m1 >>
rect 255 246 256 247 
<< m1 >>
rect 262 246 263 247 
<< m2 >>
rect 262 246 263 247 
<< pdiffusion >>
rect 264 246 265 247 
<< pdiffusion >>
rect 265 246 266 247 
<< pdiffusion >>
rect 266 246 267 247 
<< pdiffusion >>
rect 267 246 268 247 
<< pdiffusion >>
rect 268 246 269 247 
<< pdiffusion >>
rect 269 246 270 247 
<< m1 >>
rect 274 246 275 247 
<< m1 >>
rect 276 246 277 247 
<< pdiffusion >>
rect 300 246 301 247 
<< pdiffusion >>
rect 301 246 302 247 
<< pdiffusion >>
rect 302 246 303 247 
<< pdiffusion >>
rect 303 246 304 247 
<< pdiffusion >>
rect 304 246 305 247 
<< pdiffusion >>
rect 305 246 306 247 
<< m1 >>
rect 307 246 308 247 
<< m2 >>
rect 308 246 309 247 
<< pdiffusion >>
rect 318 246 319 247 
<< pdiffusion >>
rect 319 246 320 247 
<< pdiffusion >>
rect 320 246 321 247 
<< pdiffusion >>
rect 321 246 322 247 
<< pdiffusion >>
rect 322 246 323 247 
<< pdiffusion >>
rect 323 246 324 247 
<< m1 >>
rect 334 246 335 247 
<< pdiffusion >>
rect 336 246 337 247 
<< m1 >>
rect 337 246 338 247 
<< pdiffusion >>
rect 337 246 338 247 
<< pdiffusion >>
rect 338 246 339 247 
<< pdiffusion >>
rect 339 246 340 247 
<< pdiffusion >>
rect 340 246 341 247 
<< pdiffusion >>
rect 341 246 342 247 
<< m1 >>
rect 346 246 347 247 
<< m1 >>
rect 352 246 353 247 
<< pdiffusion >>
rect 372 246 373 247 
<< pdiffusion >>
rect 373 246 374 247 
<< pdiffusion >>
rect 374 246 375 247 
<< pdiffusion >>
rect 375 246 376 247 
<< pdiffusion >>
rect 376 246 377 247 
<< pdiffusion >>
rect 377 246 378 247 
<< m1 >>
rect 379 246 380 247 
<< m2 >>
rect 380 246 381 247 
<< pdiffusion >>
rect 390 246 391 247 
<< pdiffusion >>
rect 391 246 392 247 
<< pdiffusion >>
rect 392 246 393 247 
<< pdiffusion >>
rect 393 246 394 247 
<< pdiffusion >>
rect 394 246 395 247 
<< pdiffusion >>
rect 395 246 396 247 
<< pdiffusion >>
rect 408 246 409 247 
<< pdiffusion >>
rect 409 246 410 247 
<< pdiffusion >>
rect 410 246 411 247 
<< pdiffusion >>
rect 411 246 412 247 
<< pdiffusion >>
rect 412 246 413 247 
<< pdiffusion >>
rect 413 246 414 247 
<< m1 >>
rect 416 246 417 247 
<< m1 >>
rect 419 246 420 247 
<< m1 >>
rect 421 246 422 247 
<< m2 >>
rect 422 246 423 247 
<< pdiffusion >>
rect 426 246 427 247 
<< pdiffusion >>
rect 427 246 428 247 
<< pdiffusion >>
rect 428 246 429 247 
<< pdiffusion >>
rect 429 246 430 247 
<< pdiffusion >>
rect 430 246 431 247 
<< pdiffusion >>
rect 431 246 432 247 
<< m1 >>
rect 434 246 435 247 
<< m1 >>
rect 442 246 443 247 
<< m2 >>
rect 442 246 443 247 
<< pdiffusion >>
rect 444 246 445 247 
<< pdiffusion >>
rect 445 246 446 247 
<< pdiffusion >>
rect 446 246 447 247 
<< pdiffusion >>
rect 447 246 448 247 
<< pdiffusion >>
rect 448 246 449 247 
<< pdiffusion >>
rect 449 246 450 247 
<< pdiffusion >>
rect 462 246 463 247 
<< pdiffusion >>
rect 463 246 464 247 
<< pdiffusion >>
rect 464 246 465 247 
<< pdiffusion >>
rect 465 246 466 247 
<< pdiffusion >>
rect 466 246 467 247 
<< pdiffusion >>
rect 467 246 468 247 
<< pdiffusion >>
rect 480 246 481 247 
<< m1 >>
rect 481 246 482 247 
<< pdiffusion >>
rect 481 246 482 247 
<< pdiffusion >>
rect 482 246 483 247 
<< pdiffusion >>
rect 483 246 484 247 
<< pdiffusion >>
rect 484 246 485 247 
<< pdiffusion >>
rect 485 246 486 247 
<< m1 >>
rect 496 246 497 247 
<< pdiffusion >>
rect 498 246 499 247 
<< m1 >>
rect 499 246 500 247 
<< pdiffusion >>
rect 499 246 500 247 
<< pdiffusion >>
rect 500 246 501 247 
<< pdiffusion >>
rect 501 246 502 247 
<< pdiffusion >>
rect 502 246 503 247 
<< pdiffusion >>
rect 503 246 504 247 
<< pdiffusion >>
rect 516 246 517 247 
<< pdiffusion >>
rect 517 246 518 247 
<< pdiffusion >>
rect 518 246 519 247 
<< pdiffusion >>
rect 519 246 520 247 
<< pdiffusion >>
rect 520 246 521 247 
<< pdiffusion >>
rect 521 246 522 247 
<< m1 >>
rect 523 246 524 247 
<< pdiffusion >>
rect 12 247 13 248 
<< pdiffusion >>
rect 13 247 14 248 
<< pdiffusion >>
rect 14 247 15 248 
<< pdiffusion >>
rect 15 247 16 248 
<< pdiffusion >>
rect 16 247 17 248 
<< pdiffusion >>
rect 17 247 18 248 
<< m1 >>
rect 19 247 20 248 
<< m1 >>
rect 22 247 23 248 
<< pdiffusion >>
rect 30 247 31 248 
<< pdiffusion >>
rect 31 247 32 248 
<< pdiffusion >>
rect 32 247 33 248 
<< pdiffusion >>
rect 33 247 34 248 
<< pdiffusion >>
rect 34 247 35 248 
<< pdiffusion >>
rect 35 247 36 248 
<< m1 >>
rect 44 247 45 248 
<< pdiffusion >>
rect 48 247 49 248 
<< pdiffusion >>
rect 49 247 50 248 
<< pdiffusion >>
rect 50 247 51 248 
<< pdiffusion >>
rect 51 247 52 248 
<< pdiffusion >>
rect 52 247 53 248 
<< pdiffusion >>
rect 53 247 54 248 
<< m1 >>
rect 55 247 56 248 
<< m2 >>
rect 56 247 57 248 
<< m1 >>
rect 64 247 65 248 
<< pdiffusion >>
rect 66 247 67 248 
<< pdiffusion >>
rect 67 247 68 248 
<< pdiffusion >>
rect 68 247 69 248 
<< pdiffusion >>
rect 69 247 70 248 
<< pdiffusion >>
rect 70 247 71 248 
<< pdiffusion >>
rect 71 247 72 248 
<< pdiffusion >>
rect 84 247 85 248 
<< pdiffusion >>
rect 85 247 86 248 
<< pdiffusion >>
rect 86 247 87 248 
<< pdiffusion >>
rect 87 247 88 248 
<< pdiffusion >>
rect 88 247 89 248 
<< pdiffusion >>
rect 89 247 90 248 
<< pdiffusion >>
rect 102 247 103 248 
<< pdiffusion >>
rect 103 247 104 248 
<< pdiffusion >>
rect 104 247 105 248 
<< pdiffusion >>
rect 105 247 106 248 
<< pdiffusion >>
rect 106 247 107 248 
<< pdiffusion >>
rect 107 247 108 248 
<< m1 >>
rect 118 247 119 248 
<< pdiffusion >>
rect 120 247 121 248 
<< pdiffusion >>
rect 121 247 122 248 
<< pdiffusion >>
rect 122 247 123 248 
<< pdiffusion >>
rect 123 247 124 248 
<< pdiffusion >>
rect 124 247 125 248 
<< pdiffusion >>
rect 125 247 126 248 
<< m1 >>
rect 127 247 128 248 
<< pdiffusion >>
rect 138 247 139 248 
<< pdiffusion >>
rect 139 247 140 248 
<< pdiffusion >>
rect 140 247 141 248 
<< pdiffusion >>
rect 141 247 142 248 
<< pdiffusion >>
rect 142 247 143 248 
<< pdiffusion >>
rect 143 247 144 248 
<< m1 >>
rect 148 247 149 248 
<< pdiffusion >>
rect 156 247 157 248 
<< pdiffusion >>
rect 157 247 158 248 
<< pdiffusion >>
rect 158 247 159 248 
<< pdiffusion >>
rect 159 247 160 248 
<< pdiffusion >>
rect 160 247 161 248 
<< pdiffusion >>
rect 161 247 162 248 
<< m1 >>
rect 163 247 164 248 
<< m2 >>
rect 171 247 172 248 
<< m1 >>
rect 172 247 173 248 
<< pdiffusion >>
rect 174 247 175 248 
<< pdiffusion >>
rect 175 247 176 248 
<< pdiffusion >>
rect 176 247 177 248 
<< pdiffusion >>
rect 177 247 178 248 
<< pdiffusion >>
rect 178 247 179 248 
<< pdiffusion >>
rect 179 247 180 248 
<< m1 >>
rect 181 247 182 248 
<< m2 >>
rect 182 247 183 248 
<< m1 >>
rect 186 247 187 248 
<< m1 >>
rect 190 247 191 248 
<< pdiffusion >>
rect 192 247 193 248 
<< pdiffusion >>
rect 193 247 194 248 
<< pdiffusion >>
rect 194 247 195 248 
<< pdiffusion >>
rect 195 247 196 248 
<< pdiffusion >>
rect 196 247 197 248 
<< pdiffusion >>
rect 197 247 198 248 
<< m1 >>
rect 207 247 208 248 
<< pdiffusion >>
rect 210 247 211 248 
<< pdiffusion >>
rect 211 247 212 248 
<< pdiffusion >>
rect 212 247 213 248 
<< pdiffusion >>
rect 213 247 214 248 
<< pdiffusion >>
rect 214 247 215 248 
<< pdiffusion >>
rect 215 247 216 248 
<< m1 >>
rect 224 247 225 248 
<< m1 >>
rect 226 247 227 248 
<< pdiffusion >>
rect 228 247 229 248 
<< pdiffusion >>
rect 229 247 230 248 
<< pdiffusion >>
rect 230 247 231 248 
<< pdiffusion >>
rect 231 247 232 248 
<< pdiffusion >>
rect 232 247 233 248 
<< pdiffusion >>
rect 233 247 234 248 
<< m1 >>
rect 235 247 236 248 
<< m1 >>
rect 237 247 238 248 
<< pdiffusion >>
rect 246 247 247 248 
<< pdiffusion >>
rect 247 247 248 248 
<< pdiffusion >>
rect 248 247 249 248 
<< pdiffusion >>
rect 249 247 250 248 
<< pdiffusion >>
rect 250 247 251 248 
<< pdiffusion >>
rect 251 247 252 248 
<< m1 >>
rect 255 247 256 248 
<< m1 >>
rect 262 247 263 248 
<< m2 >>
rect 262 247 263 248 
<< pdiffusion >>
rect 264 247 265 248 
<< pdiffusion >>
rect 265 247 266 248 
<< pdiffusion >>
rect 266 247 267 248 
<< pdiffusion >>
rect 267 247 268 248 
<< pdiffusion >>
rect 268 247 269 248 
<< pdiffusion >>
rect 269 247 270 248 
<< m1 >>
rect 274 247 275 248 
<< m1 >>
rect 276 247 277 248 
<< pdiffusion >>
rect 300 247 301 248 
<< pdiffusion >>
rect 301 247 302 248 
<< pdiffusion >>
rect 302 247 303 248 
<< pdiffusion >>
rect 303 247 304 248 
<< pdiffusion >>
rect 304 247 305 248 
<< pdiffusion >>
rect 305 247 306 248 
<< m1 >>
rect 307 247 308 248 
<< m2 >>
rect 308 247 309 248 
<< pdiffusion >>
rect 318 247 319 248 
<< pdiffusion >>
rect 319 247 320 248 
<< pdiffusion >>
rect 320 247 321 248 
<< pdiffusion >>
rect 321 247 322 248 
<< pdiffusion >>
rect 322 247 323 248 
<< pdiffusion >>
rect 323 247 324 248 
<< m1 >>
rect 334 247 335 248 
<< pdiffusion >>
rect 336 247 337 248 
<< pdiffusion >>
rect 337 247 338 248 
<< pdiffusion >>
rect 338 247 339 248 
<< pdiffusion >>
rect 339 247 340 248 
<< pdiffusion >>
rect 340 247 341 248 
<< pdiffusion >>
rect 341 247 342 248 
<< m1 >>
rect 346 247 347 248 
<< m1 >>
rect 352 247 353 248 
<< pdiffusion >>
rect 372 247 373 248 
<< pdiffusion >>
rect 373 247 374 248 
<< pdiffusion >>
rect 374 247 375 248 
<< pdiffusion >>
rect 375 247 376 248 
<< pdiffusion >>
rect 376 247 377 248 
<< pdiffusion >>
rect 377 247 378 248 
<< m1 >>
rect 379 247 380 248 
<< m2 >>
rect 380 247 381 248 
<< pdiffusion >>
rect 390 247 391 248 
<< pdiffusion >>
rect 391 247 392 248 
<< pdiffusion >>
rect 392 247 393 248 
<< pdiffusion >>
rect 393 247 394 248 
<< pdiffusion >>
rect 394 247 395 248 
<< pdiffusion >>
rect 395 247 396 248 
<< pdiffusion >>
rect 408 247 409 248 
<< pdiffusion >>
rect 409 247 410 248 
<< pdiffusion >>
rect 410 247 411 248 
<< pdiffusion >>
rect 411 247 412 248 
<< pdiffusion >>
rect 412 247 413 248 
<< pdiffusion >>
rect 413 247 414 248 
<< m1 >>
rect 416 247 417 248 
<< m1 >>
rect 419 247 420 248 
<< m1 >>
rect 421 247 422 248 
<< m2 >>
rect 422 247 423 248 
<< pdiffusion >>
rect 426 247 427 248 
<< pdiffusion >>
rect 427 247 428 248 
<< pdiffusion >>
rect 428 247 429 248 
<< pdiffusion >>
rect 429 247 430 248 
<< pdiffusion >>
rect 430 247 431 248 
<< pdiffusion >>
rect 431 247 432 248 
<< m1 >>
rect 434 247 435 248 
<< m1 >>
rect 442 247 443 248 
<< m2 >>
rect 442 247 443 248 
<< pdiffusion >>
rect 444 247 445 248 
<< pdiffusion >>
rect 445 247 446 248 
<< pdiffusion >>
rect 446 247 447 248 
<< pdiffusion >>
rect 447 247 448 248 
<< pdiffusion >>
rect 448 247 449 248 
<< pdiffusion >>
rect 449 247 450 248 
<< pdiffusion >>
rect 462 247 463 248 
<< pdiffusion >>
rect 463 247 464 248 
<< pdiffusion >>
rect 464 247 465 248 
<< pdiffusion >>
rect 465 247 466 248 
<< pdiffusion >>
rect 466 247 467 248 
<< pdiffusion >>
rect 467 247 468 248 
<< pdiffusion >>
rect 480 247 481 248 
<< pdiffusion >>
rect 481 247 482 248 
<< pdiffusion >>
rect 482 247 483 248 
<< pdiffusion >>
rect 483 247 484 248 
<< pdiffusion >>
rect 484 247 485 248 
<< pdiffusion >>
rect 485 247 486 248 
<< m1 >>
rect 496 247 497 248 
<< pdiffusion >>
rect 498 247 499 248 
<< pdiffusion >>
rect 499 247 500 248 
<< pdiffusion >>
rect 500 247 501 248 
<< pdiffusion >>
rect 501 247 502 248 
<< pdiffusion >>
rect 502 247 503 248 
<< pdiffusion >>
rect 503 247 504 248 
<< pdiffusion >>
rect 516 247 517 248 
<< pdiffusion >>
rect 517 247 518 248 
<< pdiffusion >>
rect 518 247 519 248 
<< pdiffusion >>
rect 519 247 520 248 
<< pdiffusion >>
rect 520 247 521 248 
<< pdiffusion >>
rect 521 247 522 248 
<< m1 >>
rect 523 247 524 248 
<< pdiffusion >>
rect 12 248 13 249 
<< pdiffusion >>
rect 13 248 14 249 
<< pdiffusion >>
rect 14 248 15 249 
<< pdiffusion >>
rect 15 248 16 249 
<< pdiffusion >>
rect 16 248 17 249 
<< pdiffusion >>
rect 17 248 18 249 
<< m1 >>
rect 19 248 20 249 
<< m1 >>
rect 22 248 23 249 
<< pdiffusion >>
rect 30 248 31 249 
<< pdiffusion >>
rect 31 248 32 249 
<< pdiffusion >>
rect 32 248 33 249 
<< pdiffusion >>
rect 33 248 34 249 
<< pdiffusion >>
rect 34 248 35 249 
<< pdiffusion >>
rect 35 248 36 249 
<< m1 >>
rect 44 248 45 249 
<< pdiffusion >>
rect 48 248 49 249 
<< pdiffusion >>
rect 49 248 50 249 
<< pdiffusion >>
rect 50 248 51 249 
<< pdiffusion >>
rect 51 248 52 249 
<< pdiffusion >>
rect 52 248 53 249 
<< pdiffusion >>
rect 53 248 54 249 
<< m1 >>
rect 55 248 56 249 
<< m2 >>
rect 56 248 57 249 
<< m1 >>
rect 64 248 65 249 
<< pdiffusion >>
rect 66 248 67 249 
<< pdiffusion >>
rect 67 248 68 249 
<< pdiffusion >>
rect 68 248 69 249 
<< pdiffusion >>
rect 69 248 70 249 
<< pdiffusion >>
rect 70 248 71 249 
<< pdiffusion >>
rect 71 248 72 249 
<< pdiffusion >>
rect 84 248 85 249 
<< pdiffusion >>
rect 85 248 86 249 
<< pdiffusion >>
rect 86 248 87 249 
<< pdiffusion >>
rect 87 248 88 249 
<< pdiffusion >>
rect 88 248 89 249 
<< pdiffusion >>
rect 89 248 90 249 
<< pdiffusion >>
rect 102 248 103 249 
<< pdiffusion >>
rect 103 248 104 249 
<< pdiffusion >>
rect 104 248 105 249 
<< pdiffusion >>
rect 105 248 106 249 
<< pdiffusion >>
rect 106 248 107 249 
<< pdiffusion >>
rect 107 248 108 249 
<< m1 >>
rect 118 248 119 249 
<< pdiffusion >>
rect 120 248 121 249 
<< pdiffusion >>
rect 121 248 122 249 
<< pdiffusion >>
rect 122 248 123 249 
<< pdiffusion >>
rect 123 248 124 249 
<< pdiffusion >>
rect 124 248 125 249 
<< pdiffusion >>
rect 125 248 126 249 
<< m1 >>
rect 127 248 128 249 
<< pdiffusion >>
rect 138 248 139 249 
<< pdiffusion >>
rect 139 248 140 249 
<< pdiffusion >>
rect 140 248 141 249 
<< pdiffusion >>
rect 141 248 142 249 
<< pdiffusion >>
rect 142 248 143 249 
<< pdiffusion >>
rect 143 248 144 249 
<< m1 >>
rect 148 248 149 249 
<< pdiffusion >>
rect 156 248 157 249 
<< pdiffusion >>
rect 157 248 158 249 
<< pdiffusion >>
rect 158 248 159 249 
<< pdiffusion >>
rect 159 248 160 249 
<< pdiffusion >>
rect 160 248 161 249 
<< pdiffusion >>
rect 161 248 162 249 
<< m1 >>
rect 163 248 164 249 
<< m2 >>
rect 171 248 172 249 
<< m1 >>
rect 172 248 173 249 
<< pdiffusion >>
rect 174 248 175 249 
<< pdiffusion >>
rect 175 248 176 249 
<< pdiffusion >>
rect 176 248 177 249 
<< pdiffusion >>
rect 177 248 178 249 
<< pdiffusion >>
rect 178 248 179 249 
<< pdiffusion >>
rect 179 248 180 249 
<< m1 >>
rect 181 248 182 249 
<< m2 >>
rect 182 248 183 249 
<< m1 >>
rect 186 248 187 249 
<< m1 >>
rect 190 248 191 249 
<< pdiffusion >>
rect 192 248 193 249 
<< pdiffusion >>
rect 193 248 194 249 
<< pdiffusion >>
rect 194 248 195 249 
<< pdiffusion >>
rect 195 248 196 249 
<< pdiffusion >>
rect 196 248 197 249 
<< pdiffusion >>
rect 197 248 198 249 
<< m1 >>
rect 207 248 208 249 
<< pdiffusion >>
rect 210 248 211 249 
<< pdiffusion >>
rect 211 248 212 249 
<< pdiffusion >>
rect 212 248 213 249 
<< pdiffusion >>
rect 213 248 214 249 
<< pdiffusion >>
rect 214 248 215 249 
<< pdiffusion >>
rect 215 248 216 249 
<< m1 >>
rect 224 248 225 249 
<< m1 >>
rect 226 248 227 249 
<< pdiffusion >>
rect 228 248 229 249 
<< pdiffusion >>
rect 229 248 230 249 
<< pdiffusion >>
rect 230 248 231 249 
<< pdiffusion >>
rect 231 248 232 249 
<< pdiffusion >>
rect 232 248 233 249 
<< pdiffusion >>
rect 233 248 234 249 
<< m1 >>
rect 235 248 236 249 
<< m1 >>
rect 237 248 238 249 
<< pdiffusion >>
rect 246 248 247 249 
<< pdiffusion >>
rect 247 248 248 249 
<< pdiffusion >>
rect 248 248 249 249 
<< pdiffusion >>
rect 249 248 250 249 
<< pdiffusion >>
rect 250 248 251 249 
<< pdiffusion >>
rect 251 248 252 249 
<< m1 >>
rect 255 248 256 249 
<< m1 >>
rect 262 248 263 249 
<< m2 >>
rect 262 248 263 249 
<< pdiffusion >>
rect 264 248 265 249 
<< pdiffusion >>
rect 265 248 266 249 
<< pdiffusion >>
rect 266 248 267 249 
<< pdiffusion >>
rect 267 248 268 249 
<< pdiffusion >>
rect 268 248 269 249 
<< pdiffusion >>
rect 269 248 270 249 
<< m1 >>
rect 274 248 275 249 
<< m1 >>
rect 276 248 277 249 
<< pdiffusion >>
rect 300 248 301 249 
<< pdiffusion >>
rect 301 248 302 249 
<< pdiffusion >>
rect 302 248 303 249 
<< pdiffusion >>
rect 303 248 304 249 
<< pdiffusion >>
rect 304 248 305 249 
<< pdiffusion >>
rect 305 248 306 249 
<< m1 >>
rect 307 248 308 249 
<< m2 >>
rect 308 248 309 249 
<< pdiffusion >>
rect 318 248 319 249 
<< pdiffusion >>
rect 319 248 320 249 
<< pdiffusion >>
rect 320 248 321 249 
<< pdiffusion >>
rect 321 248 322 249 
<< pdiffusion >>
rect 322 248 323 249 
<< pdiffusion >>
rect 323 248 324 249 
<< m1 >>
rect 334 248 335 249 
<< pdiffusion >>
rect 336 248 337 249 
<< pdiffusion >>
rect 337 248 338 249 
<< pdiffusion >>
rect 338 248 339 249 
<< pdiffusion >>
rect 339 248 340 249 
<< pdiffusion >>
rect 340 248 341 249 
<< pdiffusion >>
rect 341 248 342 249 
<< m1 >>
rect 346 248 347 249 
<< m1 >>
rect 352 248 353 249 
<< pdiffusion >>
rect 372 248 373 249 
<< pdiffusion >>
rect 373 248 374 249 
<< pdiffusion >>
rect 374 248 375 249 
<< pdiffusion >>
rect 375 248 376 249 
<< pdiffusion >>
rect 376 248 377 249 
<< pdiffusion >>
rect 377 248 378 249 
<< m1 >>
rect 379 248 380 249 
<< m2 >>
rect 380 248 381 249 
<< pdiffusion >>
rect 390 248 391 249 
<< pdiffusion >>
rect 391 248 392 249 
<< pdiffusion >>
rect 392 248 393 249 
<< pdiffusion >>
rect 393 248 394 249 
<< pdiffusion >>
rect 394 248 395 249 
<< pdiffusion >>
rect 395 248 396 249 
<< pdiffusion >>
rect 408 248 409 249 
<< pdiffusion >>
rect 409 248 410 249 
<< pdiffusion >>
rect 410 248 411 249 
<< pdiffusion >>
rect 411 248 412 249 
<< pdiffusion >>
rect 412 248 413 249 
<< pdiffusion >>
rect 413 248 414 249 
<< m1 >>
rect 416 248 417 249 
<< m1 >>
rect 419 248 420 249 
<< m1 >>
rect 421 248 422 249 
<< m2 >>
rect 422 248 423 249 
<< pdiffusion >>
rect 426 248 427 249 
<< pdiffusion >>
rect 427 248 428 249 
<< pdiffusion >>
rect 428 248 429 249 
<< pdiffusion >>
rect 429 248 430 249 
<< pdiffusion >>
rect 430 248 431 249 
<< pdiffusion >>
rect 431 248 432 249 
<< m1 >>
rect 434 248 435 249 
<< m1 >>
rect 442 248 443 249 
<< m2 >>
rect 442 248 443 249 
<< pdiffusion >>
rect 444 248 445 249 
<< pdiffusion >>
rect 445 248 446 249 
<< pdiffusion >>
rect 446 248 447 249 
<< pdiffusion >>
rect 447 248 448 249 
<< pdiffusion >>
rect 448 248 449 249 
<< pdiffusion >>
rect 449 248 450 249 
<< pdiffusion >>
rect 462 248 463 249 
<< pdiffusion >>
rect 463 248 464 249 
<< pdiffusion >>
rect 464 248 465 249 
<< pdiffusion >>
rect 465 248 466 249 
<< pdiffusion >>
rect 466 248 467 249 
<< pdiffusion >>
rect 467 248 468 249 
<< pdiffusion >>
rect 480 248 481 249 
<< pdiffusion >>
rect 481 248 482 249 
<< pdiffusion >>
rect 482 248 483 249 
<< pdiffusion >>
rect 483 248 484 249 
<< pdiffusion >>
rect 484 248 485 249 
<< pdiffusion >>
rect 485 248 486 249 
<< m1 >>
rect 496 248 497 249 
<< pdiffusion >>
rect 498 248 499 249 
<< pdiffusion >>
rect 499 248 500 249 
<< pdiffusion >>
rect 500 248 501 249 
<< pdiffusion >>
rect 501 248 502 249 
<< pdiffusion >>
rect 502 248 503 249 
<< pdiffusion >>
rect 503 248 504 249 
<< pdiffusion >>
rect 516 248 517 249 
<< pdiffusion >>
rect 517 248 518 249 
<< pdiffusion >>
rect 518 248 519 249 
<< pdiffusion >>
rect 519 248 520 249 
<< pdiffusion >>
rect 520 248 521 249 
<< pdiffusion >>
rect 521 248 522 249 
<< m1 >>
rect 523 248 524 249 
<< pdiffusion >>
rect 12 249 13 250 
<< pdiffusion >>
rect 13 249 14 250 
<< pdiffusion >>
rect 14 249 15 250 
<< pdiffusion >>
rect 15 249 16 250 
<< pdiffusion >>
rect 16 249 17 250 
<< pdiffusion >>
rect 17 249 18 250 
<< m1 >>
rect 19 249 20 250 
<< m1 >>
rect 22 249 23 250 
<< pdiffusion >>
rect 30 249 31 250 
<< pdiffusion >>
rect 31 249 32 250 
<< pdiffusion >>
rect 32 249 33 250 
<< pdiffusion >>
rect 33 249 34 250 
<< pdiffusion >>
rect 34 249 35 250 
<< pdiffusion >>
rect 35 249 36 250 
<< m1 >>
rect 44 249 45 250 
<< pdiffusion >>
rect 48 249 49 250 
<< pdiffusion >>
rect 49 249 50 250 
<< pdiffusion >>
rect 50 249 51 250 
<< pdiffusion >>
rect 51 249 52 250 
<< pdiffusion >>
rect 52 249 53 250 
<< pdiffusion >>
rect 53 249 54 250 
<< m1 >>
rect 55 249 56 250 
<< m2 >>
rect 56 249 57 250 
<< m1 >>
rect 64 249 65 250 
<< pdiffusion >>
rect 66 249 67 250 
<< pdiffusion >>
rect 67 249 68 250 
<< pdiffusion >>
rect 68 249 69 250 
<< pdiffusion >>
rect 69 249 70 250 
<< pdiffusion >>
rect 70 249 71 250 
<< pdiffusion >>
rect 71 249 72 250 
<< pdiffusion >>
rect 84 249 85 250 
<< pdiffusion >>
rect 85 249 86 250 
<< pdiffusion >>
rect 86 249 87 250 
<< pdiffusion >>
rect 87 249 88 250 
<< pdiffusion >>
rect 88 249 89 250 
<< pdiffusion >>
rect 89 249 90 250 
<< pdiffusion >>
rect 102 249 103 250 
<< pdiffusion >>
rect 103 249 104 250 
<< pdiffusion >>
rect 104 249 105 250 
<< pdiffusion >>
rect 105 249 106 250 
<< pdiffusion >>
rect 106 249 107 250 
<< pdiffusion >>
rect 107 249 108 250 
<< m1 >>
rect 118 249 119 250 
<< pdiffusion >>
rect 120 249 121 250 
<< pdiffusion >>
rect 121 249 122 250 
<< pdiffusion >>
rect 122 249 123 250 
<< pdiffusion >>
rect 123 249 124 250 
<< pdiffusion >>
rect 124 249 125 250 
<< pdiffusion >>
rect 125 249 126 250 
<< m1 >>
rect 127 249 128 250 
<< pdiffusion >>
rect 138 249 139 250 
<< pdiffusion >>
rect 139 249 140 250 
<< pdiffusion >>
rect 140 249 141 250 
<< pdiffusion >>
rect 141 249 142 250 
<< pdiffusion >>
rect 142 249 143 250 
<< pdiffusion >>
rect 143 249 144 250 
<< m1 >>
rect 148 249 149 250 
<< pdiffusion >>
rect 156 249 157 250 
<< pdiffusion >>
rect 157 249 158 250 
<< pdiffusion >>
rect 158 249 159 250 
<< pdiffusion >>
rect 159 249 160 250 
<< pdiffusion >>
rect 160 249 161 250 
<< pdiffusion >>
rect 161 249 162 250 
<< m1 >>
rect 163 249 164 250 
<< m2 >>
rect 171 249 172 250 
<< m1 >>
rect 172 249 173 250 
<< pdiffusion >>
rect 174 249 175 250 
<< pdiffusion >>
rect 175 249 176 250 
<< pdiffusion >>
rect 176 249 177 250 
<< pdiffusion >>
rect 177 249 178 250 
<< pdiffusion >>
rect 178 249 179 250 
<< pdiffusion >>
rect 179 249 180 250 
<< m1 >>
rect 181 249 182 250 
<< m2 >>
rect 182 249 183 250 
<< m1 >>
rect 186 249 187 250 
<< m1 >>
rect 190 249 191 250 
<< pdiffusion >>
rect 192 249 193 250 
<< pdiffusion >>
rect 193 249 194 250 
<< pdiffusion >>
rect 194 249 195 250 
<< pdiffusion >>
rect 195 249 196 250 
<< pdiffusion >>
rect 196 249 197 250 
<< pdiffusion >>
rect 197 249 198 250 
<< m1 >>
rect 207 249 208 250 
<< pdiffusion >>
rect 210 249 211 250 
<< pdiffusion >>
rect 211 249 212 250 
<< pdiffusion >>
rect 212 249 213 250 
<< pdiffusion >>
rect 213 249 214 250 
<< pdiffusion >>
rect 214 249 215 250 
<< pdiffusion >>
rect 215 249 216 250 
<< m1 >>
rect 224 249 225 250 
<< m1 >>
rect 226 249 227 250 
<< pdiffusion >>
rect 228 249 229 250 
<< pdiffusion >>
rect 229 249 230 250 
<< pdiffusion >>
rect 230 249 231 250 
<< pdiffusion >>
rect 231 249 232 250 
<< pdiffusion >>
rect 232 249 233 250 
<< pdiffusion >>
rect 233 249 234 250 
<< m1 >>
rect 235 249 236 250 
<< m1 >>
rect 237 249 238 250 
<< pdiffusion >>
rect 246 249 247 250 
<< pdiffusion >>
rect 247 249 248 250 
<< pdiffusion >>
rect 248 249 249 250 
<< pdiffusion >>
rect 249 249 250 250 
<< pdiffusion >>
rect 250 249 251 250 
<< pdiffusion >>
rect 251 249 252 250 
<< m1 >>
rect 255 249 256 250 
<< m1 >>
rect 262 249 263 250 
<< m2 >>
rect 262 249 263 250 
<< pdiffusion >>
rect 264 249 265 250 
<< pdiffusion >>
rect 265 249 266 250 
<< pdiffusion >>
rect 266 249 267 250 
<< pdiffusion >>
rect 267 249 268 250 
<< pdiffusion >>
rect 268 249 269 250 
<< pdiffusion >>
rect 269 249 270 250 
<< m1 >>
rect 274 249 275 250 
<< m1 >>
rect 276 249 277 250 
<< pdiffusion >>
rect 300 249 301 250 
<< pdiffusion >>
rect 301 249 302 250 
<< pdiffusion >>
rect 302 249 303 250 
<< pdiffusion >>
rect 303 249 304 250 
<< pdiffusion >>
rect 304 249 305 250 
<< pdiffusion >>
rect 305 249 306 250 
<< m1 >>
rect 307 249 308 250 
<< m2 >>
rect 308 249 309 250 
<< pdiffusion >>
rect 318 249 319 250 
<< pdiffusion >>
rect 319 249 320 250 
<< pdiffusion >>
rect 320 249 321 250 
<< pdiffusion >>
rect 321 249 322 250 
<< pdiffusion >>
rect 322 249 323 250 
<< pdiffusion >>
rect 323 249 324 250 
<< m1 >>
rect 334 249 335 250 
<< pdiffusion >>
rect 336 249 337 250 
<< pdiffusion >>
rect 337 249 338 250 
<< pdiffusion >>
rect 338 249 339 250 
<< pdiffusion >>
rect 339 249 340 250 
<< pdiffusion >>
rect 340 249 341 250 
<< pdiffusion >>
rect 341 249 342 250 
<< m1 >>
rect 346 249 347 250 
<< m1 >>
rect 352 249 353 250 
<< pdiffusion >>
rect 372 249 373 250 
<< pdiffusion >>
rect 373 249 374 250 
<< pdiffusion >>
rect 374 249 375 250 
<< pdiffusion >>
rect 375 249 376 250 
<< pdiffusion >>
rect 376 249 377 250 
<< pdiffusion >>
rect 377 249 378 250 
<< m1 >>
rect 379 249 380 250 
<< m2 >>
rect 380 249 381 250 
<< pdiffusion >>
rect 390 249 391 250 
<< pdiffusion >>
rect 391 249 392 250 
<< pdiffusion >>
rect 392 249 393 250 
<< pdiffusion >>
rect 393 249 394 250 
<< pdiffusion >>
rect 394 249 395 250 
<< pdiffusion >>
rect 395 249 396 250 
<< pdiffusion >>
rect 408 249 409 250 
<< pdiffusion >>
rect 409 249 410 250 
<< pdiffusion >>
rect 410 249 411 250 
<< pdiffusion >>
rect 411 249 412 250 
<< pdiffusion >>
rect 412 249 413 250 
<< pdiffusion >>
rect 413 249 414 250 
<< m1 >>
rect 416 249 417 250 
<< m1 >>
rect 419 249 420 250 
<< m1 >>
rect 421 249 422 250 
<< m2 >>
rect 422 249 423 250 
<< pdiffusion >>
rect 426 249 427 250 
<< pdiffusion >>
rect 427 249 428 250 
<< pdiffusion >>
rect 428 249 429 250 
<< pdiffusion >>
rect 429 249 430 250 
<< pdiffusion >>
rect 430 249 431 250 
<< pdiffusion >>
rect 431 249 432 250 
<< m1 >>
rect 434 249 435 250 
<< m1 >>
rect 442 249 443 250 
<< m2 >>
rect 442 249 443 250 
<< pdiffusion >>
rect 444 249 445 250 
<< pdiffusion >>
rect 445 249 446 250 
<< pdiffusion >>
rect 446 249 447 250 
<< pdiffusion >>
rect 447 249 448 250 
<< pdiffusion >>
rect 448 249 449 250 
<< pdiffusion >>
rect 449 249 450 250 
<< pdiffusion >>
rect 462 249 463 250 
<< pdiffusion >>
rect 463 249 464 250 
<< pdiffusion >>
rect 464 249 465 250 
<< pdiffusion >>
rect 465 249 466 250 
<< pdiffusion >>
rect 466 249 467 250 
<< pdiffusion >>
rect 467 249 468 250 
<< pdiffusion >>
rect 480 249 481 250 
<< pdiffusion >>
rect 481 249 482 250 
<< pdiffusion >>
rect 482 249 483 250 
<< pdiffusion >>
rect 483 249 484 250 
<< pdiffusion >>
rect 484 249 485 250 
<< pdiffusion >>
rect 485 249 486 250 
<< m1 >>
rect 496 249 497 250 
<< pdiffusion >>
rect 498 249 499 250 
<< pdiffusion >>
rect 499 249 500 250 
<< pdiffusion >>
rect 500 249 501 250 
<< pdiffusion >>
rect 501 249 502 250 
<< pdiffusion >>
rect 502 249 503 250 
<< pdiffusion >>
rect 503 249 504 250 
<< pdiffusion >>
rect 516 249 517 250 
<< pdiffusion >>
rect 517 249 518 250 
<< pdiffusion >>
rect 518 249 519 250 
<< pdiffusion >>
rect 519 249 520 250 
<< pdiffusion >>
rect 520 249 521 250 
<< pdiffusion >>
rect 521 249 522 250 
<< m1 >>
rect 523 249 524 250 
<< pdiffusion >>
rect 12 250 13 251 
<< pdiffusion >>
rect 13 250 14 251 
<< pdiffusion >>
rect 14 250 15 251 
<< pdiffusion >>
rect 15 250 16 251 
<< pdiffusion >>
rect 16 250 17 251 
<< pdiffusion >>
rect 17 250 18 251 
<< m1 >>
rect 19 250 20 251 
<< m1 >>
rect 22 250 23 251 
<< pdiffusion >>
rect 30 250 31 251 
<< pdiffusion >>
rect 31 250 32 251 
<< pdiffusion >>
rect 32 250 33 251 
<< pdiffusion >>
rect 33 250 34 251 
<< pdiffusion >>
rect 34 250 35 251 
<< pdiffusion >>
rect 35 250 36 251 
<< m1 >>
rect 44 250 45 251 
<< pdiffusion >>
rect 48 250 49 251 
<< pdiffusion >>
rect 49 250 50 251 
<< pdiffusion >>
rect 50 250 51 251 
<< pdiffusion >>
rect 51 250 52 251 
<< pdiffusion >>
rect 52 250 53 251 
<< pdiffusion >>
rect 53 250 54 251 
<< m1 >>
rect 55 250 56 251 
<< m2 >>
rect 56 250 57 251 
<< m1 >>
rect 64 250 65 251 
<< pdiffusion >>
rect 66 250 67 251 
<< pdiffusion >>
rect 67 250 68 251 
<< pdiffusion >>
rect 68 250 69 251 
<< pdiffusion >>
rect 69 250 70 251 
<< pdiffusion >>
rect 70 250 71 251 
<< pdiffusion >>
rect 71 250 72 251 
<< pdiffusion >>
rect 84 250 85 251 
<< pdiffusion >>
rect 85 250 86 251 
<< pdiffusion >>
rect 86 250 87 251 
<< pdiffusion >>
rect 87 250 88 251 
<< pdiffusion >>
rect 88 250 89 251 
<< pdiffusion >>
rect 89 250 90 251 
<< pdiffusion >>
rect 102 250 103 251 
<< pdiffusion >>
rect 103 250 104 251 
<< pdiffusion >>
rect 104 250 105 251 
<< pdiffusion >>
rect 105 250 106 251 
<< pdiffusion >>
rect 106 250 107 251 
<< pdiffusion >>
rect 107 250 108 251 
<< m1 >>
rect 118 250 119 251 
<< pdiffusion >>
rect 120 250 121 251 
<< pdiffusion >>
rect 121 250 122 251 
<< pdiffusion >>
rect 122 250 123 251 
<< pdiffusion >>
rect 123 250 124 251 
<< pdiffusion >>
rect 124 250 125 251 
<< pdiffusion >>
rect 125 250 126 251 
<< m1 >>
rect 127 250 128 251 
<< pdiffusion >>
rect 138 250 139 251 
<< pdiffusion >>
rect 139 250 140 251 
<< pdiffusion >>
rect 140 250 141 251 
<< pdiffusion >>
rect 141 250 142 251 
<< pdiffusion >>
rect 142 250 143 251 
<< pdiffusion >>
rect 143 250 144 251 
<< m1 >>
rect 148 250 149 251 
<< pdiffusion >>
rect 156 250 157 251 
<< pdiffusion >>
rect 157 250 158 251 
<< pdiffusion >>
rect 158 250 159 251 
<< pdiffusion >>
rect 159 250 160 251 
<< pdiffusion >>
rect 160 250 161 251 
<< pdiffusion >>
rect 161 250 162 251 
<< m1 >>
rect 163 250 164 251 
<< m2 >>
rect 171 250 172 251 
<< m1 >>
rect 172 250 173 251 
<< pdiffusion >>
rect 174 250 175 251 
<< pdiffusion >>
rect 175 250 176 251 
<< pdiffusion >>
rect 176 250 177 251 
<< pdiffusion >>
rect 177 250 178 251 
<< pdiffusion >>
rect 178 250 179 251 
<< pdiffusion >>
rect 179 250 180 251 
<< m1 >>
rect 181 250 182 251 
<< m2 >>
rect 182 250 183 251 
<< m1 >>
rect 186 250 187 251 
<< m1 >>
rect 190 250 191 251 
<< pdiffusion >>
rect 192 250 193 251 
<< pdiffusion >>
rect 193 250 194 251 
<< pdiffusion >>
rect 194 250 195 251 
<< pdiffusion >>
rect 195 250 196 251 
<< pdiffusion >>
rect 196 250 197 251 
<< pdiffusion >>
rect 197 250 198 251 
<< m1 >>
rect 207 250 208 251 
<< pdiffusion >>
rect 210 250 211 251 
<< pdiffusion >>
rect 211 250 212 251 
<< pdiffusion >>
rect 212 250 213 251 
<< pdiffusion >>
rect 213 250 214 251 
<< pdiffusion >>
rect 214 250 215 251 
<< pdiffusion >>
rect 215 250 216 251 
<< m1 >>
rect 224 250 225 251 
<< m1 >>
rect 226 250 227 251 
<< pdiffusion >>
rect 228 250 229 251 
<< pdiffusion >>
rect 229 250 230 251 
<< pdiffusion >>
rect 230 250 231 251 
<< pdiffusion >>
rect 231 250 232 251 
<< pdiffusion >>
rect 232 250 233 251 
<< pdiffusion >>
rect 233 250 234 251 
<< m1 >>
rect 235 250 236 251 
<< m1 >>
rect 237 250 238 251 
<< pdiffusion >>
rect 246 250 247 251 
<< pdiffusion >>
rect 247 250 248 251 
<< pdiffusion >>
rect 248 250 249 251 
<< pdiffusion >>
rect 249 250 250 251 
<< pdiffusion >>
rect 250 250 251 251 
<< pdiffusion >>
rect 251 250 252 251 
<< m1 >>
rect 255 250 256 251 
<< m1 >>
rect 262 250 263 251 
<< m2 >>
rect 262 250 263 251 
<< pdiffusion >>
rect 264 250 265 251 
<< pdiffusion >>
rect 265 250 266 251 
<< pdiffusion >>
rect 266 250 267 251 
<< pdiffusion >>
rect 267 250 268 251 
<< pdiffusion >>
rect 268 250 269 251 
<< pdiffusion >>
rect 269 250 270 251 
<< m1 >>
rect 274 250 275 251 
<< m1 >>
rect 276 250 277 251 
<< pdiffusion >>
rect 300 250 301 251 
<< pdiffusion >>
rect 301 250 302 251 
<< pdiffusion >>
rect 302 250 303 251 
<< pdiffusion >>
rect 303 250 304 251 
<< pdiffusion >>
rect 304 250 305 251 
<< pdiffusion >>
rect 305 250 306 251 
<< m1 >>
rect 307 250 308 251 
<< m2 >>
rect 308 250 309 251 
<< pdiffusion >>
rect 318 250 319 251 
<< pdiffusion >>
rect 319 250 320 251 
<< pdiffusion >>
rect 320 250 321 251 
<< pdiffusion >>
rect 321 250 322 251 
<< pdiffusion >>
rect 322 250 323 251 
<< pdiffusion >>
rect 323 250 324 251 
<< m1 >>
rect 334 250 335 251 
<< pdiffusion >>
rect 336 250 337 251 
<< pdiffusion >>
rect 337 250 338 251 
<< pdiffusion >>
rect 338 250 339 251 
<< pdiffusion >>
rect 339 250 340 251 
<< pdiffusion >>
rect 340 250 341 251 
<< pdiffusion >>
rect 341 250 342 251 
<< m1 >>
rect 346 250 347 251 
<< m1 >>
rect 352 250 353 251 
<< pdiffusion >>
rect 372 250 373 251 
<< pdiffusion >>
rect 373 250 374 251 
<< pdiffusion >>
rect 374 250 375 251 
<< pdiffusion >>
rect 375 250 376 251 
<< pdiffusion >>
rect 376 250 377 251 
<< pdiffusion >>
rect 377 250 378 251 
<< m1 >>
rect 379 250 380 251 
<< m2 >>
rect 380 250 381 251 
<< pdiffusion >>
rect 390 250 391 251 
<< pdiffusion >>
rect 391 250 392 251 
<< pdiffusion >>
rect 392 250 393 251 
<< pdiffusion >>
rect 393 250 394 251 
<< pdiffusion >>
rect 394 250 395 251 
<< pdiffusion >>
rect 395 250 396 251 
<< pdiffusion >>
rect 408 250 409 251 
<< pdiffusion >>
rect 409 250 410 251 
<< pdiffusion >>
rect 410 250 411 251 
<< pdiffusion >>
rect 411 250 412 251 
<< pdiffusion >>
rect 412 250 413 251 
<< pdiffusion >>
rect 413 250 414 251 
<< m1 >>
rect 416 250 417 251 
<< m1 >>
rect 419 250 420 251 
<< m1 >>
rect 421 250 422 251 
<< m2 >>
rect 422 250 423 251 
<< pdiffusion >>
rect 426 250 427 251 
<< pdiffusion >>
rect 427 250 428 251 
<< pdiffusion >>
rect 428 250 429 251 
<< pdiffusion >>
rect 429 250 430 251 
<< pdiffusion >>
rect 430 250 431 251 
<< pdiffusion >>
rect 431 250 432 251 
<< m1 >>
rect 434 250 435 251 
<< m1 >>
rect 442 250 443 251 
<< m2 >>
rect 442 250 443 251 
<< pdiffusion >>
rect 444 250 445 251 
<< pdiffusion >>
rect 445 250 446 251 
<< pdiffusion >>
rect 446 250 447 251 
<< pdiffusion >>
rect 447 250 448 251 
<< pdiffusion >>
rect 448 250 449 251 
<< pdiffusion >>
rect 449 250 450 251 
<< pdiffusion >>
rect 462 250 463 251 
<< pdiffusion >>
rect 463 250 464 251 
<< pdiffusion >>
rect 464 250 465 251 
<< pdiffusion >>
rect 465 250 466 251 
<< pdiffusion >>
rect 466 250 467 251 
<< pdiffusion >>
rect 467 250 468 251 
<< pdiffusion >>
rect 480 250 481 251 
<< pdiffusion >>
rect 481 250 482 251 
<< pdiffusion >>
rect 482 250 483 251 
<< pdiffusion >>
rect 483 250 484 251 
<< pdiffusion >>
rect 484 250 485 251 
<< pdiffusion >>
rect 485 250 486 251 
<< m1 >>
rect 496 250 497 251 
<< pdiffusion >>
rect 498 250 499 251 
<< pdiffusion >>
rect 499 250 500 251 
<< pdiffusion >>
rect 500 250 501 251 
<< pdiffusion >>
rect 501 250 502 251 
<< pdiffusion >>
rect 502 250 503 251 
<< pdiffusion >>
rect 503 250 504 251 
<< pdiffusion >>
rect 516 250 517 251 
<< pdiffusion >>
rect 517 250 518 251 
<< pdiffusion >>
rect 518 250 519 251 
<< pdiffusion >>
rect 519 250 520 251 
<< pdiffusion >>
rect 520 250 521 251 
<< pdiffusion >>
rect 521 250 522 251 
<< m1 >>
rect 523 250 524 251 
<< pdiffusion >>
rect 12 251 13 252 
<< pdiffusion >>
rect 13 251 14 252 
<< pdiffusion >>
rect 14 251 15 252 
<< pdiffusion >>
rect 15 251 16 252 
<< pdiffusion >>
rect 16 251 17 252 
<< pdiffusion >>
rect 17 251 18 252 
<< m1 >>
rect 19 251 20 252 
<< m1 >>
rect 22 251 23 252 
<< pdiffusion >>
rect 30 251 31 252 
<< pdiffusion >>
rect 31 251 32 252 
<< pdiffusion >>
rect 32 251 33 252 
<< pdiffusion >>
rect 33 251 34 252 
<< pdiffusion >>
rect 34 251 35 252 
<< pdiffusion >>
rect 35 251 36 252 
<< m1 >>
rect 44 251 45 252 
<< pdiffusion >>
rect 48 251 49 252 
<< pdiffusion >>
rect 49 251 50 252 
<< pdiffusion >>
rect 50 251 51 252 
<< pdiffusion >>
rect 51 251 52 252 
<< m1 >>
rect 52 251 53 252 
<< pdiffusion >>
rect 52 251 53 252 
<< pdiffusion >>
rect 53 251 54 252 
<< m1 >>
rect 55 251 56 252 
<< m2 >>
rect 56 251 57 252 
<< m1 >>
rect 64 251 65 252 
<< pdiffusion >>
rect 66 251 67 252 
<< pdiffusion >>
rect 67 251 68 252 
<< pdiffusion >>
rect 68 251 69 252 
<< pdiffusion >>
rect 69 251 70 252 
<< pdiffusion >>
rect 70 251 71 252 
<< pdiffusion >>
rect 71 251 72 252 
<< pdiffusion >>
rect 84 251 85 252 
<< pdiffusion >>
rect 85 251 86 252 
<< pdiffusion >>
rect 86 251 87 252 
<< pdiffusion >>
rect 87 251 88 252 
<< pdiffusion >>
rect 88 251 89 252 
<< pdiffusion >>
rect 89 251 90 252 
<< pdiffusion >>
rect 102 251 103 252 
<< pdiffusion >>
rect 103 251 104 252 
<< pdiffusion >>
rect 104 251 105 252 
<< pdiffusion >>
rect 105 251 106 252 
<< pdiffusion >>
rect 106 251 107 252 
<< pdiffusion >>
rect 107 251 108 252 
<< m1 >>
rect 118 251 119 252 
<< pdiffusion >>
rect 120 251 121 252 
<< pdiffusion >>
rect 121 251 122 252 
<< pdiffusion >>
rect 122 251 123 252 
<< pdiffusion >>
rect 123 251 124 252 
<< pdiffusion >>
rect 124 251 125 252 
<< pdiffusion >>
rect 125 251 126 252 
<< m1 >>
rect 127 251 128 252 
<< pdiffusion >>
rect 138 251 139 252 
<< pdiffusion >>
rect 139 251 140 252 
<< pdiffusion >>
rect 140 251 141 252 
<< pdiffusion >>
rect 141 251 142 252 
<< m1 >>
rect 142 251 143 252 
<< pdiffusion >>
rect 142 251 143 252 
<< pdiffusion >>
rect 143 251 144 252 
<< m1 >>
rect 148 251 149 252 
<< pdiffusion >>
rect 156 251 157 252 
<< pdiffusion >>
rect 157 251 158 252 
<< pdiffusion >>
rect 158 251 159 252 
<< pdiffusion >>
rect 159 251 160 252 
<< pdiffusion >>
rect 160 251 161 252 
<< pdiffusion >>
rect 161 251 162 252 
<< m1 >>
rect 163 251 164 252 
<< m2 >>
rect 171 251 172 252 
<< m1 >>
rect 172 251 173 252 
<< pdiffusion >>
rect 174 251 175 252 
<< pdiffusion >>
rect 175 251 176 252 
<< pdiffusion >>
rect 176 251 177 252 
<< pdiffusion >>
rect 177 251 178 252 
<< pdiffusion >>
rect 178 251 179 252 
<< pdiffusion >>
rect 179 251 180 252 
<< m1 >>
rect 181 251 182 252 
<< m2 >>
rect 182 251 183 252 
<< m1 >>
rect 186 251 187 252 
<< m1 >>
rect 190 251 191 252 
<< pdiffusion >>
rect 192 251 193 252 
<< pdiffusion >>
rect 193 251 194 252 
<< pdiffusion >>
rect 194 251 195 252 
<< pdiffusion >>
rect 195 251 196 252 
<< pdiffusion >>
rect 196 251 197 252 
<< pdiffusion >>
rect 197 251 198 252 
<< m1 >>
rect 207 251 208 252 
<< pdiffusion >>
rect 210 251 211 252 
<< m1 >>
rect 211 251 212 252 
<< pdiffusion >>
rect 211 251 212 252 
<< pdiffusion >>
rect 212 251 213 252 
<< pdiffusion >>
rect 213 251 214 252 
<< m1 >>
rect 214 251 215 252 
<< pdiffusion >>
rect 214 251 215 252 
<< pdiffusion >>
rect 215 251 216 252 
<< m1 >>
rect 224 251 225 252 
<< m2 >>
rect 224 251 225 252 
<< m2c >>
rect 224 251 225 252 
<< m1 >>
rect 224 251 225 252 
<< m2 >>
rect 224 251 225 252 
<< m2 >>
rect 225 251 226 252 
<< m1 >>
rect 226 251 227 252 
<< m2 >>
rect 226 251 227 252 
<< pdiffusion >>
rect 228 251 229 252 
<< pdiffusion >>
rect 229 251 230 252 
<< pdiffusion >>
rect 230 251 231 252 
<< pdiffusion >>
rect 231 251 232 252 
<< m1 >>
rect 232 251 233 252 
<< pdiffusion >>
rect 232 251 233 252 
<< pdiffusion >>
rect 233 251 234 252 
<< m1 >>
rect 235 251 236 252 
<< m1 >>
rect 237 251 238 252 
<< pdiffusion >>
rect 246 251 247 252 
<< m1 >>
rect 247 251 248 252 
<< pdiffusion >>
rect 247 251 248 252 
<< pdiffusion >>
rect 248 251 249 252 
<< pdiffusion >>
rect 249 251 250 252 
<< m1 >>
rect 250 251 251 252 
<< pdiffusion >>
rect 250 251 251 252 
<< pdiffusion >>
rect 251 251 252 252 
<< m1 >>
rect 255 251 256 252 
<< m1 >>
rect 262 251 263 252 
<< m2 >>
rect 262 251 263 252 
<< pdiffusion >>
rect 264 251 265 252 
<< m1 >>
rect 265 251 266 252 
<< pdiffusion >>
rect 265 251 266 252 
<< pdiffusion >>
rect 266 251 267 252 
<< pdiffusion >>
rect 267 251 268 252 
<< pdiffusion >>
rect 268 251 269 252 
<< pdiffusion >>
rect 269 251 270 252 
<< m1 >>
rect 274 251 275 252 
<< m1 >>
rect 276 251 277 252 
<< pdiffusion >>
rect 300 251 301 252 
<< pdiffusion >>
rect 301 251 302 252 
<< pdiffusion >>
rect 302 251 303 252 
<< pdiffusion >>
rect 303 251 304 252 
<< pdiffusion >>
rect 304 251 305 252 
<< pdiffusion >>
rect 305 251 306 252 
<< m1 >>
rect 307 251 308 252 
<< m2 >>
rect 308 251 309 252 
<< pdiffusion >>
rect 318 251 319 252 
<< pdiffusion >>
rect 319 251 320 252 
<< pdiffusion >>
rect 320 251 321 252 
<< pdiffusion >>
rect 321 251 322 252 
<< pdiffusion >>
rect 322 251 323 252 
<< pdiffusion >>
rect 323 251 324 252 
<< m1 >>
rect 334 251 335 252 
<< pdiffusion >>
rect 336 251 337 252 
<< m1 >>
rect 337 251 338 252 
<< pdiffusion >>
rect 337 251 338 252 
<< pdiffusion >>
rect 338 251 339 252 
<< pdiffusion >>
rect 339 251 340 252 
<< pdiffusion >>
rect 340 251 341 252 
<< pdiffusion >>
rect 341 251 342 252 
<< m1 >>
rect 346 251 347 252 
<< m1 >>
rect 352 251 353 252 
<< pdiffusion >>
rect 372 251 373 252 
<< pdiffusion >>
rect 373 251 374 252 
<< pdiffusion >>
rect 374 251 375 252 
<< pdiffusion >>
rect 375 251 376 252 
<< pdiffusion >>
rect 376 251 377 252 
<< pdiffusion >>
rect 377 251 378 252 
<< m1 >>
rect 379 251 380 252 
<< m2 >>
rect 380 251 381 252 
<< pdiffusion >>
rect 390 251 391 252 
<< pdiffusion >>
rect 391 251 392 252 
<< pdiffusion >>
rect 392 251 393 252 
<< pdiffusion >>
rect 393 251 394 252 
<< pdiffusion >>
rect 394 251 395 252 
<< pdiffusion >>
rect 395 251 396 252 
<< pdiffusion >>
rect 408 251 409 252 
<< m1 >>
rect 409 251 410 252 
<< pdiffusion >>
rect 409 251 410 252 
<< pdiffusion >>
rect 410 251 411 252 
<< pdiffusion >>
rect 411 251 412 252 
<< m1 >>
rect 412 251 413 252 
<< pdiffusion >>
rect 412 251 413 252 
<< pdiffusion >>
rect 413 251 414 252 
<< m1 >>
rect 416 251 417 252 
<< m1 >>
rect 419 251 420 252 
<< m1 >>
rect 421 251 422 252 
<< m2 >>
rect 422 251 423 252 
<< pdiffusion >>
rect 426 251 427 252 
<< pdiffusion >>
rect 427 251 428 252 
<< pdiffusion >>
rect 428 251 429 252 
<< pdiffusion >>
rect 429 251 430 252 
<< m1 >>
rect 430 251 431 252 
<< pdiffusion >>
rect 430 251 431 252 
<< pdiffusion >>
rect 431 251 432 252 
<< m1 >>
rect 434 251 435 252 
<< m2 >>
rect 434 251 435 252 
<< m2c >>
rect 434 251 435 252 
<< m1 >>
rect 434 251 435 252 
<< m2 >>
rect 434 251 435 252 
<< m1 >>
rect 442 251 443 252 
<< m2 >>
rect 442 251 443 252 
<< pdiffusion >>
rect 444 251 445 252 
<< pdiffusion >>
rect 445 251 446 252 
<< pdiffusion >>
rect 446 251 447 252 
<< pdiffusion >>
rect 447 251 448 252 
<< pdiffusion >>
rect 448 251 449 252 
<< pdiffusion >>
rect 449 251 450 252 
<< pdiffusion >>
rect 462 251 463 252 
<< pdiffusion >>
rect 463 251 464 252 
<< pdiffusion >>
rect 464 251 465 252 
<< pdiffusion >>
rect 465 251 466 252 
<< pdiffusion >>
rect 466 251 467 252 
<< pdiffusion >>
rect 467 251 468 252 
<< pdiffusion >>
rect 480 251 481 252 
<< pdiffusion >>
rect 481 251 482 252 
<< pdiffusion >>
rect 482 251 483 252 
<< pdiffusion >>
rect 483 251 484 252 
<< pdiffusion >>
rect 484 251 485 252 
<< pdiffusion >>
rect 485 251 486 252 
<< m1 >>
rect 496 251 497 252 
<< pdiffusion >>
rect 498 251 499 252 
<< pdiffusion >>
rect 499 251 500 252 
<< pdiffusion >>
rect 500 251 501 252 
<< pdiffusion >>
rect 501 251 502 252 
<< pdiffusion >>
rect 502 251 503 252 
<< pdiffusion >>
rect 503 251 504 252 
<< pdiffusion >>
rect 516 251 517 252 
<< pdiffusion >>
rect 517 251 518 252 
<< pdiffusion >>
rect 518 251 519 252 
<< pdiffusion >>
rect 519 251 520 252 
<< pdiffusion >>
rect 520 251 521 252 
<< pdiffusion >>
rect 521 251 522 252 
<< m1 >>
rect 523 251 524 252 
<< m1 >>
rect 19 252 20 253 
<< m1 >>
rect 22 252 23 253 
<< m1 >>
rect 44 252 45 253 
<< m1 >>
rect 52 252 53 253 
<< m1 >>
rect 55 252 56 253 
<< m2 >>
rect 56 252 57 253 
<< m1 >>
rect 64 252 65 253 
<< m1 >>
rect 118 252 119 253 
<< m1 >>
rect 127 252 128 253 
<< m1 >>
rect 142 252 143 253 
<< m1 >>
rect 148 252 149 253 
<< m1 >>
rect 163 252 164 253 
<< m2 >>
rect 171 252 172 253 
<< m1 >>
rect 172 252 173 253 
<< m1 >>
rect 181 252 182 253 
<< m2 >>
rect 182 252 183 253 
<< m1 >>
rect 186 252 187 253 
<< m1 >>
rect 190 252 191 253 
<< m1 >>
rect 207 252 208 253 
<< m1 >>
rect 211 252 212 253 
<< m1 >>
rect 214 252 215 253 
<< m1 >>
rect 226 252 227 253 
<< m2 >>
rect 226 252 227 253 
<< m1 >>
rect 232 252 233 253 
<< m1 >>
rect 235 252 236 253 
<< m1 >>
rect 237 252 238 253 
<< m1 >>
rect 247 252 248 253 
<< m1 >>
rect 250 252 251 253 
<< m1 >>
rect 255 252 256 253 
<< m1 >>
rect 262 252 263 253 
<< m2 >>
rect 262 252 263 253 
<< m1 >>
rect 265 252 266 253 
<< m1 >>
rect 274 252 275 253 
<< m1 >>
rect 276 252 277 253 
<< m1 >>
rect 307 252 308 253 
<< m2 >>
rect 308 252 309 253 
<< m1 >>
rect 334 252 335 253 
<< m1 >>
rect 337 252 338 253 
<< m1 >>
rect 346 252 347 253 
<< m1 >>
rect 352 252 353 253 
<< m1 >>
rect 379 252 380 253 
<< m2 >>
rect 380 252 381 253 
<< m1 >>
rect 409 252 410 253 
<< m1 >>
rect 412 252 413 253 
<< m1 >>
rect 416 252 417 253 
<< m1 >>
rect 419 252 420 253 
<< m1 >>
rect 421 252 422 253 
<< m2 >>
rect 422 252 423 253 
<< m1 >>
rect 430 252 431 253 
<< m2 >>
rect 434 252 435 253 
<< m1 >>
rect 442 252 443 253 
<< m2 >>
rect 442 252 443 253 
<< m1 >>
rect 496 252 497 253 
<< m1 >>
rect 523 252 524 253 
<< m1 >>
rect 19 253 20 254 
<< m1 >>
rect 22 253 23 254 
<< m1 >>
rect 44 253 45 254 
<< m1 >>
rect 52 253 53 254 
<< m1 >>
rect 53 253 54 254 
<< m2 >>
rect 53 253 54 254 
<< m2c >>
rect 53 253 54 254 
<< m1 >>
rect 53 253 54 254 
<< m2 >>
rect 53 253 54 254 
<< m2 >>
rect 54 253 55 254 
<< m1 >>
rect 55 253 56 254 
<< m2 >>
rect 55 253 56 254 
<< m2 >>
rect 56 253 57 254 
<< m1 >>
rect 64 253 65 254 
<< m1 >>
rect 118 253 119 254 
<< m1 >>
rect 127 253 128 254 
<< m1 >>
rect 142 253 143 254 
<< m1 >>
rect 148 253 149 254 
<< m1 >>
rect 163 253 164 254 
<< m2 >>
rect 171 253 172 254 
<< m1 >>
rect 172 253 173 254 
<< m1 >>
rect 179 253 180 254 
<< m2 >>
rect 179 253 180 254 
<< m2c >>
rect 179 253 180 254 
<< m1 >>
rect 179 253 180 254 
<< m2 >>
rect 179 253 180 254 
<< m2 >>
rect 180 253 181 254 
<< m1 >>
rect 181 253 182 254 
<< m2 >>
rect 181 253 182 254 
<< m2 >>
rect 182 253 183 254 
<< m1 >>
rect 186 253 187 254 
<< m1 >>
rect 190 253 191 254 
<< m1 >>
rect 207 253 208 254 
<< m1 >>
rect 211 253 212 254 
<< m1 >>
rect 214 253 215 254 
<< m1 >>
rect 215 253 216 254 
<< m1 >>
rect 216 253 217 254 
<< m1 >>
rect 217 253 218 254 
<< m1 >>
rect 218 253 219 254 
<< m1 >>
rect 219 253 220 254 
<< m1 >>
rect 220 253 221 254 
<< m1 >>
rect 221 253 222 254 
<< m1 >>
rect 222 253 223 254 
<< m1 >>
rect 223 253 224 254 
<< m1 >>
rect 224 253 225 254 
<< m1 >>
rect 225 253 226 254 
<< m1 >>
rect 226 253 227 254 
<< m2 >>
rect 226 253 227 254 
<< m1 >>
rect 232 253 233 254 
<< m1 >>
rect 235 253 236 254 
<< m1 >>
rect 237 253 238 254 
<< m1 >>
rect 247 253 248 254 
<< m1 >>
rect 250 253 251 254 
<< m1 >>
rect 255 253 256 254 
<< m1 >>
rect 262 253 263 254 
<< m2 >>
rect 262 253 263 254 
<< m1 >>
rect 265 253 266 254 
<< m1 >>
rect 274 253 275 254 
<< m1 >>
rect 276 253 277 254 
<< m1 >>
rect 307 253 308 254 
<< m2 >>
rect 308 253 309 254 
<< m1 >>
rect 334 253 335 254 
<< m1 >>
rect 337 253 338 254 
<< m1 >>
rect 346 253 347 254 
<< m1 >>
rect 352 253 353 254 
<< m1 >>
rect 377 253 378 254 
<< m2 >>
rect 377 253 378 254 
<< m2c >>
rect 377 253 378 254 
<< m1 >>
rect 377 253 378 254 
<< m2 >>
rect 377 253 378 254 
<< m2 >>
rect 378 253 379 254 
<< m1 >>
rect 379 253 380 254 
<< m2 >>
rect 379 253 380 254 
<< m2 >>
rect 380 253 381 254 
<< m1 >>
rect 409 253 410 254 
<< m1 >>
rect 412 253 413 254 
<< m2 >>
rect 413 253 414 254 
<< m1 >>
rect 414 253 415 254 
<< m2 >>
rect 414 253 415 254 
<< m2c >>
rect 414 253 415 254 
<< m1 >>
rect 414 253 415 254 
<< m2 >>
rect 414 253 415 254 
<< m2 >>
rect 415 253 416 254 
<< m1 >>
rect 416 253 417 254 
<< m2 >>
rect 416 253 417 254 
<< m2 >>
rect 417 253 418 254 
<< m2 >>
rect 418 253 419 254 
<< m1 >>
rect 419 253 420 254 
<< m2 >>
rect 419 253 420 254 
<< m2 >>
rect 420 253 421 254 
<< m1 >>
rect 421 253 422 254 
<< m2 >>
rect 421 253 422 254 
<< m2 >>
rect 422 253 423 254 
<< m1 >>
rect 430 253 431 254 
<< m2 >>
rect 431 253 432 254 
<< m1 >>
rect 432 253 433 254 
<< m2 >>
rect 432 253 433 254 
<< m2c >>
rect 432 253 433 254 
<< m1 >>
rect 432 253 433 254 
<< m2 >>
rect 432 253 433 254 
<< m1 >>
rect 433 253 434 254 
<< m1 >>
rect 434 253 435 254 
<< m2 >>
rect 434 253 435 254 
<< m1 >>
rect 435 253 436 254 
<< m1 >>
rect 436 253 437 254 
<< m1 >>
rect 437 253 438 254 
<< m1 >>
rect 438 253 439 254 
<< m1 >>
rect 439 253 440 254 
<< m1 >>
rect 440 253 441 254 
<< m1 >>
rect 441 253 442 254 
<< m1 >>
rect 442 253 443 254 
<< m2 >>
rect 442 253 443 254 
<< m1 >>
rect 496 253 497 254 
<< m1 >>
rect 523 253 524 254 
<< m1 >>
rect 19 254 20 255 
<< m1 >>
rect 22 254 23 255 
<< m1 >>
rect 44 254 45 255 
<< m1 >>
rect 55 254 56 255 
<< m1 >>
rect 64 254 65 255 
<< m1 >>
rect 118 254 119 255 
<< m1 >>
rect 127 254 128 255 
<< m1 >>
rect 142 254 143 255 
<< m1 >>
rect 148 254 149 255 
<< m1 >>
rect 163 254 164 255 
<< m2 >>
rect 171 254 172 255 
<< m1 >>
rect 172 254 173 255 
<< m1 >>
rect 177 254 178 255 
<< m1 >>
rect 178 254 179 255 
<< m1 >>
rect 179 254 180 255 
<< m1 >>
rect 181 254 182 255 
<< m1 >>
rect 186 254 187 255 
<< m1 >>
rect 190 254 191 255 
<< m1 >>
rect 207 254 208 255 
<< m1 >>
rect 211 254 212 255 
<< m2 >>
rect 226 254 227 255 
<< m2 >>
rect 227 254 228 255 
<< m1 >>
rect 228 254 229 255 
<< m2 >>
rect 228 254 229 255 
<< m1 >>
rect 232 254 233 255 
<< m1 >>
rect 235 254 236 255 
<< m1 >>
rect 237 254 238 255 
<< m1 >>
rect 247 254 248 255 
<< m1 >>
rect 250 254 251 255 
<< m1 >>
rect 255 254 256 255 
<< m1 >>
rect 262 254 263 255 
<< m2 >>
rect 262 254 263 255 
<< m1 >>
rect 265 254 266 255 
<< m1 >>
rect 266 254 267 255 
<< m1 >>
rect 267 254 268 255 
<< m1 >>
rect 268 254 269 255 
<< m1 >>
rect 269 254 270 255 
<< m1 >>
rect 270 254 271 255 
<< m1 >>
rect 271 254 272 255 
<< m1 >>
rect 272 254 273 255 
<< m1 >>
rect 273 254 274 255 
<< m1 >>
rect 274 254 275 255 
<< m1 >>
rect 276 254 277 255 
<< m1 >>
rect 307 254 308 255 
<< m2 >>
rect 308 254 309 255 
<< m1 >>
rect 309 254 310 255 
<< m2 >>
rect 309 254 310 255 
<< m2c >>
rect 309 254 310 255 
<< m1 >>
rect 309 254 310 255 
<< m2 >>
rect 309 254 310 255 
<< m1 >>
rect 310 254 311 255 
<< m1 >>
rect 311 254 312 255 
<< m1 >>
rect 312 254 313 255 
<< m1 >>
rect 313 254 314 255 
<< m1 >>
rect 314 254 315 255 
<< m1 >>
rect 315 254 316 255 
<< m1 >>
rect 316 254 317 255 
<< m1 >>
rect 317 254 318 255 
<< m1 >>
rect 318 254 319 255 
<< m2 >>
rect 318 254 319 255 
<< m2c >>
rect 318 254 319 255 
<< m1 >>
rect 318 254 319 255 
<< m2 >>
rect 318 254 319 255 
<< m1 >>
rect 334 254 335 255 
<< m1 >>
rect 337 254 338 255 
<< m1 >>
rect 338 254 339 255 
<< m1 >>
rect 339 254 340 255 
<< m1 >>
rect 340 254 341 255 
<< m1 >>
rect 341 254 342 255 
<< m1 >>
rect 342 254 343 255 
<< m1 >>
rect 346 254 347 255 
<< m1 >>
rect 352 254 353 255 
<< m1 >>
rect 376 254 377 255 
<< m1 >>
rect 377 254 378 255 
<< m1 >>
rect 379 254 380 255 
<< m1 >>
rect 392 254 393 255 
<< m2 >>
rect 392 254 393 255 
<< m2c >>
rect 392 254 393 255 
<< m1 >>
rect 392 254 393 255 
<< m2 >>
rect 392 254 393 255 
<< m1 >>
rect 393 254 394 255 
<< m1 >>
rect 394 254 395 255 
<< m1 >>
rect 395 254 396 255 
<< m1 >>
rect 396 254 397 255 
<< m1 >>
rect 397 254 398 255 
<< m1 >>
rect 398 254 399 255 
<< m1 >>
rect 399 254 400 255 
<< m1 >>
rect 400 254 401 255 
<< m1 >>
rect 401 254 402 255 
<< m1 >>
rect 402 254 403 255 
<< m1 >>
rect 403 254 404 255 
<< m1 >>
rect 404 254 405 255 
<< m1 >>
rect 405 254 406 255 
<< m1 >>
rect 406 254 407 255 
<< m1 >>
rect 407 254 408 255 
<< m1 >>
rect 408 254 409 255 
<< m1 >>
rect 409 254 410 255 
<< m1 >>
rect 412 254 413 255 
<< m2 >>
rect 412 254 413 255 
<< m2 >>
rect 413 254 414 255 
<< m1 >>
rect 416 254 417 255 
<< m1 >>
rect 419 254 420 255 
<< m1 >>
rect 421 254 422 255 
<< m1 >>
rect 428 254 429 255 
<< m2 >>
rect 428 254 429 255 
<< m2c >>
rect 428 254 429 255 
<< m1 >>
rect 428 254 429 255 
<< m2 >>
rect 428 254 429 255 
<< m1 >>
rect 429 254 430 255 
<< m1 >>
rect 430 254 431 255 
<< m2 >>
rect 431 254 432 255 
<< m2 >>
rect 434 254 435 255 
<< m2 >>
rect 442 254 443 255 
<< m1 >>
rect 484 254 485 255 
<< m1 >>
rect 485 254 486 255 
<< m1 >>
rect 486 254 487 255 
<< m1 >>
rect 487 254 488 255 
<< m1 >>
rect 488 254 489 255 
<< m1 >>
rect 489 254 490 255 
<< m1 >>
rect 490 254 491 255 
<< m1 >>
rect 491 254 492 255 
<< m1 >>
rect 492 254 493 255 
<< m1 >>
rect 493 254 494 255 
<< m1 >>
rect 494 254 495 255 
<< m1 >>
rect 495 254 496 255 
<< m1 >>
rect 496 254 497 255 
<< m1 >>
rect 523 254 524 255 
<< m1 >>
rect 19 255 20 256 
<< m1 >>
rect 22 255 23 256 
<< m1 >>
rect 44 255 45 256 
<< m1 >>
rect 55 255 56 256 
<< m1 >>
rect 64 255 65 256 
<< m1 >>
rect 118 255 119 256 
<< m1 >>
rect 127 255 128 256 
<< m1 >>
rect 142 255 143 256 
<< m1 >>
rect 148 255 149 256 
<< m1 >>
rect 163 255 164 256 
<< m2 >>
rect 171 255 172 256 
<< m1 >>
rect 172 255 173 256 
<< m1 >>
rect 177 255 178 256 
<< m1 >>
rect 181 255 182 256 
<< m1 >>
rect 186 255 187 256 
<< m1 >>
rect 190 255 191 256 
<< m1 >>
rect 207 255 208 256 
<< m1 >>
rect 211 255 212 256 
<< m1 >>
rect 228 255 229 256 
<< m2 >>
rect 228 255 229 256 
<< m2c >>
rect 228 255 229 256 
<< m1 >>
rect 228 255 229 256 
<< m2 >>
rect 228 255 229 256 
<< m1 >>
rect 232 255 233 256 
<< m1 >>
rect 235 255 236 256 
<< m1 >>
rect 237 255 238 256 
<< m1 >>
rect 247 255 248 256 
<< m1 >>
rect 250 255 251 256 
<< m1 >>
rect 251 255 252 256 
<< m1 >>
rect 252 255 253 256 
<< m1 >>
rect 253 255 254 256 
<< m2 >>
rect 253 255 254 256 
<< m2c >>
rect 253 255 254 256 
<< m1 >>
rect 253 255 254 256 
<< m2 >>
rect 253 255 254 256 
<< m2 >>
rect 254 255 255 256 
<< m1 >>
rect 255 255 256 256 
<< m2 >>
rect 255 255 256 256 
<< m2 >>
rect 256 255 257 256 
<< m1 >>
rect 257 255 258 256 
<< m2 >>
rect 257 255 258 256 
<< m2c >>
rect 257 255 258 256 
<< m1 >>
rect 257 255 258 256 
<< m2 >>
rect 257 255 258 256 
<< m1 >>
rect 258 255 259 256 
<< m1 >>
rect 259 255 260 256 
<< m1 >>
rect 262 255 263 256 
<< m2 >>
rect 262 255 263 256 
<< m1 >>
rect 276 255 277 256 
<< m2 >>
rect 276 255 277 256 
<< m2c >>
rect 276 255 277 256 
<< m1 >>
rect 276 255 277 256 
<< m2 >>
rect 276 255 277 256 
<< m1 >>
rect 307 255 308 256 
<< m2 >>
rect 318 255 319 256 
<< m1 >>
rect 334 255 335 256 
<< m1 >>
rect 342 255 343 256 
<< m1 >>
rect 346 255 347 256 
<< m1 >>
rect 352 255 353 256 
<< m1 >>
rect 376 255 377 256 
<< m1 >>
rect 379 255 380 256 
<< m2 >>
rect 392 255 393 256 
<< m1 >>
rect 412 255 413 256 
<< m2 >>
rect 412 255 413 256 
<< m1 >>
rect 416 255 417 256 
<< m1 >>
rect 419 255 420 256 
<< m1 >>
rect 421 255 422 256 
<< m2 >>
rect 428 255 429 256 
<< m2 >>
rect 431 255 432 256 
<< m1 >>
rect 434 255 435 256 
<< m2 >>
rect 434 255 435 256 
<< m2c >>
rect 434 255 435 256 
<< m1 >>
rect 434 255 435 256 
<< m2 >>
rect 434 255 435 256 
<< m1 >>
rect 435 255 436 256 
<< m1 >>
rect 436 255 437 256 
<< m1 >>
rect 437 255 438 256 
<< m1 >>
rect 442 255 443 256 
<< m2 >>
rect 442 255 443 256 
<< m2c >>
rect 442 255 443 256 
<< m1 >>
rect 442 255 443 256 
<< m2 >>
rect 442 255 443 256 
<< m1 >>
rect 484 255 485 256 
<< m1 >>
rect 523 255 524 256 
<< m1 >>
rect 19 256 20 257 
<< m1 >>
rect 22 256 23 257 
<< m1 >>
rect 44 256 45 257 
<< m1 >>
rect 55 256 56 257 
<< m1 >>
rect 64 256 65 257 
<< m1 >>
rect 118 256 119 257 
<< m1 >>
rect 127 256 128 257 
<< m1 >>
rect 128 256 129 257 
<< m1 >>
rect 129 256 130 257 
<< m1 >>
rect 130 256 131 257 
<< m1 >>
rect 131 256 132 257 
<< m1 >>
rect 132 256 133 257 
<< m1 >>
rect 133 256 134 257 
<< m1 >>
rect 134 256 135 257 
<< m1 >>
rect 135 256 136 257 
<< m1 >>
rect 136 256 137 257 
<< m1 >>
rect 137 256 138 257 
<< m1 >>
rect 138 256 139 257 
<< m1 >>
rect 139 256 140 257 
<< m1 >>
rect 140 256 141 257 
<< m1 >>
rect 141 256 142 257 
<< m1 >>
rect 142 256 143 257 
<< m1 >>
rect 148 256 149 257 
<< m1 >>
rect 163 256 164 257 
<< m2 >>
rect 171 256 172 257 
<< m1 >>
rect 172 256 173 257 
<< m1 >>
rect 177 256 178 257 
<< m1 >>
rect 181 256 182 257 
<< m1 >>
rect 186 256 187 257 
<< m1 >>
rect 190 256 191 257 
<< m1 >>
rect 207 256 208 257 
<< m1 >>
rect 211 256 212 257 
<< m2 >>
rect 228 256 229 257 
<< m1 >>
rect 232 256 233 257 
<< m1 >>
rect 235 256 236 257 
<< m1 >>
rect 237 256 238 257 
<< m1 >>
rect 247 256 248 257 
<< m1 >>
rect 255 256 256 257 
<< m1 >>
rect 259 256 260 257 
<< m1 >>
rect 262 256 263 257 
<< m2 >>
rect 262 256 263 257 
<< m2 >>
rect 264 256 265 257 
<< m2 >>
rect 265 256 266 257 
<< m2 >>
rect 266 256 267 257 
<< m2 >>
rect 267 256 268 257 
<< m2 >>
rect 268 256 269 257 
<< m2 >>
rect 269 256 270 257 
<< m2 >>
rect 270 256 271 257 
<< m2 >>
rect 271 256 272 257 
<< m2 >>
rect 272 256 273 257 
<< m2 >>
rect 273 256 274 257 
<< m2 >>
rect 274 256 275 257 
<< m2 >>
rect 275 256 276 257 
<< m2 >>
rect 276 256 277 257 
<< m1 >>
rect 280 256 281 257 
<< m1 >>
rect 281 256 282 257 
<< m1 >>
rect 282 256 283 257 
<< m1 >>
rect 283 256 284 257 
<< m1 >>
rect 284 256 285 257 
<< m1 >>
rect 285 256 286 257 
<< m1 >>
rect 286 256 287 257 
<< m1 >>
rect 287 256 288 257 
<< m1 >>
rect 288 256 289 257 
<< m1 >>
rect 289 256 290 257 
<< m1 >>
rect 290 256 291 257 
<< m1 >>
rect 291 256 292 257 
<< m1 >>
rect 292 256 293 257 
<< m1 >>
rect 293 256 294 257 
<< m1 >>
rect 294 256 295 257 
<< m1 >>
rect 295 256 296 257 
<< m1 >>
rect 296 256 297 257 
<< m1 >>
rect 297 256 298 257 
<< m1 >>
rect 298 256 299 257 
<< m1 >>
rect 299 256 300 257 
<< m1 >>
rect 300 256 301 257 
<< m1 >>
rect 301 256 302 257 
<< m1 >>
rect 302 256 303 257 
<< m1 >>
rect 303 256 304 257 
<< m1 >>
rect 304 256 305 257 
<< m1 >>
rect 305 256 306 257 
<< m2 >>
rect 305 256 306 257 
<< m2c >>
rect 305 256 306 257 
<< m1 >>
rect 305 256 306 257 
<< m2 >>
rect 305 256 306 257 
<< m2 >>
rect 306 256 307 257 
<< m1 >>
rect 307 256 308 257 
<< m2 >>
rect 307 256 308 257 
<< m2 >>
rect 308 256 309 257 
<< m1 >>
rect 309 256 310 257 
<< m2 >>
rect 309 256 310 257 
<< m2c >>
rect 309 256 310 257 
<< m1 >>
rect 309 256 310 257 
<< m2 >>
rect 309 256 310 257 
<< m1 >>
rect 310 256 311 257 
<< m1 >>
rect 311 256 312 257 
<< m1 >>
rect 312 256 313 257 
<< m1 >>
rect 313 256 314 257 
<< m1 >>
rect 314 256 315 257 
<< m1 >>
rect 315 256 316 257 
<< m1 >>
rect 316 256 317 257 
<< m1 >>
rect 317 256 318 257 
<< m1 >>
rect 318 256 319 257 
<< m2 >>
rect 318 256 319 257 
<< m1 >>
rect 319 256 320 257 
<< m1 >>
rect 320 256 321 257 
<< m1 >>
rect 321 256 322 257 
<< m1 >>
rect 322 256 323 257 
<< m1 >>
rect 323 256 324 257 
<< m1 >>
rect 324 256 325 257 
<< m1 >>
rect 325 256 326 257 
<< m1 >>
rect 326 256 327 257 
<< m1 >>
rect 327 256 328 257 
<< m1 >>
rect 328 256 329 257 
<< m1 >>
rect 329 256 330 257 
<< m1 >>
rect 330 256 331 257 
<< m1 >>
rect 331 256 332 257 
<< m1 >>
rect 332 256 333 257 
<< m1 >>
rect 333 256 334 257 
<< m1 >>
rect 334 256 335 257 
<< m1 >>
rect 342 256 343 257 
<< m1 >>
rect 346 256 347 257 
<< m1 >>
rect 352 256 353 257 
<< m1 >>
rect 376 256 377 257 
<< m1 >>
rect 379 256 380 257 
<< m1 >>
rect 380 256 381 257 
<< m1 >>
rect 381 256 382 257 
<< m1 >>
rect 382 256 383 257 
<< m1 >>
rect 383 256 384 257 
<< m1 >>
rect 384 256 385 257 
<< m1 >>
rect 385 256 386 257 
<< m1 >>
rect 386 256 387 257 
<< m1 >>
rect 387 256 388 257 
<< m1 >>
rect 388 256 389 257 
<< m1 >>
rect 389 256 390 257 
<< m1 >>
rect 390 256 391 257 
<< m1 >>
rect 391 256 392 257 
<< m1 >>
rect 392 256 393 257 
<< m2 >>
rect 392 256 393 257 
<< m1 >>
rect 393 256 394 257 
<< m1 >>
rect 394 256 395 257 
<< m1 >>
rect 395 256 396 257 
<< m1 >>
rect 396 256 397 257 
<< m1 >>
rect 397 256 398 257 
<< m1 >>
rect 398 256 399 257 
<< m1 >>
rect 399 256 400 257 
<< m1 >>
rect 400 256 401 257 
<< m1 >>
rect 401 256 402 257 
<< m1 >>
rect 402 256 403 257 
<< m1 >>
rect 403 256 404 257 
<< m1 >>
rect 404 256 405 257 
<< m1 >>
rect 405 256 406 257 
<< m1 >>
rect 406 256 407 257 
<< m1 >>
rect 407 256 408 257 
<< m1 >>
rect 408 256 409 257 
<< m1 >>
rect 409 256 410 257 
<< m1 >>
rect 410 256 411 257 
<< m1 >>
rect 411 256 412 257 
<< m1 >>
rect 412 256 413 257 
<< m2 >>
rect 412 256 413 257 
<< m1 >>
rect 416 256 417 257 
<< m1 >>
rect 419 256 420 257 
<< m1 >>
rect 421 256 422 257 
<< m1 >>
rect 422 256 423 257 
<< m1 >>
rect 423 256 424 257 
<< m1 >>
rect 424 256 425 257 
<< m1 >>
rect 425 256 426 257 
<< m1 >>
rect 426 256 427 257 
<< m1 >>
rect 427 256 428 257 
<< m1 >>
rect 428 256 429 257 
<< m2 >>
rect 428 256 429 257 
<< m1 >>
rect 429 256 430 257 
<< m1 >>
rect 430 256 431 257 
<< m2 >>
rect 431 256 432 257 
<< m1 >>
rect 437 256 438 257 
<< m1 >>
rect 442 256 443 257 
<< m1 >>
rect 484 256 485 257 
<< m1 >>
rect 523 256 524 257 
<< m1 >>
rect 19 257 20 258 
<< m1 >>
rect 22 257 23 258 
<< m1 >>
rect 44 257 45 258 
<< m1 >>
rect 55 257 56 258 
<< m1 >>
rect 64 257 65 258 
<< m1 >>
rect 118 257 119 258 
<< m2 >>
rect 118 257 119 258 
<< m2c >>
rect 118 257 119 258 
<< m1 >>
rect 118 257 119 258 
<< m2 >>
rect 118 257 119 258 
<< m1 >>
rect 148 257 149 258 
<< m1 >>
rect 163 257 164 258 
<< m2 >>
rect 163 257 164 258 
<< m2c >>
rect 163 257 164 258 
<< m1 >>
rect 163 257 164 258 
<< m2 >>
rect 163 257 164 258 
<< m2 >>
rect 171 257 172 258 
<< m1 >>
rect 172 257 173 258 
<< m1 >>
rect 177 257 178 258 
<< m2 >>
rect 177 257 178 258 
<< m2c >>
rect 177 257 178 258 
<< m1 >>
rect 177 257 178 258 
<< m2 >>
rect 177 257 178 258 
<< m1 >>
rect 181 257 182 258 
<< m1 >>
rect 186 257 187 258 
<< m2 >>
rect 186 257 187 258 
<< m2c >>
rect 186 257 187 258 
<< m1 >>
rect 186 257 187 258 
<< m2 >>
rect 186 257 187 258 
<< m1 >>
rect 190 257 191 258 
<< m2 >>
rect 190 257 191 258 
<< m2c >>
rect 190 257 191 258 
<< m1 >>
rect 190 257 191 258 
<< m2 >>
rect 190 257 191 258 
<< m1 >>
rect 207 257 208 258 
<< m2 >>
rect 207 257 208 258 
<< m2c >>
rect 207 257 208 258 
<< m1 >>
rect 207 257 208 258 
<< m2 >>
rect 207 257 208 258 
<< m1 >>
rect 211 257 212 258 
<< m2 >>
rect 211 257 212 258 
<< m2c >>
rect 211 257 212 258 
<< m1 >>
rect 211 257 212 258 
<< m2 >>
rect 211 257 212 258 
<< m1 >>
rect 219 257 220 258 
<< m2 >>
rect 219 257 220 258 
<< m2c >>
rect 219 257 220 258 
<< m1 >>
rect 219 257 220 258 
<< m2 >>
rect 219 257 220 258 
<< m1 >>
rect 220 257 221 258 
<< m1 >>
rect 221 257 222 258 
<< m1 >>
rect 222 257 223 258 
<< m1 >>
rect 223 257 224 258 
<< m1 >>
rect 224 257 225 258 
<< m1 >>
rect 225 257 226 258 
<< m1 >>
rect 226 257 227 258 
<< m1 >>
rect 227 257 228 258 
<< m1 >>
rect 228 257 229 258 
<< m2 >>
rect 228 257 229 258 
<< m1 >>
rect 229 257 230 258 
<< m1 >>
rect 230 257 231 258 
<< m1 >>
rect 231 257 232 258 
<< m1 >>
rect 232 257 233 258 
<< m1 >>
rect 235 257 236 258 
<< m1 >>
rect 237 257 238 258 
<< m1 >>
rect 247 257 248 258 
<< m1 >>
rect 248 257 249 258 
<< m1 >>
rect 249 257 250 258 
<< m1 >>
rect 250 257 251 258 
<< m1 >>
rect 251 257 252 258 
<< m1 >>
rect 252 257 253 258 
<< m1 >>
rect 253 257 254 258 
<< m2 >>
rect 253 257 254 258 
<< m2c >>
rect 253 257 254 258 
<< m1 >>
rect 253 257 254 258 
<< m2 >>
rect 253 257 254 258 
<< m1 >>
rect 255 257 256 258 
<< m2 >>
rect 255 257 256 258 
<< m2c >>
rect 255 257 256 258 
<< m1 >>
rect 255 257 256 258 
<< m2 >>
rect 255 257 256 258 
<< m1 >>
rect 259 257 260 258 
<< m2 >>
rect 259 257 260 258 
<< m2c >>
rect 259 257 260 258 
<< m1 >>
rect 259 257 260 258 
<< m2 >>
rect 259 257 260 258 
<< m1 >>
rect 262 257 263 258 
<< m2 >>
rect 262 257 263 258 
<< m1 >>
rect 263 257 264 258 
<< m1 >>
rect 264 257 265 258 
<< m2 >>
rect 264 257 265 258 
<< m1 >>
rect 265 257 266 258 
<< m1 >>
rect 266 257 267 258 
<< m1 >>
rect 267 257 268 258 
<< m1 >>
rect 268 257 269 258 
<< m1 >>
rect 269 257 270 258 
<< m1 >>
rect 270 257 271 258 
<< m1 >>
rect 271 257 272 258 
<< m1 >>
rect 272 257 273 258 
<< m1 >>
rect 273 257 274 258 
<< m1 >>
rect 274 257 275 258 
<< m1 >>
rect 275 257 276 258 
<< m1 >>
rect 276 257 277 258 
<< m1 >>
rect 277 257 278 258 
<< m1 >>
rect 278 257 279 258 
<< m2 >>
rect 278 257 279 258 
<< m2c >>
rect 278 257 279 258 
<< m1 >>
rect 278 257 279 258 
<< m2 >>
rect 278 257 279 258 
<< m2 >>
rect 279 257 280 258 
<< m1 >>
rect 280 257 281 258 
<< m2 >>
rect 280 257 281 258 
<< m2 >>
rect 281 257 282 258 
<< m2 >>
rect 282 257 283 258 
<< m2 >>
rect 283 257 284 258 
<< m2 >>
rect 284 257 285 258 
<< m2 >>
rect 285 257 286 258 
<< m2 >>
rect 286 257 287 258 
<< m2 >>
rect 287 257 288 258 
<< m2 >>
rect 288 257 289 258 
<< m2 >>
rect 289 257 290 258 
<< m2 >>
rect 290 257 291 258 
<< m2 >>
rect 291 257 292 258 
<< m2 >>
rect 292 257 293 258 
<< m2 >>
rect 293 257 294 258 
<< m2 >>
rect 294 257 295 258 
<< m2 >>
rect 295 257 296 258 
<< m2 >>
rect 296 257 297 258 
<< m2 >>
rect 297 257 298 258 
<< m2 >>
rect 298 257 299 258 
<< m2 >>
rect 299 257 300 258 
<< m2 >>
rect 300 257 301 258 
<< m2 >>
rect 301 257 302 258 
<< m2 >>
rect 302 257 303 258 
<< m2 >>
rect 303 257 304 258 
<< m1 >>
rect 307 257 308 258 
<< m2 >>
rect 318 257 319 258 
<< m2 >>
rect 319 257 320 258 
<< m2 >>
rect 320 257 321 258 
<< m2 >>
rect 321 257 322 258 
<< m2 >>
rect 322 257 323 258 
<< m2 >>
rect 323 257 324 258 
<< m2 >>
rect 324 257 325 258 
<< m2 >>
rect 325 257 326 258 
<< m2 >>
rect 326 257 327 258 
<< m2 >>
rect 327 257 328 258 
<< m2 >>
rect 328 257 329 258 
<< m2 >>
rect 329 257 330 258 
<< m2 >>
rect 330 257 331 258 
<< m2 >>
rect 331 257 332 258 
<< m2 >>
rect 332 257 333 258 
<< m2 >>
rect 333 257 334 258 
<< m2 >>
rect 334 257 335 258 
<< m2 >>
rect 335 257 336 258 
<< m1 >>
rect 342 257 343 258 
<< m2 >>
rect 342 257 343 258 
<< m2c >>
rect 342 257 343 258 
<< m1 >>
rect 342 257 343 258 
<< m2 >>
rect 342 257 343 258 
<< m1 >>
rect 346 257 347 258 
<< m2 >>
rect 346 257 347 258 
<< m2c >>
rect 346 257 347 258 
<< m1 >>
rect 346 257 347 258 
<< m2 >>
rect 346 257 347 258 
<< m1 >>
rect 352 257 353 258 
<< m1 >>
rect 353 257 354 258 
<< m1 >>
rect 354 257 355 258 
<< m1 >>
rect 355 257 356 258 
<< m1 >>
rect 356 257 357 258 
<< m1 >>
rect 357 257 358 258 
<< m1 >>
rect 358 257 359 258 
<< m1 >>
rect 359 257 360 258 
<< m1 >>
rect 360 257 361 258 
<< m1 >>
rect 361 257 362 258 
<< m1 >>
rect 362 257 363 258 
<< m1 >>
rect 363 257 364 258 
<< m1 >>
rect 364 257 365 258 
<< m1 >>
rect 365 257 366 258 
<< m1 >>
rect 366 257 367 258 
<< m2 >>
rect 366 257 367 258 
<< m2c >>
rect 366 257 367 258 
<< m1 >>
rect 366 257 367 258 
<< m2 >>
rect 366 257 367 258 
<< m1 >>
rect 376 257 377 258 
<< m2 >>
rect 376 257 377 258 
<< m2c >>
rect 376 257 377 258 
<< m1 >>
rect 376 257 377 258 
<< m2 >>
rect 376 257 377 258 
<< m2 >>
rect 378 257 379 258 
<< m2 >>
rect 379 257 380 258 
<< m2 >>
rect 380 257 381 258 
<< m2 >>
rect 381 257 382 258 
<< m2 >>
rect 382 257 383 258 
<< m2 >>
rect 383 257 384 258 
<< m2 >>
rect 384 257 385 258 
<< m2 >>
rect 385 257 386 258 
<< m2 >>
rect 386 257 387 258 
<< m2 >>
rect 387 257 388 258 
<< m2 >>
rect 388 257 389 258 
<< m2 >>
rect 389 257 390 258 
<< m2 >>
rect 390 257 391 258 
<< m2 >>
rect 391 257 392 258 
<< m2 >>
rect 392 257 393 258 
<< m2 >>
rect 412 257 413 258 
<< m2 >>
rect 415 257 416 258 
<< m1 >>
rect 416 257 417 258 
<< m2 >>
rect 416 257 417 258 
<< m2 >>
rect 417 257 418 258 
<< m2 >>
rect 418 257 419 258 
<< m1 >>
rect 419 257 420 258 
<< m2 >>
rect 419 257 420 258 
<< m2 >>
rect 420 257 421 258 
<< m2 >>
rect 421 257 422 258 
<< m2 >>
rect 422 257 423 258 
<< m2 >>
rect 423 257 424 258 
<< m2 >>
rect 424 257 425 258 
<< m2 >>
rect 425 257 426 258 
<< m2 >>
rect 426 257 427 258 
<< m2 >>
rect 427 257 428 258 
<< m2 >>
rect 428 257 429 258 
<< m1 >>
rect 430 257 431 258 
<< m2 >>
rect 431 257 432 258 
<< m1 >>
rect 437 257 438 258 
<< m1 >>
rect 442 257 443 258 
<< m1 >>
rect 484 257 485 258 
<< m1 >>
rect 523 257 524 258 
<< m1 >>
rect 19 258 20 259 
<< m1 >>
rect 22 258 23 259 
<< m1 >>
rect 44 258 45 259 
<< m1 >>
rect 55 258 56 259 
<< m1 >>
rect 64 258 65 259 
<< m2 >>
rect 92 258 93 259 
<< m2 >>
rect 93 258 94 259 
<< m2 >>
rect 94 258 95 259 
<< m2 >>
rect 95 258 96 259 
<< m2 >>
rect 96 258 97 259 
<< m2 >>
rect 97 258 98 259 
<< m2 >>
rect 98 258 99 259 
<< m2 >>
rect 99 258 100 259 
<< m2 >>
rect 100 258 101 259 
<< m2 >>
rect 101 258 102 259 
<< m2 >>
rect 102 258 103 259 
<< m2 >>
rect 103 258 104 259 
<< m2 >>
rect 104 258 105 259 
<< m2 >>
rect 105 258 106 259 
<< m2 >>
rect 106 258 107 259 
<< m2 >>
rect 107 258 108 259 
<< m2 >>
rect 108 258 109 259 
<< m2 >>
rect 109 258 110 259 
<< m2 >>
rect 110 258 111 259 
<< m2 >>
rect 111 258 112 259 
<< m2 >>
rect 112 258 113 259 
<< m2 >>
rect 113 258 114 259 
<< m2 >>
rect 114 258 115 259 
<< m2 >>
rect 115 258 116 259 
<< m2 >>
rect 116 258 117 259 
<< m2 >>
rect 117 258 118 259 
<< m2 >>
rect 118 258 119 259 
<< m1 >>
rect 148 258 149 259 
<< m2 >>
rect 163 258 164 259 
<< m2 >>
rect 171 258 172 259 
<< m1 >>
rect 172 258 173 259 
<< m2 >>
rect 177 258 178 259 
<< m1 >>
rect 181 258 182 259 
<< m2 >>
rect 186 258 187 259 
<< m2 >>
rect 190 258 191 259 
<< m2 >>
rect 192 258 193 259 
<< m2 >>
rect 193 258 194 259 
<< m2 >>
rect 194 258 195 259 
<< m2 >>
rect 195 258 196 259 
<< m2 >>
rect 196 258 197 259 
<< m2 >>
rect 197 258 198 259 
<< m2 >>
rect 198 258 199 259 
<< m2 >>
rect 199 258 200 259 
<< m2 >>
rect 200 258 201 259 
<< m2 >>
rect 201 258 202 259 
<< m2 >>
rect 202 258 203 259 
<< m2 >>
rect 203 258 204 259 
<< m2 >>
rect 204 258 205 259 
<< m2 >>
rect 205 258 206 259 
<< m2 >>
rect 206 258 207 259 
<< m2 >>
rect 207 258 208 259 
<< m2 >>
rect 211 258 212 259 
<< m2 >>
rect 212 258 213 259 
<< m2 >>
rect 213 258 214 259 
<< m2 >>
rect 214 258 215 259 
<< m2 >>
rect 215 258 216 259 
<< m2 >>
rect 216 258 217 259 
<< m2 >>
rect 217 258 218 259 
<< m2 >>
rect 219 258 220 259 
<< m2 >>
rect 228 258 229 259 
<< m1 >>
rect 235 258 236 259 
<< m1 >>
rect 237 258 238 259 
<< m2 >>
rect 253 258 254 259 
<< m2 >>
rect 255 258 256 259 
<< m2 >>
rect 259 258 260 259 
<< m2 >>
rect 262 258 263 259 
<< m2 >>
rect 264 258 265 259 
<< m1 >>
rect 280 258 281 259 
<< m2 >>
rect 303 258 304 259 
<< m1 >>
rect 307 258 308 259 
<< m2 >>
rect 335 258 336 259 
<< m2 >>
rect 342 258 343 259 
<< m2 >>
rect 346 258 347 259 
<< m2 >>
rect 366 258 367 259 
<< m2 >>
rect 372 258 373 259 
<< m2 >>
rect 373 258 374 259 
<< m2 >>
rect 374 258 375 259 
<< m2 >>
rect 375 258 376 259 
<< m2 >>
rect 376 258 377 259 
<< m1 >>
rect 378 258 379 259 
<< m2 >>
rect 378 258 379 259 
<< m2c >>
rect 378 258 379 259 
<< m1 >>
rect 378 258 379 259 
<< m2 >>
rect 378 258 379 259 
<< m1 >>
rect 386 258 387 259 
<< m1 >>
rect 387 258 388 259 
<< m1 >>
rect 388 258 389 259 
<< m1 >>
rect 389 258 390 259 
<< m1 >>
rect 390 258 391 259 
<< m1 >>
rect 391 258 392 259 
<< m1 >>
rect 392 258 393 259 
<< m1 >>
rect 393 258 394 259 
<< m1 >>
rect 394 258 395 259 
<< m1 >>
rect 395 258 396 259 
<< m2 >>
rect 395 258 396 259 
<< m2c >>
rect 395 258 396 259 
<< m1 >>
rect 395 258 396 259 
<< m2 >>
rect 395 258 396 259 
<< m2 >>
rect 396 258 397 259 
<< m2 >>
rect 397 258 398 259 
<< m2 >>
rect 398 258 399 259 
<< m2 >>
rect 399 258 400 259 
<< m2 >>
rect 400 258 401 259 
<< m2 >>
rect 401 258 402 259 
<< m2 >>
rect 402 258 403 259 
<< m2 >>
rect 403 258 404 259 
<< m2 >>
rect 404 258 405 259 
<< m2 >>
rect 405 258 406 259 
<< m2 >>
rect 406 258 407 259 
<< m2 >>
rect 407 258 408 259 
<< m2 >>
rect 408 258 409 259 
<< m2 >>
rect 409 258 410 259 
<< m2 >>
rect 410 258 411 259 
<< m2 >>
rect 411 258 412 259 
<< m2 >>
rect 412 258 413 259 
<< m2 >>
rect 415 258 416 259 
<< m1 >>
rect 416 258 417 259 
<< m1 >>
rect 419 258 420 259 
<< m1 >>
rect 430 258 431 259 
<< m2 >>
rect 431 258 432 259 
<< m1 >>
rect 437 258 438 259 
<< m1 >>
rect 442 258 443 259 
<< m1 >>
rect 484 258 485 259 
<< m1 >>
rect 523 258 524 259 
<< m1 >>
rect 19 259 20 260 
<< m1 >>
rect 22 259 23 260 
<< m1 >>
rect 44 259 45 260 
<< m1 >>
rect 55 259 56 260 
<< m1 >>
rect 64 259 65 260 
<< m1 >>
rect 91 259 92 260 
<< m1 >>
rect 92 259 93 260 
<< m2 >>
rect 92 259 93 260 
<< m1 >>
rect 93 259 94 260 
<< m1 >>
rect 94 259 95 260 
<< m1 >>
rect 95 259 96 260 
<< m1 >>
rect 96 259 97 260 
<< m1 >>
rect 97 259 98 260 
<< m1 >>
rect 98 259 99 260 
<< m1 >>
rect 99 259 100 260 
<< m1 >>
rect 100 259 101 260 
<< m1 >>
rect 101 259 102 260 
<< m1 >>
rect 102 259 103 260 
<< m1 >>
rect 103 259 104 260 
<< m1 >>
rect 104 259 105 260 
<< m1 >>
rect 105 259 106 260 
<< m1 >>
rect 106 259 107 260 
<< m1 >>
rect 107 259 108 260 
<< m1 >>
rect 108 259 109 260 
<< m1 >>
rect 109 259 110 260 
<< m1 >>
rect 110 259 111 260 
<< m1 >>
rect 111 259 112 260 
<< m1 >>
rect 112 259 113 260 
<< m1 >>
rect 113 259 114 260 
<< m1 >>
rect 114 259 115 260 
<< m1 >>
rect 115 259 116 260 
<< m1 >>
rect 116 259 117 260 
<< m1 >>
rect 117 259 118 260 
<< m1 >>
rect 118 259 119 260 
<< m2 >>
rect 118 259 119 260 
<< m1 >>
rect 119 259 120 260 
<< m2 >>
rect 119 259 120 260 
<< m1 >>
rect 120 259 121 260 
<< m2 >>
rect 120 259 121 260 
<< m1 >>
rect 121 259 122 260 
<< m2 >>
rect 121 259 122 260 
<< m1 >>
rect 122 259 123 260 
<< m2 >>
rect 122 259 123 260 
<< m1 >>
rect 123 259 124 260 
<< m2 >>
rect 123 259 124 260 
<< m1 >>
rect 124 259 125 260 
<< m2 >>
rect 124 259 125 260 
<< m1 >>
rect 125 259 126 260 
<< m2 >>
rect 125 259 126 260 
<< m1 >>
rect 126 259 127 260 
<< m2 >>
rect 126 259 127 260 
<< m1 >>
rect 127 259 128 260 
<< m2 >>
rect 127 259 128 260 
<< m1 >>
rect 128 259 129 260 
<< m2 >>
rect 128 259 129 260 
<< m1 >>
rect 129 259 130 260 
<< m2 >>
rect 129 259 130 260 
<< m1 >>
rect 130 259 131 260 
<< m2 >>
rect 130 259 131 260 
<< m1 >>
rect 131 259 132 260 
<< m2 >>
rect 131 259 132 260 
<< m1 >>
rect 132 259 133 260 
<< m2 >>
rect 132 259 133 260 
<< m1 >>
rect 133 259 134 260 
<< m2 >>
rect 133 259 134 260 
<< m1 >>
rect 134 259 135 260 
<< m2 >>
rect 134 259 135 260 
<< m1 >>
rect 135 259 136 260 
<< m2 >>
rect 135 259 136 260 
<< m1 >>
rect 136 259 137 260 
<< m2 >>
rect 136 259 137 260 
<< m1 >>
rect 137 259 138 260 
<< m2 >>
rect 137 259 138 260 
<< m1 >>
rect 138 259 139 260 
<< m2 >>
rect 138 259 139 260 
<< m1 >>
rect 139 259 140 260 
<< m2 >>
rect 139 259 140 260 
<< m1 >>
rect 140 259 141 260 
<< m2 >>
rect 140 259 141 260 
<< m1 >>
rect 141 259 142 260 
<< m2 >>
rect 141 259 142 260 
<< m1 >>
rect 142 259 143 260 
<< m2 >>
rect 142 259 143 260 
<< m2 >>
rect 143 259 144 260 
<< m1 >>
rect 144 259 145 260 
<< m2 >>
rect 144 259 145 260 
<< m2c >>
rect 144 259 145 260 
<< m1 >>
rect 144 259 145 260 
<< m2 >>
rect 144 259 145 260 
<< m1 >>
rect 145 259 146 260 
<< m1 >>
rect 146 259 147 260 
<< m2 >>
rect 146 259 147 260 
<< m2c >>
rect 146 259 147 260 
<< m1 >>
rect 146 259 147 260 
<< m2 >>
rect 146 259 147 260 
<< m2 >>
rect 147 259 148 260 
<< m1 >>
rect 148 259 149 260 
<< m2 >>
rect 148 259 149 260 
<< m2 >>
rect 149 259 150 260 
<< m1 >>
rect 150 259 151 260 
<< m2 >>
rect 150 259 151 260 
<< m1 >>
rect 151 259 152 260 
<< m2 >>
rect 151 259 152 260 
<< m1 >>
rect 152 259 153 260 
<< m2 >>
rect 152 259 153 260 
<< m1 >>
rect 153 259 154 260 
<< m2 >>
rect 153 259 154 260 
<< m1 >>
rect 154 259 155 260 
<< m2 >>
rect 154 259 155 260 
<< m1 >>
rect 155 259 156 260 
<< m2 >>
rect 155 259 156 260 
<< m1 >>
rect 156 259 157 260 
<< m2 >>
rect 156 259 157 260 
<< m1 >>
rect 157 259 158 260 
<< m2 >>
rect 157 259 158 260 
<< m1 >>
rect 158 259 159 260 
<< m2 >>
rect 158 259 159 260 
<< m1 >>
rect 159 259 160 260 
<< m1 >>
rect 160 259 161 260 
<< m1 >>
rect 161 259 162 260 
<< m1 >>
rect 162 259 163 260 
<< m1 >>
rect 163 259 164 260 
<< m2 >>
rect 163 259 164 260 
<< m1 >>
rect 164 259 165 260 
<< m1 >>
rect 165 259 166 260 
<< m1 >>
rect 166 259 167 260 
<< m1 >>
rect 167 259 168 260 
<< m1 >>
rect 168 259 169 260 
<< m1 >>
rect 169 259 170 260 
<< m1 >>
rect 170 259 171 260 
<< m2 >>
rect 170 259 171 260 
<< m2c >>
rect 170 259 171 260 
<< m1 >>
rect 170 259 171 260 
<< m2 >>
rect 170 259 171 260 
<< m2 >>
rect 171 259 172 260 
<< m1 >>
rect 172 259 173 260 
<< m1 >>
rect 173 259 174 260 
<< m1 >>
rect 174 259 175 260 
<< m1 >>
rect 175 259 176 260 
<< m1 >>
rect 176 259 177 260 
<< m1 >>
rect 177 259 178 260 
<< m2 >>
rect 177 259 178 260 
<< m1 >>
rect 178 259 179 260 
<< m1 >>
rect 179 259 180 260 
<< m2 >>
rect 179 259 180 260 
<< m2c >>
rect 179 259 180 260 
<< m1 >>
rect 179 259 180 260 
<< m2 >>
rect 179 259 180 260 
<< m2 >>
rect 180 259 181 260 
<< m1 >>
rect 181 259 182 260 
<< m2 >>
rect 181 259 182 260 
<< m2 >>
rect 182 259 183 260 
<< m1 >>
rect 183 259 184 260 
<< m2 >>
rect 183 259 184 260 
<< m2c >>
rect 183 259 184 260 
<< m1 >>
rect 183 259 184 260 
<< m2 >>
rect 183 259 184 260 
<< m1 >>
rect 184 259 185 260 
<< m1 >>
rect 185 259 186 260 
<< m1 >>
rect 186 259 187 260 
<< m2 >>
rect 186 259 187 260 
<< m1 >>
rect 187 259 188 260 
<< m1 >>
rect 188 259 189 260 
<< m1 >>
rect 189 259 190 260 
<< m1 >>
rect 190 259 191 260 
<< m2 >>
rect 190 259 191 260 
<< m1 >>
rect 191 259 192 260 
<< m1 >>
rect 192 259 193 260 
<< m2 >>
rect 192 259 193 260 
<< m1 >>
rect 193 259 194 260 
<< m1 >>
rect 194 259 195 260 
<< m1 >>
rect 195 259 196 260 
<< m1 >>
rect 196 259 197 260 
<< m1 >>
rect 197 259 198 260 
<< m1 >>
rect 198 259 199 260 
<< m1 >>
rect 199 259 200 260 
<< m1 >>
rect 200 259 201 260 
<< m1 >>
rect 201 259 202 260 
<< m1 >>
rect 202 259 203 260 
<< m1 >>
rect 203 259 204 260 
<< m1 >>
rect 204 259 205 260 
<< m1 >>
rect 205 259 206 260 
<< m1 >>
rect 206 259 207 260 
<< m1 >>
rect 207 259 208 260 
<< m1 >>
rect 208 259 209 260 
<< m1 >>
rect 209 259 210 260 
<< m1 >>
rect 210 259 211 260 
<< m1 >>
rect 211 259 212 260 
<< m1 >>
rect 212 259 213 260 
<< m1 >>
rect 213 259 214 260 
<< m1 >>
rect 214 259 215 260 
<< m1 >>
rect 215 259 216 260 
<< m1 >>
rect 216 259 217 260 
<< m1 >>
rect 217 259 218 260 
<< m2 >>
rect 217 259 218 260 
<< m1 >>
rect 218 259 219 260 
<< m1 >>
rect 219 259 220 260 
<< m2 >>
rect 219 259 220 260 
<< m1 >>
rect 220 259 221 260 
<< m1 >>
rect 221 259 222 260 
<< m1 >>
rect 222 259 223 260 
<< m1 >>
rect 223 259 224 260 
<< m1 >>
rect 224 259 225 260 
<< m1 >>
rect 225 259 226 260 
<< m1 >>
rect 226 259 227 260 
<< m1 >>
rect 227 259 228 260 
<< m1 >>
rect 228 259 229 260 
<< m2 >>
rect 228 259 229 260 
<< m1 >>
rect 229 259 230 260 
<< m2 >>
rect 229 259 230 260 
<< m1 >>
rect 230 259 231 260 
<< m2 >>
rect 230 259 231 260 
<< m1 >>
rect 231 259 232 260 
<< m2 >>
rect 231 259 232 260 
<< m1 >>
rect 232 259 233 260 
<< m1 >>
rect 233 259 234 260 
<< m2 >>
rect 233 259 234 260 
<< m2c >>
rect 233 259 234 260 
<< m1 >>
rect 233 259 234 260 
<< m2 >>
rect 233 259 234 260 
<< m2 >>
rect 234 259 235 260 
<< m1 >>
rect 235 259 236 260 
<< m2 >>
rect 235 259 236 260 
<< m2 >>
rect 236 259 237 260 
<< m1 >>
rect 237 259 238 260 
<< m2 >>
rect 237 259 238 260 
<< m2 >>
rect 238 259 239 260 
<< m1 >>
rect 239 259 240 260 
<< m2 >>
rect 239 259 240 260 
<< m2c >>
rect 239 259 240 260 
<< m1 >>
rect 239 259 240 260 
<< m2 >>
rect 239 259 240 260 
<< m1 >>
rect 240 259 241 260 
<< m1 >>
rect 241 259 242 260 
<< m1 >>
rect 242 259 243 260 
<< m1 >>
rect 243 259 244 260 
<< m1 >>
rect 244 259 245 260 
<< m1 >>
rect 245 259 246 260 
<< m1 >>
rect 246 259 247 260 
<< m1 >>
rect 247 259 248 260 
<< m1 >>
rect 248 259 249 260 
<< m1 >>
rect 249 259 250 260 
<< m1 >>
rect 250 259 251 260 
<< m1 >>
rect 251 259 252 260 
<< m1 >>
rect 252 259 253 260 
<< m1 >>
rect 253 259 254 260 
<< m2 >>
rect 253 259 254 260 
<< m1 >>
rect 254 259 255 260 
<< m1 >>
rect 255 259 256 260 
<< m2 >>
rect 255 259 256 260 
<< m1 >>
rect 256 259 257 260 
<< m1 >>
rect 257 259 258 260 
<< m1 >>
rect 258 259 259 260 
<< m1 >>
rect 259 259 260 260 
<< m2 >>
rect 259 259 260 260 
<< m1 >>
rect 260 259 261 260 
<< m1 >>
rect 261 259 262 260 
<< m1 >>
rect 262 259 263 260 
<< m2 >>
rect 262 259 263 260 
<< m1 >>
rect 263 259 264 260 
<< m1 >>
rect 264 259 265 260 
<< m2 >>
rect 264 259 265 260 
<< m1 >>
rect 265 259 266 260 
<< m1 >>
rect 266 259 267 260 
<< m1 >>
rect 267 259 268 260 
<< m1 >>
rect 268 259 269 260 
<< m1 >>
rect 269 259 270 260 
<< m1 >>
rect 270 259 271 260 
<< m1 >>
rect 271 259 272 260 
<< m1 >>
rect 272 259 273 260 
<< m1 >>
rect 273 259 274 260 
<< m1 >>
rect 274 259 275 260 
<< m1 >>
rect 275 259 276 260 
<< m1 >>
rect 276 259 277 260 
<< m1 >>
rect 277 259 278 260 
<< m1 >>
rect 278 259 279 260 
<< m2 >>
rect 278 259 279 260 
<< m2c >>
rect 278 259 279 260 
<< m1 >>
rect 278 259 279 260 
<< m2 >>
rect 278 259 279 260 
<< m2 >>
rect 279 259 280 260 
<< m1 >>
rect 280 259 281 260 
<< m2 >>
rect 280 259 281 260 
<< m2 >>
rect 281 259 282 260 
<< m1 >>
rect 282 259 283 260 
<< m2 >>
rect 282 259 283 260 
<< m2c >>
rect 282 259 283 260 
<< m1 >>
rect 282 259 283 260 
<< m2 >>
rect 282 259 283 260 
<< m1 >>
rect 283 259 284 260 
<< m1 >>
rect 284 259 285 260 
<< m1 >>
rect 285 259 286 260 
<< m1 >>
rect 286 259 287 260 
<< m1 >>
rect 287 259 288 260 
<< m1 >>
rect 288 259 289 260 
<< m1 >>
rect 289 259 290 260 
<< m1 >>
rect 290 259 291 260 
<< m1 >>
rect 291 259 292 260 
<< m1 >>
rect 292 259 293 260 
<< m1 >>
rect 293 259 294 260 
<< m1 >>
rect 294 259 295 260 
<< m1 >>
rect 295 259 296 260 
<< m1 >>
rect 296 259 297 260 
<< m1 >>
rect 297 259 298 260 
<< m1 >>
rect 298 259 299 260 
<< m1 >>
rect 299 259 300 260 
<< m1 >>
rect 300 259 301 260 
<< m1 >>
rect 301 259 302 260 
<< m1 >>
rect 302 259 303 260 
<< m1 >>
rect 303 259 304 260 
<< m2 >>
rect 303 259 304 260 
<< m1 >>
rect 304 259 305 260 
<< m1 >>
rect 305 259 306 260 
<< m2 >>
rect 305 259 306 260 
<< m2c >>
rect 305 259 306 260 
<< m1 >>
rect 305 259 306 260 
<< m2 >>
rect 305 259 306 260 
<< m2 >>
rect 306 259 307 260 
<< m1 >>
rect 307 259 308 260 
<< m2 >>
rect 307 259 308 260 
<< m2 >>
rect 308 259 309 260 
<< m1 >>
rect 309 259 310 260 
<< m2 >>
rect 309 259 310 260 
<< m1 >>
rect 310 259 311 260 
<< m2 >>
rect 310 259 311 260 
<< m1 >>
rect 311 259 312 260 
<< m2 >>
rect 311 259 312 260 
<< m1 >>
rect 312 259 313 260 
<< m2 >>
rect 312 259 313 260 
<< m1 >>
rect 313 259 314 260 
<< m2 >>
rect 313 259 314 260 
<< m1 >>
rect 314 259 315 260 
<< m2 >>
rect 314 259 315 260 
<< m1 >>
rect 315 259 316 260 
<< m2 >>
rect 315 259 316 260 
<< m1 >>
rect 316 259 317 260 
<< m2 >>
rect 316 259 317 260 
<< m1 >>
rect 317 259 318 260 
<< m2 >>
rect 317 259 318 260 
<< m1 >>
rect 318 259 319 260 
<< m2 >>
rect 318 259 319 260 
<< m1 >>
rect 319 259 320 260 
<< m2 >>
rect 319 259 320 260 
<< m1 >>
rect 320 259 321 260 
<< m2 >>
rect 320 259 321 260 
<< m1 >>
rect 321 259 322 260 
<< m2 >>
rect 321 259 322 260 
<< m1 >>
rect 322 259 323 260 
<< m2 >>
rect 322 259 323 260 
<< m1 >>
rect 323 259 324 260 
<< m1 >>
rect 324 259 325 260 
<< m1 >>
rect 325 259 326 260 
<< m1 >>
rect 326 259 327 260 
<< m1 >>
rect 327 259 328 260 
<< m1 >>
rect 328 259 329 260 
<< m1 >>
rect 329 259 330 260 
<< m1 >>
rect 330 259 331 260 
<< m1 >>
rect 331 259 332 260 
<< m1 >>
rect 332 259 333 260 
<< m1 >>
rect 333 259 334 260 
<< m1 >>
rect 334 259 335 260 
<< m1 >>
rect 335 259 336 260 
<< m2 >>
rect 335 259 336 260 
<< m1 >>
rect 336 259 337 260 
<< m2 >>
rect 336 259 337 260 
<< m1 >>
rect 337 259 338 260 
<< m2 >>
rect 337 259 338 260 
<< m1 >>
rect 338 259 339 260 
<< m2 >>
rect 338 259 339 260 
<< m1 >>
rect 339 259 340 260 
<< m2 >>
rect 339 259 340 260 
<< m1 >>
rect 340 259 341 260 
<< m2 >>
rect 340 259 341 260 
<< m1 >>
rect 341 259 342 260 
<< m1 >>
rect 342 259 343 260 
<< m2 >>
rect 342 259 343 260 
<< m1 >>
rect 343 259 344 260 
<< m1 >>
rect 344 259 345 260 
<< m1 >>
rect 345 259 346 260 
<< m1 >>
rect 346 259 347 260 
<< m2 >>
rect 346 259 347 260 
<< m1 >>
rect 347 259 348 260 
<< m1 >>
rect 348 259 349 260 
<< m1 >>
rect 349 259 350 260 
<< m1 >>
rect 350 259 351 260 
<< m1 >>
rect 351 259 352 260 
<< m1 >>
rect 352 259 353 260 
<< m1 >>
rect 353 259 354 260 
<< m1 >>
rect 354 259 355 260 
<< m1 >>
rect 355 259 356 260 
<< m1 >>
rect 356 259 357 260 
<< m1 >>
rect 357 259 358 260 
<< m1 >>
rect 358 259 359 260 
<< m1 >>
rect 359 259 360 260 
<< m1 >>
rect 360 259 361 260 
<< m1 >>
rect 361 259 362 260 
<< m1 >>
rect 362 259 363 260 
<< m1 >>
rect 363 259 364 260 
<< m1 >>
rect 364 259 365 260 
<< m1 >>
rect 365 259 366 260 
<< m1 >>
rect 366 259 367 260 
<< m2 >>
rect 366 259 367 260 
<< m1 >>
rect 367 259 368 260 
<< m1 >>
rect 368 259 369 260 
<< m1 >>
rect 369 259 370 260 
<< m1 >>
rect 370 259 371 260 
<< m1 >>
rect 371 259 372 260 
<< m1 >>
rect 372 259 373 260 
<< m2 >>
rect 372 259 373 260 
<< m1 >>
rect 373 259 374 260 
<< m1 >>
rect 374 259 375 260 
<< m1 >>
rect 375 259 376 260 
<< m1 >>
rect 376 259 377 260 
<< m1 >>
rect 377 259 378 260 
<< m1 >>
rect 378 259 379 260 
<< m1 >>
rect 386 259 387 260 
<< m1 >>
rect 397 259 398 260 
<< m1 >>
rect 398 259 399 260 
<< m1 >>
rect 399 259 400 260 
<< m1 >>
rect 400 259 401 260 
<< m1 >>
rect 401 259 402 260 
<< m1 >>
rect 402 259 403 260 
<< m1 >>
rect 403 259 404 260 
<< m1 >>
rect 404 259 405 260 
<< m1 >>
rect 405 259 406 260 
<< m1 >>
rect 406 259 407 260 
<< m1 >>
rect 407 259 408 260 
<< m1 >>
rect 408 259 409 260 
<< m1 >>
rect 409 259 410 260 
<< m1 >>
rect 410 259 411 260 
<< m1 >>
rect 411 259 412 260 
<< m1 >>
rect 412 259 413 260 
<< m1 >>
rect 413 259 414 260 
<< m1 >>
rect 414 259 415 260 
<< m2 >>
rect 414 259 415 260 
<< m2c >>
rect 414 259 415 260 
<< m1 >>
rect 414 259 415 260 
<< m2 >>
rect 414 259 415 260 
<< m2 >>
rect 415 259 416 260 
<< m1 >>
rect 416 259 417 260 
<< m1 >>
rect 419 259 420 260 
<< m2 >>
rect 420 259 421 260 
<< m1 >>
rect 421 259 422 260 
<< m2 >>
rect 421 259 422 260 
<< m2c >>
rect 421 259 422 260 
<< m1 >>
rect 421 259 422 260 
<< m2 >>
rect 421 259 422 260 
<< m1 >>
rect 422 259 423 260 
<< m1 >>
rect 423 259 424 260 
<< m1 >>
rect 424 259 425 260 
<< m1 >>
rect 425 259 426 260 
<< m1 >>
rect 426 259 427 260 
<< m1 >>
rect 427 259 428 260 
<< m1 >>
rect 428 259 429 260 
<< m2 >>
rect 428 259 429 260 
<< m2c >>
rect 428 259 429 260 
<< m1 >>
rect 428 259 429 260 
<< m2 >>
rect 428 259 429 260 
<< m2 >>
rect 429 259 430 260 
<< m1 >>
rect 430 259 431 260 
<< m2 >>
rect 430 259 431 260 
<< m2 >>
rect 431 259 432 260 
<< m1 >>
rect 437 259 438 260 
<< m1 >>
rect 442 259 443 260 
<< m1 >>
rect 484 259 485 260 
<< m1 >>
rect 523 259 524 260 
<< m1 >>
rect 19 260 20 261 
<< m1 >>
rect 22 260 23 261 
<< m1 >>
rect 44 260 45 261 
<< m1 >>
rect 55 260 56 261 
<< m1 >>
rect 64 260 65 261 
<< m1 >>
rect 91 260 92 261 
<< m2 >>
rect 92 260 93 261 
<< m2 >>
rect 109 260 110 261 
<< m2 >>
rect 110 260 111 261 
<< m2 >>
rect 111 260 112 261 
<< m2 >>
rect 112 260 113 261 
<< m2 >>
rect 113 260 114 261 
<< m2 >>
rect 114 260 115 261 
<< m2 >>
rect 115 260 116 261 
<< m2 >>
rect 116 260 117 261 
<< m2 >>
rect 117 260 118 261 
<< m2 >>
rect 118 260 119 261 
<< m1 >>
rect 142 260 143 261 
<< m1 >>
rect 148 260 149 261 
<< m1 >>
rect 150 260 151 261 
<< m2 >>
rect 158 260 159 261 
<< m2 >>
rect 163 260 164 261 
<< m2 >>
rect 177 260 178 261 
<< m1 >>
rect 181 260 182 261 
<< m2 >>
rect 186 260 187 261 
<< m2 >>
rect 190 260 191 261 
<< m2 >>
rect 192 260 193 261 
<< m2 >>
rect 217 260 218 261 
<< m2 >>
rect 219 260 220 261 
<< m2 >>
rect 231 260 232 261 
<< m1 >>
rect 235 260 236 261 
<< m1 >>
rect 237 260 238 261 
<< m2 >>
rect 253 260 254 261 
<< m2 >>
rect 255 260 256 261 
<< m2 >>
rect 259 260 260 261 
<< m2 >>
rect 262 260 263 261 
<< m2 >>
rect 264 260 265 261 
<< m1 >>
rect 280 260 281 261 
<< m2 >>
rect 303 260 304 261 
<< m1 >>
rect 307 260 308 261 
<< m1 >>
rect 309 260 310 261 
<< m2 >>
rect 322 260 323 261 
<< m2 >>
rect 340 260 341 261 
<< m2 >>
rect 342 260 343 261 
<< m2 >>
rect 346 260 347 261 
<< m2 >>
rect 366 260 367 261 
<< m2 >>
rect 372 260 373 261 
<< m1 >>
rect 386 260 387 261 
<< m1 >>
rect 397 260 398 261 
<< m1 >>
rect 416 260 417 261 
<< m1 >>
rect 419 260 420 261 
<< m2 >>
rect 420 260 421 261 
<< m1 >>
rect 430 260 431 261 
<< m1 >>
rect 437 260 438 261 
<< m1 >>
rect 442 260 443 261 
<< m1 >>
rect 484 260 485 261 
<< m1 >>
rect 523 260 524 261 
<< m1 >>
rect 19 261 20 262 
<< m1 >>
rect 22 261 23 262 
<< m1 >>
rect 44 261 45 262 
<< m1 >>
rect 55 261 56 262 
<< m1 >>
rect 64 261 65 262 
<< m1 >>
rect 91 261 92 262 
<< m2 >>
rect 92 261 93 262 
<< m1 >>
rect 109 261 110 262 
<< m2 >>
rect 109 261 110 262 
<< m2c >>
rect 109 261 110 262 
<< m1 >>
rect 109 261 110 262 
<< m2 >>
rect 109 261 110 262 
<< m2 >>
rect 141 261 142 262 
<< m1 >>
rect 142 261 143 262 
<< m2 >>
rect 142 261 143 262 
<< m2 >>
rect 143 261 144 262 
<< m1 >>
rect 144 261 145 262 
<< m2 >>
rect 144 261 145 262 
<< m2c >>
rect 144 261 145 262 
<< m1 >>
rect 144 261 145 262 
<< m2 >>
rect 144 261 145 262 
<< m1 >>
rect 145 261 146 262 
<< m1 >>
rect 146 261 147 262 
<< m2 >>
rect 146 261 147 262 
<< m2c >>
rect 146 261 147 262 
<< m1 >>
rect 146 261 147 262 
<< m2 >>
rect 146 261 147 262 
<< m2 >>
rect 147 261 148 262 
<< m1 >>
rect 148 261 149 262 
<< m2 >>
rect 148 261 149 262 
<< m2 >>
rect 149 261 150 262 
<< m1 >>
rect 150 261 151 262 
<< m2 >>
rect 150 261 151 262 
<< m2c >>
rect 150 261 151 262 
<< m1 >>
rect 150 261 151 262 
<< m2 >>
rect 150 261 151 262 
<< m1 >>
rect 158 261 159 262 
<< m2 >>
rect 158 261 159 262 
<< m2c >>
rect 158 261 159 262 
<< m1 >>
rect 158 261 159 262 
<< m2 >>
rect 158 261 159 262 
<< m1 >>
rect 159 261 160 262 
<< m1 >>
rect 160 261 161 262 
<< m1 >>
rect 163 261 164 262 
<< m2 >>
rect 163 261 164 262 
<< m2c >>
rect 163 261 164 262 
<< m1 >>
rect 163 261 164 262 
<< m2 >>
rect 163 261 164 262 
<< m1 >>
rect 177 261 178 262 
<< m2 >>
rect 177 261 178 262 
<< m2c >>
rect 177 261 178 262 
<< m1 >>
rect 177 261 178 262 
<< m2 >>
rect 177 261 178 262 
<< m1 >>
rect 178 261 179 262 
<< m1 >>
rect 181 261 182 262 
<< m2 >>
rect 182 261 183 262 
<< m1 >>
rect 183 261 184 262 
<< m2 >>
rect 183 261 184 262 
<< m2c >>
rect 183 261 184 262 
<< m1 >>
rect 183 261 184 262 
<< m2 >>
rect 183 261 184 262 
<< m1 >>
rect 184 261 185 262 
<< m1 >>
rect 185 261 186 262 
<< m1 >>
rect 186 261 187 262 
<< m2 >>
rect 186 261 187 262 
<< m1 >>
rect 187 261 188 262 
<< m1 >>
rect 188 261 189 262 
<< m1 >>
rect 189 261 190 262 
<< m1 >>
rect 190 261 191 262 
<< m2 >>
rect 190 261 191 262 
<< m1 >>
rect 191 261 192 262 
<< m1 >>
rect 192 261 193 262 
<< m2 >>
rect 192 261 193 262 
<< m2c >>
rect 192 261 193 262 
<< m1 >>
rect 192 261 193 262 
<< m2 >>
rect 192 261 193 262 
<< m2 >>
rect 217 261 218 262 
<< m1 >>
rect 219 261 220 262 
<< m2 >>
rect 219 261 220 262 
<< m2c >>
rect 219 261 220 262 
<< m1 >>
rect 219 261 220 262 
<< m2 >>
rect 219 261 220 262 
<< m2 >>
rect 231 261 232 262 
<< m2 >>
rect 232 261 233 262 
<< m2 >>
rect 233 261 234 262 
<< m2 >>
rect 234 261 235 262 
<< m1 >>
rect 235 261 236 262 
<< m2 >>
rect 235 261 236 262 
<< m2 >>
rect 236 261 237 262 
<< m1 >>
rect 237 261 238 262 
<< m2 >>
rect 237 261 238 262 
<< m2 >>
rect 238 261 239 262 
<< m1 >>
rect 253 261 254 262 
<< m2 >>
rect 253 261 254 262 
<< m2c >>
rect 253 261 254 262 
<< m1 >>
rect 253 261 254 262 
<< m2 >>
rect 253 261 254 262 
<< m1 >>
rect 255 261 256 262 
<< m2 >>
rect 255 261 256 262 
<< m2c >>
rect 255 261 256 262 
<< m1 >>
rect 255 261 256 262 
<< m2 >>
rect 255 261 256 262 
<< m1 >>
rect 259 261 260 262 
<< m2 >>
rect 259 261 260 262 
<< m2c >>
rect 259 261 260 262 
<< m1 >>
rect 259 261 260 262 
<< m2 >>
rect 259 261 260 262 
<< m1 >>
rect 262 261 263 262 
<< m2 >>
rect 262 261 263 262 
<< m1 >>
rect 263 261 264 262 
<< m1 >>
rect 264 261 265 262 
<< m2 >>
rect 264 261 265 262 
<< m2c >>
rect 264 261 265 262 
<< m1 >>
rect 264 261 265 262 
<< m2 >>
rect 264 261 265 262 
<< m1 >>
rect 280 261 281 262 
<< m1 >>
rect 283 261 284 262 
<< m1 >>
rect 284 261 285 262 
<< m1 >>
rect 285 261 286 262 
<< m1 >>
rect 286 261 287 262 
<< m1 >>
rect 287 261 288 262 
<< m1 >>
rect 303 261 304 262 
<< m2 >>
rect 303 261 304 262 
<< m2c >>
rect 303 261 304 262 
<< m1 >>
rect 303 261 304 262 
<< m2 >>
rect 303 261 304 262 
<< m1 >>
rect 304 261 305 262 
<< m1 >>
rect 305 261 306 262 
<< m1 >>
rect 307 261 308 262 
<< m1 >>
rect 309 261 310 262 
<< m1 >>
rect 322 261 323 262 
<< m2 >>
rect 322 261 323 262 
<< m2c >>
rect 322 261 323 262 
<< m1 >>
rect 322 261 323 262 
<< m2 >>
rect 322 261 323 262 
<< m1 >>
rect 340 261 341 262 
<< m2 >>
rect 340 261 341 262 
<< m2c >>
rect 340 261 341 262 
<< m1 >>
rect 340 261 341 262 
<< m2 >>
rect 340 261 341 262 
<< m1 >>
rect 342 261 343 262 
<< m2 >>
rect 342 261 343 262 
<< m2c >>
rect 342 261 343 262 
<< m1 >>
rect 342 261 343 262 
<< m2 >>
rect 342 261 343 262 
<< m1 >>
rect 343 261 344 262 
<< m1 >>
rect 344 261 345 262 
<< m1 >>
rect 346 261 347 262 
<< m2 >>
rect 346 261 347 262 
<< m2c >>
rect 346 261 347 262 
<< m1 >>
rect 346 261 347 262 
<< m2 >>
rect 346 261 347 262 
<< m1 >>
rect 358 261 359 262 
<< m1 >>
rect 359 261 360 262 
<< m1 >>
rect 360 261 361 262 
<< m1 >>
rect 361 261 362 262 
<< m1 >>
rect 362 261 363 262 
<< m1 >>
rect 363 261 364 262 
<< m1 >>
rect 364 261 365 262 
<< m1 >>
rect 365 261 366 262 
<< m1 >>
rect 366 261 367 262 
<< m2 >>
rect 366 261 367 262 
<< m1 >>
rect 367 261 368 262 
<< m1 >>
rect 368 261 369 262 
<< m2 >>
rect 368 261 369 262 
<< m2c >>
rect 368 261 369 262 
<< m1 >>
rect 368 261 369 262 
<< m2 >>
rect 368 261 369 262 
<< m2 >>
rect 369 261 370 262 
<< m2 >>
rect 370 261 371 262 
<< m2 >>
rect 371 261 372 262 
<< m2 >>
rect 372 261 373 262 
<< m1 >>
rect 386 261 387 262 
<< m1 >>
rect 397 261 398 262 
<< m1 >>
rect 416 261 417 262 
<< m1 >>
rect 419 261 420 262 
<< m2 >>
rect 420 261 421 262 
<< m1 >>
rect 430 261 431 262 
<< m1 >>
rect 437 261 438 262 
<< m1 >>
rect 442 261 443 262 
<< m1 >>
rect 484 261 485 262 
<< m1 >>
rect 523 261 524 262 
<< m1 >>
rect 19 262 20 263 
<< m1 >>
rect 22 262 23 263 
<< m1 >>
rect 44 262 45 263 
<< m1 >>
rect 55 262 56 263 
<< m1 >>
rect 64 262 65 263 
<< m1 >>
rect 91 262 92 263 
<< m2 >>
rect 92 262 93 263 
<< m1 >>
rect 109 262 110 263 
<< m1 >>
rect 139 262 140 263 
<< m1 >>
rect 140 262 141 263 
<< m2 >>
rect 140 262 141 263 
<< m2c >>
rect 140 262 141 263 
<< m1 >>
rect 140 262 141 263 
<< m2 >>
rect 140 262 141 263 
<< m2 >>
rect 141 262 142 263 
<< m1 >>
rect 142 262 143 263 
<< m1 >>
rect 148 262 149 263 
<< m1 >>
rect 160 262 161 263 
<< m1 >>
rect 163 262 164 263 
<< m1 >>
rect 178 262 179 263 
<< m1 >>
rect 181 262 182 263 
<< m2 >>
rect 182 262 183 263 
<< m2 >>
rect 186 262 187 263 
<< m2 >>
rect 190 262 191 263 
<< m1 >>
rect 196 262 197 263 
<< m1 >>
rect 197 262 198 263 
<< m1 >>
rect 198 262 199 263 
<< m1 >>
rect 199 262 200 263 
<< m1 >>
rect 214 262 215 263 
<< m1 >>
rect 215 262 216 263 
<< m1 >>
rect 216 262 217 263 
<< m1 >>
rect 217 262 218 263 
<< m2 >>
rect 217 262 218 263 
<< m1 >>
rect 219 262 220 263 
<< m1 >>
rect 232 262 233 263 
<< m1 >>
rect 233 262 234 263 
<< m1 >>
rect 234 262 235 263 
<< m1 >>
rect 235 262 236 263 
<< m1 >>
rect 237 262 238 263 
<< m2 >>
rect 238 262 239 263 
<< m1 >>
rect 253 262 254 263 
<< m1 >>
rect 255 262 256 263 
<< m1 >>
rect 259 262 260 263 
<< m1 >>
rect 262 262 263 263 
<< m2 >>
rect 262 262 263 263 
<< m1 >>
rect 280 262 281 263 
<< m1 >>
rect 283 262 284 263 
<< m1 >>
rect 287 262 288 263 
<< m2 >>
rect 287 262 288 263 
<< m2c >>
rect 287 262 288 263 
<< m1 >>
rect 287 262 288 263 
<< m2 >>
rect 287 262 288 263 
<< m2 >>
rect 288 262 289 263 
<< m1 >>
rect 289 262 290 263 
<< m2 >>
rect 289 262 290 263 
<< m1 >>
rect 290 262 291 263 
<< m1 >>
rect 291 262 292 263 
<< m1 >>
rect 292 262 293 263 
<< m1 >>
rect 293 262 294 263 
<< m1 >>
rect 294 262 295 263 
<< m1 >>
rect 295 262 296 263 
<< m1 >>
rect 296 262 297 263 
<< m1 >>
rect 297 262 298 263 
<< m1 >>
rect 298 262 299 263 
<< m1 >>
rect 299 262 300 263 
<< m1 >>
rect 300 262 301 263 
<< m1 >>
rect 301 262 302 263 
<< m1 >>
rect 305 262 306 263 
<< m2 >>
rect 305 262 306 263 
<< m2c >>
rect 305 262 306 263 
<< m1 >>
rect 305 262 306 263 
<< m2 >>
rect 305 262 306 263 
<< m2 >>
rect 306 262 307 263 
<< m1 >>
rect 307 262 308 263 
<< m2 >>
rect 307 262 308 263 
<< m2 >>
rect 308 262 309 263 
<< m1 >>
rect 309 262 310 263 
<< m2 >>
rect 309 262 310 263 
<< m2 >>
rect 310 262 311 263 
<< m1 >>
rect 322 262 323 263 
<< m1 >>
rect 340 262 341 263 
<< m1 >>
rect 344 262 345 263 
<< m1 >>
rect 346 262 347 263 
<< m1 >>
rect 358 262 359 263 
<< m2 >>
rect 366 262 367 263 
<< m1 >>
rect 370 262 371 263 
<< m1 >>
rect 371 262 372 263 
<< m1 >>
rect 372 262 373 263 
<< m1 >>
rect 373 262 374 263 
<< m1 >>
rect 386 262 387 263 
<< m1 >>
rect 388 262 389 263 
<< m1 >>
rect 389 262 390 263 
<< m1 >>
rect 390 262 391 263 
<< m1 >>
rect 391 262 392 263 
<< m1 >>
rect 397 262 398 263 
<< m1 >>
rect 416 262 417 263 
<< m1 >>
rect 419 262 420 263 
<< m2 >>
rect 420 262 421 263 
<< m1 >>
rect 430 262 431 263 
<< m1 >>
rect 437 262 438 263 
<< m1 >>
rect 442 262 443 263 
<< m1 >>
rect 484 262 485 263 
<< m1 >>
rect 523 262 524 263 
<< m1 >>
rect 19 263 20 264 
<< m1 >>
rect 22 263 23 264 
<< m1 >>
rect 44 263 45 264 
<< m1 >>
rect 55 263 56 264 
<< m1 >>
rect 64 263 65 264 
<< m1 >>
rect 91 263 92 264 
<< m2 >>
rect 92 263 93 264 
<< m1 >>
rect 109 263 110 264 
<< m1 >>
rect 139 263 140 264 
<< m1 >>
rect 142 263 143 264 
<< m1 >>
rect 148 263 149 264 
<< m1 >>
rect 160 263 161 264 
<< m1 >>
rect 163 263 164 264 
<< m1 >>
rect 178 263 179 264 
<< m1 >>
rect 181 263 182 264 
<< m2 >>
rect 182 263 183 264 
<< m1 >>
rect 186 263 187 264 
<< m2 >>
rect 186 263 187 264 
<< m2c >>
rect 186 263 187 264 
<< m1 >>
rect 186 263 187 264 
<< m2 >>
rect 186 263 187 264 
<< m1 >>
rect 190 263 191 264 
<< m2 >>
rect 190 263 191 264 
<< m2c >>
rect 190 263 191 264 
<< m1 >>
rect 190 263 191 264 
<< m2 >>
rect 190 263 191 264 
<< m1 >>
rect 196 263 197 264 
<< m1 >>
rect 199 263 200 264 
<< m1 >>
rect 214 263 215 264 
<< m1 >>
rect 217 263 218 264 
<< m2 >>
rect 217 263 218 264 
<< m1 >>
rect 219 263 220 264 
<< m1 >>
rect 232 263 233 264 
<< m1 >>
rect 237 263 238 264 
<< m2 >>
rect 238 263 239 264 
<< m1 >>
rect 253 263 254 264 
<< m1 >>
rect 255 263 256 264 
<< m1 >>
rect 259 263 260 264 
<< m1 >>
rect 262 263 263 264 
<< m2 >>
rect 262 263 263 264 
<< m1 >>
rect 280 263 281 264 
<< m1 >>
rect 283 263 284 264 
<< m1 >>
rect 289 263 290 264 
<< m2 >>
rect 289 263 290 264 
<< m1 >>
rect 301 263 302 264 
<< m1 >>
rect 307 263 308 264 
<< m1 >>
rect 309 263 310 264 
<< m2 >>
rect 310 263 311 264 
<< m1 >>
rect 322 263 323 264 
<< m1 >>
rect 340 263 341 264 
<< m1 >>
rect 344 263 345 264 
<< m1 >>
rect 346 263 347 264 
<< m1 >>
rect 358 263 359 264 
<< m1 >>
rect 366 263 367 264 
<< m2 >>
rect 366 263 367 264 
<< m2c >>
rect 366 263 367 264 
<< m1 >>
rect 366 263 367 264 
<< m2 >>
rect 366 263 367 264 
<< m1 >>
rect 370 263 371 264 
<< m1 >>
rect 373 263 374 264 
<< m1 >>
rect 386 263 387 264 
<< m1 >>
rect 388 263 389 264 
<< m1 >>
rect 391 263 392 264 
<< m1 >>
rect 397 263 398 264 
<< m1 >>
rect 416 263 417 264 
<< m1 >>
rect 419 263 420 264 
<< m2 >>
rect 420 263 421 264 
<< m1 >>
rect 430 263 431 264 
<< m1 >>
rect 437 263 438 264 
<< m1 >>
rect 442 263 443 264 
<< m1 >>
rect 484 263 485 264 
<< m1 >>
rect 523 263 524 264 
<< pdiffusion >>
rect 12 264 13 265 
<< pdiffusion >>
rect 13 264 14 265 
<< pdiffusion >>
rect 14 264 15 265 
<< pdiffusion >>
rect 15 264 16 265 
<< pdiffusion >>
rect 16 264 17 265 
<< pdiffusion >>
rect 17 264 18 265 
<< m1 >>
rect 19 264 20 265 
<< m1 >>
rect 22 264 23 265 
<< m1 >>
rect 44 264 45 265 
<< pdiffusion >>
rect 48 264 49 265 
<< pdiffusion >>
rect 49 264 50 265 
<< pdiffusion >>
rect 50 264 51 265 
<< pdiffusion >>
rect 51 264 52 265 
<< pdiffusion >>
rect 52 264 53 265 
<< pdiffusion >>
rect 53 264 54 265 
<< m1 >>
rect 55 264 56 265 
<< m1 >>
rect 64 264 65 265 
<< pdiffusion >>
rect 66 264 67 265 
<< pdiffusion >>
rect 67 264 68 265 
<< pdiffusion >>
rect 68 264 69 265 
<< pdiffusion >>
rect 69 264 70 265 
<< pdiffusion >>
rect 70 264 71 265 
<< pdiffusion >>
rect 71 264 72 265 
<< pdiffusion >>
rect 84 264 85 265 
<< pdiffusion >>
rect 85 264 86 265 
<< pdiffusion >>
rect 86 264 87 265 
<< pdiffusion >>
rect 87 264 88 265 
<< pdiffusion >>
rect 88 264 89 265 
<< pdiffusion >>
rect 89 264 90 265 
<< m1 >>
rect 91 264 92 265 
<< m2 >>
rect 92 264 93 265 
<< pdiffusion >>
rect 102 264 103 265 
<< pdiffusion >>
rect 103 264 104 265 
<< pdiffusion >>
rect 104 264 105 265 
<< pdiffusion >>
rect 105 264 106 265 
<< pdiffusion >>
rect 106 264 107 265 
<< pdiffusion >>
rect 107 264 108 265 
<< m1 >>
rect 109 264 110 265 
<< pdiffusion >>
rect 120 264 121 265 
<< pdiffusion >>
rect 121 264 122 265 
<< pdiffusion >>
rect 122 264 123 265 
<< pdiffusion >>
rect 123 264 124 265 
<< pdiffusion >>
rect 124 264 125 265 
<< pdiffusion >>
rect 125 264 126 265 
<< pdiffusion >>
rect 138 264 139 265 
<< m1 >>
rect 139 264 140 265 
<< pdiffusion >>
rect 139 264 140 265 
<< pdiffusion >>
rect 140 264 141 265 
<< pdiffusion >>
rect 141 264 142 265 
<< m1 >>
rect 142 264 143 265 
<< pdiffusion >>
rect 142 264 143 265 
<< pdiffusion >>
rect 143 264 144 265 
<< m1 >>
rect 148 264 149 265 
<< pdiffusion >>
rect 156 264 157 265 
<< pdiffusion >>
rect 157 264 158 265 
<< pdiffusion >>
rect 158 264 159 265 
<< pdiffusion >>
rect 159 264 160 265 
<< m1 >>
rect 160 264 161 265 
<< pdiffusion >>
rect 160 264 161 265 
<< pdiffusion >>
rect 161 264 162 265 
<< m1 >>
rect 163 264 164 265 
<< pdiffusion >>
rect 174 264 175 265 
<< pdiffusion >>
rect 175 264 176 265 
<< pdiffusion >>
rect 176 264 177 265 
<< pdiffusion >>
rect 177 264 178 265 
<< m1 >>
rect 178 264 179 265 
<< pdiffusion >>
rect 178 264 179 265 
<< pdiffusion >>
rect 179 264 180 265 
<< m1 >>
rect 181 264 182 265 
<< m2 >>
rect 182 264 183 265 
<< m1 >>
rect 186 264 187 265 
<< m1 >>
rect 190 264 191 265 
<< pdiffusion >>
rect 192 264 193 265 
<< pdiffusion >>
rect 193 264 194 265 
<< pdiffusion >>
rect 194 264 195 265 
<< pdiffusion >>
rect 195 264 196 265 
<< m1 >>
rect 196 264 197 265 
<< pdiffusion >>
rect 196 264 197 265 
<< pdiffusion >>
rect 197 264 198 265 
<< m1 >>
rect 199 264 200 265 
<< pdiffusion >>
rect 210 264 211 265 
<< pdiffusion >>
rect 211 264 212 265 
<< pdiffusion >>
rect 212 264 213 265 
<< pdiffusion >>
rect 213 264 214 265 
<< m1 >>
rect 214 264 215 265 
<< pdiffusion >>
rect 214 264 215 265 
<< pdiffusion >>
rect 215 264 216 265 
<< m1 >>
rect 217 264 218 265 
<< m2 >>
rect 217 264 218 265 
<< m1 >>
rect 219 264 220 265 
<< pdiffusion >>
rect 228 264 229 265 
<< pdiffusion >>
rect 229 264 230 265 
<< pdiffusion >>
rect 230 264 231 265 
<< pdiffusion >>
rect 231 264 232 265 
<< m1 >>
rect 232 264 233 265 
<< pdiffusion >>
rect 232 264 233 265 
<< pdiffusion >>
rect 233 264 234 265 
<< m1 >>
rect 237 264 238 265 
<< m2 >>
rect 238 264 239 265 
<< pdiffusion >>
rect 246 264 247 265 
<< pdiffusion >>
rect 247 264 248 265 
<< pdiffusion >>
rect 248 264 249 265 
<< pdiffusion >>
rect 249 264 250 265 
<< pdiffusion >>
rect 250 264 251 265 
<< pdiffusion >>
rect 251 264 252 265 
<< m1 >>
rect 253 264 254 265 
<< m1 >>
rect 255 264 256 265 
<< m1 >>
rect 259 264 260 265 
<< m1 >>
rect 262 264 263 265 
<< m2 >>
rect 262 264 263 265 
<< pdiffusion >>
rect 264 264 265 265 
<< pdiffusion >>
rect 265 264 266 265 
<< pdiffusion >>
rect 266 264 267 265 
<< pdiffusion >>
rect 267 264 268 265 
<< pdiffusion >>
rect 268 264 269 265 
<< pdiffusion >>
rect 269 264 270 265 
<< m1 >>
rect 280 264 281 265 
<< pdiffusion >>
rect 282 264 283 265 
<< m1 >>
rect 283 264 284 265 
<< pdiffusion >>
rect 283 264 284 265 
<< pdiffusion >>
rect 284 264 285 265 
<< pdiffusion >>
rect 285 264 286 265 
<< pdiffusion >>
rect 286 264 287 265 
<< pdiffusion >>
rect 287 264 288 265 
<< m1 >>
rect 289 264 290 265 
<< m2 >>
rect 289 264 290 265 
<< pdiffusion >>
rect 300 264 301 265 
<< m1 >>
rect 301 264 302 265 
<< pdiffusion >>
rect 301 264 302 265 
<< pdiffusion >>
rect 302 264 303 265 
<< pdiffusion >>
rect 303 264 304 265 
<< pdiffusion >>
rect 304 264 305 265 
<< pdiffusion >>
rect 305 264 306 265 
<< m1 >>
rect 307 264 308 265 
<< m1 >>
rect 309 264 310 265 
<< m2 >>
rect 310 264 311 265 
<< pdiffusion >>
rect 318 264 319 265 
<< pdiffusion >>
rect 319 264 320 265 
<< pdiffusion >>
rect 320 264 321 265 
<< pdiffusion >>
rect 321 264 322 265 
<< m1 >>
rect 322 264 323 265 
<< pdiffusion >>
rect 322 264 323 265 
<< pdiffusion >>
rect 323 264 324 265 
<< pdiffusion >>
rect 336 264 337 265 
<< pdiffusion >>
rect 337 264 338 265 
<< pdiffusion >>
rect 338 264 339 265 
<< pdiffusion >>
rect 339 264 340 265 
<< m1 >>
rect 340 264 341 265 
<< pdiffusion >>
rect 340 264 341 265 
<< pdiffusion >>
rect 341 264 342 265 
<< m1 >>
rect 344 264 345 265 
<< m1 >>
rect 346 264 347 265 
<< pdiffusion >>
rect 354 264 355 265 
<< pdiffusion >>
rect 355 264 356 265 
<< pdiffusion >>
rect 356 264 357 265 
<< pdiffusion >>
rect 357 264 358 265 
<< m1 >>
rect 358 264 359 265 
<< pdiffusion >>
rect 358 264 359 265 
<< pdiffusion >>
rect 359 264 360 265 
<< m1 >>
rect 366 264 367 265 
<< m1 >>
rect 370 264 371 265 
<< pdiffusion >>
rect 372 264 373 265 
<< m1 >>
rect 373 264 374 265 
<< pdiffusion >>
rect 373 264 374 265 
<< pdiffusion >>
rect 374 264 375 265 
<< pdiffusion >>
rect 375 264 376 265 
<< pdiffusion >>
rect 376 264 377 265 
<< pdiffusion >>
rect 377 264 378 265 
<< m1 >>
rect 386 264 387 265 
<< m1 >>
rect 388 264 389 265 
<< pdiffusion >>
rect 390 264 391 265 
<< m1 >>
rect 391 264 392 265 
<< pdiffusion >>
rect 391 264 392 265 
<< pdiffusion >>
rect 392 264 393 265 
<< pdiffusion >>
rect 393 264 394 265 
<< pdiffusion >>
rect 394 264 395 265 
<< pdiffusion >>
rect 395 264 396 265 
<< m1 >>
rect 397 264 398 265 
<< pdiffusion >>
rect 408 264 409 265 
<< pdiffusion >>
rect 409 264 410 265 
<< pdiffusion >>
rect 410 264 411 265 
<< pdiffusion >>
rect 411 264 412 265 
<< pdiffusion >>
rect 412 264 413 265 
<< pdiffusion >>
rect 413 264 414 265 
<< m1 >>
rect 416 264 417 265 
<< m1 >>
rect 419 264 420 265 
<< m2 >>
rect 420 264 421 265 
<< pdiffusion >>
rect 426 264 427 265 
<< pdiffusion >>
rect 427 264 428 265 
<< pdiffusion >>
rect 428 264 429 265 
<< pdiffusion >>
rect 429 264 430 265 
<< m1 >>
rect 430 264 431 265 
<< pdiffusion >>
rect 430 264 431 265 
<< pdiffusion >>
rect 431 264 432 265 
<< m1 >>
rect 437 264 438 265 
<< m1 >>
rect 442 264 443 265 
<< pdiffusion >>
rect 444 264 445 265 
<< pdiffusion >>
rect 445 264 446 265 
<< pdiffusion >>
rect 446 264 447 265 
<< pdiffusion >>
rect 447 264 448 265 
<< pdiffusion >>
rect 448 264 449 265 
<< pdiffusion >>
rect 449 264 450 265 
<< pdiffusion >>
rect 462 264 463 265 
<< pdiffusion >>
rect 463 264 464 265 
<< pdiffusion >>
rect 464 264 465 265 
<< pdiffusion >>
rect 465 264 466 265 
<< pdiffusion >>
rect 466 264 467 265 
<< pdiffusion >>
rect 467 264 468 265 
<< pdiffusion >>
rect 480 264 481 265 
<< pdiffusion >>
rect 481 264 482 265 
<< pdiffusion >>
rect 482 264 483 265 
<< pdiffusion >>
rect 483 264 484 265 
<< m1 >>
rect 484 264 485 265 
<< pdiffusion >>
rect 484 264 485 265 
<< pdiffusion >>
rect 485 264 486 265 
<< pdiffusion >>
rect 498 264 499 265 
<< pdiffusion >>
rect 499 264 500 265 
<< pdiffusion >>
rect 500 264 501 265 
<< pdiffusion >>
rect 501 264 502 265 
<< pdiffusion >>
rect 502 264 503 265 
<< pdiffusion >>
rect 503 264 504 265 
<< pdiffusion >>
rect 516 264 517 265 
<< pdiffusion >>
rect 517 264 518 265 
<< pdiffusion >>
rect 518 264 519 265 
<< pdiffusion >>
rect 519 264 520 265 
<< pdiffusion >>
rect 520 264 521 265 
<< pdiffusion >>
rect 521 264 522 265 
<< m1 >>
rect 523 264 524 265 
<< pdiffusion >>
rect 12 265 13 266 
<< pdiffusion >>
rect 13 265 14 266 
<< pdiffusion >>
rect 14 265 15 266 
<< pdiffusion >>
rect 15 265 16 266 
<< pdiffusion >>
rect 16 265 17 266 
<< pdiffusion >>
rect 17 265 18 266 
<< m1 >>
rect 19 265 20 266 
<< m1 >>
rect 22 265 23 266 
<< m1 >>
rect 44 265 45 266 
<< pdiffusion >>
rect 48 265 49 266 
<< pdiffusion >>
rect 49 265 50 266 
<< pdiffusion >>
rect 50 265 51 266 
<< pdiffusion >>
rect 51 265 52 266 
<< pdiffusion >>
rect 52 265 53 266 
<< pdiffusion >>
rect 53 265 54 266 
<< m1 >>
rect 55 265 56 266 
<< m1 >>
rect 64 265 65 266 
<< pdiffusion >>
rect 66 265 67 266 
<< pdiffusion >>
rect 67 265 68 266 
<< pdiffusion >>
rect 68 265 69 266 
<< pdiffusion >>
rect 69 265 70 266 
<< pdiffusion >>
rect 70 265 71 266 
<< pdiffusion >>
rect 71 265 72 266 
<< pdiffusion >>
rect 84 265 85 266 
<< pdiffusion >>
rect 85 265 86 266 
<< pdiffusion >>
rect 86 265 87 266 
<< pdiffusion >>
rect 87 265 88 266 
<< pdiffusion >>
rect 88 265 89 266 
<< pdiffusion >>
rect 89 265 90 266 
<< m1 >>
rect 91 265 92 266 
<< m2 >>
rect 92 265 93 266 
<< pdiffusion >>
rect 102 265 103 266 
<< pdiffusion >>
rect 103 265 104 266 
<< pdiffusion >>
rect 104 265 105 266 
<< pdiffusion >>
rect 105 265 106 266 
<< pdiffusion >>
rect 106 265 107 266 
<< pdiffusion >>
rect 107 265 108 266 
<< m1 >>
rect 109 265 110 266 
<< pdiffusion >>
rect 120 265 121 266 
<< pdiffusion >>
rect 121 265 122 266 
<< pdiffusion >>
rect 122 265 123 266 
<< pdiffusion >>
rect 123 265 124 266 
<< pdiffusion >>
rect 124 265 125 266 
<< pdiffusion >>
rect 125 265 126 266 
<< pdiffusion >>
rect 138 265 139 266 
<< pdiffusion >>
rect 139 265 140 266 
<< pdiffusion >>
rect 140 265 141 266 
<< pdiffusion >>
rect 141 265 142 266 
<< pdiffusion >>
rect 142 265 143 266 
<< pdiffusion >>
rect 143 265 144 266 
<< m1 >>
rect 148 265 149 266 
<< pdiffusion >>
rect 156 265 157 266 
<< pdiffusion >>
rect 157 265 158 266 
<< pdiffusion >>
rect 158 265 159 266 
<< pdiffusion >>
rect 159 265 160 266 
<< pdiffusion >>
rect 160 265 161 266 
<< pdiffusion >>
rect 161 265 162 266 
<< m1 >>
rect 163 265 164 266 
<< pdiffusion >>
rect 174 265 175 266 
<< pdiffusion >>
rect 175 265 176 266 
<< pdiffusion >>
rect 176 265 177 266 
<< pdiffusion >>
rect 177 265 178 266 
<< pdiffusion >>
rect 178 265 179 266 
<< pdiffusion >>
rect 179 265 180 266 
<< m1 >>
rect 181 265 182 266 
<< m2 >>
rect 182 265 183 266 
<< m1 >>
rect 186 265 187 266 
<< m1 >>
rect 190 265 191 266 
<< pdiffusion >>
rect 192 265 193 266 
<< pdiffusion >>
rect 193 265 194 266 
<< pdiffusion >>
rect 194 265 195 266 
<< pdiffusion >>
rect 195 265 196 266 
<< pdiffusion >>
rect 196 265 197 266 
<< pdiffusion >>
rect 197 265 198 266 
<< m1 >>
rect 199 265 200 266 
<< pdiffusion >>
rect 210 265 211 266 
<< pdiffusion >>
rect 211 265 212 266 
<< pdiffusion >>
rect 212 265 213 266 
<< pdiffusion >>
rect 213 265 214 266 
<< pdiffusion >>
rect 214 265 215 266 
<< pdiffusion >>
rect 215 265 216 266 
<< m1 >>
rect 217 265 218 266 
<< m2 >>
rect 217 265 218 266 
<< m1 >>
rect 219 265 220 266 
<< pdiffusion >>
rect 228 265 229 266 
<< pdiffusion >>
rect 229 265 230 266 
<< pdiffusion >>
rect 230 265 231 266 
<< pdiffusion >>
rect 231 265 232 266 
<< pdiffusion >>
rect 232 265 233 266 
<< pdiffusion >>
rect 233 265 234 266 
<< m1 >>
rect 237 265 238 266 
<< m2 >>
rect 238 265 239 266 
<< pdiffusion >>
rect 246 265 247 266 
<< pdiffusion >>
rect 247 265 248 266 
<< pdiffusion >>
rect 248 265 249 266 
<< pdiffusion >>
rect 249 265 250 266 
<< pdiffusion >>
rect 250 265 251 266 
<< pdiffusion >>
rect 251 265 252 266 
<< m1 >>
rect 253 265 254 266 
<< m1 >>
rect 255 265 256 266 
<< m1 >>
rect 259 265 260 266 
<< m1 >>
rect 262 265 263 266 
<< m2 >>
rect 262 265 263 266 
<< pdiffusion >>
rect 264 265 265 266 
<< pdiffusion >>
rect 265 265 266 266 
<< pdiffusion >>
rect 266 265 267 266 
<< pdiffusion >>
rect 267 265 268 266 
<< pdiffusion >>
rect 268 265 269 266 
<< pdiffusion >>
rect 269 265 270 266 
<< m1 >>
rect 280 265 281 266 
<< pdiffusion >>
rect 282 265 283 266 
<< pdiffusion >>
rect 283 265 284 266 
<< pdiffusion >>
rect 284 265 285 266 
<< pdiffusion >>
rect 285 265 286 266 
<< pdiffusion >>
rect 286 265 287 266 
<< pdiffusion >>
rect 287 265 288 266 
<< m1 >>
rect 289 265 290 266 
<< m2 >>
rect 289 265 290 266 
<< pdiffusion >>
rect 300 265 301 266 
<< pdiffusion >>
rect 301 265 302 266 
<< pdiffusion >>
rect 302 265 303 266 
<< pdiffusion >>
rect 303 265 304 266 
<< pdiffusion >>
rect 304 265 305 266 
<< pdiffusion >>
rect 305 265 306 266 
<< m1 >>
rect 307 265 308 266 
<< m1 >>
rect 309 265 310 266 
<< m2 >>
rect 310 265 311 266 
<< pdiffusion >>
rect 318 265 319 266 
<< pdiffusion >>
rect 319 265 320 266 
<< pdiffusion >>
rect 320 265 321 266 
<< pdiffusion >>
rect 321 265 322 266 
<< pdiffusion >>
rect 322 265 323 266 
<< pdiffusion >>
rect 323 265 324 266 
<< pdiffusion >>
rect 336 265 337 266 
<< pdiffusion >>
rect 337 265 338 266 
<< pdiffusion >>
rect 338 265 339 266 
<< pdiffusion >>
rect 339 265 340 266 
<< pdiffusion >>
rect 340 265 341 266 
<< pdiffusion >>
rect 341 265 342 266 
<< m1 >>
rect 344 265 345 266 
<< m1 >>
rect 346 265 347 266 
<< pdiffusion >>
rect 354 265 355 266 
<< pdiffusion >>
rect 355 265 356 266 
<< pdiffusion >>
rect 356 265 357 266 
<< pdiffusion >>
rect 357 265 358 266 
<< pdiffusion >>
rect 358 265 359 266 
<< pdiffusion >>
rect 359 265 360 266 
<< m1 >>
rect 366 265 367 266 
<< m1 >>
rect 370 265 371 266 
<< pdiffusion >>
rect 372 265 373 266 
<< pdiffusion >>
rect 373 265 374 266 
<< pdiffusion >>
rect 374 265 375 266 
<< pdiffusion >>
rect 375 265 376 266 
<< pdiffusion >>
rect 376 265 377 266 
<< pdiffusion >>
rect 377 265 378 266 
<< m1 >>
rect 386 265 387 266 
<< m1 >>
rect 388 265 389 266 
<< pdiffusion >>
rect 390 265 391 266 
<< pdiffusion >>
rect 391 265 392 266 
<< pdiffusion >>
rect 392 265 393 266 
<< pdiffusion >>
rect 393 265 394 266 
<< pdiffusion >>
rect 394 265 395 266 
<< pdiffusion >>
rect 395 265 396 266 
<< m1 >>
rect 397 265 398 266 
<< pdiffusion >>
rect 408 265 409 266 
<< pdiffusion >>
rect 409 265 410 266 
<< pdiffusion >>
rect 410 265 411 266 
<< pdiffusion >>
rect 411 265 412 266 
<< pdiffusion >>
rect 412 265 413 266 
<< pdiffusion >>
rect 413 265 414 266 
<< m1 >>
rect 416 265 417 266 
<< m1 >>
rect 419 265 420 266 
<< m2 >>
rect 420 265 421 266 
<< pdiffusion >>
rect 426 265 427 266 
<< pdiffusion >>
rect 427 265 428 266 
<< pdiffusion >>
rect 428 265 429 266 
<< pdiffusion >>
rect 429 265 430 266 
<< pdiffusion >>
rect 430 265 431 266 
<< pdiffusion >>
rect 431 265 432 266 
<< m1 >>
rect 437 265 438 266 
<< m1 >>
rect 442 265 443 266 
<< pdiffusion >>
rect 444 265 445 266 
<< pdiffusion >>
rect 445 265 446 266 
<< pdiffusion >>
rect 446 265 447 266 
<< pdiffusion >>
rect 447 265 448 266 
<< pdiffusion >>
rect 448 265 449 266 
<< pdiffusion >>
rect 449 265 450 266 
<< pdiffusion >>
rect 462 265 463 266 
<< pdiffusion >>
rect 463 265 464 266 
<< pdiffusion >>
rect 464 265 465 266 
<< pdiffusion >>
rect 465 265 466 266 
<< pdiffusion >>
rect 466 265 467 266 
<< pdiffusion >>
rect 467 265 468 266 
<< pdiffusion >>
rect 480 265 481 266 
<< pdiffusion >>
rect 481 265 482 266 
<< pdiffusion >>
rect 482 265 483 266 
<< pdiffusion >>
rect 483 265 484 266 
<< pdiffusion >>
rect 484 265 485 266 
<< pdiffusion >>
rect 485 265 486 266 
<< pdiffusion >>
rect 498 265 499 266 
<< pdiffusion >>
rect 499 265 500 266 
<< pdiffusion >>
rect 500 265 501 266 
<< pdiffusion >>
rect 501 265 502 266 
<< pdiffusion >>
rect 502 265 503 266 
<< pdiffusion >>
rect 503 265 504 266 
<< pdiffusion >>
rect 516 265 517 266 
<< pdiffusion >>
rect 517 265 518 266 
<< pdiffusion >>
rect 518 265 519 266 
<< pdiffusion >>
rect 519 265 520 266 
<< pdiffusion >>
rect 520 265 521 266 
<< pdiffusion >>
rect 521 265 522 266 
<< m1 >>
rect 523 265 524 266 
<< pdiffusion >>
rect 12 266 13 267 
<< pdiffusion >>
rect 13 266 14 267 
<< pdiffusion >>
rect 14 266 15 267 
<< pdiffusion >>
rect 15 266 16 267 
<< pdiffusion >>
rect 16 266 17 267 
<< pdiffusion >>
rect 17 266 18 267 
<< m1 >>
rect 19 266 20 267 
<< m1 >>
rect 22 266 23 267 
<< m1 >>
rect 44 266 45 267 
<< pdiffusion >>
rect 48 266 49 267 
<< pdiffusion >>
rect 49 266 50 267 
<< pdiffusion >>
rect 50 266 51 267 
<< pdiffusion >>
rect 51 266 52 267 
<< pdiffusion >>
rect 52 266 53 267 
<< pdiffusion >>
rect 53 266 54 267 
<< m1 >>
rect 55 266 56 267 
<< m1 >>
rect 64 266 65 267 
<< pdiffusion >>
rect 66 266 67 267 
<< pdiffusion >>
rect 67 266 68 267 
<< pdiffusion >>
rect 68 266 69 267 
<< pdiffusion >>
rect 69 266 70 267 
<< pdiffusion >>
rect 70 266 71 267 
<< pdiffusion >>
rect 71 266 72 267 
<< pdiffusion >>
rect 84 266 85 267 
<< pdiffusion >>
rect 85 266 86 267 
<< pdiffusion >>
rect 86 266 87 267 
<< pdiffusion >>
rect 87 266 88 267 
<< pdiffusion >>
rect 88 266 89 267 
<< pdiffusion >>
rect 89 266 90 267 
<< m1 >>
rect 91 266 92 267 
<< m2 >>
rect 92 266 93 267 
<< pdiffusion >>
rect 102 266 103 267 
<< pdiffusion >>
rect 103 266 104 267 
<< pdiffusion >>
rect 104 266 105 267 
<< pdiffusion >>
rect 105 266 106 267 
<< pdiffusion >>
rect 106 266 107 267 
<< pdiffusion >>
rect 107 266 108 267 
<< m1 >>
rect 109 266 110 267 
<< pdiffusion >>
rect 120 266 121 267 
<< pdiffusion >>
rect 121 266 122 267 
<< pdiffusion >>
rect 122 266 123 267 
<< pdiffusion >>
rect 123 266 124 267 
<< pdiffusion >>
rect 124 266 125 267 
<< pdiffusion >>
rect 125 266 126 267 
<< pdiffusion >>
rect 138 266 139 267 
<< pdiffusion >>
rect 139 266 140 267 
<< pdiffusion >>
rect 140 266 141 267 
<< pdiffusion >>
rect 141 266 142 267 
<< pdiffusion >>
rect 142 266 143 267 
<< pdiffusion >>
rect 143 266 144 267 
<< m1 >>
rect 148 266 149 267 
<< pdiffusion >>
rect 156 266 157 267 
<< pdiffusion >>
rect 157 266 158 267 
<< pdiffusion >>
rect 158 266 159 267 
<< pdiffusion >>
rect 159 266 160 267 
<< pdiffusion >>
rect 160 266 161 267 
<< pdiffusion >>
rect 161 266 162 267 
<< m1 >>
rect 163 266 164 267 
<< pdiffusion >>
rect 174 266 175 267 
<< pdiffusion >>
rect 175 266 176 267 
<< pdiffusion >>
rect 176 266 177 267 
<< pdiffusion >>
rect 177 266 178 267 
<< pdiffusion >>
rect 178 266 179 267 
<< pdiffusion >>
rect 179 266 180 267 
<< m1 >>
rect 181 266 182 267 
<< m2 >>
rect 182 266 183 267 
<< m1 >>
rect 186 266 187 267 
<< m1 >>
rect 190 266 191 267 
<< pdiffusion >>
rect 192 266 193 267 
<< pdiffusion >>
rect 193 266 194 267 
<< pdiffusion >>
rect 194 266 195 267 
<< pdiffusion >>
rect 195 266 196 267 
<< pdiffusion >>
rect 196 266 197 267 
<< pdiffusion >>
rect 197 266 198 267 
<< m1 >>
rect 199 266 200 267 
<< pdiffusion >>
rect 210 266 211 267 
<< pdiffusion >>
rect 211 266 212 267 
<< pdiffusion >>
rect 212 266 213 267 
<< pdiffusion >>
rect 213 266 214 267 
<< pdiffusion >>
rect 214 266 215 267 
<< pdiffusion >>
rect 215 266 216 267 
<< m1 >>
rect 217 266 218 267 
<< m2 >>
rect 217 266 218 267 
<< m1 >>
rect 219 266 220 267 
<< pdiffusion >>
rect 228 266 229 267 
<< pdiffusion >>
rect 229 266 230 267 
<< pdiffusion >>
rect 230 266 231 267 
<< pdiffusion >>
rect 231 266 232 267 
<< pdiffusion >>
rect 232 266 233 267 
<< pdiffusion >>
rect 233 266 234 267 
<< m1 >>
rect 237 266 238 267 
<< m2 >>
rect 238 266 239 267 
<< pdiffusion >>
rect 246 266 247 267 
<< pdiffusion >>
rect 247 266 248 267 
<< pdiffusion >>
rect 248 266 249 267 
<< pdiffusion >>
rect 249 266 250 267 
<< pdiffusion >>
rect 250 266 251 267 
<< pdiffusion >>
rect 251 266 252 267 
<< m1 >>
rect 253 266 254 267 
<< m1 >>
rect 255 266 256 267 
<< m1 >>
rect 259 266 260 267 
<< m1 >>
rect 262 266 263 267 
<< m2 >>
rect 262 266 263 267 
<< pdiffusion >>
rect 264 266 265 267 
<< pdiffusion >>
rect 265 266 266 267 
<< pdiffusion >>
rect 266 266 267 267 
<< pdiffusion >>
rect 267 266 268 267 
<< pdiffusion >>
rect 268 266 269 267 
<< pdiffusion >>
rect 269 266 270 267 
<< m1 >>
rect 280 266 281 267 
<< pdiffusion >>
rect 282 266 283 267 
<< pdiffusion >>
rect 283 266 284 267 
<< pdiffusion >>
rect 284 266 285 267 
<< pdiffusion >>
rect 285 266 286 267 
<< pdiffusion >>
rect 286 266 287 267 
<< pdiffusion >>
rect 287 266 288 267 
<< m1 >>
rect 289 266 290 267 
<< m2 >>
rect 289 266 290 267 
<< pdiffusion >>
rect 300 266 301 267 
<< pdiffusion >>
rect 301 266 302 267 
<< pdiffusion >>
rect 302 266 303 267 
<< pdiffusion >>
rect 303 266 304 267 
<< pdiffusion >>
rect 304 266 305 267 
<< pdiffusion >>
rect 305 266 306 267 
<< m1 >>
rect 307 266 308 267 
<< m1 >>
rect 309 266 310 267 
<< m2 >>
rect 310 266 311 267 
<< pdiffusion >>
rect 318 266 319 267 
<< pdiffusion >>
rect 319 266 320 267 
<< pdiffusion >>
rect 320 266 321 267 
<< pdiffusion >>
rect 321 266 322 267 
<< pdiffusion >>
rect 322 266 323 267 
<< pdiffusion >>
rect 323 266 324 267 
<< pdiffusion >>
rect 336 266 337 267 
<< pdiffusion >>
rect 337 266 338 267 
<< pdiffusion >>
rect 338 266 339 267 
<< pdiffusion >>
rect 339 266 340 267 
<< pdiffusion >>
rect 340 266 341 267 
<< pdiffusion >>
rect 341 266 342 267 
<< m1 >>
rect 344 266 345 267 
<< m1 >>
rect 346 266 347 267 
<< pdiffusion >>
rect 354 266 355 267 
<< pdiffusion >>
rect 355 266 356 267 
<< pdiffusion >>
rect 356 266 357 267 
<< pdiffusion >>
rect 357 266 358 267 
<< pdiffusion >>
rect 358 266 359 267 
<< pdiffusion >>
rect 359 266 360 267 
<< m1 >>
rect 366 266 367 267 
<< m1 >>
rect 370 266 371 267 
<< pdiffusion >>
rect 372 266 373 267 
<< pdiffusion >>
rect 373 266 374 267 
<< pdiffusion >>
rect 374 266 375 267 
<< pdiffusion >>
rect 375 266 376 267 
<< pdiffusion >>
rect 376 266 377 267 
<< pdiffusion >>
rect 377 266 378 267 
<< m1 >>
rect 386 266 387 267 
<< m1 >>
rect 388 266 389 267 
<< pdiffusion >>
rect 390 266 391 267 
<< pdiffusion >>
rect 391 266 392 267 
<< pdiffusion >>
rect 392 266 393 267 
<< pdiffusion >>
rect 393 266 394 267 
<< pdiffusion >>
rect 394 266 395 267 
<< pdiffusion >>
rect 395 266 396 267 
<< m1 >>
rect 397 266 398 267 
<< pdiffusion >>
rect 408 266 409 267 
<< pdiffusion >>
rect 409 266 410 267 
<< pdiffusion >>
rect 410 266 411 267 
<< pdiffusion >>
rect 411 266 412 267 
<< pdiffusion >>
rect 412 266 413 267 
<< pdiffusion >>
rect 413 266 414 267 
<< m1 >>
rect 416 266 417 267 
<< m1 >>
rect 419 266 420 267 
<< m2 >>
rect 420 266 421 267 
<< pdiffusion >>
rect 426 266 427 267 
<< pdiffusion >>
rect 427 266 428 267 
<< pdiffusion >>
rect 428 266 429 267 
<< pdiffusion >>
rect 429 266 430 267 
<< pdiffusion >>
rect 430 266 431 267 
<< pdiffusion >>
rect 431 266 432 267 
<< m1 >>
rect 437 266 438 267 
<< m1 >>
rect 442 266 443 267 
<< pdiffusion >>
rect 444 266 445 267 
<< pdiffusion >>
rect 445 266 446 267 
<< pdiffusion >>
rect 446 266 447 267 
<< pdiffusion >>
rect 447 266 448 267 
<< pdiffusion >>
rect 448 266 449 267 
<< pdiffusion >>
rect 449 266 450 267 
<< pdiffusion >>
rect 462 266 463 267 
<< pdiffusion >>
rect 463 266 464 267 
<< pdiffusion >>
rect 464 266 465 267 
<< pdiffusion >>
rect 465 266 466 267 
<< pdiffusion >>
rect 466 266 467 267 
<< pdiffusion >>
rect 467 266 468 267 
<< pdiffusion >>
rect 480 266 481 267 
<< pdiffusion >>
rect 481 266 482 267 
<< pdiffusion >>
rect 482 266 483 267 
<< pdiffusion >>
rect 483 266 484 267 
<< pdiffusion >>
rect 484 266 485 267 
<< pdiffusion >>
rect 485 266 486 267 
<< pdiffusion >>
rect 498 266 499 267 
<< pdiffusion >>
rect 499 266 500 267 
<< pdiffusion >>
rect 500 266 501 267 
<< pdiffusion >>
rect 501 266 502 267 
<< pdiffusion >>
rect 502 266 503 267 
<< pdiffusion >>
rect 503 266 504 267 
<< pdiffusion >>
rect 516 266 517 267 
<< pdiffusion >>
rect 517 266 518 267 
<< pdiffusion >>
rect 518 266 519 267 
<< pdiffusion >>
rect 519 266 520 267 
<< pdiffusion >>
rect 520 266 521 267 
<< pdiffusion >>
rect 521 266 522 267 
<< m1 >>
rect 523 266 524 267 
<< pdiffusion >>
rect 12 267 13 268 
<< pdiffusion >>
rect 13 267 14 268 
<< pdiffusion >>
rect 14 267 15 268 
<< pdiffusion >>
rect 15 267 16 268 
<< pdiffusion >>
rect 16 267 17 268 
<< pdiffusion >>
rect 17 267 18 268 
<< m1 >>
rect 19 267 20 268 
<< m1 >>
rect 22 267 23 268 
<< m1 >>
rect 44 267 45 268 
<< pdiffusion >>
rect 48 267 49 268 
<< pdiffusion >>
rect 49 267 50 268 
<< pdiffusion >>
rect 50 267 51 268 
<< pdiffusion >>
rect 51 267 52 268 
<< pdiffusion >>
rect 52 267 53 268 
<< pdiffusion >>
rect 53 267 54 268 
<< m1 >>
rect 55 267 56 268 
<< m1 >>
rect 64 267 65 268 
<< pdiffusion >>
rect 66 267 67 268 
<< pdiffusion >>
rect 67 267 68 268 
<< pdiffusion >>
rect 68 267 69 268 
<< pdiffusion >>
rect 69 267 70 268 
<< pdiffusion >>
rect 70 267 71 268 
<< pdiffusion >>
rect 71 267 72 268 
<< pdiffusion >>
rect 84 267 85 268 
<< pdiffusion >>
rect 85 267 86 268 
<< pdiffusion >>
rect 86 267 87 268 
<< pdiffusion >>
rect 87 267 88 268 
<< pdiffusion >>
rect 88 267 89 268 
<< pdiffusion >>
rect 89 267 90 268 
<< m1 >>
rect 91 267 92 268 
<< m2 >>
rect 92 267 93 268 
<< pdiffusion >>
rect 102 267 103 268 
<< pdiffusion >>
rect 103 267 104 268 
<< pdiffusion >>
rect 104 267 105 268 
<< pdiffusion >>
rect 105 267 106 268 
<< pdiffusion >>
rect 106 267 107 268 
<< pdiffusion >>
rect 107 267 108 268 
<< m1 >>
rect 109 267 110 268 
<< pdiffusion >>
rect 120 267 121 268 
<< pdiffusion >>
rect 121 267 122 268 
<< pdiffusion >>
rect 122 267 123 268 
<< pdiffusion >>
rect 123 267 124 268 
<< pdiffusion >>
rect 124 267 125 268 
<< pdiffusion >>
rect 125 267 126 268 
<< pdiffusion >>
rect 138 267 139 268 
<< pdiffusion >>
rect 139 267 140 268 
<< pdiffusion >>
rect 140 267 141 268 
<< pdiffusion >>
rect 141 267 142 268 
<< pdiffusion >>
rect 142 267 143 268 
<< pdiffusion >>
rect 143 267 144 268 
<< m1 >>
rect 148 267 149 268 
<< pdiffusion >>
rect 156 267 157 268 
<< pdiffusion >>
rect 157 267 158 268 
<< pdiffusion >>
rect 158 267 159 268 
<< pdiffusion >>
rect 159 267 160 268 
<< pdiffusion >>
rect 160 267 161 268 
<< pdiffusion >>
rect 161 267 162 268 
<< m1 >>
rect 163 267 164 268 
<< pdiffusion >>
rect 174 267 175 268 
<< pdiffusion >>
rect 175 267 176 268 
<< pdiffusion >>
rect 176 267 177 268 
<< pdiffusion >>
rect 177 267 178 268 
<< pdiffusion >>
rect 178 267 179 268 
<< pdiffusion >>
rect 179 267 180 268 
<< m1 >>
rect 181 267 182 268 
<< m2 >>
rect 182 267 183 268 
<< m1 >>
rect 186 267 187 268 
<< m1 >>
rect 190 267 191 268 
<< pdiffusion >>
rect 192 267 193 268 
<< pdiffusion >>
rect 193 267 194 268 
<< pdiffusion >>
rect 194 267 195 268 
<< pdiffusion >>
rect 195 267 196 268 
<< pdiffusion >>
rect 196 267 197 268 
<< pdiffusion >>
rect 197 267 198 268 
<< m1 >>
rect 199 267 200 268 
<< pdiffusion >>
rect 210 267 211 268 
<< pdiffusion >>
rect 211 267 212 268 
<< pdiffusion >>
rect 212 267 213 268 
<< pdiffusion >>
rect 213 267 214 268 
<< pdiffusion >>
rect 214 267 215 268 
<< pdiffusion >>
rect 215 267 216 268 
<< m1 >>
rect 217 267 218 268 
<< m2 >>
rect 217 267 218 268 
<< m1 >>
rect 219 267 220 268 
<< pdiffusion >>
rect 228 267 229 268 
<< pdiffusion >>
rect 229 267 230 268 
<< pdiffusion >>
rect 230 267 231 268 
<< pdiffusion >>
rect 231 267 232 268 
<< pdiffusion >>
rect 232 267 233 268 
<< pdiffusion >>
rect 233 267 234 268 
<< m1 >>
rect 237 267 238 268 
<< m2 >>
rect 238 267 239 268 
<< pdiffusion >>
rect 246 267 247 268 
<< pdiffusion >>
rect 247 267 248 268 
<< pdiffusion >>
rect 248 267 249 268 
<< pdiffusion >>
rect 249 267 250 268 
<< pdiffusion >>
rect 250 267 251 268 
<< pdiffusion >>
rect 251 267 252 268 
<< m1 >>
rect 253 267 254 268 
<< m1 >>
rect 255 267 256 268 
<< m1 >>
rect 259 267 260 268 
<< m1 >>
rect 262 267 263 268 
<< m2 >>
rect 262 267 263 268 
<< pdiffusion >>
rect 264 267 265 268 
<< pdiffusion >>
rect 265 267 266 268 
<< pdiffusion >>
rect 266 267 267 268 
<< pdiffusion >>
rect 267 267 268 268 
<< pdiffusion >>
rect 268 267 269 268 
<< pdiffusion >>
rect 269 267 270 268 
<< m1 >>
rect 280 267 281 268 
<< pdiffusion >>
rect 282 267 283 268 
<< pdiffusion >>
rect 283 267 284 268 
<< pdiffusion >>
rect 284 267 285 268 
<< pdiffusion >>
rect 285 267 286 268 
<< pdiffusion >>
rect 286 267 287 268 
<< pdiffusion >>
rect 287 267 288 268 
<< m1 >>
rect 289 267 290 268 
<< m2 >>
rect 289 267 290 268 
<< pdiffusion >>
rect 300 267 301 268 
<< pdiffusion >>
rect 301 267 302 268 
<< pdiffusion >>
rect 302 267 303 268 
<< pdiffusion >>
rect 303 267 304 268 
<< pdiffusion >>
rect 304 267 305 268 
<< pdiffusion >>
rect 305 267 306 268 
<< m1 >>
rect 307 267 308 268 
<< m1 >>
rect 309 267 310 268 
<< m2 >>
rect 310 267 311 268 
<< pdiffusion >>
rect 318 267 319 268 
<< pdiffusion >>
rect 319 267 320 268 
<< pdiffusion >>
rect 320 267 321 268 
<< pdiffusion >>
rect 321 267 322 268 
<< pdiffusion >>
rect 322 267 323 268 
<< pdiffusion >>
rect 323 267 324 268 
<< pdiffusion >>
rect 336 267 337 268 
<< pdiffusion >>
rect 337 267 338 268 
<< pdiffusion >>
rect 338 267 339 268 
<< pdiffusion >>
rect 339 267 340 268 
<< pdiffusion >>
rect 340 267 341 268 
<< pdiffusion >>
rect 341 267 342 268 
<< m1 >>
rect 344 267 345 268 
<< m1 >>
rect 346 267 347 268 
<< pdiffusion >>
rect 354 267 355 268 
<< pdiffusion >>
rect 355 267 356 268 
<< pdiffusion >>
rect 356 267 357 268 
<< pdiffusion >>
rect 357 267 358 268 
<< pdiffusion >>
rect 358 267 359 268 
<< pdiffusion >>
rect 359 267 360 268 
<< m1 >>
rect 366 267 367 268 
<< m1 >>
rect 370 267 371 268 
<< pdiffusion >>
rect 372 267 373 268 
<< pdiffusion >>
rect 373 267 374 268 
<< pdiffusion >>
rect 374 267 375 268 
<< pdiffusion >>
rect 375 267 376 268 
<< pdiffusion >>
rect 376 267 377 268 
<< pdiffusion >>
rect 377 267 378 268 
<< m1 >>
rect 386 267 387 268 
<< m1 >>
rect 388 267 389 268 
<< pdiffusion >>
rect 390 267 391 268 
<< pdiffusion >>
rect 391 267 392 268 
<< pdiffusion >>
rect 392 267 393 268 
<< pdiffusion >>
rect 393 267 394 268 
<< pdiffusion >>
rect 394 267 395 268 
<< pdiffusion >>
rect 395 267 396 268 
<< m1 >>
rect 397 267 398 268 
<< pdiffusion >>
rect 408 267 409 268 
<< pdiffusion >>
rect 409 267 410 268 
<< pdiffusion >>
rect 410 267 411 268 
<< pdiffusion >>
rect 411 267 412 268 
<< pdiffusion >>
rect 412 267 413 268 
<< pdiffusion >>
rect 413 267 414 268 
<< m1 >>
rect 416 267 417 268 
<< m1 >>
rect 419 267 420 268 
<< m2 >>
rect 420 267 421 268 
<< pdiffusion >>
rect 426 267 427 268 
<< pdiffusion >>
rect 427 267 428 268 
<< pdiffusion >>
rect 428 267 429 268 
<< pdiffusion >>
rect 429 267 430 268 
<< pdiffusion >>
rect 430 267 431 268 
<< pdiffusion >>
rect 431 267 432 268 
<< m1 >>
rect 437 267 438 268 
<< m1 >>
rect 442 267 443 268 
<< pdiffusion >>
rect 444 267 445 268 
<< pdiffusion >>
rect 445 267 446 268 
<< pdiffusion >>
rect 446 267 447 268 
<< pdiffusion >>
rect 447 267 448 268 
<< pdiffusion >>
rect 448 267 449 268 
<< pdiffusion >>
rect 449 267 450 268 
<< pdiffusion >>
rect 462 267 463 268 
<< pdiffusion >>
rect 463 267 464 268 
<< pdiffusion >>
rect 464 267 465 268 
<< pdiffusion >>
rect 465 267 466 268 
<< pdiffusion >>
rect 466 267 467 268 
<< pdiffusion >>
rect 467 267 468 268 
<< pdiffusion >>
rect 480 267 481 268 
<< pdiffusion >>
rect 481 267 482 268 
<< pdiffusion >>
rect 482 267 483 268 
<< pdiffusion >>
rect 483 267 484 268 
<< pdiffusion >>
rect 484 267 485 268 
<< pdiffusion >>
rect 485 267 486 268 
<< pdiffusion >>
rect 498 267 499 268 
<< pdiffusion >>
rect 499 267 500 268 
<< pdiffusion >>
rect 500 267 501 268 
<< pdiffusion >>
rect 501 267 502 268 
<< pdiffusion >>
rect 502 267 503 268 
<< pdiffusion >>
rect 503 267 504 268 
<< pdiffusion >>
rect 516 267 517 268 
<< pdiffusion >>
rect 517 267 518 268 
<< pdiffusion >>
rect 518 267 519 268 
<< pdiffusion >>
rect 519 267 520 268 
<< pdiffusion >>
rect 520 267 521 268 
<< pdiffusion >>
rect 521 267 522 268 
<< m1 >>
rect 523 267 524 268 
<< pdiffusion >>
rect 12 268 13 269 
<< pdiffusion >>
rect 13 268 14 269 
<< pdiffusion >>
rect 14 268 15 269 
<< pdiffusion >>
rect 15 268 16 269 
<< pdiffusion >>
rect 16 268 17 269 
<< pdiffusion >>
rect 17 268 18 269 
<< m1 >>
rect 19 268 20 269 
<< m1 >>
rect 22 268 23 269 
<< m1 >>
rect 44 268 45 269 
<< pdiffusion >>
rect 48 268 49 269 
<< pdiffusion >>
rect 49 268 50 269 
<< pdiffusion >>
rect 50 268 51 269 
<< pdiffusion >>
rect 51 268 52 269 
<< pdiffusion >>
rect 52 268 53 269 
<< pdiffusion >>
rect 53 268 54 269 
<< m1 >>
rect 55 268 56 269 
<< m1 >>
rect 64 268 65 269 
<< pdiffusion >>
rect 66 268 67 269 
<< pdiffusion >>
rect 67 268 68 269 
<< pdiffusion >>
rect 68 268 69 269 
<< pdiffusion >>
rect 69 268 70 269 
<< pdiffusion >>
rect 70 268 71 269 
<< pdiffusion >>
rect 71 268 72 269 
<< pdiffusion >>
rect 84 268 85 269 
<< pdiffusion >>
rect 85 268 86 269 
<< pdiffusion >>
rect 86 268 87 269 
<< pdiffusion >>
rect 87 268 88 269 
<< pdiffusion >>
rect 88 268 89 269 
<< pdiffusion >>
rect 89 268 90 269 
<< m1 >>
rect 91 268 92 269 
<< m2 >>
rect 92 268 93 269 
<< pdiffusion >>
rect 102 268 103 269 
<< pdiffusion >>
rect 103 268 104 269 
<< pdiffusion >>
rect 104 268 105 269 
<< pdiffusion >>
rect 105 268 106 269 
<< pdiffusion >>
rect 106 268 107 269 
<< pdiffusion >>
rect 107 268 108 269 
<< m1 >>
rect 109 268 110 269 
<< pdiffusion >>
rect 120 268 121 269 
<< pdiffusion >>
rect 121 268 122 269 
<< pdiffusion >>
rect 122 268 123 269 
<< pdiffusion >>
rect 123 268 124 269 
<< pdiffusion >>
rect 124 268 125 269 
<< pdiffusion >>
rect 125 268 126 269 
<< pdiffusion >>
rect 138 268 139 269 
<< pdiffusion >>
rect 139 268 140 269 
<< pdiffusion >>
rect 140 268 141 269 
<< pdiffusion >>
rect 141 268 142 269 
<< pdiffusion >>
rect 142 268 143 269 
<< pdiffusion >>
rect 143 268 144 269 
<< m1 >>
rect 148 268 149 269 
<< pdiffusion >>
rect 156 268 157 269 
<< pdiffusion >>
rect 157 268 158 269 
<< pdiffusion >>
rect 158 268 159 269 
<< pdiffusion >>
rect 159 268 160 269 
<< pdiffusion >>
rect 160 268 161 269 
<< pdiffusion >>
rect 161 268 162 269 
<< m1 >>
rect 163 268 164 269 
<< pdiffusion >>
rect 174 268 175 269 
<< pdiffusion >>
rect 175 268 176 269 
<< pdiffusion >>
rect 176 268 177 269 
<< pdiffusion >>
rect 177 268 178 269 
<< pdiffusion >>
rect 178 268 179 269 
<< pdiffusion >>
rect 179 268 180 269 
<< m1 >>
rect 181 268 182 269 
<< m2 >>
rect 182 268 183 269 
<< m1 >>
rect 186 268 187 269 
<< m1 >>
rect 190 268 191 269 
<< pdiffusion >>
rect 192 268 193 269 
<< pdiffusion >>
rect 193 268 194 269 
<< pdiffusion >>
rect 194 268 195 269 
<< pdiffusion >>
rect 195 268 196 269 
<< pdiffusion >>
rect 196 268 197 269 
<< pdiffusion >>
rect 197 268 198 269 
<< m1 >>
rect 199 268 200 269 
<< pdiffusion >>
rect 210 268 211 269 
<< pdiffusion >>
rect 211 268 212 269 
<< pdiffusion >>
rect 212 268 213 269 
<< pdiffusion >>
rect 213 268 214 269 
<< pdiffusion >>
rect 214 268 215 269 
<< pdiffusion >>
rect 215 268 216 269 
<< m1 >>
rect 217 268 218 269 
<< m2 >>
rect 217 268 218 269 
<< m1 >>
rect 219 268 220 269 
<< pdiffusion >>
rect 228 268 229 269 
<< pdiffusion >>
rect 229 268 230 269 
<< pdiffusion >>
rect 230 268 231 269 
<< pdiffusion >>
rect 231 268 232 269 
<< pdiffusion >>
rect 232 268 233 269 
<< pdiffusion >>
rect 233 268 234 269 
<< m1 >>
rect 237 268 238 269 
<< m2 >>
rect 238 268 239 269 
<< pdiffusion >>
rect 246 268 247 269 
<< pdiffusion >>
rect 247 268 248 269 
<< pdiffusion >>
rect 248 268 249 269 
<< pdiffusion >>
rect 249 268 250 269 
<< pdiffusion >>
rect 250 268 251 269 
<< pdiffusion >>
rect 251 268 252 269 
<< m1 >>
rect 253 268 254 269 
<< m1 >>
rect 255 268 256 269 
<< m1 >>
rect 259 268 260 269 
<< m1 >>
rect 262 268 263 269 
<< m2 >>
rect 262 268 263 269 
<< pdiffusion >>
rect 264 268 265 269 
<< pdiffusion >>
rect 265 268 266 269 
<< pdiffusion >>
rect 266 268 267 269 
<< pdiffusion >>
rect 267 268 268 269 
<< pdiffusion >>
rect 268 268 269 269 
<< pdiffusion >>
rect 269 268 270 269 
<< m1 >>
rect 280 268 281 269 
<< pdiffusion >>
rect 282 268 283 269 
<< pdiffusion >>
rect 283 268 284 269 
<< pdiffusion >>
rect 284 268 285 269 
<< pdiffusion >>
rect 285 268 286 269 
<< pdiffusion >>
rect 286 268 287 269 
<< pdiffusion >>
rect 287 268 288 269 
<< m1 >>
rect 289 268 290 269 
<< m2 >>
rect 289 268 290 269 
<< pdiffusion >>
rect 300 268 301 269 
<< pdiffusion >>
rect 301 268 302 269 
<< pdiffusion >>
rect 302 268 303 269 
<< pdiffusion >>
rect 303 268 304 269 
<< pdiffusion >>
rect 304 268 305 269 
<< pdiffusion >>
rect 305 268 306 269 
<< m1 >>
rect 307 268 308 269 
<< m1 >>
rect 309 268 310 269 
<< m2 >>
rect 310 268 311 269 
<< pdiffusion >>
rect 318 268 319 269 
<< pdiffusion >>
rect 319 268 320 269 
<< pdiffusion >>
rect 320 268 321 269 
<< pdiffusion >>
rect 321 268 322 269 
<< pdiffusion >>
rect 322 268 323 269 
<< pdiffusion >>
rect 323 268 324 269 
<< pdiffusion >>
rect 336 268 337 269 
<< pdiffusion >>
rect 337 268 338 269 
<< pdiffusion >>
rect 338 268 339 269 
<< pdiffusion >>
rect 339 268 340 269 
<< pdiffusion >>
rect 340 268 341 269 
<< pdiffusion >>
rect 341 268 342 269 
<< m1 >>
rect 344 268 345 269 
<< m1 >>
rect 346 268 347 269 
<< pdiffusion >>
rect 354 268 355 269 
<< pdiffusion >>
rect 355 268 356 269 
<< pdiffusion >>
rect 356 268 357 269 
<< pdiffusion >>
rect 357 268 358 269 
<< pdiffusion >>
rect 358 268 359 269 
<< pdiffusion >>
rect 359 268 360 269 
<< m1 >>
rect 366 268 367 269 
<< m1 >>
rect 370 268 371 269 
<< pdiffusion >>
rect 372 268 373 269 
<< pdiffusion >>
rect 373 268 374 269 
<< pdiffusion >>
rect 374 268 375 269 
<< pdiffusion >>
rect 375 268 376 269 
<< pdiffusion >>
rect 376 268 377 269 
<< pdiffusion >>
rect 377 268 378 269 
<< m1 >>
rect 386 268 387 269 
<< m1 >>
rect 388 268 389 269 
<< pdiffusion >>
rect 390 268 391 269 
<< pdiffusion >>
rect 391 268 392 269 
<< pdiffusion >>
rect 392 268 393 269 
<< pdiffusion >>
rect 393 268 394 269 
<< pdiffusion >>
rect 394 268 395 269 
<< pdiffusion >>
rect 395 268 396 269 
<< m1 >>
rect 397 268 398 269 
<< pdiffusion >>
rect 408 268 409 269 
<< pdiffusion >>
rect 409 268 410 269 
<< pdiffusion >>
rect 410 268 411 269 
<< pdiffusion >>
rect 411 268 412 269 
<< pdiffusion >>
rect 412 268 413 269 
<< pdiffusion >>
rect 413 268 414 269 
<< m1 >>
rect 416 268 417 269 
<< m1 >>
rect 419 268 420 269 
<< m2 >>
rect 420 268 421 269 
<< pdiffusion >>
rect 426 268 427 269 
<< pdiffusion >>
rect 427 268 428 269 
<< pdiffusion >>
rect 428 268 429 269 
<< pdiffusion >>
rect 429 268 430 269 
<< pdiffusion >>
rect 430 268 431 269 
<< pdiffusion >>
rect 431 268 432 269 
<< m1 >>
rect 437 268 438 269 
<< m2 >>
rect 437 268 438 269 
<< m2c >>
rect 437 268 438 269 
<< m1 >>
rect 437 268 438 269 
<< m2 >>
rect 437 268 438 269 
<< m1 >>
rect 442 268 443 269 
<< pdiffusion >>
rect 444 268 445 269 
<< pdiffusion >>
rect 445 268 446 269 
<< pdiffusion >>
rect 446 268 447 269 
<< pdiffusion >>
rect 447 268 448 269 
<< pdiffusion >>
rect 448 268 449 269 
<< pdiffusion >>
rect 449 268 450 269 
<< pdiffusion >>
rect 462 268 463 269 
<< pdiffusion >>
rect 463 268 464 269 
<< pdiffusion >>
rect 464 268 465 269 
<< pdiffusion >>
rect 465 268 466 269 
<< pdiffusion >>
rect 466 268 467 269 
<< pdiffusion >>
rect 467 268 468 269 
<< pdiffusion >>
rect 480 268 481 269 
<< pdiffusion >>
rect 481 268 482 269 
<< pdiffusion >>
rect 482 268 483 269 
<< pdiffusion >>
rect 483 268 484 269 
<< pdiffusion >>
rect 484 268 485 269 
<< pdiffusion >>
rect 485 268 486 269 
<< pdiffusion >>
rect 498 268 499 269 
<< pdiffusion >>
rect 499 268 500 269 
<< pdiffusion >>
rect 500 268 501 269 
<< pdiffusion >>
rect 501 268 502 269 
<< pdiffusion >>
rect 502 268 503 269 
<< pdiffusion >>
rect 503 268 504 269 
<< pdiffusion >>
rect 516 268 517 269 
<< pdiffusion >>
rect 517 268 518 269 
<< pdiffusion >>
rect 518 268 519 269 
<< pdiffusion >>
rect 519 268 520 269 
<< pdiffusion >>
rect 520 268 521 269 
<< pdiffusion >>
rect 521 268 522 269 
<< m1 >>
rect 523 268 524 269 
<< pdiffusion >>
rect 12 269 13 270 
<< pdiffusion >>
rect 13 269 14 270 
<< pdiffusion >>
rect 14 269 15 270 
<< pdiffusion >>
rect 15 269 16 270 
<< pdiffusion >>
rect 16 269 17 270 
<< pdiffusion >>
rect 17 269 18 270 
<< m1 >>
rect 19 269 20 270 
<< m1 >>
rect 22 269 23 270 
<< m1 >>
rect 44 269 45 270 
<< pdiffusion >>
rect 48 269 49 270 
<< pdiffusion >>
rect 49 269 50 270 
<< pdiffusion >>
rect 50 269 51 270 
<< pdiffusion >>
rect 51 269 52 270 
<< pdiffusion >>
rect 52 269 53 270 
<< pdiffusion >>
rect 53 269 54 270 
<< m1 >>
rect 55 269 56 270 
<< m1 >>
rect 64 269 65 270 
<< pdiffusion >>
rect 66 269 67 270 
<< pdiffusion >>
rect 67 269 68 270 
<< pdiffusion >>
rect 68 269 69 270 
<< pdiffusion >>
rect 69 269 70 270 
<< pdiffusion >>
rect 70 269 71 270 
<< pdiffusion >>
rect 71 269 72 270 
<< pdiffusion >>
rect 84 269 85 270 
<< pdiffusion >>
rect 85 269 86 270 
<< pdiffusion >>
rect 86 269 87 270 
<< pdiffusion >>
rect 87 269 88 270 
<< pdiffusion >>
rect 88 269 89 270 
<< pdiffusion >>
rect 89 269 90 270 
<< m1 >>
rect 91 269 92 270 
<< m2 >>
rect 92 269 93 270 
<< pdiffusion >>
rect 102 269 103 270 
<< pdiffusion >>
rect 103 269 104 270 
<< pdiffusion >>
rect 104 269 105 270 
<< pdiffusion >>
rect 105 269 106 270 
<< pdiffusion >>
rect 106 269 107 270 
<< pdiffusion >>
rect 107 269 108 270 
<< m1 >>
rect 109 269 110 270 
<< pdiffusion >>
rect 120 269 121 270 
<< pdiffusion >>
rect 121 269 122 270 
<< pdiffusion >>
rect 122 269 123 270 
<< pdiffusion >>
rect 123 269 124 270 
<< pdiffusion >>
rect 124 269 125 270 
<< pdiffusion >>
rect 125 269 126 270 
<< pdiffusion >>
rect 138 269 139 270 
<< pdiffusion >>
rect 139 269 140 270 
<< pdiffusion >>
rect 140 269 141 270 
<< pdiffusion >>
rect 141 269 142 270 
<< pdiffusion >>
rect 142 269 143 270 
<< pdiffusion >>
rect 143 269 144 270 
<< m1 >>
rect 148 269 149 270 
<< pdiffusion >>
rect 156 269 157 270 
<< pdiffusion >>
rect 157 269 158 270 
<< pdiffusion >>
rect 158 269 159 270 
<< pdiffusion >>
rect 159 269 160 270 
<< pdiffusion >>
rect 160 269 161 270 
<< pdiffusion >>
rect 161 269 162 270 
<< m1 >>
rect 163 269 164 270 
<< pdiffusion >>
rect 174 269 175 270 
<< pdiffusion >>
rect 175 269 176 270 
<< pdiffusion >>
rect 176 269 177 270 
<< pdiffusion >>
rect 177 269 178 270 
<< pdiffusion >>
rect 178 269 179 270 
<< pdiffusion >>
rect 179 269 180 270 
<< m1 >>
rect 181 269 182 270 
<< m2 >>
rect 182 269 183 270 
<< m1 >>
rect 186 269 187 270 
<< m1 >>
rect 190 269 191 270 
<< pdiffusion >>
rect 192 269 193 270 
<< pdiffusion >>
rect 193 269 194 270 
<< pdiffusion >>
rect 194 269 195 270 
<< pdiffusion >>
rect 195 269 196 270 
<< pdiffusion >>
rect 196 269 197 270 
<< pdiffusion >>
rect 197 269 198 270 
<< m1 >>
rect 199 269 200 270 
<< pdiffusion >>
rect 210 269 211 270 
<< pdiffusion >>
rect 211 269 212 270 
<< pdiffusion >>
rect 212 269 213 270 
<< pdiffusion >>
rect 213 269 214 270 
<< pdiffusion >>
rect 214 269 215 270 
<< pdiffusion >>
rect 215 269 216 270 
<< m1 >>
rect 217 269 218 270 
<< m2 >>
rect 217 269 218 270 
<< m1 >>
rect 219 269 220 270 
<< pdiffusion >>
rect 228 269 229 270 
<< pdiffusion >>
rect 229 269 230 270 
<< pdiffusion >>
rect 230 269 231 270 
<< m1 >>
rect 231 269 232 270 
<< m2 >>
rect 231 269 232 270 
<< m2c >>
rect 231 269 232 270 
<< m1 >>
rect 231 269 232 270 
<< m2 >>
rect 231 269 232 270 
<< pdiffusion >>
rect 231 269 232 270 
<< m1 >>
rect 232 269 233 270 
<< pdiffusion >>
rect 232 269 233 270 
<< pdiffusion >>
rect 233 269 234 270 
<< m1 >>
rect 237 269 238 270 
<< m2 >>
rect 238 269 239 270 
<< pdiffusion >>
rect 246 269 247 270 
<< m1 >>
rect 247 269 248 270 
<< pdiffusion >>
rect 247 269 248 270 
<< pdiffusion >>
rect 248 269 249 270 
<< pdiffusion >>
rect 249 269 250 270 
<< pdiffusion >>
rect 250 269 251 270 
<< pdiffusion >>
rect 251 269 252 270 
<< m1 >>
rect 253 269 254 270 
<< m1 >>
rect 255 269 256 270 
<< m1 >>
rect 259 269 260 270 
<< m1 >>
rect 262 269 263 270 
<< m2 >>
rect 262 269 263 270 
<< pdiffusion >>
rect 264 269 265 270 
<< pdiffusion >>
rect 265 269 266 270 
<< pdiffusion >>
rect 266 269 267 270 
<< pdiffusion >>
rect 267 269 268 270 
<< m1 >>
rect 268 269 269 270 
<< pdiffusion >>
rect 268 269 269 270 
<< pdiffusion >>
rect 269 269 270 270 
<< m1 >>
rect 280 269 281 270 
<< pdiffusion >>
rect 282 269 283 270 
<< pdiffusion >>
rect 283 269 284 270 
<< pdiffusion >>
rect 284 269 285 270 
<< pdiffusion >>
rect 285 269 286 270 
<< m1 >>
rect 286 269 287 270 
<< pdiffusion >>
rect 286 269 287 270 
<< pdiffusion >>
rect 287 269 288 270 
<< m1 >>
rect 289 269 290 270 
<< m2 >>
rect 289 269 290 270 
<< pdiffusion >>
rect 300 269 301 270 
<< pdiffusion >>
rect 301 269 302 270 
<< pdiffusion >>
rect 302 269 303 270 
<< pdiffusion >>
rect 303 269 304 270 
<< pdiffusion >>
rect 304 269 305 270 
<< pdiffusion >>
rect 305 269 306 270 
<< m1 >>
rect 307 269 308 270 
<< m1 >>
rect 309 269 310 270 
<< m2 >>
rect 310 269 311 270 
<< pdiffusion >>
rect 318 269 319 270 
<< pdiffusion >>
rect 319 269 320 270 
<< pdiffusion >>
rect 320 269 321 270 
<< pdiffusion >>
rect 321 269 322 270 
<< m1 >>
rect 322 269 323 270 
<< pdiffusion >>
rect 322 269 323 270 
<< pdiffusion >>
rect 323 269 324 270 
<< pdiffusion >>
rect 336 269 337 270 
<< pdiffusion >>
rect 337 269 338 270 
<< pdiffusion >>
rect 338 269 339 270 
<< pdiffusion >>
rect 339 269 340 270 
<< m1 >>
rect 340 269 341 270 
<< pdiffusion >>
rect 340 269 341 270 
<< pdiffusion >>
rect 341 269 342 270 
<< m1 >>
rect 344 269 345 270 
<< m1 >>
rect 346 269 347 270 
<< pdiffusion >>
rect 354 269 355 270 
<< pdiffusion >>
rect 355 269 356 270 
<< pdiffusion >>
rect 356 269 357 270 
<< pdiffusion >>
rect 357 269 358 270 
<< pdiffusion >>
rect 358 269 359 270 
<< pdiffusion >>
rect 359 269 360 270 
<< m1 >>
rect 366 269 367 270 
<< m1 >>
rect 370 269 371 270 
<< pdiffusion >>
rect 372 269 373 270 
<< pdiffusion >>
rect 373 269 374 270 
<< pdiffusion >>
rect 374 269 375 270 
<< pdiffusion >>
rect 375 269 376 270 
<< pdiffusion >>
rect 376 269 377 270 
<< pdiffusion >>
rect 377 269 378 270 
<< m1 >>
rect 386 269 387 270 
<< m1 >>
rect 388 269 389 270 
<< pdiffusion >>
rect 390 269 391 270 
<< m1 >>
rect 391 269 392 270 
<< pdiffusion >>
rect 391 269 392 270 
<< pdiffusion >>
rect 392 269 393 270 
<< pdiffusion >>
rect 393 269 394 270 
<< pdiffusion >>
rect 394 269 395 270 
<< pdiffusion >>
rect 395 269 396 270 
<< m1 >>
rect 397 269 398 270 
<< pdiffusion >>
rect 408 269 409 270 
<< pdiffusion >>
rect 409 269 410 270 
<< pdiffusion >>
rect 410 269 411 270 
<< pdiffusion >>
rect 411 269 412 270 
<< pdiffusion >>
rect 412 269 413 270 
<< pdiffusion >>
rect 413 269 414 270 
<< m1 >>
rect 416 269 417 270 
<< m1 >>
rect 419 269 420 270 
<< m2 >>
rect 420 269 421 270 
<< pdiffusion >>
rect 426 269 427 270 
<< pdiffusion >>
rect 427 269 428 270 
<< pdiffusion >>
rect 428 269 429 270 
<< pdiffusion >>
rect 429 269 430 270 
<< m1 >>
rect 430 269 431 270 
<< pdiffusion >>
rect 430 269 431 270 
<< pdiffusion >>
rect 431 269 432 270 
<< m2 >>
rect 437 269 438 270 
<< m1 >>
rect 442 269 443 270 
<< pdiffusion >>
rect 444 269 445 270 
<< pdiffusion >>
rect 445 269 446 270 
<< pdiffusion >>
rect 446 269 447 270 
<< pdiffusion >>
rect 447 269 448 270 
<< pdiffusion >>
rect 448 269 449 270 
<< pdiffusion >>
rect 449 269 450 270 
<< pdiffusion >>
rect 462 269 463 270 
<< pdiffusion >>
rect 463 269 464 270 
<< pdiffusion >>
rect 464 269 465 270 
<< pdiffusion >>
rect 465 269 466 270 
<< pdiffusion >>
rect 466 269 467 270 
<< pdiffusion >>
rect 467 269 468 270 
<< pdiffusion >>
rect 480 269 481 270 
<< pdiffusion >>
rect 481 269 482 270 
<< pdiffusion >>
rect 482 269 483 270 
<< pdiffusion >>
rect 483 269 484 270 
<< pdiffusion >>
rect 484 269 485 270 
<< pdiffusion >>
rect 485 269 486 270 
<< pdiffusion >>
rect 498 269 499 270 
<< pdiffusion >>
rect 499 269 500 270 
<< pdiffusion >>
rect 500 269 501 270 
<< pdiffusion >>
rect 501 269 502 270 
<< pdiffusion >>
rect 502 269 503 270 
<< pdiffusion >>
rect 503 269 504 270 
<< pdiffusion >>
rect 516 269 517 270 
<< pdiffusion >>
rect 517 269 518 270 
<< pdiffusion >>
rect 518 269 519 270 
<< pdiffusion >>
rect 519 269 520 270 
<< pdiffusion >>
rect 520 269 521 270 
<< pdiffusion >>
rect 521 269 522 270 
<< m1 >>
rect 523 269 524 270 
<< m1 >>
rect 19 270 20 271 
<< m1 >>
rect 22 270 23 271 
<< m1 >>
rect 44 270 45 271 
<< m1 >>
rect 55 270 56 271 
<< m1 >>
rect 64 270 65 271 
<< m1 >>
rect 91 270 92 271 
<< m2 >>
rect 92 270 93 271 
<< m1 >>
rect 109 270 110 271 
<< m1 >>
rect 148 270 149 271 
<< m1 >>
rect 163 270 164 271 
<< m1 >>
rect 181 270 182 271 
<< m2 >>
rect 182 270 183 271 
<< m1 >>
rect 186 270 187 271 
<< m1 >>
rect 190 270 191 271 
<< m1 >>
rect 199 270 200 271 
<< m1 >>
rect 217 270 218 271 
<< m2 >>
rect 217 270 218 271 
<< m1 >>
rect 219 270 220 271 
<< m1 >>
rect 232 270 233 271 
<< m2 >>
rect 232 270 233 271 
<< m1 >>
rect 237 270 238 271 
<< m2 >>
rect 238 270 239 271 
<< m1 >>
rect 247 270 248 271 
<< m1 >>
rect 253 270 254 271 
<< m2 >>
rect 253 270 254 271 
<< m2c >>
rect 253 270 254 271 
<< m1 >>
rect 253 270 254 271 
<< m2 >>
rect 253 270 254 271 
<< m1 >>
rect 255 270 256 271 
<< m2 >>
rect 255 270 256 271 
<< m2c >>
rect 255 270 256 271 
<< m1 >>
rect 255 270 256 271 
<< m2 >>
rect 255 270 256 271 
<< m1 >>
rect 259 270 260 271 
<< m2 >>
rect 259 270 260 271 
<< m2c >>
rect 259 270 260 271 
<< m1 >>
rect 259 270 260 271 
<< m2 >>
rect 259 270 260 271 
<< m1 >>
rect 262 270 263 271 
<< m2 >>
rect 262 270 263 271 
<< m1 >>
rect 268 270 269 271 
<< m1 >>
rect 280 270 281 271 
<< m1 >>
rect 286 270 287 271 
<< m1 >>
rect 289 270 290 271 
<< m2 >>
rect 289 270 290 271 
<< m1 >>
rect 307 270 308 271 
<< m1 >>
rect 309 270 310 271 
<< m2 >>
rect 310 270 311 271 
<< m1 >>
rect 322 270 323 271 
<< m1 >>
rect 340 270 341 271 
<< m1 >>
rect 344 270 345 271 
<< m1 >>
rect 346 270 347 271 
<< m1 >>
rect 366 270 367 271 
<< m1 >>
rect 370 270 371 271 
<< m1 >>
rect 386 270 387 271 
<< m1 >>
rect 388 270 389 271 
<< m1 >>
rect 391 270 392 271 
<< m1 >>
rect 397 270 398 271 
<< m1 >>
rect 416 270 417 271 
<< m1 >>
rect 419 270 420 271 
<< m2 >>
rect 420 270 421 271 
<< m1 >>
rect 430 270 431 271 
<< m2 >>
rect 434 270 435 271 
<< m1 >>
rect 435 270 436 271 
<< m2 >>
rect 435 270 436 271 
<< m2c >>
rect 435 270 436 271 
<< m1 >>
rect 435 270 436 271 
<< m2 >>
rect 435 270 436 271 
<< m1 >>
rect 436 270 437 271 
<< m1 >>
rect 437 270 438 271 
<< m2 >>
rect 437 270 438 271 
<< m1 >>
rect 438 270 439 271 
<< m1 >>
rect 439 270 440 271 
<< m1 >>
rect 440 270 441 271 
<< m1 >>
rect 441 270 442 271 
<< m1 >>
rect 442 270 443 271 
<< m1 >>
rect 523 270 524 271 
<< m1 >>
rect 19 271 20 272 
<< m1 >>
rect 22 271 23 272 
<< m1 >>
rect 44 271 45 272 
<< m1 >>
rect 55 271 56 272 
<< m1 >>
rect 64 271 65 272 
<< m1 >>
rect 89 271 90 272 
<< m2 >>
rect 89 271 90 272 
<< m2c >>
rect 89 271 90 272 
<< m1 >>
rect 89 271 90 272 
<< m2 >>
rect 89 271 90 272 
<< m2 >>
rect 90 271 91 272 
<< m1 >>
rect 91 271 92 272 
<< m2 >>
rect 91 271 92 272 
<< m2 >>
rect 92 271 93 272 
<< m1 >>
rect 109 271 110 272 
<< m1 >>
rect 148 271 149 272 
<< m1 >>
rect 163 271 164 272 
<< m1 >>
rect 181 271 182 272 
<< m2 >>
rect 182 271 183 272 
<< m1 >>
rect 186 271 187 272 
<< m1 >>
rect 190 271 191 272 
<< m1 >>
rect 199 271 200 272 
<< m1 >>
rect 215 271 216 272 
<< m2 >>
rect 215 271 216 272 
<< m2c >>
rect 215 271 216 272 
<< m1 >>
rect 215 271 216 272 
<< m2 >>
rect 215 271 216 272 
<< m2 >>
rect 216 271 217 272 
<< m1 >>
rect 217 271 218 272 
<< m2 >>
rect 217 271 218 272 
<< m1 >>
rect 219 271 220 272 
<< m2 >>
rect 232 271 233 272 
<< m1 >>
rect 237 271 238 272 
<< m2 >>
rect 238 271 239 272 
<< m1 >>
rect 247 271 248 272 
<< m2 >>
rect 253 271 254 272 
<< m2 >>
rect 255 271 256 272 
<< m2 >>
rect 259 271 260 272 
<< m1 >>
rect 262 271 263 272 
<< m2 >>
rect 262 271 263 272 
<< m1 >>
rect 268 271 269 272 
<< m1 >>
rect 269 271 270 272 
<< m1 >>
rect 270 271 271 272 
<< m2 >>
rect 270 271 271 272 
<< m1 >>
rect 271 271 272 272 
<< m2 >>
rect 271 271 272 272 
<< m1 >>
rect 272 271 273 272 
<< m2 >>
rect 272 271 273 272 
<< m1 >>
rect 273 271 274 272 
<< m2 >>
rect 273 271 274 272 
<< m1 >>
rect 274 271 275 272 
<< m2 >>
rect 274 271 275 272 
<< m1 >>
rect 275 271 276 272 
<< m2 >>
rect 275 271 276 272 
<< m1 >>
rect 276 271 277 272 
<< m2 >>
rect 276 271 277 272 
<< m1 >>
rect 277 271 278 272 
<< m1 >>
rect 278 271 279 272 
<< m2 >>
rect 278 271 279 272 
<< m2c >>
rect 278 271 279 272 
<< m1 >>
rect 278 271 279 272 
<< m2 >>
rect 278 271 279 272 
<< m2 >>
rect 279 271 280 272 
<< m1 >>
rect 280 271 281 272 
<< m2 >>
rect 280 271 281 272 
<< m1 >>
rect 286 271 287 272 
<< m1 >>
rect 289 271 290 272 
<< m2 >>
rect 289 271 290 272 
<< m1 >>
rect 307 271 308 272 
<< m1 >>
rect 309 271 310 272 
<< m2 >>
rect 310 271 311 272 
<< m1 >>
rect 322 271 323 272 
<< m1 >>
rect 340 271 341 272 
<< m1 >>
rect 344 271 345 272 
<< m1 >>
rect 346 271 347 272 
<< m1 >>
rect 366 271 367 272 
<< m1 >>
rect 370 271 371 272 
<< m1 >>
rect 386 271 387 272 
<< m1 >>
rect 388 271 389 272 
<< m1 >>
rect 391 271 392 272 
<< m1 >>
rect 397 271 398 272 
<< m1 >>
rect 416 271 417 272 
<< m1 >>
rect 419 271 420 272 
<< m2 >>
rect 420 271 421 272 
<< m1 >>
rect 430 271 431 272 
<< m1 >>
rect 431 271 432 272 
<< m1 >>
rect 432 271 433 272 
<< m1 >>
rect 433 271 434 272 
<< m2 >>
rect 434 271 435 272 
<< m2 >>
rect 437 271 438 272 
<< m1 >>
rect 523 271 524 272 
<< m1 >>
rect 19 272 20 273 
<< m1 >>
rect 22 272 23 273 
<< m1 >>
rect 44 272 45 273 
<< m1 >>
rect 55 272 56 273 
<< m1 >>
rect 64 272 65 273 
<< m1 >>
rect 89 272 90 273 
<< m1 >>
rect 91 272 92 273 
<< m1 >>
rect 109 272 110 273 
<< m1 >>
rect 148 272 149 273 
<< m1 >>
rect 163 272 164 273 
<< m2 >>
rect 163 272 164 273 
<< m2c >>
rect 163 272 164 273 
<< m1 >>
rect 163 272 164 273 
<< m2 >>
rect 163 272 164 273 
<< m1 >>
rect 176 272 177 273 
<< m2 >>
rect 176 272 177 273 
<< m2c >>
rect 176 272 177 273 
<< m1 >>
rect 176 272 177 273 
<< m2 >>
rect 176 272 177 273 
<< m2 >>
rect 177 272 178 273 
<< m1 >>
rect 178 272 179 273 
<< m2 >>
rect 178 272 179 273 
<< m1 >>
rect 179 272 180 273 
<< m2 >>
rect 179 272 180 273 
<< m1 >>
rect 180 272 181 273 
<< m2 >>
rect 180 272 181 273 
<< m1 >>
rect 181 272 182 273 
<< m2 >>
rect 181 272 182 273 
<< m2 >>
rect 182 272 183 273 
<< m1 >>
rect 186 272 187 273 
<< m2 >>
rect 186 272 187 273 
<< m2c >>
rect 186 272 187 273 
<< m1 >>
rect 186 272 187 273 
<< m2 >>
rect 186 272 187 273 
<< m1 >>
rect 190 272 191 273 
<< m1 >>
rect 199 272 200 273 
<< m1 >>
rect 215 272 216 273 
<< m1 >>
rect 217 272 218 273 
<< m1 >>
rect 219 272 220 273 
<< m2 >>
rect 219 272 220 273 
<< m2c >>
rect 219 272 220 273 
<< m1 >>
rect 219 272 220 273 
<< m2 >>
rect 219 272 220 273 
<< m1 >>
rect 230 272 231 273 
<< m2 >>
rect 230 272 231 273 
<< m2c >>
rect 230 272 231 273 
<< m1 >>
rect 230 272 231 273 
<< m2 >>
rect 230 272 231 273 
<< m1 >>
rect 231 272 232 273 
<< m1 >>
rect 232 272 233 273 
<< m2 >>
rect 232 272 233 273 
<< m1 >>
rect 233 272 234 273 
<< m1 >>
rect 234 272 235 273 
<< m1 >>
rect 235 272 236 273 
<< m1 >>
rect 236 272 237 273 
<< m1 >>
rect 237 272 238 273 
<< m2 >>
rect 238 272 239 273 
<< m1 >>
rect 247 272 248 273 
<< m1 >>
rect 248 272 249 273 
<< m1 >>
rect 249 272 250 273 
<< m1 >>
rect 250 272 251 273 
<< m1 >>
rect 251 272 252 273 
<< m1 >>
rect 252 272 253 273 
<< m1 >>
rect 253 272 254 273 
<< m2 >>
rect 253 272 254 273 
<< m1 >>
rect 254 272 255 273 
<< m1 >>
rect 255 272 256 273 
<< m2 >>
rect 255 272 256 273 
<< m1 >>
rect 256 272 257 273 
<< m1 >>
rect 257 272 258 273 
<< m1 >>
rect 258 272 259 273 
<< m1 >>
rect 259 272 260 273 
<< m2 >>
rect 259 272 260 273 
<< m1 >>
rect 260 272 261 273 
<< m1 >>
rect 261 272 262 273 
<< m1 >>
rect 262 272 263 273 
<< m2 >>
rect 262 272 263 273 
<< m2 >>
rect 270 272 271 273 
<< m2 >>
rect 276 272 277 273 
<< m1 >>
rect 280 272 281 273 
<< m2 >>
rect 280 272 281 273 
<< m1 >>
rect 286 272 287 273 
<< m1 >>
rect 289 272 290 273 
<< m2 >>
rect 289 272 290 273 
<< m1 >>
rect 307 272 308 273 
<< m1 >>
rect 309 272 310 273 
<< m2 >>
rect 310 272 311 273 
<< m1 >>
rect 322 272 323 273 
<< m1 >>
rect 340 272 341 273 
<< m1 >>
rect 344 272 345 273 
<< m2 >>
rect 344 272 345 273 
<< m2c >>
rect 344 272 345 273 
<< m1 >>
rect 344 272 345 273 
<< m2 >>
rect 344 272 345 273 
<< m1 >>
rect 346 272 347 273 
<< m2 >>
rect 346 272 347 273 
<< m2c >>
rect 346 272 347 273 
<< m1 >>
rect 346 272 347 273 
<< m2 >>
rect 346 272 347 273 
<< m1 >>
rect 366 272 367 273 
<< m2 >>
rect 366 272 367 273 
<< m2c >>
rect 366 272 367 273 
<< m1 >>
rect 366 272 367 273 
<< m2 >>
rect 366 272 367 273 
<< m1 >>
rect 370 272 371 273 
<< m1 >>
rect 386 272 387 273 
<< m1 >>
rect 388 272 389 273 
<< m1 >>
rect 391 272 392 273 
<< m1 >>
rect 392 272 393 273 
<< m1 >>
rect 393 272 394 273 
<< m1 >>
rect 394 272 395 273 
<< m1 >>
rect 395 272 396 273 
<< m1 >>
rect 396 272 397 273 
<< m1 >>
rect 397 272 398 273 
<< m1 >>
rect 416 272 417 273 
<< m1 >>
rect 419 272 420 273 
<< m2 >>
rect 420 272 421 273 
<< m1 >>
rect 433 272 434 273 
<< m2 >>
rect 434 272 435 273 
<< m1 >>
rect 437 272 438 273 
<< m2 >>
rect 437 272 438 273 
<< m2c >>
rect 437 272 438 273 
<< m1 >>
rect 437 272 438 273 
<< m2 >>
rect 437 272 438 273 
<< m1 >>
rect 523 272 524 273 
<< m1 >>
rect 19 273 20 274 
<< m1 >>
rect 22 273 23 274 
<< m1 >>
rect 44 273 45 274 
<< m1 >>
rect 55 273 56 274 
<< m1 >>
rect 64 273 65 274 
<< m1 >>
rect 89 273 90 274 
<< m1 >>
rect 91 273 92 274 
<< m1 >>
rect 109 273 110 274 
<< m1 >>
rect 148 273 149 274 
<< m2 >>
rect 163 273 164 274 
<< m1 >>
rect 176 273 177 274 
<< m1 >>
rect 178 273 179 274 
<< m2 >>
rect 186 273 187 274 
<< m1 >>
rect 190 273 191 274 
<< m1 >>
rect 199 273 200 274 
<< m2 >>
rect 214 273 215 274 
<< m1 >>
rect 215 273 216 274 
<< m2 >>
rect 215 273 216 274 
<< m2 >>
rect 216 273 217 274 
<< m1 >>
rect 217 273 218 274 
<< m2 >>
rect 217 273 218 274 
<< m2 >>
rect 218 273 219 274 
<< m2 >>
rect 219 273 220 274 
<< m2 >>
rect 230 273 231 274 
<< m2 >>
rect 232 273 233 274 
<< m2 >>
rect 238 273 239 274 
<< m2 >>
rect 253 273 254 274 
<< m2 >>
rect 255 273 256 274 
<< m2 >>
rect 259 273 260 274 
<< m2 >>
rect 262 273 263 274 
<< m2 >>
rect 270 273 271 274 
<< m2 >>
rect 272 273 273 274 
<< m1 >>
rect 273 273 274 274 
<< m2 >>
rect 273 273 274 274 
<< m2c >>
rect 273 273 274 274 
<< m1 >>
rect 273 273 274 274 
<< m2 >>
rect 273 273 274 274 
<< m1 >>
rect 274 273 275 274 
<< m1 >>
rect 275 273 276 274 
<< m1 >>
rect 276 273 277 274 
<< m2 >>
rect 276 273 277 274 
<< m1 >>
rect 277 273 278 274 
<< m1 >>
rect 278 273 279 274 
<< m1 >>
rect 279 273 280 274 
<< m1 >>
rect 280 273 281 274 
<< m2 >>
rect 280 273 281 274 
<< m1 >>
rect 286 273 287 274 
<< m1 >>
rect 289 273 290 274 
<< m2 >>
rect 289 273 290 274 
<< m1 >>
rect 307 273 308 274 
<< m1 >>
rect 309 273 310 274 
<< m2 >>
rect 310 273 311 274 
<< m1 >>
rect 322 273 323 274 
<< m1 >>
rect 340 273 341 274 
<< m2 >>
rect 344 273 345 274 
<< m2 >>
rect 346 273 347 274 
<< m2 >>
rect 366 273 367 274 
<< m1 >>
rect 370 273 371 274 
<< m2 >>
rect 380 273 381 274 
<< m1 >>
rect 381 273 382 274 
<< m2 >>
rect 381 273 382 274 
<< m2c >>
rect 381 273 382 274 
<< m1 >>
rect 381 273 382 274 
<< m2 >>
rect 381 273 382 274 
<< m1 >>
rect 382 273 383 274 
<< m1 >>
rect 383 273 384 274 
<< m1 >>
rect 384 273 385 274 
<< m1 >>
rect 385 273 386 274 
<< m1 >>
rect 386 273 387 274 
<< m1 >>
rect 388 273 389 274 
<< m1 >>
rect 416 273 417 274 
<< m1 >>
rect 419 273 420 274 
<< m2 >>
rect 420 273 421 274 
<< m1 >>
rect 431 273 432 274 
<< m2 >>
rect 431 273 432 274 
<< m2c >>
rect 431 273 432 274 
<< m1 >>
rect 431 273 432 274 
<< m2 >>
rect 431 273 432 274 
<< m2 >>
rect 432 273 433 274 
<< m1 >>
rect 433 273 434 274 
<< m2 >>
rect 433 273 434 274 
<< m2 >>
rect 434 273 435 274 
<< m1 >>
rect 437 273 438 274 
<< m1 >>
rect 523 273 524 274 
<< m1 >>
rect 19 274 20 275 
<< m1 >>
rect 22 274 23 275 
<< m1 >>
rect 44 274 45 275 
<< m1 >>
rect 55 274 56 275 
<< m1 >>
rect 64 274 65 275 
<< m1 >>
rect 89 274 90 275 
<< m1 >>
rect 91 274 92 275 
<< m1 >>
rect 109 274 110 275 
<< m1 >>
rect 148 274 149 275 
<< m2 >>
rect 149 274 150 275 
<< m1 >>
rect 150 274 151 275 
<< m2 >>
rect 150 274 151 275 
<< m2c >>
rect 150 274 151 275 
<< m1 >>
rect 150 274 151 275 
<< m2 >>
rect 150 274 151 275 
<< m1 >>
rect 151 274 152 275 
<< m1 >>
rect 152 274 153 275 
<< m1 >>
rect 153 274 154 275 
<< m1 >>
rect 154 274 155 275 
<< m2 >>
rect 154 274 155 275 
<< m2c >>
rect 154 274 155 275 
<< m1 >>
rect 154 274 155 275 
<< m2 >>
rect 154 274 155 275 
<< m2 >>
rect 155 274 156 275 
<< m1 >>
rect 156 274 157 275 
<< m2 >>
rect 156 274 157 275 
<< m1 >>
rect 157 274 158 275 
<< m2 >>
rect 157 274 158 275 
<< m1 >>
rect 158 274 159 275 
<< m2 >>
rect 158 274 159 275 
<< m1 >>
rect 159 274 160 275 
<< m2 >>
rect 159 274 160 275 
<< m1 >>
rect 160 274 161 275 
<< m2 >>
rect 160 274 161 275 
<< m1 >>
rect 161 274 162 275 
<< m2 >>
rect 161 274 162 275 
<< m1 >>
rect 162 274 163 275 
<< m2 >>
rect 162 274 163 275 
<< m1 >>
rect 163 274 164 275 
<< m2 >>
rect 163 274 164 275 
<< m1 >>
rect 164 274 165 275 
<< m1 >>
rect 165 274 166 275 
<< m1 >>
rect 166 274 167 275 
<< m1 >>
rect 167 274 168 275 
<< m1 >>
rect 168 274 169 275 
<< m1 >>
rect 169 274 170 275 
<< m1 >>
rect 170 274 171 275 
<< m1 >>
rect 171 274 172 275 
<< m1 >>
rect 172 274 173 275 
<< m1 >>
rect 173 274 174 275 
<< m1 >>
rect 174 274 175 275 
<< m1 >>
rect 175 274 176 275 
<< m1 >>
rect 176 274 177 275 
<< m1 >>
rect 178 274 179 275 
<< m2 >>
rect 179 274 180 275 
<< m1 >>
rect 180 274 181 275 
<< m2 >>
rect 180 274 181 275 
<< m2c >>
rect 180 274 181 275 
<< m1 >>
rect 180 274 181 275 
<< m2 >>
rect 180 274 181 275 
<< m1 >>
rect 181 274 182 275 
<< m1 >>
rect 182 274 183 275 
<< m1 >>
rect 183 274 184 275 
<< m1 >>
rect 184 274 185 275 
<< m1 >>
rect 185 274 186 275 
<< m1 >>
rect 186 274 187 275 
<< m2 >>
rect 186 274 187 275 
<< m1 >>
rect 187 274 188 275 
<< m1 >>
rect 188 274 189 275 
<< m1 >>
rect 189 274 190 275 
<< m1 >>
rect 190 274 191 275 
<< m1 >>
rect 199 274 200 275 
<< m1 >>
rect 200 274 201 275 
<< m1 >>
rect 201 274 202 275 
<< m1 >>
rect 202 274 203 275 
<< m1 >>
rect 203 274 204 275 
<< m1 >>
rect 204 274 205 275 
<< m1 >>
rect 205 274 206 275 
<< m1 >>
rect 206 274 207 275 
<< m1 >>
rect 207 274 208 275 
<< m1 >>
rect 208 274 209 275 
<< m1 >>
rect 209 274 210 275 
<< m1 >>
rect 210 274 211 275 
<< m1 >>
rect 211 274 212 275 
<< m1 >>
rect 212 274 213 275 
<< m1 >>
rect 213 274 214 275 
<< m2 >>
rect 213 274 214 275 
<< m2c >>
rect 213 274 214 275 
<< m1 >>
rect 213 274 214 275 
<< m2 >>
rect 213 274 214 275 
<< m2 >>
rect 214 274 215 275 
<< m1 >>
rect 215 274 216 275 
<< m1 >>
rect 217 274 218 275 
<< m1 >>
rect 218 274 219 275 
<< m1 >>
rect 219 274 220 275 
<< m1 >>
rect 220 274 221 275 
<< m1 >>
rect 221 274 222 275 
<< m1 >>
rect 222 274 223 275 
<< m1 >>
rect 223 274 224 275 
<< m1 >>
rect 224 274 225 275 
<< m1 >>
rect 225 274 226 275 
<< m1 >>
rect 226 274 227 275 
<< m1 >>
rect 227 274 228 275 
<< m1 >>
rect 228 274 229 275 
<< m1 >>
rect 229 274 230 275 
<< m1 >>
rect 230 274 231 275 
<< m2 >>
rect 230 274 231 275 
<< m1 >>
rect 231 274 232 275 
<< m1 >>
rect 232 274 233 275 
<< m2 >>
rect 232 274 233 275 
<< m1 >>
rect 233 274 234 275 
<< m1 >>
rect 234 274 235 275 
<< m1 >>
rect 235 274 236 275 
<< m1 >>
rect 236 274 237 275 
<< m1 >>
rect 237 274 238 275 
<< m1 >>
rect 238 274 239 275 
<< m2 >>
rect 238 274 239 275 
<< m1 >>
rect 239 274 240 275 
<< m1 >>
rect 240 274 241 275 
<< m1 >>
rect 241 274 242 275 
<< m1 >>
rect 242 274 243 275 
<< m1 >>
rect 243 274 244 275 
<< m1 >>
rect 244 274 245 275 
<< m1 >>
rect 245 274 246 275 
<< m1 >>
rect 246 274 247 275 
<< m1 >>
rect 247 274 248 275 
<< m1 >>
rect 248 274 249 275 
<< m1 >>
rect 249 274 250 275 
<< m1 >>
rect 250 274 251 275 
<< m1 >>
rect 251 274 252 275 
<< m1 >>
rect 252 274 253 275 
<< m1 >>
rect 253 274 254 275 
<< m2 >>
rect 253 274 254 275 
<< m1 >>
rect 254 274 255 275 
<< m1 >>
rect 255 274 256 275 
<< m2 >>
rect 255 274 256 275 
<< m1 >>
rect 256 274 257 275 
<< m1 >>
rect 257 274 258 275 
<< m1 >>
rect 258 274 259 275 
<< m1 >>
rect 259 274 260 275 
<< m2 >>
rect 259 274 260 275 
<< m1 >>
rect 260 274 261 275 
<< m1 >>
rect 261 274 262 275 
<< m1 >>
rect 262 274 263 275 
<< m2 >>
rect 262 274 263 275 
<< m1 >>
rect 263 274 264 275 
<< m2 >>
rect 263 274 264 275 
<< m1 >>
rect 264 274 265 275 
<< m2 >>
rect 264 274 265 275 
<< m1 >>
rect 265 274 266 275 
<< m2 >>
rect 265 274 266 275 
<< m1 >>
rect 266 274 267 275 
<< m2 >>
rect 266 274 267 275 
<< m1 >>
rect 267 274 268 275 
<< m2 >>
rect 267 274 268 275 
<< m1 >>
rect 268 274 269 275 
<< m2 >>
rect 268 274 269 275 
<< m1 >>
rect 269 274 270 275 
<< m2 >>
rect 269 274 270 275 
<< m1 >>
rect 270 274 271 275 
<< m2 >>
rect 270 274 271 275 
<< m1 >>
rect 271 274 272 275 
<< m2 >>
rect 272 274 273 275 
<< m2 >>
rect 276 274 277 275 
<< m2 >>
rect 280 274 281 275 
<< m1 >>
rect 286 274 287 275 
<< m1 >>
rect 289 274 290 275 
<< m2 >>
rect 289 274 290 275 
<< m1 >>
rect 307 274 308 275 
<< m1 >>
rect 309 274 310 275 
<< m2 >>
rect 310 274 311 275 
<< m1 >>
rect 322 274 323 275 
<< m1 >>
rect 323 274 324 275 
<< m1 >>
rect 324 274 325 275 
<< m1 >>
rect 325 274 326 275 
<< m1 >>
rect 326 274 327 275 
<< m1 >>
rect 327 274 328 275 
<< m1 >>
rect 328 274 329 275 
<< m1 >>
rect 329 274 330 275 
<< m1 >>
rect 330 274 331 275 
<< m1 >>
rect 331 274 332 275 
<< m1 >>
rect 332 274 333 275 
<< m1 >>
rect 333 274 334 275 
<< m1 >>
rect 334 274 335 275 
<< m1 >>
rect 335 274 336 275 
<< m1 >>
rect 336 274 337 275 
<< m1 >>
rect 337 274 338 275 
<< m1 >>
rect 338 274 339 275 
<< m2 >>
rect 338 274 339 275 
<< m2c >>
rect 338 274 339 275 
<< m1 >>
rect 338 274 339 275 
<< m2 >>
rect 338 274 339 275 
<< m2 >>
rect 339 274 340 275 
<< m1 >>
rect 340 274 341 275 
<< m2 >>
rect 340 274 341 275 
<< m2 >>
rect 341 274 342 275 
<< m1 >>
rect 342 274 343 275 
<< m2 >>
rect 342 274 343 275 
<< m2c >>
rect 342 274 343 275 
<< m1 >>
rect 342 274 343 275 
<< m2 >>
rect 342 274 343 275 
<< m1 >>
rect 343 274 344 275 
<< m1 >>
rect 344 274 345 275 
<< m2 >>
rect 344 274 345 275 
<< m1 >>
rect 345 274 346 275 
<< m1 >>
rect 346 274 347 275 
<< m2 >>
rect 346 274 347 275 
<< m1 >>
rect 347 274 348 275 
<< m1 >>
rect 348 274 349 275 
<< m1 >>
rect 349 274 350 275 
<< m1 >>
rect 350 274 351 275 
<< m1 >>
rect 351 274 352 275 
<< m1 >>
rect 352 274 353 275 
<< m1 >>
rect 353 274 354 275 
<< m1 >>
rect 354 274 355 275 
<< m1 >>
rect 355 274 356 275 
<< m1 >>
rect 356 274 357 275 
<< m1 >>
rect 357 274 358 275 
<< m1 >>
rect 358 274 359 275 
<< m1 >>
rect 359 274 360 275 
<< m1 >>
rect 360 274 361 275 
<< m1 >>
rect 361 274 362 275 
<< m1 >>
rect 362 274 363 275 
<< m1 >>
rect 363 274 364 275 
<< m1 >>
rect 364 274 365 275 
<< m1 >>
rect 365 274 366 275 
<< m1 >>
rect 366 274 367 275 
<< m2 >>
rect 366 274 367 275 
<< m1 >>
rect 367 274 368 275 
<< m1 >>
rect 368 274 369 275 
<< m2 >>
rect 368 274 369 275 
<< m2c >>
rect 368 274 369 275 
<< m1 >>
rect 368 274 369 275 
<< m2 >>
rect 368 274 369 275 
<< m2 >>
rect 369 274 370 275 
<< m1 >>
rect 370 274 371 275 
<< m2 >>
rect 370 274 371 275 
<< m2 >>
rect 371 274 372 275 
<< m1 >>
rect 372 274 373 275 
<< m2 >>
rect 372 274 373 275 
<< m2c >>
rect 372 274 373 275 
<< m1 >>
rect 372 274 373 275 
<< m2 >>
rect 372 274 373 275 
<< m1 >>
rect 373 274 374 275 
<< m1 >>
rect 374 274 375 275 
<< m1 >>
rect 375 274 376 275 
<< m1 >>
rect 376 274 377 275 
<< m1 >>
rect 377 274 378 275 
<< m1 >>
rect 378 274 379 275 
<< m1 >>
rect 379 274 380 275 
<< m2 >>
rect 380 274 381 275 
<< m1 >>
rect 388 274 389 275 
<< m1 >>
rect 416 274 417 275 
<< m1 >>
rect 419 274 420 275 
<< m2 >>
rect 420 274 421 275 
<< m1 >>
rect 427 274 428 275 
<< m1 >>
rect 428 274 429 275 
<< m1 >>
rect 429 274 430 275 
<< m1 >>
rect 430 274 431 275 
<< m1 >>
rect 431 274 432 275 
<< m1 >>
rect 433 274 434 275 
<< m1 >>
rect 437 274 438 275 
<< m1 >>
rect 523 274 524 275 
<< m1 >>
rect 19 275 20 276 
<< m1 >>
rect 22 275 23 276 
<< m1 >>
rect 44 275 45 276 
<< m1 >>
rect 55 275 56 276 
<< m1 >>
rect 64 275 65 276 
<< m1 >>
rect 89 275 90 276 
<< m1 >>
rect 91 275 92 276 
<< m1 >>
rect 109 275 110 276 
<< m1 >>
rect 148 275 149 276 
<< m2 >>
rect 149 275 150 276 
<< m1 >>
rect 156 275 157 276 
<< m1 >>
rect 178 275 179 276 
<< m2 >>
rect 179 275 180 276 
<< m2 >>
rect 186 275 187 276 
<< m1 >>
rect 215 275 216 276 
<< m2 >>
rect 217 275 218 276 
<< m2 >>
rect 218 275 219 276 
<< m2 >>
rect 219 275 220 276 
<< m2 >>
rect 220 275 221 276 
<< m2 >>
rect 221 275 222 276 
<< m2 >>
rect 222 275 223 276 
<< m2 >>
rect 223 275 224 276 
<< m2 >>
rect 224 275 225 276 
<< m2 >>
rect 225 275 226 276 
<< m2 >>
rect 226 275 227 276 
<< m2 >>
rect 227 275 228 276 
<< m2 >>
rect 228 275 229 276 
<< m2 >>
rect 229 275 230 276 
<< m2 >>
rect 230 275 231 276 
<< m2 >>
rect 232 275 233 276 
<< m2 >>
rect 238 275 239 276 
<< m2 >>
rect 239 275 240 276 
<< m2 >>
rect 240 275 241 276 
<< m2 >>
rect 241 275 242 276 
<< m2 >>
rect 242 275 243 276 
<< m2 >>
rect 243 275 244 276 
<< m2 >>
rect 244 275 245 276 
<< m2 >>
rect 245 275 246 276 
<< m2 >>
rect 246 275 247 276 
<< m2 >>
rect 247 275 248 276 
<< m2 >>
rect 253 275 254 276 
<< m2 >>
rect 255 275 256 276 
<< m2 >>
rect 259 275 260 276 
<< m1 >>
rect 271 275 272 276 
<< m2 >>
rect 272 275 273 276 
<< m1 >>
rect 276 275 277 276 
<< m2 >>
rect 276 275 277 276 
<< m2c >>
rect 276 275 277 276 
<< m1 >>
rect 276 275 277 276 
<< m2 >>
rect 276 275 277 276 
<< m1 >>
rect 280 275 281 276 
<< m2 >>
rect 280 275 281 276 
<< m2c >>
rect 280 275 281 276 
<< m1 >>
rect 280 275 281 276 
<< m2 >>
rect 280 275 281 276 
<< m1 >>
rect 286 275 287 276 
<< m1 >>
rect 289 275 290 276 
<< m2 >>
rect 289 275 290 276 
<< m1 >>
rect 307 275 308 276 
<< m1 >>
rect 309 275 310 276 
<< m2 >>
rect 310 275 311 276 
<< m1 >>
rect 340 275 341 276 
<< m2 >>
rect 344 275 345 276 
<< m2 >>
rect 346 275 347 276 
<< m2 >>
rect 366 275 367 276 
<< m1 >>
rect 370 275 371 276 
<< m1 >>
rect 379 275 380 276 
<< m2 >>
rect 380 275 381 276 
<< m1 >>
rect 388 275 389 276 
<< m1 >>
rect 416 275 417 276 
<< m1 >>
rect 419 275 420 276 
<< m2 >>
rect 420 275 421 276 
<< m1 >>
rect 427 275 428 276 
<< m1 >>
rect 433 275 434 276 
<< m1 >>
rect 437 275 438 276 
<< m1 >>
rect 523 275 524 276 
<< m1 >>
rect 19 276 20 277 
<< m1 >>
rect 22 276 23 277 
<< m1 >>
rect 44 276 45 277 
<< m1 >>
rect 55 276 56 277 
<< m1 >>
rect 64 276 65 277 
<< m1 >>
rect 89 276 90 277 
<< m1 >>
rect 91 276 92 277 
<< m1 >>
rect 109 276 110 277 
<< m1 >>
rect 148 276 149 277 
<< m2 >>
rect 149 276 150 277 
<< m1 >>
rect 156 276 157 277 
<< m1 >>
rect 172 276 173 277 
<< m1 >>
rect 173 276 174 277 
<< m1 >>
rect 174 276 175 277 
<< m1 >>
rect 175 276 176 277 
<< m1 >>
rect 176 276 177 277 
<< m2 >>
rect 176 276 177 277 
<< m2c >>
rect 176 276 177 277 
<< m1 >>
rect 176 276 177 277 
<< m2 >>
rect 176 276 177 277 
<< m2 >>
rect 177 276 178 277 
<< m1 >>
rect 178 276 179 277 
<< m2 >>
rect 178 276 179 277 
<< m2 >>
rect 179 276 180 277 
<< m1 >>
rect 186 276 187 277 
<< m2 >>
rect 186 276 187 277 
<< m2c >>
rect 186 276 187 277 
<< m1 >>
rect 186 276 187 277 
<< m2 >>
rect 186 276 187 277 
<< m1 >>
rect 215 276 216 277 
<< m1 >>
rect 217 276 218 277 
<< m2 >>
rect 217 276 218 277 
<< m2c >>
rect 217 276 218 277 
<< m1 >>
rect 217 276 218 277 
<< m2 >>
rect 217 276 218 277 
<< m1 >>
rect 226 276 227 277 
<< m1 >>
rect 227 276 228 277 
<< m1 >>
rect 228 276 229 277 
<< m1 >>
rect 229 276 230 277 
<< m1 >>
rect 230 276 231 277 
<< m1 >>
rect 231 276 232 277 
<< m1 >>
rect 232 276 233 277 
<< m2 >>
rect 232 276 233 277 
<< m2c >>
rect 232 276 233 277 
<< m1 >>
rect 232 276 233 277 
<< m2 >>
rect 232 276 233 277 
<< m1 >>
rect 247 276 248 277 
<< m2 >>
rect 247 276 248 277 
<< m2c >>
rect 247 276 248 277 
<< m1 >>
rect 247 276 248 277 
<< m2 >>
rect 247 276 248 277 
<< m1 >>
rect 253 276 254 277 
<< m2 >>
rect 253 276 254 277 
<< m2c >>
rect 253 276 254 277 
<< m1 >>
rect 253 276 254 277 
<< m2 >>
rect 253 276 254 277 
<< m2 >>
rect 255 276 256 277 
<< m2 >>
rect 259 276 260 277 
<< m1 >>
rect 271 276 272 277 
<< m2 >>
rect 272 276 273 277 
<< m1 >>
rect 276 276 277 277 
<< m1 >>
rect 280 276 281 277 
<< m1 >>
rect 286 276 287 277 
<< m1 >>
rect 289 276 290 277 
<< m2 >>
rect 289 276 290 277 
<< m1 >>
rect 307 276 308 277 
<< m1 >>
rect 309 276 310 277 
<< m2 >>
rect 310 276 311 277 
<< m1 >>
rect 340 276 341 277 
<< m1 >>
rect 344 276 345 277 
<< m2 >>
rect 344 276 345 277 
<< m2c >>
rect 344 276 345 277 
<< m1 >>
rect 344 276 345 277 
<< m2 >>
rect 344 276 345 277 
<< m1 >>
rect 346 276 347 277 
<< m2 >>
rect 346 276 347 277 
<< m1 >>
rect 358 276 359 277 
<< m1 >>
rect 359 276 360 277 
<< m1 >>
rect 360 276 361 277 
<< m1 >>
rect 361 276 362 277 
<< m1 >>
rect 362 276 363 277 
<< m1 >>
rect 363 276 364 277 
<< m1 >>
rect 364 276 365 277 
<< m1 >>
rect 365 276 366 277 
<< m1 >>
rect 366 276 367 277 
<< m2 >>
rect 366 276 367 277 
<< m1 >>
rect 367 276 368 277 
<< m1 >>
rect 368 276 369 277 
<< m2 >>
rect 368 276 369 277 
<< m2c >>
rect 368 276 369 277 
<< m1 >>
rect 368 276 369 277 
<< m2 >>
rect 368 276 369 277 
<< m2 >>
rect 369 276 370 277 
<< m1 >>
rect 370 276 371 277 
<< m2 >>
rect 370 276 371 277 
<< m2 >>
rect 371 276 372 277 
<< m1 >>
rect 372 276 373 277 
<< m2 >>
rect 372 276 373 277 
<< m2c >>
rect 372 276 373 277 
<< m1 >>
rect 372 276 373 277 
<< m2 >>
rect 372 276 373 277 
<< m1 >>
rect 373 276 374 277 
<< m1 >>
rect 374 276 375 277 
<< m1 >>
rect 375 276 376 277 
<< m1 >>
rect 376 276 377 277 
<< m1 >>
rect 377 276 378 277 
<< m2 >>
rect 377 276 378 277 
<< m2c >>
rect 377 276 378 277 
<< m1 >>
rect 377 276 378 277 
<< m2 >>
rect 377 276 378 277 
<< m2 >>
rect 378 276 379 277 
<< m1 >>
rect 379 276 380 277 
<< m2 >>
rect 379 276 380 277 
<< m2 >>
rect 380 276 381 277 
<< m1 >>
rect 388 276 389 277 
<< m1 >>
rect 416 276 417 277 
<< m1 >>
rect 419 276 420 277 
<< m2 >>
rect 420 276 421 277 
<< m1 >>
rect 427 276 428 277 
<< m1 >>
rect 433 276 434 277 
<< m1 >>
rect 437 276 438 277 
<< m1 >>
rect 523 276 524 277 
<< m1 >>
rect 19 277 20 278 
<< m1 >>
rect 22 277 23 278 
<< m1 >>
rect 44 277 45 278 
<< m1 >>
rect 55 277 56 278 
<< m1 >>
rect 64 277 65 278 
<< m1 >>
rect 89 277 90 278 
<< m1 >>
rect 91 277 92 278 
<< m1 >>
rect 109 277 110 278 
<< m1 >>
rect 148 277 149 278 
<< m2 >>
rect 149 277 150 278 
<< m1 >>
rect 156 277 157 278 
<< m1 >>
rect 172 277 173 278 
<< m1 >>
rect 178 277 179 278 
<< m1 >>
rect 186 277 187 278 
<< m1 >>
rect 215 277 216 278 
<< m1 >>
rect 217 277 218 278 
<< m1 >>
rect 226 277 227 278 
<< m1 >>
rect 247 277 248 278 
<< m1 >>
rect 253 277 254 278 
<< m1 >>
rect 255 277 256 278 
<< m2 >>
rect 255 277 256 278 
<< m1 >>
rect 256 277 257 278 
<< m1 >>
rect 257 277 258 278 
<< m1 >>
rect 258 277 259 278 
<< m1 >>
rect 259 277 260 278 
<< m2 >>
rect 259 277 260 278 
<< m1 >>
rect 260 277 261 278 
<< m1 >>
rect 261 277 262 278 
<< m1 >>
rect 262 277 263 278 
<< m1 >>
rect 263 277 264 278 
<< m1 >>
rect 264 277 265 278 
<< m1 >>
rect 265 277 266 278 
<< m1 >>
rect 266 277 267 278 
<< m1 >>
rect 267 277 268 278 
<< m1 >>
rect 268 277 269 278 
<< m1 >>
rect 271 277 272 278 
<< m2 >>
rect 272 277 273 278 
<< m1 >>
rect 276 277 277 278 
<< m1 >>
rect 278 277 279 278 
<< m2 >>
rect 278 277 279 278 
<< m2c >>
rect 278 277 279 278 
<< m1 >>
rect 278 277 279 278 
<< m2 >>
rect 278 277 279 278 
<< m2 >>
rect 279 277 280 278 
<< m1 >>
rect 280 277 281 278 
<< m2 >>
rect 280 277 281 278 
<< m2 >>
rect 281 277 282 278 
<< m1 >>
rect 282 277 283 278 
<< m2 >>
rect 282 277 283 278 
<< m2c >>
rect 282 277 283 278 
<< m1 >>
rect 282 277 283 278 
<< m2 >>
rect 282 277 283 278 
<< m1 >>
rect 283 277 284 278 
<< m1 >>
rect 284 277 285 278 
<< m1 >>
rect 285 277 286 278 
<< m1 >>
rect 286 277 287 278 
<< m1 >>
rect 289 277 290 278 
<< m2 >>
rect 289 277 290 278 
<< m1 >>
rect 307 277 308 278 
<< m1 >>
rect 309 277 310 278 
<< m2 >>
rect 310 277 311 278 
<< m1 >>
rect 340 277 341 278 
<< m1 >>
rect 344 277 345 278 
<< m2 >>
rect 344 277 345 278 
<< m1 >>
rect 346 277 347 278 
<< m2 >>
rect 346 277 347 278 
<< m2c >>
rect 346 277 347 278 
<< m1 >>
rect 346 277 347 278 
<< m2 >>
rect 346 277 347 278 
<< m1 >>
rect 358 277 359 278 
<< m2 >>
rect 366 277 367 278 
<< m1 >>
rect 370 277 371 278 
<< m1 >>
rect 379 277 380 278 
<< m1 >>
rect 388 277 389 278 
<< m1 >>
rect 416 277 417 278 
<< m1 >>
rect 419 277 420 278 
<< m2 >>
rect 420 277 421 278 
<< m1 >>
rect 427 277 428 278 
<< m1 >>
rect 433 277 434 278 
<< m1 >>
rect 437 277 438 278 
<< m1 >>
rect 523 277 524 278 
<< m1 >>
rect 19 278 20 279 
<< m1 >>
rect 22 278 23 279 
<< m1 >>
rect 44 278 45 279 
<< m1 >>
rect 55 278 56 279 
<< m1 >>
rect 64 278 65 279 
<< m1 >>
rect 89 278 90 279 
<< m1 >>
rect 91 278 92 279 
<< m1 >>
rect 109 278 110 279 
<< m1 >>
rect 148 278 149 279 
<< m2 >>
rect 149 278 150 279 
<< m1 >>
rect 156 278 157 279 
<< m2 >>
rect 156 278 157 279 
<< m2c >>
rect 156 278 157 279 
<< m1 >>
rect 156 278 157 279 
<< m2 >>
rect 156 278 157 279 
<< m1 >>
rect 172 278 173 279 
<< m1 >>
rect 178 278 179 279 
<< m1 >>
rect 186 278 187 279 
<< m1 >>
rect 215 278 216 279 
<< m2 >>
rect 215 278 216 279 
<< m2c >>
rect 215 278 216 279 
<< m1 >>
rect 215 278 216 279 
<< m2 >>
rect 215 278 216 279 
<< m2 >>
rect 216 278 217 279 
<< m1 >>
rect 217 278 218 279 
<< m2 >>
rect 217 278 218 279 
<< m1 >>
rect 226 278 227 279 
<< m1 >>
rect 247 278 248 279 
<< m1 >>
rect 253 278 254 279 
<< m1 >>
rect 255 278 256 279 
<< m2 >>
rect 255 278 256 279 
<< m2 >>
rect 259 278 260 279 
<< m1 >>
rect 268 278 269 279 
<< m1 >>
rect 271 278 272 279 
<< m2 >>
rect 272 278 273 279 
<< m1 >>
rect 276 278 277 279 
<< m1 >>
rect 278 278 279 279 
<< m1 >>
rect 280 278 281 279 
<< m1 >>
rect 289 278 290 279 
<< m2 >>
rect 289 278 290 279 
<< m1 >>
rect 307 278 308 279 
<< m1 >>
rect 309 278 310 279 
<< m2 >>
rect 310 278 311 279 
<< m1 >>
rect 340 278 341 279 
<< m2 >>
rect 344 278 345 279 
<< m2 >>
rect 346 278 347 279 
<< m1 >>
rect 358 278 359 279 
<< m1 >>
rect 366 278 367 279 
<< m2 >>
rect 366 278 367 279 
<< m2c >>
rect 366 278 367 279 
<< m1 >>
rect 366 278 367 279 
<< m2 >>
rect 366 278 367 279 
<< m1 >>
rect 370 278 371 279 
<< m1 >>
rect 379 278 380 279 
<< m1 >>
rect 388 278 389 279 
<< m1 >>
rect 416 278 417 279 
<< m1 >>
rect 419 278 420 279 
<< m2 >>
rect 420 278 421 279 
<< m1 >>
rect 427 278 428 279 
<< m1 >>
rect 433 278 434 279 
<< m1 >>
rect 437 278 438 279 
<< m1 >>
rect 523 278 524 279 
<< m1 >>
rect 19 279 20 280 
<< m1 >>
rect 22 279 23 280 
<< m1 >>
rect 44 279 45 280 
<< m1 >>
rect 55 279 56 280 
<< m1 >>
rect 64 279 65 280 
<< m1 >>
rect 89 279 90 280 
<< m1 >>
rect 91 279 92 280 
<< m1 >>
rect 109 279 110 280 
<< m1 >>
rect 148 279 149 280 
<< m2 >>
rect 149 279 150 280 
<< m2 >>
rect 151 279 152 280 
<< m2 >>
rect 152 279 153 280 
<< m2 >>
rect 153 279 154 280 
<< m2 >>
rect 154 279 155 280 
<< m2 >>
rect 155 279 156 280 
<< m2 >>
rect 156 279 157 280 
<< m1 >>
rect 172 279 173 280 
<< m1 >>
rect 178 279 179 280 
<< m1 >>
rect 186 279 187 280 
<< m1 >>
rect 217 279 218 280 
<< m2 >>
rect 217 279 218 280 
<< m1 >>
rect 226 279 227 280 
<< m1 >>
rect 247 279 248 280 
<< m1 >>
rect 253 279 254 280 
<< m1 >>
rect 255 279 256 280 
<< m2 >>
rect 255 279 256 280 
<< m2 >>
rect 256 279 257 280 
<< m1 >>
rect 257 279 258 280 
<< m2 >>
rect 257 279 258 280 
<< m2c >>
rect 257 279 258 280 
<< m1 >>
rect 257 279 258 280 
<< m2 >>
rect 257 279 258 280 
<< m1 >>
rect 259 279 260 280 
<< m2 >>
rect 259 279 260 280 
<< m2c >>
rect 259 279 260 280 
<< m1 >>
rect 259 279 260 280 
<< m2 >>
rect 259 279 260 280 
<< m1 >>
rect 268 279 269 280 
<< m1 >>
rect 271 279 272 280 
<< m2 >>
rect 272 279 273 280 
<< m1 >>
rect 276 279 277 280 
<< m1 >>
rect 278 279 279 280 
<< m1 >>
rect 280 279 281 280 
<< m1 >>
rect 289 279 290 280 
<< m2 >>
rect 289 279 290 280 
<< m1 >>
rect 301 279 302 280 
<< m1 >>
rect 302 279 303 280 
<< m1 >>
rect 303 279 304 280 
<< m1 >>
rect 304 279 305 280 
<< m1 >>
rect 305 279 306 280 
<< m1 >>
rect 306 279 307 280 
<< m1 >>
rect 307 279 308 280 
<< m1 >>
rect 309 279 310 280 
<< m2 >>
rect 310 279 311 280 
<< m1 >>
rect 340 279 341 280 
<< m1 >>
rect 341 279 342 280 
<< m1 >>
rect 342 279 343 280 
<< m1 >>
rect 343 279 344 280 
<< m1 >>
rect 344 279 345 280 
<< m2 >>
rect 344 279 345 280 
<< m1 >>
rect 345 279 346 280 
<< m1 >>
rect 346 279 347 280 
<< m2 >>
rect 346 279 347 280 
<< m1 >>
rect 347 279 348 280 
<< m1 >>
rect 348 279 349 280 
<< m1 >>
rect 349 279 350 280 
<< m1 >>
rect 350 279 351 280 
<< m1 >>
rect 351 279 352 280 
<< m1 >>
rect 352 279 353 280 
<< m1 >>
rect 358 279 359 280 
<< m1 >>
rect 366 279 367 280 
<< m1 >>
rect 370 279 371 280 
<< m1 >>
rect 379 279 380 280 
<< m1 >>
rect 388 279 389 280 
<< m1 >>
rect 416 279 417 280 
<< m1 >>
rect 419 279 420 280 
<< m2 >>
rect 420 279 421 280 
<< m1 >>
rect 427 279 428 280 
<< m1 >>
rect 433 279 434 280 
<< m1 >>
rect 437 279 438 280 
<< m1 >>
rect 523 279 524 280 
<< m1 >>
rect 19 280 20 281 
<< m1 >>
rect 22 280 23 281 
<< m1 >>
rect 44 280 45 281 
<< m1 >>
rect 55 280 56 281 
<< m1 >>
rect 64 280 65 281 
<< m1 >>
rect 89 280 90 281 
<< m1 >>
rect 91 280 92 281 
<< m1 >>
rect 109 280 110 281 
<< m1 >>
rect 148 280 149 281 
<< m2 >>
rect 149 280 150 281 
<< m1 >>
rect 150 280 151 281 
<< m1 >>
rect 151 280 152 281 
<< m2 >>
rect 151 280 152 281 
<< m1 >>
rect 152 280 153 281 
<< m1 >>
rect 153 280 154 281 
<< m1 >>
rect 154 280 155 281 
<< m1 >>
rect 155 280 156 281 
<< m1 >>
rect 156 280 157 281 
<< m1 >>
rect 157 280 158 281 
<< m1 >>
rect 172 280 173 281 
<< m1 >>
rect 178 280 179 281 
<< m1 >>
rect 186 280 187 281 
<< m1 >>
rect 217 280 218 281 
<< m2 >>
rect 217 280 218 281 
<< m1 >>
rect 226 280 227 281 
<< m1 >>
rect 232 280 233 281 
<< m1 >>
rect 233 280 234 281 
<< m1 >>
rect 234 280 235 281 
<< m1 >>
rect 235 280 236 281 
<< m1 >>
rect 236 280 237 281 
<< m1 >>
rect 237 280 238 281 
<< m1 >>
rect 238 280 239 281 
<< m1 >>
rect 239 280 240 281 
<< m1 >>
rect 240 280 241 281 
<< m1 >>
rect 241 280 242 281 
<< m1 >>
rect 242 280 243 281 
<< m1 >>
rect 243 280 244 281 
<< m1 >>
rect 244 280 245 281 
<< m1 >>
rect 247 280 248 281 
<< m1 >>
rect 253 280 254 281 
<< m1 >>
rect 255 280 256 281 
<< m1 >>
rect 257 280 258 281 
<< m1 >>
rect 259 280 260 281 
<< m1 >>
rect 268 280 269 281 
<< m1 >>
rect 271 280 272 281 
<< m2 >>
rect 272 280 273 281 
<< m1 >>
rect 276 280 277 281 
<< m2 >>
rect 276 280 277 281 
<< m2c >>
rect 276 280 277 281 
<< m1 >>
rect 276 280 277 281 
<< m2 >>
rect 276 280 277 281 
<< m2 >>
rect 277 280 278 281 
<< m1 >>
rect 278 280 279 281 
<< m2 >>
rect 278 280 279 281 
<< m2 >>
rect 279 280 280 281 
<< m1 >>
rect 280 280 281 281 
<< m2 >>
rect 280 280 281 281 
<< m2 >>
rect 281 280 282 281 
<< m1 >>
rect 282 280 283 281 
<< m2 >>
rect 282 280 283 281 
<< m2c >>
rect 282 280 283 281 
<< m1 >>
rect 282 280 283 281 
<< m2 >>
rect 282 280 283 281 
<< m1 >>
rect 283 280 284 281 
<< m1 >>
rect 289 280 290 281 
<< m2 >>
rect 289 280 290 281 
<< m1 >>
rect 301 280 302 281 
<< m1 >>
rect 309 280 310 281 
<< m2 >>
rect 310 280 311 281 
<< m1 >>
rect 322 280 323 281 
<< m1 >>
rect 323 280 324 281 
<< m1 >>
rect 324 280 325 281 
<< m1 >>
rect 325 280 326 281 
<< m2 >>
rect 344 280 345 281 
<< m2 >>
rect 346 280 347 281 
<< m1 >>
rect 352 280 353 281 
<< m2 >>
rect 352 280 353 281 
<< m2 >>
rect 353 280 354 281 
<< m1 >>
rect 354 280 355 281 
<< m2 >>
rect 354 280 355 281 
<< m2c >>
rect 354 280 355 281 
<< m1 >>
rect 354 280 355 281 
<< m2 >>
rect 354 280 355 281 
<< m1 >>
rect 355 280 356 281 
<< m1 >>
rect 358 280 359 281 
<< m1 >>
rect 366 280 367 281 
<< m1 >>
rect 370 280 371 281 
<< m1 >>
rect 379 280 380 281 
<< m1 >>
rect 388 280 389 281 
<< m1 >>
rect 406 280 407 281 
<< m1 >>
rect 407 280 408 281 
<< m1 >>
rect 408 280 409 281 
<< m1 >>
rect 409 280 410 281 
<< m1 >>
rect 416 280 417 281 
<< m1 >>
rect 419 280 420 281 
<< m2 >>
rect 420 280 421 281 
<< m1 >>
rect 427 280 428 281 
<< m1 >>
rect 433 280 434 281 
<< m1 >>
rect 437 280 438 281 
<< m1 >>
rect 484 280 485 281 
<< m1 >>
rect 485 280 486 281 
<< m1 >>
rect 486 280 487 281 
<< m1 >>
rect 487 280 488 281 
<< m1 >>
rect 523 280 524 281 
<< m1 >>
rect 19 281 20 282 
<< m1 >>
rect 22 281 23 282 
<< m1 >>
rect 44 281 45 282 
<< m1 >>
rect 55 281 56 282 
<< m1 >>
rect 64 281 65 282 
<< m1 >>
rect 89 281 90 282 
<< m1 >>
rect 91 281 92 282 
<< m1 >>
rect 109 281 110 282 
<< m1 >>
rect 148 281 149 282 
<< m2 >>
rect 149 281 150 282 
<< m1 >>
rect 150 281 151 282 
<< m2 >>
rect 151 281 152 282 
<< m1 >>
rect 157 281 158 282 
<< m1 >>
rect 172 281 173 282 
<< m1 >>
rect 178 281 179 282 
<< m1 >>
rect 186 281 187 282 
<< m1 >>
rect 217 281 218 282 
<< m2 >>
rect 217 281 218 282 
<< m1 >>
rect 226 281 227 282 
<< m1 >>
rect 232 281 233 282 
<< m1 >>
rect 244 281 245 282 
<< m1 >>
rect 247 281 248 282 
<< m1 >>
rect 253 281 254 282 
<< m1 >>
rect 255 281 256 282 
<< m1 >>
rect 257 281 258 282 
<< m1 >>
rect 259 281 260 282 
<< m1 >>
rect 268 281 269 282 
<< m1 >>
rect 271 281 272 282 
<< m2 >>
rect 272 281 273 282 
<< m1 >>
rect 278 281 279 282 
<< m1 >>
rect 280 281 281 282 
<< m1 >>
rect 283 281 284 282 
<< m1 >>
rect 289 281 290 282 
<< m2 >>
rect 289 281 290 282 
<< m1 >>
rect 301 281 302 282 
<< m1 >>
rect 309 281 310 282 
<< m2 >>
rect 310 281 311 282 
<< m1 >>
rect 322 281 323 282 
<< m1 >>
rect 325 281 326 282 
<< m1 >>
rect 344 281 345 282 
<< m2 >>
rect 344 281 345 282 
<< m2c >>
rect 344 281 345 282 
<< m1 >>
rect 344 281 345 282 
<< m2 >>
rect 344 281 345 282 
<< m1 >>
rect 346 281 347 282 
<< m2 >>
rect 346 281 347 282 
<< m2c >>
rect 346 281 347 282 
<< m1 >>
rect 346 281 347 282 
<< m2 >>
rect 346 281 347 282 
<< m1 >>
rect 348 281 349 282 
<< m1 >>
rect 349 281 350 282 
<< m1 >>
rect 350 281 351 282 
<< m2 >>
rect 350 281 351 282 
<< m2c >>
rect 350 281 351 282 
<< m1 >>
rect 350 281 351 282 
<< m2 >>
rect 350 281 351 282 
<< m2 >>
rect 351 281 352 282 
<< m1 >>
rect 352 281 353 282 
<< m2 >>
rect 352 281 353 282 
<< m1 >>
rect 355 281 356 282 
<< m1 >>
rect 358 281 359 282 
<< m1 >>
rect 366 281 367 282 
<< m1 >>
rect 370 281 371 282 
<< m1 >>
rect 379 281 380 282 
<< m1 >>
rect 388 281 389 282 
<< m1 >>
rect 406 281 407 282 
<< m1 >>
rect 409 281 410 282 
<< m1 >>
rect 416 281 417 282 
<< m1 >>
rect 419 281 420 282 
<< m2 >>
rect 420 281 421 282 
<< m1 >>
rect 427 281 428 282 
<< m1 >>
rect 433 281 434 282 
<< m1 >>
rect 437 281 438 282 
<< m1 >>
rect 484 281 485 282 
<< m1 >>
rect 487 281 488 282 
<< m1 >>
rect 523 281 524 282 
<< pdiffusion >>
rect 12 282 13 283 
<< pdiffusion >>
rect 13 282 14 283 
<< pdiffusion >>
rect 14 282 15 283 
<< pdiffusion >>
rect 15 282 16 283 
<< pdiffusion >>
rect 16 282 17 283 
<< pdiffusion >>
rect 17 282 18 283 
<< m1 >>
rect 19 282 20 283 
<< m1 >>
rect 22 282 23 283 
<< pdiffusion >>
rect 30 282 31 283 
<< pdiffusion >>
rect 31 282 32 283 
<< pdiffusion >>
rect 32 282 33 283 
<< pdiffusion >>
rect 33 282 34 283 
<< pdiffusion >>
rect 34 282 35 283 
<< pdiffusion >>
rect 35 282 36 283 
<< m1 >>
rect 44 282 45 283 
<< pdiffusion >>
rect 48 282 49 283 
<< pdiffusion >>
rect 49 282 50 283 
<< pdiffusion >>
rect 50 282 51 283 
<< pdiffusion >>
rect 51 282 52 283 
<< pdiffusion >>
rect 52 282 53 283 
<< pdiffusion >>
rect 53 282 54 283 
<< m1 >>
rect 55 282 56 283 
<< m1 >>
rect 64 282 65 283 
<< pdiffusion >>
rect 66 282 67 283 
<< pdiffusion >>
rect 67 282 68 283 
<< pdiffusion >>
rect 68 282 69 283 
<< pdiffusion >>
rect 69 282 70 283 
<< pdiffusion >>
rect 70 282 71 283 
<< pdiffusion >>
rect 71 282 72 283 
<< m1 >>
rect 89 282 90 283 
<< m1 >>
rect 91 282 92 283 
<< pdiffusion >>
rect 102 282 103 283 
<< pdiffusion >>
rect 103 282 104 283 
<< pdiffusion >>
rect 104 282 105 283 
<< pdiffusion >>
rect 105 282 106 283 
<< pdiffusion >>
rect 106 282 107 283 
<< pdiffusion >>
rect 107 282 108 283 
<< m1 >>
rect 109 282 110 283 
<< pdiffusion >>
rect 120 282 121 283 
<< pdiffusion >>
rect 121 282 122 283 
<< pdiffusion >>
rect 122 282 123 283 
<< pdiffusion >>
rect 123 282 124 283 
<< pdiffusion >>
rect 124 282 125 283 
<< pdiffusion >>
rect 125 282 126 283 
<< pdiffusion >>
rect 138 282 139 283 
<< pdiffusion >>
rect 139 282 140 283 
<< pdiffusion >>
rect 140 282 141 283 
<< pdiffusion >>
rect 141 282 142 283 
<< pdiffusion >>
rect 142 282 143 283 
<< pdiffusion >>
rect 143 282 144 283 
<< m1 >>
rect 148 282 149 283 
<< m2 >>
rect 149 282 150 283 
<< m1 >>
rect 150 282 151 283 
<< m2 >>
rect 151 282 152 283 
<< pdiffusion >>
rect 156 282 157 283 
<< m1 >>
rect 157 282 158 283 
<< pdiffusion >>
rect 157 282 158 283 
<< pdiffusion >>
rect 158 282 159 283 
<< pdiffusion >>
rect 159 282 160 283 
<< pdiffusion >>
rect 160 282 161 283 
<< pdiffusion >>
rect 161 282 162 283 
<< m1 >>
rect 172 282 173 283 
<< pdiffusion >>
rect 174 282 175 283 
<< pdiffusion >>
rect 175 282 176 283 
<< pdiffusion >>
rect 176 282 177 283 
<< pdiffusion >>
rect 177 282 178 283 
<< m1 >>
rect 178 282 179 283 
<< pdiffusion >>
rect 178 282 179 283 
<< pdiffusion >>
rect 179 282 180 283 
<< m1 >>
rect 186 282 187 283 
<< pdiffusion >>
rect 192 282 193 283 
<< pdiffusion >>
rect 193 282 194 283 
<< pdiffusion >>
rect 194 282 195 283 
<< pdiffusion >>
rect 195 282 196 283 
<< pdiffusion >>
rect 196 282 197 283 
<< pdiffusion >>
rect 197 282 198 283 
<< pdiffusion >>
rect 210 282 211 283 
<< pdiffusion >>
rect 211 282 212 283 
<< pdiffusion >>
rect 212 282 213 283 
<< pdiffusion >>
rect 213 282 214 283 
<< pdiffusion >>
rect 214 282 215 283 
<< pdiffusion >>
rect 215 282 216 283 
<< m1 >>
rect 217 282 218 283 
<< m2 >>
rect 217 282 218 283 
<< m1 >>
rect 226 282 227 283 
<< pdiffusion >>
rect 228 282 229 283 
<< pdiffusion >>
rect 229 282 230 283 
<< pdiffusion >>
rect 230 282 231 283 
<< pdiffusion >>
rect 231 282 232 283 
<< m1 >>
rect 232 282 233 283 
<< pdiffusion >>
rect 232 282 233 283 
<< pdiffusion >>
rect 233 282 234 283 
<< m1 >>
rect 244 282 245 283 
<< pdiffusion >>
rect 246 282 247 283 
<< m1 >>
rect 247 282 248 283 
<< pdiffusion >>
rect 247 282 248 283 
<< pdiffusion >>
rect 248 282 249 283 
<< pdiffusion >>
rect 249 282 250 283 
<< pdiffusion >>
rect 250 282 251 283 
<< pdiffusion >>
rect 251 282 252 283 
<< m1 >>
rect 253 282 254 283 
<< m1 >>
rect 255 282 256 283 
<< m1 >>
rect 257 282 258 283 
<< m1 >>
rect 259 282 260 283 
<< pdiffusion >>
rect 264 282 265 283 
<< pdiffusion >>
rect 265 282 266 283 
<< pdiffusion >>
rect 266 282 267 283 
<< pdiffusion >>
rect 267 282 268 283 
<< m1 >>
rect 268 282 269 283 
<< pdiffusion >>
rect 268 282 269 283 
<< pdiffusion >>
rect 269 282 270 283 
<< m1 >>
rect 271 282 272 283 
<< m2 >>
rect 272 282 273 283 
<< m1 >>
rect 278 282 279 283 
<< m1 >>
rect 280 282 281 283 
<< pdiffusion >>
rect 282 282 283 283 
<< m1 >>
rect 283 282 284 283 
<< pdiffusion >>
rect 283 282 284 283 
<< pdiffusion >>
rect 284 282 285 283 
<< pdiffusion >>
rect 285 282 286 283 
<< pdiffusion >>
rect 286 282 287 283 
<< pdiffusion >>
rect 287 282 288 283 
<< m1 >>
rect 289 282 290 283 
<< m2 >>
rect 289 282 290 283 
<< pdiffusion >>
rect 300 282 301 283 
<< m1 >>
rect 301 282 302 283 
<< pdiffusion >>
rect 301 282 302 283 
<< pdiffusion >>
rect 302 282 303 283 
<< pdiffusion >>
rect 303 282 304 283 
<< pdiffusion >>
rect 304 282 305 283 
<< pdiffusion >>
rect 305 282 306 283 
<< m1 >>
rect 309 282 310 283 
<< m2 >>
rect 310 282 311 283 
<< pdiffusion >>
rect 318 282 319 283 
<< pdiffusion >>
rect 319 282 320 283 
<< pdiffusion >>
rect 320 282 321 283 
<< pdiffusion >>
rect 321 282 322 283 
<< m1 >>
rect 322 282 323 283 
<< pdiffusion >>
rect 322 282 323 283 
<< pdiffusion >>
rect 323 282 324 283 
<< m1 >>
rect 325 282 326 283 
<< pdiffusion >>
rect 336 282 337 283 
<< pdiffusion >>
rect 337 282 338 283 
<< pdiffusion >>
rect 338 282 339 283 
<< pdiffusion >>
rect 339 282 340 283 
<< pdiffusion >>
rect 340 282 341 283 
<< pdiffusion >>
rect 341 282 342 283 
<< m1 >>
rect 344 282 345 283 
<< m1 >>
rect 346 282 347 283 
<< m1 >>
rect 348 282 349 283 
<< m1 >>
rect 352 282 353 283 
<< pdiffusion >>
rect 354 282 355 283 
<< m1 >>
rect 355 282 356 283 
<< pdiffusion >>
rect 355 282 356 283 
<< pdiffusion >>
rect 356 282 357 283 
<< pdiffusion >>
rect 357 282 358 283 
<< m1 >>
rect 358 282 359 283 
<< pdiffusion >>
rect 358 282 359 283 
<< pdiffusion >>
rect 359 282 360 283 
<< m1 >>
rect 366 282 367 283 
<< m1 >>
rect 370 282 371 283 
<< pdiffusion >>
rect 372 282 373 283 
<< pdiffusion >>
rect 373 282 374 283 
<< pdiffusion >>
rect 374 282 375 283 
<< pdiffusion >>
rect 375 282 376 283 
<< pdiffusion >>
rect 376 282 377 283 
<< pdiffusion >>
rect 377 282 378 283 
<< m1 >>
rect 379 282 380 283 
<< m1 >>
rect 388 282 389 283 
<< pdiffusion >>
rect 390 282 391 283 
<< pdiffusion >>
rect 391 282 392 283 
<< pdiffusion >>
rect 392 282 393 283 
<< pdiffusion >>
rect 393 282 394 283 
<< pdiffusion >>
rect 394 282 395 283 
<< pdiffusion >>
rect 395 282 396 283 
<< m1 >>
rect 406 282 407 283 
<< pdiffusion >>
rect 408 282 409 283 
<< m1 >>
rect 409 282 410 283 
<< pdiffusion >>
rect 409 282 410 283 
<< pdiffusion >>
rect 410 282 411 283 
<< pdiffusion >>
rect 411 282 412 283 
<< pdiffusion >>
rect 412 282 413 283 
<< pdiffusion >>
rect 413 282 414 283 
<< m1 >>
rect 416 282 417 283 
<< m1 >>
rect 419 282 420 283 
<< m2 >>
rect 420 282 421 283 
<< pdiffusion >>
rect 426 282 427 283 
<< m1 >>
rect 427 282 428 283 
<< pdiffusion >>
rect 427 282 428 283 
<< pdiffusion >>
rect 428 282 429 283 
<< pdiffusion >>
rect 429 282 430 283 
<< pdiffusion >>
rect 430 282 431 283 
<< pdiffusion >>
rect 431 282 432 283 
<< m1 >>
rect 433 282 434 283 
<< m1 >>
rect 437 282 438 283 
<< pdiffusion >>
rect 444 282 445 283 
<< pdiffusion >>
rect 445 282 446 283 
<< pdiffusion >>
rect 446 282 447 283 
<< pdiffusion >>
rect 447 282 448 283 
<< pdiffusion >>
rect 448 282 449 283 
<< pdiffusion >>
rect 449 282 450 283 
<< pdiffusion >>
rect 462 282 463 283 
<< pdiffusion >>
rect 463 282 464 283 
<< pdiffusion >>
rect 464 282 465 283 
<< pdiffusion >>
rect 465 282 466 283 
<< pdiffusion >>
rect 466 282 467 283 
<< pdiffusion >>
rect 467 282 468 283 
<< pdiffusion >>
rect 480 282 481 283 
<< pdiffusion >>
rect 481 282 482 283 
<< pdiffusion >>
rect 482 282 483 283 
<< pdiffusion >>
rect 483 282 484 283 
<< m1 >>
rect 484 282 485 283 
<< pdiffusion >>
rect 484 282 485 283 
<< pdiffusion >>
rect 485 282 486 283 
<< m1 >>
rect 487 282 488 283 
<< pdiffusion >>
rect 498 282 499 283 
<< pdiffusion >>
rect 499 282 500 283 
<< pdiffusion >>
rect 500 282 501 283 
<< pdiffusion >>
rect 501 282 502 283 
<< pdiffusion >>
rect 502 282 503 283 
<< pdiffusion >>
rect 503 282 504 283 
<< pdiffusion >>
rect 516 282 517 283 
<< pdiffusion >>
rect 517 282 518 283 
<< pdiffusion >>
rect 518 282 519 283 
<< pdiffusion >>
rect 519 282 520 283 
<< pdiffusion >>
rect 520 282 521 283 
<< pdiffusion >>
rect 521 282 522 283 
<< m1 >>
rect 523 282 524 283 
<< pdiffusion >>
rect 12 283 13 284 
<< pdiffusion >>
rect 13 283 14 284 
<< pdiffusion >>
rect 14 283 15 284 
<< pdiffusion >>
rect 15 283 16 284 
<< pdiffusion >>
rect 16 283 17 284 
<< pdiffusion >>
rect 17 283 18 284 
<< m1 >>
rect 19 283 20 284 
<< m1 >>
rect 22 283 23 284 
<< pdiffusion >>
rect 30 283 31 284 
<< pdiffusion >>
rect 31 283 32 284 
<< pdiffusion >>
rect 32 283 33 284 
<< pdiffusion >>
rect 33 283 34 284 
<< pdiffusion >>
rect 34 283 35 284 
<< pdiffusion >>
rect 35 283 36 284 
<< m1 >>
rect 44 283 45 284 
<< pdiffusion >>
rect 48 283 49 284 
<< pdiffusion >>
rect 49 283 50 284 
<< pdiffusion >>
rect 50 283 51 284 
<< pdiffusion >>
rect 51 283 52 284 
<< pdiffusion >>
rect 52 283 53 284 
<< pdiffusion >>
rect 53 283 54 284 
<< m1 >>
rect 55 283 56 284 
<< m1 >>
rect 64 283 65 284 
<< pdiffusion >>
rect 66 283 67 284 
<< pdiffusion >>
rect 67 283 68 284 
<< pdiffusion >>
rect 68 283 69 284 
<< pdiffusion >>
rect 69 283 70 284 
<< pdiffusion >>
rect 70 283 71 284 
<< pdiffusion >>
rect 71 283 72 284 
<< m1 >>
rect 89 283 90 284 
<< m1 >>
rect 91 283 92 284 
<< pdiffusion >>
rect 102 283 103 284 
<< pdiffusion >>
rect 103 283 104 284 
<< pdiffusion >>
rect 104 283 105 284 
<< pdiffusion >>
rect 105 283 106 284 
<< pdiffusion >>
rect 106 283 107 284 
<< pdiffusion >>
rect 107 283 108 284 
<< m1 >>
rect 109 283 110 284 
<< pdiffusion >>
rect 120 283 121 284 
<< pdiffusion >>
rect 121 283 122 284 
<< pdiffusion >>
rect 122 283 123 284 
<< pdiffusion >>
rect 123 283 124 284 
<< pdiffusion >>
rect 124 283 125 284 
<< pdiffusion >>
rect 125 283 126 284 
<< pdiffusion >>
rect 138 283 139 284 
<< pdiffusion >>
rect 139 283 140 284 
<< pdiffusion >>
rect 140 283 141 284 
<< pdiffusion >>
rect 141 283 142 284 
<< pdiffusion >>
rect 142 283 143 284 
<< pdiffusion >>
rect 143 283 144 284 
<< m1 >>
rect 148 283 149 284 
<< m2 >>
rect 149 283 150 284 
<< m1 >>
rect 150 283 151 284 
<< m2 >>
rect 151 283 152 284 
<< pdiffusion >>
rect 156 283 157 284 
<< pdiffusion >>
rect 157 283 158 284 
<< pdiffusion >>
rect 158 283 159 284 
<< pdiffusion >>
rect 159 283 160 284 
<< pdiffusion >>
rect 160 283 161 284 
<< pdiffusion >>
rect 161 283 162 284 
<< m1 >>
rect 172 283 173 284 
<< pdiffusion >>
rect 174 283 175 284 
<< pdiffusion >>
rect 175 283 176 284 
<< pdiffusion >>
rect 176 283 177 284 
<< pdiffusion >>
rect 177 283 178 284 
<< pdiffusion >>
rect 178 283 179 284 
<< pdiffusion >>
rect 179 283 180 284 
<< m1 >>
rect 186 283 187 284 
<< pdiffusion >>
rect 192 283 193 284 
<< pdiffusion >>
rect 193 283 194 284 
<< pdiffusion >>
rect 194 283 195 284 
<< pdiffusion >>
rect 195 283 196 284 
<< pdiffusion >>
rect 196 283 197 284 
<< pdiffusion >>
rect 197 283 198 284 
<< pdiffusion >>
rect 210 283 211 284 
<< pdiffusion >>
rect 211 283 212 284 
<< pdiffusion >>
rect 212 283 213 284 
<< pdiffusion >>
rect 213 283 214 284 
<< pdiffusion >>
rect 214 283 215 284 
<< pdiffusion >>
rect 215 283 216 284 
<< m1 >>
rect 217 283 218 284 
<< m2 >>
rect 217 283 218 284 
<< m1 >>
rect 226 283 227 284 
<< pdiffusion >>
rect 228 283 229 284 
<< pdiffusion >>
rect 229 283 230 284 
<< pdiffusion >>
rect 230 283 231 284 
<< pdiffusion >>
rect 231 283 232 284 
<< pdiffusion >>
rect 232 283 233 284 
<< pdiffusion >>
rect 233 283 234 284 
<< m1 >>
rect 244 283 245 284 
<< pdiffusion >>
rect 246 283 247 284 
<< pdiffusion >>
rect 247 283 248 284 
<< pdiffusion >>
rect 248 283 249 284 
<< pdiffusion >>
rect 249 283 250 284 
<< pdiffusion >>
rect 250 283 251 284 
<< pdiffusion >>
rect 251 283 252 284 
<< m1 >>
rect 253 283 254 284 
<< m1 >>
rect 255 283 256 284 
<< m1 >>
rect 257 283 258 284 
<< m1 >>
rect 259 283 260 284 
<< pdiffusion >>
rect 264 283 265 284 
<< pdiffusion >>
rect 265 283 266 284 
<< pdiffusion >>
rect 266 283 267 284 
<< pdiffusion >>
rect 267 283 268 284 
<< pdiffusion >>
rect 268 283 269 284 
<< pdiffusion >>
rect 269 283 270 284 
<< m1 >>
rect 271 283 272 284 
<< m2 >>
rect 272 283 273 284 
<< m1 >>
rect 278 283 279 284 
<< m1 >>
rect 280 283 281 284 
<< pdiffusion >>
rect 282 283 283 284 
<< pdiffusion >>
rect 283 283 284 284 
<< pdiffusion >>
rect 284 283 285 284 
<< pdiffusion >>
rect 285 283 286 284 
<< pdiffusion >>
rect 286 283 287 284 
<< pdiffusion >>
rect 287 283 288 284 
<< m1 >>
rect 289 283 290 284 
<< m2 >>
rect 289 283 290 284 
<< pdiffusion >>
rect 300 283 301 284 
<< pdiffusion >>
rect 301 283 302 284 
<< pdiffusion >>
rect 302 283 303 284 
<< pdiffusion >>
rect 303 283 304 284 
<< pdiffusion >>
rect 304 283 305 284 
<< pdiffusion >>
rect 305 283 306 284 
<< m1 >>
rect 309 283 310 284 
<< m2 >>
rect 310 283 311 284 
<< pdiffusion >>
rect 318 283 319 284 
<< pdiffusion >>
rect 319 283 320 284 
<< pdiffusion >>
rect 320 283 321 284 
<< pdiffusion >>
rect 321 283 322 284 
<< pdiffusion >>
rect 322 283 323 284 
<< pdiffusion >>
rect 323 283 324 284 
<< m1 >>
rect 325 283 326 284 
<< pdiffusion >>
rect 336 283 337 284 
<< pdiffusion >>
rect 337 283 338 284 
<< pdiffusion >>
rect 338 283 339 284 
<< pdiffusion >>
rect 339 283 340 284 
<< pdiffusion >>
rect 340 283 341 284 
<< pdiffusion >>
rect 341 283 342 284 
<< m1 >>
rect 344 283 345 284 
<< m1 >>
rect 346 283 347 284 
<< m1 >>
rect 348 283 349 284 
<< m1 >>
rect 352 283 353 284 
<< pdiffusion >>
rect 354 283 355 284 
<< pdiffusion >>
rect 355 283 356 284 
<< pdiffusion >>
rect 356 283 357 284 
<< pdiffusion >>
rect 357 283 358 284 
<< pdiffusion >>
rect 358 283 359 284 
<< pdiffusion >>
rect 359 283 360 284 
<< m1 >>
rect 366 283 367 284 
<< m1 >>
rect 370 283 371 284 
<< pdiffusion >>
rect 372 283 373 284 
<< pdiffusion >>
rect 373 283 374 284 
<< pdiffusion >>
rect 374 283 375 284 
<< pdiffusion >>
rect 375 283 376 284 
<< pdiffusion >>
rect 376 283 377 284 
<< pdiffusion >>
rect 377 283 378 284 
<< m1 >>
rect 379 283 380 284 
<< m1 >>
rect 388 283 389 284 
<< pdiffusion >>
rect 390 283 391 284 
<< pdiffusion >>
rect 391 283 392 284 
<< pdiffusion >>
rect 392 283 393 284 
<< pdiffusion >>
rect 393 283 394 284 
<< pdiffusion >>
rect 394 283 395 284 
<< pdiffusion >>
rect 395 283 396 284 
<< m1 >>
rect 406 283 407 284 
<< pdiffusion >>
rect 408 283 409 284 
<< pdiffusion >>
rect 409 283 410 284 
<< pdiffusion >>
rect 410 283 411 284 
<< pdiffusion >>
rect 411 283 412 284 
<< pdiffusion >>
rect 412 283 413 284 
<< pdiffusion >>
rect 413 283 414 284 
<< m1 >>
rect 416 283 417 284 
<< m1 >>
rect 419 283 420 284 
<< m2 >>
rect 420 283 421 284 
<< pdiffusion >>
rect 426 283 427 284 
<< pdiffusion >>
rect 427 283 428 284 
<< pdiffusion >>
rect 428 283 429 284 
<< pdiffusion >>
rect 429 283 430 284 
<< pdiffusion >>
rect 430 283 431 284 
<< pdiffusion >>
rect 431 283 432 284 
<< m1 >>
rect 433 283 434 284 
<< m1 >>
rect 437 283 438 284 
<< pdiffusion >>
rect 444 283 445 284 
<< pdiffusion >>
rect 445 283 446 284 
<< pdiffusion >>
rect 446 283 447 284 
<< pdiffusion >>
rect 447 283 448 284 
<< pdiffusion >>
rect 448 283 449 284 
<< pdiffusion >>
rect 449 283 450 284 
<< pdiffusion >>
rect 462 283 463 284 
<< pdiffusion >>
rect 463 283 464 284 
<< pdiffusion >>
rect 464 283 465 284 
<< pdiffusion >>
rect 465 283 466 284 
<< pdiffusion >>
rect 466 283 467 284 
<< pdiffusion >>
rect 467 283 468 284 
<< pdiffusion >>
rect 480 283 481 284 
<< pdiffusion >>
rect 481 283 482 284 
<< pdiffusion >>
rect 482 283 483 284 
<< pdiffusion >>
rect 483 283 484 284 
<< pdiffusion >>
rect 484 283 485 284 
<< pdiffusion >>
rect 485 283 486 284 
<< m1 >>
rect 487 283 488 284 
<< pdiffusion >>
rect 498 283 499 284 
<< pdiffusion >>
rect 499 283 500 284 
<< pdiffusion >>
rect 500 283 501 284 
<< pdiffusion >>
rect 501 283 502 284 
<< pdiffusion >>
rect 502 283 503 284 
<< pdiffusion >>
rect 503 283 504 284 
<< pdiffusion >>
rect 516 283 517 284 
<< pdiffusion >>
rect 517 283 518 284 
<< pdiffusion >>
rect 518 283 519 284 
<< pdiffusion >>
rect 519 283 520 284 
<< pdiffusion >>
rect 520 283 521 284 
<< pdiffusion >>
rect 521 283 522 284 
<< m1 >>
rect 523 283 524 284 
<< pdiffusion >>
rect 12 284 13 285 
<< pdiffusion >>
rect 13 284 14 285 
<< pdiffusion >>
rect 14 284 15 285 
<< pdiffusion >>
rect 15 284 16 285 
<< pdiffusion >>
rect 16 284 17 285 
<< pdiffusion >>
rect 17 284 18 285 
<< m1 >>
rect 19 284 20 285 
<< m1 >>
rect 22 284 23 285 
<< pdiffusion >>
rect 30 284 31 285 
<< pdiffusion >>
rect 31 284 32 285 
<< pdiffusion >>
rect 32 284 33 285 
<< pdiffusion >>
rect 33 284 34 285 
<< pdiffusion >>
rect 34 284 35 285 
<< pdiffusion >>
rect 35 284 36 285 
<< m1 >>
rect 44 284 45 285 
<< pdiffusion >>
rect 48 284 49 285 
<< pdiffusion >>
rect 49 284 50 285 
<< pdiffusion >>
rect 50 284 51 285 
<< pdiffusion >>
rect 51 284 52 285 
<< pdiffusion >>
rect 52 284 53 285 
<< pdiffusion >>
rect 53 284 54 285 
<< m1 >>
rect 55 284 56 285 
<< m1 >>
rect 64 284 65 285 
<< pdiffusion >>
rect 66 284 67 285 
<< pdiffusion >>
rect 67 284 68 285 
<< pdiffusion >>
rect 68 284 69 285 
<< pdiffusion >>
rect 69 284 70 285 
<< pdiffusion >>
rect 70 284 71 285 
<< pdiffusion >>
rect 71 284 72 285 
<< m1 >>
rect 89 284 90 285 
<< m1 >>
rect 91 284 92 285 
<< pdiffusion >>
rect 102 284 103 285 
<< pdiffusion >>
rect 103 284 104 285 
<< pdiffusion >>
rect 104 284 105 285 
<< pdiffusion >>
rect 105 284 106 285 
<< pdiffusion >>
rect 106 284 107 285 
<< pdiffusion >>
rect 107 284 108 285 
<< m1 >>
rect 109 284 110 285 
<< pdiffusion >>
rect 120 284 121 285 
<< pdiffusion >>
rect 121 284 122 285 
<< pdiffusion >>
rect 122 284 123 285 
<< pdiffusion >>
rect 123 284 124 285 
<< pdiffusion >>
rect 124 284 125 285 
<< pdiffusion >>
rect 125 284 126 285 
<< pdiffusion >>
rect 138 284 139 285 
<< pdiffusion >>
rect 139 284 140 285 
<< pdiffusion >>
rect 140 284 141 285 
<< pdiffusion >>
rect 141 284 142 285 
<< pdiffusion >>
rect 142 284 143 285 
<< pdiffusion >>
rect 143 284 144 285 
<< m1 >>
rect 148 284 149 285 
<< m2 >>
rect 149 284 150 285 
<< m1 >>
rect 150 284 151 285 
<< m2 >>
rect 151 284 152 285 
<< pdiffusion >>
rect 156 284 157 285 
<< pdiffusion >>
rect 157 284 158 285 
<< pdiffusion >>
rect 158 284 159 285 
<< pdiffusion >>
rect 159 284 160 285 
<< pdiffusion >>
rect 160 284 161 285 
<< pdiffusion >>
rect 161 284 162 285 
<< m1 >>
rect 172 284 173 285 
<< pdiffusion >>
rect 174 284 175 285 
<< pdiffusion >>
rect 175 284 176 285 
<< pdiffusion >>
rect 176 284 177 285 
<< pdiffusion >>
rect 177 284 178 285 
<< pdiffusion >>
rect 178 284 179 285 
<< pdiffusion >>
rect 179 284 180 285 
<< m1 >>
rect 186 284 187 285 
<< pdiffusion >>
rect 192 284 193 285 
<< pdiffusion >>
rect 193 284 194 285 
<< pdiffusion >>
rect 194 284 195 285 
<< pdiffusion >>
rect 195 284 196 285 
<< pdiffusion >>
rect 196 284 197 285 
<< pdiffusion >>
rect 197 284 198 285 
<< pdiffusion >>
rect 210 284 211 285 
<< pdiffusion >>
rect 211 284 212 285 
<< pdiffusion >>
rect 212 284 213 285 
<< pdiffusion >>
rect 213 284 214 285 
<< pdiffusion >>
rect 214 284 215 285 
<< pdiffusion >>
rect 215 284 216 285 
<< m1 >>
rect 217 284 218 285 
<< m2 >>
rect 217 284 218 285 
<< m1 >>
rect 226 284 227 285 
<< pdiffusion >>
rect 228 284 229 285 
<< pdiffusion >>
rect 229 284 230 285 
<< pdiffusion >>
rect 230 284 231 285 
<< pdiffusion >>
rect 231 284 232 285 
<< pdiffusion >>
rect 232 284 233 285 
<< pdiffusion >>
rect 233 284 234 285 
<< m1 >>
rect 244 284 245 285 
<< pdiffusion >>
rect 246 284 247 285 
<< pdiffusion >>
rect 247 284 248 285 
<< pdiffusion >>
rect 248 284 249 285 
<< pdiffusion >>
rect 249 284 250 285 
<< pdiffusion >>
rect 250 284 251 285 
<< pdiffusion >>
rect 251 284 252 285 
<< m1 >>
rect 253 284 254 285 
<< m1 >>
rect 255 284 256 285 
<< m1 >>
rect 257 284 258 285 
<< m1 >>
rect 259 284 260 285 
<< pdiffusion >>
rect 264 284 265 285 
<< pdiffusion >>
rect 265 284 266 285 
<< pdiffusion >>
rect 266 284 267 285 
<< pdiffusion >>
rect 267 284 268 285 
<< pdiffusion >>
rect 268 284 269 285 
<< pdiffusion >>
rect 269 284 270 285 
<< m1 >>
rect 271 284 272 285 
<< m2 >>
rect 272 284 273 285 
<< m1 >>
rect 278 284 279 285 
<< m1 >>
rect 280 284 281 285 
<< pdiffusion >>
rect 282 284 283 285 
<< pdiffusion >>
rect 283 284 284 285 
<< pdiffusion >>
rect 284 284 285 285 
<< pdiffusion >>
rect 285 284 286 285 
<< pdiffusion >>
rect 286 284 287 285 
<< pdiffusion >>
rect 287 284 288 285 
<< m1 >>
rect 289 284 290 285 
<< m2 >>
rect 289 284 290 285 
<< pdiffusion >>
rect 300 284 301 285 
<< pdiffusion >>
rect 301 284 302 285 
<< pdiffusion >>
rect 302 284 303 285 
<< pdiffusion >>
rect 303 284 304 285 
<< pdiffusion >>
rect 304 284 305 285 
<< pdiffusion >>
rect 305 284 306 285 
<< m1 >>
rect 309 284 310 285 
<< m2 >>
rect 310 284 311 285 
<< pdiffusion >>
rect 318 284 319 285 
<< pdiffusion >>
rect 319 284 320 285 
<< pdiffusion >>
rect 320 284 321 285 
<< pdiffusion >>
rect 321 284 322 285 
<< pdiffusion >>
rect 322 284 323 285 
<< pdiffusion >>
rect 323 284 324 285 
<< m1 >>
rect 325 284 326 285 
<< pdiffusion >>
rect 336 284 337 285 
<< pdiffusion >>
rect 337 284 338 285 
<< pdiffusion >>
rect 338 284 339 285 
<< pdiffusion >>
rect 339 284 340 285 
<< pdiffusion >>
rect 340 284 341 285 
<< pdiffusion >>
rect 341 284 342 285 
<< m1 >>
rect 344 284 345 285 
<< m1 >>
rect 346 284 347 285 
<< m1 >>
rect 348 284 349 285 
<< m1 >>
rect 352 284 353 285 
<< pdiffusion >>
rect 354 284 355 285 
<< pdiffusion >>
rect 355 284 356 285 
<< pdiffusion >>
rect 356 284 357 285 
<< pdiffusion >>
rect 357 284 358 285 
<< pdiffusion >>
rect 358 284 359 285 
<< pdiffusion >>
rect 359 284 360 285 
<< m1 >>
rect 366 284 367 285 
<< m1 >>
rect 370 284 371 285 
<< pdiffusion >>
rect 372 284 373 285 
<< pdiffusion >>
rect 373 284 374 285 
<< pdiffusion >>
rect 374 284 375 285 
<< pdiffusion >>
rect 375 284 376 285 
<< pdiffusion >>
rect 376 284 377 285 
<< pdiffusion >>
rect 377 284 378 285 
<< m1 >>
rect 379 284 380 285 
<< m1 >>
rect 388 284 389 285 
<< pdiffusion >>
rect 390 284 391 285 
<< pdiffusion >>
rect 391 284 392 285 
<< pdiffusion >>
rect 392 284 393 285 
<< pdiffusion >>
rect 393 284 394 285 
<< pdiffusion >>
rect 394 284 395 285 
<< pdiffusion >>
rect 395 284 396 285 
<< m1 >>
rect 406 284 407 285 
<< pdiffusion >>
rect 408 284 409 285 
<< pdiffusion >>
rect 409 284 410 285 
<< pdiffusion >>
rect 410 284 411 285 
<< pdiffusion >>
rect 411 284 412 285 
<< pdiffusion >>
rect 412 284 413 285 
<< pdiffusion >>
rect 413 284 414 285 
<< m1 >>
rect 416 284 417 285 
<< m1 >>
rect 419 284 420 285 
<< m2 >>
rect 420 284 421 285 
<< pdiffusion >>
rect 426 284 427 285 
<< pdiffusion >>
rect 427 284 428 285 
<< pdiffusion >>
rect 428 284 429 285 
<< pdiffusion >>
rect 429 284 430 285 
<< pdiffusion >>
rect 430 284 431 285 
<< pdiffusion >>
rect 431 284 432 285 
<< m1 >>
rect 433 284 434 285 
<< m1 >>
rect 437 284 438 285 
<< pdiffusion >>
rect 444 284 445 285 
<< pdiffusion >>
rect 445 284 446 285 
<< pdiffusion >>
rect 446 284 447 285 
<< pdiffusion >>
rect 447 284 448 285 
<< pdiffusion >>
rect 448 284 449 285 
<< pdiffusion >>
rect 449 284 450 285 
<< pdiffusion >>
rect 462 284 463 285 
<< pdiffusion >>
rect 463 284 464 285 
<< pdiffusion >>
rect 464 284 465 285 
<< pdiffusion >>
rect 465 284 466 285 
<< pdiffusion >>
rect 466 284 467 285 
<< pdiffusion >>
rect 467 284 468 285 
<< pdiffusion >>
rect 480 284 481 285 
<< pdiffusion >>
rect 481 284 482 285 
<< pdiffusion >>
rect 482 284 483 285 
<< pdiffusion >>
rect 483 284 484 285 
<< pdiffusion >>
rect 484 284 485 285 
<< pdiffusion >>
rect 485 284 486 285 
<< m1 >>
rect 487 284 488 285 
<< pdiffusion >>
rect 498 284 499 285 
<< pdiffusion >>
rect 499 284 500 285 
<< pdiffusion >>
rect 500 284 501 285 
<< pdiffusion >>
rect 501 284 502 285 
<< pdiffusion >>
rect 502 284 503 285 
<< pdiffusion >>
rect 503 284 504 285 
<< pdiffusion >>
rect 516 284 517 285 
<< pdiffusion >>
rect 517 284 518 285 
<< pdiffusion >>
rect 518 284 519 285 
<< pdiffusion >>
rect 519 284 520 285 
<< pdiffusion >>
rect 520 284 521 285 
<< pdiffusion >>
rect 521 284 522 285 
<< m1 >>
rect 523 284 524 285 
<< pdiffusion >>
rect 12 285 13 286 
<< pdiffusion >>
rect 13 285 14 286 
<< pdiffusion >>
rect 14 285 15 286 
<< pdiffusion >>
rect 15 285 16 286 
<< pdiffusion >>
rect 16 285 17 286 
<< pdiffusion >>
rect 17 285 18 286 
<< m1 >>
rect 19 285 20 286 
<< m1 >>
rect 22 285 23 286 
<< pdiffusion >>
rect 30 285 31 286 
<< pdiffusion >>
rect 31 285 32 286 
<< pdiffusion >>
rect 32 285 33 286 
<< pdiffusion >>
rect 33 285 34 286 
<< pdiffusion >>
rect 34 285 35 286 
<< pdiffusion >>
rect 35 285 36 286 
<< m1 >>
rect 44 285 45 286 
<< pdiffusion >>
rect 48 285 49 286 
<< pdiffusion >>
rect 49 285 50 286 
<< pdiffusion >>
rect 50 285 51 286 
<< pdiffusion >>
rect 51 285 52 286 
<< pdiffusion >>
rect 52 285 53 286 
<< pdiffusion >>
rect 53 285 54 286 
<< m1 >>
rect 55 285 56 286 
<< m1 >>
rect 64 285 65 286 
<< pdiffusion >>
rect 66 285 67 286 
<< pdiffusion >>
rect 67 285 68 286 
<< pdiffusion >>
rect 68 285 69 286 
<< pdiffusion >>
rect 69 285 70 286 
<< pdiffusion >>
rect 70 285 71 286 
<< pdiffusion >>
rect 71 285 72 286 
<< m1 >>
rect 89 285 90 286 
<< m1 >>
rect 91 285 92 286 
<< pdiffusion >>
rect 102 285 103 286 
<< pdiffusion >>
rect 103 285 104 286 
<< pdiffusion >>
rect 104 285 105 286 
<< pdiffusion >>
rect 105 285 106 286 
<< pdiffusion >>
rect 106 285 107 286 
<< pdiffusion >>
rect 107 285 108 286 
<< m1 >>
rect 109 285 110 286 
<< pdiffusion >>
rect 120 285 121 286 
<< pdiffusion >>
rect 121 285 122 286 
<< pdiffusion >>
rect 122 285 123 286 
<< pdiffusion >>
rect 123 285 124 286 
<< pdiffusion >>
rect 124 285 125 286 
<< pdiffusion >>
rect 125 285 126 286 
<< pdiffusion >>
rect 138 285 139 286 
<< pdiffusion >>
rect 139 285 140 286 
<< pdiffusion >>
rect 140 285 141 286 
<< pdiffusion >>
rect 141 285 142 286 
<< pdiffusion >>
rect 142 285 143 286 
<< pdiffusion >>
rect 143 285 144 286 
<< m1 >>
rect 148 285 149 286 
<< m2 >>
rect 149 285 150 286 
<< m1 >>
rect 150 285 151 286 
<< m2 >>
rect 151 285 152 286 
<< pdiffusion >>
rect 156 285 157 286 
<< pdiffusion >>
rect 157 285 158 286 
<< pdiffusion >>
rect 158 285 159 286 
<< pdiffusion >>
rect 159 285 160 286 
<< pdiffusion >>
rect 160 285 161 286 
<< pdiffusion >>
rect 161 285 162 286 
<< m1 >>
rect 172 285 173 286 
<< pdiffusion >>
rect 174 285 175 286 
<< pdiffusion >>
rect 175 285 176 286 
<< pdiffusion >>
rect 176 285 177 286 
<< pdiffusion >>
rect 177 285 178 286 
<< pdiffusion >>
rect 178 285 179 286 
<< pdiffusion >>
rect 179 285 180 286 
<< m1 >>
rect 186 285 187 286 
<< pdiffusion >>
rect 192 285 193 286 
<< pdiffusion >>
rect 193 285 194 286 
<< pdiffusion >>
rect 194 285 195 286 
<< pdiffusion >>
rect 195 285 196 286 
<< pdiffusion >>
rect 196 285 197 286 
<< pdiffusion >>
rect 197 285 198 286 
<< pdiffusion >>
rect 210 285 211 286 
<< pdiffusion >>
rect 211 285 212 286 
<< pdiffusion >>
rect 212 285 213 286 
<< pdiffusion >>
rect 213 285 214 286 
<< pdiffusion >>
rect 214 285 215 286 
<< pdiffusion >>
rect 215 285 216 286 
<< m1 >>
rect 217 285 218 286 
<< m2 >>
rect 217 285 218 286 
<< m1 >>
rect 226 285 227 286 
<< pdiffusion >>
rect 228 285 229 286 
<< pdiffusion >>
rect 229 285 230 286 
<< pdiffusion >>
rect 230 285 231 286 
<< pdiffusion >>
rect 231 285 232 286 
<< pdiffusion >>
rect 232 285 233 286 
<< pdiffusion >>
rect 233 285 234 286 
<< m1 >>
rect 244 285 245 286 
<< pdiffusion >>
rect 246 285 247 286 
<< pdiffusion >>
rect 247 285 248 286 
<< pdiffusion >>
rect 248 285 249 286 
<< pdiffusion >>
rect 249 285 250 286 
<< pdiffusion >>
rect 250 285 251 286 
<< pdiffusion >>
rect 251 285 252 286 
<< m1 >>
rect 253 285 254 286 
<< m1 >>
rect 255 285 256 286 
<< m1 >>
rect 257 285 258 286 
<< m1 >>
rect 259 285 260 286 
<< pdiffusion >>
rect 264 285 265 286 
<< pdiffusion >>
rect 265 285 266 286 
<< pdiffusion >>
rect 266 285 267 286 
<< pdiffusion >>
rect 267 285 268 286 
<< pdiffusion >>
rect 268 285 269 286 
<< pdiffusion >>
rect 269 285 270 286 
<< m1 >>
rect 271 285 272 286 
<< m2 >>
rect 272 285 273 286 
<< m1 >>
rect 278 285 279 286 
<< m1 >>
rect 280 285 281 286 
<< pdiffusion >>
rect 282 285 283 286 
<< pdiffusion >>
rect 283 285 284 286 
<< pdiffusion >>
rect 284 285 285 286 
<< pdiffusion >>
rect 285 285 286 286 
<< pdiffusion >>
rect 286 285 287 286 
<< pdiffusion >>
rect 287 285 288 286 
<< m1 >>
rect 289 285 290 286 
<< m2 >>
rect 289 285 290 286 
<< pdiffusion >>
rect 300 285 301 286 
<< pdiffusion >>
rect 301 285 302 286 
<< pdiffusion >>
rect 302 285 303 286 
<< pdiffusion >>
rect 303 285 304 286 
<< pdiffusion >>
rect 304 285 305 286 
<< pdiffusion >>
rect 305 285 306 286 
<< m1 >>
rect 309 285 310 286 
<< m2 >>
rect 310 285 311 286 
<< pdiffusion >>
rect 318 285 319 286 
<< pdiffusion >>
rect 319 285 320 286 
<< pdiffusion >>
rect 320 285 321 286 
<< pdiffusion >>
rect 321 285 322 286 
<< pdiffusion >>
rect 322 285 323 286 
<< pdiffusion >>
rect 323 285 324 286 
<< m1 >>
rect 325 285 326 286 
<< pdiffusion >>
rect 336 285 337 286 
<< pdiffusion >>
rect 337 285 338 286 
<< pdiffusion >>
rect 338 285 339 286 
<< pdiffusion >>
rect 339 285 340 286 
<< pdiffusion >>
rect 340 285 341 286 
<< pdiffusion >>
rect 341 285 342 286 
<< m1 >>
rect 344 285 345 286 
<< m1 >>
rect 346 285 347 286 
<< m1 >>
rect 348 285 349 286 
<< m1 >>
rect 352 285 353 286 
<< pdiffusion >>
rect 354 285 355 286 
<< pdiffusion >>
rect 355 285 356 286 
<< pdiffusion >>
rect 356 285 357 286 
<< pdiffusion >>
rect 357 285 358 286 
<< pdiffusion >>
rect 358 285 359 286 
<< pdiffusion >>
rect 359 285 360 286 
<< m1 >>
rect 366 285 367 286 
<< m1 >>
rect 370 285 371 286 
<< pdiffusion >>
rect 372 285 373 286 
<< pdiffusion >>
rect 373 285 374 286 
<< pdiffusion >>
rect 374 285 375 286 
<< pdiffusion >>
rect 375 285 376 286 
<< pdiffusion >>
rect 376 285 377 286 
<< pdiffusion >>
rect 377 285 378 286 
<< m1 >>
rect 379 285 380 286 
<< m1 >>
rect 388 285 389 286 
<< pdiffusion >>
rect 390 285 391 286 
<< pdiffusion >>
rect 391 285 392 286 
<< pdiffusion >>
rect 392 285 393 286 
<< pdiffusion >>
rect 393 285 394 286 
<< pdiffusion >>
rect 394 285 395 286 
<< pdiffusion >>
rect 395 285 396 286 
<< m1 >>
rect 406 285 407 286 
<< pdiffusion >>
rect 408 285 409 286 
<< pdiffusion >>
rect 409 285 410 286 
<< pdiffusion >>
rect 410 285 411 286 
<< pdiffusion >>
rect 411 285 412 286 
<< pdiffusion >>
rect 412 285 413 286 
<< pdiffusion >>
rect 413 285 414 286 
<< m1 >>
rect 416 285 417 286 
<< m1 >>
rect 419 285 420 286 
<< m2 >>
rect 420 285 421 286 
<< pdiffusion >>
rect 426 285 427 286 
<< pdiffusion >>
rect 427 285 428 286 
<< pdiffusion >>
rect 428 285 429 286 
<< pdiffusion >>
rect 429 285 430 286 
<< pdiffusion >>
rect 430 285 431 286 
<< pdiffusion >>
rect 431 285 432 286 
<< m1 >>
rect 433 285 434 286 
<< m1 >>
rect 437 285 438 286 
<< pdiffusion >>
rect 444 285 445 286 
<< pdiffusion >>
rect 445 285 446 286 
<< pdiffusion >>
rect 446 285 447 286 
<< pdiffusion >>
rect 447 285 448 286 
<< pdiffusion >>
rect 448 285 449 286 
<< pdiffusion >>
rect 449 285 450 286 
<< pdiffusion >>
rect 462 285 463 286 
<< pdiffusion >>
rect 463 285 464 286 
<< pdiffusion >>
rect 464 285 465 286 
<< pdiffusion >>
rect 465 285 466 286 
<< pdiffusion >>
rect 466 285 467 286 
<< pdiffusion >>
rect 467 285 468 286 
<< pdiffusion >>
rect 480 285 481 286 
<< pdiffusion >>
rect 481 285 482 286 
<< pdiffusion >>
rect 482 285 483 286 
<< pdiffusion >>
rect 483 285 484 286 
<< pdiffusion >>
rect 484 285 485 286 
<< pdiffusion >>
rect 485 285 486 286 
<< m1 >>
rect 487 285 488 286 
<< pdiffusion >>
rect 498 285 499 286 
<< pdiffusion >>
rect 499 285 500 286 
<< pdiffusion >>
rect 500 285 501 286 
<< pdiffusion >>
rect 501 285 502 286 
<< pdiffusion >>
rect 502 285 503 286 
<< pdiffusion >>
rect 503 285 504 286 
<< pdiffusion >>
rect 516 285 517 286 
<< pdiffusion >>
rect 517 285 518 286 
<< pdiffusion >>
rect 518 285 519 286 
<< pdiffusion >>
rect 519 285 520 286 
<< pdiffusion >>
rect 520 285 521 286 
<< pdiffusion >>
rect 521 285 522 286 
<< m1 >>
rect 523 285 524 286 
<< pdiffusion >>
rect 12 286 13 287 
<< pdiffusion >>
rect 13 286 14 287 
<< pdiffusion >>
rect 14 286 15 287 
<< pdiffusion >>
rect 15 286 16 287 
<< pdiffusion >>
rect 16 286 17 287 
<< pdiffusion >>
rect 17 286 18 287 
<< m1 >>
rect 19 286 20 287 
<< m1 >>
rect 22 286 23 287 
<< pdiffusion >>
rect 30 286 31 287 
<< pdiffusion >>
rect 31 286 32 287 
<< pdiffusion >>
rect 32 286 33 287 
<< pdiffusion >>
rect 33 286 34 287 
<< pdiffusion >>
rect 34 286 35 287 
<< pdiffusion >>
rect 35 286 36 287 
<< m1 >>
rect 44 286 45 287 
<< pdiffusion >>
rect 48 286 49 287 
<< pdiffusion >>
rect 49 286 50 287 
<< pdiffusion >>
rect 50 286 51 287 
<< pdiffusion >>
rect 51 286 52 287 
<< pdiffusion >>
rect 52 286 53 287 
<< pdiffusion >>
rect 53 286 54 287 
<< m1 >>
rect 55 286 56 287 
<< m1 >>
rect 64 286 65 287 
<< pdiffusion >>
rect 66 286 67 287 
<< pdiffusion >>
rect 67 286 68 287 
<< pdiffusion >>
rect 68 286 69 287 
<< pdiffusion >>
rect 69 286 70 287 
<< pdiffusion >>
rect 70 286 71 287 
<< pdiffusion >>
rect 71 286 72 287 
<< m1 >>
rect 89 286 90 287 
<< m1 >>
rect 91 286 92 287 
<< pdiffusion >>
rect 102 286 103 287 
<< pdiffusion >>
rect 103 286 104 287 
<< pdiffusion >>
rect 104 286 105 287 
<< pdiffusion >>
rect 105 286 106 287 
<< pdiffusion >>
rect 106 286 107 287 
<< pdiffusion >>
rect 107 286 108 287 
<< m1 >>
rect 109 286 110 287 
<< pdiffusion >>
rect 120 286 121 287 
<< pdiffusion >>
rect 121 286 122 287 
<< pdiffusion >>
rect 122 286 123 287 
<< pdiffusion >>
rect 123 286 124 287 
<< pdiffusion >>
rect 124 286 125 287 
<< pdiffusion >>
rect 125 286 126 287 
<< pdiffusion >>
rect 138 286 139 287 
<< pdiffusion >>
rect 139 286 140 287 
<< pdiffusion >>
rect 140 286 141 287 
<< pdiffusion >>
rect 141 286 142 287 
<< pdiffusion >>
rect 142 286 143 287 
<< pdiffusion >>
rect 143 286 144 287 
<< m1 >>
rect 148 286 149 287 
<< m2 >>
rect 149 286 150 287 
<< m1 >>
rect 150 286 151 287 
<< m2 >>
rect 151 286 152 287 
<< pdiffusion >>
rect 156 286 157 287 
<< pdiffusion >>
rect 157 286 158 287 
<< pdiffusion >>
rect 158 286 159 287 
<< pdiffusion >>
rect 159 286 160 287 
<< pdiffusion >>
rect 160 286 161 287 
<< pdiffusion >>
rect 161 286 162 287 
<< m1 >>
rect 172 286 173 287 
<< pdiffusion >>
rect 174 286 175 287 
<< pdiffusion >>
rect 175 286 176 287 
<< pdiffusion >>
rect 176 286 177 287 
<< pdiffusion >>
rect 177 286 178 287 
<< pdiffusion >>
rect 178 286 179 287 
<< pdiffusion >>
rect 179 286 180 287 
<< m1 >>
rect 186 286 187 287 
<< pdiffusion >>
rect 192 286 193 287 
<< pdiffusion >>
rect 193 286 194 287 
<< pdiffusion >>
rect 194 286 195 287 
<< pdiffusion >>
rect 195 286 196 287 
<< pdiffusion >>
rect 196 286 197 287 
<< pdiffusion >>
rect 197 286 198 287 
<< pdiffusion >>
rect 210 286 211 287 
<< pdiffusion >>
rect 211 286 212 287 
<< pdiffusion >>
rect 212 286 213 287 
<< pdiffusion >>
rect 213 286 214 287 
<< pdiffusion >>
rect 214 286 215 287 
<< pdiffusion >>
rect 215 286 216 287 
<< m1 >>
rect 217 286 218 287 
<< m2 >>
rect 217 286 218 287 
<< m1 >>
rect 226 286 227 287 
<< pdiffusion >>
rect 228 286 229 287 
<< pdiffusion >>
rect 229 286 230 287 
<< pdiffusion >>
rect 230 286 231 287 
<< pdiffusion >>
rect 231 286 232 287 
<< pdiffusion >>
rect 232 286 233 287 
<< pdiffusion >>
rect 233 286 234 287 
<< m1 >>
rect 244 286 245 287 
<< pdiffusion >>
rect 246 286 247 287 
<< pdiffusion >>
rect 247 286 248 287 
<< pdiffusion >>
rect 248 286 249 287 
<< pdiffusion >>
rect 249 286 250 287 
<< pdiffusion >>
rect 250 286 251 287 
<< pdiffusion >>
rect 251 286 252 287 
<< m1 >>
rect 253 286 254 287 
<< m1 >>
rect 255 286 256 287 
<< m1 >>
rect 257 286 258 287 
<< m1 >>
rect 259 286 260 287 
<< pdiffusion >>
rect 264 286 265 287 
<< pdiffusion >>
rect 265 286 266 287 
<< pdiffusion >>
rect 266 286 267 287 
<< pdiffusion >>
rect 267 286 268 287 
<< pdiffusion >>
rect 268 286 269 287 
<< pdiffusion >>
rect 269 286 270 287 
<< m1 >>
rect 271 286 272 287 
<< m2 >>
rect 272 286 273 287 
<< m1 >>
rect 278 286 279 287 
<< m1 >>
rect 280 286 281 287 
<< pdiffusion >>
rect 282 286 283 287 
<< pdiffusion >>
rect 283 286 284 287 
<< pdiffusion >>
rect 284 286 285 287 
<< pdiffusion >>
rect 285 286 286 287 
<< pdiffusion >>
rect 286 286 287 287 
<< pdiffusion >>
rect 287 286 288 287 
<< m1 >>
rect 289 286 290 287 
<< m2 >>
rect 289 286 290 287 
<< pdiffusion >>
rect 300 286 301 287 
<< pdiffusion >>
rect 301 286 302 287 
<< pdiffusion >>
rect 302 286 303 287 
<< pdiffusion >>
rect 303 286 304 287 
<< pdiffusion >>
rect 304 286 305 287 
<< pdiffusion >>
rect 305 286 306 287 
<< m1 >>
rect 309 286 310 287 
<< m2 >>
rect 310 286 311 287 
<< pdiffusion >>
rect 318 286 319 287 
<< pdiffusion >>
rect 319 286 320 287 
<< pdiffusion >>
rect 320 286 321 287 
<< pdiffusion >>
rect 321 286 322 287 
<< pdiffusion >>
rect 322 286 323 287 
<< pdiffusion >>
rect 323 286 324 287 
<< m1 >>
rect 325 286 326 287 
<< pdiffusion >>
rect 336 286 337 287 
<< pdiffusion >>
rect 337 286 338 287 
<< pdiffusion >>
rect 338 286 339 287 
<< pdiffusion >>
rect 339 286 340 287 
<< pdiffusion >>
rect 340 286 341 287 
<< pdiffusion >>
rect 341 286 342 287 
<< m1 >>
rect 344 286 345 287 
<< m1 >>
rect 346 286 347 287 
<< m1 >>
rect 348 286 349 287 
<< m1 >>
rect 352 286 353 287 
<< pdiffusion >>
rect 354 286 355 287 
<< pdiffusion >>
rect 355 286 356 287 
<< pdiffusion >>
rect 356 286 357 287 
<< pdiffusion >>
rect 357 286 358 287 
<< pdiffusion >>
rect 358 286 359 287 
<< pdiffusion >>
rect 359 286 360 287 
<< m1 >>
rect 366 286 367 287 
<< m1 >>
rect 370 286 371 287 
<< pdiffusion >>
rect 372 286 373 287 
<< pdiffusion >>
rect 373 286 374 287 
<< pdiffusion >>
rect 374 286 375 287 
<< pdiffusion >>
rect 375 286 376 287 
<< pdiffusion >>
rect 376 286 377 287 
<< pdiffusion >>
rect 377 286 378 287 
<< m1 >>
rect 379 286 380 287 
<< m1 >>
rect 388 286 389 287 
<< pdiffusion >>
rect 390 286 391 287 
<< pdiffusion >>
rect 391 286 392 287 
<< pdiffusion >>
rect 392 286 393 287 
<< pdiffusion >>
rect 393 286 394 287 
<< pdiffusion >>
rect 394 286 395 287 
<< pdiffusion >>
rect 395 286 396 287 
<< m1 >>
rect 406 286 407 287 
<< pdiffusion >>
rect 408 286 409 287 
<< pdiffusion >>
rect 409 286 410 287 
<< pdiffusion >>
rect 410 286 411 287 
<< pdiffusion >>
rect 411 286 412 287 
<< pdiffusion >>
rect 412 286 413 287 
<< pdiffusion >>
rect 413 286 414 287 
<< m1 >>
rect 416 286 417 287 
<< m1 >>
rect 419 286 420 287 
<< m2 >>
rect 420 286 421 287 
<< pdiffusion >>
rect 426 286 427 287 
<< pdiffusion >>
rect 427 286 428 287 
<< pdiffusion >>
rect 428 286 429 287 
<< pdiffusion >>
rect 429 286 430 287 
<< pdiffusion >>
rect 430 286 431 287 
<< pdiffusion >>
rect 431 286 432 287 
<< m1 >>
rect 433 286 434 287 
<< m1 >>
rect 437 286 438 287 
<< pdiffusion >>
rect 444 286 445 287 
<< pdiffusion >>
rect 445 286 446 287 
<< pdiffusion >>
rect 446 286 447 287 
<< pdiffusion >>
rect 447 286 448 287 
<< pdiffusion >>
rect 448 286 449 287 
<< pdiffusion >>
rect 449 286 450 287 
<< pdiffusion >>
rect 462 286 463 287 
<< pdiffusion >>
rect 463 286 464 287 
<< pdiffusion >>
rect 464 286 465 287 
<< pdiffusion >>
rect 465 286 466 287 
<< pdiffusion >>
rect 466 286 467 287 
<< pdiffusion >>
rect 467 286 468 287 
<< pdiffusion >>
rect 480 286 481 287 
<< pdiffusion >>
rect 481 286 482 287 
<< pdiffusion >>
rect 482 286 483 287 
<< pdiffusion >>
rect 483 286 484 287 
<< pdiffusion >>
rect 484 286 485 287 
<< pdiffusion >>
rect 485 286 486 287 
<< m1 >>
rect 487 286 488 287 
<< pdiffusion >>
rect 498 286 499 287 
<< pdiffusion >>
rect 499 286 500 287 
<< pdiffusion >>
rect 500 286 501 287 
<< pdiffusion >>
rect 501 286 502 287 
<< pdiffusion >>
rect 502 286 503 287 
<< pdiffusion >>
rect 503 286 504 287 
<< pdiffusion >>
rect 516 286 517 287 
<< pdiffusion >>
rect 517 286 518 287 
<< pdiffusion >>
rect 518 286 519 287 
<< pdiffusion >>
rect 519 286 520 287 
<< pdiffusion >>
rect 520 286 521 287 
<< pdiffusion >>
rect 521 286 522 287 
<< m1 >>
rect 523 286 524 287 
<< pdiffusion >>
rect 12 287 13 288 
<< pdiffusion >>
rect 13 287 14 288 
<< pdiffusion >>
rect 14 287 15 288 
<< pdiffusion >>
rect 15 287 16 288 
<< pdiffusion >>
rect 16 287 17 288 
<< pdiffusion >>
rect 17 287 18 288 
<< m1 >>
rect 19 287 20 288 
<< m1 >>
rect 22 287 23 288 
<< pdiffusion >>
rect 30 287 31 288 
<< pdiffusion >>
rect 31 287 32 288 
<< pdiffusion >>
rect 32 287 33 288 
<< pdiffusion >>
rect 33 287 34 288 
<< pdiffusion >>
rect 34 287 35 288 
<< pdiffusion >>
rect 35 287 36 288 
<< m1 >>
rect 44 287 45 288 
<< pdiffusion >>
rect 48 287 49 288 
<< m1 >>
rect 49 287 50 288 
<< pdiffusion >>
rect 49 287 50 288 
<< pdiffusion >>
rect 50 287 51 288 
<< m1 >>
rect 51 287 52 288 
<< m2 >>
rect 51 287 52 288 
<< m2c >>
rect 51 287 52 288 
<< m1 >>
rect 51 287 52 288 
<< m2 >>
rect 51 287 52 288 
<< pdiffusion >>
rect 51 287 52 288 
<< m1 >>
rect 52 287 53 288 
<< pdiffusion >>
rect 52 287 53 288 
<< pdiffusion >>
rect 53 287 54 288 
<< m1 >>
rect 55 287 56 288 
<< m1 >>
rect 64 287 65 288 
<< pdiffusion >>
rect 66 287 67 288 
<< pdiffusion >>
rect 67 287 68 288 
<< pdiffusion >>
rect 68 287 69 288 
<< pdiffusion >>
rect 69 287 70 288 
<< pdiffusion >>
rect 70 287 71 288 
<< pdiffusion >>
rect 71 287 72 288 
<< m1 >>
rect 89 287 90 288 
<< m1 >>
rect 91 287 92 288 
<< pdiffusion >>
rect 102 287 103 288 
<< pdiffusion >>
rect 103 287 104 288 
<< pdiffusion >>
rect 104 287 105 288 
<< pdiffusion >>
rect 105 287 106 288 
<< pdiffusion >>
rect 106 287 107 288 
<< pdiffusion >>
rect 107 287 108 288 
<< m1 >>
rect 109 287 110 288 
<< pdiffusion >>
rect 120 287 121 288 
<< pdiffusion >>
rect 121 287 122 288 
<< pdiffusion >>
rect 122 287 123 288 
<< pdiffusion >>
rect 123 287 124 288 
<< pdiffusion >>
rect 124 287 125 288 
<< pdiffusion >>
rect 125 287 126 288 
<< pdiffusion >>
rect 138 287 139 288 
<< pdiffusion >>
rect 139 287 140 288 
<< pdiffusion >>
rect 140 287 141 288 
<< pdiffusion >>
rect 141 287 142 288 
<< pdiffusion >>
rect 142 287 143 288 
<< pdiffusion >>
rect 143 287 144 288 
<< m1 >>
rect 148 287 149 288 
<< m2 >>
rect 149 287 150 288 
<< m1 >>
rect 150 287 151 288 
<< m2 >>
rect 151 287 152 288 
<< pdiffusion >>
rect 156 287 157 288 
<< pdiffusion >>
rect 157 287 158 288 
<< pdiffusion >>
rect 158 287 159 288 
<< pdiffusion >>
rect 159 287 160 288 
<< m1 >>
rect 160 287 161 288 
<< pdiffusion >>
rect 160 287 161 288 
<< pdiffusion >>
rect 161 287 162 288 
<< m1 >>
rect 172 287 173 288 
<< pdiffusion >>
rect 174 287 175 288 
<< m1 >>
rect 175 287 176 288 
<< pdiffusion >>
rect 175 287 176 288 
<< pdiffusion >>
rect 176 287 177 288 
<< pdiffusion >>
rect 177 287 178 288 
<< pdiffusion >>
rect 178 287 179 288 
<< pdiffusion >>
rect 179 287 180 288 
<< m1 >>
rect 186 287 187 288 
<< pdiffusion >>
rect 192 287 193 288 
<< pdiffusion >>
rect 193 287 194 288 
<< pdiffusion >>
rect 194 287 195 288 
<< pdiffusion >>
rect 195 287 196 288 
<< pdiffusion >>
rect 196 287 197 288 
<< pdiffusion >>
rect 197 287 198 288 
<< pdiffusion >>
rect 210 287 211 288 
<< m1 >>
rect 211 287 212 288 
<< pdiffusion >>
rect 211 287 212 288 
<< pdiffusion >>
rect 212 287 213 288 
<< pdiffusion >>
rect 213 287 214 288 
<< pdiffusion >>
rect 214 287 215 288 
<< pdiffusion >>
rect 215 287 216 288 
<< m1 >>
rect 217 287 218 288 
<< m2 >>
rect 217 287 218 288 
<< m1 >>
rect 226 287 227 288 
<< pdiffusion >>
rect 228 287 229 288 
<< pdiffusion >>
rect 229 287 230 288 
<< pdiffusion >>
rect 230 287 231 288 
<< pdiffusion >>
rect 231 287 232 288 
<< m1 >>
rect 232 287 233 288 
<< pdiffusion >>
rect 232 287 233 288 
<< pdiffusion >>
rect 233 287 234 288 
<< m1 >>
rect 244 287 245 288 
<< pdiffusion >>
rect 246 287 247 288 
<< pdiffusion >>
rect 247 287 248 288 
<< pdiffusion >>
rect 248 287 249 288 
<< pdiffusion >>
rect 249 287 250 288 
<< m1 >>
rect 250 287 251 288 
<< pdiffusion >>
rect 250 287 251 288 
<< pdiffusion >>
rect 251 287 252 288 
<< m1 >>
rect 253 287 254 288 
<< m1 >>
rect 255 287 256 288 
<< m1 >>
rect 257 287 258 288 
<< m1 >>
rect 259 287 260 288 
<< pdiffusion >>
rect 264 287 265 288 
<< pdiffusion >>
rect 265 287 266 288 
<< pdiffusion >>
rect 266 287 267 288 
<< pdiffusion >>
rect 267 287 268 288 
<< m1 >>
rect 268 287 269 288 
<< pdiffusion >>
rect 268 287 269 288 
<< pdiffusion >>
rect 269 287 270 288 
<< m1 >>
rect 271 287 272 288 
<< m2 >>
rect 272 287 273 288 
<< m1 >>
rect 278 287 279 288 
<< m1 >>
rect 280 287 281 288 
<< pdiffusion >>
rect 282 287 283 288 
<< m1 >>
rect 283 287 284 288 
<< pdiffusion >>
rect 283 287 284 288 
<< pdiffusion >>
rect 284 287 285 288 
<< pdiffusion >>
rect 285 287 286 288 
<< pdiffusion >>
rect 286 287 287 288 
<< pdiffusion >>
rect 287 287 288 288 
<< m1 >>
rect 289 287 290 288 
<< m2 >>
rect 289 287 290 288 
<< pdiffusion >>
rect 300 287 301 288 
<< pdiffusion >>
rect 301 287 302 288 
<< pdiffusion >>
rect 302 287 303 288 
<< pdiffusion >>
rect 303 287 304 288 
<< m1 >>
rect 304 287 305 288 
<< pdiffusion >>
rect 304 287 305 288 
<< pdiffusion >>
rect 305 287 306 288 
<< m1 >>
rect 309 287 310 288 
<< m2 >>
rect 310 287 311 288 
<< pdiffusion >>
rect 318 287 319 288 
<< pdiffusion >>
rect 319 287 320 288 
<< pdiffusion >>
rect 320 287 321 288 
<< pdiffusion >>
rect 321 287 322 288 
<< pdiffusion >>
rect 322 287 323 288 
<< pdiffusion >>
rect 323 287 324 288 
<< m1 >>
rect 325 287 326 288 
<< pdiffusion >>
rect 336 287 337 288 
<< pdiffusion >>
rect 337 287 338 288 
<< pdiffusion >>
rect 338 287 339 288 
<< pdiffusion >>
rect 339 287 340 288 
<< m1 >>
rect 340 287 341 288 
<< pdiffusion >>
rect 340 287 341 288 
<< pdiffusion >>
rect 341 287 342 288 
<< m1 >>
rect 344 287 345 288 
<< m1 >>
rect 346 287 347 288 
<< m1 >>
rect 348 287 349 288 
<< m1 >>
rect 352 287 353 288 
<< pdiffusion >>
rect 354 287 355 288 
<< pdiffusion >>
rect 355 287 356 288 
<< pdiffusion >>
rect 356 287 357 288 
<< pdiffusion >>
rect 357 287 358 288 
<< pdiffusion >>
rect 358 287 359 288 
<< pdiffusion >>
rect 359 287 360 288 
<< m1 >>
rect 366 287 367 288 
<< m1 >>
rect 370 287 371 288 
<< pdiffusion >>
rect 372 287 373 288 
<< pdiffusion >>
rect 373 287 374 288 
<< pdiffusion >>
rect 374 287 375 288 
<< pdiffusion >>
rect 375 287 376 288 
<< pdiffusion >>
rect 376 287 377 288 
<< pdiffusion >>
rect 377 287 378 288 
<< m1 >>
rect 379 287 380 288 
<< m1 >>
rect 388 287 389 288 
<< pdiffusion >>
rect 390 287 391 288 
<< pdiffusion >>
rect 391 287 392 288 
<< pdiffusion >>
rect 392 287 393 288 
<< pdiffusion >>
rect 393 287 394 288 
<< pdiffusion >>
rect 394 287 395 288 
<< pdiffusion >>
rect 395 287 396 288 
<< m1 >>
rect 406 287 407 288 
<< pdiffusion >>
rect 408 287 409 288 
<< m1 >>
rect 409 287 410 288 
<< pdiffusion >>
rect 409 287 410 288 
<< pdiffusion >>
rect 410 287 411 288 
<< pdiffusion >>
rect 411 287 412 288 
<< m1 >>
rect 412 287 413 288 
<< pdiffusion >>
rect 412 287 413 288 
<< pdiffusion >>
rect 413 287 414 288 
<< m1 >>
rect 416 287 417 288 
<< m1 >>
rect 419 287 420 288 
<< m2 >>
rect 420 287 421 288 
<< pdiffusion >>
rect 426 287 427 288 
<< pdiffusion >>
rect 427 287 428 288 
<< pdiffusion >>
rect 428 287 429 288 
<< pdiffusion >>
rect 429 287 430 288 
<< m1 >>
rect 430 287 431 288 
<< pdiffusion >>
rect 430 287 431 288 
<< pdiffusion >>
rect 431 287 432 288 
<< m1 >>
rect 433 287 434 288 
<< m1 >>
rect 437 287 438 288 
<< pdiffusion >>
rect 444 287 445 288 
<< pdiffusion >>
rect 445 287 446 288 
<< pdiffusion >>
rect 446 287 447 288 
<< pdiffusion >>
rect 447 287 448 288 
<< pdiffusion >>
rect 448 287 449 288 
<< pdiffusion >>
rect 449 287 450 288 
<< pdiffusion >>
rect 462 287 463 288 
<< pdiffusion >>
rect 463 287 464 288 
<< pdiffusion >>
rect 464 287 465 288 
<< pdiffusion >>
rect 465 287 466 288 
<< pdiffusion >>
rect 466 287 467 288 
<< pdiffusion >>
rect 467 287 468 288 
<< pdiffusion >>
rect 480 287 481 288 
<< pdiffusion >>
rect 481 287 482 288 
<< pdiffusion >>
rect 482 287 483 288 
<< pdiffusion >>
rect 483 287 484 288 
<< pdiffusion >>
rect 484 287 485 288 
<< pdiffusion >>
rect 485 287 486 288 
<< m1 >>
rect 487 287 488 288 
<< pdiffusion >>
rect 498 287 499 288 
<< pdiffusion >>
rect 499 287 500 288 
<< pdiffusion >>
rect 500 287 501 288 
<< pdiffusion >>
rect 501 287 502 288 
<< pdiffusion >>
rect 502 287 503 288 
<< pdiffusion >>
rect 503 287 504 288 
<< pdiffusion >>
rect 516 287 517 288 
<< pdiffusion >>
rect 517 287 518 288 
<< pdiffusion >>
rect 518 287 519 288 
<< pdiffusion >>
rect 519 287 520 288 
<< pdiffusion >>
rect 520 287 521 288 
<< pdiffusion >>
rect 521 287 522 288 
<< m1 >>
rect 523 287 524 288 
<< m1 >>
rect 19 288 20 289 
<< m1 >>
rect 22 288 23 289 
<< m1 >>
rect 44 288 45 289 
<< m1 >>
rect 49 288 50 289 
<< m1 >>
rect 52 288 53 289 
<< m2 >>
rect 52 288 53 289 
<< m1 >>
rect 55 288 56 289 
<< m2 >>
rect 55 288 56 289 
<< m2c >>
rect 55 288 56 289 
<< m1 >>
rect 55 288 56 289 
<< m2 >>
rect 55 288 56 289 
<< m1 >>
rect 64 288 65 289 
<< m1 >>
rect 89 288 90 289 
<< m1 >>
rect 91 288 92 289 
<< m1 >>
rect 109 288 110 289 
<< m1 >>
rect 148 288 149 289 
<< m2 >>
rect 149 288 150 289 
<< m1 >>
rect 150 288 151 289 
<< m2 >>
rect 151 288 152 289 
<< m1 >>
rect 160 288 161 289 
<< m1 >>
rect 172 288 173 289 
<< m1 >>
rect 175 288 176 289 
<< m1 >>
rect 186 288 187 289 
<< m1 >>
rect 211 288 212 289 
<< m1 >>
rect 217 288 218 289 
<< m2 >>
rect 217 288 218 289 
<< m1 >>
rect 226 288 227 289 
<< m1 >>
rect 232 288 233 289 
<< m1 >>
rect 244 288 245 289 
<< m1 >>
rect 250 288 251 289 
<< m1 >>
rect 253 288 254 289 
<< m1 >>
rect 255 288 256 289 
<< m1 >>
rect 257 288 258 289 
<< m1 >>
rect 259 288 260 289 
<< m1 >>
rect 268 288 269 289 
<< m1 >>
rect 271 288 272 289 
<< m2 >>
rect 272 288 273 289 
<< m1 >>
rect 278 288 279 289 
<< m1 >>
rect 280 288 281 289 
<< m1 >>
rect 283 288 284 289 
<< m1 >>
rect 289 288 290 289 
<< m2 >>
rect 289 288 290 289 
<< m1 >>
rect 304 288 305 289 
<< m1 >>
rect 309 288 310 289 
<< m2 >>
rect 310 288 311 289 
<< m1 >>
rect 325 288 326 289 
<< m1 >>
rect 340 288 341 289 
<< m1 >>
rect 344 288 345 289 
<< m1 >>
rect 346 288 347 289 
<< m1 >>
rect 348 288 349 289 
<< m1 >>
rect 352 288 353 289 
<< m1 >>
rect 366 288 367 289 
<< m1 >>
rect 370 288 371 289 
<< m1 >>
rect 379 288 380 289 
<< m1 >>
rect 388 288 389 289 
<< m1 >>
rect 406 288 407 289 
<< m1 >>
rect 409 288 410 289 
<< m1 >>
rect 412 288 413 289 
<< m1 >>
rect 416 288 417 289 
<< m1 >>
rect 419 288 420 289 
<< m2 >>
rect 420 288 421 289 
<< m1 >>
rect 430 288 431 289 
<< m1 >>
rect 433 288 434 289 
<< m1 >>
rect 437 288 438 289 
<< m1 >>
rect 487 288 488 289 
<< m1 >>
rect 523 288 524 289 
<< m1 >>
rect 19 289 20 290 
<< m1 >>
rect 22 289 23 290 
<< m1 >>
rect 44 289 45 290 
<< m1 >>
rect 49 289 50 290 
<< m2 >>
rect 52 289 53 290 
<< m2 >>
rect 55 289 56 290 
<< m1 >>
rect 64 289 65 290 
<< m1 >>
rect 89 289 90 290 
<< m1 >>
rect 91 289 92 290 
<< m1 >>
rect 109 289 110 290 
<< m1 >>
rect 148 289 149 290 
<< m2 >>
rect 149 289 150 290 
<< m1 >>
rect 150 289 151 290 
<< m2 >>
rect 151 289 152 290 
<< m1 >>
rect 160 289 161 290 
<< m1 >>
rect 161 289 162 290 
<< m1 >>
rect 162 289 163 290 
<< m1 >>
rect 163 289 164 290 
<< m1 >>
rect 164 289 165 290 
<< m1 >>
rect 165 289 166 290 
<< m1 >>
rect 166 289 167 290 
<< m1 >>
rect 167 289 168 290 
<< m1 >>
rect 168 289 169 290 
<< m1 >>
rect 169 289 170 290 
<< m1 >>
rect 170 289 171 290 
<< m1 >>
rect 171 289 172 290 
<< m1 >>
rect 172 289 173 290 
<< m1 >>
rect 175 289 176 290 
<< m1 >>
rect 186 289 187 290 
<< m1 >>
rect 208 289 209 290 
<< m1 >>
rect 209 289 210 290 
<< m1 >>
rect 210 289 211 290 
<< m1 >>
rect 211 289 212 290 
<< m1 >>
rect 217 289 218 290 
<< m2 >>
rect 217 289 218 290 
<< m1 >>
rect 226 289 227 290 
<< m1 >>
rect 232 289 233 290 
<< m1 >>
rect 244 289 245 290 
<< m1 >>
rect 250 289 251 290 
<< m1 >>
rect 251 289 252 290 
<< m1 >>
rect 252 289 253 290 
<< m1 >>
rect 253 289 254 290 
<< m1 >>
rect 255 289 256 290 
<< m1 >>
rect 257 289 258 290 
<< m1 >>
rect 259 289 260 290 
<< m1 >>
rect 268 289 269 290 
<< m1 >>
rect 269 289 270 290 
<< m2 >>
rect 269 289 270 290 
<< m2c >>
rect 269 289 270 290 
<< m1 >>
rect 269 289 270 290 
<< m2 >>
rect 269 289 270 290 
<< m2 >>
rect 270 289 271 290 
<< m1 >>
rect 271 289 272 290 
<< m2 >>
rect 271 289 272 290 
<< m2 >>
rect 272 289 273 290 
<< m1 >>
rect 278 289 279 290 
<< m1 >>
rect 280 289 281 290 
<< m1 >>
rect 283 289 284 290 
<< m1 >>
rect 284 289 285 290 
<< m1 >>
rect 289 289 290 290 
<< m2 >>
rect 289 289 290 290 
<< m1 >>
rect 304 289 305 290 
<< m1 >>
rect 305 289 306 290 
<< m1 >>
rect 306 289 307 290 
<< m1 >>
rect 307 289 308 290 
<< m1 >>
rect 309 289 310 290 
<< m2 >>
rect 310 289 311 290 
<< m1 >>
rect 325 289 326 290 
<< m1 >>
rect 340 289 341 290 
<< m1 >>
rect 344 289 345 290 
<< m1 >>
rect 346 289 347 290 
<< m1 >>
rect 348 289 349 290 
<< m1 >>
rect 352 289 353 290 
<< m1 >>
rect 366 289 367 290 
<< m1 >>
rect 370 289 371 290 
<< m1 >>
rect 379 289 380 290 
<< m1 >>
rect 388 289 389 290 
<< m1 >>
rect 406 289 407 290 
<< m1 >>
rect 407 289 408 290 
<< m2 >>
rect 407 289 408 290 
<< m2c >>
rect 407 289 408 290 
<< m1 >>
rect 407 289 408 290 
<< m2 >>
rect 407 289 408 290 
<< m2 >>
rect 408 289 409 290 
<< m1 >>
rect 409 289 410 290 
<< m1 >>
rect 412 289 413 290 
<< m1 >>
rect 413 289 414 290 
<< m1 >>
rect 414 289 415 290 
<< m2 >>
rect 414 289 415 290 
<< m2c >>
rect 414 289 415 290 
<< m1 >>
rect 414 289 415 290 
<< m2 >>
rect 414 289 415 290 
<< m2 >>
rect 415 289 416 290 
<< m1 >>
rect 416 289 417 290 
<< m2 >>
rect 416 289 417 290 
<< m2 >>
rect 417 289 418 290 
<< m2 >>
rect 418 289 419 290 
<< m1 >>
rect 419 289 420 290 
<< m2 >>
rect 419 289 420 290 
<< m2 >>
rect 420 289 421 290 
<< m1 >>
rect 430 289 431 290 
<< m1 >>
rect 433 289 434 290 
<< m1 >>
rect 437 289 438 290 
<< m1 >>
rect 487 289 488 290 
<< m1 >>
rect 523 289 524 290 
<< m1 >>
rect 19 290 20 291 
<< m1 >>
rect 22 290 23 291 
<< m1 >>
rect 44 290 45 291 
<< m1 >>
rect 49 290 50 291 
<< m1 >>
rect 50 290 51 291 
<< m1 >>
rect 51 290 52 291 
<< m1 >>
rect 52 290 53 291 
<< m2 >>
rect 52 290 53 291 
<< m1 >>
rect 53 290 54 291 
<< m1 >>
rect 54 290 55 291 
<< m1 >>
rect 55 290 56 291 
<< m2 >>
rect 55 290 56 291 
<< m1 >>
rect 56 290 57 291 
<< m1 >>
rect 57 290 58 291 
<< m1 >>
rect 58 290 59 291 
<< m1 >>
rect 59 290 60 291 
<< m1 >>
rect 60 290 61 291 
<< m1 >>
rect 61 290 62 291 
<< m1 >>
rect 62 290 63 291 
<< m1 >>
rect 63 290 64 291 
<< m1 >>
rect 64 290 65 291 
<< m1 >>
rect 89 290 90 291 
<< m1 >>
rect 91 290 92 291 
<< m1 >>
rect 109 290 110 291 
<< m1 >>
rect 148 290 149 291 
<< m2 >>
rect 149 290 150 291 
<< m1 >>
rect 150 290 151 291 
<< m2 >>
rect 151 290 152 291 
<< m1 >>
rect 175 290 176 291 
<< m1 >>
rect 186 290 187 291 
<< m1 >>
rect 208 290 209 291 
<< m1 >>
rect 217 290 218 291 
<< m2 >>
rect 217 290 218 291 
<< m1 >>
rect 226 290 227 291 
<< m1 >>
rect 232 290 233 291 
<< m1 >>
rect 244 290 245 291 
<< m2 >>
rect 249 290 250 291 
<< m2 >>
rect 250 290 251 291 
<< m2 >>
rect 251 290 252 291 
<< m2 >>
rect 252 290 253 291 
<< m2 >>
rect 253 290 254 291 
<< m2 >>
rect 254 290 255 291 
<< m1 >>
rect 255 290 256 291 
<< m2 >>
rect 255 290 256 291 
<< m2 >>
rect 256 290 257 291 
<< m1 >>
rect 257 290 258 291 
<< m2 >>
rect 257 290 258 291 
<< m2 >>
rect 258 290 259 291 
<< m1 >>
rect 259 290 260 291 
<< m2 >>
rect 259 290 260 291 
<< m2c >>
rect 259 290 260 291 
<< m1 >>
rect 259 290 260 291 
<< m2 >>
rect 259 290 260 291 
<< m1 >>
rect 271 290 272 291 
<< m1 >>
rect 278 290 279 291 
<< m1 >>
rect 280 290 281 291 
<< m1 >>
rect 284 290 285 291 
<< m2 >>
rect 284 290 285 291 
<< m2c >>
rect 284 290 285 291 
<< m1 >>
rect 284 290 285 291 
<< m2 >>
rect 284 290 285 291 
<< m1 >>
rect 289 290 290 291 
<< m2 >>
rect 289 290 290 291 
<< m1 >>
rect 307 290 308 291 
<< m1 >>
rect 309 290 310 291 
<< m2 >>
rect 310 290 311 291 
<< m1 >>
rect 325 290 326 291 
<< m1 >>
rect 340 290 341 291 
<< m1 >>
rect 344 290 345 291 
<< m1 >>
rect 346 290 347 291 
<< m1 >>
rect 348 290 349 291 
<< m1 >>
rect 352 290 353 291 
<< m1 >>
rect 366 290 367 291 
<< m1 >>
rect 370 290 371 291 
<< m1 >>
rect 379 290 380 291 
<< m1 >>
rect 388 290 389 291 
<< m2 >>
rect 408 290 409 291 
<< m1 >>
rect 409 290 410 291 
<< m1 >>
rect 416 290 417 291 
<< m1 >>
rect 419 290 420 291 
<< m1 >>
rect 430 290 431 291 
<< m1 >>
rect 433 290 434 291 
<< m1 >>
rect 437 290 438 291 
<< m1 >>
rect 487 290 488 291 
<< m1 >>
rect 523 290 524 291 
<< m1 >>
rect 19 291 20 292 
<< m1 >>
rect 22 291 23 292 
<< m1 >>
rect 44 291 45 292 
<< m2 >>
rect 52 291 53 292 
<< m2 >>
rect 55 291 56 292 
<< m1 >>
rect 89 291 90 292 
<< m1 >>
rect 91 291 92 292 
<< m1 >>
rect 109 291 110 292 
<< m1 >>
rect 148 291 149 292 
<< m2 >>
rect 149 291 150 292 
<< m1 >>
rect 150 291 151 292 
<< m2 >>
rect 151 291 152 292 
<< m1 >>
rect 175 291 176 292 
<< m1 >>
rect 186 291 187 292 
<< m1 >>
rect 208 291 209 292 
<< m1 >>
rect 217 291 218 292 
<< m2 >>
rect 217 291 218 292 
<< m1 >>
rect 226 291 227 292 
<< m1 >>
rect 232 291 233 292 
<< m1 >>
rect 244 291 245 292 
<< m1 >>
rect 249 291 250 292 
<< m2 >>
rect 249 291 250 292 
<< m2c >>
rect 249 291 250 292 
<< m1 >>
rect 249 291 250 292 
<< m2 >>
rect 249 291 250 292 
<< m1 >>
rect 255 291 256 292 
<< m1 >>
rect 257 291 258 292 
<< m1 >>
rect 271 291 272 292 
<< m1 >>
rect 278 291 279 292 
<< m1 >>
rect 280 291 281 292 
<< m2 >>
rect 284 291 285 292 
<< m1 >>
rect 289 291 290 292 
<< m2 >>
rect 289 291 290 292 
<< m1 >>
rect 307 291 308 292 
<< m1 >>
rect 309 291 310 292 
<< m2 >>
rect 310 291 311 292 
<< m1 >>
rect 325 291 326 292 
<< m1 >>
rect 340 291 341 292 
<< m1 >>
rect 344 291 345 292 
<< m1 >>
rect 346 291 347 292 
<< m1 >>
rect 348 291 349 292 
<< m1 >>
rect 352 291 353 292 
<< m1 >>
rect 366 291 367 292 
<< m1 >>
rect 370 291 371 292 
<< m1 >>
rect 379 291 380 292 
<< m1 >>
rect 388 291 389 292 
<< m2 >>
rect 408 291 409 292 
<< m1 >>
rect 409 291 410 292 
<< m1 >>
rect 416 291 417 292 
<< m1 >>
rect 419 291 420 292 
<< m1 >>
rect 430 291 431 292 
<< m1 >>
rect 433 291 434 292 
<< m1 >>
rect 437 291 438 292 
<< m1 >>
rect 487 291 488 292 
<< m1 >>
rect 523 291 524 292 
<< m1 >>
rect 19 292 20 293 
<< m1 >>
rect 22 292 23 293 
<< m1 >>
rect 44 292 45 293 
<< m1 >>
rect 46 292 47 293 
<< m1 >>
rect 47 292 48 293 
<< m1 >>
rect 48 292 49 293 
<< m1 >>
rect 49 292 50 293 
<< m1 >>
rect 50 292 51 293 
<< m1 >>
rect 51 292 52 293 
<< m1 >>
rect 52 292 53 293 
<< m2 >>
rect 52 292 53 293 
<< m2c >>
rect 52 292 53 293 
<< m1 >>
rect 52 292 53 293 
<< m2 >>
rect 52 292 53 293 
<< m1 >>
rect 55 292 56 293 
<< m2 >>
rect 55 292 56 293 
<< m2c >>
rect 55 292 56 293 
<< m1 >>
rect 55 292 56 293 
<< m2 >>
rect 55 292 56 293 
<< m1 >>
rect 89 292 90 293 
<< m1 >>
rect 91 292 92 293 
<< m1 >>
rect 93 292 94 293 
<< m1 >>
rect 94 292 95 293 
<< m1 >>
rect 95 292 96 293 
<< m1 >>
rect 96 292 97 293 
<< m1 >>
rect 97 292 98 293 
<< m1 >>
rect 98 292 99 293 
<< m1 >>
rect 99 292 100 293 
<< m1 >>
rect 100 292 101 293 
<< m1 >>
rect 101 292 102 293 
<< m1 >>
rect 102 292 103 293 
<< m1 >>
rect 103 292 104 293 
<< m1 >>
rect 104 292 105 293 
<< m1 >>
rect 105 292 106 293 
<< m1 >>
rect 106 292 107 293 
<< m1 >>
rect 107 292 108 293 
<< m1 >>
rect 108 292 109 293 
<< m1 >>
rect 109 292 110 293 
<< m1 >>
rect 148 292 149 293 
<< m2 >>
rect 149 292 150 293 
<< m1 >>
rect 150 292 151 293 
<< m2 >>
rect 151 292 152 293 
<< m1 >>
rect 175 292 176 293 
<< m1 >>
rect 186 292 187 293 
<< m1 >>
rect 208 292 209 293 
<< m1 >>
rect 217 292 218 293 
<< m2 >>
rect 217 292 218 293 
<< m1 >>
rect 226 292 227 293 
<< m1 >>
rect 232 292 233 293 
<< m1 >>
rect 244 292 245 293 
<< m1 >>
rect 249 292 250 293 
<< m1 >>
rect 255 292 256 293 
<< m1 >>
rect 257 292 258 293 
<< m1 >>
rect 258 292 259 293 
<< m1 >>
rect 259 292 260 293 
<< m1 >>
rect 260 292 261 293 
<< m1 >>
rect 261 292 262 293 
<< m1 >>
rect 262 292 263 293 
<< m1 >>
rect 263 292 264 293 
<< m1 >>
rect 264 292 265 293 
<< m1 >>
rect 265 292 266 293 
<< m1 >>
rect 266 292 267 293 
<< m1 >>
rect 267 292 268 293 
<< m1 >>
rect 268 292 269 293 
<< m1 >>
rect 269 292 270 293 
<< m2 >>
rect 269 292 270 293 
<< m2c >>
rect 269 292 270 293 
<< m1 >>
rect 269 292 270 293 
<< m2 >>
rect 269 292 270 293 
<< m2 >>
rect 270 292 271 293 
<< m1 >>
rect 271 292 272 293 
<< m2 >>
rect 271 292 272 293 
<< m2 >>
rect 272 292 273 293 
<< m1 >>
rect 273 292 274 293 
<< m2 >>
rect 273 292 274 293 
<< m2c >>
rect 273 292 274 293 
<< m1 >>
rect 273 292 274 293 
<< m2 >>
rect 273 292 274 293 
<< m1 >>
rect 274 292 275 293 
<< m1 >>
rect 275 292 276 293 
<< m1 >>
rect 276 292 277 293 
<< m2 >>
rect 276 292 277 293 
<< m2c >>
rect 276 292 277 293 
<< m1 >>
rect 276 292 277 293 
<< m2 >>
rect 276 292 277 293 
<< m2 >>
rect 277 292 278 293 
<< m1 >>
rect 278 292 279 293 
<< m2 >>
rect 278 292 279 293 
<< m2 >>
rect 279 292 280 293 
<< m1 >>
rect 280 292 281 293 
<< m2 >>
rect 280 292 281 293 
<< m2 >>
rect 281 292 282 293 
<< m1 >>
rect 282 292 283 293 
<< m2 >>
rect 282 292 283 293 
<< m2c >>
rect 282 292 283 293 
<< m1 >>
rect 282 292 283 293 
<< m2 >>
rect 282 292 283 293 
<< m1 >>
rect 283 292 284 293 
<< m1 >>
rect 284 292 285 293 
<< m2 >>
rect 284 292 285 293 
<< m1 >>
rect 285 292 286 293 
<< m1 >>
rect 286 292 287 293 
<< m1 >>
rect 287 292 288 293 
<< m2 >>
rect 287 292 288 293 
<< m2c >>
rect 287 292 288 293 
<< m1 >>
rect 287 292 288 293 
<< m2 >>
rect 287 292 288 293 
<< m2 >>
rect 288 292 289 293 
<< m1 >>
rect 289 292 290 293 
<< m2 >>
rect 289 292 290 293 
<< m1 >>
rect 307 292 308 293 
<< m1 >>
rect 309 292 310 293 
<< m2 >>
rect 310 292 311 293 
<< m1 >>
rect 325 292 326 293 
<< m1 >>
rect 326 292 327 293 
<< m1 >>
rect 327 292 328 293 
<< m1 >>
rect 328 292 329 293 
<< m1 >>
rect 329 292 330 293 
<< m1 >>
rect 330 292 331 293 
<< m1 >>
rect 331 292 332 293 
<< m1 >>
rect 332 292 333 293 
<< m1 >>
rect 333 292 334 293 
<< m1 >>
rect 334 292 335 293 
<< m1 >>
rect 335 292 336 293 
<< m1 >>
rect 336 292 337 293 
<< m1 >>
rect 337 292 338 293 
<< m1 >>
rect 338 292 339 293 
<< m2 >>
rect 338 292 339 293 
<< m2c >>
rect 338 292 339 293 
<< m1 >>
rect 338 292 339 293 
<< m2 >>
rect 338 292 339 293 
<< m2 >>
rect 339 292 340 293 
<< m1 >>
rect 340 292 341 293 
<< m2 >>
rect 340 292 341 293 
<< m2 >>
rect 341 292 342 293 
<< m1 >>
rect 342 292 343 293 
<< m2 >>
rect 342 292 343 293 
<< m2c >>
rect 342 292 343 293 
<< m1 >>
rect 342 292 343 293 
<< m2 >>
rect 342 292 343 293 
<< m2 >>
rect 343 292 344 293 
<< m1 >>
rect 344 292 345 293 
<< m2 >>
rect 344 292 345 293 
<< m2 >>
rect 345 292 346 293 
<< m1 >>
rect 346 292 347 293 
<< m2 >>
rect 346 292 347 293 
<< m2c >>
rect 346 292 347 293 
<< m1 >>
rect 346 292 347 293 
<< m2 >>
rect 346 292 347 293 
<< m1 >>
rect 348 292 349 293 
<< m1 >>
rect 352 292 353 293 
<< m1 >>
rect 366 292 367 293 
<< m1 >>
rect 370 292 371 293 
<< m1 >>
rect 379 292 380 293 
<< m1 >>
rect 388 292 389 293 
<< m1 >>
rect 389 292 390 293 
<< m1 >>
rect 390 292 391 293 
<< m1 >>
rect 391 292 392 293 
<< m1 >>
rect 392 292 393 293 
<< m1 >>
rect 393 292 394 293 
<< m1 >>
rect 394 292 395 293 
<< m2 >>
rect 408 292 409 293 
<< m1 >>
rect 409 292 410 293 
<< m2 >>
rect 409 292 410 293 
<< m2 >>
rect 410 292 411 293 
<< m1 >>
rect 411 292 412 293 
<< m2 >>
rect 411 292 412 293 
<< m2c >>
rect 411 292 412 293 
<< m1 >>
rect 411 292 412 293 
<< m2 >>
rect 411 292 412 293 
<< m1 >>
rect 412 292 413 293 
<< m1 >>
rect 413 292 414 293 
<< m1 >>
rect 414 292 415 293 
<< m2 >>
rect 414 292 415 293 
<< m2c >>
rect 414 292 415 293 
<< m1 >>
rect 414 292 415 293 
<< m2 >>
rect 414 292 415 293 
<< m2 >>
rect 415 292 416 293 
<< m1 >>
rect 416 292 417 293 
<< m1 >>
rect 419 292 420 293 
<< m1 >>
rect 430 292 431 293 
<< m1 >>
rect 433 292 434 293 
<< m1 >>
rect 437 292 438 293 
<< m1 >>
rect 487 292 488 293 
<< m1 >>
rect 523 292 524 293 
<< m1 >>
rect 19 293 20 294 
<< m1 >>
rect 22 293 23 294 
<< m1 >>
rect 44 293 45 294 
<< m1 >>
rect 46 293 47 294 
<< m1 >>
rect 55 293 56 294 
<< m1 >>
rect 89 293 90 294 
<< m2 >>
rect 89 293 90 294 
<< m2c >>
rect 89 293 90 294 
<< m1 >>
rect 89 293 90 294 
<< m2 >>
rect 89 293 90 294 
<< m1 >>
rect 91 293 92 294 
<< m2 >>
rect 91 293 92 294 
<< m2c >>
rect 91 293 92 294 
<< m1 >>
rect 91 293 92 294 
<< m2 >>
rect 91 293 92 294 
<< m1 >>
rect 93 293 94 294 
<< m2 >>
rect 93 293 94 294 
<< m2c >>
rect 93 293 94 294 
<< m1 >>
rect 93 293 94 294 
<< m2 >>
rect 93 293 94 294 
<< m2 >>
rect 146 293 147 294 
<< m2 >>
rect 147 293 148 294 
<< m1 >>
rect 148 293 149 294 
<< m2 >>
rect 148 293 149 294 
<< m2 >>
rect 149 293 150 294 
<< m1 >>
rect 150 293 151 294 
<< m2 >>
rect 151 293 152 294 
<< m1 >>
rect 175 293 176 294 
<< m1 >>
rect 186 293 187 294 
<< m1 >>
rect 208 293 209 294 
<< m1 >>
rect 217 293 218 294 
<< m2 >>
rect 217 293 218 294 
<< m1 >>
rect 226 293 227 294 
<< m1 >>
rect 232 293 233 294 
<< m1 >>
rect 244 293 245 294 
<< m1 >>
rect 249 293 250 294 
<< m1 >>
rect 255 293 256 294 
<< m1 >>
rect 271 293 272 294 
<< m1 >>
rect 278 293 279 294 
<< m1 >>
rect 280 293 281 294 
<< m2 >>
rect 284 293 285 294 
<< m1 >>
rect 289 293 290 294 
<< m1 >>
rect 307 293 308 294 
<< m1 >>
rect 309 293 310 294 
<< m2 >>
rect 310 293 311 294 
<< m1 >>
rect 340 293 341 294 
<< m1 >>
rect 344 293 345 294 
<< m1 >>
rect 348 293 349 294 
<< m1 >>
rect 352 293 353 294 
<< m1 >>
rect 366 293 367 294 
<< m1 >>
rect 367 293 368 294 
<< m1 >>
rect 368 293 369 294 
<< m2 >>
rect 368 293 369 294 
<< m2c >>
rect 368 293 369 294 
<< m1 >>
rect 368 293 369 294 
<< m2 >>
rect 368 293 369 294 
<< m2 >>
rect 369 293 370 294 
<< m1 >>
rect 370 293 371 294 
<< m2 >>
rect 370 293 371 294 
<< m2 >>
rect 371 293 372 294 
<< m1 >>
rect 372 293 373 294 
<< m2 >>
rect 372 293 373 294 
<< m2c >>
rect 372 293 373 294 
<< m1 >>
rect 372 293 373 294 
<< m2 >>
rect 372 293 373 294 
<< m1 >>
rect 373 293 374 294 
<< m1 >>
rect 374 293 375 294 
<< m1 >>
rect 375 293 376 294 
<< m1 >>
rect 376 293 377 294 
<< m1 >>
rect 377 293 378 294 
<< m2 >>
rect 377 293 378 294 
<< m2c >>
rect 377 293 378 294 
<< m1 >>
rect 377 293 378 294 
<< m2 >>
rect 377 293 378 294 
<< m2 >>
rect 378 293 379 294 
<< m1 >>
rect 379 293 380 294 
<< m2 >>
rect 379 293 380 294 
<< m2 >>
rect 380 293 381 294 
<< m1 >>
rect 394 293 395 294 
<< m1 >>
rect 409 293 410 294 
<< m2 >>
rect 415 293 416 294 
<< m1 >>
rect 416 293 417 294 
<< m1 >>
rect 419 293 420 294 
<< m2 >>
rect 419 293 420 294 
<< m2c >>
rect 419 293 420 294 
<< m1 >>
rect 419 293 420 294 
<< m2 >>
rect 419 293 420 294 
<< m1 >>
rect 430 293 431 294 
<< m1 >>
rect 433 293 434 294 
<< m1 >>
rect 437 293 438 294 
<< m1 >>
rect 487 293 488 294 
<< m1 >>
rect 523 293 524 294 
<< m1 >>
rect 19 294 20 295 
<< m1 >>
rect 22 294 23 295 
<< m1 >>
rect 44 294 45 295 
<< m1 >>
rect 46 294 47 295 
<< m1 >>
rect 55 294 56 295 
<< m2 >>
rect 74 294 75 295 
<< m2 >>
rect 75 294 76 295 
<< m2 >>
rect 76 294 77 295 
<< m2 >>
rect 77 294 78 295 
<< m2 >>
rect 78 294 79 295 
<< m2 >>
rect 79 294 80 295 
<< m2 >>
rect 80 294 81 295 
<< m2 >>
rect 81 294 82 295 
<< m2 >>
rect 82 294 83 295 
<< m2 >>
rect 83 294 84 295 
<< m2 >>
rect 84 294 85 295 
<< m2 >>
rect 85 294 86 295 
<< m2 >>
rect 86 294 87 295 
<< m2 >>
rect 87 294 88 295 
<< m2 >>
rect 88 294 89 295 
<< m2 >>
rect 89 294 90 295 
<< m2 >>
rect 91 294 92 295 
<< m2 >>
rect 93 294 94 295 
<< m2 >>
rect 107 294 108 295 
<< m1 >>
rect 108 294 109 295 
<< m2 >>
rect 108 294 109 295 
<< m2c >>
rect 108 294 109 295 
<< m1 >>
rect 108 294 109 295 
<< m2 >>
rect 108 294 109 295 
<< m1 >>
rect 109 294 110 295 
<< m1 >>
rect 110 294 111 295 
<< m1 >>
rect 111 294 112 295 
<< m1 >>
rect 112 294 113 295 
<< m1 >>
rect 113 294 114 295 
<< m1 >>
rect 114 294 115 295 
<< m1 >>
rect 115 294 116 295 
<< m1 >>
rect 116 294 117 295 
<< m1 >>
rect 117 294 118 295 
<< m1 >>
rect 118 294 119 295 
<< m1 >>
rect 119 294 120 295 
<< m1 >>
rect 120 294 121 295 
<< m1 >>
rect 121 294 122 295 
<< m1 >>
rect 122 294 123 295 
<< m1 >>
rect 123 294 124 295 
<< m1 >>
rect 124 294 125 295 
<< m1 >>
rect 125 294 126 295 
<< m1 >>
rect 126 294 127 295 
<< m1 >>
rect 127 294 128 295 
<< m1 >>
rect 128 294 129 295 
<< m1 >>
rect 129 294 130 295 
<< m1 >>
rect 130 294 131 295 
<< m1 >>
rect 131 294 132 295 
<< m1 >>
rect 132 294 133 295 
<< m1 >>
rect 133 294 134 295 
<< m1 >>
rect 134 294 135 295 
<< m1 >>
rect 135 294 136 295 
<< m1 >>
rect 136 294 137 295 
<< m1 >>
rect 137 294 138 295 
<< m1 >>
rect 138 294 139 295 
<< m1 >>
rect 139 294 140 295 
<< m1 >>
rect 140 294 141 295 
<< m1 >>
rect 141 294 142 295 
<< m1 >>
rect 142 294 143 295 
<< m1 >>
rect 143 294 144 295 
<< m1 >>
rect 144 294 145 295 
<< m1 >>
rect 145 294 146 295 
<< m1 >>
rect 146 294 147 295 
<< m2 >>
rect 146 294 147 295 
<< m1 >>
rect 147 294 148 295 
<< m1 >>
rect 148 294 149 295 
<< m1 >>
rect 150 294 151 295 
<< m2 >>
rect 151 294 152 295 
<< m1 >>
rect 175 294 176 295 
<< m1 >>
rect 186 294 187 295 
<< m1 >>
rect 208 294 209 295 
<< m1 >>
rect 217 294 218 295 
<< m2 >>
rect 217 294 218 295 
<< m1 >>
rect 226 294 227 295 
<< m1 >>
rect 232 294 233 295 
<< m1 >>
rect 244 294 245 295 
<< m1 >>
rect 249 294 250 295 
<< m1 >>
rect 255 294 256 295 
<< m1 >>
rect 271 294 272 295 
<< m1 >>
rect 278 294 279 295 
<< m1 >>
rect 280 294 281 295 
<< m2 >>
rect 284 294 285 295 
<< m1 >>
rect 289 294 290 295 
<< m1 >>
rect 307 294 308 295 
<< m1 >>
rect 309 294 310 295 
<< m2 >>
rect 310 294 311 295 
<< m1 >>
rect 340 294 341 295 
<< m1 >>
rect 344 294 345 295 
<< m1 >>
rect 348 294 349 295 
<< m1 >>
rect 352 294 353 295 
<< m1 >>
rect 370 294 371 295 
<< m1 >>
rect 379 294 380 295 
<< m2 >>
rect 380 294 381 295 
<< m1 >>
rect 394 294 395 295 
<< m1 >>
rect 409 294 410 295 
<< m2 >>
rect 415 294 416 295 
<< m1 >>
rect 416 294 417 295 
<< m2 >>
rect 419 294 420 295 
<< m1 >>
rect 430 294 431 295 
<< m1 >>
rect 433 294 434 295 
<< m1 >>
rect 437 294 438 295 
<< m1 >>
rect 487 294 488 295 
<< m1 >>
rect 523 294 524 295 
<< m1 >>
rect 19 295 20 296 
<< m1 >>
rect 22 295 23 296 
<< m1 >>
rect 44 295 45 296 
<< m1 >>
rect 46 295 47 296 
<< m1 >>
rect 55 295 56 296 
<< m1 >>
rect 73 295 74 296 
<< m1 >>
rect 74 295 75 296 
<< m2 >>
rect 74 295 75 296 
<< m1 >>
rect 75 295 76 296 
<< m1 >>
rect 76 295 77 296 
<< m1 >>
rect 77 295 78 296 
<< m1 >>
rect 78 295 79 296 
<< m1 >>
rect 79 295 80 296 
<< m1 >>
rect 80 295 81 296 
<< m1 >>
rect 81 295 82 296 
<< m1 >>
rect 82 295 83 296 
<< m1 >>
rect 83 295 84 296 
<< m1 >>
rect 84 295 85 296 
<< m1 >>
rect 85 295 86 296 
<< m1 >>
rect 86 295 87 296 
<< m1 >>
rect 87 295 88 296 
<< m1 >>
rect 88 295 89 296 
<< m1 >>
rect 89 295 90 296 
<< m1 >>
rect 90 295 91 296 
<< m1 >>
rect 91 295 92 296 
<< m2 >>
rect 91 295 92 296 
<< m1 >>
rect 92 295 93 296 
<< m1 >>
rect 93 295 94 296 
<< m2 >>
rect 93 295 94 296 
<< m1 >>
rect 94 295 95 296 
<< m1 >>
rect 95 295 96 296 
<< m1 >>
rect 96 295 97 296 
<< m1 >>
rect 97 295 98 296 
<< m1 >>
rect 98 295 99 296 
<< m1 >>
rect 99 295 100 296 
<< m1 >>
rect 100 295 101 296 
<< m1 >>
rect 101 295 102 296 
<< m1 >>
rect 102 295 103 296 
<< m1 >>
rect 103 295 104 296 
<< m1 >>
rect 104 295 105 296 
<< m1 >>
rect 105 295 106 296 
<< m1 >>
rect 106 295 107 296 
<< m2 >>
rect 107 295 108 296 
<< m2 >>
rect 146 295 147 296 
<< m1 >>
rect 150 295 151 296 
<< m2 >>
rect 151 295 152 296 
<< m1 >>
rect 175 295 176 296 
<< m1 >>
rect 176 295 177 296 
<< m1 >>
rect 177 295 178 296 
<< m1 >>
rect 178 295 179 296 
<< m1 >>
rect 179 295 180 296 
<< m1 >>
rect 180 295 181 296 
<< m1 >>
rect 181 295 182 296 
<< m1 >>
rect 186 295 187 296 
<< m1 >>
rect 208 295 209 296 
<< m1 >>
rect 217 295 218 296 
<< m2 >>
rect 217 295 218 296 
<< m1 >>
rect 226 295 227 296 
<< m1 >>
rect 232 295 233 296 
<< m1 >>
rect 244 295 245 296 
<< m1 >>
rect 246 295 247 296 
<< m1 >>
rect 247 295 248 296 
<< m1 >>
rect 248 295 249 296 
<< m1 >>
rect 249 295 250 296 
<< m1 >>
rect 255 295 256 296 
<< m1 >>
rect 271 295 272 296 
<< m1 >>
rect 278 295 279 296 
<< m1 >>
rect 280 295 281 296 
<< m1 >>
rect 282 295 283 296 
<< m1 >>
rect 283 295 284 296 
<< m1 >>
rect 284 295 285 296 
<< m2 >>
rect 284 295 285 296 
<< m1 >>
rect 285 295 286 296 
<< m1 >>
rect 286 295 287 296 
<< m1 >>
rect 287 295 288 296 
<< m1 >>
rect 288 295 289 296 
<< m1 >>
rect 289 295 290 296 
<< m1 >>
rect 307 295 308 296 
<< m1 >>
rect 309 295 310 296 
<< m2 >>
rect 310 295 311 296 
<< m2 >>
rect 333 295 334 296 
<< m1 >>
rect 334 295 335 296 
<< m2 >>
rect 334 295 335 296 
<< m1 >>
rect 335 295 336 296 
<< m2 >>
rect 335 295 336 296 
<< m1 >>
rect 336 295 337 296 
<< m2 >>
rect 336 295 337 296 
<< m1 >>
rect 337 295 338 296 
<< m2 >>
rect 337 295 338 296 
<< m1 >>
rect 338 295 339 296 
<< m2 >>
rect 338 295 339 296 
<< m1 >>
rect 339 295 340 296 
<< m2 >>
rect 339 295 340 296 
<< m1 >>
rect 340 295 341 296 
<< m2 >>
rect 340 295 341 296 
<< m2 >>
rect 341 295 342 296 
<< m1 >>
rect 342 295 343 296 
<< m2 >>
rect 342 295 343 296 
<< m2c >>
rect 342 295 343 296 
<< m1 >>
rect 342 295 343 296 
<< m2 >>
rect 342 295 343 296 
<< m2 >>
rect 343 295 344 296 
<< m1 >>
rect 344 295 345 296 
<< m2 >>
rect 344 295 345 296 
<< m2 >>
rect 345 295 346 296 
<< m1 >>
rect 346 295 347 296 
<< m2 >>
rect 346 295 347 296 
<< m2c >>
rect 346 295 347 296 
<< m1 >>
rect 346 295 347 296 
<< m2 >>
rect 346 295 347 296 
<< m2 >>
rect 347 295 348 296 
<< m1 >>
rect 348 295 349 296 
<< m2 >>
rect 348 295 349 296 
<< m2 >>
rect 349 295 350 296 
<< m1 >>
rect 350 295 351 296 
<< m2 >>
rect 350 295 351 296 
<< m2c >>
rect 350 295 351 296 
<< m1 >>
rect 350 295 351 296 
<< m2 >>
rect 350 295 351 296 
<< m2 >>
rect 351 295 352 296 
<< m1 >>
rect 352 295 353 296 
<< m2 >>
rect 352 295 353 296 
<< m2 >>
rect 353 295 354 296 
<< m1 >>
rect 354 295 355 296 
<< m2 >>
rect 354 295 355 296 
<< m2c >>
rect 354 295 355 296 
<< m1 >>
rect 354 295 355 296 
<< m2 >>
rect 354 295 355 296 
<< m1 >>
rect 355 295 356 296 
<< m1 >>
rect 366 295 367 296 
<< m1 >>
rect 367 295 368 296 
<< m1 >>
rect 368 295 369 296 
<< m2 >>
rect 368 295 369 296 
<< m2c >>
rect 368 295 369 296 
<< m1 >>
rect 368 295 369 296 
<< m2 >>
rect 368 295 369 296 
<< m2 >>
rect 369 295 370 296 
<< m1 >>
rect 370 295 371 296 
<< m2 >>
rect 370 295 371 296 
<< m2 >>
rect 371 295 372 296 
<< m1 >>
rect 372 295 373 296 
<< m2 >>
rect 372 295 373 296 
<< m2c >>
rect 372 295 373 296 
<< m1 >>
rect 372 295 373 296 
<< m2 >>
rect 372 295 373 296 
<< m1 >>
rect 373 295 374 296 
<< m1 >>
rect 374 295 375 296 
<< m1 >>
rect 375 295 376 296 
<< m1 >>
rect 376 295 377 296 
<< m1 >>
rect 379 295 380 296 
<< m2 >>
rect 380 295 381 296 
<< m1 >>
rect 381 295 382 296 
<< m1 >>
rect 382 295 383 296 
<< m1 >>
rect 383 295 384 296 
<< m1 >>
rect 384 295 385 296 
<< m1 >>
rect 385 295 386 296 
<< m1 >>
rect 386 295 387 296 
<< m1 >>
rect 387 295 388 296 
<< m1 >>
rect 388 295 389 296 
<< m1 >>
rect 389 295 390 296 
<< m1 >>
rect 390 295 391 296 
<< m1 >>
rect 391 295 392 296 
<< m1 >>
rect 392 295 393 296 
<< m2 >>
rect 392 295 393 296 
<< m2c >>
rect 392 295 393 296 
<< m1 >>
rect 392 295 393 296 
<< m2 >>
rect 392 295 393 296 
<< m2 >>
rect 393 295 394 296 
<< m1 >>
rect 394 295 395 296 
<< m2 >>
rect 394 295 395 296 
<< m2 >>
rect 395 295 396 296 
<< m1 >>
rect 396 295 397 296 
<< m2 >>
rect 396 295 397 296 
<< m2c >>
rect 396 295 397 296 
<< m1 >>
rect 396 295 397 296 
<< m2 >>
rect 396 295 397 296 
<< m1 >>
rect 397 295 398 296 
<< m1 >>
rect 398 295 399 296 
<< m1 >>
rect 399 295 400 296 
<< m1 >>
rect 400 295 401 296 
<< m1 >>
rect 401 295 402 296 
<< m1 >>
rect 402 295 403 296 
<< m1 >>
rect 403 295 404 296 
<< m1 >>
rect 404 295 405 296 
<< m1 >>
rect 405 295 406 296 
<< m1 >>
rect 406 295 407 296 
<< m1 >>
rect 407 295 408 296 
<< m1 >>
rect 408 295 409 296 
<< m1 >>
rect 409 295 410 296 
<< m2 >>
rect 415 295 416 296 
<< m1 >>
rect 416 295 417 296 
<< m2 >>
rect 416 295 417 296 
<< m2 >>
rect 417 295 418 296 
<< m1 >>
rect 418 295 419 296 
<< m2 >>
rect 418 295 419 296 
<< m2c >>
rect 418 295 419 296 
<< m1 >>
rect 418 295 419 296 
<< m2 >>
rect 418 295 419 296 
<< m2 >>
rect 419 295 420 296 
<< m1 >>
rect 420 295 421 296 
<< m1 >>
rect 421 295 422 296 
<< m1 >>
rect 422 295 423 296 
<< m1 >>
rect 423 295 424 296 
<< m1 >>
rect 424 295 425 296 
<< m1 >>
rect 425 295 426 296 
<< m1 >>
rect 426 295 427 296 
<< m1 >>
rect 427 295 428 296 
<< m1 >>
rect 428 295 429 296 
<< m1 >>
rect 429 295 430 296 
<< m1 >>
rect 430 295 431 296 
<< m1 >>
rect 433 295 434 296 
<< m1 >>
rect 437 295 438 296 
<< m2 >>
rect 437 295 438 296 
<< m2c >>
rect 437 295 438 296 
<< m1 >>
rect 437 295 438 296 
<< m2 >>
rect 437 295 438 296 
<< m1 >>
rect 487 295 488 296 
<< m1 >>
rect 523 295 524 296 
<< m1 >>
rect 19 296 20 297 
<< m1 >>
rect 22 296 23 297 
<< m1 >>
rect 44 296 45 297 
<< m1 >>
rect 46 296 47 297 
<< m1 >>
rect 55 296 56 297 
<< m1 >>
rect 73 296 74 297 
<< m2 >>
rect 74 296 75 297 
<< m2 >>
rect 91 296 92 297 
<< m2 >>
rect 93 296 94 297 
<< m1 >>
rect 106 296 107 297 
<< m2 >>
rect 107 296 108 297 
<< m1 >>
rect 146 296 147 297 
<< m2 >>
rect 146 296 147 297 
<< m2c >>
rect 146 296 147 297 
<< m1 >>
rect 146 296 147 297 
<< m2 >>
rect 146 296 147 297 
<< m1 >>
rect 148 296 149 297 
<< m2 >>
rect 148 296 149 297 
<< m2c >>
rect 148 296 149 297 
<< m1 >>
rect 148 296 149 297 
<< m2 >>
rect 148 296 149 297 
<< m2 >>
rect 149 296 150 297 
<< m1 >>
rect 150 296 151 297 
<< m2 >>
rect 150 296 151 297 
<< m2 >>
rect 151 296 152 297 
<< m1 >>
rect 181 296 182 297 
<< m1 >>
rect 186 296 187 297 
<< m1 >>
rect 208 296 209 297 
<< m1 >>
rect 217 296 218 297 
<< m2 >>
rect 217 296 218 297 
<< m1 >>
rect 226 296 227 297 
<< m1 >>
rect 232 296 233 297 
<< m1 >>
rect 244 296 245 297 
<< m1 >>
rect 246 296 247 297 
<< m1 >>
rect 255 296 256 297 
<< m1 >>
rect 271 296 272 297 
<< m1 >>
rect 278 296 279 297 
<< m1 >>
rect 280 296 281 297 
<< m1 >>
rect 282 296 283 297 
<< m2 >>
rect 284 296 285 297 
<< m1 >>
rect 307 296 308 297 
<< m1 >>
rect 309 296 310 297 
<< m2 >>
rect 310 296 311 297 
<< m2 >>
rect 333 296 334 297 
<< m1 >>
rect 334 296 335 297 
<< m1 >>
rect 344 296 345 297 
<< m1 >>
rect 348 296 349 297 
<< m1 >>
rect 352 296 353 297 
<< m1 >>
rect 355 296 356 297 
<< m1 >>
rect 366 296 367 297 
<< m1 >>
rect 370 296 371 297 
<< m1 >>
rect 376 296 377 297 
<< m1 >>
rect 379 296 380 297 
<< m2 >>
rect 380 296 381 297 
<< m1 >>
rect 381 296 382 297 
<< m1 >>
rect 394 296 395 297 
<< m1 >>
rect 416 296 417 297 
<< m1 >>
rect 418 296 419 297 
<< m2 >>
rect 419 296 420 297 
<< m1 >>
rect 420 296 421 297 
<< m1 >>
rect 433 296 434 297 
<< m2 >>
rect 437 296 438 297 
<< m1 >>
rect 487 296 488 297 
<< m1 >>
rect 523 296 524 297 
<< m1 >>
rect 19 297 20 298 
<< m1 >>
rect 22 297 23 298 
<< m1 >>
rect 44 297 45 298 
<< m1 >>
rect 46 297 47 298 
<< m1 >>
rect 55 297 56 298 
<< m1 >>
rect 73 297 74 298 
<< m2 >>
rect 74 297 75 298 
<< m1 >>
rect 91 297 92 298 
<< m2 >>
rect 91 297 92 298 
<< m2c >>
rect 91 297 92 298 
<< m1 >>
rect 91 297 92 298 
<< m2 >>
rect 91 297 92 298 
<< m1 >>
rect 93 297 94 298 
<< m2 >>
rect 93 297 94 298 
<< m2c >>
rect 93 297 94 298 
<< m1 >>
rect 93 297 94 298 
<< m2 >>
rect 93 297 94 298 
<< m1 >>
rect 103 297 104 298 
<< m1 >>
rect 104 297 105 298 
<< m2 >>
rect 104 297 105 298 
<< m2c >>
rect 104 297 105 298 
<< m1 >>
rect 104 297 105 298 
<< m2 >>
rect 104 297 105 298 
<< m2 >>
rect 105 297 106 298 
<< m1 >>
rect 106 297 107 298 
<< m2 >>
rect 106 297 107 298 
<< m2 >>
rect 107 297 108 298 
<< m1 >>
rect 146 297 147 298 
<< m1 >>
rect 148 297 149 298 
<< m1 >>
rect 150 297 151 298 
<< m1 >>
rect 181 297 182 298 
<< m1 >>
rect 186 297 187 298 
<< m1 >>
rect 208 297 209 298 
<< m1 >>
rect 211 297 212 298 
<< m1 >>
rect 212 297 213 298 
<< m1 >>
rect 213 297 214 298 
<< m1 >>
rect 214 297 215 298 
<< m1 >>
rect 215 297 216 298 
<< m1 >>
rect 216 297 217 298 
<< m1 >>
rect 217 297 218 298 
<< m2 >>
rect 217 297 218 298 
<< m1 >>
rect 226 297 227 298 
<< m1 >>
rect 232 297 233 298 
<< m1 >>
rect 233 297 234 298 
<< m1 >>
rect 234 297 235 298 
<< m1 >>
rect 235 297 236 298 
<< m1 >>
rect 236 297 237 298 
<< m1 >>
rect 237 297 238 298 
<< m1 >>
rect 244 297 245 298 
<< m1 >>
rect 246 297 247 298 
<< m1 >>
rect 255 297 256 298 
<< m1 >>
rect 271 297 272 298 
<< m1 >>
rect 278 297 279 298 
<< m1 >>
rect 280 297 281 298 
<< m1 >>
rect 282 297 283 298 
<< m1 >>
rect 284 297 285 298 
<< m2 >>
rect 284 297 285 298 
<< m2c >>
rect 284 297 285 298 
<< m1 >>
rect 284 297 285 298 
<< m2 >>
rect 284 297 285 298 
<< m1 >>
rect 285 297 286 298 
<< m1 >>
rect 286 297 287 298 
<< m1 >>
rect 307 297 308 298 
<< m1 >>
rect 309 297 310 298 
<< m2 >>
rect 310 297 311 298 
<< m2 >>
rect 333 297 334 298 
<< m1 >>
rect 334 297 335 298 
<< m1 >>
rect 344 297 345 298 
<< m1 >>
rect 348 297 349 298 
<< m1 >>
rect 352 297 353 298 
<< m1 >>
rect 355 297 356 298 
<< m1 >>
rect 366 297 367 298 
<< m1 >>
rect 370 297 371 298 
<< m1 >>
rect 376 297 377 298 
<< m1 >>
rect 379 297 380 298 
<< m2 >>
rect 380 297 381 298 
<< m1 >>
rect 381 297 382 298 
<< m1 >>
rect 391 297 392 298 
<< m1 >>
rect 392 297 393 298 
<< m2 >>
rect 392 297 393 298 
<< m2c >>
rect 392 297 393 298 
<< m1 >>
rect 392 297 393 298 
<< m2 >>
rect 392 297 393 298 
<< m2 >>
rect 393 297 394 298 
<< m1 >>
rect 394 297 395 298 
<< m2 >>
rect 394 297 395 298 
<< m2 >>
rect 395 297 396 298 
<< m1 >>
rect 416 297 417 298 
<< m1 >>
rect 418 297 419 298 
<< m2 >>
rect 419 297 420 298 
<< m1 >>
rect 420 297 421 298 
<< m2 >>
rect 420 297 421 298 
<< m2 >>
rect 421 297 422 298 
<< m1 >>
rect 422 297 423 298 
<< m2 >>
rect 422 297 423 298 
<< m2c >>
rect 422 297 423 298 
<< m1 >>
rect 422 297 423 298 
<< m2 >>
rect 422 297 423 298 
<< m1 >>
rect 427 297 428 298 
<< m1 >>
rect 428 297 429 298 
<< m1 >>
rect 429 297 430 298 
<< m1 >>
rect 430 297 431 298 
<< m1 >>
rect 431 297 432 298 
<< m2 >>
rect 431 297 432 298 
<< m2c >>
rect 431 297 432 298 
<< m1 >>
rect 431 297 432 298 
<< m2 >>
rect 431 297 432 298 
<< m2 >>
rect 432 297 433 298 
<< m1 >>
rect 433 297 434 298 
<< m2 >>
rect 433 297 434 298 
<< m2 >>
rect 434 297 435 298 
<< m1 >>
rect 435 297 436 298 
<< m2 >>
rect 435 297 436 298 
<< m2c >>
rect 435 297 436 298 
<< m1 >>
rect 435 297 436 298 
<< m2 >>
rect 435 297 436 298 
<< m1 >>
rect 436 297 437 298 
<< m1 >>
rect 437 297 438 298 
<< m2 >>
rect 437 297 438 298 
<< m1 >>
rect 487 297 488 298 
<< m1 >>
rect 523 297 524 298 
<< m1 >>
rect 19 298 20 299 
<< m1 >>
rect 22 298 23 299 
<< m1 >>
rect 44 298 45 299 
<< m1 >>
rect 46 298 47 299 
<< m2 >>
rect 46 298 47 299 
<< m2 >>
rect 47 298 48 299 
<< m1 >>
rect 48 298 49 299 
<< m2 >>
rect 48 298 49 299 
<< m2c >>
rect 48 298 49 299 
<< m1 >>
rect 48 298 49 299 
<< m2 >>
rect 48 298 49 299 
<< m1 >>
rect 49 298 50 299 
<< m1 >>
rect 55 298 56 299 
<< m1 >>
rect 73 298 74 299 
<< m2 >>
rect 74 298 75 299 
<< m1 >>
rect 91 298 92 299 
<< m1 >>
rect 93 298 94 299 
<< m1 >>
rect 103 298 104 299 
<< m1 >>
rect 106 298 107 299 
<< m1 >>
rect 146 298 147 299 
<< m1 >>
rect 148 298 149 299 
<< m1 >>
rect 150 298 151 299 
<< m1 >>
rect 181 298 182 299 
<< m1 >>
rect 186 298 187 299 
<< m1 >>
rect 208 298 209 299 
<< m1 >>
rect 211 298 212 299 
<< m2 >>
rect 217 298 218 299 
<< m1 >>
rect 226 298 227 299 
<< m1 >>
rect 237 298 238 299 
<< m2 >>
rect 243 298 244 299 
<< m1 >>
rect 244 298 245 299 
<< m2 >>
rect 244 298 245 299 
<< m2 >>
rect 245 298 246 299 
<< m1 >>
rect 246 298 247 299 
<< m2 >>
rect 246 298 247 299 
<< m2c >>
rect 246 298 247 299 
<< m1 >>
rect 246 298 247 299 
<< m2 >>
rect 246 298 247 299 
<< m1 >>
rect 255 298 256 299 
<< m1 >>
rect 271 298 272 299 
<< m2 >>
rect 277 298 278 299 
<< m1 >>
rect 278 298 279 299 
<< m2 >>
rect 278 298 279 299 
<< m2 >>
rect 279 298 280 299 
<< m1 >>
rect 280 298 281 299 
<< m2 >>
rect 280 298 281 299 
<< m2 >>
rect 281 298 282 299 
<< m1 >>
rect 282 298 283 299 
<< m2 >>
rect 282 298 283 299 
<< m2c >>
rect 282 298 283 299 
<< m1 >>
rect 282 298 283 299 
<< m2 >>
rect 282 298 283 299 
<< m1 >>
rect 286 298 287 299 
<< m1 >>
rect 307 298 308 299 
<< m1 >>
rect 309 298 310 299 
<< m2 >>
rect 310 298 311 299 
<< m2 >>
rect 333 298 334 299 
<< m1 >>
rect 334 298 335 299 
<< m1 >>
rect 340 298 341 299 
<< m1 >>
rect 341 298 342 299 
<< m1 >>
rect 342 298 343 299 
<< m2 >>
rect 342 298 343 299 
<< m2c >>
rect 342 298 343 299 
<< m1 >>
rect 342 298 343 299 
<< m2 >>
rect 342 298 343 299 
<< m2 >>
rect 343 298 344 299 
<< m1 >>
rect 344 298 345 299 
<< m2 >>
rect 344 298 345 299 
<< m2 >>
rect 345 298 346 299 
<< m1 >>
rect 348 298 349 299 
<< m1 >>
rect 352 298 353 299 
<< m1 >>
rect 355 298 356 299 
<< m1 >>
rect 366 298 367 299 
<< m1 >>
rect 370 298 371 299 
<< m1 >>
rect 376 298 377 299 
<< m1 >>
rect 379 298 380 299 
<< m2 >>
rect 380 298 381 299 
<< m1 >>
rect 381 298 382 299 
<< m1 >>
rect 391 298 392 299 
<< m1 >>
rect 394 298 395 299 
<< m2 >>
rect 395 298 396 299 
<< m1 >>
rect 396 298 397 299 
<< m2 >>
rect 396 298 397 299 
<< m2c >>
rect 396 298 397 299 
<< m1 >>
rect 396 298 397 299 
<< m2 >>
rect 396 298 397 299 
<< m1 >>
rect 397 298 398 299 
<< m1 >>
rect 398 298 399 299 
<< m1 >>
rect 399 298 400 299 
<< m1 >>
rect 400 298 401 299 
<< m1 >>
rect 401 298 402 299 
<< m1 >>
rect 402 298 403 299 
<< m1 >>
rect 403 298 404 299 
<< m1 >>
rect 404 298 405 299 
<< m1 >>
rect 405 298 406 299 
<< m1 >>
rect 406 298 407 299 
<< m1 >>
rect 416 298 417 299 
<< m1 >>
rect 418 298 419 299 
<< m1 >>
rect 420 298 421 299 
<< m1 >>
rect 422 298 423 299 
<< m1 >>
rect 427 298 428 299 
<< m1 >>
rect 433 298 434 299 
<< m1 >>
rect 437 298 438 299 
<< m2 >>
rect 437 298 438 299 
<< m1 >>
rect 487 298 488 299 
<< m1 >>
rect 523 298 524 299 
<< m1 >>
rect 19 299 20 300 
<< m1 >>
rect 22 299 23 300 
<< m1 >>
rect 44 299 45 300 
<< m1 >>
rect 46 299 47 300 
<< m2 >>
rect 46 299 47 300 
<< m1 >>
rect 49 299 50 300 
<< m1 >>
rect 55 299 56 300 
<< m1 >>
rect 73 299 74 300 
<< m2 >>
rect 74 299 75 300 
<< m1 >>
rect 91 299 92 300 
<< m1 >>
rect 93 299 94 300 
<< m1 >>
rect 103 299 104 300 
<< m1 >>
rect 106 299 107 300 
<< m1 >>
rect 146 299 147 300 
<< m1 >>
rect 148 299 149 300 
<< m1 >>
rect 150 299 151 300 
<< m1 >>
rect 181 299 182 300 
<< m1 >>
rect 186 299 187 300 
<< m1 >>
rect 208 299 209 300 
<< m1 >>
rect 211 299 212 300 
<< m1 >>
rect 217 299 218 300 
<< m2 >>
rect 217 299 218 300 
<< m2c >>
rect 217 299 218 300 
<< m1 >>
rect 217 299 218 300 
<< m2 >>
rect 217 299 218 300 
<< m1 >>
rect 226 299 227 300 
<< m1 >>
rect 237 299 238 300 
<< m2 >>
rect 243 299 244 300 
<< m1 >>
rect 244 299 245 300 
<< m1 >>
rect 255 299 256 300 
<< m1 >>
rect 271 299 272 300 
<< m2 >>
rect 277 299 278 300 
<< m1 >>
rect 278 299 279 300 
<< m1 >>
rect 280 299 281 300 
<< m1 >>
rect 286 299 287 300 
<< m1 >>
rect 307 299 308 300 
<< m1 >>
rect 309 299 310 300 
<< m2 >>
rect 310 299 311 300 
<< m2 >>
rect 333 299 334 300 
<< m1 >>
rect 334 299 335 300 
<< m1 >>
rect 340 299 341 300 
<< m1 >>
rect 344 299 345 300 
<< m2 >>
rect 345 299 346 300 
<< m1 >>
rect 348 299 349 300 
<< m1 >>
rect 352 299 353 300 
<< m1 >>
rect 355 299 356 300 
<< m1 >>
rect 366 299 367 300 
<< m1 >>
rect 370 299 371 300 
<< m1 >>
rect 376 299 377 300 
<< m1 >>
rect 379 299 380 300 
<< m2 >>
rect 380 299 381 300 
<< m1 >>
rect 381 299 382 300 
<< m1 >>
rect 391 299 392 300 
<< m1 >>
rect 394 299 395 300 
<< m1 >>
rect 406 299 407 300 
<< m1 >>
rect 416 299 417 300 
<< m1 >>
rect 418 299 419 300 
<< m2 >>
rect 418 299 419 300 
<< m2c >>
rect 418 299 419 300 
<< m1 >>
rect 418 299 419 300 
<< m2 >>
rect 418 299 419 300 
<< m2 >>
rect 419 299 420 300 
<< m1 >>
rect 420 299 421 300 
<< m1 >>
rect 422 299 423 300 
<< m1 >>
rect 427 299 428 300 
<< m1 >>
rect 433 299 434 300 
<< m2 >>
rect 434 299 435 300 
<< m1 >>
rect 435 299 436 300 
<< m2 >>
rect 435 299 436 300 
<< m2c >>
rect 435 299 436 300 
<< m1 >>
rect 435 299 436 300 
<< m2 >>
rect 435 299 436 300 
<< m2 >>
rect 436 299 437 300 
<< m1 >>
rect 437 299 438 300 
<< m2 >>
rect 437 299 438 300 
<< m1 >>
rect 487 299 488 300 
<< m1 >>
rect 523 299 524 300 
<< pdiffusion >>
rect 12 300 13 301 
<< pdiffusion >>
rect 13 300 14 301 
<< pdiffusion >>
rect 14 300 15 301 
<< pdiffusion >>
rect 15 300 16 301 
<< pdiffusion >>
rect 16 300 17 301 
<< pdiffusion >>
rect 17 300 18 301 
<< m1 >>
rect 19 300 20 301 
<< m1 >>
rect 22 300 23 301 
<< pdiffusion >>
rect 30 300 31 301 
<< pdiffusion >>
rect 31 300 32 301 
<< pdiffusion >>
rect 32 300 33 301 
<< pdiffusion >>
rect 33 300 34 301 
<< pdiffusion >>
rect 34 300 35 301 
<< pdiffusion >>
rect 35 300 36 301 
<< m1 >>
rect 44 300 45 301 
<< m1 >>
rect 46 300 47 301 
<< m2 >>
rect 46 300 47 301 
<< pdiffusion >>
rect 48 300 49 301 
<< m1 >>
rect 49 300 50 301 
<< pdiffusion >>
rect 49 300 50 301 
<< pdiffusion >>
rect 50 300 51 301 
<< pdiffusion >>
rect 51 300 52 301 
<< pdiffusion >>
rect 52 300 53 301 
<< pdiffusion >>
rect 53 300 54 301 
<< m1 >>
rect 55 300 56 301 
<< pdiffusion >>
rect 66 300 67 301 
<< pdiffusion >>
rect 67 300 68 301 
<< pdiffusion >>
rect 68 300 69 301 
<< pdiffusion >>
rect 69 300 70 301 
<< pdiffusion >>
rect 70 300 71 301 
<< pdiffusion >>
rect 71 300 72 301 
<< m1 >>
rect 73 300 74 301 
<< m2 >>
rect 74 300 75 301 
<< pdiffusion >>
rect 84 300 85 301 
<< pdiffusion >>
rect 85 300 86 301 
<< pdiffusion >>
rect 86 300 87 301 
<< pdiffusion >>
rect 87 300 88 301 
<< pdiffusion >>
rect 88 300 89 301 
<< pdiffusion >>
rect 89 300 90 301 
<< m1 >>
rect 91 300 92 301 
<< m1 >>
rect 93 300 94 301 
<< pdiffusion >>
rect 102 300 103 301 
<< m1 >>
rect 103 300 104 301 
<< pdiffusion >>
rect 103 300 104 301 
<< pdiffusion >>
rect 104 300 105 301 
<< pdiffusion >>
rect 105 300 106 301 
<< m1 >>
rect 106 300 107 301 
<< pdiffusion >>
rect 106 300 107 301 
<< pdiffusion >>
rect 107 300 108 301 
<< pdiffusion >>
rect 120 300 121 301 
<< pdiffusion >>
rect 121 300 122 301 
<< pdiffusion >>
rect 122 300 123 301 
<< pdiffusion >>
rect 123 300 124 301 
<< pdiffusion >>
rect 124 300 125 301 
<< pdiffusion >>
rect 125 300 126 301 
<< pdiffusion >>
rect 138 300 139 301 
<< pdiffusion >>
rect 139 300 140 301 
<< pdiffusion >>
rect 140 300 141 301 
<< pdiffusion >>
rect 141 300 142 301 
<< pdiffusion >>
rect 142 300 143 301 
<< pdiffusion >>
rect 143 300 144 301 
<< m1 >>
rect 146 300 147 301 
<< m1 >>
rect 148 300 149 301 
<< m1 >>
rect 150 300 151 301 
<< pdiffusion >>
rect 156 300 157 301 
<< pdiffusion >>
rect 157 300 158 301 
<< pdiffusion >>
rect 158 300 159 301 
<< pdiffusion >>
rect 159 300 160 301 
<< pdiffusion >>
rect 160 300 161 301 
<< pdiffusion >>
rect 161 300 162 301 
<< pdiffusion >>
rect 174 300 175 301 
<< pdiffusion >>
rect 175 300 176 301 
<< pdiffusion >>
rect 176 300 177 301 
<< pdiffusion >>
rect 177 300 178 301 
<< pdiffusion >>
rect 178 300 179 301 
<< pdiffusion >>
rect 179 300 180 301 
<< m1 >>
rect 181 300 182 301 
<< m1 >>
rect 186 300 187 301 
<< pdiffusion >>
rect 192 300 193 301 
<< pdiffusion >>
rect 193 300 194 301 
<< pdiffusion >>
rect 194 300 195 301 
<< pdiffusion >>
rect 195 300 196 301 
<< pdiffusion >>
rect 196 300 197 301 
<< pdiffusion >>
rect 197 300 198 301 
<< m1 >>
rect 208 300 209 301 
<< pdiffusion >>
rect 210 300 211 301 
<< m1 >>
rect 211 300 212 301 
<< pdiffusion >>
rect 211 300 212 301 
<< pdiffusion >>
rect 212 300 213 301 
<< pdiffusion >>
rect 213 300 214 301 
<< pdiffusion >>
rect 214 300 215 301 
<< pdiffusion >>
rect 215 300 216 301 
<< m1 >>
rect 217 300 218 301 
<< m1 >>
rect 226 300 227 301 
<< pdiffusion >>
rect 228 300 229 301 
<< pdiffusion >>
rect 229 300 230 301 
<< pdiffusion >>
rect 230 300 231 301 
<< pdiffusion >>
rect 231 300 232 301 
<< pdiffusion >>
rect 232 300 233 301 
<< pdiffusion >>
rect 233 300 234 301 
<< m1 >>
rect 237 300 238 301 
<< m2 >>
rect 243 300 244 301 
<< m1 >>
rect 244 300 245 301 
<< pdiffusion >>
rect 246 300 247 301 
<< pdiffusion >>
rect 247 300 248 301 
<< pdiffusion >>
rect 248 300 249 301 
<< pdiffusion >>
rect 249 300 250 301 
<< pdiffusion >>
rect 250 300 251 301 
<< pdiffusion >>
rect 251 300 252 301 
<< m1 >>
rect 255 300 256 301 
<< pdiffusion >>
rect 264 300 265 301 
<< pdiffusion >>
rect 265 300 266 301 
<< pdiffusion >>
rect 266 300 267 301 
<< pdiffusion >>
rect 267 300 268 301 
<< pdiffusion >>
rect 268 300 269 301 
<< pdiffusion >>
rect 269 300 270 301 
<< m1 >>
rect 271 300 272 301 
<< m2 >>
rect 277 300 278 301 
<< m1 >>
rect 278 300 279 301 
<< m1 >>
rect 280 300 281 301 
<< pdiffusion >>
rect 282 300 283 301 
<< pdiffusion >>
rect 283 300 284 301 
<< pdiffusion >>
rect 284 300 285 301 
<< pdiffusion >>
rect 285 300 286 301 
<< m1 >>
rect 286 300 287 301 
<< pdiffusion >>
rect 286 300 287 301 
<< pdiffusion >>
rect 287 300 288 301 
<< pdiffusion >>
rect 300 300 301 301 
<< pdiffusion >>
rect 301 300 302 301 
<< pdiffusion >>
rect 302 300 303 301 
<< pdiffusion >>
rect 303 300 304 301 
<< pdiffusion >>
rect 304 300 305 301 
<< pdiffusion >>
rect 305 300 306 301 
<< m1 >>
rect 307 300 308 301 
<< m1 >>
rect 309 300 310 301 
<< m2 >>
rect 310 300 311 301 
<< pdiffusion >>
rect 318 300 319 301 
<< pdiffusion >>
rect 319 300 320 301 
<< pdiffusion >>
rect 320 300 321 301 
<< pdiffusion >>
rect 321 300 322 301 
<< pdiffusion >>
rect 322 300 323 301 
<< pdiffusion >>
rect 323 300 324 301 
<< m2 >>
rect 333 300 334 301 
<< m1 >>
rect 334 300 335 301 
<< pdiffusion >>
rect 336 300 337 301 
<< pdiffusion >>
rect 337 300 338 301 
<< pdiffusion >>
rect 338 300 339 301 
<< pdiffusion >>
rect 339 300 340 301 
<< m1 >>
rect 340 300 341 301 
<< pdiffusion >>
rect 340 300 341 301 
<< pdiffusion >>
rect 341 300 342 301 
<< m1 >>
rect 344 300 345 301 
<< m2 >>
rect 345 300 346 301 
<< m1 >>
rect 348 300 349 301 
<< m1 >>
rect 352 300 353 301 
<< pdiffusion >>
rect 354 300 355 301 
<< m1 >>
rect 355 300 356 301 
<< pdiffusion >>
rect 355 300 356 301 
<< pdiffusion >>
rect 356 300 357 301 
<< pdiffusion >>
rect 357 300 358 301 
<< pdiffusion >>
rect 358 300 359 301 
<< pdiffusion >>
rect 359 300 360 301 
<< m1 >>
rect 366 300 367 301 
<< m1 >>
rect 370 300 371 301 
<< pdiffusion >>
rect 372 300 373 301 
<< pdiffusion >>
rect 373 300 374 301 
<< pdiffusion >>
rect 374 300 375 301 
<< pdiffusion >>
rect 375 300 376 301 
<< m1 >>
rect 376 300 377 301 
<< pdiffusion >>
rect 376 300 377 301 
<< pdiffusion >>
rect 377 300 378 301 
<< m1 >>
rect 379 300 380 301 
<< m2 >>
rect 380 300 381 301 
<< m1 >>
rect 381 300 382 301 
<< pdiffusion >>
rect 390 300 391 301 
<< m1 >>
rect 391 300 392 301 
<< pdiffusion >>
rect 391 300 392 301 
<< pdiffusion >>
rect 392 300 393 301 
<< pdiffusion >>
rect 393 300 394 301 
<< m1 >>
rect 394 300 395 301 
<< pdiffusion >>
rect 394 300 395 301 
<< pdiffusion >>
rect 395 300 396 301 
<< m1 >>
rect 406 300 407 301 
<< pdiffusion >>
rect 408 300 409 301 
<< pdiffusion >>
rect 409 300 410 301 
<< pdiffusion >>
rect 410 300 411 301 
<< pdiffusion >>
rect 411 300 412 301 
<< pdiffusion >>
rect 412 300 413 301 
<< pdiffusion >>
rect 413 300 414 301 
<< m1 >>
rect 416 300 417 301 
<< m2 >>
rect 419 300 420 301 
<< m1 >>
rect 420 300 421 301 
<< m1 >>
rect 422 300 423 301 
<< pdiffusion >>
rect 426 300 427 301 
<< m1 >>
rect 427 300 428 301 
<< pdiffusion >>
rect 427 300 428 301 
<< pdiffusion >>
rect 428 300 429 301 
<< pdiffusion >>
rect 429 300 430 301 
<< pdiffusion >>
rect 430 300 431 301 
<< pdiffusion >>
rect 431 300 432 301 
<< m1 >>
rect 433 300 434 301 
<< m2 >>
rect 434 300 435 301 
<< m1 >>
rect 437 300 438 301 
<< pdiffusion >>
rect 444 300 445 301 
<< pdiffusion >>
rect 445 300 446 301 
<< pdiffusion >>
rect 446 300 447 301 
<< pdiffusion >>
rect 447 300 448 301 
<< pdiffusion >>
rect 448 300 449 301 
<< pdiffusion >>
rect 449 300 450 301 
<< pdiffusion >>
rect 462 300 463 301 
<< pdiffusion >>
rect 463 300 464 301 
<< pdiffusion >>
rect 464 300 465 301 
<< pdiffusion >>
rect 465 300 466 301 
<< pdiffusion >>
rect 466 300 467 301 
<< pdiffusion >>
rect 467 300 468 301 
<< pdiffusion >>
rect 480 300 481 301 
<< pdiffusion >>
rect 481 300 482 301 
<< pdiffusion >>
rect 482 300 483 301 
<< pdiffusion >>
rect 483 300 484 301 
<< pdiffusion >>
rect 484 300 485 301 
<< pdiffusion >>
rect 485 300 486 301 
<< m1 >>
rect 487 300 488 301 
<< pdiffusion >>
rect 498 300 499 301 
<< pdiffusion >>
rect 499 300 500 301 
<< pdiffusion >>
rect 500 300 501 301 
<< pdiffusion >>
rect 501 300 502 301 
<< pdiffusion >>
rect 502 300 503 301 
<< pdiffusion >>
rect 503 300 504 301 
<< m1 >>
rect 523 300 524 301 
<< pdiffusion >>
rect 12 301 13 302 
<< pdiffusion >>
rect 13 301 14 302 
<< pdiffusion >>
rect 14 301 15 302 
<< pdiffusion >>
rect 15 301 16 302 
<< pdiffusion >>
rect 16 301 17 302 
<< pdiffusion >>
rect 17 301 18 302 
<< m1 >>
rect 19 301 20 302 
<< m1 >>
rect 22 301 23 302 
<< pdiffusion >>
rect 30 301 31 302 
<< pdiffusion >>
rect 31 301 32 302 
<< pdiffusion >>
rect 32 301 33 302 
<< pdiffusion >>
rect 33 301 34 302 
<< pdiffusion >>
rect 34 301 35 302 
<< pdiffusion >>
rect 35 301 36 302 
<< m1 >>
rect 44 301 45 302 
<< m1 >>
rect 46 301 47 302 
<< m2 >>
rect 46 301 47 302 
<< pdiffusion >>
rect 48 301 49 302 
<< pdiffusion >>
rect 49 301 50 302 
<< pdiffusion >>
rect 50 301 51 302 
<< pdiffusion >>
rect 51 301 52 302 
<< pdiffusion >>
rect 52 301 53 302 
<< pdiffusion >>
rect 53 301 54 302 
<< m1 >>
rect 55 301 56 302 
<< pdiffusion >>
rect 66 301 67 302 
<< pdiffusion >>
rect 67 301 68 302 
<< pdiffusion >>
rect 68 301 69 302 
<< pdiffusion >>
rect 69 301 70 302 
<< pdiffusion >>
rect 70 301 71 302 
<< pdiffusion >>
rect 71 301 72 302 
<< m1 >>
rect 73 301 74 302 
<< m2 >>
rect 74 301 75 302 
<< pdiffusion >>
rect 84 301 85 302 
<< pdiffusion >>
rect 85 301 86 302 
<< pdiffusion >>
rect 86 301 87 302 
<< pdiffusion >>
rect 87 301 88 302 
<< pdiffusion >>
rect 88 301 89 302 
<< pdiffusion >>
rect 89 301 90 302 
<< m1 >>
rect 91 301 92 302 
<< m1 >>
rect 93 301 94 302 
<< pdiffusion >>
rect 102 301 103 302 
<< pdiffusion >>
rect 103 301 104 302 
<< pdiffusion >>
rect 104 301 105 302 
<< pdiffusion >>
rect 105 301 106 302 
<< pdiffusion >>
rect 106 301 107 302 
<< pdiffusion >>
rect 107 301 108 302 
<< pdiffusion >>
rect 120 301 121 302 
<< pdiffusion >>
rect 121 301 122 302 
<< pdiffusion >>
rect 122 301 123 302 
<< pdiffusion >>
rect 123 301 124 302 
<< pdiffusion >>
rect 124 301 125 302 
<< pdiffusion >>
rect 125 301 126 302 
<< pdiffusion >>
rect 138 301 139 302 
<< pdiffusion >>
rect 139 301 140 302 
<< pdiffusion >>
rect 140 301 141 302 
<< pdiffusion >>
rect 141 301 142 302 
<< pdiffusion >>
rect 142 301 143 302 
<< pdiffusion >>
rect 143 301 144 302 
<< m1 >>
rect 146 301 147 302 
<< m1 >>
rect 148 301 149 302 
<< m1 >>
rect 150 301 151 302 
<< pdiffusion >>
rect 156 301 157 302 
<< pdiffusion >>
rect 157 301 158 302 
<< pdiffusion >>
rect 158 301 159 302 
<< pdiffusion >>
rect 159 301 160 302 
<< pdiffusion >>
rect 160 301 161 302 
<< pdiffusion >>
rect 161 301 162 302 
<< pdiffusion >>
rect 174 301 175 302 
<< pdiffusion >>
rect 175 301 176 302 
<< pdiffusion >>
rect 176 301 177 302 
<< pdiffusion >>
rect 177 301 178 302 
<< pdiffusion >>
rect 178 301 179 302 
<< pdiffusion >>
rect 179 301 180 302 
<< m1 >>
rect 181 301 182 302 
<< m1 >>
rect 186 301 187 302 
<< pdiffusion >>
rect 192 301 193 302 
<< pdiffusion >>
rect 193 301 194 302 
<< pdiffusion >>
rect 194 301 195 302 
<< pdiffusion >>
rect 195 301 196 302 
<< pdiffusion >>
rect 196 301 197 302 
<< pdiffusion >>
rect 197 301 198 302 
<< m1 >>
rect 208 301 209 302 
<< pdiffusion >>
rect 210 301 211 302 
<< pdiffusion >>
rect 211 301 212 302 
<< pdiffusion >>
rect 212 301 213 302 
<< pdiffusion >>
rect 213 301 214 302 
<< pdiffusion >>
rect 214 301 215 302 
<< pdiffusion >>
rect 215 301 216 302 
<< m1 >>
rect 217 301 218 302 
<< m2 >>
rect 218 301 219 302 
<< m1 >>
rect 219 301 220 302 
<< m2 >>
rect 219 301 220 302 
<< m2c >>
rect 219 301 220 302 
<< m1 >>
rect 219 301 220 302 
<< m2 >>
rect 219 301 220 302 
<< m1 >>
rect 220 301 221 302 
<< m1 >>
rect 221 301 222 302 
<< m1 >>
rect 222 301 223 302 
<< m1 >>
rect 223 301 224 302 
<< m1 >>
rect 224 301 225 302 
<< m1 >>
rect 225 301 226 302 
<< m1 >>
rect 226 301 227 302 
<< pdiffusion >>
rect 228 301 229 302 
<< pdiffusion >>
rect 229 301 230 302 
<< pdiffusion >>
rect 230 301 231 302 
<< pdiffusion >>
rect 231 301 232 302 
<< pdiffusion >>
rect 232 301 233 302 
<< pdiffusion >>
rect 233 301 234 302 
<< m1 >>
rect 237 301 238 302 
<< m2 >>
rect 243 301 244 302 
<< m1 >>
rect 244 301 245 302 
<< pdiffusion >>
rect 246 301 247 302 
<< pdiffusion >>
rect 247 301 248 302 
<< pdiffusion >>
rect 248 301 249 302 
<< pdiffusion >>
rect 249 301 250 302 
<< pdiffusion >>
rect 250 301 251 302 
<< pdiffusion >>
rect 251 301 252 302 
<< m1 >>
rect 255 301 256 302 
<< pdiffusion >>
rect 264 301 265 302 
<< pdiffusion >>
rect 265 301 266 302 
<< pdiffusion >>
rect 266 301 267 302 
<< pdiffusion >>
rect 267 301 268 302 
<< pdiffusion >>
rect 268 301 269 302 
<< pdiffusion >>
rect 269 301 270 302 
<< m1 >>
rect 271 301 272 302 
<< m2 >>
rect 277 301 278 302 
<< m1 >>
rect 278 301 279 302 
<< m1 >>
rect 280 301 281 302 
<< pdiffusion >>
rect 282 301 283 302 
<< pdiffusion >>
rect 283 301 284 302 
<< pdiffusion >>
rect 284 301 285 302 
<< pdiffusion >>
rect 285 301 286 302 
<< pdiffusion >>
rect 286 301 287 302 
<< pdiffusion >>
rect 287 301 288 302 
<< pdiffusion >>
rect 300 301 301 302 
<< pdiffusion >>
rect 301 301 302 302 
<< pdiffusion >>
rect 302 301 303 302 
<< pdiffusion >>
rect 303 301 304 302 
<< pdiffusion >>
rect 304 301 305 302 
<< pdiffusion >>
rect 305 301 306 302 
<< m1 >>
rect 307 301 308 302 
<< m1 >>
rect 309 301 310 302 
<< m2 >>
rect 310 301 311 302 
<< pdiffusion >>
rect 318 301 319 302 
<< pdiffusion >>
rect 319 301 320 302 
<< pdiffusion >>
rect 320 301 321 302 
<< pdiffusion >>
rect 321 301 322 302 
<< pdiffusion >>
rect 322 301 323 302 
<< pdiffusion >>
rect 323 301 324 302 
<< m2 >>
rect 333 301 334 302 
<< m1 >>
rect 334 301 335 302 
<< pdiffusion >>
rect 336 301 337 302 
<< pdiffusion >>
rect 337 301 338 302 
<< pdiffusion >>
rect 338 301 339 302 
<< pdiffusion >>
rect 339 301 340 302 
<< pdiffusion >>
rect 340 301 341 302 
<< pdiffusion >>
rect 341 301 342 302 
<< m1 >>
rect 344 301 345 302 
<< m2 >>
rect 345 301 346 302 
<< m1 >>
rect 348 301 349 302 
<< m1 >>
rect 352 301 353 302 
<< pdiffusion >>
rect 354 301 355 302 
<< pdiffusion >>
rect 355 301 356 302 
<< pdiffusion >>
rect 356 301 357 302 
<< pdiffusion >>
rect 357 301 358 302 
<< pdiffusion >>
rect 358 301 359 302 
<< pdiffusion >>
rect 359 301 360 302 
<< m1 >>
rect 366 301 367 302 
<< m1 >>
rect 370 301 371 302 
<< pdiffusion >>
rect 372 301 373 302 
<< pdiffusion >>
rect 373 301 374 302 
<< pdiffusion >>
rect 374 301 375 302 
<< pdiffusion >>
rect 375 301 376 302 
<< pdiffusion >>
rect 376 301 377 302 
<< pdiffusion >>
rect 377 301 378 302 
<< m1 >>
rect 379 301 380 302 
<< m2 >>
rect 380 301 381 302 
<< m1 >>
rect 381 301 382 302 
<< pdiffusion >>
rect 390 301 391 302 
<< pdiffusion >>
rect 391 301 392 302 
<< pdiffusion >>
rect 392 301 393 302 
<< pdiffusion >>
rect 393 301 394 302 
<< pdiffusion >>
rect 394 301 395 302 
<< pdiffusion >>
rect 395 301 396 302 
<< m1 >>
rect 406 301 407 302 
<< pdiffusion >>
rect 408 301 409 302 
<< pdiffusion >>
rect 409 301 410 302 
<< pdiffusion >>
rect 410 301 411 302 
<< pdiffusion >>
rect 411 301 412 302 
<< pdiffusion >>
rect 412 301 413 302 
<< pdiffusion >>
rect 413 301 414 302 
<< m1 >>
rect 416 301 417 302 
<< m2 >>
rect 419 301 420 302 
<< m1 >>
rect 420 301 421 302 
<< m1 >>
rect 422 301 423 302 
<< pdiffusion >>
rect 426 301 427 302 
<< pdiffusion >>
rect 427 301 428 302 
<< pdiffusion >>
rect 428 301 429 302 
<< pdiffusion >>
rect 429 301 430 302 
<< pdiffusion >>
rect 430 301 431 302 
<< pdiffusion >>
rect 431 301 432 302 
<< m1 >>
rect 433 301 434 302 
<< m2 >>
rect 434 301 435 302 
<< m1 >>
rect 437 301 438 302 
<< pdiffusion >>
rect 444 301 445 302 
<< pdiffusion >>
rect 445 301 446 302 
<< pdiffusion >>
rect 446 301 447 302 
<< pdiffusion >>
rect 447 301 448 302 
<< pdiffusion >>
rect 448 301 449 302 
<< pdiffusion >>
rect 449 301 450 302 
<< pdiffusion >>
rect 462 301 463 302 
<< pdiffusion >>
rect 463 301 464 302 
<< pdiffusion >>
rect 464 301 465 302 
<< pdiffusion >>
rect 465 301 466 302 
<< pdiffusion >>
rect 466 301 467 302 
<< pdiffusion >>
rect 467 301 468 302 
<< pdiffusion >>
rect 480 301 481 302 
<< pdiffusion >>
rect 481 301 482 302 
<< pdiffusion >>
rect 482 301 483 302 
<< pdiffusion >>
rect 483 301 484 302 
<< pdiffusion >>
rect 484 301 485 302 
<< pdiffusion >>
rect 485 301 486 302 
<< m1 >>
rect 487 301 488 302 
<< pdiffusion >>
rect 498 301 499 302 
<< pdiffusion >>
rect 499 301 500 302 
<< pdiffusion >>
rect 500 301 501 302 
<< pdiffusion >>
rect 501 301 502 302 
<< pdiffusion >>
rect 502 301 503 302 
<< pdiffusion >>
rect 503 301 504 302 
<< m1 >>
rect 523 301 524 302 
<< pdiffusion >>
rect 12 302 13 303 
<< pdiffusion >>
rect 13 302 14 303 
<< pdiffusion >>
rect 14 302 15 303 
<< pdiffusion >>
rect 15 302 16 303 
<< pdiffusion >>
rect 16 302 17 303 
<< pdiffusion >>
rect 17 302 18 303 
<< m1 >>
rect 19 302 20 303 
<< m1 >>
rect 22 302 23 303 
<< pdiffusion >>
rect 30 302 31 303 
<< pdiffusion >>
rect 31 302 32 303 
<< pdiffusion >>
rect 32 302 33 303 
<< pdiffusion >>
rect 33 302 34 303 
<< pdiffusion >>
rect 34 302 35 303 
<< pdiffusion >>
rect 35 302 36 303 
<< m1 >>
rect 44 302 45 303 
<< m1 >>
rect 46 302 47 303 
<< m2 >>
rect 46 302 47 303 
<< pdiffusion >>
rect 48 302 49 303 
<< pdiffusion >>
rect 49 302 50 303 
<< pdiffusion >>
rect 50 302 51 303 
<< pdiffusion >>
rect 51 302 52 303 
<< pdiffusion >>
rect 52 302 53 303 
<< pdiffusion >>
rect 53 302 54 303 
<< m1 >>
rect 55 302 56 303 
<< pdiffusion >>
rect 66 302 67 303 
<< pdiffusion >>
rect 67 302 68 303 
<< pdiffusion >>
rect 68 302 69 303 
<< pdiffusion >>
rect 69 302 70 303 
<< pdiffusion >>
rect 70 302 71 303 
<< pdiffusion >>
rect 71 302 72 303 
<< m1 >>
rect 73 302 74 303 
<< m2 >>
rect 74 302 75 303 
<< pdiffusion >>
rect 84 302 85 303 
<< pdiffusion >>
rect 85 302 86 303 
<< pdiffusion >>
rect 86 302 87 303 
<< pdiffusion >>
rect 87 302 88 303 
<< pdiffusion >>
rect 88 302 89 303 
<< pdiffusion >>
rect 89 302 90 303 
<< m1 >>
rect 91 302 92 303 
<< m1 >>
rect 93 302 94 303 
<< pdiffusion >>
rect 102 302 103 303 
<< pdiffusion >>
rect 103 302 104 303 
<< pdiffusion >>
rect 104 302 105 303 
<< pdiffusion >>
rect 105 302 106 303 
<< pdiffusion >>
rect 106 302 107 303 
<< pdiffusion >>
rect 107 302 108 303 
<< pdiffusion >>
rect 120 302 121 303 
<< pdiffusion >>
rect 121 302 122 303 
<< pdiffusion >>
rect 122 302 123 303 
<< pdiffusion >>
rect 123 302 124 303 
<< pdiffusion >>
rect 124 302 125 303 
<< pdiffusion >>
rect 125 302 126 303 
<< pdiffusion >>
rect 138 302 139 303 
<< pdiffusion >>
rect 139 302 140 303 
<< pdiffusion >>
rect 140 302 141 303 
<< pdiffusion >>
rect 141 302 142 303 
<< pdiffusion >>
rect 142 302 143 303 
<< pdiffusion >>
rect 143 302 144 303 
<< m1 >>
rect 146 302 147 303 
<< m1 >>
rect 148 302 149 303 
<< m1 >>
rect 150 302 151 303 
<< pdiffusion >>
rect 156 302 157 303 
<< pdiffusion >>
rect 157 302 158 303 
<< pdiffusion >>
rect 158 302 159 303 
<< pdiffusion >>
rect 159 302 160 303 
<< pdiffusion >>
rect 160 302 161 303 
<< pdiffusion >>
rect 161 302 162 303 
<< pdiffusion >>
rect 174 302 175 303 
<< pdiffusion >>
rect 175 302 176 303 
<< pdiffusion >>
rect 176 302 177 303 
<< pdiffusion >>
rect 177 302 178 303 
<< pdiffusion >>
rect 178 302 179 303 
<< pdiffusion >>
rect 179 302 180 303 
<< m1 >>
rect 181 302 182 303 
<< m1 >>
rect 186 302 187 303 
<< pdiffusion >>
rect 192 302 193 303 
<< pdiffusion >>
rect 193 302 194 303 
<< pdiffusion >>
rect 194 302 195 303 
<< pdiffusion >>
rect 195 302 196 303 
<< pdiffusion >>
rect 196 302 197 303 
<< pdiffusion >>
rect 197 302 198 303 
<< m1 >>
rect 208 302 209 303 
<< pdiffusion >>
rect 210 302 211 303 
<< pdiffusion >>
rect 211 302 212 303 
<< pdiffusion >>
rect 212 302 213 303 
<< pdiffusion >>
rect 213 302 214 303 
<< pdiffusion >>
rect 214 302 215 303 
<< pdiffusion >>
rect 215 302 216 303 
<< m1 >>
rect 217 302 218 303 
<< m2 >>
rect 218 302 219 303 
<< pdiffusion >>
rect 228 302 229 303 
<< pdiffusion >>
rect 229 302 230 303 
<< pdiffusion >>
rect 230 302 231 303 
<< pdiffusion >>
rect 231 302 232 303 
<< pdiffusion >>
rect 232 302 233 303 
<< pdiffusion >>
rect 233 302 234 303 
<< m1 >>
rect 237 302 238 303 
<< m2 >>
rect 243 302 244 303 
<< m1 >>
rect 244 302 245 303 
<< pdiffusion >>
rect 246 302 247 303 
<< pdiffusion >>
rect 247 302 248 303 
<< pdiffusion >>
rect 248 302 249 303 
<< pdiffusion >>
rect 249 302 250 303 
<< pdiffusion >>
rect 250 302 251 303 
<< pdiffusion >>
rect 251 302 252 303 
<< m1 >>
rect 255 302 256 303 
<< pdiffusion >>
rect 264 302 265 303 
<< pdiffusion >>
rect 265 302 266 303 
<< pdiffusion >>
rect 266 302 267 303 
<< pdiffusion >>
rect 267 302 268 303 
<< pdiffusion >>
rect 268 302 269 303 
<< pdiffusion >>
rect 269 302 270 303 
<< m1 >>
rect 271 302 272 303 
<< m2 >>
rect 277 302 278 303 
<< m1 >>
rect 278 302 279 303 
<< m1 >>
rect 280 302 281 303 
<< pdiffusion >>
rect 282 302 283 303 
<< pdiffusion >>
rect 283 302 284 303 
<< pdiffusion >>
rect 284 302 285 303 
<< pdiffusion >>
rect 285 302 286 303 
<< pdiffusion >>
rect 286 302 287 303 
<< pdiffusion >>
rect 287 302 288 303 
<< pdiffusion >>
rect 300 302 301 303 
<< pdiffusion >>
rect 301 302 302 303 
<< pdiffusion >>
rect 302 302 303 303 
<< pdiffusion >>
rect 303 302 304 303 
<< pdiffusion >>
rect 304 302 305 303 
<< pdiffusion >>
rect 305 302 306 303 
<< m1 >>
rect 307 302 308 303 
<< m1 >>
rect 309 302 310 303 
<< m2 >>
rect 310 302 311 303 
<< pdiffusion >>
rect 318 302 319 303 
<< pdiffusion >>
rect 319 302 320 303 
<< pdiffusion >>
rect 320 302 321 303 
<< pdiffusion >>
rect 321 302 322 303 
<< pdiffusion >>
rect 322 302 323 303 
<< pdiffusion >>
rect 323 302 324 303 
<< m2 >>
rect 333 302 334 303 
<< m1 >>
rect 334 302 335 303 
<< pdiffusion >>
rect 336 302 337 303 
<< pdiffusion >>
rect 337 302 338 303 
<< pdiffusion >>
rect 338 302 339 303 
<< pdiffusion >>
rect 339 302 340 303 
<< pdiffusion >>
rect 340 302 341 303 
<< pdiffusion >>
rect 341 302 342 303 
<< m1 >>
rect 344 302 345 303 
<< m2 >>
rect 345 302 346 303 
<< m1 >>
rect 348 302 349 303 
<< m1 >>
rect 352 302 353 303 
<< pdiffusion >>
rect 354 302 355 303 
<< pdiffusion >>
rect 355 302 356 303 
<< pdiffusion >>
rect 356 302 357 303 
<< pdiffusion >>
rect 357 302 358 303 
<< pdiffusion >>
rect 358 302 359 303 
<< pdiffusion >>
rect 359 302 360 303 
<< m1 >>
rect 366 302 367 303 
<< m1 >>
rect 370 302 371 303 
<< pdiffusion >>
rect 372 302 373 303 
<< pdiffusion >>
rect 373 302 374 303 
<< pdiffusion >>
rect 374 302 375 303 
<< pdiffusion >>
rect 375 302 376 303 
<< pdiffusion >>
rect 376 302 377 303 
<< pdiffusion >>
rect 377 302 378 303 
<< m1 >>
rect 379 302 380 303 
<< m2 >>
rect 380 302 381 303 
<< m1 >>
rect 381 302 382 303 
<< pdiffusion >>
rect 390 302 391 303 
<< pdiffusion >>
rect 391 302 392 303 
<< pdiffusion >>
rect 392 302 393 303 
<< pdiffusion >>
rect 393 302 394 303 
<< pdiffusion >>
rect 394 302 395 303 
<< pdiffusion >>
rect 395 302 396 303 
<< m1 >>
rect 406 302 407 303 
<< pdiffusion >>
rect 408 302 409 303 
<< pdiffusion >>
rect 409 302 410 303 
<< pdiffusion >>
rect 410 302 411 303 
<< pdiffusion >>
rect 411 302 412 303 
<< pdiffusion >>
rect 412 302 413 303 
<< pdiffusion >>
rect 413 302 414 303 
<< m1 >>
rect 416 302 417 303 
<< m2 >>
rect 419 302 420 303 
<< m1 >>
rect 420 302 421 303 
<< m1 >>
rect 422 302 423 303 
<< pdiffusion >>
rect 426 302 427 303 
<< pdiffusion >>
rect 427 302 428 303 
<< pdiffusion >>
rect 428 302 429 303 
<< pdiffusion >>
rect 429 302 430 303 
<< pdiffusion >>
rect 430 302 431 303 
<< pdiffusion >>
rect 431 302 432 303 
<< m1 >>
rect 433 302 434 303 
<< m2 >>
rect 434 302 435 303 
<< m1 >>
rect 437 302 438 303 
<< pdiffusion >>
rect 444 302 445 303 
<< pdiffusion >>
rect 445 302 446 303 
<< pdiffusion >>
rect 446 302 447 303 
<< pdiffusion >>
rect 447 302 448 303 
<< pdiffusion >>
rect 448 302 449 303 
<< pdiffusion >>
rect 449 302 450 303 
<< pdiffusion >>
rect 462 302 463 303 
<< pdiffusion >>
rect 463 302 464 303 
<< pdiffusion >>
rect 464 302 465 303 
<< pdiffusion >>
rect 465 302 466 303 
<< pdiffusion >>
rect 466 302 467 303 
<< pdiffusion >>
rect 467 302 468 303 
<< pdiffusion >>
rect 480 302 481 303 
<< pdiffusion >>
rect 481 302 482 303 
<< pdiffusion >>
rect 482 302 483 303 
<< pdiffusion >>
rect 483 302 484 303 
<< pdiffusion >>
rect 484 302 485 303 
<< pdiffusion >>
rect 485 302 486 303 
<< m1 >>
rect 487 302 488 303 
<< pdiffusion >>
rect 498 302 499 303 
<< pdiffusion >>
rect 499 302 500 303 
<< pdiffusion >>
rect 500 302 501 303 
<< pdiffusion >>
rect 501 302 502 303 
<< pdiffusion >>
rect 502 302 503 303 
<< pdiffusion >>
rect 503 302 504 303 
<< m1 >>
rect 523 302 524 303 
<< pdiffusion >>
rect 12 303 13 304 
<< pdiffusion >>
rect 13 303 14 304 
<< pdiffusion >>
rect 14 303 15 304 
<< pdiffusion >>
rect 15 303 16 304 
<< pdiffusion >>
rect 16 303 17 304 
<< pdiffusion >>
rect 17 303 18 304 
<< m1 >>
rect 19 303 20 304 
<< m1 >>
rect 22 303 23 304 
<< pdiffusion >>
rect 30 303 31 304 
<< pdiffusion >>
rect 31 303 32 304 
<< pdiffusion >>
rect 32 303 33 304 
<< pdiffusion >>
rect 33 303 34 304 
<< pdiffusion >>
rect 34 303 35 304 
<< pdiffusion >>
rect 35 303 36 304 
<< m1 >>
rect 44 303 45 304 
<< m1 >>
rect 46 303 47 304 
<< m2 >>
rect 46 303 47 304 
<< pdiffusion >>
rect 48 303 49 304 
<< pdiffusion >>
rect 49 303 50 304 
<< pdiffusion >>
rect 50 303 51 304 
<< pdiffusion >>
rect 51 303 52 304 
<< pdiffusion >>
rect 52 303 53 304 
<< pdiffusion >>
rect 53 303 54 304 
<< m1 >>
rect 55 303 56 304 
<< pdiffusion >>
rect 66 303 67 304 
<< pdiffusion >>
rect 67 303 68 304 
<< pdiffusion >>
rect 68 303 69 304 
<< pdiffusion >>
rect 69 303 70 304 
<< pdiffusion >>
rect 70 303 71 304 
<< pdiffusion >>
rect 71 303 72 304 
<< m1 >>
rect 73 303 74 304 
<< m2 >>
rect 74 303 75 304 
<< pdiffusion >>
rect 84 303 85 304 
<< pdiffusion >>
rect 85 303 86 304 
<< pdiffusion >>
rect 86 303 87 304 
<< pdiffusion >>
rect 87 303 88 304 
<< pdiffusion >>
rect 88 303 89 304 
<< pdiffusion >>
rect 89 303 90 304 
<< m1 >>
rect 91 303 92 304 
<< m1 >>
rect 93 303 94 304 
<< pdiffusion >>
rect 102 303 103 304 
<< pdiffusion >>
rect 103 303 104 304 
<< pdiffusion >>
rect 104 303 105 304 
<< pdiffusion >>
rect 105 303 106 304 
<< pdiffusion >>
rect 106 303 107 304 
<< pdiffusion >>
rect 107 303 108 304 
<< pdiffusion >>
rect 120 303 121 304 
<< pdiffusion >>
rect 121 303 122 304 
<< pdiffusion >>
rect 122 303 123 304 
<< pdiffusion >>
rect 123 303 124 304 
<< pdiffusion >>
rect 124 303 125 304 
<< pdiffusion >>
rect 125 303 126 304 
<< pdiffusion >>
rect 138 303 139 304 
<< pdiffusion >>
rect 139 303 140 304 
<< pdiffusion >>
rect 140 303 141 304 
<< pdiffusion >>
rect 141 303 142 304 
<< pdiffusion >>
rect 142 303 143 304 
<< pdiffusion >>
rect 143 303 144 304 
<< m1 >>
rect 146 303 147 304 
<< m1 >>
rect 148 303 149 304 
<< m1 >>
rect 150 303 151 304 
<< pdiffusion >>
rect 156 303 157 304 
<< pdiffusion >>
rect 157 303 158 304 
<< pdiffusion >>
rect 158 303 159 304 
<< pdiffusion >>
rect 159 303 160 304 
<< pdiffusion >>
rect 160 303 161 304 
<< pdiffusion >>
rect 161 303 162 304 
<< pdiffusion >>
rect 174 303 175 304 
<< pdiffusion >>
rect 175 303 176 304 
<< pdiffusion >>
rect 176 303 177 304 
<< pdiffusion >>
rect 177 303 178 304 
<< pdiffusion >>
rect 178 303 179 304 
<< pdiffusion >>
rect 179 303 180 304 
<< m1 >>
rect 181 303 182 304 
<< m1 >>
rect 186 303 187 304 
<< pdiffusion >>
rect 192 303 193 304 
<< pdiffusion >>
rect 193 303 194 304 
<< pdiffusion >>
rect 194 303 195 304 
<< pdiffusion >>
rect 195 303 196 304 
<< pdiffusion >>
rect 196 303 197 304 
<< pdiffusion >>
rect 197 303 198 304 
<< m1 >>
rect 208 303 209 304 
<< pdiffusion >>
rect 210 303 211 304 
<< pdiffusion >>
rect 211 303 212 304 
<< pdiffusion >>
rect 212 303 213 304 
<< pdiffusion >>
rect 213 303 214 304 
<< pdiffusion >>
rect 214 303 215 304 
<< pdiffusion >>
rect 215 303 216 304 
<< m1 >>
rect 217 303 218 304 
<< m2 >>
rect 218 303 219 304 
<< pdiffusion >>
rect 228 303 229 304 
<< pdiffusion >>
rect 229 303 230 304 
<< pdiffusion >>
rect 230 303 231 304 
<< pdiffusion >>
rect 231 303 232 304 
<< pdiffusion >>
rect 232 303 233 304 
<< pdiffusion >>
rect 233 303 234 304 
<< m1 >>
rect 237 303 238 304 
<< m2 >>
rect 237 303 238 304 
<< m2c >>
rect 237 303 238 304 
<< m1 >>
rect 237 303 238 304 
<< m2 >>
rect 237 303 238 304 
<< m2 >>
rect 243 303 244 304 
<< m1 >>
rect 244 303 245 304 
<< pdiffusion >>
rect 246 303 247 304 
<< pdiffusion >>
rect 247 303 248 304 
<< pdiffusion >>
rect 248 303 249 304 
<< pdiffusion >>
rect 249 303 250 304 
<< pdiffusion >>
rect 250 303 251 304 
<< pdiffusion >>
rect 251 303 252 304 
<< m1 >>
rect 255 303 256 304 
<< pdiffusion >>
rect 264 303 265 304 
<< pdiffusion >>
rect 265 303 266 304 
<< pdiffusion >>
rect 266 303 267 304 
<< pdiffusion >>
rect 267 303 268 304 
<< pdiffusion >>
rect 268 303 269 304 
<< pdiffusion >>
rect 269 303 270 304 
<< m1 >>
rect 271 303 272 304 
<< m2 >>
rect 277 303 278 304 
<< m1 >>
rect 278 303 279 304 
<< m1 >>
rect 280 303 281 304 
<< pdiffusion >>
rect 282 303 283 304 
<< pdiffusion >>
rect 283 303 284 304 
<< pdiffusion >>
rect 284 303 285 304 
<< pdiffusion >>
rect 285 303 286 304 
<< pdiffusion >>
rect 286 303 287 304 
<< pdiffusion >>
rect 287 303 288 304 
<< pdiffusion >>
rect 300 303 301 304 
<< pdiffusion >>
rect 301 303 302 304 
<< pdiffusion >>
rect 302 303 303 304 
<< pdiffusion >>
rect 303 303 304 304 
<< pdiffusion >>
rect 304 303 305 304 
<< pdiffusion >>
rect 305 303 306 304 
<< m1 >>
rect 307 303 308 304 
<< m1 >>
rect 309 303 310 304 
<< m2 >>
rect 310 303 311 304 
<< pdiffusion >>
rect 318 303 319 304 
<< pdiffusion >>
rect 319 303 320 304 
<< pdiffusion >>
rect 320 303 321 304 
<< pdiffusion >>
rect 321 303 322 304 
<< pdiffusion >>
rect 322 303 323 304 
<< pdiffusion >>
rect 323 303 324 304 
<< m2 >>
rect 333 303 334 304 
<< m1 >>
rect 334 303 335 304 
<< pdiffusion >>
rect 336 303 337 304 
<< pdiffusion >>
rect 337 303 338 304 
<< pdiffusion >>
rect 338 303 339 304 
<< pdiffusion >>
rect 339 303 340 304 
<< pdiffusion >>
rect 340 303 341 304 
<< pdiffusion >>
rect 341 303 342 304 
<< m1 >>
rect 344 303 345 304 
<< m2 >>
rect 345 303 346 304 
<< m1 >>
rect 348 303 349 304 
<< m1 >>
rect 352 303 353 304 
<< pdiffusion >>
rect 354 303 355 304 
<< pdiffusion >>
rect 355 303 356 304 
<< pdiffusion >>
rect 356 303 357 304 
<< pdiffusion >>
rect 357 303 358 304 
<< pdiffusion >>
rect 358 303 359 304 
<< pdiffusion >>
rect 359 303 360 304 
<< m1 >>
rect 366 303 367 304 
<< m1 >>
rect 370 303 371 304 
<< pdiffusion >>
rect 372 303 373 304 
<< pdiffusion >>
rect 373 303 374 304 
<< pdiffusion >>
rect 374 303 375 304 
<< pdiffusion >>
rect 375 303 376 304 
<< pdiffusion >>
rect 376 303 377 304 
<< pdiffusion >>
rect 377 303 378 304 
<< m1 >>
rect 379 303 380 304 
<< m2 >>
rect 380 303 381 304 
<< m1 >>
rect 381 303 382 304 
<< pdiffusion >>
rect 390 303 391 304 
<< pdiffusion >>
rect 391 303 392 304 
<< pdiffusion >>
rect 392 303 393 304 
<< pdiffusion >>
rect 393 303 394 304 
<< pdiffusion >>
rect 394 303 395 304 
<< pdiffusion >>
rect 395 303 396 304 
<< m1 >>
rect 406 303 407 304 
<< pdiffusion >>
rect 408 303 409 304 
<< pdiffusion >>
rect 409 303 410 304 
<< pdiffusion >>
rect 410 303 411 304 
<< pdiffusion >>
rect 411 303 412 304 
<< pdiffusion >>
rect 412 303 413 304 
<< pdiffusion >>
rect 413 303 414 304 
<< m1 >>
rect 416 303 417 304 
<< m2 >>
rect 419 303 420 304 
<< m1 >>
rect 420 303 421 304 
<< m1 >>
rect 422 303 423 304 
<< pdiffusion >>
rect 426 303 427 304 
<< pdiffusion >>
rect 427 303 428 304 
<< pdiffusion >>
rect 428 303 429 304 
<< pdiffusion >>
rect 429 303 430 304 
<< pdiffusion >>
rect 430 303 431 304 
<< pdiffusion >>
rect 431 303 432 304 
<< m1 >>
rect 433 303 434 304 
<< m2 >>
rect 434 303 435 304 
<< m1 >>
rect 437 303 438 304 
<< pdiffusion >>
rect 444 303 445 304 
<< pdiffusion >>
rect 445 303 446 304 
<< pdiffusion >>
rect 446 303 447 304 
<< pdiffusion >>
rect 447 303 448 304 
<< pdiffusion >>
rect 448 303 449 304 
<< pdiffusion >>
rect 449 303 450 304 
<< pdiffusion >>
rect 462 303 463 304 
<< pdiffusion >>
rect 463 303 464 304 
<< pdiffusion >>
rect 464 303 465 304 
<< pdiffusion >>
rect 465 303 466 304 
<< pdiffusion >>
rect 466 303 467 304 
<< pdiffusion >>
rect 467 303 468 304 
<< pdiffusion >>
rect 480 303 481 304 
<< pdiffusion >>
rect 481 303 482 304 
<< pdiffusion >>
rect 482 303 483 304 
<< pdiffusion >>
rect 483 303 484 304 
<< pdiffusion >>
rect 484 303 485 304 
<< pdiffusion >>
rect 485 303 486 304 
<< m1 >>
rect 487 303 488 304 
<< pdiffusion >>
rect 498 303 499 304 
<< pdiffusion >>
rect 499 303 500 304 
<< pdiffusion >>
rect 500 303 501 304 
<< pdiffusion >>
rect 501 303 502 304 
<< pdiffusion >>
rect 502 303 503 304 
<< pdiffusion >>
rect 503 303 504 304 
<< m1 >>
rect 523 303 524 304 
<< pdiffusion >>
rect 12 304 13 305 
<< pdiffusion >>
rect 13 304 14 305 
<< pdiffusion >>
rect 14 304 15 305 
<< pdiffusion >>
rect 15 304 16 305 
<< pdiffusion >>
rect 16 304 17 305 
<< pdiffusion >>
rect 17 304 18 305 
<< m1 >>
rect 19 304 20 305 
<< m1 >>
rect 22 304 23 305 
<< pdiffusion >>
rect 30 304 31 305 
<< pdiffusion >>
rect 31 304 32 305 
<< pdiffusion >>
rect 32 304 33 305 
<< pdiffusion >>
rect 33 304 34 305 
<< pdiffusion >>
rect 34 304 35 305 
<< pdiffusion >>
rect 35 304 36 305 
<< m1 >>
rect 44 304 45 305 
<< m1 >>
rect 46 304 47 305 
<< m2 >>
rect 46 304 47 305 
<< pdiffusion >>
rect 48 304 49 305 
<< pdiffusion >>
rect 49 304 50 305 
<< pdiffusion >>
rect 50 304 51 305 
<< pdiffusion >>
rect 51 304 52 305 
<< pdiffusion >>
rect 52 304 53 305 
<< pdiffusion >>
rect 53 304 54 305 
<< m1 >>
rect 55 304 56 305 
<< pdiffusion >>
rect 66 304 67 305 
<< pdiffusion >>
rect 67 304 68 305 
<< pdiffusion >>
rect 68 304 69 305 
<< pdiffusion >>
rect 69 304 70 305 
<< pdiffusion >>
rect 70 304 71 305 
<< pdiffusion >>
rect 71 304 72 305 
<< m1 >>
rect 73 304 74 305 
<< m2 >>
rect 74 304 75 305 
<< pdiffusion >>
rect 84 304 85 305 
<< pdiffusion >>
rect 85 304 86 305 
<< pdiffusion >>
rect 86 304 87 305 
<< pdiffusion >>
rect 87 304 88 305 
<< pdiffusion >>
rect 88 304 89 305 
<< pdiffusion >>
rect 89 304 90 305 
<< m1 >>
rect 91 304 92 305 
<< m1 >>
rect 93 304 94 305 
<< pdiffusion >>
rect 102 304 103 305 
<< pdiffusion >>
rect 103 304 104 305 
<< pdiffusion >>
rect 104 304 105 305 
<< pdiffusion >>
rect 105 304 106 305 
<< pdiffusion >>
rect 106 304 107 305 
<< pdiffusion >>
rect 107 304 108 305 
<< pdiffusion >>
rect 120 304 121 305 
<< pdiffusion >>
rect 121 304 122 305 
<< pdiffusion >>
rect 122 304 123 305 
<< pdiffusion >>
rect 123 304 124 305 
<< pdiffusion >>
rect 124 304 125 305 
<< pdiffusion >>
rect 125 304 126 305 
<< pdiffusion >>
rect 138 304 139 305 
<< pdiffusion >>
rect 139 304 140 305 
<< pdiffusion >>
rect 140 304 141 305 
<< pdiffusion >>
rect 141 304 142 305 
<< pdiffusion >>
rect 142 304 143 305 
<< pdiffusion >>
rect 143 304 144 305 
<< m1 >>
rect 146 304 147 305 
<< m1 >>
rect 148 304 149 305 
<< m1 >>
rect 150 304 151 305 
<< pdiffusion >>
rect 156 304 157 305 
<< pdiffusion >>
rect 157 304 158 305 
<< pdiffusion >>
rect 158 304 159 305 
<< pdiffusion >>
rect 159 304 160 305 
<< pdiffusion >>
rect 160 304 161 305 
<< pdiffusion >>
rect 161 304 162 305 
<< pdiffusion >>
rect 174 304 175 305 
<< pdiffusion >>
rect 175 304 176 305 
<< pdiffusion >>
rect 176 304 177 305 
<< pdiffusion >>
rect 177 304 178 305 
<< pdiffusion >>
rect 178 304 179 305 
<< pdiffusion >>
rect 179 304 180 305 
<< m1 >>
rect 181 304 182 305 
<< m1 >>
rect 186 304 187 305 
<< pdiffusion >>
rect 192 304 193 305 
<< pdiffusion >>
rect 193 304 194 305 
<< pdiffusion >>
rect 194 304 195 305 
<< pdiffusion >>
rect 195 304 196 305 
<< pdiffusion >>
rect 196 304 197 305 
<< pdiffusion >>
rect 197 304 198 305 
<< m1 >>
rect 208 304 209 305 
<< pdiffusion >>
rect 210 304 211 305 
<< pdiffusion >>
rect 211 304 212 305 
<< pdiffusion >>
rect 212 304 213 305 
<< pdiffusion >>
rect 213 304 214 305 
<< pdiffusion >>
rect 214 304 215 305 
<< pdiffusion >>
rect 215 304 216 305 
<< m1 >>
rect 217 304 218 305 
<< m2 >>
rect 218 304 219 305 
<< pdiffusion >>
rect 228 304 229 305 
<< pdiffusion >>
rect 229 304 230 305 
<< pdiffusion >>
rect 230 304 231 305 
<< pdiffusion >>
rect 231 304 232 305 
<< pdiffusion >>
rect 232 304 233 305 
<< pdiffusion >>
rect 233 304 234 305 
<< m2 >>
rect 237 304 238 305 
<< m2 >>
rect 243 304 244 305 
<< m1 >>
rect 244 304 245 305 
<< pdiffusion >>
rect 246 304 247 305 
<< pdiffusion >>
rect 247 304 248 305 
<< pdiffusion >>
rect 248 304 249 305 
<< pdiffusion >>
rect 249 304 250 305 
<< pdiffusion >>
rect 250 304 251 305 
<< pdiffusion >>
rect 251 304 252 305 
<< m1 >>
rect 255 304 256 305 
<< pdiffusion >>
rect 264 304 265 305 
<< pdiffusion >>
rect 265 304 266 305 
<< pdiffusion >>
rect 266 304 267 305 
<< pdiffusion >>
rect 267 304 268 305 
<< pdiffusion >>
rect 268 304 269 305 
<< pdiffusion >>
rect 269 304 270 305 
<< m1 >>
rect 271 304 272 305 
<< m2 >>
rect 277 304 278 305 
<< m1 >>
rect 278 304 279 305 
<< m1 >>
rect 280 304 281 305 
<< pdiffusion >>
rect 282 304 283 305 
<< pdiffusion >>
rect 283 304 284 305 
<< pdiffusion >>
rect 284 304 285 305 
<< pdiffusion >>
rect 285 304 286 305 
<< pdiffusion >>
rect 286 304 287 305 
<< pdiffusion >>
rect 287 304 288 305 
<< pdiffusion >>
rect 300 304 301 305 
<< pdiffusion >>
rect 301 304 302 305 
<< pdiffusion >>
rect 302 304 303 305 
<< pdiffusion >>
rect 303 304 304 305 
<< pdiffusion >>
rect 304 304 305 305 
<< pdiffusion >>
rect 305 304 306 305 
<< m1 >>
rect 307 304 308 305 
<< m1 >>
rect 309 304 310 305 
<< m2 >>
rect 310 304 311 305 
<< pdiffusion >>
rect 318 304 319 305 
<< pdiffusion >>
rect 319 304 320 305 
<< pdiffusion >>
rect 320 304 321 305 
<< pdiffusion >>
rect 321 304 322 305 
<< pdiffusion >>
rect 322 304 323 305 
<< pdiffusion >>
rect 323 304 324 305 
<< m2 >>
rect 333 304 334 305 
<< m1 >>
rect 334 304 335 305 
<< pdiffusion >>
rect 336 304 337 305 
<< pdiffusion >>
rect 337 304 338 305 
<< pdiffusion >>
rect 338 304 339 305 
<< pdiffusion >>
rect 339 304 340 305 
<< pdiffusion >>
rect 340 304 341 305 
<< pdiffusion >>
rect 341 304 342 305 
<< m1 >>
rect 344 304 345 305 
<< m2 >>
rect 345 304 346 305 
<< m1 >>
rect 348 304 349 305 
<< m1 >>
rect 352 304 353 305 
<< pdiffusion >>
rect 354 304 355 305 
<< pdiffusion >>
rect 355 304 356 305 
<< pdiffusion >>
rect 356 304 357 305 
<< pdiffusion >>
rect 357 304 358 305 
<< pdiffusion >>
rect 358 304 359 305 
<< pdiffusion >>
rect 359 304 360 305 
<< m1 >>
rect 366 304 367 305 
<< m1 >>
rect 370 304 371 305 
<< pdiffusion >>
rect 372 304 373 305 
<< pdiffusion >>
rect 373 304 374 305 
<< pdiffusion >>
rect 374 304 375 305 
<< pdiffusion >>
rect 375 304 376 305 
<< pdiffusion >>
rect 376 304 377 305 
<< pdiffusion >>
rect 377 304 378 305 
<< m1 >>
rect 379 304 380 305 
<< m2 >>
rect 380 304 381 305 
<< m1 >>
rect 381 304 382 305 
<< pdiffusion >>
rect 390 304 391 305 
<< pdiffusion >>
rect 391 304 392 305 
<< pdiffusion >>
rect 392 304 393 305 
<< pdiffusion >>
rect 393 304 394 305 
<< pdiffusion >>
rect 394 304 395 305 
<< pdiffusion >>
rect 395 304 396 305 
<< m1 >>
rect 406 304 407 305 
<< pdiffusion >>
rect 408 304 409 305 
<< pdiffusion >>
rect 409 304 410 305 
<< pdiffusion >>
rect 410 304 411 305 
<< pdiffusion >>
rect 411 304 412 305 
<< pdiffusion >>
rect 412 304 413 305 
<< pdiffusion >>
rect 413 304 414 305 
<< m1 >>
rect 416 304 417 305 
<< m2 >>
rect 419 304 420 305 
<< m1 >>
rect 420 304 421 305 
<< m1 >>
rect 422 304 423 305 
<< pdiffusion >>
rect 426 304 427 305 
<< pdiffusion >>
rect 427 304 428 305 
<< pdiffusion >>
rect 428 304 429 305 
<< pdiffusion >>
rect 429 304 430 305 
<< pdiffusion >>
rect 430 304 431 305 
<< pdiffusion >>
rect 431 304 432 305 
<< m1 >>
rect 433 304 434 305 
<< m2 >>
rect 434 304 435 305 
<< m1 >>
rect 437 304 438 305 
<< pdiffusion >>
rect 444 304 445 305 
<< pdiffusion >>
rect 445 304 446 305 
<< pdiffusion >>
rect 446 304 447 305 
<< pdiffusion >>
rect 447 304 448 305 
<< pdiffusion >>
rect 448 304 449 305 
<< pdiffusion >>
rect 449 304 450 305 
<< pdiffusion >>
rect 462 304 463 305 
<< pdiffusion >>
rect 463 304 464 305 
<< pdiffusion >>
rect 464 304 465 305 
<< pdiffusion >>
rect 465 304 466 305 
<< pdiffusion >>
rect 466 304 467 305 
<< pdiffusion >>
rect 467 304 468 305 
<< pdiffusion >>
rect 480 304 481 305 
<< pdiffusion >>
rect 481 304 482 305 
<< pdiffusion >>
rect 482 304 483 305 
<< pdiffusion >>
rect 483 304 484 305 
<< pdiffusion >>
rect 484 304 485 305 
<< pdiffusion >>
rect 485 304 486 305 
<< m1 >>
rect 487 304 488 305 
<< pdiffusion >>
rect 498 304 499 305 
<< pdiffusion >>
rect 499 304 500 305 
<< pdiffusion >>
rect 500 304 501 305 
<< pdiffusion >>
rect 501 304 502 305 
<< pdiffusion >>
rect 502 304 503 305 
<< pdiffusion >>
rect 503 304 504 305 
<< m1 >>
rect 523 304 524 305 
<< pdiffusion >>
rect 12 305 13 306 
<< pdiffusion >>
rect 13 305 14 306 
<< pdiffusion >>
rect 14 305 15 306 
<< pdiffusion >>
rect 15 305 16 306 
<< pdiffusion >>
rect 16 305 17 306 
<< pdiffusion >>
rect 17 305 18 306 
<< m1 >>
rect 19 305 20 306 
<< m1 >>
rect 22 305 23 306 
<< pdiffusion >>
rect 30 305 31 306 
<< pdiffusion >>
rect 31 305 32 306 
<< pdiffusion >>
rect 32 305 33 306 
<< pdiffusion >>
rect 33 305 34 306 
<< pdiffusion >>
rect 34 305 35 306 
<< pdiffusion >>
rect 35 305 36 306 
<< m1 >>
rect 44 305 45 306 
<< m1 >>
rect 46 305 47 306 
<< m2 >>
rect 46 305 47 306 
<< pdiffusion >>
rect 48 305 49 306 
<< pdiffusion >>
rect 49 305 50 306 
<< pdiffusion >>
rect 50 305 51 306 
<< pdiffusion >>
rect 51 305 52 306 
<< pdiffusion >>
rect 52 305 53 306 
<< pdiffusion >>
rect 53 305 54 306 
<< m1 >>
rect 55 305 56 306 
<< pdiffusion >>
rect 66 305 67 306 
<< pdiffusion >>
rect 67 305 68 306 
<< pdiffusion >>
rect 68 305 69 306 
<< pdiffusion >>
rect 69 305 70 306 
<< pdiffusion >>
rect 70 305 71 306 
<< pdiffusion >>
rect 71 305 72 306 
<< m1 >>
rect 73 305 74 306 
<< m2 >>
rect 74 305 75 306 
<< pdiffusion >>
rect 84 305 85 306 
<< m1 >>
rect 85 305 86 306 
<< pdiffusion >>
rect 85 305 86 306 
<< pdiffusion >>
rect 86 305 87 306 
<< pdiffusion >>
rect 87 305 88 306 
<< pdiffusion >>
rect 88 305 89 306 
<< pdiffusion >>
rect 89 305 90 306 
<< m1 >>
rect 91 305 92 306 
<< m1 >>
rect 93 305 94 306 
<< pdiffusion >>
rect 102 305 103 306 
<< m1 >>
rect 103 305 104 306 
<< pdiffusion >>
rect 103 305 104 306 
<< pdiffusion >>
rect 104 305 105 306 
<< pdiffusion >>
rect 105 305 106 306 
<< pdiffusion >>
rect 106 305 107 306 
<< pdiffusion >>
rect 107 305 108 306 
<< pdiffusion >>
rect 120 305 121 306 
<< pdiffusion >>
rect 121 305 122 306 
<< pdiffusion >>
rect 122 305 123 306 
<< pdiffusion >>
rect 123 305 124 306 
<< pdiffusion >>
rect 124 305 125 306 
<< pdiffusion >>
rect 125 305 126 306 
<< pdiffusion >>
rect 138 305 139 306 
<< pdiffusion >>
rect 139 305 140 306 
<< pdiffusion >>
rect 140 305 141 306 
<< pdiffusion >>
rect 141 305 142 306 
<< pdiffusion >>
rect 142 305 143 306 
<< pdiffusion >>
rect 143 305 144 306 
<< m1 >>
rect 146 305 147 306 
<< m1 >>
rect 148 305 149 306 
<< m1 >>
rect 150 305 151 306 
<< pdiffusion >>
rect 156 305 157 306 
<< pdiffusion >>
rect 157 305 158 306 
<< pdiffusion >>
rect 158 305 159 306 
<< pdiffusion >>
rect 159 305 160 306 
<< pdiffusion >>
rect 160 305 161 306 
<< pdiffusion >>
rect 161 305 162 306 
<< pdiffusion >>
rect 174 305 175 306 
<< pdiffusion >>
rect 175 305 176 306 
<< pdiffusion >>
rect 176 305 177 306 
<< pdiffusion >>
rect 177 305 178 306 
<< m1 >>
rect 178 305 179 306 
<< pdiffusion >>
rect 178 305 179 306 
<< pdiffusion >>
rect 179 305 180 306 
<< m1 >>
rect 181 305 182 306 
<< m1 >>
rect 186 305 187 306 
<< pdiffusion >>
rect 192 305 193 306 
<< m1 >>
rect 193 305 194 306 
<< pdiffusion >>
rect 193 305 194 306 
<< pdiffusion >>
rect 194 305 195 306 
<< pdiffusion >>
rect 195 305 196 306 
<< pdiffusion >>
rect 196 305 197 306 
<< pdiffusion >>
rect 197 305 198 306 
<< m1 >>
rect 208 305 209 306 
<< pdiffusion >>
rect 210 305 211 306 
<< m1 >>
rect 211 305 212 306 
<< pdiffusion >>
rect 211 305 212 306 
<< pdiffusion >>
rect 212 305 213 306 
<< pdiffusion >>
rect 213 305 214 306 
<< pdiffusion >>
rect 214 305 215 306 
<< pdiffusion >>
rect 215 305 216 306 
<< m1 >>
rect 217 305 218 306 
<< m2 >>
rect 218 305 219 306 
<< pdiffusion >>
rect 228 305 229 306 
<< m1 >>
rect 229 305 230 306 
<< pdiffusion >>
rect 229 305 230 306 
<< pdiffusion >>
rect 230 305 231 306 
<< pdiffusion >>
rect 231 305 232 306 
<< m1 >>
rect 232 305 233 306 
<< pdiffusion >>
rect 232 305 233 306 
<< pdiffusion >>
rect 233 305 234 306 
<< m1 >>
rect 235 305 236 306 
<< m2 >>
rect 235 305 236 306 
<< m2c >>
rect 235 305 236 306 
<< m1 >>
rect 235 305 236 306 
<< m2 >>
rect 235 305 236 306 
<< m1 >>
rect 236 305 237 306 
<< m1 >>
rect 237 305 238 306 
<< m2 >>
rect 237 305 238 306 
<< m1 >>
rect 238 305 239 306 
<< m1 >>
rect 239 305 240 306 
<< m1 >>
rect 240 305 241 306 
<< m1 >>
rect 241 305 242 306 
<< m1 >>
rect 242 305 243 306 
<< m2 >>
rect 242 305 243 306 
<< m2c >>
rect 242 305 243 306 
<< m1 >>
rect 242 305 243 306 
<< m2 >>
rect 242 305 243 306 
<< m2 >>
rect 243 305 244 306 
<< m1 >>
rect 244 305 245 306 
<< pdiffusion >>
rect 246 305 247 306 
<< pdiffusion >>
rect 247 305 248 306 
<< pdiffusion >>
rect 248 305 249 306 
<< pdiffusion >>
rect 249 305 250 306 
<< m1 >>
rect 250 305 251 306 
<< pdiffusion >>
rect 250 305 251 306 
<< pdiffusion >>
rect 251 305 252 306 
<< m1 >>
rect 255 305 256 306 
<< pdiffusion >>
rect 264 305 265 306 
<< pdiffusion >>
rect 265 305 266 306 
<< pdiffusion >>
rect 266 305 267 306 
<< pdiffusion >>
rect 267 305 268 306 
<< pdiffusion >>
rect 268 305 269 306 
<< pdiffusion >>
rect 269 305 270 306 
<< m1 >>
rect 271 305 272 306 
<< m2 >>
rect 277 305 278 306 
<< m1 >>
rect 278 305 279 306 
<< m1 >>
rect 280 305 281 306 
<< pdiffusion >>
rect 282 305 283 306 
<< pdiffusion >>
rect 283 305 284 306 
<< pdiffusion >>
rect 284 305 285 306 
<< pdiffusion >>
rect 285 305 286 306 
<< pdiffusion >>
rect 286 305 287 306 
<< pdiffusion >>
rect 287 305 288 306 
<< pdiffusion >>
rect 300 305 301 306 
<< pdiffusion >>
rect 301 305 302 306 
<< pdiffusion >>
rect 302 305 303 306 
<< pdiffusion >>
rect 303 305 304 306 
<< pdiffusion >>
rect 304 305 305 306 
<< pdiffusion >>
rect 305 305 306 306 
<< m1 >>
rect 307 305 308 306 
<< m1 >>
rect 309 305 310 306 
<< m2 >>
rect 310 305 311 306 
<< pdiffusion >>
rect 318 305 319 306 
<< pdiffusion >>
rect 319 305 320 306 
<< pdiffusion >>
rect 320 305 321 306 
<< pdiffusion >>
rect 321 305 322 306 
<< m1 >>
rect 322 305 323 306 
<< pdiffusion >>
rect 322 305 323 306 
<< pdiffusion >>
rect 323 305 324 306 
<< m2 >>
rect 333 305 334 306 
<< m1 >>
rect 334 305 335 306 
<< pdiffusion >>
rect 336 305 337 306 
<< pdiffusion >>
rect 337 305 338 306 
<< pdiffusion >>
rect 338 305 339 306 
<< pdiffusion >>
rect 339 305 340 306 
<< pdiffusion >>
rect 340 305 341 306 
<< pdiffusion >>
rect 341 305 342 306 
<< m1 >>
rect 344 305 345 306 
<< m2 >>
rect 345 305 346 306 
<< m1 >>
rect 348 305 349 306 
<< m1 >>
rect 352 305 353 306 
<< pdiffusion >>
rect 354 305 355 306 
<< pdiffusion >>
rect 355 305 356 306 
<< pdiffusion >>
rect 356 305 357 306 
<< pdiffusion >>
rect 357 305 358 306 
<< pdiffusion >>
rect 358 305 359 306 
<< pdiffusion >>
rect 359 305 360 306 
<< m1 >>
rect 366 305 367 306 
<< m1 >>
rect 370 305 371 306 
<< pdiffusion >>
rect 372 305 373 306 
<< pdiffusion >>
rect 373 305 374 306 
<< pdiffusion >>
rect 374 305 375 306 
<< pdiffusion >>
rect 375 305 376 306 
<< pdiffusion >>
rect 376 305 377 306 
<< pdiffusion >>
rect 377 305 378 306 
<< m1 >>
rect 379 305 380 306 
<< m2 >>
rect 380 305 381 306 
<< m1 >>
rect 381 305 382 306 
<< pdiffusion >>
rect 390 305 391 306 
<< pdiffusion >>
rect 391 305 392 306 
<< pdiffusion >>
rect 392 305 393 306 
<< pdiffusion >>
rect 393 305 394 306 
<< pdiffusion >>
rect 394 305 395 306 
<< pdiffusion >>
rect 395 305 396 306 
<< m1 >>
rect 406 305 407 306 
<< pdiffusion >>
rect 408 305 409 306 
<< pdiffusion >>
rect 409 305 410 306 
<< pdiffusion >>
rect 410 305 411 306 
<< pdiffusion >>
rect 411 305 412 306 
<< pdiffusion >>
rect 412 305 413 306 
<< pdiffusion >>
rect 413 305 414 306 
<< m1 >>
rect 416 305 417 306 
<< m2 >>
rect 419 305 420 306 
<< m1 >>
rect 420 305 421 306 
<< m1 >>
rect 422 305 423 306 
<< pdiffusion >>
rect 426 305 427 306 
<< m1 >>
rect 427 305 428 306 
<< pdiffusion >>
rect 427 305 428 306 
<< pdiffusion >>
rect 428 305 429 306 
<< pdiffusion >>
rect 429 305 430 306 
<< pdiffusion >>
rect 430 305 431 306 
<< pdiffusion >>
rect 431 305 432 306 
<< m1 >>
rect 433 305 434 306 
<< m2 >>
rect 434 305 435 306 
<< m1 >>
rect 437 305 438 306 
<< pdiffusion >>
rect 444 305 445 306 
<< pdiffusion >>
rect 445 305 446 306 
<< pdiffusion >>
rect 446 305 447 306 
<< pdiffusion >>
rect 447 305 448 306 
<< pdiffusion >>
rect 448 305 449 306 
<< pdiffusion >>
rect 449 305 450 306 
<< pdiffusion >>
rect 462 305 463 306 
<< pdiffusion >>
rect 463 305 464 306 
<< pdiffusion >>
rect 464 305 465 306 
<< pdiffusion >>
rect 465 305 466 306 
<< pdiffusion >>
rect 466 305 467 306 
<< pdiffusion >>
rect 467 305 468 306 
<< pdiffusion >>
rect 480 305 481 306 
<< pdiffusion >>
rect 481 305 482 306 
<< pdiffusion >>
rect 482 305 483 306 
<< pdiffusion >>
rect 483 305 484 306 
<< pdiffusion >>
rect 484 305 485 306 
<< pdiffusion >>
rect 485 305 486 306 
<< m1 >>
rect 487 305 488 306 
<< pdiffusion >>
rect 498 305 499 306 
<< pdiffusion >>
rect 499 305 500 306 
<< pdiffusion >>
rect 500 305 501 306 
<< pdiffusion >>
rect 501 305 502 306 
<< pdiffusion >>
rect 502 305 503 306 
<< pdiffusion >>
rect 503 305 504 306 
<< m1 >>
rect 523 305 524 306 
<< m1 >>
rect 19 306 20 307 
<< m1 >>
rect 22 306 23 307 
<< m1 >>
rect 44 306 45 307 
<< m1 >>
rect 46 306 47 307 
<< m2 >>
rect 46 306 47 307 
<< m1 >>
rect 55 306 56 307 
<< m1 >>
rect 73 306 74 307 
<< m2 >>
rect 74 306 75 307 
<< m1 >>
rect 85 306 86 307 
<< m1 >>
rect 91 306 92 307 
<< m1 >>
rect 93 306 94 307 
<< m1 >>
rect 103 306 104 307 
<< m1 >>
rect 146 306 147 307 
<< m1 >>
rect 148 306 149 307 
<< m1 >>
rect 150 306 151 307 
<< m1 >>
rect 178 306 179 307 
<< m1 >>
rect 181 306 182 307 
<< m1 >>
rect 186 306 187 307 
<< m1 >>
rect 193 306 194 307 
<< m1 >>
rect 208 306 209 307 
<< m1 >>
rect 211 306 212 307 
<< m1 >>
rect 217 306 218 307 
<< m2 >>
rect 218 306 219 307 
<< m1 >>
rect 229 306 230 307 
<< m1 >>
rect 232 306 233 307 
<< m2 >>
rect 235 306 236 307 
<< m2 >>
rect 237 306 238 307 
<< m1 >>
rect 244 306 245 307 
<< m1 >>
rect 250 306 251 307 
<< m1 >>
rect 255 306 256 307 
<< m1 >>
rect 271 306 272 307 
<< m1 >>
rect 273 306 274 307 
<< m1 >>
rect 274 306 275 307 
<< m1 >>
rect 275 306 276 307 
<< m1 >>
rect 276 306 277 307 
<< m2 >>
rect 276 306 277 307 
<< m2c >>
rect 276 306 277 307 
<< m1 >>
rect 276 306 277 307 
<< m2 >>
rect 276 306 277 307 
<< m2 >>
rect 277 306 278 307 
<< m1 >>
rect 278 306 279 307 
<< m1 >>
rect 280 306 281 307 
<< m1 >>
rect 307 306 308 307 
<< m2 >>
rect 307 306 308 307 
<< m2c >>
rect 307 306 308 307 
<< m1 >>
rect 307 306 308 307 
<< m2 >>
rect 307 306 308 307 
<< m1 >>
rect 309 306 310 307 
<< m2 >>
rect 310 306 311 307 
<< m1 >>
rect 322 306 323 307 
<< m2 >>
rect 333 306 334 307 
<< m1 >>
rect 334 306 335 307 
<< m1 >>
rect 344 306 345 307 
<< m2 >>
rect 345 306 346 307 
<< m1 >>
rect 346 306 347 307 
<< m2 >>
rect 346 306 347 307 
<< m2c >>
rect 346 306 347 307 
<< m1 >>
rect 346 306 347 307 
<< m2 >>
rect 346 306 347 307 
<< m1 >>
rect 348 306 349 307 
<< m1 >>
rect 352 306 353 307 
<< m1 >>
rect 366 306 367 307 
<< m1 >>
rect 370 306 371 307 
<< m1 >>
rect 379 306 380 307 
<< m2 >>
rect 380 306 381 307 
<< m1 >>
rect 381 306 382 307 
<< m2 >>
rect 381 306 382 307 
<< m2 >>
rect 382 306 383 307 
<< m1 >>
rect 383 306 384 307 
<< m2 >>
rect 383 306 384 307 
<< m2c >>
rect 383 306 384 307 
<< m1 >>
rect 383 306 384 307 
<< m2 >>
rect 383 306 384 307 
<< m1 >>
rect 384 306 385 307 
<< m1 >>
rect 385 306 386 307 
<< m1 >>
rect 386 306 387 307 
<< m1 >>
rect 387 306 388 307 
<< m1 >>
rect 388 306 389 307 
<< m1 >>
rect 406 306 407 307 
<< m1 >>
rect 416 306 417 307 
<< m2 >>
rect 419 306 420 307 
<< m1 >>
rect 420 306 421 307 
<< m2 >>
rect 420 306 421 307 
<< m2 >>
rect 421 306 422 307 
<< m1 >>
rect 422 306 423 307 
<< m2 >>
rect 422 306 423 307 
<< m2 >>
rect 423 306 424 307 
<< m2 >>
rect 424 306 425 307 
<< m1 >>
rect 427 306 428 307 
<< m1 >>
rect 433 306 434 307 
<< m2 >>
rect 434 306 435 307 
<< m1 >>
rect 437 306 438 307 
<< m1 >>
rect 487 306 488 307 
<< m1 >>
rect 523 306 524 307 
<< m1 >>
rect 19 307 20 308 
<< m1 >>
rect 22 307 23 308 
<< m1 >>
rect 44 307 45 308 
<< m1 >>
rect 46 307 47 308 
<< m2 >>
rect 46 307 47 308 
<< m1 >>
rect 55 307 56 308 
<< m1 >>
rect 73 307 74 308 
<< m2 >>
rect 74 307 75 308 
<< m1 >>
rect 85 307 86 308 
<< m1 >>
rect 91 307 92 308 
<< m1 >>
rect 93 307 94 308 
<< m1 >>
rect 100 307 101 308 
<< m1 >>
rect 101 307 102 308 
<< m1 >>
rect 102 307 103 308 
<< m1 >>
rect 103 307 104 308 
<< m1 >>
rect 146 307 147 308 
<< m1 >>
rect 148 307 149 308 
<< m1 >>
rect 150 307 151 308 
<< m1 >>
rect 178 307 179 308 
<< m1 >>
rect 181 307 182 308 
<< m1 >>
rect 186 307 187 308 
<< m1 >>
rect 193 307 194 308 
<< m2 >>
rect 207 307 208 308 
<< m1 >>
rect 208 307 209 308 
<< m2 >>
rect 208 307 209 308 
<< m2 >>
rect 209 307 210 308 
<< m1 >>
rect 210 307 211 308 
<< m2 >>
rect 210 307 211 308 
<< m2c >>
rect 210 307 211 308 
<< m1 >>
rect 210 307 211 308 
<< m2 >>
rect 210 307 211 308 
<< m1 >>
rect 211 307 212 308 
<< m1 >>
rect 217 307 218 308 
<< m2 >>
rect 218 307 219 308 
<< m1 >>
rect 229 307 230 308 
<< m1 >>
rect 232 307 233 308 
<< m1 >>
rect 233 307 234 308 
<< m1 >>
rect 234 307 235 308 
<< m1 >>
rect 235 307 236 308 
<< m2 >>
rect 235 307 236 308 
<< m1 >>
rect 236 307 237 308 
<< m1 >>
rect 237 307 238 308 
<< m2 >>
rect 237 307 238 308 
<< m1 >>
rect 238 307 239 308 
<< m1 >>
rect 239 307 240 308 
<< m1 >>
rect 240 307 241 308 
<< m1 >>
rect 241 307 242 308 
<< m1 >>
rect 242 307 243 308 
<< m2 >>
rect 242 307 243 308 
<< m2c >>
rect 242 307 243 308 
<< m1 >>
rect 242 307 243 308 
<< m2 >>
rect 242 307 243 308 
<< m2 >>
rect 243 307 244 308 
<< m1 >>
rect 244 307 245 308 
<< m2 >>
rect 244 307 245 308 
<< m2 >>
rect 245 307 246 308 
<< m1 >>
rect 246 307 247 308 
<< m2 >>
rect 246 307 247 308 
<< m2c >>
rect 246 307 247 308 
<< m1 >>
rect 246 307 247 308 
<< m2 >>
rect 246 307 247 308 
<< m1 >>
rect 250 307 251 308 
<< m1 >>
rect 251 307 252 308 
<< m1 >>
rect 252 307 253 308 
<< m1 >>
rect 253 307 254 308 
<< m1 >>
rect 255 307 256 308 
<< m1 >>
rect 271 307 272 308 
<< m1 >>
rect 273 307 274 308 
<< m1 >>
rect 278 307 279 308 
<< m1 >>
rect 280 307 281 308 
<< m2 >>
rect 307 307 308 308 
<< m1 >>
rect 309 307 310 308 
<< m2 >>
rect 310 307 311 308 
<< m1 >>
rect 322 307 323 308 
<< m1 >>
rect 323 307 324 308 
<< m1 >>
rect 324 307 325 308 
<< m1 >>
rect 325 307 326 308 
<< m1 >>
rect 326 307 327 308 
<< m1 >>
rect 327 307 328 308 
<< m1 >>
rect 328 307 329 308 
<< m1 >>
rect 329 307 330 308 
<< m1 >>
rect 330 307 331 308 
<< m1 >>
rect 331 307 332 308 
<< m1 >>
rect 332 307 333 308 
<< m2 >>
rect 332 307 333 308 
<< m2c >>
rect 332 307 333 308 
<< m1 >>
rect 332 307 333 308 
<< m2 >>
rect 332 307 333 308 
<< m2 >>
rect 333 307 334 308 
<< m1 >>
rect 334 307 335 308 
<< m1 >>
rect 344 307 345 308 
<< m1 >>
rect 346 307 347 308 
<< m1 >>
rect 348 307 349 308 
<< m1 >>
rect 352 307 353 308 
<< m1 >>
rect 366 307 367 308 
<< m1 >>
rect 370 307 371 308 
<< m1 >>
rect 379 307 380 308 
<< m1 >>
rect 381 307 382 308 
<< m1 >>
rect 388 307 389 308 
<< m1 >>
rect 406 307 407 308 
<< m1 >>
rect 416 307 417 308 
<< m1 >>
rect 420 307 421 308 
<< m1 >>
rect 422 307 423 308 
<< m1 >>
rect 423 307 424 308 
<< m1 >>
rect 424 307 425 308 
<< m2 >>
rect 424 307 425 308 
<< m1 >>
rect 425 307 426 308 
<< m1 >>
rect 426 307 427 308 
<< m1 >>
rect 427 307 428 308 
<< m1 >>
rect 431 307 432 308 
<< m2 >>
rect 431 307 432 308 
<< m2c >>
rect 431 307 432 308 
<< m1 >>
rect 431 307 432 308 
<< m2 >>
rect 431 307 432 308 
<< m2 >>
rect 432 307 433 308 
<< m1 >>
rect 433 307 434 308 
<< m2 >>
rect 433 307 434 308 
<< m2 >>
rect 434 307 435 308 
<< m1 >>
rect 437 307 438 308 
<< m1 >>
rect 487 307 488 308 
<< m1 >>
rect 523 307 524 308 
<< m1 >>
rect 19 308 20 309 
<< m1 >>
rect 22 308 23 309 
<< m1 >>
rect 44 308 45 309 
<< m1 >>
rect 46 308 47 309 
<< m2 >>
rect 46 308 47 309 
<< m1 >>
rect 55 308 56 309 
<< m1 >>
rect 73 308 74 309 
<< m2 >>
rect 74 308 75 309 
<< m1 >>
rect 85 308 86 309 
<< m1 >>
rect 86 308 87 309 
<< m1 >>
rect 87 308 88 309 
<< m1 >>
rect 88 308 89 309 
<< m1 >>
rect 89 308 90 309 
<< m1 >>
rect 90 308 91 309 
<< m1 >>
rect 91 308 92 309 
<< m1 >>
rect 93 308 94 309 
<< m1 >>
rect 100 308 101 309 
<< m1 >>
rect 146 308 147 309 
<< m2 >>
rect 146 308 147 309 
<< m2c >>
rect 146 308 147 309 
<< m1 >>
rect 146 308 147 309 
<< m2 >>
rect 146 308 147 309 
<< m1 >>
rect 148 308 149 309 
<< m2 >>
rect 148 308 149 309 
<< m2c >>
rect 148 308 149 309 
<< m1 >>
rect 148 308 149 309 
<< m2 >>
rect 148 308 149 309 
<< m1 >>
rect 150 308 151 309 
<< m2 >>
rect 150 308 151 309 
<< m2c >>
rect 150 308 151 309 
<< m1 >>
rect 150 308 151 309 
<< m2 >>
rect 150 308 151 309 
<< m1 >>
rect 178 308 179 309 
<< m2 >>
rect 178 308 179 309 
<< m2c >>
rect 178 308 179 309 
<< m1 >>
rect 178 308 179 309 
<< m2 >>
rect 178 308 179 309 
<< m1 >>
rect 180 308 181 309 
<< m2 >>
rect 180 308 181 309 
<< m2c >>
rect 180 308 181 309 
<< m1 >>
rect 180 308 181 309 
<< m2 >>
rect 180 308 181 309 
<< m1 >>
rect 181 308 182 309 
<< m1 >>
rect 186 308 187 309 
<< m2 >>
rect 186 308 187 309 
<< m2c >>
rect 186 308 187 309 
<< m1 >>
rect 186 308 187 309 
<< m2 >>
rect 186 308 187 309 
<< m1 >>
rect 193 308 194 309 
<< m2 >>
rect 207 308 208 309 
<< m1 >>
rect 208 308 209 309 
<< m1 >>
rect 217 308 218 309 
<< m2 >>
rect 218 308 219 309 
<< m1 >>
rect 229 308 230 309 
<< m2 >>
rect 230 308 231 309 
<< m2 >>
rect 231 308 232 309 
<< m2 >>
rect 232 308 233 309 
<< m2 >>
rect 233 308 234 309 
<< m2 >>
rect 234 308 235 309 
<< m2 >>
rect 235 308 236 309 
<< m2 >>
rect 237 308 238 309 
<< m1 >>
rect 244 308 245 309 
<< m1 >>
rect 246 308 247 309 
<< m2 >>
rect 249 308 250 309 
<< m2 >>
rect 250 308 251 309 
<< m2 >>
rect 251 308 252 309 
<< m2 >>
rect 252 308 253 309 
<< m1 >>
rect 253 308 254 309 
<< m2 >>
rect 253 308 254 309 
<< m2 >>
rect 254 308 255 309 
<< m1 >>
rect 255 308 256 309 
<< m2 >>
rect 255 308 256 309 
<< m2c >>
rect 255 308 256 309 
<< m1 >>
rect 255 308 256 309 
<< m2 >>
rect 255 308 256 309 
<< m1 >>
rect 266 308 267 309 
<< m2 >>
rect 266 308 267 309 
<< m2c >>
rect 266 308 267 309 
<< m1 >>
rect 266 308 267 309 
<< m2 >>
rect 266 308 267 309 
<< m1 >>
rect 267 308 268 309 
<< m1 >>
rect 268 308 269 309 
<< m1 >>
rect 269 308 270 309 
<< m2 >>
rect 269 308 270 309 
<< m2c >>
rect 269 308 270 309 
<< m1 >>
rect 269 308 270 309 
<< m2 >>
rect 269 308 270 309 
<< m2 >>
rect 270 308 271 309 
<< m1 >>
rect 271 308 272 309 
<< m2 >>
rect 271 308 272 309 
<< m2 >>
rect 272 308 273 309 
<< m1 >>
rect 273 308 274 309 
<< m2 >>
rect 273 308 274 309 
<< m2c >>
rect 273 308 274 309 
<< m1 >>
rect 273 308 274 309 
<< m2 >>
rect 273 308 274 309 
<< m1 >>
rect 278 308 279 309 
<< m2 >>
rect 278 308 279 309 
<< m2c >>
rect 278 308 279 309 
<< m1 >>
rect 278 308 279 309 
<< m2 >>
rect 278 308 279 309 
<< m1 >>
rect 280 308 281 309 
<< m2 >>
rect 280 308 281 309 
<< m2c >>
rect 280 308 281 309 
<< m1 >>
rect 280 308 281 309 
<< m2 >>
rect 280 308 281 309 
<< m1 >>
rect 302 308 303 309 
<< m2 >>
rect 302 308 303 309 
<< m2c >>
rect 302 308 303 309 
<< m1 >>
rect 302 308 303 309 
<< m2 >>
rect 302 308 303 309 
<< m1 >>
rect 303 308 304 309 
<< m1 >>
rect 304 308 305 309 
<< m1 >>
rect 305 308 306 309 
<< m1 >>
rect 306 308 307 309 
<< m1 >>
rect 307 308 308 309 
<< m2 >>
rect 307 308 308 309 
<< m1 >>
rect 308 308 309 309 
<< m1 >>
rect 309 308 310 309 
<< m2 >>
rect 310 308 311 309 
<< m1 >>
rect 334 308 335 309 
<< m1 >>
rect 344 308 345 309 
<< m2 >>
rect 344 308 345 309 
<< m2c >>
rect 344 308 345 309 
<< m1 >>
rect 344 308 345 309 
<< m2 >>
rect 344 308 345 309 
<< m1 >>
rect 346 308 347 309 
<< m2 >>
rect 346 308 347 309 
<< m2c >>
rect 346 308 347 309 
<< m1 >>
rect 346 308 347 309 
<< m2 >>
rect 346 308 347 309 
<< m1 >>
rect 348 308 349 309 
<< m2 >>
rect 348 308 349 309 
<< m2c >>
rect 348 308 349 309 
<< m1 >>
rect 348 308 349 309 
<< m2 >>
rect 348 308 349 309 
<< m1 >>
rect 352 308 353 309 
<< m1 >>
rect 366 308 367 309 
<< m2 >>
rect 366 308 367 309 
<< m2c >>
rect 366 308 367 309 
<< m1 >>
rect 366 308 367 309 
<< m2 >>
rect 366 308 367 309 
<< m1 >>
rect 370 308 371 309 
<< m1 >>
rect 374 308 375 309 
<< m2 >>
rect 374 308 375 309 
<< m2c >>
rect 374 308 375 309 
<< m1 >>
rect 374 308 375 309 
<< m2 >>
rect 374 308 375 309 
<< m1 >>
rect 375 308 376 309 
<< m1 >>
rect 376 308 377 309 
<< m1 >>
rect 377 308 378 309 
<< m2 >>
rect 377 308 378 309 
<< m2c >>
rect 377 308 378 309 
<< m1 >>
rect 377 308 378 309 
<< m2 >>
rect 377 308 378 309 
<< m2 >>
rect 378 308 379 309 
<< m1 >>
rect 379 308 380 309 
<< m2 >>
rect 379 308 380 309 
<< m2 >>
rect 380 308 381 309 
<< m1 >>
rect 381 308 382 309 
<< m2 >>
rect 381 308 382 309 
<< m2c >>
rect 381 308 382 309 
<< m1 >>
rect 381 308 382 309 
<< m2 >>
rect 381 308 382 309 
<< m1 >>
rect 388 308 389 309 
<< m1 >>
rect 389 308 390 309 
<< m1 >>
rect 390 308 391 309 
<< m2 >>
rect 390 308 391 309 
<< m2c >>
rect 390 308 391 309 
<< m1 >>
rect 390 308 391 309 
<< m2 >>
rect 390 308 391 309 
<< m1 >>
rect 406 308 407 309 
<< m1 >>
rect 416 308 417 309 
<< m1 >>
rect 420 308 421 309 
<< m2 >>
rect 424 308 425 309 
<< m1 >>
rect 429 308 430 309 
<< m2 >>
rect 429 308 430 309 
<< m2c >>
rect 429 308 430 309 
<< m1 >>
rect 429 308 430 309 
<< m2 >>
rect 429 308 430 309 
<< m1 >>
rect 430 308 431 309 
<< m1 >>
rect 431 308 432 309 
<< m1 >>
rect 433 308 434 309 
<< m1 >>
rect 437 308 438 309 
<< m1 >>
rect 487 308 488 309 
<< m1 >>
rect 523 308 524 309 
<< m1 >>
rect 19 309 20 310 
<< m1 >>
rect 22 309 23 310 
<< m1 >>
rect 44 309 45 310 
<< m1 >>
rect 46 309 47 310 
<< m2 >>
rect 46 309 47 310 
<< m1 >>
rect 55 309 56 310 
<< m1 >>
rect 73 309 74 310 
<< m2 >>
rect 74 309 75 310 
<< m1 >>
rect 93 309 94 310 
<< m1 >>
rect 100 309 101 310 
<< m2 >>
rect 146 309 147 310 
<< m2 >>
rect 148 309 149 310 
<< m2 >>
rect 150 309 151 310 
<< m2 >>
rect 178 309 179 310 
<< m2 >>
rect 180 309 181 310 
<< m2 >>
rect 186 309 187 310 
<< m1 >>
rect 193 309 194 310 
<< m2 >>
rect 207 309 208 310 
<< m1 >>
rect 208 309 209 310 
<< m1 >>
rect 217 309 218 310 
<< m2 >>
rect 218 309 219 310 
<< m1 >>
rect 229 309 230 310 
<< m2 >>
rect 230 309 231 310 
<< m1 >>
rect 237 309 238 310 
<< m2 >>
rect 237 309 238 310 
<< m2c >>
rect 237 309 238 310 
<< m1 >>
rect 237 309 238 310 
<< m2 >>
rect 237 309 238 310 
<< m1 >>
rect 244 309 245 310 
<< m1 >>
rect 246 309 247 310 
<< m2 >>
rect 249 309 250 310 
<< m1 >>
rect 253 309 254 310 
<< m2 >>
rect 266 309 267 310 
<< m1 >>
rect 271 309 272 310 
<< m2 >>
rect 278 309 279 310 
<< m2 >>
rect 280 309 281 310 
<< m2 >>
rect 302 309 303 310 
<< m2 >>
rect 307 309 308 310 
<< m2 >>
rect 310 309 311 310 
<< m1 >>
rect 334 309 335 310 
<< m2 >>
rect 344 309 345 310 
<< m2 >>
rect 346 309 347 310 
<< m2 >>
rect 348 309 349 310 
<< m1 >>
rect 352 309 353 310 
<< m2 >>
rect 366 309 367 310 
<< m1 >>
rect 370 309 371 310 
<< m2 >>
rect 374 309 375 310 
<< m1 >>
rect 379 309 380 310 
<< m2 >>
rect 390 309 391 310 
<< m1 >>
rect 406 309 407 310 
<< m1 >>
rect 416 309 417 310 
<< m1 >>
rect 420 309 421 310 
<< m2 >>
rect 424 309 425 310 
<< m2 >>
rect 429 309 430 310 
<< m1 >>
rect 433 309 434 310 
<< m1 >>
rect 437 309 438 310 
<< m1 >>
rect 487 309 488 310 
<< m1 >>
rect 523 309 524 310 
<< m1 >>
rect 19 310 20 311 
<< m1 >>
rect 22 310 23 311 
<< m1 >>
rect 44 310 45 311 
<< m1 >>
rect 46 310 47 311 
<< m2 >>
rect 46 310 47 311 
<< m1 >>
rect 55 310 56 311 
<< m1 >>
rect 73 310 74 311 
<< m2 >>
rect 74 310 75 311 
<< m1 >>
rect 93 310 94 311 
<< m1 >>
rect 100 310 101 311 
<< m1 >>
rect 121 310 122 311 
<< m1 >>
rect 122 310 123 311 
<< m1 >>
rect 123 310 124 311 
<< m1 >>
rect 124 310 125 311 
<< m1 >>
rect 125 310 126 311 
<< m1 >>
rect 126 310 127 311 
<< m1 >>
rect 127 310 128 311 
<< m1 >>
rect 128 310 129 311 
<< m1 >>
rect 129 310 130 311 
<< m1 >>
rect 130 310 131 311 
<< m1 >>
rect 131 310 132 311 
<< m1 >>
rect 132 310 133 311 
<< m1 >>
rect 133 310 134 311 
<< m1 >>
rect 134 310 135 311 
<< m1 >>
rect 135 310 136 311 
<< m1 >>
rect 136 310 137 311 
<< m1 >>
rect 137 310 138 311 
<< m1 >>
rect 138 310 139 311 
<< m1 >>
rect 139 310 140 311 
<< m1 >>
rect 140 310 141 311 
<< m1 >>
rect 141 310 142 311 
<< m1 >>
rect 142 310 143 311 
<< m1 >>
rect 143 310 144 311 
<< m1 >>
rect 144 310 145 311 
<< m1 >>
rect 145 310 146 311 
<< m1 >>
rect 146 310 147 311 
<< m2 >>
rect 146 310 147 311 
<< m1 >>
rect 147 310 148 311 
<< m1 >>
rect 148 310 149 311 
<< m2 >>
rect 148 310 149 311 
<< m1 >>
rect 149 310 150 311 
<< m1 >>
rect 150 310 151 311 
<< m2 >>
rect 150 310 151 311 
<< m1 >>
rect 151 310 152 311 
<< m1 >>
rect 152 310 153 311 
<< m2 >>
rect 152 310 153 311 
<< m2c >>
rect 152 310 153 311 
<< m1 >>
rect 152 310 153 311 
<< m2 >>
rect 152 310 153 311 
<< m2 >>
rect 153 310 154 311 
<< m1 >>
rect 154 310 155 311 
<< m2 >>
rect 154 310 155 311 
<< m1 >>
rect 155 310 156 311 
<< m2 >>
rect 155 310 156 311 
<< m1 >>
rect 156 310 157 311 
<< m2 >>
rect 156 310 157 311 
<< m1 >>
rect 157 310 158 311 
<< m2 >>
rect 157 310 158 311 
<< m1 >>
rect 158 310 159 311 
<< m2 >>
rect 158 310 159 311 
<< m1 >>
rect 159 310 160 311 
<< m2 >>
rect 159 310 160 311 
<< m1 >>
rect 160 310 161 311 
<< m2 >>
rect 160 310 161 311 
<< m1 >>
rect 161 310 162 311 
<< m2 >>
rect 161 310 162 311 
<< m1 >>
rect 162 310 163 311 
<< m2 >>
rect 162 310 163 311 
<< m1 >>
rect 163 310 164 311 
<< m2 >>
rect 163 310 164 311 
<< m1 >>
rect 164 310 165 311 
<< m2 >>
rect 164 310 165 311 
<< m1 >>
rect 165 310 166 311 
<< m2 >>
rect 165 310 166 311 
<< m1 >>
rect 166 310 167 311 
<< m2 >>
rect 166 310 167 311 
<< m1 >>
rect 167 310 168 311 
<< m2 >>
rect 167 310 168 311 
<< m1 >>
rect 168 310 169 311 
<< m2 >>
rect 168 310 169 311 
<< m1 >>
rect 169 310 170 311 
<< m2 >>
rect 169 310 170 311 
<< m1 >>
rect 170 310 171 311 
<< m2 >>
rect 170 310 171 311 
<< m1 >>
rect 171 310 172 311 
<< m2 >>
rect 171 310 172 311 
<< m1 >>
rect 172 310 173 311 
<< m2 >>
rect 172 310 173 311 
<< m1 >>
rect 173 310 174 311 
<< m2 >>
rect 173 310 174 311 
<< m1 >>
rect 174 310 175 311 
<< m2 >>
rect 174 310 175 311 
<< m1 >>
rect 175 310 176 311 
<< m2 >>
rect 175 310 176 311 
<< m1 >>
rect 176 310 177 311 
<< m2 >>
rect 176 310 177 311 
<< m1 >>
rect 177 310 178 311 
<< m2 >>
rect 177 310 178 311 
<< m1 >>
rect 178 310 179 311 
<< m2 >>
rect 178 310 179 311 
<< m1 >>
rect 179 310 180 311 
<< m1 >>
rect 180 310 181 311 
<< m2 >>
rect 180 310 181 311 
<< m1 >>
rect 181 310 182 311 
<< m1 >>
rect 182 310 183 311 
<< m1 >>
rect 183 310 184 311 
<< m1 >>
rect 184 310 185 311 
<< m1 >>
rect 185 310 186 311 
<< m1 >>
rect 186 310 187 311 
<< m2 >>
rect 186 310 187 311 
<< m1 >>
rect 187 310 188 311 
<< m1 >>
rect 188 310 189 311 
<< m1 >>
rect 189 310 190 311 
<< m1 >>
rect 190 310 191 311 
<< m1 >>
rect 191 310 192 311 
<< m1 >>
rect 192 310 193 311 
<< m1 >>
rect 193 310 194 311 
<< m2 >>
rect 207 310 208 311 
<< m1 >>
rect 208 310 209 311 
<< m1 >>
rect 217 310 218 311 
<< m2 >>
rect 218 310 219 311 
<< m1 >>
rect 229 310 230 311 
<< m2 >>
rect 230 310 231 311 
<< m1 >>
rect 237 310 238 311 
<< m1 >>
rect 244 310 245 311 
<< m1 >>
rect 246 310 247 311 
<< m1 >>
rect 247 310 248 311 
<< m1 >>
rect 248 310 249 311 
<< m1 >>
rect 249 310 250 311 
<< m2 >>
rect 249 310 250 311 
<< m1 >>
rect 250 310 251 311 
<< m1 >>
rect 251 310 252 311 
<< m2 >>
rect 251 310 252 311 
<< m2c >>
rect 251 310 252 311 
<< m1 >>
rect 251 310 252 311 
<< m2 >>
rect 251 310 252 311 
<< m2 >>
rect 252 310 253 311 
<< m1 >>
rect 253 310 254 311 
<< m2 >>
rect 253 310 254 311 
<< m2 >>
rect 254 310 255 311 
<< m1 >>
rect 255 310 256 311 
<< m2 >>
rect 255 310 256 311 
<< m2c >>
rect 255 310 256 311 
<< m1 >>
rect 255 310 256 311 
<< m2 >>
rect 255 310 256 311 
<< m1 >>
rect 256 310 257 311 
<< m1 >>
rect 257 310 258 311 
<< m1 >>
rect 258 310 259 311 
<< m1 >>
rect 259 310 260 311 
<< m1 >>
rect 260 310 261 311 
<< m1 >>
rect 261 310 262 311 
<< m1 >>
rect 262 310 263 311 
<< m1 >>
rect 263 310 264 311 
<< m1 >>
rect 264 310 265 311 
<< m1 >>
rect 265 310 266 311 
<< m1 >>
rect 266 310 267 311 
<< m2 >>
rect 266 310 267 311 
<< m1 >>
rect 267 310 268 311 
<< m1 >>
rect 268 310 269 311 
<< m1 >>
rect 269 310 270 311 
<< m2 >>
rect 269 310 270 311 
<< m2c >>
rect 269 310 270 311 
<< m1 >>
rect 269 310 270 311 
<< m2 >>
rect 269 310 270 311 
<< m2 >>
rect 270 310 271 311 
<< m1 >>
rect 271 310 272 311 
<< m2 >>
rect 271 310 272 311 
<< m2 >>
rect 272 310 273 311 
<< m1 >>
rect 273 310 274 311 
<< m2 >>
rect 273 310 274 311 
<< m2c >>
rect 273 310 274 311 
<< m1 >>
rect 273 310 274 311 
<< m2 >>
rect 273 310 274 311 
<< m1 >>
rect 274 310 275 311 
<< m1 >>
rect 275 310 276 311 
<< m1 >>
rect 276 310 277 311 
<< m1 >>
rect 277 310 278 311 
<< m1 >>
rect 278 310 279 311 
<< m2 >>
rect 278 310 279 311 
<< m1 >>
rect 279 310 280 311 
<< m1 >>
rect 280 310 281 311 
<< m2 >>
rect 280 310 281 311 
<< m1 >>
rect 281 310 282 311 
<< m1 >>
rect 282 310 283 311 
<< m1 >>
rect 283 310 284 311 
<< m1 >>
rect 284 310 285 311 
<< m1 >>
rect 285 310 286 311 
<< m1 >>
rect 286 310 287 311 
<< m1 >>
rect 287 310 288 311 
<< m1 >>
rect 288 310 289 311 
<< m1 >>
rect 289 310 290 311 
<< m1 >>
rect 290 310 291 311 
<< m1 >>
rect 291 310 292 311 
<< m1 >>
rect 292 310 293 311 
<< m1 >>
rect 293 310 294 311 
<< m1 >>
rect 294 310 295 311 
<< m1 >>
rect 295 310 296 311 
<< m1 >>
rect 296 310 297 311 
<< m1 >>
rect 297 310 298 311 
<< m1 >>
rect 298 310 299 311 
<< m1 >>
rect 299 310 300 311 
<< m1 >>
rect 300 310 301 311 
<< m1 >>
rect 301 310 302 311 
<< m1 >>
rect 302 310 303 311 
<< m2 >>
rect 302 310 303 311 
<< m1 >>
rect 303 310 304 311 
<< m1 >>
rect 304 310 305 311 
<< m1 >>
rect 305 310 306 311 
<< m1 >>
rect 306 310 307 311 
<< m1 >>
rect 307 310 308 311 
<< m2 >>
rect 307 310 308 311 
<< m1 >>
rect 308 310 309 311 
<< m1 >>
rect 309 310 310 311 
<< m1 >>
rect 310 310 311 311 
<< m2 >>
rect 310 310 311 311 
<< m1 >>
rect 311 310 312 311 
<< m1 >>
rect 312 310 313 311 
<< m1 >>
rect 313 310 314 311 
<< m1 >>
rect 314 310 315 311 
<< m1 >>
rect 315 310 316 311 
<< m1 >>
rect 316 310 317 311 
<< m1 >>
rect 317 310 318 311 
<< m1 >>
rect 318 310 319 311 
<< m1 >>
rect 319 310 320 311 
<< m1 >>
rect 320 310 321 311 
<< m1 >>
rect 321 310 322 311 
<< m1 >>
rect 322 310 323 311 
<< m1 >>
rect 323 310 324 311 
<< m1 >>
rect 324 310 325 311 
<< m1 >>
rect 325 310 326 311 
<< m1 >>
rect 326 310 327 311 
<< m1 >>
rect 327 310 328 311 
<< m1 >>
rect 328 310 329 311 
<< m1 >>
rect 329 310 330 311 
<< m1 >>
rect 330 310 331 311 
<< m1 >>
rect 331 310 332 311 
<< m1 >>
rect 332 310 333 311 
<< m2 >>
rect 332 310 333 311 
<< m2c >>
rect 332 310 333 311 
<< m1 >>
rect 332 310 333 311 
<< m2 >>
rect 332 310 333 311 
<< m2 >>
rect 333 310 334 311 
<< m1 >>
rect 334 310 335 311 
<< m2 >>
rect 334 310 335 311 
<< m2 >>
rect 335 310 336 311 
<< m1 >>
rect 336 310 337 311 
<< m2 >>
rect 336 310 337 311 
<< m2c >>
rect 336 310 337 311 
<< m1 >>
rect 336 310 337 311 
<< m2 >>
rect 336 310 337 311 
<< m1 >>
rect 337 310 338 311 
<< m1 >>
rect 338 310 339 311 
<< m1 >>
rect 339 310 340 311 
<< m1 >>
rect 340 310 341 311 
<< m1 >>
rect 341 310 342 311 
<< m1 >>
rect 342 310 343 311 
<< m1 >>
rect 343 310 344 311 
<< m1 >>
rect 344 310 345 311 
<< m2 >>
rect 344 310 345 311 
<< m1 >>
rect 345 310 346 311 
<< m1 >>
rect 346 310 347 311 
<< m2 >>
rect 346 310 347 311 
<< m1 >>
rect 347 310 348 311 
<< m1 >>
rect 348 310 349 311 
<< m2 >>
rect 348 310 349 311 
<< m1 >>
rect 349 310 350 311 
<< m1 >>
rect 350 310 351 311 
<< m2 >>
rect 350 310 351 311 
<< m2c >>
rect 350 310 351 311 
<< m1 >>
rect 350 310 351 311 
<< m2 >>
rect 350 310 351 311 
<< m2 >>
rect 351 310 352 311 
<< m1 >>
rect 352 310 353 311 
<< m2 >>
rect 352 310 353 311 
<< m2 >>
rect 353 310 354 311 
<< m1 >>
rect 354 310 355 311 
<< m2 >>
rect 354 310 355 311 
<< m2c >>
rect 354 310 355 311 
<< m1 >>
rect 354 310 355 311 
<< m2 >>
rect 354 310 355 311 
<< m1 >>
rect 355 310 356 311 
<< m1 >>
rect 356 310 357 311 
<< m1 >>
rect 357 310 358 311 
<< m1 >>
rect 358 310 359 311 
<< m1 >>
rect 359 310 360 311 
<< m1 >>
rect 360 310 361 311 
<< m1 >>
rect 361 310 362 311 
<< m1 >>
rect 362 310 363 311 
<< m1 >>
rect 363 310 364 311 
<< m1 >>
rect 364 310 365 311 
<< m1 >>
rect 365 310 366 311 
<< m1 >>
rect 366 310 367 311 
<< m2 >>
rect 366 310 367 311 
<< m1 >>
rect 367 310 368 311 
<< m1 >>
rect 368 310 369 311 
<< m2 >>
rect 368 310 369 311 
<< m2c >>
rect 368 310 369 311 
<< m1 >>
rect 368 310 369 311 
<< m2 >>
rect 368 310 369 311 
<< m2 >>
rect 369 310 370 311 
<< m1 >>
rect 370 310 371 311 
<< m2 >>
rect 370 310 371 311 
<< m2 >>
rect 371 310 372 311 
<< m1 >>
rect 372 310 373 311 
<< m2 >>
rect 372 310 373 311 
<< m2c >>
rect 372 310 373 311 
<< m1 >>
rect 372 310 373 311 
<< m2 >>
rect 372 310 373 311 
<< m1 >>
rect 373 310 374 311 
<< m1 >>
rect 374 310 375 311 
<< m2 >>
rect 374 310 375 311 
<< m1 >>
rect 375 310 376 311 
<< m1 >>
rect 376 310 377 311 
<< m1 >>
rect 377 310 378 311 
<< m2 >>
rect 377 310 378 311 
<< m2c >>
rect 377 310 378 311 
<< m1 >>
rect 377 310 378 311 
<< m2 >>
rect 377 310 378 311 
<< m2 >>
rect 378 310 379 311 
<< m1 >>
rect 379 310 380 311 
<< m2 >>
rect 379 310 380 311 
<< m2 >>
rect 380 310 381 311 
<< m1 >>
rect 381 310 382 311 
<< m2 >>
rect 381 310 382 311 
<< m2c >>
rect 381 310 382 311 
<< m1 >>
rect 381 310 382 311 
<< m2 >>
rect 381 310 382 311 
<< m1 >>
rect 382 310 383 311 
<< m1 >>
rect 383 310 384 311 
<< m1 >>
rect 384 310 385 311 
<< m1 >>
rect 385 310 386 311 
<< m1 >>
rect 386 310 387 311 
<< m1 >>
rect 387 310 388 311 
<< m1 >>
rect 388 310 389 311 
<< m1 >>
rect 389 310 390 311 
<< m1 >>
rect 390 310 391 311 
<< m2 >>
rect 390 310 391 311 
<< m1 >>
rect 391 310 392 311 
<< m1 >>
rect 392 310 393 311 
<< m1 >>
rect 393 310 394 311 
<< m1 >>
rect 394 310 395 311 
<< m1 >>
rect 395 310 396 311 
<< m1 >>
rect 396 310 397 311 
<< m1 >>
rect 397 310 398 311 
<< m1 >>
rect 398 310 399 311 
<< m1 >>
rect 399 310 400 311 
<< m1 >>
rect 400 310 401 311 
<< m1 >>
rect 401 310 402 311 
<< m1 >>
rect 402 310 403 311 
<< m1 >>
rect 403 310 404 311 
<< m1 >>
rect 404 310 405 311 
<< m2 >>
rect 404 310 405 311 
<< m2c >>
rect 404 310 405 311 
<< m1 >>
rect 404 310 405 311 
<< m2 >>
rect 404 310 405 311 
<< m2 >>
rect 405 310 406 311 
<< m1 >>
rect 406 310 407 311 
<< m2 >>
rect 406 310 407 311 
<< m2 >>
rect 407 310 408 311 
<< m1 >>
rect 408 310 409 311 
<< m2 >>
rect 408 310 409 311 
<< m2c >>
rect 408 310 409 311 
<< m1 >>
rect 408 310 409 311 
<< m2 >>
rect 408 310 409 311 
<< m1 >>
rect 409 310 410 311 
<< m1 >>
rect 410 310 411 311 
<< m1 >>
rect 411 310 412 311 
<< m1 >>
rect 412 310 413 311 
<< m1 >>
rect 413 310 414 311 
<< m1 >>
rect 414 310 415 311 
<< m2 >>
rect 414 310 415 311 
<< m2c >>
rect 414 310 415 311 
<< m1 >>
rect 414 310 415 311 
<< m2 >>
rect 414 310 415 311 
<< m2 >>
rect 415 310 416 311 
<< m1 >>
rect 416 310 417 311 
<< m2 >>
rect 416 310 417 311 
<< m2 >>
rect 417 310 418 311 
<< m1 >>
rect 418 310 419 311 
<< m2 >>
rect 418 310 419 311 
<< m2c >>
rect 418 310 419 311 
<< m1 >>
rect 418 310 419 311 
<< m2 >>
rect 418 310 419 311 
<< m2 >>
rect 419 310 420 311 
<< m1 >>
rect 420 310 421 311 
<< m2 >>
rect 420 310 421 311 
<< m2 >>
rect 421 310 422 311 
<< m1 >>
rect 422 310 423 311 
<< m2 >>
rect 422 310 423 311 
<< m2c >>
rect 422 310 423 311 
<< m1 >>
rect 422 310 423 311 
<< m2 >>
rect 422 310 423 311 
<< m1 >>
rect 423 310 424 311 
<< m1 >>
rect 424 310 425 311 
<< m2 >>
rect 424 310 425 311 
<< m1 >>
rect 425 310 426 311 
<< m1 >>
rect 426 310 427 311 
<< m2 >>
rect 426 310 427 311 
<< m1 >>
rect 427 310 428 311 
<< m2 >>
rect 427 310 428 311 
<< m1 >>
rect 428 310 429 311 
<< m2 >>
rect 428 310 429 311 
<< m1 >>
rect 429 310 430 311 
<< m2 >>
rect 429 310 430 311 
<< m1 >>
rect 430 310 431 311 
<< m1 >>
rect 431 310 432 311 
<< m2 >>
rect 431 310 432 311 
<< m2c >>
rect 431 310 432 311 
<< m1 >>
rect 431 310 432 311 
<< m2 >>
rect 431 310 432 311 
<< m2 >>
rect 432 310 433 311 
<< m1 >>
rect 433 310 434 311 
<< m2 >>
rect 433 310 434 311 
<< m2 >>
rect 434 310 435 311 
<< m1 >>
rect 435 310 436 311 
<< m2 >>
rect 435 310 436 311 
<< m2c >>
rect 435 310 436 311 
<< m1 >>
rect 435 310 436 311 
<< m2 >>
rect 435 310 436 311 
<< m1 >>
rect 437 310 438 311 
<< m1 >>
rect 487 310 488 311 
<< m1 >>
rect 523 310 524 311 
<< m1 >>
rect 19 311 20 312 
<< m1 >>
rect 22 311 23 312 
<< m1 >>
rect 44 311 45 312 
<< m1 >>
rect 46 311 47 312 
<< m2 >>
rect 46 311 47 312 
<< m1 >>
rect 55 311 56 312 
<< m1 >>
rect 73 311 74 312 
<< m2 >>
rect 74 311 75 312 
<< m1 >>
rect 93 311 94 312 
<< m1 >>
rect 100 311 101 312 
<< m1 >>
rect 121 311 122 312 
<< m2 >>
rect 146 311 147 312 
<< m2 >>
rect 148 311 149 312 
<< m2 >>
rect 150 311 151 312 
<< m1 >>
rect 154 311 155 312 
<< m2 >>
rect 180 311 181 312 
<< m2 >>
rect 186 311 187 312 
<< m2 >>
rect 207 311 208 312 
<< m1 >>
rect 208 311 209 312 
<< m1 >>
rect 217 311 218 312 
<< m2 >>
rect 218 311 219 312 
<< m1 >>
rect 229 311 230 312 
<< m2 >>
rect 230 311 231 312 
<< m1 >>
rect 237 311 238 312 
<< m2 >>
rect 243 311 244 312 
<< m1 >>
rect 244 311 245 312 
<< m2 >>
rect 244 311 245 312 
<< m2 >>
rect 245 311 246 312 
<< m2 >>
rect 246 311 247 312 
<< m2 >>
rect 247 311 248 312 
<< m2 >>
rect 248 311 249 312 
<< m2 >>
rect 249 311 250 312 
<< m1 >>
rect 253 311 254 312 
<< m2 >>
rect 257 311 258 312 
<< m2 >>
rect 258 311 259 312 
<< m2 >>
rect 259 311 260 312 
<< m2 >>
rect 260 311 261 312 
<< m2 >>
rect 261 311 262 312 
<< m2 >>
rect 262 311 263 312 
<< m2 >>
rect 263 311 264 312 
<< m2 >>
rect 264 311 265 312 
<< m2 >>
rect 265 311 266 312 
<< m2 >>
rect 266 311 267 312 
<< m1 >>
rect 271 311 272 312 
<< m2 >>
rect 278 311 279 312 
<< m2 >>
rect 280 311 281 312 
<< m2 >>
rect 282 311 283 312 
<< m2 >>
rect 283 311 284 312 
<< m2 >>
rect 284 311 285 312 
<< m2 >>
rect 285 311 286 312 
<< m2 >>
rect 286 311 287 312 
<< m2 >>
rect 287 311 288 312 
<< m2 >>
rect 288 311 289 312 
<< m2 >>
rect 289 311 290 312 
<< m2 >>
rect 290 311 291 312 
<< m2 >>
rect 291 311 292 312 
<< m2 >>
rect 292 311 293 312 
<< m2 >>
rect 293 311 294 312 
<< m2 >>
rect 294 311 295 312 
<< m2 >>
rect 295 311 296 312 
<< m2 >>
rect 296 311 297 312 
<< m2 >>
rect 297 311 298 312 
<< m2 >>
rect 298 311 299 312 
<< m2 >>
rect 299 311 300 312 
<< m2 >>
rect 300 311 301 312 
<< m2 >>
rect 301 311 302 312 
<< m2 >>
rect 302 311 303 312 
<< m2 >>
rect 307 311 308 312 
<< m2 >>
rect 310 311 311 312 
<< m2 >>
rect 311 311 312 312 
<< m2 >>
rect 312 311 313 312 
<< m2 >>
rect 313 311 314 312 
<< m2 >>
rect 314 311 315 312 
<< m2 >>
rect 315 311 316 312 
<< m2 >>
rect 316 311 317 312 
<< m2 >>
rect 317 311 318 312 
<< m2 >>
rect 318 311 319 312 
<< m2 >>
rect 319 311 320 312 
<< m2 >>
rect 320 311 321 312 
<< m2 >>
rect 321 311 322 312 
<< m2 >>
rect 322 311 323 312 
<< m2 >>
rect 323 311 324 312 
<< m2 >>
rect 324 311 325 312 
<< m2 >>
rect 325 311 326 312 
<< m2 >>
rect 326 311 327 312 
<< m2 >>
rect 327 311 328 312 
<< m2 >>
rect 328 311 329 312 
<< m2 >>
rect 329 311 330 312 
<< m2 >>
rect 330 311 331 312 
<< m1 >>
rect 334 311 335 312 
<< m2 >>
rect 344 311 345 312 
<< m2 >>
rect 346 311 347 312 
<< m2 >>
rect 348 311 349 312 
<< m1 >>
rect 352 311 353 312 
<< m2 >>
rect 366 311 367 312 
<< m1 >>
rect 370 311 371 312 
<< m2 >>
rect 374 311 375 312 
<< m1 >>
rect 379 311 380 312 
<< m2 >>
rect 390 311 391 312 
<< m2 >>
rect 391 311 392 312 
<< m2 >>
rect 392 311 393 312 
<< m2 >>
rect 393 311 394 312 
<< m2 >>
rect 394 311 395 312 
<< m2 >>
rect 395 311 396 312 
<< m2 >>
rect 396 311 397 312 
<< m2 >>
rect 397 311 398 312 
<< m2 >>
rect 398 311 399 312 
<< m2 >>
rect 399 311 400 312 
<< m2 >>
rect 400 311 401 312 
<< m2 >>
rect 401 311 402 312 
<< m2 >>
rect 402 311 403 312 
<< m1 >>
rect 406 311 407 312 
<< m1 >>
rect 416 311 417 312 
<< m1 >>
rect 420 311 421 312 
<< m2 >>
rect 424 311 425 312 
<< m2 >>
rect 426 311 427 312 
<< m1 >>
rect 433 311 434 312 
<< m1 >>
rect 435 311 436 312 
<< m1 >>
rect 437 311 438 312 
<< m1 >>
rect 487 311 488 312 
<< m1 >>
rect 523 311 524 312 
<< m1 >>
rect 19 312 20 313 
<< m1 >>
rect 22 312 23 313 
<< m1 >>
rect 44 312 45 313 
<< m1 >>
rect 46 312 47 313 
<< m2 >>
rect 46 312 47 313 
<< m1 >>
rect 55 312 56 313 
<< m1 >>
rect 73 312 74 313 
<< m2 >>
rect 74 312 75 313 
<< m1 >>
rect 93 312 94 313 
<< m1 >>
rect 100 312 101 313 
<< m1 >>
rect 121 312 122 313 
<< m1 >>
rect 136 312 137 313 
<< m1 >>
rect 137 312 138 313 
<< m1 >>
rect 138 312 139 313 
<< m1 >>
rect 139 312 140 313 
<< m1 >>
rect 140 312 141 313 
<< m1 >>
rect 141 312 142 313 
<< m1 >>
rect 142 312 143 313 
<< m1 >>
rect 143 312 144 313 
<< m1 >>
rect 144 312 145 313 
<< m1 >>
rect 145 312 146 313 
<< m1 >>
rect 146 312 147 313 
<< m2 >>
rect 146 312 147 313 
<< m2c >>
rect 146 312 147 313 
<< m1 >>
rect 146 312 147 313 
<< m2 >>
rect 146 312 147 313 
<< m1 >>
rect 148 312 149 313 
<< m2 >>
rect 148 312 149 313 
<< m2c >>
rect 148 312 149 313 
<< m1 >>
rect 148 312 149 313 
<< m2 >>
rect 148 312 149 313 
<< m1 >>
rect 150 312 151 313 
<< m2 >>
rect 150 312 151 313 
<< m2c >>
rect 150 312 151 313 
<< m1 >>
rect 150 312 151 313 
<< m2 >>
rect 150 312 151 313 
<< m1 >>
rect 154 312 155 313 
<< m1 >>
rect 180 312 181 313 
<< m2 >>
rect 180 312 181 313 
<< m2c >>
rect 180 312 181 313 
<< m1 >>
rect 180 312 181 313 
<< m2 >>
rect 180 312 181 313 
<< m1 >>
rect 186 312 187 313 
<< m2 >>
rect 186 312 187 313 
<< m2c >>
rect 186 312 187 313 
<< m1 >>
rect 186 312 187 313 
<< m2 >>
rect 186 312 187 313 
<< m2 >>
rect 207 312 208 313 
<< m1 >>
rect 208 312 209 313 
<< m1 >>
rect 217 312 218 313 
<< m2 >>
rect 218 312 219 313 
<< m1 >>
rect 229 312 230 313 
<< m2 >>
rect 230 312 231 313 
<< m1 >>
rect 237 312 238 313 
<< m2 >>
rect 243 312 244 313 
<< m1 >>
rect 244 312 245 313 
<< m1 >>
rect 253 312 254 313 
<< m1 >>
rect 257 312 258 313 
<< m2 >>
rect 257 312 258 313 
<< m2c >>
rect 257 312 258 313 
<< m1 >>
rect 257 312 258 313 
<< m2 >>
rect 257 312 258 313 
<< m1 >>
rect 271 312 272 313 
<< m1 >>
rect 276 312 277 313 
<< m1 >>
rect 277 312 278 313 
<< m1 >>
rect 278 312 279 313 
<< m2 >>
rect 278 312 279 313 
<< m2c >>
rect 278 312 279 313 
<< m1 >>
rect 278 312 279 313 
<< m2 >>
rect 278 312 279 313 
<< m1 >>
rect 280 312 281 313 
<< m2 >>
rect 280 312 281 313 
<< m2c >>
rect 280 312 281 313 
<< m1 >>
rect 280 312 281 313 
<< m2 >>
rect 280 312 281 313 
<< m1 >>
rect 282 312 283 313 
<< m2 >>
rect 282 312 283 313 
<< m2c >>
rect 282 312 283 313 
<< m1 >>
rect 282 312 283 313 
<< m2 >>
rect 282 312 283 313 
<< m1 >>
rect 307 312 308 313 
<< m2 >>
rect 307 312 308 313 
<< m2c >>
rect 307 312 308 313 
<< m1 >>
rect 307 312 308 313 
<< m2 >>
rect 307 312 308 313 
<< m1 >>
rect 330 312 331 313 
<< m2 >>
rect 330 312 331 313 
<< m2c >>
rect 330 312 331 313 
<< m1 >>
rect 330 312 331 313 
<< m2 >>
rect 330 312 331 313 
<< m1 >>
rect 334 312 335 313 
<< m2 >>
rect 344 312 345 313 
<< m2 >>
rect 346 312 347 313 
<< m2 >>
rect 348 312 349 313 
<< m1 >>
rect 352 312 353 313 
<< m1 >>
rect 366 312 367 313 
<< m2 >>
rect 366 312 367 313 
<< m2c >>
rect 366 312 367 313 
<< m1 >>
rect 366 312 367 313 
<< m2 >>
rect 366 312 367 313 
<< m1 >>
rect 370 312 371 313 
<< m1 >>
rect 374 312 375 313 
<< m2 >>
rect 374 312 375 313 
<< m2c >>
rect 374 312 375 313 
<< m1 >>
rect 374 312 375 313 
<< m2 >>
rect 374 312 375 313 
<< m1 >>
rect 379 312 380 313 
<< m1 >>
rect 402 312 403 313 
<< m2 >>
rect 402 312 403 313 
<< m2c >>
rect 402 312 403 313 
<< m1 >>
rect 402 312 403 313 
<< m2 >>
rect 402 312 403 313 
<< m1 >>
rect 406 312 407 313 
<< m1 >>
rect 416 312 417 313 
<< m1 >>
rect 420 312 421 313 
<< m1 >>
rect 424 312 425 313 
<< m2 >>
rect 424 312 425 313 
<< m2c >>
rect 424 312 425 313 
<< m1 >>
rect 424 312 425 313 
<< m2 >>
rect 424 312 425 313 
<< m1 >>
rect 425 312 426 313 
<< m1 >>
rect 426 312 427 313 
<< m2 >>
rect 426 312 427 313 
<< m1 >>
rect 427 312 428 313 
<< m1 >>
rect 428 312 429 313 
<< m1 >>
rect 429 312 430 313 
<< m1 >>
rect 430 312 431 313 
<< m1 >>
rect 431 312 432 313 
<< m2 >>
rect 431 312 432 313 
<< m2c >>
rect 431 312 432 313 
<< m1 >>
rect 431 312 432 313 
<< m2 >>
rect 431 312 432 313 
<< m2 >>
rect 432 312 433 313 
<< m1 >>
rect 433 312 434 313 
<< m2 >>
rect 433 312 434 313 
<< m2 >>
rect 434 312 435 313 
<< m1 >>
rect 435 312 436 313 
<< m2 >>
rect 435 312 436 313 
<< m2 >>
rect 436 312 437 313 
<< m1 >>
rect 437 312 438 313 
<< m2 >>
rect 437 312 438 313 
<< m2 >>
rect 438 312 439 313 
<< m1 >>
rect 439 312 440 313 
<< m2 >>
rect 439 312 440 313 
<< m2c >>
rect 439 312 440 313 
<< m1 >>
rect 439 312 440 313 
<< m2 >>
rect 439 312 440 313 
<< m1 >>
rect 487 312 488 313 
<< m1 >>
rect 523 312 524 313 
<< m1 >>
rect 19 313 20 314 
<< m1 >>
rect 22 313 23 314 
<< m1 >>
rect 44 313 45 314 
<< m1 >>
rect 46 313 47 314 
<< m2 >>
rect 46 313 47 314 
<< m1 >>
rect 55 313 56 314 
<< m1 >>
rect 73 313 74 314 
<< m2 >>
rect 74 313 75 314 
<< m1 >>
rect 93 313 94 314 
<< m1 >>
rect 100 313 101 314 
<< m1 >>
rect 121 313 122 314 
<< m1 >>
rect 136 313 137 314 
<< m1 >>
rect 148 313 149 314 
<< m1 >>
rect 150 313 151 314 
<< m1 >>
rect 152 313 153 314 
<< m2 >>
rect 152 313 153 314 
<< m2c >>
rect 152 313 153 314 
<< m1 >>
rect 152 313 153 314 
<< m2 >>
rect 152 313 153 314 
<< m2 >>
rect 153 313 154 314 
<< m1 >>
rect 154 313 155 314 
<< m2 >>
rect 154 313 155 314 
<< m2 >>
rect 155 313 156 314 
<< m1 >>
rect 156 313 157 314 
<< m2 >>
rect 156 313 157 314 
<< m1 >>
rect 157 313 158 314 
<< m2 >>
rect 157 313 158 314 
<< m2c >>
rect 157 313 158 314 
<< m1 >>
rect 157 313 158 314 
<< m2 >>
rect 157 313 158 314 
<< m2 >>
rect 158 313 159 314 
<< m1 >>
rect 159 313 160 314 
<< m2 >>
rect 159 313 160 314 
<< m1 >>
rect 160 313 161 314 
<< m2 >>
rect 160 313 161 314 
<< m1 >>
rect 161 313 162 314 
<< m2 >>
rect 161 313 162 314 
<< m1 >>
rect 162 313 163 314 
<< m2 >>
rect 162 313 163 314 
<< m1 >>
rect 163 313 164 314 
<< m2 >>
rect 163 313 164 314 
<< m1 >>
rect 164 313 165 314 
<< m2 >>
rect 164 313 165 314 
<< m1 >>
rect 165 313 166 314 
<< m2 >>
rect 165 313 166 314 
<< m1 >>
rect 166 313 167 314 
<< m2 >>
rect 166 313 167 314 
<< m1 >>
rect 167 313 168 314 
<< m2 >>
rect 167 313 168 314 
<< m1 >>
rect 168 313 169 314 
<< m2 >>
rect 168 313 169 314 
<< m1 >>
rect 169 313 170 314 
<< m2 >>
rect 169 313 170 314 
<< m1 >>
rect 170 313 171 314 
<< m2 >>
rect 170 313 171 314 
<< m1 >>
rect 171 313 172 314 
<< m2 >>
rect 171 313 172 314 
<< m1 >>
rect 172 313 173 314 
<< m2 >>
rect 172 313 173 314 
<< m1 >>
rect 173 313 174 314 
<< m2 >>
rect 173 313 174 314 
<< m1 >>
rect 174 313 175 314 
<< m2 >>
rect 174 313 175 314 
<< m1 >>
rect 175 313 176 314 
<< m2 >>
rect 175 313 176 314 
<< m1 >>
rect 176 313 177 314 
<< m2 >>
rect 176 313 177 314 
<< m1 >>
rect 177 313 178 314 
<< m2 >>
rect 177 313 178 314 
<< m1 >>
rect 178 313 179 314 
<< m2 >>
rect 178 313 179 314 
<< m1 >>
rect 179 313 180 314 
<< m1 >>
rect 180 313 181 314 
<< m1 >>
rect 186 313 187 314 
<< m2 >>
rect 207 313 208 314 
<< m1 >>
rect 208 313 209 314 
<< m1 >>
rect 217 313 218 314 
<< m2 >>
rect 218 313 219 314 
<< m1 >>
rect 223 313 224 314 
<< m1 >>
rect 224 313 225 314 
<< m1 >>
rect 225 313 226 314 
<< m2 >>
rect 225 313 226 314 
<< m1 >>
rect 226 313 227 314 
<< m2 >>
rect 226 313 227 314 
<< m1 >>
rect 227 313 228 314 
<< m2 >>
rect 227 313 228 314 
<< m1 >>
rect 228 313 229 314 
<< m2 >>
rect 228 313 229 314 
<< m1 >>
rect 229 313 230 314 
<< m2 >>
rect 229 313 230 314 
<< m2 >>
rect 230 313 231 314 
<< m1 >>
rect 237 313 238 314 
<< m2 >>
rect 243 313 244 314 
<< m1 >>
rect 244 313 245 314 
<< m1 >>
rect 253 313 254 314 
<< m1 >>
rect 257 313 258 314 
<< m1 >>
rect 271 313 272 314 
<< m1 >>
rect 276 313 277 314 
<< m1 >>
rect 280 313 281 314 
<< m1 >>
rect 282 313 283 314 
<< m1 >>
rect 307 313 308 314 
<< m1 >>
rect 330 313 331 314 
<< m1 >>
rect 331 313 332 314 
<< m1 >>
rect 332 313 333 314 
<< m2 >>
rect 332 313 333 314 
<< m2c >>
rect 332 313 333 314 
<< m1 >>
rect 332 313 333 314 
<< m2 >>
rect 332 313 333 314 
<< m2 >>
rect 333 313 334 314 
<< m1 >>
rect 334 313 335 314 
<< m2 >>
rect 334 313 335 314 
<< m2 >>
rect 335 313 336 314 
<< m1 >>
rect 336 313 337 314 
<< m2 >>
rect 336 313 337 314 
<< m2c >>
rect 336 313 337 314 
<< m1 >>
rect 336 313 337 314 
<< m2 >>
rect 336 313 337 314 
<< m1 >>
rect 337 313 338 314 
<< m1 >>
rect 338 313 339 314 
<< m1 >>
rect 339 313 340 314 
<< m1 >>
rect 340 313 341 314 
<< m1 >>
rect 341 313 342 314 
<< m1 >>
rect 342 313 343 314 
<< m1 >>
rect 343 313 344 314 
<< m1 >>
rect 344 313 345 314 
<< m2 >>
rect 344 313 345 314 
<< m1 >>
rect 345 313 346 314 
<< m1 >>
rect 346 313 347 314 
<< m2 >>
rect 346 313 347 314 
<< m1 >>
rect 347 313 348 314 
<< m1 >>
rect 348 313 349 314 
<< m2 >>
rect 348 313 349 314 
<< m1 >>
rect 349 313 350 314 
<< m1 >>
rect 350 313 351 314 
<< m1 >>
rect 352 313 353 314 
<< m1 >>
rect 366 313 367 314 
<< m1 >>
rect 370 313 371 314 
<< m1 >>
rect 372 313 373 314 
<< m1 >>
rect 373 313 374 314 
<< m1 >>
rect 374 313 375 314 
<< m1 >>
rect 379 313 380 314 
<< m1 >>
rect 402 313 403 314 
<< m1 >>
rect 403 313 404 314 
<< m1 >>
rect 404 313 405 314 
<< m2 >>
rect 404 313 405 314 
<< m2c >>
rect 404 313 405 314 
<< m1 >>
rect 404 313 405 314 
<< m2 >>
rect 404 313 405 314 
<< m2 >>
rect 405 313 406 314 
<< m1 >>
rect 406 313 407 314 
<< m2 >>
rect 406 313 407 314 
<< m1 >>
rect 407 313 408 314 
<< m2 >>
rect 407 313 408 314 
<< m1 >>
rect 408 313 409 314 
<< m2 >>
rect 408 313 409 314 
<< m1 >>
rect 409 313 410 314 
<< m2 >>
rect 409 313 410 314 
<< m1 >>
rect 410 313 411 314 
<< m2 >>
rect 410 313 411 314 
<< m1 >>
rect 411 313 412 314 
<< m2 >>
rect 411 313 412 314 
<< m1 >>
rect 412 313 413 314 
<< m2 >>
rect 412 313 413 314 
<< m1 >>
rect 413 313 414 314 
<< m2 >>
rect 413 313 414 314 
<< m1 >>
rect 414 313 415 314 
<< m2 >>
rect 414 313 415 314 
<< m2 >>
rect 415 313 416 314 
<< m1 >>
rect 416 313 417 314 
<< m2 >>
rect 416 313 417 314 
<< m2 >>
rect 417 313 418 314 
<< m1 >>
rect 420 313 421 314 
<< m2 >>
rect 426 313 427 314 
<< m1 >>
rect 433 313 434 314 
<< m1 >>
rect 435 313 436 314 
<< m1 >>
rect 437 313 438 314 
<< m1 >>
rect 439 313 440 314 
<< m1 >>
rect 487 313 488 314 
<< m1 >>
rect 523 313 524 314 
<< m1 >>
rect 19 314 20 315 
<< m1 >>
rect 22 314 23 315 
<< m2 >>
rect 22 314 23 315 
<< m2c >>
rect 22 314 23 315 
<< m1 >>
rect 22 314 23 315 
<< m2 >>
rect 22 314 23 315 
<< m1 >>
rect 44 314 45 315 
<< m1 >>
rect 46 314 47 315 
<< m2 >>
rect 46 314 47 315 
<< m1 >>
rect 55 314 56 315 
<< m1 >>
rect 73 314 74 315 
<< m2 >>
rect 74 314 75 315 
<< m1 >>
rect 93 314 94 315 
<< m1 >>
rect 100 314 101 315 
<< m1 >>
rect 121 314 122 315 
<< m1 >>
rect 136 314 137 315 
<< m1 >>
rect 148 314 149 315 
<< m1 >>
rect 150 314 151 315 
<< m2 >>
rect 151 314 152 315 
<< m1 >>
rect 152 314 153 315 
<< m2 >>
rect 152 314 153 315 
<< m1 >>
rect 154 314 155 315 
<< m1 >>
rect 159 314 160 315 
<< m2 >>
rect 178 314 179 315 
<< m2 >>
rect 179 314 180 315 
<< m2 >>
rect 180 314 181 315 
<< m2 >>
rect 181 314 182 315 
<< m1 >>
rect 182 314 183 315 
<< m2 >>
rect 182 314 183 315 
<< m2c >>
rect 182 314 183 315 
<< m1 >>
rect 182 314 183 315 
<< m2 >>
rect 182 314 183 315 
<< m1 >>
rect 183 314 184 315 
<< m1 >>
rect 184 314 185 315 
<< m1 >>
rect 185 314 186 315 
<< m1 >>
rect 186 314 187 315 
<< m2 >>
rect 207 314 208 315 
<< m1 >>
rect 208 314 209 315 
<< m1 >>
rect 217 314 218 315 
<< m2 >>
rect 218 314 219 315 
<< m1 >>
rect 223 314 224 315 
<< m2 >>
rect 225 314 226 315 
<< m1 >>
rect 237 314 238 315 
<< m2 >>
rect 243 314 244 315 
<< m1 >>
rect 244 314 245 315 
<< m1 >>
rect 253 314 254 315 
<< m1 >>
rect 257 314 258 315 
<< m1 >>
rect 271 314 272 315 
<< m1 >>
rect 276 314 277 315 
<< m1 >>
rect 280 314 281 315 
<< m1 >>
rect 282 314 283 315 
<< m1 >>
rect 307 314 308 315 
<< m1 >>
rect 334 314 335 315 
<< m2 >>
rect 344 314 345 315 
<< m2 >>
rect 346 314 347 315 
<< m2 >>
rect 348 314 349 315 
<< m1 >>
rect 350 314 351 315 
<< m1 >>
rect 352 314 353 315 
<< m1 >>
rect 366 314 367 315 
<< m1 >>
rect 370 314 371 315 
<< m1 >>
rect 372 314 373 315 
<< m1 >>
rect 379 314 380 315 
<< m1 >>
rect 414 314 415 315 
<< m1 >>
rect 416 314 417 315 
<< m2 >>
rect 417 314 418 315 
<< m1 >>
rect 418 314 419 315 
<< m2 >>
rect 418 314 419 315 
<< m2c >>
rect 418 314 419 315 
<< m1 >>
rect 418 314 419 315 
<< m2 >>
rect 418 314 419 315 
<< m2 >>
rect 419 314 420 315 
<< m1 >>
rect 420 314 421 315 
<< m2 >>
rect 420 314 421 315 
<< m2 >>
rect 421 314 422 315 
<< m1 >>
rect 422 314 423 315 
<< m2 >>
rect 422 314 423 315 
<< m2c >>
rect 422 314 423 315 
<< m1 >>
rect 422 314 423 315 
<< m2 >>
rect 422 314 423 315 
<< m1 >>
rect 423 314 424 315 
<< m1 >>
rect 424 314 425 315 
<< m1 >>
rect 425 314 426 315 
<< m1 >>
rect 426 314 427 315 
<< m2 >>
rect 426 314 427 315 
<< m2c >>
rect 426 314 427 315 
<< m1 >>
rect 426 314 427 315 
<< m2 >>
rect 426 314 427 315 
<< m1 >>
rect 433 314 434 315 
<< m1 >>
rect 435 314 436 315 
<< m1 >>
rect 437 314 438 315 
<< m1 >>
rect 439 314 440 315 
<< m1 >>
rect 487 314 488 315 
<< m1 >>
rect 523 314 524 315 
<< m1 >>
rect 19 315 20 316 
<< m2 >>
rect 22 315 23 316 
<< m1 >>
rect 44 315 45 316 
<< m1 >>
rect 46 315 47 316 
<< m2 >>
rect 46 315 47 316 
<< m1 >>
rect 55 315 56 316 
<< m1 >>
rect 73 315 74 316 
<< m2 >>
rect 74 315 75 316 
<< m1 >>
rect 93 315 94 316 
<< m1 >>
rect 100 315 101 316 
<< m1 >>
rect 121 315 122 316 
<< m1 >>
rect 136 315 137 316 
<< m1 >>
rect 148 315 149 316 
<< m1 >>
rect 150 315 151 316 
<< m2 >>
rect 151 315 152 316 
<< m1 >>
rect 154 315 155 316 
<< m1 >>
rect 159 315 160 316 
<< m2 >>
rect 207 315 208 316 
<< m1 >>
rect 208 315 209 316 
<< m1 >>
rect 217 315 218 316 
<< m2 >>
rect 218 315 219 316 
<< m1 >>
rect 223 315 224 316 
<< m1 >>
rect 225 315 226 316 
<< m2 >>
rect 225 315 226 316 
<< m2c >>
rect 225 315 226 316 
<< m1 >>
rect 225 315 226 316 
<< m2 >>
rect 225 315 226 316 
<< m1 >>
rect 237 315 238 316 
<< m2 >>
rect 243 315 244 316 
<< m1 >>
rect 244 315 245 316 
<< m1 >>
rect 253 315 254 316 
<< m1 >>
rect 257 315 258 316 
<< m1 >>
rect 271 315 272 316 
<< m1 >>
rect 276 315 277 316 
<< m1 >>
rect 280 315 281 316 
<< m1 >>
rect 282 315 283 316 
<< m1 >>
rect 307 315 308 316 
<< m1 >>
rect 334 315 335 316 
<< m1 >>
rect 344 315 345 316 
<< m2 >>
rect 344 315 345 316 
<< m2c >>
rect 344 315 345 316 
<< m1 >>
rect 344 315 345 316 
<< m2 >>
rect 344 315 345 316 
<< m2 >>
rect 346 315 347 316 
<< m1 >>
rect 347 315 348 316 
<< m1 >>
rect 348 315 349 316 
<< m2 >>
rect 348 315 349 316 
<< m2c >>
rect 348 315 349 316 
<< m1 >>
rect 348 315 349 316 
<< m2 >>
rect 348 315 349 316 
<< m1 >>
rect 350 315 351 316 
<< m1 >>
rect 352 315 353 316 
<< m1 >>
rect 366 315 367 316 
<< m1 >>
rect 370 315 371 316 
<< m1 >>
rect 372 315 373 316 
<< m1 >>
rect 379 315 380 316 
<< m1 >>
rect 414 315 415 316 
<< m1 >>
rect 416 315 417 316 
<< m1 >>
rect 420 315 421 316 
<< m1 >>
rect 433 315 434 316 
<< m1 >>
rect 435 315 436 316 
<< m1 >>
rect 437 315 438 316 
<< m1 >>
rect 439 315 440 316 
<< m1 >>
rect 487 315 488 316 
<< m1 >>
rect 523 315 524 316 
<< m1 >>
rect 19 316 20 317 
<< m2 >>
rect 22 316 23 317 
<< m1 >>
rect 23 316 24 317 
<< m1 >>
rect 24 316 25 317 
<< m1 >>
rect 25 316 26 317 
<< m1 >>
rect 26 316 27 317 
<< m1 >>
rect 27 316 28 317 
<< m1 >>
rect 28 316 29 317 
<< m1 >>
rect 29 316 30 317 
<< m1 >>
rect 30 316 31 317 
<< m1 >>
rect 31 316 32 317 
<< m1 >>
rect 44 316 45 317 
<< m1 >>
rect 46 316 47 317 
<< m2 >>
rect 46 316 47 317 
<< m1 >>
rect 55 316 56 317 
<< m1 >>
rect 73 316 74 317 
<< m2 >>
rect 74 316 75 317 
<< m1 >>
rect 93 316 94 317 
<< m1 >>
rect 100 316 101 317 
<< m1 >>
rect 121 316 122 317 
<< m1 >>
rect 136 316 137 317 
<< m1 >>
rect 148 316 149 317 
<< m1 >>
rect 150 316 151 317 
<< m2 >>
rect 151 316 152 317 
<< m1 >>
rect 154 316 155 317 
<< m1 >>
rect 159 316 160 317 
<< m2 >>
rect 207 316 208 317 
<< m1 >>
rect 208 316 209 317 
<< m1 >>
rect 217 316 218 317 
<< m2 >>
rect 218 316 219 317 
<< m1 >>
rect 223 316 224 317 
<< m1 >>
rect 225 316 226 317 
<< m1 >>
rect 237 316 238 317 
<< m2 >>
rect 243 316 244 317 
<< m1 >>
rect 244 316 245 317 
<< m1 >>
rect 253 316 254 317 
<< m1 >>
rect 257 316 258 317 
<< m1 >>
rect 271 316 272 317 
<< m1 >>
rect 276 316 277 317 
<< m2 >>
rect 279 316 280 317 
<< m1 >>
rect 280 316 281 317 
<< m2 >>
rect 280 316 281 317 
<< m2 >>
rect 281 316 282 317 
<< m1 >>
rect 282 316 283 317 
<< m2 >>
rect 282 316 283 317 
<< m2c >>
rect 282 316 283 317 
<< m1 >>
rect 282 316 283 317 
<< m2 >>
rect 282 316 283 317 
<< m1 >>
rect 307 316 308 317 
<< m1 >>
rect 334 316 335 317 
<< m1 >>
rect 344 316 345 317 
<< m2 >>
rect 346 316 347 317 
<< m1 >>
rect 347 316 348 317 
<< m1 >>
rect 350 316 351 317 
<< m1 >>
rect 352 316 353 317 
<< m1 >>
rect 366 316 367 317 
<< m2 >>
rect 369 316 370 317 
<< m1 >>
rect 370 316 371 317 
<< m2 >>
rect 370 316 371 317 
<< m2 >>
rect 371 316 372 317 
<< m1 >>
rect 372 316 373 317 
<< m2 >>
rect 372 316 373 317 
<< m2c >>
rect 372 316 373 317 
<< m1 >>
rect 372 316 373 317 
<< m2 >>
rect 372 316 373 317 
<< m1 >>
rect 379 316 380 317 
<< m1 >>
rect 414 316 415 317 
<< m2 >>
rect 414 316 415 317 
<< m2c >>
rect 414 316 415 317 
<< m1 >>
rect 414 316 415 317 
<< m2 >>
rect 414 316 415 317 
<< m2 >>
rect 415 316 416 317 
<< m1 >>
rect 416 316 417 317 
<< m2 >>
rect 416 316 417 317 
<< m2 >>
rect 417 316 418 317 
<< m1 >>
rect 420 316 421 317 
<< m1 >>
rect 424 316 425 317 
<< m1 >>
rect 425 316 426 317 
<< m1 >>
rect 426 316 427 317 
<< m1 >>
rect 427 316 428 317 
<< m1 >>
rect 433 316 434 317 
<< m1 >>
rect 435 316 436 317 
<< m1 >>
rect 437 316 438 317 
<< m1 >>
rect 439 316 440 317 
<< m1 >>
rect 487 316 488 317 
<< m1 >>
rect 523 316 524 317 
<< m1 >>
rect 19 317 20 318 
<< m2 >>
rect 22 317 23 318 
<< m1 >>
rect 23 317 24 318 
<< m1 >>
rect 31 317 32 318 
<< m1 >>
rect 44 317 45 318 
<< m1 >>
rect 46 317 47 318 
<< m2 >>
rect 46 317 47 318 
<< m1 >>
rect 55 317 56 318 
<< m1 >>
rect 73 317 74 318 
<< m2 >>
rect 74 317 75 318 
<< m1 >>
rect 93 317 94 318 
<< m1 >>
rect 100 317 101 318 
<< m1 >>
rect 121 317 122 318 
<< m1 >>
rect 136 317 137 318 
<< m1 >>
rect 148 317 149 318 
<< m1 >>
rect 150 317 151 318 
<< m2 >>
rect 151 317 152 318 
<< m1 >>
rect 154 317 155 318 
<< m1 >>
rect 159 317 160 318 
<< m2 >>
rect 207 317 208 318 
<< m1 >>
rect 208 317 209 318 
<< m1 >>
rect 217 317 218 318 
<< m2 >>
rect 218 317 219 318 
<< m1 >>
rect 223 317 224 318 
<< m1 >>
rect 225 317 226 318 
<< m1 >>
rect 237 317 238 318 
<< m2 >>
rect 243 317 244 318 
<< m1 >>
rect 244 317 245 318 
<< m1 >>
rect 253 317 254 318 
<< m1 >>
rect 257 317 258 318 
<< m1 >>
rect 271 317 272 318 
<< m1 >>
rect 276 317 277 318 
<< m2 >>
rect 279 317 280 318 
<< m1 >>
rect 280 317 281 318 
<< m1 >>
rect 307 317 308 318 
<< m1 >>
rect 334 317 335 318 
<< m1 >>
rect 344 317 345 318 
<< m2 >>
rect 346 317 347 318 
<< m1 >>
rect 347 317 348 318 
<< m1 >>
rect 350 317 351 318 
<< m1 >>
rect 352 317 353 318 
<< m1 >>
rect 366 317 367 318 
<< m2 >>
rect 369 317 370 318 
<< m1 >>
rect 370 317 371 318 
<< m1 >>
rect 379 317 380 318 
<< m1 >>
rect 416 317 417 318 
<< m2 >>
rect 417 317 418 318 
<< m1 >>
rect 420 317 421 318 
<< m1 >>
rect 424 317 425 318 
<< m1 >>
rect 427 317 428 318 
<< m1 >>
rect 433 317 434 318 
<< m1 >>
rect 435 317 436 318 
<< m1 >>
rect 437 317 438 318 
<< m1 >>
rect 439 317 440 318 
<< m1 >>
rect 487 317 488 318 
<< m1 >>
rect 523 317 524 318 
<< pdiffusion >>
rect 12 318 13 319 
<< pdiffusion >>
rect 13 318 14 319 
<< pdiffusion >>
rect 14 318 15 319 
<< pdiffusion >>
rect 15 318 16 319 
<< pdiffusion >>
rect 16 318 17 319 
<< pdiffusion >>
rect 17 318 18 319 
<< m1 >>
rect 19 318 20 319 
<< m2 >>
rect 22 318 23 319 
<< m1 >>
rect 23 318 24 319 
<< m2 >>
rect 23 318 24 319 
<< m2 >>
rect 24 318 25 319 
<< m1 >>
rect 25 318 26 319 
<< m2 >>
rect 25 318 26 319 
<< m2c >>
rect 25 318 26 319 
<< m1 >>
rect 25 318 26 319 
<< m2 >>
rect 25 318 26 319 
<< pdiffusion >>
rect 30 318 31 319 
<< m1 >>
rect 31 318 32 319 
<< pdiffusion >>
rect 31 318 32 319 
<< pdiffusion >>
rect 32 318 33 319 
<< pdiffusion >>
rect 33 318 34 319 
<< pdiffusion >>
rect 34 318 35 319 
<< pdiffusion >>
rect 35 318 36 319 
<< m1 >>
rect 44 318 45 319 
<< m1 >>
rect 46 318 47 319 
<< m2 >>
rect 46 318 47 319 
<< pdiffusion >>
rect 48 318 49 319 
<< pdiffusion >>
rect 49 318 50 319 
<< pdiffusion >>
rect 50 318 51 319 
<< pdiffusion >>
rect 51 318 52 319 
<< pdiffusion >>
rect 52 318 53 319 
<< pdiffusion >>
rect 53 318 54 319 
<< m1 >>
rect 55 318 56 319 
<< pdiffusion >>
rect 66 318 67 319 
<< pdiffusion >>
rect 67 318 68 319 
<< pdiffusion >>
rect 68 318 69 319 
<< pdiffusion >>
rect 69 318 70 319 
<< pdiffusion >>
rect 70 318 71 319 
<< pdiffusion >>
rect 71 318 72 319 
<< m1 >>
rect 73 318 74 319 
<< m2 >>
rect 74 318 75 319 
<< pdiffusion >>
rect 84 318 85 319 
<< pdiffusion >>
rect 85 318 86 319 
<< pdiffusion >>
rect 86 318 87 319 
<< pdiffusion >>
rect 87 318 88 319 
<< pdiffusion >>
rect 88 318 89 319 
<< pdiffusion >>
rect 89 318 90 319 
<< m1 >>
rect 93 318 94 319 
<< m1 >>
rect 100 318 101 319 
<< pdiffusion >>
rect 102 318 103 319 
<< pdiffusion >>
rect 103 318 104 319 
<< pdiffusion >>
rect 104 318 105 319 
<< pdiffusion >>
rect 105 318 106 319 
<< pdiffusion >>
rect 106 318 107 319 
<< pdiffusion >>
rect 107 318 108 319 
<< pdiffusion >>
rect 120 318 121 319 
<< m1 >>
rect 121 318 122 319 
<< pdiffusion >>
rect 121 318 122 319 
<< pdiffusion >>
rect 122 318 123 319 
<< pdiffusion >>
rect 123 318 124 319 
<< pdiffusion >>
rect 124 318 125 319 
<< pdiffusion >>
rect 125 318 126 319 
<< m1 >>
rect 136 318 137 319 
<< pdiffusion >>
rect 138 318 139 319 
<< pdiffusion >>
rect 139 318 140 319 
<< pdiffusion >>
rect 140 318 141 319 
<< pdiffusion >>
rect 141 318 142 319 
<< pdiffusion >>
rect 142 318 143 319 
<< pdiffusion >>
rect 143 318 144 319 
<< m1 >>
rect 148 318 149 319 
<< m1 >>
rect 150 318 151 319 
<< m2 >>
rect 151 318 152 319 
<< m1 >>
rect 154 318 155 319 
<< m1 >>
rect 159 318 160 319 
<< pdiffusion >>
rect 174 318 175 319 
<< pdiffusion >>
rect 175 318 176 319 
<< pdiffusion >>
rect 176 318 177 319 
<< pdiffusion >>
rect 177 318 178 319 
<< pdiffusion >>
rect 178 318 179 319 
<< pdiffusion >>
rect 179 318 180 319 
<< pdiffusion >>
rect 192 318 193 319 
<< pdiffusion >>
rect 193 318 194 319 
<< pdiffusion >>
rect 194 318 195 319 
<< pdiffusion >>
rect 195 318 196 319 
<< pdiffusion >>
rect 196 318 197 319 
<< pdiffusion >>
rect 197 318 198 319 
<< m2 >>
rect 207 318 208 319 
<< m1 >>
rect 208 318 209 319 
<< pdiffusion >>
rect 210 318 211 319 
<< pdiffusion >>
rect 211 318 212 319 
<< pdiffusion >>
rect 212 318 213 319 
<< pdiffusion >>
rect 213 318 214 319 
<< pdiffusion >>
rect 214 318 215 319 
<< pdiffusion >>
rect 215 318 216 319 
<< m1 >>
rect 217 318 218 319 
<< m2 >>
rect 218 318 219 319 
<< m1 >>
rect 223 318 224 319 
<< m1 >>
rect 225 318 226 319 
<< pdiffusion >>
rect 228 318 229 319 
<< pdiffusion >>
rect 229 318 230 319 
<< pdiffusion >>
rect 230 318 231 319 
<< pdiffusion >>
rect 231 318 232 319 
<< pdiffusion >>
rect 232 318 233 319 
<< pdiffusion >>
rect 233 318 234 319 
<< m1 >>
rect 237 318 238 319 
<< m2 >>
rect 243 318 244 319 
<< m1 >>
rect 244 318 245 319 
<< pdiffusion >>
rect 246 318 247 319 
<< pdiffusion >>
rect 247 318 248 319 
<< pdiffusion >>
rect 248 318 249 319 
<< pdiffusion >>
rect 249 318 250 319 
<< pdiffusion >>
rect 250 318 251 319 
<< pdiffusion >>
rect 251 318 252 319 
<< m1 >>
rect 253 318 254 319 
<< m1 >>
rect 257 318 258 319 
<< pdiffusion >>
rect 264 318 265 319 
<< pdiffusion >>
rect 265 318 266 319 
<< pdiffusion >>
rect 266 318 267 319 
<< pdiffusion >>
rect 267 318 268 319 
<< pdiffusion >>
rect 268 318 269 319 
<< pdiffusion >>
rect 269 318 270 319 
<< m1 >>
rect 271 318 272 319 
<< m1 >>
rect 276 318 277 319 
<< m2 >>
rect 279 318 280 319 
<< m1 >>
rect 280 318 281 319 
<< pdiffusion >>
rect 282 318 283 319 
<< pdiffusion >>
rect 283 318 284 319 
<< pdiffusion >>
rect 284 318 285 319 
<< pdiffusion >>
rect 285 318 286 319 
<< pdiffusion >>
rect 286 318 287 319 
<< pdiffusion >>
rect 287 318 288 319 
<< pdiffusion >>
rect 300 318 301 319 
<< pdiffusion >>
rect 301 318 302 319 
<< pdiffusion >>
rect 302 318 303 319 
<< pdiffusion >>
rect 303 318 304 319 
<< pdiffusion >>
rect 304 318 305 319 
<< pdiffusion >>
rect 305 318 306 319 
<< m1 >>
rect 307 318 308 319 
<< pdiffusion >>
rect 318 318 319 319 
<< pdiffusion >>
rect 319 318 320 319 
<< pdiffusion >>
rect 320 318 321 319 
<< pdiffusion >>
rect 321 318 322 319 
<< pdiffusion >>
rect 322 318 323 319 
<< pdiffusion >>
rect 323 318 324 319 
<< m1 >>
rect 334 318 335 319 
<< pdiffusion >>
rect 336 318 337 319 
<< pdiffusion >>
rect 337 318 338 319 
<< pdiffusion >>
rect 338 318 339 319 
<< pdiffusion >>
rect 339 318 340 319 
<< pdiffusion >>
rect 340 318 341 319 
<< pdiffusion >>
rect 341 318 342 319 
<< m1 >>
rect 344 318 345 319 
<< m2 >>
rect 346 318 347 319 
<< m1 >>
rect 347 318 348 319 
<< m1 >>
rect 350 318 351 319 
<< m1 >>
rect 352 318 353 319 
<< m1 >>
rect 366 318 367 319 
<< m2 >>
rect 369 318 370 319 
<< m1 >>
rect 370 318 371 319 
<< pdiffusion >>
rect 372 318 373 319 
<< pdiffusion >>
rect 373 318 374 319 
<< pdiffusion >>
rect 374 318 375 319 
<< pdiffusion >>
rect 375 318 376 319 
<< pdiffusion >>
rect 376 318 377 319 
<< pdiffusion >>
rect 377 318 378 319 
<< m1 >>
rect 379 318 380 319 
<< pdiffusion >>
rect 390 318 391 319 
<< pdiffusion >>
rect 391 318 392 319 
<< pdiffusion >>
rect 392 318 393 319 
<< pdiffusion >>
rect 393 318 394 319 
<< pdiffusion >>
rect 394 318 395 319 
<< pdiffusion >>
rect 395 318 396 319 
<< pdiffusion >>
rect 408 318 409 319 
<< pdiffusion >>
rect 409 318 410 319 
<< pdiffusion >>
rect 410 318 411 319 
<< pdiffusion >>
rect 411 318 412 319 
<< pdiffusion >>
rect 412 318 413 319 
<< pdiffusion >>
rect 413 318 414 319 
<< m1 >>
rect 416 318 417 319 
<< m2 >>
rect 417 318 418 319 
<< m1 >>
rect 420 318 421 319 
<< m1 >>
rect 424 318 425 319 
<< pdiffusion >>
rect 426 318 427 319 
<< m1 >>
rect 427 318 428 319 
<< pdiffusion >>
rect 427 318 428 319 
<< pdiffusion >>
rect 428 318 429 319 
<< pdiffusion >>
rect 429 318 430 319 
<< pdiffusion >>
rect 430 318 431 319 
<< pdiffusion >>
rect 431 318 432 319 
<< m1 >>
rect 433 318 434 319 
<< m1 >>
rect 435 318 436 319 
<< m1 >>
rect 437 318 438 319 
<< m1 >>
rect 439 318 440 319 
<< pdiffusion >>
rect 444 318 445 319 
<< pdiffusion >>
rect 445 318 446 319 
<< pdiffusion >>
rect 446 318 447 319 
<< pdiffusion >>
rect 447 318 448 319 
<< pdiffusion >>
rect 448 318 449 319 
<< pdiffusion >>
rect 449 318 450 319 
<< pdiffusion >>
rect 462 318 463 319 
<< pdiffusion >>
rect 463 318 464 319 
<< pdiffusion >>
rect 464 318 465 319 
<< pdiffusion >>
rect 465 318 466 319 
<< pdiffusion >>
rect 466 318 467 319 
<< pdiffusion >>
rect 467 318 468 319 
<< pdiffusion >>
rect 480 318 481 319 
<< pdiffusion >>
rect 481 318 482 319 
<< pdiffusion >>
rect 482 318 483 319 
<< pdiffusion >>
rect 483 318 484 319 
<< pdiffusion >>
rect 484 318 485 319 
<< pdiffusion >>
rect 485 318 486 319 
<< m1 >>
rect 487 318 488 319 
<< pdiffusion >>
rect 498 318 499 319 
<< pdiffusion >>
rect 499 318 500 319 
<< pdiffusion >>
rect 500 318 501 319 
<< pdiffusion >>
rect 501 318 502 319 
<< pdiffusion >>
rect 502 318 503 319 
<< pdiffusion >>
rect 503 318 504 319 
<< pdiffusion >>
rect 516 318 517 319 
<< pdiffusion >>
rect 517 318 518 319 
<< pdiffusion >>
rect 518 318 519 319 
<< pdiffusion >>
rect 519 318 520 319 
<< pdiffusion >>
rect 520 318 521 319 
<< pdiffusion >>
rect 521 318 522 319 
<< m1 >>
rect 523 318 524 319 
<< pdiffusion >>
rect 12 319 13 320 
<< pdiffusion >>
rect 13 319 14 320 
<< pdiffusion >>
rect 14 319 15 320 
<< pdiffusion >>
rect 15 319 16 320 
<< pdiffusion >>
rect 16 319 17 320 
<< pdiffusion >>
rect 17 319 18 320 
<< m1 >>
rect 19 319 20 320 
<< m1 >>
rect 23 319 24 320 
<< m1 >>
rect 25 319 26 320 
<< pdiffusion >>
rect 30 319 31 320 
<< pdiffusion >>
rect 31 319 32 320 
<< pdiffusion >>
rect 32 319 33 320 
<< pdiffusion >>
rect 33 319 34 320 
<< pdiffusion >>
rect 34 319 35 320 
<< pdiffusion >>
rect 35 319 36 320 
<< m1 >>
rect 44 319 45 320 
<< m1 >>
rect 46 319 47 320 
<< m2 >>
rect 46 319 47 320 
<< pdiffusion >>
rect 48 319 49 320 
<< pdiffusion >>
rect 49 319 50 320 
<< pdiffusion >>
rect 50 319 51 320 
<< pdiffusion >>
rect 51 319 52 320 
<< pdiffusion >>
rect 52 319 53 320 
<< pdiffusion >>
rect 53 319 54 320 
<< m1 >>
rect 55 319 56 320 
<< pdiffusion >>
rect 66 319 67 320 
<< pdiffusion >>
rect 67 319 68 320 
<< pdiffusion >>
rect 68 319 69 320 
<< pdiffusion >>
rect 69 319 70 320 
<< pdiffusion >>
rect 70 319 71 320 
<< pdiffusion >>
rect 71 319 72 320 
<< m1 >>
rect 73 319 74 320 
<< m2 >>
rect 74 319 75 320 
<< pdiffusion >>
rect 84 319 85 320 
<< pdiffusion >>
rect 85 319 86 320 
<< pdiffusion >>
rect 86 319 87 320 
<< pdiffusion >>
rect 87 319 88 320 
<< pdiffusion >>
rect 88 319 89 320 
<< pdiffusion >>
rect 89 319 90 320 
<< m1 >>
rect 93 319 94 320 
<< m1 >>
rect 100 319 101 320 
<< pdiffusion >>
rect 102 319 103 320 
<< pdiffusion >>
rect 103 319 104 320 
<< pdiffusion >>
rect 104 319 105 320 
<< pdiffusion >>
rect 105 319 106 320 
<< pdiffusion >>
rect 106 319 107 320 
<< pdiffusion >>
rect 107 319 108 320 
<< pdiffusion >>
rect 120 319 121 320 
<< pdiffusion >>
rect 121 319 122 320 
<< pdiffusion >>
rect 122 319 123 320 
<< pdiffusion >>
rect 123 319 124 320 
<< pdiffusion >>
rect 124 319 125 320 
<< pdiffusion >>
rect 125 319 126 320 
<< m1 >>
rect 136 319 137 320 
<< pdiffusion >>
rect 138 319 139 320 
<< pdiffusion >>
rect 139 319 140 320 
<< pdiffusion >>
rect 140 319 141 320 
<< pdiffusion >>
rect 141 319 142 320 
<< pdiffusion >>
rect 142 319 143 320 
<< pdiffusion >>
rect 143 319 144 320 
<< m1 >>
rect 148 319 149 320 
<< m1 >>
rect 150 319 151 320 
<< m2 >>
rect 151 319 152 320 
<< m1 >>
rect 154 319 155 320 
<< m1 >>
rect 159 319 160 320 
<< pdiffusion >>
rect 174 319 175 320 
<< pdiffusion >>
rect 175 319 176 320 
<< pdiffusion >>
rect 176 319 177 320 
<< pdiffusion >>
rect 177 319 178 320 
<< pdiffusion >>
rect 178 319 179 320 
<< pdiffusion >>
rect 179 319 180 320 
<< pdiffusion >>
rect 192 319 193 320 
<< pdiffusion >>
rect 193 319 194 320 
<< pdiffusion >>
rect 194 319 195 320 
<< pdiffusion >>
rect 195 319 196 320 
<< pdiffusion >>
rect 196 319 197 320 
<< pdiffusion >>
rect 197 319 198 320 
<< m2 >>
rect 207 319 208 320 
<< m1 >>
rect 208 319 209 320 
<< pdiffusion >>
rect 210 319 211 320 
<< pdiffusion >>
rect 211 319 212 320 
<< pdiffusion >>
rect 212 319 213 320 
<< pdiffusion >>
rect 213 319 214 320 
<< pdiffusion >>
rect 214 319 215 320 
<< pdiffusion >>
rect 215 319 216 320 
<< m1 >>
rect 217 319 218 320 
<< m2 >>
rect 218 319 219 320 
<< m1 >>
rect 223 319 224 320 
<< m1 >>
rect 225 319 226 320 
<< pdiffusion >>
rect 228 319 229 320 
<< pdiffusion >>
rect 229 319 230 320 
<< pdiffusion >>
rect 230 319 231 320 
<< pdiffusion >>
rect 231 319 232 320 
<< pdiffusion >>
rect 232 319 233 320 
<< pdiffusion >>
rect 233 319 234 320 
<< m1 >>
rect 237 319 238 320 
<< m2 >>
rect 243 319 244 320 
<< m1 >>
rect 244 319 245 320 
<< pdiffusion >>
rect 246 319 247 320 
<< pdiffusion >>
rect 247 319 248 320 
<< pdiffusion >>
rect 248 319 249 320 
<< pdiffusion >>
rect 249 319 250 320 
<< pdiffusion >>
rect 250 319 251 320 
<< pdiffusion >>
rect 251 319 252 320 
<< m1 >>
rect 253 319 254 320 
<< m1 >>
rect 257 319 258 320 
<< pdiffusion >>
rect 264 319 265 320 
<< pdiffusion >>
rect 265 319 266 320 
<< pdiffusion >>
rect 266 319 267 320 
<< pdiffusion >>
rect 267 319 268 320 
<< pdiffusion >>
rect 268 319 269 320 
<< pdiffusion >>
rect 269 319 270 320 
<< m1 >>
rect 271 319 272 320 
<< m1 >>
rect 276 319 277 320 
<< m2 >>
rect 276 319 277 320 
<< m2c >>
rect 276 319 277 320 
<< m1 >>
rect 276 319 277 320 
<< m2 >>
rect 276 319 277 320 
<< m2 >>
rect 279 319 280 320 
<< m1 >>
rect 280 319 281 320 
<< pdiffusion >>
rect 282 319 283 320 
<< pdiffusion >>
rect 283 319 284 320 
<< pdiffusion >>
rect 284 319 285 320 
<< pdiffusion >>
rect 285 319 286 320 
<< pdiffusion >>
rect 286 319 287 320 
<< pdiffusion >>
rect 287 319 288 320 
<< pdiffusion >>
rect 300 319 301 320 
<< pdiffusion >>
rect 301 319 302 320 
<< pdiffusion >>
rect 302 319 303 320 
<< pdiffusion >>
rect 303 319 304 320 
<< pdiffusion >>
rect 304 319 305 320 
<< pdiffusion >>
rect 305 319 306 320 
<< m1 >>
rect 307 319 308 320 
<< pdiffusion >>
rect 318 319 319 320 
<< pdiffusion >>
rect 319 319 320 320 
<< pdiffusion >>
rect 320 319 321 320 
<< pdiffusion >>
rect 321 319 322 320 
<< pdiffusion >>
rect 322 319 323 320 
<< pdiffusion >>
rect 323 319 324 320 
<< m1 >>
rect 334 319 335 320 
<< pdiffusion >>
rect 336 319 337 320 
<< pdiffusion >>
rect 337 319 338 320 
<< pdiffusion >>
rect 338 319 339 320 
<< pdiffusion >>
rect 339 319 340 320 
<< pdiffusion >>
rect 340 319 341 320 
<< pdiffusion >>
rect 341 319 342 320 
<< m1 >>
rect 344 319 345 320 
<< m2 >>
rect 346 319 347 320 
<< m1 >>
rect 347 319 348 320 
<< m1 >>
rect 350 319 351 320 
<< m1 >>
rect 352 319 353 320 
<< m1 >>
rect 366 319 367 320 
<< m2 >>
rect 369 319 370 320 
<< m1 >>
rect 370 319 371 320 
<< pdiffusion >>
rect 372 319 373 320 
<< pdiffusion >>
rect 373 319 374 320 
<< pdiffusion >>
rect 374 319 375 320 
<< pdiffusion >>
rect 375 319 376 320 
<< pdiffusion >>
rect 376 319 377 320 
<< pdiffusion >>
rect 377 319 378 320 
<< m1 >>
rect 379 319 380 320 
<< pdiffusion >>
rect 390 319 391 320 
<< pdiffusion >>
rect 391 319 392 320 
<< pdiffusion >>
rect 392 319 393 320 
<< pdiffusion >>
rect 393 319 394 320 
<< pdiffusion >>
rect 394 319 395 320 
<< pdiffusion >>
rect 395 319 396 320 
<< pdiffusion >>
rect 408 319 409 320 
<< pdiffusion >>
rect 409 319 410 320 
<< pdiffusion >>
rect 410 319 411 320 
<< pdiffusion >>
rect 411 319 412 320 
<< pdiffusion >>
rect 412 319 413 320 
<< pdiffusion >>
rect 413 319 414 320 
<< m1 >>
rect 416 319 417 320 
<< m2 >>
rect 417 319 418 320 
<< m1 >>
rect 420 319 421 320 
<< m1 >>
rect 424 319 425 320 
<< pdiffusion >>
rect 426 319 427 320 
<< pdiffusion >>
rect 427 319 428 320 
<< pdiffusion >>
rect 428 319 429 320 
<< pdiffusion >>
rect 429 319 430 320 
<< pdiffusion >>
rect 430 319 431 320 
<< pdiffusion >>
rect 431 319 432 320 
<< m1 >>
rect 433 319 434 320 
<< m1 >>
rect 435 319 436 320 
<< m1 >>
rect 437 319 438 320 
<< m1 >>
rect 439 319 440 320 
<< pdiffusion >>
rect 444 319 445 320 
<< pdiffusion >>
rect 445 319 446 320 
<< pdiffusion >>
rect 446 319 447 320 
<< pdiffusion >>
rect 447 319 448 320 
<< pdiffusion >>
rect 448 319 449 320 
<< pdiffusion >>
rect 449 319 450 320 
<< pdiffusion >>
rect 462 319 463 320 
<< pdiffusion >>
rect 463 319 464 320 
<< pdiffusion >>
rect 464 319 465 320 
<< pdiffusion >>
rect 465 319 466 320 
<< pdiffusion >>
rect 466 319 467 320 
<< pdiffusion >>
rect 467 319 468 320 
<< pdiffusion >>
rect 480 319 481 320 
<< pdiffusion >>
rect 481 319 482 320 
<< pdiffusion >>
rect 482 319 483 320 
<< pdiffusion >>
rect 483 319 484 320 
<< pdiffusion >>
rect 484 319 485 320 
<< pdiffusion >>
rect 485 319 486 320 
<< m1 >>
rect 487 319 488 320 
<< pdiffusion >>
rect 498 319 499 320 
<< pdiffusion >>
rect 499 319 500 320 
<< pdiffusion >>
rect 500 319 501 320 
<< pdiffusion >>
rect 501 319 502 320 
<< pdiffusion >>
rect 502 319 503 320 
<< pdiffusion >>
rect 503 319 504 320 
<< pdiffusion >>
rect 516 319 517 320 
<< pdiffusion >>
rect 517 319 518 320 
<< pdiffusion >>
rect 518 319 519 320 
<< pdiffusion >>
rect 519 319 520 320 
<< pdiffusion >>
rect 520 319 521 320 
<< pdiffusion >>
rect 521 319 522 320 
<< m1 >>
rect 523 319 524 320 
<< pdiffusion >>
rect 12 320 13 321 
<< pdiffusion >>
rect 13 320 14 321 
<< pdiffusion >>
rect 14 320 15 321 
<< pdiffusion >>
rect 15 320 16 321 
<< pdiffusion >>
rect 16 320 17 321 
<< pdiffusion >>
rect 17 320 18 321 
<< m1 >>
rect 19 320 20 321 
<< m1 >>
rect 23 320 24 321 
<< m1 >>
rect 25 320 26 321 
<< pdiffusion >>
rect 30 320 31 321 
<< pdiffusion >>
rect 31 320 32 321 
<< pdiffusion >>
rect 32 320 33 321 
<< pdiffusion >>
rect 33 320 34 321 
<< pdiffusion >>
rect 34 320 35 321 
<< pdiffusion >>
rect 35 320 36 321 
<< m1 >>
rect 44 320 45 321 
<< m1 >>
rect 46 320 47 321 
<< m2 >>
rect 46 320 47 321 
<< pdiffusion >>
rect 48 320 49 321 
<< pdiffusion >>
rect 49 320 50 321 
<< pdiffusion >>
rect 50 320 51 321 
<< pdiffusion >>
rect 51 320 52 321 
<< pdiffusion >>
rect 52 320 53 321 
<< pdiffusion >>
rect 53 320 54 321 
<< m1 >>
rect 55 320 56 321 
<< pdiffusion >>
rect 66 320 67 321 
<< pdiffusion >>
rect 67 320 68 321 
<< pdiffusion >>
rect 68 320 69 321 
<< pdiffusion >>
rect 69 320 70 321 
<< pdiffusion >>
rect 70 320 71 321 
<< pdiffusion >>
rect 71 320 72 321 
<< m1 >>
rect 73 320 74 321 
<< m2 >>
rect 74 320 75 321 
<< pdiffusion >>
rect 84 320 85 321 
<< pdiffusion >>
rect 85 320 86 321 
<< pdiffusion >>
rect 86 320 87 321 
<< pdiffusion >>
rect 87 320 88 321 
<< pdiffusion >>
rect 88 320 89 321 
<< pdiffusion >>
rect 89 320 90 321 
<< m1 >>
rect 93 320 94 321 
<< m1 >>
rect 100 320 101 321 
<< pdiffusion >>
rect 102 320 103 321 
<< pdiffusion >>
rect 103 320 104 321 
<< pdiffusion >>
rect 104 320 105 321 
<< pdiffusion >>
rect 105 320 106 321 
<< pdiffusion >>
rect 106 320 107 321 
<< pdiffusion >>
rect 107 320 108 321 
<< pdiffusion >>
rect 120 320 121 321 
<< pdiffusion >>
rect 121 320 122 321 
<< pdiffusion >>
rect 122 320 123 321 
<< pdiffusion >>
rect 123 320 124 321 
<< pdiffusion >>
rect 124 320 125 321 
<< pdiffusion >>
rect 125 320 126 321 
<< m1 >>
rect 136 320 137 321 
<< pdiffusion >>
rect 138 320 139 321 
<< pdiffusion >>
rect 139 320 140 321 
<< pdiffusion >>
rect 140 320 141 321 
<< pdiffusion >>
rect 141 320 142 321 
<< pdiffusion >>
rect 142 320 143 321 
<< pdiffusion >>
rect 143 320 144 321 
<< m1 >>
rect 148 320 149 321 
<< m1 >>
rect 150 320 151 321 
<< m2 >>
rect 151 320 152 321 
<< m1 >>
rect 154 320 155 321 
<< m1 >>
rect 159 320 160 321 
<< pdiffusion >>
rect 174 320 175 321 
<< pdiffusion >>
rect 175 320 176 321 
<< pdiffusion >>
rect 176 320 177 321 
<< pdiffusion >>
rect 177 320 178 321 
<< pdiffusion >>
rect 178 320 179 321 
<< pdiffusion >>
rect 179 320 180 321 
<< pdiffusion >>
rect 192 320 193 321 
<< pdiffusion >>
rect 193 320 194 321 
<< pdiffusion >>
rect 194 320 195 321 
<< pdiffusion >>
rect 195 320 196 321 
<< pdiffusion >>
rect 196 320 197 321 
<< pdiffusion >>
rect 197 320 198 321 
<< m2 >>
rect 207 320 208 321 
<< m1 >>
rect 208 320 209 321 
<< pdiffusion >>
rect 210 320 211 321 
<< pdiffusion >>
rect 211 320 212 321 
<< pdiffusion >>
rect 212 320 213 321 
<< pdiffusion >>
rect 213 320 214 321 
<< pdiffusion >>
rect 214 320 215 321 
<< pdiffusion >>
rect 215 320 216 321 
<< m1 >>
rect 217 320 218 321 
<< m2 >>
rect 218 320 219 321 
<< m1 >>
rect 223 320 224 321 
<< m1 >>
rect 225 320 226 321 
<< pdiffusion >>
rect 228 320 229 321 
<< pdiffusion >>
rect 229 320 230 321 
<< pdiffusion >>
rect 230 320 231 321 
<< pdiffusion >>
rect 231 320 232 321 
<< pdiffusion >>
rect 232 320 233 321 
<< pdiffusion >>
rect 233 320 234 321 
<< m1 >>
rect 237 320 238 321 
<< m2 >>
rect 243 320 244 321 
<< m1 >>
rect 244 320 245 321 
<< pdiffusion >>
rect 246 320 247 321 
<< pdiffusion >>
rect 247 320 248 321 
<< pdiffusion >>
rect 248 320 249 321 
<< pdiffusion >>
rect 249 320 250 321 
<< pdiffusion >>
rect 250 320 251 321 
<< pdiffusion >>
rect 251 320 252 321 
<< m1 >>
rect 253 320 254 321 
<< m1 >>
rect 257 320 258 321 
<< pdiffusion >>
rect 264 320 265 321 
<< pdiffusion >>
rect 265 320 266 321 
<< pdiffusion >>
rect 266 320 267 321 
<< pdiffusion >>
rect 267 320 268 321 
<< pdiffusion >>
rect 268 320 269 321 
<< pdiffusion >>
rect 269 320 270 321 
<< m1 >>
rect 271 320 272 321 
<< m2 >>
rect 276 320 277 321 
<< m2 >>
rect 279 320 280 321 
<< m1 >>
rect 280 320 281 321 
<< pdiffusion >>
rect 282 320 283 321 
<< pdiffusion >>
rect 283 320 284 321 
<< pdiffusion >>
rect 284 320 285 321 
<< pdiffusion >>
rect 285 320 286 321 
<< pdiffusion >>
rect 286 320 287 321 
<< pdiffusion >>
rect 287 320 288 321 
<< pdiffusion >>
rect 300 320 301 321 
<< pdiffusion >>
rect 301 320 302 321 
<< pdiffusion >>
rect 302 320 303 321 
<< pdiffusion >>
rect 303 320 304 321 
<< pdiffusion >>
rect 304 320 305 321 
<< pdiffusion >>
rect 305 320 306 321 
<< m1 >>
rect 307 320 308 321 
<< pdiffusion >>
rect 318 320 319 321 
<< pdiffusion >>
rect 319 320 320 321 
<< pdiffusion >>
rect 320 320 321 321 
<< pdiffusion >>
rect 321 320 322 321 
<< pdiffusion >>
rect 322 320 323 321 
<< pdiffusion >>
rect 323 320 324 321 
<< m1 >>
rect 334 320 335 321 
<< pdiffusion >>
rect 336 320 337 321 
<< pdiffusion >>
rect 337 320 338 321 
<< pdiffusion >>
rect 338 320 339 321 
<< pdiffusion >>
rect 339 320 340 321 
<< pdiffusion >>
rect 340 320 341 321 
<< pdiffusion >>
rect 341 320 342 321 
<< m1 >>
rect 344 320 345 321 
<< m2 >>
rect 346 320 347 321 
<< m1 >>
rect 347 320 348 321 
<< m1 >>
rect 350 320 351 321 
<< m1 >>
rect 352 320 353 321 
<< m1 >>
rect 366 320 367 321 
<< m2 >>
rect 369 320 370 321 
<< m1 >>
rect 370 320 371 321 
<< pdiffusion >>
rect 372 320 373 321 
<< pdiffusion >>
rect 373 320 374 321 
<< pdiffusion >>
rect 374 320 375 321 
<< pdiffusion >>
rect 375 320 376 321 
<< pdiffusion >>
rect 376 320 377 321 
<< pdiffusion >>
rect 377 320 378 321 
<< m1 >>
rect 379 320 380 321 
<< pdiffusion >>
rect 390 320 391 321 
<< pdiffusion >>
rect 391 320 392 321 
<< pdiffusion >>
rect 392 320 393 321 
<< pdiffusion >>
rect 393 320 394 321 
<< pdiffusion >>
rect 394 320 395 321 
<< pdiffusion >>
rect 395 320 396 321 
<< pdiffusion >>
rect 408 320 409 321 
<< pdiffusion >>
rect 409 320 410 321 
<< pdiffusion >>
rect 410 320 411 321 
<< pdiffusion >>
rect 411 320 412 321 
<< pdiffusion >>
rect 412 320 413 321 
<< pdiffusion >>
rect 413 320 414 321 
<< m1 >>
rect 416 320 417 321 
<< m2 >>
rect 417 320 418 321 
<< m1 >>
rect 420 320 421 321 
<< m1 >>
rect 424 320 425 321 
<< pdiffusion >>
rect 426 320 427 321 
<< pdiffusion >>
rect 427 320 428 321 
<< pdiffusion >>
rect 428 320 429 321 
<< pdiffusion >>
rect 429 320 430 321 
<< pdiffusion >>
rect 430 320 431 321 
<< pdiffusion >>
rect 431 320 432 321 
<< m1 >>
rect 433 320 434 321 
<< m1 >>
rect 435 320 436 321 
<< m1 >>
rect 437 320 438 321 
<< m1 >>
rect 439 320 440 321 
<< pdiffusion >>
rect 444 320 445 321 
<< pdiffusion >>
rect 445 320 446 321 
<< pdiffusion >>
rect 446 320 447 321 
<< pdiffusion >>
rect 447 320 448 321 
<< pdiffusion >>
rect 448 320 449 321 
<< pdiffusion >>
rect 449 320 450 321 
<< pdiffusion >>
rect 462 320 463 321 
<< pdiffusion >>
rect 463 320 464 321 
<< pdiffusion >>
rect 464 320 465 321 
<< pdiffusion >>
rect 465 320 466 321 
<< pdiffusion >>
rect 466 320 467 321 
<< pdiffusion >>
rect 467 320 468 321 
<< pdiffusion >>
rect 480 320 481 321 
<< pdiffusion >>
rect 481 320 482 321 
<< pdiffusion >>
rect 482 320 483 321 
<< pdiffusion >>
rect 483 320 484 321 
<< pdiffusion >>
rect 484 320 485 321 
<< pdiffusion >>
rect 485 320 486 321 
<< m1 >>
rect 487 320 488 321 
<< pdiffusion >>
rect 498 320 499 321 
<< pdiffusion >>
rect 499 320 500 321 
<< pdiffusion >>
rect 500 320 501 321 
<< pdiffusion >>
rect 501 320 502 321 
<< pdiffusion >>
rect 502 320 503 321 
<< pdiffusion >>
rect 503 320 504 321 
<< pdiffusion >>
rect 516 320 517 321 
<< pdiffusion >>
rect 517 320 518 321 
<< pdiffusion >>
rect 518 320 519 321 
<< pdiffusion >>
rect 519 320 520 321 
<< pdiffusion >>
rect 520 320 521 321 
<< pdiffusion >>
rect 521 320 522 321 
<< m1 >>
rect 523 320 524 321 
<< pdiffusion >>
rect 12 321 13 322 
<< pdiffusion >>
rect 13 321 14 322 
<< pdiffusion >>
rect 14 321 15 322 
<< pdiffusion >>
rect 15 321 16 322 
<< pdiffusion >>
rect 16 321 17 322 
<< pdiffusion >>
rect 17 321 18 322 
<< m1 >>
rect 19 321 20 322 
<< m1 >>
rect 23 321 24 322 
<< m1 >>
rect 25 321 26 322 
<< pdiffusion >>
rect 30 321 31 322 
<< pdiffusion >>
rect 31 321 32 322 
<< pdiffusion >>
rect 32 321 33 322 
<< pdiffusion >>
rect 33 321 34 322 
<< pdiffusion >>
rect 34 321 35 322 
<< pdiffusion >>
rect 35 321 36 322 
<< m1 >>
rect 44 321 45 322 
<< m1 >>
rect 46 321 47 322 
<< m2 >>
rect 46 321 47 322 
<< pdiffusion >>
rect 48 321 49 322 
<< pdiffusion >>
rect 49 321 50 322 
<< pdiffusion >>
rect 50 321 51 322 
<< pdiffusion >>
rect 51 321 52 322 
<< pdiffusion >>
rect 52 321 53 322 
<< pdiffusion >>
rect 53 321 54 322 
<< m1 >>
rect 55 321 56 322 
<< pdiffusion >>
rect 66 321 67 322 
<< pdiffusion >>
rect 67 321 68 322 
<< pdiffusion >>
rect 68 321 69 322 
<< pdiffusion >>
rect 69 321 70 322 
<< pdiffusion >>
rect 70 321 71 322 
<< pdiffusion >>
rect 71 321 72 322 
<< m1 >>
rect 73 321 74 322 
<< m2 >>
rect 74 321 75 322 
<< pdiffusion >>
rect 84 321 85 322 
<< pdiffusion >>
rect 85 321 86 322 
<< pdiffusion >>
rect 86 321 87 322 
<< pdiffusion >>
rect 87 321 88 322 
<< pdiffusion >>
rect 88 321 89 322 
<< pdiffusion >>
rect 89 321 90 322 
<< m1 >>
rect 93 321 94 322 
<< m1 >>
rect 100 321 101 322 
<< pdiffusion >>
rect 102 321 103 322 
<< pdiffusion >>
rect 103 321 104 322 
<< pdiffusion >>
rect 104 321 105 322 
<< pdiffusion >>
rect 105 321 106 322 
<< pdiffusion >>
rect 106 321 107 322 
<< pdiffusion >>
rect 107 321 108 322 
<< pdiffusion >>
rect 120 321 121 322 
<< pdiffusion >>
rect 121 321 122 322 
<< pdiffusion >>
rect 122 321 123 322 
<< pdiffusion >>
rect 123 321 124 322 
<< pdiffusion >>
rect 124 321 125 322 
<< pdiffusion >>
rect 125 321 126 322 
<< m1 >>
rect 136 321 137 322 
<< pdiffusion >>
rect 138 321 139 322 
<< pdiffusion >>
rect 139 321 140 322 
<< pdiffusion >>
rect 140 321 141 322 
<< pdiffusion >>
rect 141 321 142 322 
<< pdiffusion >>
rect 142 321 143 322 
<< pdiffusion >>
rect 143 321 144 322 
<< m1 >>
rect 148 321 149 322 
<< m1 >>
rect 150 321 151 322 
<< m2 >>
rect 151 321 152 322 
<< m1 >>
rect 154 321 155 322 
<< m1 >>
rect 159 321 160 322 
<< pdiffusion >>
rect 174 321 175 322 
<< pdiffusion >>
rect 175 321 176 322 
<< pdiffusion >>
rect 176 321 177 322 
<< pdiffusion >>
rect 177 321 178 322 
<< pdiffusion >>
rect 178 321 179 322 
<< pdiffusion >>
rect 179 321 180 322 
<< pdiffusion >>
rect 192 321 193 322 
<< pdiffusion >>
rect 193 321 194 322 
<< pdiffusion >>
rect 194 321 195 322 
<< pdiffusion >>
rect 195 321 196 322 
<< pdiffusion >>
rect 196 321 197 322 
<< pdiffusion >>
rect 197 321 198 322 
<< m2 >>
rect 207 321 208 322 
<< m1 >>
rect 208 321 209 322 
<< pdiffusion >>
rect 210 321 211 322 
<< pdiffusion >>
rect 211 321 212 322 
<< pdiffusion >>
rect 212 321 213 322 
<< pdiffusion >>
rect 213 321 214 322 
<< pdiffusion >>
rect 214 321 215 322 
<< pdiffusion >>
rect 215 321 216 322 
<< m1 >>
rect 217 321 218 322 
<< m2 >>
rect 218 321 219 322 
<< m1 >>
rect 223 321 224 322 
<< m1 >>
rect 225 321 226 322 
<< pdiffusion >>
rect 228 321 229 322 
<< pdiffusion >>
rect 229 321 230 322 
<< pdiffusion >>
rect 230 321 231 322 
<< pdiffusion >>
rect 231 321 232 322 
<< pdiffusion >>
rect 232 321 233 322 
<< pdiffusion >>
rect 233 321 234 322 
<< m1 >>
rect 237 321 238 322 
<< m2 >>
rect 243 321 244 322 
<< m1 >>
rect 244 321 245 322 
<< pdiffusion >>
rect 246 321 247 322 
<< pdiffusion >>
rect 247 321 248 322 
<< pdiffusion >>
rect 248 321 249 322 
<< pdiffusion >>
rect 249 321 250 322 
<< pdiffusion >>
rect 250 321 251 322 
<< pdiffusion >>
rect 251 321 252 322 
<< m1 >>
rect 253 321 254 322 
<< m1 >>
rect 257 321 258 322 
<< pdiffusion >>
rect 264 321 265 322 
<< pdiffusion >>
rect 265 321 266 322 
<< pdiffusion >>
rect 266 321 267 322 
<< pdiffusion >>
rect 267 321 268 322 
<< pdiffusion >>
rect 268 321 269 322 
<< pdiffusion >>
rect 269 321 270 322 
<< m1 >>
rect 271 321 272 322 
<< m1 >>
rect 273 321 274 322 
<< m1 >>
rect 274 321 275 322 
<< m1 >>
rect 275 321 276 322 
<< m1 >>
rect 276 321 277 322 
<< m2 >>
rect 276 321 277 322 
<< m1 >>
rect 277 321 278 322 
<< m1 >>
rect 278 321 279 322 
<< m2 >>
rect 278 321 279 322 
<< m2c >>
rect 278 321 279 322 
<< m1 >>
rect 278 321 279 322 
<< m2 >>
rect 278 321 279 322 
<< m2 >>
rect 279 321 280 322 
<< m1 >>
rect 280 321 281 322 
<< pdiffusion >>
rect 282 321 283 322 
<< pdiffusion >>
rect 283 321 284 322 
<< pdiffusion >>
rect 284 321 285 322 
<< pdiffusion >>
rect 285 321 286 322 
<< pdiffusion >>
rect 286 321 287 322 
<< pdiffusion >>
rect 287 321 288 322 
<< pdiffusion >>
rect 300 321 301 322 
<< pdiffusion >>
rect 301 321 302 322 
<< pdiffusion >>
rect 302 321 303 322 
<< pdiffusion >>
rect 303 321 304 322 
<< pdiffusion >>
rect 304 321 305 322 
<< pdiffusion >>
rect 305 321 306 322 
<< m1 >>
rect 307 321 308 322 
<< pdiffusion >>
rect 318 321 319 322 
<< pdiffusion >>
rect 319 321 320 322 
<< pdiffusion >>
rect 320 321 321 322 
<< pdiffusion >>
rect 321 321 322 322 
<< pdiffusion >>
rect 322 321 323 322 
<< pdiffusion >>
rect 323 321 324 322 
<< m1 >>
rect 334 321 335 322 
<< pdiffusion >>
rect 336 321 337 322 
<< pdiffusion >>
rect 337 321 338 322 
<< pdiffusion >>
rect 338 321 339 322 
<< pdiffusion >>
rect 339 321 340 322 
<< pdiffusion >>
rect 340 321 341 322 
<< pdiffusion >>
rect 341 321 342 322 
<< m1 >>
rect 344 321 345 322 
<< m2 >>
rect 346 321 347 322 
<< m1 >>
rect 347 321 348 322 
<< m1 >>
rect 350 321 351 322 
<< m1 >>
rect 352 321 353 322 
<< m1 >>
rect 366 321 367 322 
<< m2 >>
rect 369 321 370 322 
<< m1 >>
rect 370 321 371 322 
<< pdiffusion >>
rect 372 321 373 322 
<< pdiffusion >>
rect 373 321 374 322 
<< pdiffusion >>
rect 374 321 375 322 
<< pdiffusion >>
rect 375 321 376 322 
<< pdiffusion >>
rect 376 321 377 322 
<< pdiffusion >>
rect 377 321 378 322 
<< m1 >>
rect 379 321 380 322 
<< pdiffusion >>
rect 390 321 391 322 
<< pdiffusion >>
rect 391 321 392 322 
<< pdiffusion >>
rect 392 321 393 322 
<< pdiffusion >>
rect 393 321 394 322 
<< pdiffusion >>
rect 394 321 395 322 
<< pdiffusion >>
rect 395 321 396 322 
<< pdiffusion >>
rect 408 321 409 322 
<< pdiffusion >>
rect 409 321 410 322 
<< pdiffusion >>
rect 410 321 411 322 
<< pdiffusion >>
rect 411 321 412 322 
<< pdiffusion >>
rect 412 321 413 322 
<< pdiffusion >>
rect 413 321 414 322 
<< m1 >>
rect 416 321 417 322 
<< m2 >>
rect 417 321 418 322 
<< m1 >>
rect 420 321 421 322 
<< m1 >>
rect 424 321 425 322 
<< pdiffusion >>
rect 426 321 427 322 
<< pdiffusion >>
rect 427 321 428 322 
<< pdiffusion >>
rect 428 321 429 322 
<< pdiffusion >>
rect 429 321 430 322 
<< pdiffusion >>
rect 430 321 431 322 
<< pdiffusion >>
rect 431 321 432 322 
<< m1 >>
rect 433 321 434 322 
<< m1 >>
rect 435 321 436 322 
<< m1 >>
rect 437 321 438 322 
<< m1 >>
rect 439 321 440 322 
<< pdiffusion >>
rect 444 321 445 322 
<< pdiffusion >>
rect 445 321 446 322 
<< pdiffusion >>
rect 446 321 447 322 
<< pdiffusion >>
rect 447 321 448 322 
<< pdiffusion >>
rect 448 321 449 322 
<< pdiffusion >>
rect 449 321 450 322 
<< pdiffusion >>
rect 462 321 463 322 
<< pdiffusion >>
rect 463 321 464 322 
<< pdiffusion >>
rect 464 321 465 322 
<< pdiffusion >>
rect 465 321 466 322 
<< pdiffusion >>
rect 466 321 467 322 
<< pdiffusion >>
rect 467 321 468 322 
<< pdiffusion >>
rect 480 321 481 322 
<< pdiffusion >>
rect 481 321 482 322 
<< pdiffusion >>
rect 482 321 483 322 
<< pdiffusion >>
rect 483 321 484 322 
<< pdiffusion >>
rect 484 321 485 322 
<< pdiffusion >>
rect 485 321 486 322 
<< m1 >>
rect 487 321 488 322 
<< pdiffusion >>
rect 498 321 499 322 
<< pdiffusion >>
rect 499 321 500 322 
<< pdiffusion >>
rect 500 321 501 322 
<< pdiffusion >>
rect 501 321 502 322 
<< pdiffusion >>
rect 502 321 503 322 
<< pdiffusion >>
rect 503 321 504 322 
<< pdiffusion >>
rect 516 321 517 322 
<< pdiffusion >>
rect 517 321 518 322 
<< pdiffusion >>
rect 518 321 519 322 
<< pdiffusion >>
rect 519 321 520 322 
<< pdiffusion >>
rect 520 321 521 322 
<< pdiffusion >>
rect 521 321 522 322 
<< m1 >>
rect 523 321 524 322 
<< pdiffusion >>
rect 12 322 13 323 
<< pdiffusion >>
rect 13 322 14 323 
<< pdiffusion >>
rect 14 322 15 323 
<< pdiffusion >>
rect 15 322 16 323 
<< pdiffusion >>
rect 16 322 17 323 
<< pdiffusion >>
rect 17 322 18 323 
<< m1 >>
rect 19 322 20 323 
<< m1 >>
rect 23 322 24 323 
<< m1 >>
rect 25 322 26 323 
<< pdiffusion >>
rect 30 322 31 323 
<< pdiffusion >>
rect 31 322 32 323 
<< pdiffusion >>
rect 32 322 33 323 
<< pdiffusion >>
rect 33 322 34 323 
<< pdiffusion >>
rect 34 322 35 323 
<< pdiffusion >>
rect 35 322 36 323 
<< m1 >>
rect 44 322 45 323 
<< m1 >>
rect 46 322 47 323 
<< m2 >>
rect 46 322 47 323 
<< pdiffusion >>
rect 48 322 49 323 
<< pdiffusion >>
rect 49 322 50 323 
<< pdiffusion >>
rect 50 322 51 323 
<< pdiffusion >>
rect 51 322 52 323 
<< pdiffusion >>
rect 52 322 53 323 
<< pdiffusion >>
rect 53 322 54 323 
<< m1 >>
rect 55 322 56 323 
<< pdiffusion >>
rect 66 322 67 323 
<< pdiffusion >>
rect 67 322 68 323 
<< pdiffusion >>
rect 68 322 69 323 
<< pdiffusion >>
rect 69 322 70 323 
<< pdiffusion >>
rect 70 322 71 323 
<< pdiffusion >>
rect 71 322 72 323 
<< m1 >>
rect 73 322 74 323 
<< m2 >>
rect 74 322 75 323 
<< pdiffusion >>
rect 84 322 85 323 
<< pdiffusion >>
rect 85 322 86 323 
<< pdiffusion >>
rect 86 322 87 323 
<< pdiffusion >>
rect 87 322 88 323 
<< pdiffusion >>
rect 88 322 89 323 
<< pdiffusion >>
rect 89 322 90 323 
<< m1 >>
rect 93 322 94 323 
<< m1 >>
rect 100 322 101 323 
<< pdiffusion >>
rect 102 322 103 323 
<< pdiffusion >>
rect 103 322 104 323 
<< pdiffusion >>
rect 104 322 105 323 
<< pdiffusion >>
rect 105 322 106 323 
<< pdiffusion >>
rect 106 322 107 323 
<< pdiffusion >>
rect 107 322 108 323 
<< pdiffusion >>
rect 120 322 121 323 
<< pdiffusion >>
rect 121 322 122 323 
<< pdiffusion >>
rect 122 322 123 323 
<< pdiffusion >>
rect 123 322 124 323 
<< pdiffusion >>
rect 124 322 125 323 
<< pdiffusion >>
rect 125 322 126 323 
<< m1 >>
rect 136 322 137 323 
<< pdiffusion >>
rect 138 322 139 323 
<< pdiffusion >>
rect 139 322 140 323 
<< pdiffusion >>
rect 140 322 141 323 
<< pdiffusion >>
rect 141 322 142 323 
<< pdiffusion >>
rect 142 322 143 323 
<< pdiffusion >>
rect 143 322 144 323 
<< m1 >>
rect 148 322 149 323 
<< m1 >>
rect 150 322 151 323 
<< m2 >>
rect 151 322 152 323 
<< m1 >>
rect 154 322 155 323 
<< m1 >>
rect 159 322 160 323 
<< pdiffusion >>
rect 174 322 175 323 
<< pdiffusion >>
rect 175 322 176 323 
<< pdiffusion >>
rect 176 322 177 323 
<< pdiffusion >>
rect 177 322 178 323 
<< pdiffusion >>
rect 178 322 179 323 
<< pdiffusion >>
rect 179 322 180 323 
<< pdiffusion >>
rect 192 322 193 323 
<< pdiffusion >>
rect 193 322 194 323 
<< pdiffusion >>
rect 194 322 195 323 
<< pdiffusion >>
rect 195 322 196 323 
<< pdiffusion >>
rect 196 322 197 323 
<< pdiffusion >>
rect 197 322 198 323 
<< m2 >>
rect 207 322 208 323 
<< m1 >>
rect 208 322 209 323 
<< pdiffusion >>
rect 210 322 211 323 
<< pdiffusion >>
rect 211 322 212 323 
<< pdiffusion >>
rect 212 322 213 323 
<< pdiffusion >>
rect 213 322 214 323 
<< pdiffusion >>
rect 214 322 215 323 
<< pdiffusion >>
rect 215 322 216 323 
<< m1 >>
rect 217 322 218 323 
<< m2 >>
rect 218 322 219 323 
<< m1 >>
rect 223 322 224 323 
<< m1 >>
rect 225 322 226 323 
<< pdiffusion >>
rect 228 322 229 323 
<< pdiffusion >>
rect 229 322 230 323 
<< pdiffusion >>
rect 230 322 231 323 
<< pdiffusion >>
rect 231 322 232 323 
<< pdiffusion >>
rect 232 322 233 323 
<< pdiffusion >>
rect 233 322 234 323 
<< m1 >>
rect 237 322 238 323 
<< m2 >>
rect 243 322 244 323 
<< m1 >>
rect 244 322 245 323 
<< pdiffusion >>
rect 246 322 247 323 
<< pdiffusion >>
rect 247 322 248 323 
<< pdiffusion >>
rect 248 322 249 323 
<< pdiffusion >>
rect 249 322 250 323 
<< pdiffusion >>
rect 250 322 251 323 
<< pdiffusion >>
rect 251 322 252 323 
<< m1 >>
rect 253 322 254 323 
<< m1 >>
rect 257 322 258 323 
<< pdiffusion >>
rect 264 322 265 323 
<< pdiffusion >>
rect 265 322 266 323 
<< pdiffusion >>
rect 266 322 267 323 
<< pdiffusion >>
rect 267 322 268 323 
<< pdiffusion >>
rect 268 322 269 323 
<< pdiffusion >>
rect 269 322 270 323 
<< m1 >>
rect 271 322 272 323 
<< m1 >>
rect 273 322 274 323 
<< m2 >>
rect 276 322 277 323 
<< m1 >>
rect 280 322 281 323 
<< pdiffusion >>
rect 282 322 283 323 
<< pdiffusion >>
rect 283 322 284 323 
<< pdiffusion >>
rect 284 322 285 323 
<< pdiffusion >>
rect 285 322 286 323 
<< pdiffusion >>
rect 286 322 287 323 
<< pdiffusion >>
rect 287 322 288 323 
<< pdiffusion >>
rect 300 322 301 323 
<< pdiffusion >>
rect 301 322 302 323 
<< pdiffusion >>
rect 302 322 303 323 
<< pdiffusion >>
rect 303 322 304 323 
<< pdiffusion >>
rect 304 322 305 323 
<< pdiffusion >>
rect 305 322 306 323 
<< m1 >>
rect 307 322 308 323 
<< pdiffusion >>
rect 318 322 319 323 
<< pdiffusion >>
rect 319 322 320 323 
<< pdiffusion >>
rect 320 322 321 323 
<< pdiffusion >>
rect 321 322 322 323 
<< pdiffusion >>
rect 322 322 323 323 
<< pdiffusion >>
rect 323 322 324 323 
<< m1 >>
rect 334 322 335 323 
<< pdiffusion >>
rect 336 322 337 323 
<< pdiffusion >>
rect 337 322 338 323 
<< pdiffusion >>
rect 338 322 339 323 
<< pdiffusion >>
rect 339 322 340 323 
<< pdiffusion >>
rect 340 322 341 323 
<< pdiffusion >>
rect 341 322 342 323 
<< m1 >>
rect 344 322 345 323 
<< m2 >>
rect 346 322 347 323 
<< m1 >>
rect 347 322 348 323 
<< m1 >>
rect 350 322 351 323 
<< m1 >>
rect 352 322 353 323 
<< m1 >>
rect 366 322 367 323 
<< m2 >>
rect 366 322 367 323 
<< m2c >>
rect 366 322 367 323 
<< m1 >>
rect 366 322 367 323 
<< m2 >>
rect 366 322 367 323 
<< m2 >>
rect 369 322 370 323 
<< m1 >>
rect 370 322 371 323 
<< pdiffusion >>
rect 372 322 373 323 
<< pdiffusion >>
rect 373 322 374 323 
<< pdiffusion >>
rect 374 322 375 323 
<< pdiffusion >>
rect 375 322 376 323 
<< pdiffusion >>
rect 376 322 377 323 
<< pdiffusion >>
rect 377 322 378 323 
<< m1 >>
rect 379 322 380 323 
<< pdiffusion >>
rect 390 322 391 323 
<< pdiffusion >>
rect 391 322 392 323 
<< pdiffusion >>
rect 392 322 393 323 
<< pdiffusion >>
rect 393 322 394 323 
<< pdiffusion >>
rect 394 322 395 323 
<< pdiffusion >>
rect 395 322 396 323 
<< pdiffusion >>
rect 408 322 409 323 
<< pdiffusion >>
rect 409 322 410 323 
<< pdiffusion >>
rect 410 322 411 323 
<< pdiffusion >>
rect 411 322 412 323 
<< pdiffusion >>
rect 412 322 413 323 
<< pdiffusion >>
rect 413 322 414 323 
<< m1 >>
rect 416 322 417 323 
<< m2 >>
rect 417 322 418 323 
<< m1 >>
rect 420 322 421 323 
<< m2 >>
rect 420 322 421 323 
<< m2c >>
rect 420 322 421 323 
<< m1 >>
rect 420 322 421 323 
<< m2 >>
rect 420 322 421 323 
<< m1 >>
rect 424 322 425 323 
<< m2 >>
rect 424 322 425 323 
<< m2c >>
rect 424 322 425 323 
<< m1 >>
rect 424 322 425 323 
<< m2 >>
rect 424 322 425 323 
<< pdiffusion >>
rect 426 322 427 323 
<< pdiffusion >>
rect 427 322 428 323 
<< pdiffusion >>
rect 428 322 429 323 
<< pdiffusion >>
rect 429 322 430 323 
<< pdiffusion >>
rect 430 322 431 323 
<< pdiffusion >>
rect 431 322 432 323 
<< m1 >>
rect 433 322 434 323 
<< m1 >>
rect 435 322 436 323 
<< m1 >>
rect 437 322 438 323 
<< m1 >>
rect 439 322 440 323 
<< pdiffusion >>
rect 444 322 445 323 
<< pdiffusion >>
rect 445 322 446 323 
<< pdiffusion >>
rect 446 322 447 323 
<< pdiffusion >>
rect 447 322 448 323 
<< pdiffusion >>
rect 448 322 449 323 
<< pdiffusion >>
rect 449 322 450 323 
<< pdiffusion >>
rect 462 322 463 323 
<< pdiffusion >>
rect 463 322 464 323 
<< pdiffusion >>
rect 464 322 465 323 
<< pdiffusion >>
rect 465 322 466 323 
<< pdiffusion >>
rect 466 322 467 323 
<< pdiffusion >>
rect 467 322 468 323 
<< pdiffusion >>
rect 480 322 481 323 
<< pdiffusion >>
rect 481 322 482 323 
<< pdiffusion >>
rect 482 322 483 323 
<< pdiffusion >>
rect 483 322 484 323 
<< pdiffusion >>
rect 484 322 485 323 
<< pdiffusion >>
rect 485 322 486 323 
<< m1 >>
rect 487 322 488 323 
<< pdiffusion >>
rect 498 322 499 323 
<< pdiffusion >>
rect 499 322 500 323 
<< pdiffusion >>
rect 500 322 501 323 
<< pdiffusion >>
rect 501 322 502 323 
<< pdiffusion >>
rect 502 322 503 323 
<< pdiffusion >>
rect 503 322 504 323 
<< pdiffusion >>
rect 516 322 517 323 
<< pdiffusion >>
rect 517 322 518 323 
<< pdiffusion >>
rect 518 322 519 323 
<< pdiffusion >>
rect 519 322 520 323 
<< pdiffusion >>
rect 520 322 521 323 
<< pdiffusion >>
rect 521 322 522 323 
<< m1 >>
rect 523 322 524 323 
<< pdiffusion >>
rect 12 323 13 324 
<< pdiffusion >>
rect 13 323 14 324 
<< pdiffusion >>
rect 14 323 15 324 
<< pdiffusion >>
rect 15 323 16 324 
<< pdiffusion >>
rect 16 323 17 324 
<< pdiffusion >>
rect 17 323 18 324 
<< m1 >>
rect 19 323 20 324 
<< m1 >>
rect 23 323 24 324 
<< m1 >>
rect 25 323 26 324 
<< pdiffusion >>
rect 30 323 31 324 
<< pdiffusion >>
rect 31 323 32 324 
<< pdiffusion >>
rect 32 323 33 324 
<< pdiffusion >>
rect 33 323 34 324 
<< m1 >>
rect 34 323 35 324 
<< pdiffusion >>
rect 34 323 35 324 
<< pdiffusion >>
rect 35 323 36 324 
<< m1 >>
rect 44 323 45 324 
<< m2 >>
rect 44 323 45 324 
<< m2c >>
rect 44 323 45 324 
<< m1 >>
rect 44 323 45 324 
<< m2 >>
rect 44 323 45 324 
<< m1 >>
rect 46 323 47 324 
<< m2 >>
rect 46 323 47 324 
<< pdiffusion >>
rect 48 323 49 324 
<< m1 >>
rect 49 323 50 324 
<< pdiffusion >>
rect 49 323 50 324 
<< pdiffusion >>
rect 50 323 51 324 
<< pdiffusion >>
rect 51 323 52 324 
<< pdiffusion >>
rect 52 323 53 324 
<< pdiffusion >>
rect 53 323 54 324 
<< m1 >>
rect 55 323 56 324 
<< pdiffusion >>
rect 66 323 67 324 
<< m1 >>
rect 67 323 68 324 
<< pdiffusion >>
rect 67 323 68 324 
<< pdiffusion >>
rect 68 323 69 324 
<< pdiffusion >>
rect 69 323 70 324 
<< m1 >>
rect 70 323 71 324 
<< pdiffusion >>
rect 70 323 71 324 
<< pdiffusion >>
rect 71 323 72 324 
<< m1 >>
rect 73 323 74 324 
<< m2 >>
rect 74 323 75 324 
<< pdiffusion >>
rect 84 323 85 324 
<< pdiffusion >>
rect 85 323 86 324 
<< pdiffusion >>
rect 86 323 87 324 
<< pdiffusion >>
rect 87 323 88 324 
<< pdiffusion >>
rect 88 323 89 324 
<< pdiffusion >>
rect 89 323 90 324 
<< m1 >>
rect 93 323 94 324 
<< m1 >>
rect 100 323 101 324 
<< pdiffusion >>
rect 102 323 103 324 
<< pdiffusion >>
rect 103 323 104 324 
<< pdiffusion >>
rect 104 323 105 324 
<< pdiffusion >>
rect 105 323 106 324 
<< pdiffusion >>
rect 106 323 107 324 
<< pdiffusion >>
rect 107 323 108 324 
<< pdiffusion >>
rect 120 323 121 324 
<< pdiffusion >>
rect 121 323 122 324 
<< pdiffusion >>
rect 122 323 123 324 
<< pdiffusion >>
rect 123 323 124 324 
<< m1 >>
rect 124 323 125 324 
<< pdiffusion >>
rect 124 323 125 324 
<< pdiffusion >>
rect 125 323 126 324 
<< m1 >>
rect 136 323 137 324 
<< pdiffusion >>
rect 138 323 139 324 
<< m1 >>
rect 139 323 140 324 
<< pdiffusion >>
rect 139 323 140 324 
<< pdiffusion >>
rect 140 323 141 324 
<< pdiffusion >>
rect 141 323 142 324 
<< pdiffusion >>
rect 142 323 143 324 
<< pdiffusion >>
rect 143 323 144 324 
<< m1 >>
rect 148 323 149 324 
<< m1 >>
rect 150 323 151 324 
<< m2 >>
rect 151 323 152 324 
<< m1 >>
rect 154 323 155 324 
<< m1 >>
rect 159 323 160 324 
<< pdiffusion >>
rect 174 323 175 324 
<< pdiffusion >>
rect 175 323 176 324 
<< pdiffusion >>
rect 176 323 177 324 
<< pdiffusion >>
rect 177 323 178 324 
<< pdiffusion >>
rect 178 323 179 324 
<< pdiffusion >>
rect 179 323 180 324 
<< pdiffusion >>
rect 192 323 193 324 
<< pdiffusion >>
rect 193 323 194 324 
<< pdiffusion >>
rect 194 323 195 324 
<< pdiffusion >>
rect 195 323 196 324 
<< pdiffusion >>
rect 196 323 197 324 
<< pdiffusion >>
rect 197 323 198 324 
<< m2 >>
rect 207 323 208 324 
<< m1 >>
rect 208 323 209 324 
<< pdiffusion >>
rect 210 323 211 324 
<< pdiffusion >>
rect 211 323 212 324 
<< pdiffusion >>
rect 212 323 213 324 
<< pdiffusion >>
rect 213 323 214 324 
<< pdiffusion >>
rect 214 323 215 324 
<< pdiffusion >>
rect 215 323 216 324 
<< m1 >>
rect 217 323 218 324 
<< m2 >>
rect 218 323 219 324 
<< m1 >>
rect 223 323 224 324 
<< m1 >>
rect 225 323 226 324 
<< pdiffusion >>
rect 228 323 229 324 
<< m1 >>
rect 229 323 230 324 
<< pdiffusion >>
rect 229 323 230 324 
<< pdiffusion >>
rect 230 323 231 324 
<< pdiffusion >>
rect 231 323 232 324 
<< pdiffusion >>
rect 232 323 233 324 
<< pdiffusion >>
rect 233 323 234 324 
<< m1 >>
rect 237 323 238 324 
<< m2 >>
rect 243 323 244 324 
<< m1 >>
rect 244 323 245 324 
<< pdiffusion >>
rect 246 323 247 324 
<< pdiffusion >>
rect 247 323 248 324 
<< pdiffusion >>
rect 248 323 249 324 
<< pdiffusion >>
rect 249 323 250 324 
<< m1 >>
rect 250 323 251 324 
<< pdiffusion >>
rect 250 323 251 324 
<< pdiffusion >>
rect 251 323 252 324 
<< m1 >>
rect 253 323 254 324 
<< m1 >>
rect 257 323 258 324 
<< pdiffusion >>
rect 264 323 265 324 
<< pdiffusion >>
rect 265 323 266 324 
<< pdiffusion >>
rect 266 323 267 324 
<< pdiffusion >>
rect 267 323 268 324 
<< pdiffusion >>
rect 268 323 269 324 
<< pdiffusion >>
rect 269 323 270 324 
<< m1 >>
rect 271 323 272 324 
<< m2 >>
rect 271 323 272 324 
<< m2 >>
rect 272 323 273 324 
<< m1 >>
rect 273 323 274 324 
<< m2 >>
rect 273 323 274 324 
<< m2c >>
rect 273 323 274 324 
<< m1 >>
rect 273 323 274 324 
<< m2 >>
rect 273 323 274 324 
<< m1 >>
rect 276 323 277 324 
<< m2 >>
rect 276 323 277 324 
<< m2c >>
rect 276 323 277 324 
<< m1 >>
rect 276 323 277 324 
<< m2 >>
rect 276 323 277 324 
<< m1 >>
rect 280 323 281 324 
<< m2 >>
rect 280 323 281 324 
<< m2c >>
rect 280 323 281 324 
<< m1 >>
rect 280 323 281 324 
<< m2 >>
rect 280 323 281 324 
<< pdiffusion >>
rect 282 323 283 324 
<< m1 >>
rect 283 323 284 324 
<< pdiffusion >>
rect 283 323 284 324 
<< pdiffusion >>
rect 284 323 285 324 
<< pdiffusion >>
rect 285 323 286 324 
<< m1 >>
rect 286 323 287 324 
<< pdiffusion >>
rect 286 323 287 324 
<< pdiffusion >>
rect 287 323 288 324 
<< pdiffusion >>
rect 300 323 301 324 
<< pdiffusion >>
rect 301 323 302 324 
<< pdiffusion >>
rect 302 323 303 324 
<< pdiffusion >>
rect 303 323 304 324 
<< pdiffusion >>
rect 304 323 305 324 
<< pdiffusion >>
rect 305 323 306 324 
<< m1 >>
rect 307 323 308 324 
<< pdiffusion >>
rect 318 323 319 324 
<< pdiffusion >>
rect 319 323 320 324 
<< pdiffusion >>
rect 320 323 321 324 
<< pdiffusion >>
rect 321 323 322 324 
<< pdiffusion >>
rect 322 323 323 324 
<< pdiffusion >>
rect 323 323 324 324 
<< m1 >>
rect 334 323 335 324 
<< pdiffusion >>
rect 336 323 337 324 
<< pdiffusion >>
rect 337 323 338 324 
<< pdiffusion >>
rect 338 323 339 324 
<< pdiffusion >>
rect 339 323 340 324 
<< m1 >>
rect 340 323 341 324 
<< pdiffusion >>
rect 340 323 341 324 
<< pdiffusion >>
rect 341 323 342 324 
<< m1 >>
rect 344 323 345 324 
<< m2 >>
rect 346 323 347 324 
<< m1 >>
rect 347 323 348 324 
<< m1 >>
rect 350 323 351 324 
<< m1 >>
rect 352 323 353 324 
<< m2 >>
rect 366 323 367 324 
<< m2 >>
rect 369 323 370 324 
<< m1 >>
rect 370 323 371 324 
<< pdiffusion >>
rect 372 323 373 324 
<< m1 >>
rect 373 323 374 324 
<< pdiffusion >>
rect 373 323 374 324 
<< pdiffusion >>
rect 374 323 375 324 
<< pdiffusion >>
rect 375 323 376 324 
<< pdiffusion >>
rect 376 323 377 324 
<< pdiffusion >>
rect 377 323 378 324 
<< m1 >>
rect 379 323 380 324 
<< pdiffusion >>
rect 390 323 391 324 
<< pdiffusion >>
rect 391 323 392 324 
<< pdiffusion >>
rect 392 323 393 324 
<< pdiffusion >>
rect 393 323 394 324 
<< pdiffusion >>
rect 394 323 395 324 
<< pdiffusion >>
rect 395 323 396 324 
<< pdiffusion >>
rect 408 323 409 324 
<< pdiffusion >>
rect 409 323 410 324 
<< pdiffusion >>
rect 410 323 411 324 
<< pdiffusion >>
rect 411 323 412 324 
<< m1 >>
rect 412 323 413 324 
<< pdiffusion >>
rect 412 323 413 324 
<< pdiffusion >>
rect 413 323 414 324 
<< m1 >>
rect 416 323 417 324 
<< m2 >>
rect 417 323 418 324 
<< m2 >>
rect 420 323 421 324 
<< m2 >>
rect 422 323 423 324 
<< m2 >>
rect 423 323 424 324 
<< m2 >>
rect 424 323 425 324 
<< pdiffusion >>
rect 426 323 427 324 
<< pdiffusion >>
rect 427 323 428 324 
<< pdiffusion >>
rect 428 323 429 324 
<< pdiffusion >>
rect 429 323 430 324 
<< m1 >>
rect 430 323 431 324 
<< pdiffusion >>
rect 430 323 431 324 
<< pdiffusion >>
rect 431 323 432 324 
<< m1 >>
rect 433 323 434 324 
<< m1 >>
rect 435 323 436 324 
<< m1 >>
rect 437 323 438 324 
<< m1 >>
rect 439 323 440 324 
<< pdiffusion >>
rect 444 323 445 324 
<< pdiffusion >>
rect 445 323 446 324 
<< pdiffusion >>
rect 446 323 447 324 
<< pdiffusion >>
rect 447 323 448 324 
<< pdiffusion >>
rect 448 323 449 324 
<< pdiffusion >>
rect 449 323 450 324 
<< pdiffusion >>
rect 462 323 463 324 
<< pdiffusion >>
rect 463 323 464 324 
<< pdiffusion >>
rect 464 323 465 324 
<< pdiffusion >>
rect 465 323 466 324 
<< pdiffusion >>
rect 466 323 467 324 
<< pdiffusion >>
rect 467 323 468 324 
<< pdiffusion >>
rect 480 323 481 324 
<< pdiffusion >>
rect 481 323 482 324 
<< pdiffusion >>
rect 482 323 483 324 
<< pdiffusion >>
rect 483 323 484 324 
<< m1 >>
rect 484 323 485 324 
<< pdiffusion >>
rect 484 323 485 324 
<< pdiffusion >>
rect 485 323 486 324 
<< m1 >>
rect 487 323 488 324 
<< pdiffusion >>
rect 498 323 499 324 
<< pdiffusion >>
rect 499 323 500 324 
<< pdiffusion >>
rect 500 323 501 324 
<< pdiffusion >>
rect 501 323 502 324 
<< pdiffusion >>
rect 502 323 503 324 
<< pdiffusion >>
rect 503 323 504 324 
<< pdiffusion >>
rect 516 323 517 324 
<< pdiffusion >>
rect 517 323 518 324 
<< pdiffusion >>
rect 518 323 519 324 
<< pdiffusion >>
rect 519 323 520 324 
<< pdiffusion >>
rect 520 323 521 324 
<< pdiffusion >>
rect 521 323 522 324 
<< m1 >>
rect 523 323 524 324 
<< m1 >>
rect 19 324 20 325 
<< m1 >>
rect 23 324 24 325 
<< m1 >>
rect 25 324 26 325 
<< m1 >>
rect 34 324 35 325 
<< m2 >>
rect 44 324 45 325 
<< m1 >>
rect 46 324 47 325 
<< m2 >>
rect 46 324 47 325 
<< m1 >>
rect 49 324 50 325 
<< m1 >>
rect 55 324 56 325 
<< m1 >>
rect 67 324 68 325 
<< m1 >>
rect 70 324 71 325 
<< m1 >>
rect 73 324 74 325 
<< m2 >>
rect 74 324 75 325 
<< m1 >>
rect 93 324 94 325 
<< m1 >>
rect 100 324 101 325 
<< m1 >>
rect 124 324 125 325 
<< m1 >>
rect 136 324 137 325 
<< m1 >>
rect 139 324 140 325 
<< m1 >>
rect 148 324 149 325 
<< m1 >>
rect 150 324 151 325 
<< m2 >>
rect 151 324 152 325 
<< m1 >>
rect 154 324 155 325 
<< m1 >>
rect 159 324 160 325 
<< m2 >>
rect 207 324 208 325 
<< m1 >>
rect 208 324 209 325 
<< m1 >>
rect 217 324 218 325 
<< m2 >>
rect 218 324 219 325 
<< m1 >>
rect 223 324 224 325 
<< m1 >>
rect 225 324 226 325 
<< m1 >>
rect 229 324 230 325 
<< m1 >>
rect 237 324 238 325 
<< m2 >>
rect 243 324 244 325 
<< m1 >>
rect 244 324 245 325 
<< m1 >>
rect 250 324 251 325 
<< m1 >>
rect 253 324 254 325 
<< m1 >>
rect 257 324 258 325 
<< m1 >>
rect 271 324 272 325 
<< m2 >>
rect 271 324 272 325 
<< m2 >>
rect 276 324 277 325 
<< m2 >>
rect 280 324 281 325 
<< m1 >>
rect 283 324 284 325 
<< m1 >>
rect 286 324 287 325 
<< m1 >>
rect 307 324 308 325 
<< m1 >>
rect 334 324 335 325 
<< m1 >>
rect 340 324 341 325 
<< m1 >>
rect 344 324 345 325 
<< m2 >>
rect 346 324 347 325 
<< m1 >>
rect 347 324 348 325 
<< m1 >>
rect 350 324 351 325 
<< m2 >>
rect 350 324 351 325 
<< m2c >>
rect 350 324 351 325 
<< m1 >>
rect 350 324 351 325 
<< m2 >>
rect 350 324 351 325 
<< m2 >>
rect 351 324 352 325 
<< m1 >>
rect 352 324 353 325 
<< m2 >>
rect 352 324 353 325 
<< m2 >>
rect 353 324 354 325 
<< m1 >>
rect 354 324 355 325 
<< m2 >>
rect 354 324 355 325 
<< m1 >>
rect 355 324 356 325 
<< m2 >>
rect 355 324 356 325 
<< m1 >>
rect 356 324 357 325 
<< m2 >>
rect 356 324 357 325 
<< m1 >>
rect 357 324 358 325 
<< m2 >>
rect 357 324 358 325 
<< m1 >>
rect 358 324 359 325 
<< m2 >>
rect 358 324 359 325 
<< m1 >>
rect 359 324 360 325 
<< m2 >>
rect 359 324 360 325 
<< m1 >>
rect 360 324 361 325 
<< m2 >>
rect 360 324 361 325 
<< m1 >>
rect 361 324 362 325 
<< m2 >>
rect 361 324 362 325 
<< m1 >>
rect 362 324 363 325 
<< m2 >>
rect 362 324 363 325 
<< m1 >>
rect 363 324 364 325 
<< m2 >>
rect 363 324 364 325 
<< m1 >>
rect 364 324 365 325 
<< m2 >>
rect 364 324 365 325 
<< m1 >>
rect 365 324 366 325 
<< m1 >>
rect 366 324 367 325 
<< m2 >>
rect 366 324 367 325 
<< m1 >>
rect 367 324 368 325 
<< m1 >>
rect 368 324 369 325 
<< m2 >>
rect 368 324 369 325 
<< m2c >>
rect 368 324 369 325 
<< m1 >>
rect 368 324 369 325 
<< m2 >>
rect 368 324 369 325 
<< m2 >>
rect 369 324 370 325 
<< m1 >>
rect 370 324 371 325 
<< m1 >>
rect 373 324 374 325 
<< m1 >>
rect 379 324 380 325 
<< m1 >>
rect 412 324 413 325 
<< m1 >>
rect 416 324 417 325 
<< m2 >>
rect 417 324 418 325 
<< m1 >>
rect 418 324 419 325 
<< m2 >>
rect 418 324 419 325 
<< m2c >>
rect 418 324 419 325 
<< m1 >>
rect 418 324 419 325 
<< m2 >>
rect 418 324 419 325 
<< m1 >>
rect 419 324 420 325 
<< m1 >>
rect 420 324 421 325 
<< m2 >>
rect 420 324 421 325 
<< m1 >>
rect 421 324 422 325 
<< m1 >>
rect 422 324 423 325 
<< m2 >>
rect 422 324 423 325 
<< m1 >>
rect 423 324 424 325 
<< m1 >>
rect 424 324 425 325 
<< m1 >>
rect 430 324 431 325 
<< m1 >>
rect 433 324 434 325 
<< m1 >>
rect 435 324 436 325 
<< m1 >>
rect 437 324 438 325 
<< m1 >>
rect 439 324 440 325 
<< m1 >>
rect 484 324 485 325 
<< m1 >>
rect 487 324 488 325 
<< m1 >>
rect 523 324 524 325 
<< m1 >>
rect 19 325 20 326 
<< m1 >>
rect 23 325 24 326 
<< m1 >>
rect 25 325 26 326 
<< m1 >>
rect 34 325 35 326 
<< m1 >>
rect 35 325 36 326 
<< m1 >>
rect 36 325 37 326 
<< m1 >>
rect 37 325 38 326 
<< m1 >>
rect 38 325 39 326 
<< m1 >>
rect 39 325 40 326 
<< m1 >>
rect 40 325 41 326 
<< m1 >>
rect 41 325 42 326 
<< m1 >>
rect 42 325 43 326 
<< m1 >>
rect 43 325 44 326 
<< m1 >>
rect 44 325 45 326 
<< m2 >>
rect 44 325 45 326 
<< m1 >>
rect 45 325 46 326 
<< m1 >>
rect 46 325 47 326 
<< m2 >>
rect 46 325 47 326 
<< m2 >>
rect 47 325 48 326 
<< m1 >>
rect 48 325 49 326 
<< m2 >>
rect 48 325 49 326 
<< m2c >>
rect 48 325 49 326 
<< m1 >>
rect 48 325 49 326 
<< m2 >>
rect 48 325 49 326 
<< m1 >>
rect 49 325 50 326 
<< m1 >>
rect 55 325 56 326 
<< m1 >>
rect 67 325 68 326 
<< m1 >>
rect 70 325 71 326 
<< m1 >>
rect 73 325 74 326 
<< m2 >>
rect 74 325 75 326 
<< m1 >>
rect 93 325 94 326 
<< m1 >>
rect 100 325 101 326 
<< m1 >>
rect 124 325 125 326 
<< m2 >>
rect 125 325 126 326 
<< m1 >>
rect 126 325 127 326 
<< m2 >>
rect 126 325 127 326 
<< m2c >>
rect 126 325 127 326 
<< m1 >>
rect 126 325 127 326 
<< m2 >>
rect 126 325 127 326 
<< m1 >>
rect 127 325 128 326 
<< m1 >>
rect 128 325 129 326 
<< m1 >>
rect 129 325 130 326 
<< m1 >>
rect 130 325 131 326 
<< m1 >>
rect 131 325 132 326 
<< m1 >>
rect 132 325 133 326 
<< m1 >>
rect 133 325 134 326 
<< m1 >>
rect 134 325 135 326 
<< m1 >>
rect 135 325 136 326 
<< m1 >>
rect 136 325 137 326 
<< m1 >>
rect 139 325 140 326 
<< m1 >>
rect 148 325 149 326 
<< m1 >>
rect 150 325 151 326 
<< m2 >>
rect 151 325 152 326 
<< m1 >>
rect 154 325 155 326 
<< m1 >>
rect 159 325 160 326 
<< m2 >>
rect 207 325 208 326 
<< m1 >>
rect 208 325 209 326 
<< m1 >>
rect 215 325 216 326 
<< m2 >>
rect 215 325 216 326 
<< m2c >>
rect 215 325 216 326 
<< m1 >>
rect 215 325 216 326 
<< m2 >>
rect 215 325 216 326 
<< m2 >>
rect 216 325 217 326 
<< m1 >>
rect 217 325 218 326 
<< m2 >>
rect 217 325 218 326 
<< m2 >>
rect 218 325 219 326 
<< m1 >>
rect 223 325 224 326 
<< m1 >>
rect 225 325 226 326 
<< m1 >>
rect 229 325 230 326 
<< m1 >>
rect 237 325 238 326 
<< m2 >>
rect 243 325 244 326 
<< m1 >>
rect 244 325 245 326 
<< m1 >>
rect 250 325 251 326 
<< m1 >>
rect 253 325 254 326 
<< m1 >>
rect 257 325 258 326 
<< m1 >>
rect 271 325 272 326 
<< m2 >>
rect 271 325 272 326 
<< m1 >>
rect 272 325 273 326 
<< m1 >>
rect 273 325 274 326 
<< m1 >>
rect 274 325 275 326 
<< m1 >>
rect 275 325 276 326 
<< m1 >>
rect 276 325 277 326 
<< m2 >>
rect 276 325 277 326 
<< m1 >>
rect 277 325 278 326 
<< m1 >>
rect 278 325 279 326 
<< m1 >>
rect 279 325 280 326 
<< m1 >>
rect 280 325 281 326 
<< m2 >>
rect 280 325 281 326 
<< m1 >>
rect 281 325 282 326 
<< m1 >>
rect 282 325 283 326 
<< m1 >>
rect 283 325 284 326 
<< m1 >>
rect 286 325 287 326 
<< m1 >>
rect 307 325 308 326 
<< m1 >>
rect 334 325 335 326 
<< m1 >>
rect 340 325 341 326 
<< m1 >>
rect 344 325 345 326 
<< m2 >>
rect 346 325 347 326 
<< m1 >>
rect 347 325 348 326 
<< m1 >>
rect 352 325 353 326 
<< m1 >>
rect 354 325 355 326 
<< m2 >>
rect 364 325 365 326 
<< m2 >>
rect 366 325 367 326 
<< m1 >>
rect 370 325 371 326 
<< m1 >>
rect 373 325 374 326 
<< m1 >>
rect 379 325 380 326 
<< m1 >>
rect 412 325 413 326 
<< m1 >>
rect 416 325 417 326 
<< m2 >>
rect 420 325 421 326 
<< m2 >>
rect 422 325 423 326 
<< m1 >>
rect 424 325 425 326 
<< m1 >>
rect 430 325 431 326 
<< m1 >>
rect 433 325 434 326 
<< m1 >>
rect 435 325 436 326 
<< m1 >>
rect 437 325 438 326 
<< m1 >>
rect 439 325 440 326 
<< m1 >>
rect 484 325 485 326 
<< m2 >>
rect 485 325 486 326 
<< m1 >>
rect 486 325 487 326 
<< m2 >>
rect 486 325 487 326 
<< m2c >>
rect 486 325 487 326 
<< m1 >>
rect 486 325 487 326 
<< m2 >>
rect 486 325 487 326 
<< m1 >>
rect 487 325 488 326 
<< m1 >>
rect 523 325 524 326 
<< m1 >>
rect 19 326 20 327 
<< m1 >>
rect 23 326 24 327 
<< m1 >>
rect 25 326 26 327 
<< m2 >>
rect 44 326 45 327 
<< m1 >>
rect 55 326 56 327 
<< m1 >>
rect 67 326 68 327 
<< m2 >>
rect 67 326 68 327 
<< m2c >>
rect 67 326 68 327 
<< m1 >>
rect 67 326 68 327 
<< m2 >>
rect 67 326 68 327 
<< m1 >>
rect 70 326 71 327 
<< m1 >>
rect 73 326 74 327 
<< m2 >>
rect 74 326 75 327 
<< m1 >>
rect 91 326 92 327 
<< m2 >>
rect 91 326 92 327 
<< m2c >>
rect 91 326 92 327 
<< m1 >>
rect 91 326 92 327 
<< m2 >>
rect 91 326 92 327 
<< m1 >>
rect 92 326 93 327 
<< m1 >>
rect 93 326 94 327 
<< m1 >>
rect 100 326 101 327 
<< m1 >>
rect 124 326 125 327 
<< m2 >>
rect 125 326 126 327 
<< m1 >>
rect 139 326 140 327 
<< m1 >>
rect 140 326 141 327 
<< m1 >>
rect 141 326 142 327 
<< m1 >>
rect 142 326 143 327 
<< m1 >>
rect 143 326 144 327 
<< m1 >>
rect 144 326 145 327 
<< m1 >>
rect 145 326 146 327 
<< m1 >>
rect 146 326 147 327 
<< m1 >>
rect 147 326 148 327 
<< m1 >>
rect 148 326 149 327 
<< m1 >>
rect 150 326 151 327 
<< m2 >>
rect 151 326 152 327 
<< m1 >>
rect 154 326 155 327 
<< m1 >>
rect 159 326 160 327 
<< m2 >>
rect 207 326 208 327 
<< m1 >>
rect 208 326 209 327 
<< m1 >>
rect 215 326 216 327 
<< m1 >>
rect 217 326 218 327 
<< m1 >>
rect 223 326 224 327 
<< m2 >>
rect 223 326 224 327 
<< m2c >>
rect 223 326 224 327 
<< m1 >>
rect 223 326 224 327 
<< m2 >>
rect 223 326 224 327 
<< m1 >>
rect 225 326 226 327 
<< m2 >>
rect 225 326 226 327 
<< m2c >>
rect 225 326 226 327 
<< m1 >>
rect 225 326 226 327 
<< m2 >>
rect 225 326 226 327 
<< m1 >>
rect 229 326 230 327 
<< m1 >>
rect 237 326 238 327 
<< m2 >>
rect 243 326 244 327 
<< m1 >>
rect 244 326 245 327 
<< m2 >>
rect 249 326 250 327 
<< m1 >>
rect 250 326 251 327 
<< m2 >>
rect 250 326 251 327 
<< m2 >>
rect 251 326 252 327 
<< m2 >>
rect 252 326 253 327 
<< m1 >>
rect 253 326 254 327 
<< m2 >>
rect 253 326 254 327 
<< m2 >>
rect 254 326 255 327 
<< m1 >>
rect 255 326 256 327 
<< m2 >>
rect 255 326 256 327 
<< m2c >>
rect 255 326 256 327 
<< m1 >>
rect 255 326 256 327 
<< m2 >>
rect 255 326 256 327 
<< m1 >>
rect 256 326 257 327 
<< m1 >>
rect 257 326 258 327 
<< m2 >>
rect 271 326 272 327 
<< m2 >>
rect 276 326 277 327 
<< m2 >>
rect 280 326 281 327 
<< m1 >>
rect 286 326 287 327 
<< m1 >>
rect 287 326 288 327 
<< m1 >>
rect 288 326 289 327 
<< m1 >>
rect 289 326 290 327 
<< m2 >>
rect 289 326 290 327 
<< m2c >>
rect 289 326 290 327 
<< m1 >>
rect 289 326 290 327 
<< m2 >>
rect 289 326 290 327 
<< m1 >>
rect 307 326 308 327 
<< m2 >>
rect 307 326 308 327 
<< m2c >>
rect 307 326 308 327 
<< m1 >>
rect 307 326 308 327 
<< m2 >>
rect 307 326 308 327 
<< m1 >>
rect 334 326 335 327 
<< m2 >>
rect 334 326 335 327 
<< m2c >>
rect 334 326 335 327 
<< m1 >>
rect 334 326 335 327 
<< m2 >>
rect 334 326 335 327 
<< m1 >>
rect 340 326 341 327 
<< m1 >>
rect 344 326 345 327 
<< m2 >>
rect 346 326 347 327 
<< m1 >>
rect 347 326 348 327 
<< m2 >>
rect 351 326 352 327 
<< m1 >>
rect 352 326 353 327 
<< m2 >>
rect 352 326 353 327 
<< m2 >>
rect 353 326 354 327 
<< m1 >>
rect 354 326 355 327 
<< m2 >>
rect 354 326 355 327 
<< m2c >>
rect 354 326 355 327 
<< m1 >>
rect 354 326 355 327 
<< m2 >>
rect 354 326 355 327 
<< m1 >>
rect 364 326 365 327 
<< m2 >>
rect 364 326 365 327 
<< m2c >>
rect 364 326 365 327 
<< m1 >>
rect 364 326 365 327 
<< m2 >>
rect 364 326 365 327 
<< m1 >>
rect 366 326 367 327 
<< m2 >>
rect 366 326 367 327 
<< m2c >>
rect 366 326 367 327 
<< m1 >>
rect 366 326 367 327 
<< m2 >>
rect 366 326 367 327 
<< m1 >>
rect 370 326 371 327 
<< m2 >>
rect 370 326 371 327 
<< m2c >>
rect 370 326 371 327 
<< m1 >>
rect 370 326 371 327 
<< m2 >>
rect 370 326 371 327 
<< m1 >>
rect 372 326 373 327 
<< m2 >>
rect 372 326 373 327 
<< m2c >>
rect 372 326 373 327 
<< m1 >>
rect 372 326 373 327 
<< m2 >>
rect 372 326 373 327 
<< m1 >>
rect 373 326 374 327 
<< m1 >>
rect 379 326 380 327 
<< m2 >>
rect 379 326 380 327 
<< m2c >>
rect 379 326 380 327 
<< m1 >>
rect 379 326 380 327 
<< m2 >>
rect 379 326 380 327 
<< m1 >>
rect 412 326 413 327 
<< m1 >>
rect 416 326 417 327 
<< m2 >>
rect 416 326 417 327 
<< m2c >>
rect 416 326 417 327 
<< m1 >>
rect 416 326 417 327 
<< m2 >>
rect 416 326 417 327 
<< m1 >>
rect 418 326 419 327 
<< m2 >>
rect 418 326 419 327 
<< m2c >>
rect 418 326 419 327 
<< m1 >>
rect 418 326 419 327 
<< m2 >>
rect 418 326 419 327 
<< m1 >>
rect 419 326 420 327 
<< m1 >>
rect 420 326 421 327 
<< m2 >>
rect 420 326 421 327 
<< m2c >>
rect 420 326 421 327 
<< m1 >>
rect 420 326 421 327 
<< m2 >>
rect 420 326 421 327 
<< m1 >>
rect 422 326 423 327 
<< m2 >>
rect 422 326 423 327 
<< m2c >>
rect 422 326 423 327 
<< m1 >>
rect 422 326 423 327 
<< m2 >>
rect 422 326 423 327 
<< m1 >>
rect 424 326 425 327 
<< m2 >>
rect 424 326 425 327 
<< m2c >>
rect 424 326 425 327 
<< m1 >>
rect 424 326 425 327 
<< m2 >>
rect 424 326 425 327 
<< m1 >>
rect 430 326 431 327 
<< m1 >>
rect 431 326 432 327 
<< m2 >>
rect 431 326 432 327 
<< m2c >>
rect 431 326 432 327 
<< m1 >>
rect 431 326 432 327 
<< m2 >>
rect 431 326 432 327 
<< m1 >>
rect 433 326 434 327 
<< m2 >>
rect 433 326 434 327 
<< m2c >>
rect 433 326 434 327 
<< m1 >>
rect 433 326 434 327 
<< m2 >>
rect 433 326 434 327 
<< m1 >>
rect 435 326 436 327 
<< m2 >>
rect 435 326 436 327 
<< m2c >>
rect 435 326 436 327 
<< m1 >>
rect 435 326 436 327 
<< m2 >>
rect 435 326 436 327 
<< m1 >>
rect 437 326 438 327 
<< m2 >>
rect 437 326 438 327 
<< m2c >>
rect 437 326 438 327 
<< m1 >>
rect 437 326 438 327 
<< m2 >>
rect 437 326 438 327 
<< m1 >>
rect 439 326 440 327 
<< m2 >>
rect 439 326 440 327 
<< m2c >>
rect 439 326 440 327 
<< m1 >>
rect 439 326 440 327 
<< m2 >>
rect 439 326 440 327 
<< m1 >>
rect 484 326 485 327 
<< m2 >>
rect 485 326 486 327 
<< m1 >>
rect 523 326 524 327 
<< m1 >>
rect 19 327 20 328 
<< m1 >>
rect 23 327 24 328 
<< m1 >>
rect 25 327 26 328 
<< m1 >>
rect 44 327 45 328 
<< m2 >>
rect 44 327 45 328 
<< m2c >>
rect 44 327 45 328 
<< m1 >>
rect 44 327 45 328 
<< m2 >>
rect 44 327 45 328 
<< m1 >>
rect 55 327 56 328 
<< m2 >>
rect 67 327 68 328 
<< m1 >>
rect 70 327 71 328 
<< m1 >>
rect 73 327 74 328 
<< m2 >>
rect 74 327 75 328 
<< m2 >>
rect 91 327 92 328 
<< m1 >>
rect 100 327 101 328 
<< m1 >>
rect 124 327 125 328 
<< m2 >>
rect 125 327 126 328 
<< m1 >>
rect 150 327 151 328 
<< m2 >>
rect 151 327 152 328 
<< m1 >>
rect 154 327 155 328 
<< m1 >>
rect 159 327 160 328 
<< m2 >>
rect 207 327 208 328 
<< m1 >>
rect 208 327 209 328 
<< m1 >>
rect 215 327 216 328 
<< m1 >>
rect 217 327 218 328 
<< m2 >>
rect 223 327 224 328 
<< m2 >>
rect 225 327 226 328 
<< m1 >>
rect 229 327 230 328 
<< m1 >>
rect 237 327 238 328 
<< m2 >>
rect 243 327 244 328 
<< m1 >>
rect 244 327 245 328 
<< m2 >>
rect 249 327 250 328 
<< m1 >>
rect 250 327 251 328 
<< m1 >>
rect 253 327 254 328 
<< m2 >>
rect 271 327 272 328 
<< m2 >>
rect 276 327 277 328 
<< m2 >>
rect 280 327 281 328 
<< m2 >>
rect 289 327 290 328 
<< m2 >>
rect 307 327 308 328 
<< m2 >>
rect 334 327 335 328 
<< m1 >>
rect 340 327 341 328 
<< m1 >>
rect 344 327 345 328 
<< m2 >>
rect 346 327 347 328 
<< m1 >>
rect 347 327 348 328 
<< m2 >>
rect 351 327 352 328 
<< m1 >>
rect 352 327 353 328 
<< m2 >>
rect 364 327 365 328 
<< m2 >>
rect 366 327 367 328 
<< m2 >>
rect 370 327 371 328 
<< m2 >>
rect 372 327 373 328 
<< m2 >>
rect 379 327 380 328 
<< m1 >>
rect 412 327 413 328 
<< m2 >>
rect 416 327 417 328 
<< m2 >>
rect 418 327 419 328 
<< m2 >>
rect 422 327 423 328 
<< m2 >>
rect 424 327 425 328 
<< m2 >>
rect 431 327 432 328 
<< m2 >>
rect 433 327 434 328 
<< m2 >>
rect 435 327 436 328 
<< m2 >>
rect 437 327 438 328 
<< m2 >>
rect 439 327 440 328 
<< m1 >>
rect 484 327 485 328 
<< m2 >>
rect 485 327 486 328 
<< m1 >>
rect 523 327 524 328 
<< m1 >>
rect 19 328 20 329 
<< m1 >>
rect 23 328 24 329 
<< m1 >>
rect 25 328 26 329 
<< m1 >>
rect 44 328 45 329 
<< m1 >>
rect 55 328 56 329 
<< m1 >>
rect 56 328 57 329 
<< m1 >>
rect 57 328 58 329 
<< m1 >>
rect 58 328 59 329 
<< m1 >>
rect 59 328 60 329 
<< m1 >>
rect 60 328 61 329 
<< m1 >>
rect 61 328 62 329 
<< m1 >>
rect 62 328 63 329 
<< m1 >>
rect 63 328 64 329 
<< m1 >>
rect 64 328 65 329 
<< m1 >>
rect 65 328 66 329 
<< m1 >>
rect 66 328 67 329 
<< m1 >>
rect 67 328 68 329 
<< m2 >>
rect 67 328 68 329 
<< m1 >>
rect 68 328 69 329 
<< m1 >>
rect 69 328 70 329 
<< m1 >>
rect 70 328 71 329 
<< m1 >>
rect 73 328 74 329 
<< m2 >>
rect 74 328 75 329 
<< m1 >>
rect 88 328 89 329 
<< m1 >>
rect 89 328 90 329 
<< m1 >>
rect 90 328 91 329 
<< m1 >>
rect 91 328 92 329 
<< m2 >>
rect 91 328 92 329 
<< m1 >>
rect 92 328 93 329 
<< m1 >>
rect 93 328 94 329 
<< m1 >>
rect 94 328 95 329 
<< m1 >>
rect 95 328 96 329 
<< m1 >>
rect 96 328 97 329 
<< m1 >>
rect 97 328 98 329 
<< m1 >>
rect 98 328 99 329 
<< m2 >>
rect 98 328 99 329 
<< m2c >>
rect 98 328 99 329 
<< m1 >>
rect 98 328 99 329 
<< m2 >>
rect 98 328 99 329 
<< m2 >>
rect 99 328 100 329 
<< m1 >>
rect 100 328 101 329 
<< m2 >>
rect 100 328 101 329 
<< m2 >>
rect 101 328 102 329 
<< m1 >>
rect 102 328 103 329 
<< m2 >>
rect 102 328 103 329 
<< m2c >>
rect 102 328 103 329 
<< m1 >>
rect 102 328 103 329 
<< m2 >>
rect 102 328 103 329 
<< m1 >>
rect 103 328 104 329 
<< m1 >>
rect 104 328 105 329 
<< m1 >>
rect 105 328 106 329 
<< m1 >>
rect 106 328 107 329 
<< m1 >>
rect 107 328 108 329 
<< m1 >>
rect 108 328 109 329 
<< m1 >>
rect 109 328 110 329 
<< m1 >>
rect 110 328 111 329 
<< m1 >>
rect 111 328 112 329 
<< m1 >>
rect 112 328 113 329 
<< m1 >>
rect 113 328 114 329 
<< m1 >>
rect 114 328 115 329 
<< m1 >>
rect 115 328 116 329 
<< m1 >>
rect 116 328 117 329 
<< m1 >>
rect 117 328 118 329 
<< m1 >>
rect 118 328 119 329 
<< m1 >>
rect 119 328 120 329 
<< m1 >>
rect 120 328 121 329 
<< m1 >>
rect 121 328 122 329 
<< m1 >>
rect 122 328 123 329 
<< m1 >>
rect 123 328 124 329 
<< m1 >>
rect 124 328 125 329 
<< m2 >>
rect 125 328 126 329 
<< m1 >>
rect 146 328 147 329 
<< m1 >>
rect 147 328 148 329 
<< m1 >>
rect 148 328 149 329 
<< m2 >>
rect 148 328 149 329 
<< m2c >>
rect 148 328 149 329 
<< m1 >>
rect 148 328 149 329 
<< m2 >>
rect 148 328 149 329 
<< m2 >>
rect 149 328 150 329 
<< m1 >>
rect 150 328 151 329 
<< m2 >>
rect 150 328 151 329 
<< m2 >>
rect 151 328 152 329 
<< m1 >>
rect 154 328 155 329 
<< m1 >>
rect 159 328 160 329 
<< m2 >>
rect 207 328 208 329 
<< m1 >>
rect 208 328 209 329 
<< m1 >>
rect 209 328 210 329 
<< m1 >>
rect 210 328 211 329 
<< m1 >>
rect 211 328 212 329 
<< m1 >>
rect 212 328 213 329 
<< m1 >>
rect 213 328 214 329 
<< m2 >>
rect 213 328 214 329 
<< m2c >>
rect 213 328 214 329 
<< m1 >>
rect 213 328 214 329 
<< m2 >>
rect 213 328 214 329 
<< m2 >>
rect 214 328 215 329 
<< m1 >>
rect 215 328 216 329 
<< m2 >>
rect 215 328 216 329 
<< m2 >>
rect 216 328 217 329 
<< m1 >>
rect 217 328 218 329 
<< m2 >>
rect 217 328 218 329 
<< m2 >>
rect 218 328 219 329 
<< m1 >>
rect 219 328 220 329 
<< m2 >>
rect 219 328 220 329 
<< m2c >>
rect 219 328 220 329 
<< m1 >>
rect 219 328 220 329 
<< m2 >>
rect 219 328 220 329 
<< m1 >>
rect 221 328 222 329 
<< m2 >>
rect 221 328 222 329 
<< m2c >>
rect 221 328 222 329 
<< m1 >>
rect 221 328 222 329 
<< m2 >>
rect 221 328 222 329 
<< m1 >>
rect 222 328 223 329 
<< m1 >>
rect 223 328 224 329 
<< m2 >>
rect 223 328 224 329 
<< m1 >>
rect 224 328 225 329 
<< m1 >>
rect 225 328 226 329 
<< m2 >>
rect 225 328 226 329 
<< m1 >>
rect 226 328 227 329 
<< m1 >>
rect 227 328 228 329 
<< m1 >>
rect 228 328 229 329 
<< m1 >>
rect 229 328 230 329 
<< m1 >>
rect 235 328 236 329 
<< m2 >>
rect 235 328 236 329 
<< m2c >>
rect 235 328 236 329 
<< m1 >>
rect 235 328 236 329 
<< m2 >>
rect 235 328 236 329 
<< m1 >>
rect 236 328 237 329 
<< m1 >>
rect 237 328 238 329 
<< m2 >>
rect 243 328 244 329 
<< m1 >>
rect 244 328 245 329 
<< m1 >>
rect 245 328 246 329 
<< m1 >>
rect 246 328 247 329 
<< m1 >>
rect 247 328 248 329 
<< m1 >>
rect 248 328 249 329 
<< m1 >>
rect 249 328 250 329 
<< m2 >>
rect 249 328 250 329 
<< m1 >>
rect 250 328 251 329 
<< m1 >>
rect 253 328 254 329 
<< m1 >>
rect 254 328 255 329 
<< m1 >>
rect 255 328 256 329 
<< m1 >>
rect 256 328 257 329 
<< m1 >>
rect 257 328 258 329 
<< m1 >>
rect 258 328 259 329 
<< m1 >>
rect 259 328 260 329 
<< m1 >>
rect 260 328 261 329 
<< m1 >>
rect 261 328 262 329 
<< m1 >>
rect 262 328 263 329 
<< m1 >>
rect 263 328 264 329 
<< m1 >>
rect 264 328 265 329 
<< m1 >>
rect 265 328 266 329 
<< m1 >>
rect 266 328 267 329 
<< m1 >>
rect 267 328 268 329 
<< m1 >>
rect 268 328 269 329 
<< m1 >>
rect 269 328 270 329 
<< m1 >>
rect 270 328 271 329 
<< m1 >>
rect 271 328 272 329 
<< m2 >>
rect 271 328 272 329 
<< m1 >>
rect 272 328 273 329 
<< m1 >>
rect 273 328 274 329 
<< m1 >>
rect 274 328 275 329 
<< m1 >>
rect 275 328 276 329 
<< m1 >>
rect 276 328 277 329 
<< m2 >>
rect 276 328 277 329 
<< m1 >>
rect 277 328 278 329 
<< m1 >>
rect 278 328 279 329 
<< m1 >>
rect 279 328 280 329 
<< m1 >>
rect 280 328 281 329 
<< m2 >>
rect 280 328 281 329 
<< m1 >>
rect 281 328 282 329 
<< m1 >>
rect 282 328 283 329 
<< m1 >>
rect 283 328 284 329 
<< m1 >>
rect 284 328 285 329 
<< m1 >>
rect 285 328 286 329 
<< m1 >>
rect 286 328 287 329 
<< m1 >>
rect 287 328 288 329 
<< m1 >>
rect 288 328 289 329 
<< m1 >>
rect 289 328 290 329 
<< m2 >>
rect 289 328 290 329 
<< m1 >>
rect 290 328 291 329 
<< m1 >>
rect 291 328 292 329 
<< m1 >>
rect 292 328 293 329 
<< m1 >>
rect 293 328 294 329 
<< m1 >>
rect 294 328 295 329 
<< m1 >>
rect 295 328 296 329 
<< m1 >>
rect 296 328 297 329 
<< m1 >>
rect 297 328 298 329 
<< m1 >>
rect 298 328 299 329 
<< m1 >>
rect 299 328 300 329 
<< m1 >>
rect 300 328 301 329 
<< m1 >>
rect 301 328 302 329 
<< m1 >>
rect 302 328 303 329 
<< m1 >>
rect 303 328 304 329 
<< m1 >>
rect 304 328 305 329 
<< m1 >>
rect 305 328 306 329 
<< m1 >>
rect 306 328 307 329 
<< m1 >>
rect 307 328 308 329 
<< m2 >>
rect 307 328 308 329 
<< m1 >>
rect 308 328 309 329 
<< m1 >>
rect 309 328 310 329 
<< m1 >>
rect 310 328 311 329 
<< m1 >>
rect 311 328 312 329 
<< m1 >>
rect 312 328 313 329 
<< m1 >>
rect 313 328 314 329 
<< m1 >>
rect 314 328 315 329 
<< m1 >>
rect 315 328 316 329 
<< m1 >>
rect 316 328 317 329 
<< m1 >>
rect 317 328 318 329 
<< m1 >>
rect 318 328 319 329 
<< m1 >>
rect 319 328 320 329 
<< m1 >>
rect 320 328 321 329 
<< m1 >>
rect 321 328 322 329 
<< m1 >>
rect 322 328 323 329 
<< m1 >>
rect 323 328 324 329 
<< m1 >>
rect 324 328 325 329 
<< m1 >>
rect 325 328 326 329 
<< m1 >>
rect 326 328 327 329 
<< m1 >>
rect 327 328 328 329 
<< m1 >>
rect 328 328 329 329 
<< m1 >>
rect 329 328 330 329 
<< m1 >>
rect 330 328 331 329 
<< m1 >>
rect 331 328 332 329 
<< m1 >>
rect 332 328 333 329 
<< m1 >>
rect 333 328 334 329 
<< m1 >>
rect 334 328 335 329 
<< m2 >>
rect 334 328 335 329 
<< m1 >>
rect 335 328 336 329 
<< m1 >>
rect 336 328 337 329 
<< m1 >>
rect 337 328 338 329 
<< m1 >>
rect 338 328 339 329 
<< m1 >>
rect 339 328 340 329 
<< m1 >>
rect 340 328 341 329 
<< m2 >>
rect 343 328 344 329 
<< m1 >>
rect 344 328 345 329 
<< m2 >>
rect 344 328 345 329 
<< m2 >>
rect 345 328 346 329 
<< m2 >>
rect 346 328 347 329 
<< m1 >>
rect 347 328 348 329 
<< m2 >>
rect 351 328 352 329 
<< m1 >>
rect 352 328 353 329 
<< m1 >>
rect 353 328 354 329 
<< m1 >>
rect 354 328 355 329 
<< m1 >>
rect 355 328 356 329 
<< m1 >>
rect 356 328 357 329 
<< m1 >>
rect 357 328 358 329 
<< m1 >>
rect 358 328 359 329 
<< m1 >>
rect 359 328 360 329 
<< m1 >>
rect 360 328 361 329 
<< m1 >>
rect 361 328 362 329 
<< m1 >>
rect 362 328 363 329 
<< m1 >>
rect 363 328 364 329 
<< m1 >>
rect 364 328 365 329 
<< m2 >>
rect 364 328 365 329 
<< m1 >>
rect 365 328 366 329 
<< m1 >>
rect 366 328 367 329 
<< m2 >>
rect 366 328 367 329 
<< m1 >>
rect 367 328 368 329 
<< m1 >>
rect 368 328 369 329 
<< m1 >>
rect 369 328 370 329 
<< m1 >>
rect 370 328 371 329 
<< m2 >>
rect 370 328 371 329 
<< m1 >>
rect 371 328 372 329 
<< m1 >>
rect 372 328 373 329 
<< m2 >>
rect 372 328 373 329 
<< m1 >>
rect 373 328 374 329 
<< m1 >>
rect 374 328 375 329 
<< m1 >>
rect 375 328 376 329 
<< m1 >>
rect 376 328 377 329 
<< m1 >>
rect 377 328 378 329 
<< m1 >>
rect 378 328 379 329 
<< m1 >>
rect 379 328 380 329 
<< m2 >>
rect 379 328 380 329 
<< m1 >>
rect 380 328 381 329 
<< m2 >>
rect 380 328 381 329 
<< m1 >>
rect 381 328 382 329 
<< m2 >>
rect 381 328 382 329 
<< m1 >>
rect 382 328 383 329 
<< m2 >>
rect 382 328 383 329 
<< m1 >>
rect 383 328 384 329 
<< m2 >>
rect 383 328 384 329 
<< m1 >>
rect 384 328 385 329 
<< m2 >>
rect 384 328 385 329 
<< m1 >>
rect 385 328 386 329 
<< m2 >>
rect 385 328 386 329 
<< m1 >>
rect 386 328 387 329 
<< m2 >>
rect 386 328 387 329 
<< m1 >>
rect 387 328 388 329 
<< m2 >>
rect 387 328 388 329 
<< m1 >>
rect 388 328 389 329 
<< m2 >>
rect 388 328 389 329 
<< m1 >>
rect 389 328 390 329 
<< m2 >>
rect 389 328 390 329 
<< m1 >>
rect 390 328 391 329 
<< m2 >>
rect 390 328 391 329 
<< m1 >>
rect 391 328 392 329 
<< m2 >>
rect 391 328 392 329 
<< m1 >>
rect 392 328 393 329 
<< m2 >>
rect 392 328 393 329 
<< m1 >>
rect 393 328 394 329 
<< m2 >>
rect 393 328 394 329 
<< m1 >>
rect 394 328 395 329 
<< m2 >>
rect 394 328 395 329 
<< m1 >>
rect 395 328 396 329 
<< m2 >>
rect 395 328 396 329 
<< m1 >>
rect 396 328 397 329 
<< m2 >>
rect 396 328 397 329 
<< m1 >>
rect 397 328 398 329 
<< m2 >>
rect 397 328 398 329 
<< m1 >>
rect 398 328 399 329 
<< m2 >>
rect 398 328 399 329 
<< m1 >>
rect 399 328 400 329 
<< m2 >>
rect 399 328 400 329 
<< m1 >>
rect 400 328 401 329 
<< m2 >>
rect 400 328 401 329 
<< m1 >>
rect 401 328 402 329 
<< m2 >>
rect 401 328 402 329 
<< m1 >>
rect 402 328 403 329 
<< m2 >>
rect 402 328 403 329 
<< m1 >>
rect 403 328 404 329 
<< m2 >>
rect 403 328 404 329 
<< m1 >>
rect 404 328 405 329 
<< m2 >>
rect 404 328 405 329 
<< m1 >>
rect 405 328 406 329 
<< m2 >>
rect 405 328 406 329 
<< m1 >>
rect 406 328 407 329 
<< m2 >>
rect 406 328 407 329 
<< m1 >>
rect 407 328 408 329 
<< m2 >>
rect 407 328 408 329 
<< m1 >>
rect 408 328 409 329 
<< m2 >>
rect 408 328 409 329 
<< m1 >>
rect 409 328 410 329 
<< m2 >>
rect 409 328 410 329 
<< m1 >>
rect 410 328 411 329 
<< m2 >>
rect 410 328 411 329 
<< m1 >>
rect 411 328 412 329 
<< m2 >>
rect 411 328 412 329 
<< m1 >>
rect 412 328 413 329 
<< m2 >>
rect 412 328 413 329 
<< m2 >>
rect 413 328 414 329 
<< m1 >>
rect 414 328 415 329 
<< m2 >>
rect 414 328 415 329 
<< m2c >>
rect 414 328 415 329 
<< m1 >>
rect 414 328 415 329 
<< m2 >>
rect 414 328 415 329 
<< m1 >>
rect 415 328 416 329 
<< m1 >>
rect 416 328 417 329 
<< m2 >>
rect 416 328 417 329 
<< m1 >>
rect 417 328 418 329 
<< m1 >>
rect 418 328 419 329 
<< m2 >>
rect 418 328 419 329 
<< m1 >>
rect 419 328 420 329 
<< m1 >>
rect 420 328 421 329 
<< m1 >>
rect 421 328 422 329 
<< m1 >>
rect 422 328 423 329 
<< m2 >>
rect 422 328 423 329 
<< m1 >>
rect 423 328 424 329 
<< m1 >>
rect 424 328 425 329 
<< m2 >>
rect 424 328 425 329 
<< m1 >>
rect 425 328 426 329 
<< m1 >>
rect 426 328 427 329 
<< m1 >>
rect 427 328 428 329 
<< m1 >>
rect 428 328 429 329 
<< m1 >>
rect 429 328 430 329 
<< m1 >>
rect 430 328 431 329 
<< m1 >>
rect 431 328 432 329 
<< m2 >>
rect 431 328 432 329 
<< m1 >>
rect 432 328 433 329 
<< m1 >>
rect 433 328 434 329 
<< m2 >>
rect 433 328 434 329 
<< m1 >>
rect 434 328 435 329 
<< m1 >>
rect 435 328 436 329 
<< m2 >>
rect 435 328 436 329 
<< m1 >>
rect 436 328 437 329 
<< m1 >>
rect 437 328 438 329 
<< m2 >>
rect 437 328 438 329 
<< m1 >>
rect 438 328 439 329 
<< m1 >>
rect 439 328 440 329 
<< m2 >>
rect 439 328 440 329 
<< m1 >>
rect 440 328 441 329 
<< m1 >>
rect 441 328 442 329 
<< m1 >>
rect 442 328 443 329 
<< m1 >>
rect 443 328 444 329 
<< m1 >>
rect 444 328 445 329 
<< m2 >>
rect 444 328 445 329 
<< m1 >>
rect 445 328 446 329 
<< m2 >>
rect 445 328 446 329 
<< m1 >>
rect 446 328 447 329 
<< m2 >>
rect 446 328 447 329 
<< m1 >>
rect 447 328 448 329 
<< m2 >>
rect 447 328 448 329 
<< m1 >>
rect 448 328 449 329 
<< m2 >>
rect 448 328 449 329 
<< m1 >>
rect 449 328 450 329 
<< m2 >>
rect 449 328 450 329 
<< m1 >>
rect 450 328 451 329 
<< m2 >>
rect 450 328 451 329 
<< m1 >>
rect 451 328 452 329 
<< m2 >>
rect 451 328 452 329 
<< m1 >>
rect 452 328 453 329 
<< m2 >>
rect 452 328 453 329 
<< m1 >>
rect 453 328 454 329 
<< m2 >>
rect 453 328 454 329 
<< m1 >>
rect 454 328 455 329 
<< m2 >>
rect 454 328 455 329 
<< m1 >>
rect 455 328 456 329 
<< m2 >>
rect 455 328 456 329 
<< m1 >>
rect 456 328 457 329 
<< m2 >>
rect 456 328 457 329 
<< m1 >>
rect 457 328 458 329 
<< m2 >>
rect 457 328 458 329 
<< m1 >>
rect 458 328 459 329 
<< m2 >>
rect 458 328 459 329 
<< m1 >>
rect 459 328 460 329 
<< m2 >>
rect 459 328 460 329 
<< m1 >>
rect 460 328 461 329 
<< m2 >>
rect 460 328 461 329 
<< m1 >>
rect 461 328 462 329 
<< m2 >>
rect 461 328 462 329 
<< m1 >>
rect 462 328 463 329 
<< m2 >>
rect 462 328 463 329 
<< m1 >>
rect 463 328 464 329 
<< m2 >>
rect 463 328 464 329 
<< m1 >>
rect 464 328 465 329 
<< m2 >>
rect 464 328 465 329 
<< m1 >>
rect 465 328 466 329 
<< m2 >>
rect 465 328 466 329 
<< m1 >>
rect 466 328 467 329 
<< m2 >>
rect 466 328 467 329 
<< m1 >>
rect 467 328 468 329 
<< m2 >>
rect 467 328 468 329 
<< m1 >>
rect 468 328 469 329 
<< m2 >>
rect 468 328 469 329 
<< m1 >>
rect 469 328 470 329 
<< m2 >>
rect 469 328 470 329 
<< m1 >>
rect 470 328 471 329 
<< m2 >>
rect 470 328 471 329 
<< m1 >>
rect 471 328 472 329 
<< m2 >>
rect 471 328 472 329 
<< m1 >>
rect 472 328 473 329 
<< m2 >>
rect 472 328 473 329 
<< m1 >>
rect 473 328 474 329 
<< m2 >>
rect 473 328 474 329 
<< m1 >>
rect 474 328 475 329 
<< m2 >>
rect 474 328 475 329 
<< m1 >>
rect 475 328 476 329 
<< m2 >>
rect 475 328 476 329 
<< m1 >>
rect 476 328 477 329 
<< m2 >>
rect 476 328 477 329 
<< m1 >>
rect 477 328 478 329 
<< m2 >>
rect 477 328 478 329 
<< m1 >>
rect 478 328 479 329 
<< m2 >>
rect 478 328 479 329 
<< m1 >>
rect 479 328 480 329 
<< m2 >>
rect 479 328 480 329 
<< m1 >>
rect 480 328 481 329 
<< m2 >>
rect 480 328 481 329 
<< m1 >>
rect 481 328 482 329 
<< m2 >>
rect 481 328 482 329 
<< m1 >>
rect 482 328 483 329 
<< m2 >>
rect 482 328 483 329 
<< m1 >>
rect 483 328 484 329 
<< m2 >>
rect 483 328 484 329 
<< m1 >>
rect 484 328 485 329 
<< m2 >>
rect 484 328 485 329 
<< m2 >>
rect 485 328 486 329 
<< m1 >>
rect 523 328 524 329 
<< m1 >>
rect 19 329 20 330 
<< m1 >>
rect 23 329 24 330 
<< m1 >>
rect 25 329 26 330 
<< m1 >>
rect 26 329 27 330 
<< m1 >>
rect 27 329 28 330 
<< m1 >>
rect 28 329 29 330 
<< m1 >>
rect 29 329 30 330 
<< m1 >>
rect 30 329 31 330 
<< m1 >>
rect 31 329 32 330 
<< m1 >>
rect 32 329 33 330 
<< m1 >>
rect 33 329 34 330 
<< m1 >>
rect 34 329 35 330 
<< m1 >>
rect 35 329 36 330 
<< m1 >>
rect 36 329 37 330 
<< m1 >>
rect 37 329 38 330 
<< m1 >>
rect 38 329 39 330 
<< m1 >>
rect 39 329 40 330 
<< m1 >>
rect 40 329 41 330 
<< m1 >>
rect 41 329 42 330 
<< m1 >>
rect 42 329 43 330 
<< m2 >>
rect 42 329 43 330 
<< m2c >>
rect 42 329 43 330 
<< m1 >>
rect 42 329 43 330 
<< m2 >>
rect 42 329 43 330 
<< m2 >>
rect 43 329 44 330 
<< m1 >>
rect 44 329 45 330 
<< m2 >>
rect 44 329 45 330 
<< m2 >>
rect 45 329 46 330 
<< m1 >>
rect 46 329 47 330 
<< m2 >>
rect 46 329 47 330 
<< m2c >>
rect 46 329 47 330 
<< m1 >>
rect 46 329 47 330 
<< m2 >>
rect 46 329 47 330 
<< m1 >>
rect 47 329 48 330 
<< m1 >>
rect 48 329 49 330 
<< m1 >>
rect 49 329 50 330 
<< m1 >>
rect 50 329 51 330 
<< m2 >>
rect 67 329 68 330 
<< m1 >>
rect 73 329 74 330 
<< m2 >>
rect 74 329 75 330 
<< m1 >>
rect 88 329 89 330 
<< m2 >>
rect 91 329 92 330 
<< m1 >>
rect 100 329 101 330 
<< m2 >>
rect 125 329 126 330 
<< m1 >>
rect 146 329 147 330 
<< m1 >>
rect 150 329 151 330 
<< m1 >>
rect 154 329 155 330 
<< m1 >>
rect 159 329 160 330 
<< m2 >>
rect 159 329 160 330 
<< m2c >>
rect 159 329 160 330 
<< m1 >>
rect 159 329 160 330 
<< m2 >>
rect 159 329 160 330 
<< m2 >>
rect 207 329 208 330 
<< m1 >>
rect 215 329 216 330 
<< m1 >>
rect 217 329 218 330 
<< m1 >>
rect 219 329 220 330 
<< m2 >>
rect 221 329 222 330 
<< m2 >>
rect 223 329 224 330 
<< m2 >>
rect 225 329 226 330 
<< m2 >>
rect 235 329 236 330 
<< m2 >>
rect 243 329 244 330 
<< m2 >>
rect 249 329 250 330 
<< m2 >>
rect 253 329 254 330 
<< m2 >>
rect 254 329 255 330 
<< m2 >>
rect 255 329 256 330 
<< m2 >>
rect 256 329 257 330 
<< m2 >>
rect 257 329 258 330 
<< m2 >>
rect 258 329 259 330 
<< m2 >>
rect 259 329 260 330 
<< m2 >>
rect 260 329 261 330 
<< m2 >>
rect 261 329 262 330 
<< m2 >>
rect 262 329 263 330 
<< m2 >>
rect 263 329 264 330 
<< m2 >>
rect 264 329 265 330 
<< m2 >>
rect 265 329 266 330 
<< m2 >>
rect 266 329 267 330 
<< m2 >>
rect 267 329 268 330 
<< m2 >>
rect 268 329 269 330 
<< m2 >>
rect 269 329 270 330 
<< m2 >>
rect 270 329 271 330 
<< m2 >>
rect 271 329 272 330 
<< m2 >>
rect 276 329 277 330 
<< m2 >>
rect 280 329 281 330 
<< m2 >>
rect 281 329 282 330 
<< m2 >>
rect 282 329 283 330 
<< m2 >>
rect 283 329 284 330 
<< m2 >>
rect 284 329 285 330 
<< m2 >>
rect 285 329 286 330 
<< m2 >>
rect 286 329 287 330 
<< m2 >>
rect 289 329 290 330 
<< m2 >>
rect 307 329 308 330 
<< m2 >>
rect 334 329 335 330 
<< m2 >>
rect 343 329 344 330 
<< m1 >>
rect 344 329 345 330 
<< m1 >>
rect 347 329 348 330 
<< m2 >>
rect 351 329 352 330 
<< m2 >>
rect 364 329 365 330 
<< m2 >>
rect 366 329 367 330 
<< m2 >>
rect 370 329 371 330 
<< m2 >>
rect 372 329 373 330 
<< m2 >>
rect 416 329 417 330 
<< m2 >>
rect 418 329 419 330 
<< m2 >>
rect 422 329 423 330 
<< m2 >>
rect 424 329 425 330 
<< m2 >>
rect 431 329 432 330 
<< m2 >>
rect 433 329 434 330 
<< m2 >>
rect 435 329 436 330 
<< m2 >>
rect 437 329 438 330 
<< m2 >>
rect 439 329 440 330 
<< m2 >>
rect 444 329 445 330 
<< m1 >>
rect 523 329 524 330 
<< m1 >>
rect 19 330 20 331 
<< m1 >>
rect 23 330 24 331 
<< m1 >>
rect 44 330 45 331 
<< m1 >>
rect 50 330 51 331 
<< m1 >>
rect 62 330 63 331 
<< m2 >>
rect 62 330 63 331 
<< m2c >>
rect 62 330 63 331 
<< m1 >>
rect 62 330 63 331 
<< m2 >>
rect 62 330 63 331 
<< m2 >>
rect 63 330 64 331 
<< m1 >>
rect 64 330 65 331 
<< m2 >>
rect 64 330 65 331 
<< m1 >>
rect 65 330 66 331 
<< m2 >>
rect 65 330 66 331 
<< m1 >>
rect 66 330 67 331 
<< m2 >>
rect 66 330 67 331 
<< m1 >>
rect 67 330 68 331 
<< m2 >>
rect 67 330 68 331 
<< m1 >>
rect 68 330 69 331 
<< m1 >>
rect 69 330 70 331 
<< m1 >>
rect 70 330 71 331 
<< m1 >>
rect 71 330 72 331 
<< m2 >>
rect 71 330 72 331 
<< m2c >>
rect 71 330 72 331 
<< m1 >>
rect 71 330 72 331 
<< m2 >>
rect 71 330 72 331 
<< m2 >>
rect 72 330 73 331 
<< m1 >>
rect 73 330 74 331 
<< m2 >>
rect 73 330 74 331 
<< m2 >>
rect 74 330 75 331 
<< m1 >>
rect 88 330 89 331 
<< m1 >>
rect 91 330 92 331 
<< m2 >>
rect 91 330 92 331 
<< m2c >>
rect 91 330 92 331 
<< m1 >>
rect 91 330 92 331 
<< m2 >>
rect 91 330 92 331 
<< m1 >>
rect 100 330 101 331 
<< m1 >>
rect 116 330 117 331 
<< m2 >>
rect 116 330 117 331 
<< m2c >>
rect 116 330 117 331 
<< m1 >>
rect 116 330 117 331 
<< m2 >>
rect 116 330 117 331 
<< m2 >>
rect 117 330 118 331 
<< m2 >>
rect 118 330 119 331 
<< m2 >>
rect 119 330 120 331 
<< m2 >>
rect 120 330 121 331 
<< m2 >>
rect 121 330 122 331 
<< m2 >>
rect 122 330 123 331 
<< m2 >>
rect 123 330 124 331 
<< m2 >>
rect 124 330 125 331 
<< m2 >>
rect 125 330 126 331 
<< m1 >>
rect 146 330 147 331 
<< m1 >>
rect 150 330 151 331 
<< m1 >>
rect 154 330 155 331 
<< m2 >>
rect 159 330 160 331 
<< m2 >>
rect 207 330 208 331 
<< m2 >>
rect 210 330 211 331 
<< m2 >>
rect 211 330 212 331 
<< m2 >>
rect 212 330 213 331 
<< m1 >>
rect 213 330 214 331 
<< m2 >>
rect 213 330 214 331 
<< m2c >>
rect 213 330 214 331 
<< m1 >>
rect 213 330 214 331 
<< m2 >>
rect 213 330 214 331 
<< m1 >>
rect 214 330 215 331 
<< m1 >>
rect 215 330 216 331 
<< m1 >>
rect 217 330 218 331 
<< m1 >>
rect 219 330 220 331 
<< m1 >>
rect 220 330 221 331 
<< m1 >>
rect 221 330 222 331 
<< m2 >>
rect 221 330 222 331 
<< m1 >>
rect 222 330 223 331 
<< m1 >>
rect 223 330 224 331 
<< m2 >>
rect 223 330 224 331 
<< m1 >>
rect 224 330 225 331 
<< m1 >>
rect 225 330 226 331 
<< m2 >>
rect 225 330 226 331 
<< m1 >>
rect 226 330 227 331 
<< m1 >>
rect 227 330 228 331 
<< m1 >>
rect 228 330 229 331 
<< m1 >>
rect 229 330 230 331 
<< m1 >>
rect 230 330 231 331 
<< m1 >>
rect 231 330 232 331 
<< m1 >>
rect 232 330 233 331 
<< m1 >>
rect 233 330 234 331 
<< m1 >>
rect 234 330 235 331 
<< m1 >>
rect 235 330 236 331 
<< m2 >>
rect 235 330 236 331 
<< m1 >>
rect 236 330 237 331 
<< m1 >>
rect 237 330 238 331 
<< m1 >>
rect 238 330 239 331 
<< m1 >>
rect 239 330 240 331 
<< m1 >>
rect 240 330 241 331 
<< m1 >>
rect 241 330 242 331 
<< m1 >>
rect 242 330 243 331 
<< m2 >>
rect 242 330 243 331 
<< m1 >>
rect 243 330 244 331 
<< m2 >>
rect 243 330 244 331 
<< m1 >>
rect 244 330 245 331 
<< m1 >>
rect 245 330 246 331 
<< m1 >>
rect 246 330 247 331 
<< m1 >>
rect 247 330 248 331 
<< m1 >>
rect 248 330 249 331 
<< m2 >>
rect 249 330 250 331 
<< m1 >>
rect 253 330 254 331 
<< m2 >>
rect 253 330 254 331 
<< m2c >>
rect 253 330 254 331 
<< m1 >>
rect 253 330 254 331 
<< m2 >>
rect 253 330 254 331 
<< m1 >>
rect 276 330 277 331 
<< m2 >>
rect 276 330 277 331 
<< m2c >>
rect 276 330 277 331 
<< m1 >>
rect 276 330 277 331 
<< m2 >>
rect 276 330 277 331 
<< m1 >>
rect 286 330 287 331 
<< m2 >>
rect 286 330 287 331 
<< m2c >>
rect 286 330 287 331 
<< m1 >>
rect 286 330 287 331 
<< m2 >>
rect 286 330 287 331 
<< m1 >>
rect 289 330 290 331 
<< m2 >>
rect 289 330 290 331 
<< m2c >>
rect 289 330 290 331 
<< m1 >>
rect 289 330 290 331 
<< m2 >>
rect 289 330 290 331 
<< m1 >>
rect 307 330 308 331 
<< m2 >>
rect 307 330 308 331 
<< m2c >>
rect 307 330 308 331 
<< m1 >>
rect 307 330 308 331 
<< m2 >>
rect 307 330 308 331 
<< m1 >>
rect 308 330 309 331 
<< m1 >>
rect 309 330 310 331 
<< m1 >>
rect 310 330 311 331 
<< m1 >>
rect 311 330 312 331 
<< m1 >>
rect 312 330 313 331 
<< m1 >>
rect 313 330 314 331 
<< m1 >>
rect 314 330 315 331 
<< m1 >>
rect 315 330 316 331 
<< m1 >>
rect 316 330 317 331 
<< m1 >>
rect 317 330 318 331 
<< m1 >>
rect 318 330 319 331 
<< m1 >>
rect 319 330 320 331 
<< m1 >>
rect 320 330 321 331 
<< m1 >>
rect 334 330 335 331 
<< m2 >>
rect 334 330 335 331 
<< m2c >>
rect 334 330 335 331 
<< m1 >>
rect 334 330 335 331 
<< m2 >>
rect 334 330 335 331 
<< m2 >>
rect 343 330 344 331 
<< m1 >>
rect 344 330 345 331 
<< m1 >>
rect 347 330 348 331 
<< m2 >>
rect 347 330 348 331 
<< m2c >>
rect 347 330 348 331 
<< m1 >>
rect 347 330 348 331 
<< m2 >>
rect 347 330 348 331 
<< m1 >>
rect 351 330 352 331 
<< m2 >>
rect 351 330 352 331 
<< m2c >>
rect 351 330 352 331 
<< m1 >>
rect 351 330 352 331 
<< m2 >>
rect 351 330 352 331 
<< m1 >>
rect 364 330 365 331 
<< m2 >>
rect 364 330 365 331 
<< m2c >>
rect 364 330 365 331 
<< m1 >>
rect 364 330 365 331 
<< m2 >>
rect 364 330 365 331 
<< m1 >>
rect 366 330 367 331 
<< m2 >>
rect 366 330 367 331 
<< m2c >>
rect 366 330 367 331 
<< m1 >>
rect 366 330 367 331 
<< m2 >>
rect 366 330 367 331 
<< m1 >>
rect 370 330 371 331 
<< m2 >>
rect 370 330 371 331 
<< m2c >>
rect 370 330 371 331 
<< m1 >>
rect 370 330 371 331 
<< m2 >>
rect 370 330 371 331 
<< m1 >>
rect 372 330 373 331 
<< m2 >>
rect 372 330 373 331 
<< m2c >>
rect 372 330 373 331 
<< m1 >>
rect 372 330 373 331 
<< m2 >>
rect 372 330 373 331 
<< m1 >>
rect 416 330 417 331 
<< m2 >>
rect 416 330 417 331 
<< m2c >>
rect 416 330 417 331 
<< m1 >>
rect 416 330 417 331 
<< m2 >>
rect 416 330 417 331 
<< m1 >>
rect 418 330 419 331 
<< m2 >>
rect 418 330 419 331 
<< m2c >>
rect 418 330 419 331 
<< m1 >>
rect 418 330 419 331 
<< m2 >>
rect 418 330 419 331 
<< m1 >>
rect 422 330 423 331 
<< m2 >>
rect 422 330 423 331 
<< m2c >>
rect 422 330 423 331 
<< m1 >>
rect 422 330 423 331 
<< m2 >>
rect 422 330 423 331 
<< m1 >>
rect 424 330 425 331 
<< m2 >>
rect 424 330 425 331 
<< m2c >>
rect 424 330 425 331 
<< m1 >>
rect 424 330 425 331 
<< m2 >>
rect 424 330 425 331 
<< m1 >>
rect 431 330 432 331 
<< m2 >>
rect 431 330 432 331 
<< m2c >>
rect 431 330 432 331 
<< m1 >>
rect 431 330 432 331 
<< m2 >>
rect 431 330 432 331 
<< m1 >>
rect 433 330 434 331 
<< m2 >>
rect 433 330 434 331 
<< m2c >>
rect 433 330 434 331 
<< m1 >>
rect 433 330 434 331 
<< m2 >>
rect 433 330 434 331 
<< m1 >>
rect 435 330 436 331 
<< m2 >>
rect 435 330 436 331 
<< m2c >>
rect 435 330 436 331 
<< m1 >>
rect 435 330 436 331 
<< m2 >>
rect 435 330 436 331 
<< m1 >>
rect 437 330 438 331 
<< m2 >>
rect 437 330 438 331 
<< m2c >>
rect 437 330 438 331 
<< m1 >>
rect 437 330 438 331 
<< m2 >>
rect 437 330 438 331 
<< m1 >>
rect 438 330 439 331 
<< m1 >>
rect 439 330 440 331 
<< m2 >>
rect 439 330 440 331 
<< m1 >>
rect 440 330 441 331 
<< m1 >>
rect 441 330 442 331 
<< m1 >>
rect 442 330 443 331 
<< m1 >>
rect 443 330 444 331 
<< m1 >>
rect 444 330 445 331 
<< m2 >>
rect 444 330 445 331 
<< m1 >>
rect 445 330 446 331 
<< m1 >>
rect 446 330 447 331 
<< m1 >>
rect 447 330 448 331 
<< m1 >>
rect 448 330 449 331 
<< m1 >>
rect 449 330 450 331 
<< m1 >>
rect 450 330 451 331 
<< m1 >>
rect 451 330 452 331 
<< m1 >>
rect 523 330 524 331 
<< m1 >>
rect 19 331 20 332 
<< m1 >>
rect 23 331 24 332 
<< m1 >>
rect 44 331 45 332 
<< m1 >>
rect 50 331 51 332 
<< m1 >>
rect 62 331 63 332 
<< m1 >>
rect 64 331 65 332 
<< m1 >>
rect 73 331 74 332 
<< m1 >>
rect 88 331 89 332 
<< m1 >>
rect 91 331 92 332 
<< m1 >>
rect 100 331 101 332 
<< m1 >>
rect 116 331 117 332 
<< m1 >>
rect 118 331 119 332 
<< m1 >>
rect 119 331 120 332 
<< m1 >>
rect 120 331 121 332 
<< m1 >>
rect 121 331 122 332 
<< m1 >>
rect 122 331 123 332 
<< m1 >>
rect 123 331 124 332 
<< m1 >>
rect 124 331 125 332 
<< m1 >>
rect 146 331 147 332 
<< m1 >>
rect 148 331 149 332 
<< m2 >>
rect 148 331 149 332 
<< m2c >>
rect 148 331 149 332 
<< m1 >>
rect 148 331 149 332 
<< m2 >>
rect 148 331 149 332 
<< m2 >>
rect 149 331 150 332 
<< m1 >>
rect 150 331 151 332 
<< m2 >>
rect 150 331 151 332 
<< m2 >>
rect 151 331 152 332 
<< m1 >>
rect 152 331 153 332 
<< m2 >>
rect 152 331 153 332 
<< m2c >>
rect 152 331 153 332 
<< m1 >>
rect 152 331 153 332 
<< m2 >>
rect 152 331 153 332 
<< m2 >>
rect 153 331 154 332 
<< m1 >>
rect 154 331 155 332 
<< m2 >>
rect 154 331 155 332 
<< m2 >>
rect 155 331 156 332 
<< m1 >>
rect 156 331 157 332 
<< m2 >>
rect 156 331 157 332 
<< m2c >>
rect 156 331 157 332 
<< m1 >>
rect 156 331 157 332 
<< m2 >>
rect 156 331 157 332 
<< m1 >>
rect 157 331 158 332 
<< m1 >>
rect 158 331 159 332 
<< m1 >>
rect 159 331 160 332 
<< m2 >>
rect 159 331 160 332 
<< m1 >>
rect 160 331 161 332 
<< m1 >>
rect 161 331 162 332 
<< m2 >>
rect 161 331 162 332 
<< m2c >>
rect 161 331 162 332 
<< m1 >>
rect 161 331 162 332 
<< m2 >>
rect 161 331 162 332 
<< m2 >>
rect 162 331 163 332 
<< m1 >>
rect 163 331 164 332 
<< m2 >>
rect 163 331 164 332 
<< m1 >>
rect 164 331 165 332 
<< m2 >>
rect 164 331 165 332 
<< m1 >>
rect 165 331 166 332 
<< m2 >>
rect 165 331 166 332 
<< m1 >>
rect 166 331 167 332 
<< m2 >>
rect 166 331 167 332 
<< m1 >>
rect 167 331 168 332 
<< m2 >>
rect 167 331 168 332 
<< m1 >>
rect 168 331 169 332 
<< m2 >>
rect 168 331 169 332 
<< m1 >>
rect 169 331 170 332 
<< m2 >>
rect 169 331 170 332 
<< m1 >>
rect 170 331 171 332 
<< m2 >>
rect 170 331 171 332 
<< m1 >>
rect 171 331 172 332 
<< m2 >>
rect 171 331 172 332 
<< m1 >>
rect 172 331 173 332 
<< m2 >>
rect 172 331 173 332 
<< m1 >>
rect 173 331 174 332 
<< m2 >>
rect 173 331 174 332 
<< m1 >>
rect 174 331 175 332 
<< m2 >>
rect 174 331 175 332 
<< m1 >>
rect 175 331 176 332 
<< m2 >>
rect 175 331 176 332 
<< m1 >>
rect 176 331 177 332 
<< m2 >>
rect 176 331 177 332 
<< m1 >>
rect 177 331 178 332 
<< m2 >>
rect 177 331 178 332 
<< m1 >>
rect 178 331 179 332 
<< m2 >>
rect 178 331 179 332 
<< m1 >>
rect 179 331 180 332 
<< m1 >>
rect 180 331 181 332 
<< m1 >>
rect 181 331 182 332 
<< m2 >>
rect 181 331 182 332 
<< m1 >>
rect 182 331 183 332 
<< m2 >>
rect 182 331 183 332 
<< m1 >>
rect 183 331 184 332 
<< m2 >>
rect 183 331 184 332 
<< m1 >>
rect 184 331 185 332 
<< m2 >>
rect 184 331 185 332 
<< m1 >>
rect 185 331 186 332 
<< m2 >>
rect 185 331 186 332 
<< m1 >>
rect 186 331 187 332 
<< m2 >>
rect 186 331 187 332 
<< m1 >>
rect 187 331 188 332 
<< m2 >>
rect 187 331 188 332 
<< m1 >>
rect 188 331 189 332 
<< m2 >>
rect 188 331 189 332 
<< m1 >>
rect 189 331 190 332 
<< m2 >>
rect 189 331 190 332 
<< m1 >>
rect 190 331 191 332 
<< m2 >>
rect 190 331 191 332 
<< m1 >>
rect 191 331 192 332 
<< m2 >>
rect 191 331 192 332 
<< m1 >>
rect 192 331 193 332 
<< m2 >>
rect 192 331 193 332 
<< m1 >>
rect 193 331 194 332 
<< m2 >>
rect 193 331 194 332 
<< m1 >>
rect 194 331 195 332 
<< m2 >>
rect 194 331 195 332 
<< m1 >>
rect 195 331 196 332 
<< m2 >>
rect 195 331 196 332 
<< m1 >>
rect 196 331 197 332 
<< m2 >>
rect 196 331 197 332 
<< m2 >>
rect 197 331 198 332 
<< m1 >>
rect 198 331 199 332 
<< m2 >>
rect 198 331 199 332 
<< m2c >>
rect 198 331 199 332 
<< m1 >>
rect 198 331 199 332 
<< m2 >>
rect 198 331 199 332 
<< m1 >>
rect 199 331 200 332 
<< m1 >>
rect 200 331 201 332 
<< m1 >>
rect 201 331 202 332 
<< m1 >>
rect 202 331 203 332 
<< m1 >>
rect 203 331 204 332 
<< m1 >>
rect 204 331 205 332 
<< m1 >>
rect 205 331 206 332 
<< m1 >>
rect 206 331 207 332 
<< m1 >>
rect 207 331 208 332 
<< m2 >>
rect 207 331 208 332 
<< m1 >>
rect 208 331 209 332 
<< m1 >>
rect 209 331 210 332 
<< m1 >>
rect 210 331 211 332 
<< m2 >>
rect 210 331 211 332 
<< m1 >>
rect 211 331 212 332 
<< m1 >>
rect 217 331 218 332 
<< m2 >>
rect 219 331 220 332 
<< m2 >>
rect 220 331 221 332 
<< m2 >>
rect 221 331 222 332 
<< m2 >>
rect 223 331 224 332 
<< m2 >>
rect 225 331 226 332 
<< m2 >>
rect 235 331 236 332 
<< m2 >>
rect 242 331 243 332 
<< m2 >>
rect 244 331 245 332 
<< m2 >>
rect 245 331 246 332 
<< m2 >>
rect 246 331 247 332 
<< m2 >>
rect 247 331 248 332 
<< m1 >>
rect 248 331 249 332 
<< m2 >>
rect 248 331 249 332 
<< m2 >>
rect 249 331 250 332 
<< m1 >>
rect 253 331 254 332 
<< m1 >>
rect 255 331 256 332 
<< m1 >>
rect 256 331 257 332 
<< m1 >>
rect 257 331 258 332 
<< m1 >>
rect 258 331 259 332 
<< m1 >>
rect 259 331 260 332 
<< m1 >>
rect 260 331 261 332 
<< m1 >>
rect 261 331 262 332 
<< m1 >>
rect 262 331 263 332 
<< m1 >>
rect 263 331 264 332 
<< m1 >>
rect 264 331 265 332 
<< m1 >>
rect 265 331 266 332 
<< m1 >>
rect 266 331 267 332 
<< m1 >>
rect 267 331 268 332 
<< m1 >>
rect 268 331 269 332 
<< m1 >>
rect 276 331 277 332 
<< m1 >>
rect 286 331 287 332 
<< m1 >>
rect 289 331 290 332 
<< m1 >>
rect 320 331 321 332 
<< m1 >>
rect 334 331 335 332 
<< m1 >>
rect 336 331 337 332 
<< m1 >>
rect 337 331 338 332 
<< m1 >>
rect 338 331 339 332 
<< m1 >>
rect 339 331 340 332 
<< m1 >>
rect 340 331 341 332 
<< m1 >>
rect 341 331 342 332 
<< m1 >>
rect 342 331 343 332 
<< m2 >>
rect 342 331 343 332 
<< m2c >>
rect 342 331 343 332 
<< m1 >>
rect 342 331 343 332 
<< m2 >>
rect 342 331 343 332 
<< m2 >>
rect 343 331 344 332 
<< m1 >>
rect 344 331 345 332 
<< m2 >>
rect 347 331 348 332 
<< m1 >>
rect 351 331 352 332 
<< m1 >>
rect 353 331 354 332 
<< m1 >>
rect 354 331 355 332 
<< m1 >>
rect 355 331 356 332 
<< m1 >>
rect 356 331 357 332 
<< m1 >>
rect 357 331 358 332 
<< m1 >>
rect 358 331 359 332 
<< m1 >>
rect 359 331 360 332 
<< m1 >>
rect 360 331 361 332 
<< m1 >>
rect 361 331 362 332 
<< m1 >>
rect 364 331 365 332 
<< m1 >>
rect 366 331 367 332 
<< m1 >>
rect 370 331 371 332 
<< m1 >>
rect 372 331 373 332 
<< m1 >>
rect 416 331 417 332 
<< m1 >>
rect 418 331 419 332 
<< m1 >>
rect 422 331 423 332 
<< m1 >>
rect 424 331 425 332 
<< m1 >>
rect 431 331 432 332 
<< m1 >>
rect 433 331 434 332 
<< m1 >>
rect 435 331 436 332 
<< m2 >>
rect 439 331 440 332 
<< m2 >>
rect 444 331 445 332 
<< m1 >>
rect 451 331 452 332 
<< m1 >>
rect 523 331 524 332 
<< m1 >>
rect 19 332 20 333 
<< m1 >>
rect 23 332 24 333 
<< m2 >>
rect 23 332 24 333 
<< m2c >>
rect 23 332 24 333 
<< m1 >>
rect 23 332 24 333 
<< m2 >>
rect 23 332 24 333 
<< m1 >>
rect 44 332 45 333 
<< m1 >>
rect 50 332 51 333 
<< m1 >>
rect 51 332 52 333 
<< m1 >>
rect 52 332 53 333 
<< m1 >>
rect 53 332 54 333 
<< m1 >>
rect 54 332 55 333 
<< m1 >>
rect 55 332 56 333 
<< m1 >>
rect 56 332 57 333 
<< m1 >>
rect 57 332 58 333 
<< m1 >>
rect 58 332 59 333 
<< m1 >>
rect 59 332 60 333 
<< m1 >>
rect 60 332 61 333 
<< m2 >>
rect 60 332 61 333 
<< m2c >>
rect 60 332 61 333 
<< m1 >>
rect 60 332 61 333 
<< m2 >>
rect 60 332 61 333 
<< m2 >>
rect 61 332 62 333 
<< m1 >>
rect 62 332 63 333 
<< m1 >>
rect 64 332 65 333 
<< m1 >>
rect 73 332 74 333 
<< m1 >>
rect 88 332 89 333 
<< m1 >>
rect 91 332 92 333 
<< m1 >>
rect 100 332 101 333 
<< m1 >>
rect 116 332 117 333 
<< m1 >>
rect 118 332 119 333 
<< m1 >>
rect 124 332 125 333 
<< m1 >>
rect 146 332 147 333 
<< m2 >>
rect 146 332 147 333 
<< m2c >>
rect 146 332 147 333 
<< m1 >>
rect 146 332 147 333 
<< m2 >>
rect 146 332 147 333 
<< m1 >>
rect 148 332 149 333 
<< m1 >>
rect 150 332 151 333 
<< m1 >>
rect 154 332 155 333 
<< m2 >>
rect 159 332 160 333 
<< m1 >>
rect 163 332 164 333 
<< m2 >>
rect 178 332 179 333 
<< m2 >>
rect 181 332 182 333 
<< m1 >>
rect 196 332 197 333 
<< m2 >>
rect 207 332 208 333 
<< m2 >>
rect 210 332 211 333 
<< m1 >>
rect 211 332 212 333 
<< m1 >>
rect 217 332 218 333 
<< m1 >>
rect 219 332 220 333 
<< m2 >>
rect 219 332 220 333 
<< m2c >>
rect 219 332 220 333 
<< m1 >>
rect 219 332 220 333 
<< m2 >>
rect 219 332 220 333 
<< m1 >>
rect 223 332 224 333 
<< m2 >>
rect 223 332 224 333 
<< m2c >>
rect 223 332 224 333 
<< m1 >>
rect 223 332 224 333 
<< m2 >>
rect 223 332 224 333 
<< m1 >>
rect 225 332 226 333 
<< m2 >>
rect 225 332 226 333 
<< m2c >>
rect 225 332 226 333 
<< m1 >>
rect 225 332 226 333 
<< m2 >>
rect 225 332 226 333 
<< m1 >>
rect 235 332 236 333 
<< m2 >>
rect 235 332 236 333 
<< m2c >>
rect 235 332 236 333 
<< m1 >>
rect 235 332 236 333 
<< m2 >>
rect 235 332 236 333 
<< m1 >>
rect 242 332 243 333 
<< m2 >>
rect 242 332 243 333 
<< m2c >>
rect 242 332 243 333 
<< m1 >>
rect 242 332 243 333 
<< m2 >>
rect 242 332 243 333 
<< m1 >>
rect 244 332 245 333 
<< m2 >>
rect 244 332 245 333 
<< m2c >>
rect 244 332 245 333 
<< m1 >>
rect 244 332 245 333 
<< m2 >>
rect 244 332 245 333 
<< m1 >>
rect 248 332 249 333 
<< m1 >>
rect 249 332 250 333 
<< m1 >>
rect 250 332 251 333 
<< m1 >>
rect 251 332 252 333 
<< m2 >>
rect 251 332 252 333 
<< m2c >>
rect 251 332 252 333 
<< m1 >>
rect 251 332 252 333 
<< m2 >>
rect 251 332 252 333 
<< m2 >>
rect 252 332 253 333 
<< m1 >>
rect 253 332 254 333 
<< m2 >>
rect 253 332 254 333 
<< m2 >>
rect 254 332 255 333 
<< m1 >>
rect 255 332 256 333 
<< m2 >>
rect 255 332 256 333 
<< m2c >>
rect 255 332 256 333 
<< m1 >>
rect 255 332 256 333 
<< m2 >>
rect 255 332 256 333 
<< m1 >>
rect 268 332 269 333 
<< m1 >>
rect 276 332 277 333 
<< m1 >>
rect 286 332 287 333 
<< m1 >>
rect 289 332 290 333 
<< m1 >>
rect 320 332 321 333 
<< m1 >>
rect 321 332 322 333 
<< m1 >>
rect 322 332 323 333 
<< m1 >>
rect 323 332 324 333 
<< m1 >>
rect 324 332 325 333 
<< m1 >>
rect 325 332 326 333 
<< m1 >>
rect 326 332 327 333 
<< m1 >>
rect 327 332 328 333 
<< m1 >>
rect 328 332 329 333 
<< m1 >>
rect 329 332 330 333 
<< m1 >>
rect 330 332 331 333 
<< m1 >>
rect 331 332 332 333 
<< m1 >>
rect 332 332 333 333 
<< m2 >>
rect 332 332 333 333 
<< m2c >>
rect 332 332 333 333 
<< m1 >>
rect 332 332 333 333 
<< m2 >>
rect 332 332 333 333 
<< m2 >>
rect 333 332 334 333 
<< m1 >>
rect 334 332 335 333 
<< m2 >>
rect 334 332 335 333 
<< m2 >>
rect 335 332 336 333 
<< m1 >>
rect 336 332 337 333 
<< m2 >>
rect 336 332 337 333 
<< m2c >>
rect 336 332 337 333 
<< m1 >>
rect 336 332 337 333 
<< m2 >>
rect 336 332 337 333 
<< m1 >>
rect 344 332 345 333 
<< m1 >>
rect 345 332 346 333 
<< m1 >>
rect 346 332 347 333 
<< m1 >>
rect 347 332 348 333 
<< m2 >>
rect 347 332 348 333 
<< m1 >>
rect 348 332 349 333 
<< m1 >>
rect 349 332 350 333 
<< m2 >>
rect 349 332 350 333 
<< m2c >>
rect 349 332 350 333 
<< m1 >>
rect 349 332 350 333 
<< m2 >>
rect 349 332 350 333 
<< m2 >>
rect 350 332 351 333 
<< m1 >>
rect 351 332 352 333 
<< m2 >>
rect 351 332 352 333 
<< m2 >>
rect 352 332 353 333 
<< m1 >>
rect 353 332 354 333 
<< m2 >>
rect 353 332 354 333 
<< m2c >>
rect 353 332 354 333 
<< m1 >>
rect 353 332 354 333 
<< m2 >>
rect 353 332 354 333 
<< m1 >>
rect 361 332 362 333 
<< m1 >>
rect 364 332 365 333 
<< m1 >>
rect 366 332 367 333 
<< m1 >>
rect 367 332 368 333 
<< m1 >>
rect 368 332 369 333 
<< m2 >>
rect 368 332 369 333 
<< m2c >>
rect 368 332 369 333 
<< m1 >>
rect 368 332 369 333 
<< m2 >>
rect 368 332 369 333 
<< m2 >>
rect 369 332 370 333 
<< m1 >>
rect 370 332 371 333 
<< m2 >>
rect 370 332 371 333 
<< m2 >>
rect 371 332 372 333 
<< m1 >>
rect 372 332 373 333 
<< m2 >>
rect 372 332 373 333 
<< m2c >>
rect 372 332 373 333 
<< m1 >>
rect 372 332 373 333 
<< m2 >>
rect 372 332 373 333 
<< m1 >>
rect 416 332 417 333 
<< m1 >>
rect 418 332 419 333 
<< m1 >>
rect 422 332 423 333 
<< m1 >>
rect 424 332 425 333 
<< m1 >>
rect 431 332 432 333 
<< m2 >>
rect 431 332 432 333 
<< m2c >>
rect 431 332 432 333 
<< m1 >>
rect 431 332 432 333 
<< m2 >>
rect 431 332 432 333 
<< m2 >>
rect 432 332 433 333 
<< m1 >>
rect 433 332 434 333 
<< m2 >>
rect 433 332 434 333 
<< m2 >>
rect 434 332 435 333 
<< m1 >>
rect 435 332 436 333 
<< m2 >>
rect 435 332 436 333 
<< m2 >>
rect 436 332 437 333 
<< m1 >>
rect 437 332 438 333 
<< m2 >>
rect 437 332 438 333 
<< m2c >>
rect 437 332 438 333 
<< m1 >>
rect 437 332 438 333 
<< m2 >>
rect 437 332 438 333 
<< m1 >>
rect 438 332 439 333 
<< m1 >>
rect 439 332 440 333 
<< m2 >>
rect 439 332 440 333 
<< m1 >>
rect 440 332 441 333 
<< m1 >>
rect 441 332 442 333 
<< m1 >>
rect 442 332 443 333 
<< m1 >>
rect 443 332 444 333 
<< m1 >>
rect 444 332 445 333 
<< m2 >>
rect 444 332 445 333 
<< m2c >>
rect 444 332 445 333 
<< m1 >>
rect 444 332 445 333 
<< m2 >>
rect 444 332 445 333 
<< m1 >>
rect 451 332 452 333 
<< m1 >>
rect 523 332 524 333 
<< m1 >>
rect 19 333 20 334 
<< m2 >>
rect 23 333 24 334 
<< m1 >>
rect 44 333 45 334 
<< m2 >>
rect 61 333 62 334 
<< m1 >>
rect 62 333 63 334 
<< m1 >>
rect 64 333 65 334 
<< m1 >>
rect 73 333 74 334 
<< m1 >>
rect 88 333 89 334 
<< m1 >>
rect 91 333 92 334 
<< m1 >>
rect 100 333 101 334 
<< m1 >>
rect 116 333 117 334 
<< m1 >>
rect 118 333 119 334 
<< m1 >>
rect 124 333 125 334 
<< m2 >>
rect 146 333 147 334 
<< m1 >>
rect 148 333 149 334 
<< m1 >>
rect 150 333 151 334 
<< m1 >>
rect 154 333 155 334 
<< m1 >>
rect 159 333 160 334 
<< m2 >>
rect 159 333 160 334 
<< m2c >>
rect 159 333 160 334 
<< m1 >>
rect 159 333 160 334 
<< m2 >>
rect 159 333 160 334 
<< m1 >>
rect 160 333 161 334 
<< m1 >>
rect 161 333 162 334 
<< m1 >>
rect 163 333 164 334 
<< m1 >>
rect 178 333 179 334 
<< m2 >>
rect 178 333 179 334 
<< m2c >>
rect 178 333 179 334 
<< m1 >>
rect 178 333 179 334 
<< m2 >>
rect 178 333 179 334 
<< m1 >>
rect 181 333 182 334 
<< m2 >>
rect 181 333 182 334 
<< m2c >>
rect 181 333 182 334 
<< m1 >>
rect 181 333 182 334 
<< m2 >>
rect 181 333 182 334 
<< m1 >>
rect 196 333 197 334 
<< m1 >>
rect 204 333 205 334 
<< m2 >>
rect 204 333 205 334 
<< m2c >>
rect 204 333 205 334 
<< m1 >>
rect 204 333 205 334 
<< m2 >>
rect 204 333 205 334 
<< m2 >>
rect 205 333 206 334 
<< m1 >>
rect 206 333 207 334 
<< m2 >>
rect 206 333 207 334 
<< m1 >>
rect 207 333 208 334 
<< m2 >>
rect 207 333 208 334 
<< m1 >>
rect 208 333 209 334 
<< m1 >>
rect 209 333 210 334 
<< m2 >>
rect 209 333 210 334 
<< m2c >>
rect 209 333 210 334 
<< m1 >>
rect 209 333 210 334 
<< m2 >>
rect 209 333 210 334 
<< m2 >>
rect 210 333 211 334 
<< m1 >>
rect 211 333 212 334 
<< m1 >>
rect 217 333 218 334 
<< m1 >>
rect 219 333 220 334 
<< m1 >>
rect 223 333 224 334 
<< m1 >>
rect 225 333 226 334 
<< m1 >>
rect 235 333 236 334 
<< m1 >>
rect 242 333 243 334 
<< m2 >>
rect 244 333 245 334 
<< m1 >>
rect 253 333 254 334 
<< m1 >>
rect 268 333 269 334 
<< m1 >>
rect 276 333 277 334 
<< m1 >>
rect 286 333 287 334 
<< m1 >>
rect 289 333 290 334 
<< m1 >>
rect 334 333 335 334 
<< m2 >>
rect 347 333 348 334 
<< m1 >>
rect 351 333 352 334 
<< m1 >>
rect 361 333 362 334 
<< m1 >>
rect 364 333 365 334 
<< m1 >>
rect 370 333 371 334 
<< m1 >>
rect 416 333 417 334 
<< m1 >>
rect 418 333 419 334 
<< m1 >>
rect 422 333 423 334 
<< m1 >>
rect 424 333 425 334 
<< m1 >>
rect 433 333 434 334 
<< m1 >>
rect 435 333 436 334 
<< m2 >>
rect 439 333 440 334 
<< m1 >>
rect 451 333 452 334 
<< m1 >>
rect 523 333 524 334 
<< m1 >>
rect 19 334 20 335 
<< m2 >>
rect 20 334 21 335 
<< m1 >>
rect 21 334 22 335 
<< m2 >>
rect 21 334 22 335 
<< m2c >>
rect 21 334 22 335 
<< m1 >>
rect 21 334 22 335 
<< m2 >>
rect 21 334 22 335 
<< m1 >>
rect 22 334 23 335 
<< m1 >>
rect 23 334 24 335 
<< m2 >>
rect 23 334 24 335 
<< m1 >>
rect 24 334 25 335 
<< m1 >>
rect 25 334 26 335 
<< m1 >>
rect 26 334 27 335 
<< m1 >>
rect 27 334 28 335 
<< m1 >>
rect 28 334 29 335 
<< m1 >>
rect 29 334 30 335 
<< m1 >>
rect 30 334 31 335 
<< m1 >>
rect 31 334 32 335 
<< m1 >>
rect 44 334 45 335 
<< m2 >>
rect 61 334 62 335 
<< m1 >>
rect 62 334 63 335 
<< m1 >>
rect 64 334 65 335 
<< m1 >>
rect 73 334 74 335 
<< m1 >>
rect 82 334 83 335 
<< m1 >>
rect 83 334 84 335 
<< m1 >>
rect 84 334 85 335 
<< m1 >>
rect 85 334 86 335 
<< m1 >>
rect 88 334 89 335 
<< m1 >>
rect 91 334 92 335 
<< m1 >>
rect 100 334 101 335 
<< m1 >>
rect 116 334 117 335 
<< m1 >>
rect 118 334 119 335 
<< m1 >>
rect 124 334 125 335 
<< m1 >>
rect 142 334 143 335 
<< m1 >>
rect 143 334 144 335 
<< m1 >>
rect 144 334 145 335 
<< m1 >>
rect 145 334 146 335 
<< m2 >>
rect 146 334 147 335 
<< m1 >>
rect 148 334 149 335 
<< m1 >>
rect 150 334 151 335 
<< m1 >>
rect 154 334 155 335 
<< m1 >>
rect 161 334 162 335 
<< m2 >>
rect 161 334 162 335 
<< m2c >>
rect 161 334 162 335 
<< m1 >>
rect 161 334 162 335 
<< m2 >>
rect 161 334 162 335 
<< m2 >>
rect 162 334 163 335 
<< m1 >>
rect 163 334 164 335 
<< m2 >>
rect 163 334 164 335 
<< m2 >>
rect 164 334 165 335 
<< m1 >>
rect 178 334 179 335 
<< m1 >>
rect 181 334 182 335 
<< m1 >>
rect 196 334 197 335 
<< m1 >>
rect 204 334 205 335 
<< m1 >>
rect 206 334 207 335 
<< m1 >>
rect 211 334 212 335 
<< m1 >>
rect 217 334 218 335 
<< m1 >>
rect 219 334 220 335 
<< m1 >>
rect 223 334 224 335 
<< m1 >>
rect 225 334 226 335 
<< m1 >>
rect 235 334 236 335 
<< m1 >>
rect 242 334 243 335 
<< m1 >>
rect 244 334 245 335 
<< m2 >>
rect 244 334 245 335 
<< m1 >>
rect 245 334 246 335 
<< m1 >>
rect 246 334 247 335 
<< m1 >>
rect 247 334 248 335 
<< m1 >>
rect 253 334 254 335 
<< m1 >>
rect 268 334 269 335 
<< m1 >>
rect 276 334 277 335 
<< m1 >>
rect 286 334 287 335 
<< m1 >>
rect 289 334 290 335 
<< m1 >>
rect 334 334 335 335 
<< m1 >>
rect 347 334 348 335 
<< m2 >>
rect 347 334 348 335 
<< m2c >>
rect 347 334 348 335 
<< m1 >>
rect 347 334 348 335 
<< m2 >>
rect 347 334 348 335 
<< m2 >>
rect 350 334 351 335 
<< m1 >>
rect 351 334 352 335 
<< m2 >>
rect 351 334 352 335 
<< m2 >>
rect 352 334 353 335 
<< m1 >>
rect 353 334 354 335 
<< m2 >>
rect 353 334 354 335 
<< m2c >>
rect 353 334 354 335 
<< m1 >>
rect 353 334 354 335 
<< m2 >>
rect 353 334 354 335 
<< m1 >>
rect 354 334 355 335 
<< m1 >>
rect 355 334 356 335 
<< m1 >>
rect 361 334 362 335 
<< m1 >>
rect 364 334 365 335 
<< m1 >>
rect 370 334 371 335 
<< m1 >>
rect 376 334 377 335 
<< m1 >>
rect 377 334 378 335 
<< m1 >>
rect 378 334 379 335 
<< m1 >>
rect 379 334 380 335 
<< m1 >>
rect 412 334 413 335 
<< m1 >>
rect 413 334 414 335 
<< m1 >>
rect 414 334 415 335 
<< m2 >>
rect 414 334 415 335 
<< m2c >>
rect 414 334 415 335 
<< m1 >>
rect 414 334 415 335 
<< m2 >>
rect 414 334 415 335 
<< m2 >>
rect 415 334 416 335 
<< m1 >>
rect 416 334 417 335 
<< m2 >>
rect 416 334 417 335 
<< m2 >>
rect 417 334 418 335 
<< m1 >>
rect 418 334 419 335 
<< m2 >>
rect 418 334 419 335 
<< m2 >>
rect 419 334 420 335 
<< m1 >>
rect 420 334 421 335 
<< m2 >>
rect 420 334 421 335 
<< m2c >>
rect 420 334 421 335 
<< m1 >>
rect 420 334 421 335 
<< m2 >>
rect 420 334 421 335 
<< m2 >>
rect 421 334 422 335 
<< m1 >>
rect 422 334 423 335 
<< m1 >>
rect 424 334 425 335 
<< m2 >>
rect 424 334 425 335 
<< m2 >>
rect 425 334 426 335 
<< m1 >>
rect 426 334 427 335 
<< m2 >>
rect 426 334 427 335 
<< m2c >>
rect 426 334 427 335 
<< m1 >>
rect 426 334 427 335 
<< m2 >>
rect 426 334 427 335 
<< m1 >>
rect 427 334 428 335 
<< m1 >>
rect 433 334 434 335 
<< m1 >>
rect 435 334 436 335 
<< m1 >>
rect 439 334 440 335 
<< m2 >>
rect 439 334 440 335 
<< m2c >>
rect 439 334 440 335 
<< m1 >>
rect 439 334 440 335 
<< m2 >>
rect 439 334 440 335 
<< m1 >>
rect 451 334 452 335 
<< m1 >>
rect 523 334 524 335 
<< m1 >>
rect 19 335 20 336 
<< m2 >>
rect 20 335 21 336 
<< m2 >>
rect 23 335 24 336 
<< m1 >>
rect 31 335 32 336 
<< m1 >>
rect 44 335 45 336 
<< m2 >>
rect 61 335 62 336 
<< m1 >>
rect 62 335 63 336 
<< m1 >>
rect 64 335 65 336 
<< m1 >>
rect 73 335 74 336 
<< m1 >>
rect 82 335 83 336 
<< m1 >>
rect 85 335 86 336 
<< m1 >>
rect 88 335 89 336 
<< m1 >>
rect 91 335 92 336 
<< m1 >>
rect 100 335 101 336 
<< m1 >>
rect 116 335 117 336 
<< m1 >>
rect 118 335 119 336 
<< m1 >>
rect 124 335 125 336 
<< m1 >>
rect 142 335 143 336 
<< m1 >>
rect 145 335 146 336 
<< m2 >>
rect 146 335 147 336 
<< m1 >>
rect 148 335 149 336 
<< m1 >>
rect 150 335 151 336 
<< m1 >>
rect 154 335 155 336 
<< m1 >>
rect 163 335 164 336 
<< m2 >>
rect 164 335 165 336 
<< m1 >>
rect 178 335 179 336 
<< m1 >>
rect 181 335 182 336 
<< m1 >>
rect 196 335 197 336 
<< m1 >>
rect 204 335 205 336 
<< m1 >>
rect 206 335 207 336 
<< m1 >>
rect 211 335 212 336 
<< m1 >>
rect 217 335 218 336 
<< m1 >>
rect 219 335 220 336 
<< m1 >>
rect 223 335 224 336 
<< m1 >>
rect 225 335 226 336 
<< m1 >>
rect 235 335 236 336 
<< m1 >>
rect 242 335 243 336 
<< m1 >>
rect 244 335 245 336 
<< m2 >>
rect 244 335 245 336 
<< m1 >>
rect 247 335 248 336 
<< m1 >>
rect 253 335 254 336 
<< m1 >>
rect 268 335 269 336 
<< m1 >>
rect 276 335 277 336 
<< m1 >>
rect 286 335 287 336 
<< m1 >>
rect 289 335 290 336 
<< m1 >>
rect 334 335 335 336 
<< m1 >>
rect 347 335 348 336 
<< m2 >>
rect 350 335 351 336 
<< m1 >>
rect 351 335 352 336 
<< m1 >>
rect 355 335 356 336 
<< m1 >>
rect 361 335 362 336 
<< m1 >>
rect 364 335 365 336 
<< m1 >>
rect 370 335 371 336 
<< m1 >>
rect 376 335 377 336 
<< m1 >>
rect 379 335 380 336 
<< m1 >>
rect 412 335 413 336 
<< m1 >>
rect 416 335 417 336 
<< m1 >>
rect 418 335 419 336 
<< m2 >>
rect 421 335 422 336 
<< m1 >>
rect 422 335 423 336 
<< m1 >>
rect 424 335 425 336 
<< m2 >>
rect 424 335 425 336 
<< m1 >>
rect 427 335 428 336 
<< m1 >>
rect 433 335 434 336 
<< m1 >>
rect 435 335 436 336 
<< m1 >>
rect 439 335 440 336 
<< m1 >>
rect 451 335 452 336 
<< m1 >>
rect 523 335 524 336 
<< pdiffusion >>
rect 12 336 13 337 
<< pdiffusion >>
rect 13 336 14 337 
<< pdiffusion >>
rect 14 336 15 337 
<< pdiffusion >>
rect 15 336 16 337 
<< pdiffusion >>
rect 16 336 17 337 
<< pdiffusion >>
rect 17 336 18 337 
<< m1 >>
rect 19 336 20 337 
<< m2 >>
rect 20 336 21 337 
<< m1 >>
rect 23 336 24 337 
<< m2 >>
rect 23 336 24 337 
<< m2c >>
rect 23 336 24 337 
<< m1 >>
rect 23 336 24 337 
<< m2 >>
rect 23 336 24 337 
<< pdiffusion >>
rect 30 336 31 337 
<< m1 >>
rect 31 336 32 337 
<< pdiffusion >>
rect 31 336 32 337 
<< pdiffusion >>
rect 32 336 33 337 
<< pdiffusion >>
rect 33 336 34 337 
<< pdiffusion >>
rect 34 336 35 337 
<< pdiffusion >>
rect 35 336 36 337 
<< m1 >>
rect 44 336 45 337 
<< pdiffusion >>
rect 48 336 49 337 
<< pdiffusion >>
rect 49 336 50 337 
<< pdiffusion >>
rect 50 336 51 337 
<< pdiffusion >>
rect 51 336 52 337 
<< pdiffusion >>
rect 52 336 53 337 
<< pdiffusion >>
rect 53 336 54 337 
<< m2 >>
rect 61 336 62 337 
<< m1 >>
rect 62 336 63 337 
<< m1 >>
rect 64 336 65 337 
<< pdiffusion >>
rect 66 336 67 337 
<< pdiffusion >>
rect 67 336 68 337 
<< pdiffusion >>
rect 68 336 69 337 
<< pdiffusion >>
rect 69 336 70 337 
<< pdiffusion >>
rect 70 336 71 337 
<< pdiffusion >>
rect 71 336 72 337 
<< m1 >>
rect 73 336 74 337 
<< m1 >>
rect 82 336 83 337 
<< pdiffusion >>
rect 84 336 85 337 
<< m1 >>
rect 85 336 86 337 
<< pdiffusion >>
rect 85 336 86 337 
<< pdiffusion >>
rect 86 336 87 337 
<< pdiffusion >>
rect 87 336 88 337 
<< m1 >>
rect 88 336 89 337 
<< pdiffusion >>
rect 88 336 89 337 
<< pdiffusion >>
rect 89 336 90 337 
<< m1 >>
rect 91 336 92 337 
<< m1 >>
rect 100 336 101 337 
<< m1 >>
rect 116 336 117 337 
<< m1 >>
rect 118 336 119 337 
<< pdiffusion >>
rect 120 336 121 337 
<< pdiffusion >>
rect 121 336 122 337 
<< pdiffusion >>
rect 122 336 123 337 
<< pdiffusion >>
rect 123 336 124 337 
<< m1 >>
rect 124 336 125 337 
<< pdiffusion >>
rect 124 336 125 337 
<< pdiffusion >>
rect 125 336 126 337 
<< pdiffusion >>
rect 138 336 139 337 
<< pdiffusion >>
rect 139 336 140 337 
<< pdiffusion >>
rect 140 336 141 337 
<< pdiffusion >>
rect 141 336 142 337 
<< m1 >>
rect 142 336 143 337 
<< pdiffusion >>
rect 142 336 143 337 
<< pdiffusion >>
rect 143 336 144 337 
<< m1 >>
rect 145 336 146 337 
<< m2 >>
rect 146 336 147 337 
<< m1 >>
rect 148 336 149 337 
<< m1 >>
rect 150 336 151 337 
<< m1 >>
rect 154 336 155 337 
<< pdiffusion >>
rect 156 336 157 337 
<< pdiffusion >>
rect 157 336 158 337 
<< pdiffusion >>
rect 158 336 159 337 
<< pdiffusion >>
rect 159 336 160 337 
<< pdiffusion >>
rect 160 336 161 337 
<< pdiffusion >>
rect 161 336 162 337 
<< m1 >>
rect 163 336 164 337 
<< m2 >>
rect 164 336 165 337 
<< pdiffusion >>
rect 174 336 175 337 
<< pdiffusion >>
rect 175 336 176 337 
<< pdiffusion >>
rect 176 336 177 337 
<< pdiffusion >>
rect 177 336 178 337 
<< m1 >>
rect 178 336 179 337 
<< pdiffusion >>
rect 178 336 179 337 
<< pdiffusion >>
rect 179 336 180 337 
<< m1 >>
rect 181 336 182 337 
<< pdiffusion >>
rect 192 336 193 337 
<< pdiffusion >>
rect 193 336 194 337 
<< pdiffusion >>
rect 194 336 195 337 
<< pdiffusion >>
rect 195 336 196 337 
<< m1 >>
rect 196 336 197 337 
<< pdiffusion >>
rect 196 336 197 337 
<< pdiffusion >>
rect 197 336 198 337 
<< m1 >>
rect 204 336 205 337 
<< m1 >>
rect 206 336 207 337 
<< pdiffusion >>
rect 210 336 211 337 
<< m1 >>
rect 211 336 212 337 
<< pdiffusion >>
rect 211 336 212 337 
<< pdiffusion >>
rect 212 336 213 337 
<< pdiffusion >>
rect 213 336 214 337 
<< pdiffusion >>
rect 214 336 215 337 
<< pdiffusion >>
rect 215 336 216 337 
<< m1 >>
rect 217 336 218 337 
<< m1 >>
rect 219 336 220 337 
<< m1 >>
rect 223 336 224 337 
<< m1 >>
rect 225 336 226 337 
<< pdiffusion >>
rect 228 336 229 337 
<< pdiffusion >>
rect 229 336 230 337 
<< pdiffusion >>
rect 230 336 231 337 
<< pdiffusion >>
rect 231 336 232 337 
<< pdiffusion >>
rect 232 336 233 337 
<< pdiffusion >>
rect 233 336 234 337 
<< m1 >>
rect 235 336 236 337 
<< m1 >>
rect 242 336 243 337 
<< m1 >>
rect 244 336 245 337 
<< m2 >>
rect 244 336 245 337 
<< pdiffusion >>
rect 246 336 247 337 
<< m1 >>
rect 247 336 248 337 
<< pdiffusion >>
rect 247 336 248 337 
<< pdiffusion >>
rect 248 336 249 337 
<< pdiffusion >>
rect 249 336 250 337 
<< pdiffusion >>
rect 250 336 251 337 
<< pdiffusion >>
rect 251 336 252 337 
<< m1 >>
rect 253 336 254 337 
<< pdiffusion >>
rect 264 336 265 337 
<< pdiffusion >>
rect 265 336 266 337 
<< pdiffusion >>
rect 266 336 267 337 
<< pdiffusion >>
rect 267 336 268 337 
<< m1 >>
rect 268 336 269 337 
<< pdiffusion >>
rect 268 336 269 337 
<< pdiffusion >>
rect 269 336 270 337 
<< m1 >>
rect 276 336 277 337 
<< pdiffusion >>
rect 282 336 283 337 
<< pdiffusion >>
rect 283 336 284 337 
<< pdiffusion >>
rect 284 336 285 337 
<< pdiffusion >>
rect 285 336 286 337 
<< m1 >>
rect 286 336 287 337 
<< pdiffusion >>
rect 286 336 287 337 
<< pdiffusion >>
rect 287 336 288 337 
<< m1 >>
rect 289 336 290 337 
<< pdiffusion >>
rect 300 336 301 337 
<< pdiffusion >>
rect 301 336 302 337 
<< pdiffusion >>
rect 302 336 303 337 
<< pdiffusion >>
rect 303 336 304 337 
<< pdiffusion >>
rect 304 336 305 337 
<< pdiffusion >>
rect 305 336 306 337 
<< pdiffusion >>
rect 318 336 319 337 
<< pdiffusion >>
rect 319 336 320 337 
<< pdiffusion >>
rect 320 336 321 337 
<< pdiffusion >>
rect 321 336 322 337 
<< pdiffusion >>
rect 322 336 323 337 
<< pdiffusion >>
rect 323 336 324 337 
<< m1 >>
rect 334 336 335 337 
<< pdiffusion >>
rect 336 336 337 337 
<< pdiffusion >>
rect 337 336 338 337 
<< pdiffusion >>
rect 338 336 339 337 
<< pdiffusion >>
rect 339 336 340 337 
<< pdiffusion >>
rect 340 336 341 337 
<< pdiffusion >>
rect 341 336 342 337 
<< m1 >>
rect 347 336 348 337 
<< m2 >>
rect 350 336 351 337 
<< m1 >>
rect 351 336 352 337 
<< pdiffusion >>
rect 354 336 355 337 
<< m1 >>
rect 355 336 356 337 
<< pdiffusion >>
rect 355 336 356 337 
<< pdiffusion >>
rect 356 336 357 337 
<< pdiffusion >>
rect 357 336 358 337 
<< pdiffusion >>
rect 358 336 359 337 
<< pdiffusion >>
rect 359 336 360 337 
<< m1 >>
rect 361 336 362 337 
<< m1 >>
rect 364 336 365 337 
<< m1 >>
rect 370 336 371 337 
<< pdiffusion >>
rect 372 336 373 337 
<< pdiffusion >>
rect 373 336 374 337 
<< pdiffusion >>
rect 374 336 375 337 
<< pdiffusion >>
rect 375 336 376 337 
<< m1 >>
rect 376 336 377 337 
<< pdiffusion >>
rect 376 336 377 337 
<< pdiffusion >>
rect 377 336 378 337 
<< m1 >>
rect 379 336 380 337 
<< pdiffusion >>
rect 390 336 391 337 
<< pdiffusion >>
rect 391 336 392 337 
<< pdiffusion >>
rect 392 336 393 337 
<< pdiffusion >>
rect 393 336 394 337 
<< pdiffusion >>
rect 394 336 395 337 
<< pdiffusion >>
rect 395 336 396 337 
<< pdiffusion >>
rect 408 336 409 337 
<< pdiffusion >>
rect 409 336 410 337 
<< pdiffusion >>
rect 410 336 411 337 
<< pdiffusion >>
rect 411 336 412 337 
<< m1 >>
rect 412 336 413 337 
<< pdiffusion >>
rect 412 336 413 337 
<< pdiffusion >>
rect 413 336 414 337 
<< m1 >>
rect 416 336 417 337 
<< m1 >>
rect 418 336 419 337 
<< m2 >>
rect 421 336 422 337 
<< m1 >>
rect 422 336 423 337 
<< m1 >>
rect 424 336 425 337 
<< m2 >>
rect 424 336 425 337 
<< pdiffusion >>
rect 426 336 427 337 
<< m1 >>
rect 427 336 428 337 
<< pdiffusion >>
rect 427 336 428 337 
<< pdiffusion >>
rect 428 336 429 337 
<< pdiffusion >>
rect 429 336 430 337 
<< pdiffusion >>
rect 430 336 431 337 
<< pdiffusion >>
rect 431 336 432 337 
<< m1 >>
rect 433 336 434 337 
<< m1 >>
rect 435 336 436 337 
<< m1 >>
rect 439 336 440 337 
<< pdiffusion >>
rect 444 336 445 337 
<< pdiffusion >>
rect 445 336 446 337 
<< pdiffusion >>
rect 446 336 447 337 
<< pdiffusion >>
rect 447 336 448 337 
<< pdiffusion >>
rect 448 336 449 337 
<< pdiffusion >>
rect 449 336 450 337 
<< m1 >>
rect 451 336 452 337 
<< pdiffusion >>
rect 462 336 463 337 
<< pdiffusion >>
rect 463 336 464 337 
<< pdiffusion >>
rect 464 336 465 337 
<< pdiffusion >>
rect 465 336 466 337 
<< pdiffusion >>
rect 466 336 467 337 
<< pdiffusion >>
rect 467 336 468 337 
<< pdiffusion >>
rect 480 336 481 337 
<< pdiffusion >>
rect 481 336 482 337 
<< pdiffusion >>
rect 482 336 483 337 
<< pdiffusion >>
rect 483 336 484 337 
<< pdiffusion >>
rect 484 336 485 337 
<< pdiffusion >>
rect 485 336 486 337 
<< pdiffusion >>
rect 498 336 499 337 
<< pdiffusion >>
rect 499 336 500 337 
<< pdiffusion >>
rect 500 336 501 337 
<< pdiffusion >>
rect 501 336 502 337 
<< pdiffusion >>
rect 502 336 503 337 
<< pdiffusion >>
rect 503 336 504 337 
<< pdiffusion >>
rect 516 336 517 337 
<< pdiffusion >>
rect 517 336 518 337 
<< pdiffusion >>
rect 518 336 519 337 
<< pdiffusion >>
rect 519 336 520 337 
<< pdiffusion >>
rect 520 336 521 337 
<< pdiffusion >>
rect 521 336 522 337 
<< m1 >>
rect 523 336 524 337 
<< pdiffusion >>
rect 12 337 13 338 
<< pdiffusion >>
rect 13 337 14 338 
<< pdiffusion >>
rect 14 337 15 338 
<< pdiffusion >>
rect 15 337 16 338 
<< pdiffusion >>
rect 16 337 17 338 
<< pdiffusion >>
rect 17 337 18 338 
<< m1 >>
rect 19 337 20 338 
<< m2 >>
rect 20 337 21 338 
<< m1 >>
rect 23 337 24 338 
<< pdiffusion >>
rect 30 337 31 338 
<< pdiffusion >>
rect 31 337 32 338 
<< pdiffusion >>
rect 32 337 33 338 
<< pdiffusion >>
rect 33 337 34 338 
<< pdiffusion >>
rect 34 337 35 338 
<< pdiffusion >>
rect 35 337 36 338 
<< m1 >>
rect 44 337 45 338 
<< pdiffusion >>
rect 48 337 49 338 
<< pdiffusion >>
rect 49 337 50 338 
<< pdiffusion >>
rect 50 337 51 338 
<< pdiffusion >>
rect 51 337 52 338 
<< pdiffusion >>
rect 52 337 53 338 
<< pdiffusion >>
rect 53 337 54 338 
<< m2 >>
rect 61 337 62 338 
<< m1 >>
rect 62 337 63 338 
<< m1 >>
rect 64 337 65 338 
<< pdiffusion >>
rect 66 337 67 338 
<< pdiffusion >>
rect 67 337 68 338 
<< pdiffusion >>
rect 68 337 69 338 
<< pdiffusion >>
rect 69 337 70 338 
<< pdiffusion >>
rect 70 337 71 338 
<< pdiffusion >>
rect 71 337 72 338 
<< m1 >>
rect 73 337 74 338 
<< m1 >>
rect 82 337 83 338 
<< pdiffusion >>
rect 84 337 85 338 
<< pdiffusion >>
rect 85 337 86 338 
<< pdiffusion >>
rect 86 337 87 338 
<< pdiffusion >>
rect 87 337 88 338 
<< pdiffusion >>
rect 88 337 89 338 
<< pdiffusion >>
rect 89 337 90 338 
<< m1 >>
rect 91 337 92 338 
<< m1 >>
rect 100 337 101 338 
<< m1 >>
rect 116 337 117 338 
<< m1 >>
rect 118 337 119 338 
<< pdiffusion >>
rect 120 337 121 338 
<< pdiffusion >>
rect 121 337 122 338 
<< pdiffusion >>
rect 122 337 123 338 
<< pdiffusion >>
rect 123 337 124 338 
<< pdiffusion >>
rect 124 337 125 338 
<< pdiffusion >>
rect 125 337 126 338 
<< pdiffusion >>
rect 138 337 139 338 
<< pdiffusion >>
rect 139 337 140 338 
<< pdiffusion >>
rect 140 337 141 338 
<< pdiffusion >>
rect 141 337 142 338 
<< pdiffusion >>
rect 142 337 143 338 
<< pdiffusion >>
rect 143 337 144 338 
<< m1 >>
rect 145 337 146 338 
<< m2 >>
rect 146 337 147 338 
<< m1 >>
rect 148 337 149 338 
<< m1 >>
rect 150 337 151 338 
<< m1 >>
rect 154 337 155 338 
<< pdiffusion >>
rect 156 337 157 338 
<< pdiffusion >>
rect 157 337 158 338 
<< pdiffusion >>
rect 158 337 159 338 
<< pdiffusion >>
rect 159 337 160 338 
<< pdiffusion >>
rect 160 337 161 338 
<< pdiffusion >>
rect 161 337 162 338 
<< m1 >>
rect 163 337 164 338 
<< m2 >>
rect 164 337 165 338 
<< pdiffusion >>
rect 174 337 175 338 
<< pdiffusion >>
rect 175 337 176 338 
<< pdiffusion >>
rect 176 337 177 338 
<< pdiffusion >>
rect 177 337 178 338 
<< pdiffusion >>
rect 178 337 179 338 
<< pdiffusion >>
rect 179 337 180 338 
<< m1 >>
rect 181 337 182 338 
<< pdiffusion >>
rect 192 337 193 338 
<< pdiffusion >>
rect 193 337 194 338 
<< pdiffusion >>
rect 194 337 195 338 
<< pdiffusion >>
rect 195 337 196 338 
<< pdiffusion >>
rect 196 337 197 338 
<< pdiffusion >>
rect 197 337 198 338 
<< m1 >>
rect 204 337 205 338 
<< m1 >>
rect 206 337 207 338 
<< pdiffusion >>
rect 210 337 211 338 
<< pdiffusion >>
rect 211 337 212 338 
<< pdiffusion >>
rect 212 337 213 338 
<< pdiffusion >>
rect 213 337 214 338 
<< pdiffusion >>
rect 214 337 215 338 
<< pdiffusion >>
rect 215 337 216 338 
<< m1 >>
rect 217 337 218 338 
<< m1 >>
rect 219 337 220 338 
<< m1 >>
rect 223 337 224 338 
<< m1 >>
rect 225 337 226 338 
<< pdiffusion >>
rect 228 337 229 338 
<< pdiffusion >>
rect 229 337 230 338 
<< pdiffusion >>
rect 230 337 231 338 
<< pdiffusion >>
rect 231 337 232 338 
<< pdiffusion >>
rect 232 337 233 338 
<< pdiffusion >>
rect 233 337 234 338 
<< m1 >>
rect 235 337 236 338 
<< m1 >>
rect 242 337 243 338 
<< m1 >>
rect 244 337 245 338 
<< m2 >>
rect 244 337 245 338 
<< pdiffusion >>
rect 246 337 247 338 
<< pdiffusion >>
rect 247 337 248 338 
<< pdiffusion >>
rect 248 337 249 338 
<< pdiffusion >>
rect 249 337 250 338 
<< pdiffusion >>
rect 250 337 251 338 
<< pdiffusion >>
rect 251 337 252 338 
<< m1 >>
rect 253 337 254 338 
<< pdiffusion >>
rect 264 337 265 338 
<< pdiffusion >>
rect 265 337 266 338 
<< pdiffusion >>
rect 266 337 267 338 
<< pdiffusion >>
rect 267 337 268 338 
<< pdiffusion >>
rect 268 337 269 338 
<< pdiffusion >>
rect 269 337 270 338 
<< m1 >>
rect 276 337 277 338 
<< pdiffusion >>
rect 282 337 283 338 
<< pdiffusion >>
rect 283 337 284 338 
<< pdiffusion >>
rect 284 337 285 338 
<< pdiffusion >>
rect 285 337 286 338 
<< pdiffusion >>
rect 286 337 287 338 
<< pdiffusion >>
rect 287 337 288 338 
<< m1 >>
rect 289 337 290 338 
<< pdiffusion >>
rect 300 337 301 338 
<< pdiffusion >>
rect 301 337 302 338 
<< pdiffusion >>
rect 302 337 303 338 
<< pdiffusion >>
rect 303 337 304 338 
<< pdiffusion >>
rect 304 337 305 338 
<< pdiffusion >>
rect 305 337 306 338 
<< pdiffusion >>
rect 318 337 319 338 
<< pdiffusion >>
rect 319 337 320 338 
<< pdiffusion >>
rect 320 337 321 338 
<< pdiffusion >>
rect 321 337 322 338 
<< pdiffusion >>
rect 322 337 323 338 
<< pdiffusion >>
rect 323 337 324 338 
<< m1 >>
rect 334 337 335 338 
<< pdiffusion >>
rect 336 337 337 338 
<< pdiffusion >>
rect 337 337 338 338 
<< pdiffusion >>
rect 338 337 339 338 
<< pdiffusion >>
rect 339 337 340 338 
<< pdiffusion >>
rect 340 337 341 338 
<< pdiffusion >>
rect 341 337 342 338 
<< m1 >>
rect 347 337 348 338 
<< m2 >>
rect 350 337 351 338 
<< m1 >>
rect 351 337 352 338 
<< pdiffusion >>
rect 354 337 355 338 
<< pdiffusion >>
rect 355 337 356 338 
<< pdiffusion >>
rect 356 337 357 338 
<< pdiffusion >>
rect 357 337 358 338 
<< pdiffusion >>
rect 358 337 359 338 
<< pdiffusion >>
rect 359 337 360 338 
<< m1 >>
rect 361 337 362 338 
<< m1 >>
rect 364 337 365 338 
<< m1 >>
rect 370 337 371 338 
<< pdiffusion >>
rect 372 337 373 338 
<< pdiffusion >>
rect 373 337 374 338 
<< pdiffusion >>
rect 374 337 375 338 
<< pdiffusion >>
rect 375 337 376 338 
<< pdiffusion >>
rect 376 337 377 338 
<< pdiffusion >>
rect 377 337 378 338 
<< m1 >>
rect 379 337 380 338 
<< pdiffusion >>
rect 390 337 391 338 
<< pdiffusion >>
rect 391 337 392 338 
<< pdiffusion >>
rect 392 337 393 338 
<< pdiffusion >>
rect 393 337 394 338 
<< pdiffusion >>
rect 394 337 395 338 
<< pdiffusion >>
rect 395 337 396 338 
<< pdiffusion >>
rect 408 337 409 338 
<< pdiffusion >>
rect 409 337 410 338 
<< pdiffusion >>
rect 410 337 411 338 
<< pdiffusion >>
rect 411 337 412 338 
<< pdiffusion >>
rect 412 337 413 338 
<< pdiffusion >>
rect 413 337 414 338 
<< m1 >>
rect 416 337 417 338 
<< m1 >>
rect 418 337 419 338 
<< m2 >>
rect 421 337 422 338 
<< m1 >>
rect 422 337 423 338 
<< m1 >>
rect 424 337 425 338 
<< m2 >>
rect 424 337 425 338 
<< pdiffusion >>
rect 426 337 427 338 
<< pdiffusion >>
rect 427 337 428 338 
<< pdiffusion >>
rect 428 337 429 338 
<< pdiffusion >>
rect 429 337 430 338 
<< pdiffusion >>
rect 430 337 431 338 
<< pdiffusion >>
rect 431 337 432 338 
<< m1 >>
rect 433 337 434 338 
<< m1 >>
rect 435 337 436 338 
<< m1 >>
rect 439 337 440 338 
<< pdiffusion >>
rect 444 337 445 338 
<< pdiffusion >>
rect 445 337 446 338 
<< pdiffusion >>
rect 446 337 447 338 
<< pdiffusion >>
rect 447 337 448 338 
<< pdiffusion >>
rect 448 337 449 338 
<< pdiffusion >>
rect 449 337 450 338 
<< m1 >>
rect 451 337 452 338 
<< pdiffusion >>
rect 462 337 463 338 
<< pdiffusion >>
rect 463 337 464 338 
<< pdiffusion >>
rect 464 337 465 338 
<< pdiffusion >>
rect 465 337 466 338 
<< pdiffusion >>
rect 466 337 467 338 
<< pdiffusion >>
rect 467 337 468 338 
<< pdiffusion >>
rect 480 337 481 338 
<< pdiffusion >>
rect 481 337 482 338 
<< pdiffusion >>
rect 482 337 483 338 
<< pdiffusion >>
rect 483 337 484 338 
<< pdiffusion >>
rect 484 337 485 338 
<< pdiffusion >>
rect 485 337 486 338 
<< pdiffusion >>
rect 498 337 499 338 
<< pdiffusion >>
rect 499 337 500 338 
<< pdiffusion >>
rect 500 337 501 338 
<< pdiffusion >>
rect 501 337 502 338 
<< pdiffusion >>
rect 502 337 503 338 
<< pdiffusion >>
rect 503 337 504 338 
<< pdiffusion >>
rect 516 337 517 338 
<< pdiffusion >>
rect 517 337 518 338 
<< pdiffusion >>
rect 518 337 519 338 
<< pdiffusion >>
rect 519 337 520 338 
<< pdiffusion >>
rect 520 337 521 338 
<< pdiffusion >>
rect 521 337 522 338 
<< m1 >>
rect 523 337 524 338 
<< pdiffusion >>
rect 12 338 13 339 
<< pdiffusion >>
rect 13 338 14 339 
<< pdiffusion >>
rect 14 338 15 339 
<< pdiffusion >>
rect 15 338 16 339 
<< pdiffusion >>
rect 16 338 17 339 
<< pdiffusion >>
rect 17 338 18 339 
<< m1 >>
rect 19 338 20 339 
<< m2 >>
rect 20 338 21 339 
<< m1 >>
rect 23 338 24 339 
<< pdiffusion >>
rect 30 338 31 339 
<< pdiffusion >>
rect 31 338 32 339 
<< pdiffusion >>
rect 32 338 33 339 
<< pdiffusion >>
rect 33 338 34 339 
<< pdiffusion >>
rect 34 338 35 339 
<< pdiffusion >>
rect 35 338 36 339 
<< m1 >>
rect 44 338 45 339 
<< pdiffusion >>
rect 48 338 49 339 
<< pdiffusion >>
rect 49 338 50 339 
<< pdiffusion >>
rect 50 338 51 339 
<< pdiffusion >>
rect 51 338 52 339 
<< pdiffusion >>
rect 52 338 53 339 
<< pdiffusion >>
rect 53 338 54 339 
<< m2 >>
rect 61 338 62 339 
<< m1 >>
rect 62 338 63 339 
<< m1 >>
rect 64 338 65 339 
<< pdiffusion >>
rect 66 338 67 339 
<< pdiffusion >>
rect 67 338 68 339 
<< pdiffusion >>
rect 68 338 69 339 
<< pdiffusion >>
rect 69 338 70 339 
<< pdiffusion >>
rect 70 338 71 339 
<< pdiffusion >>
rect 71 338 72 339 
<< m1 >>
rect 73 338 74 339 
<< m1 >>
rect 82 338 83 339 
<< pdiffusion >>
rect 84 338 85 339 
<< pdiffusion >>
rect 85 338 86 339 
<< pdiffusion >>
rect 86 338 87 339 
<< pdiffusion >>
rect 87 338 88 339 
<< pdiffusion >>
rect 88 338 89 339 
<< pdiffusion >>
rect 89 338 90 339 
<< m1 >>
rect 91 338 92 339 
<< m1 >>
rect 100 338 101 339 
<< m1 >>
rect 116 338 117 339 
<< m1 >>
rect 118 338 119 339 
<< pdiffusion >>
rect 120 338 121 339 
<< pdiffusion >>
rect 121 338 122 339 
<< pdiffusion >>
rect 122 338 123 339 
<< pdiffusion >>
rect 123 338 124 339 
<< pdiffusion >>
rect 124 338 125 339 
<< pdiffusion >>
rect 125 338 126 339 
<< pdiffusion >>
rect 138 338 139 339 
<< pdiffusion >>
rect 139 338 140 339 
<< pdiffusion >>
rect 140 338 141 339 
<< pdiffusion >>
rect 141 338 142 339 
<< pdiffusion >>
rect 142 338 143 339 
<< pdiffusion >>
rect 143 338 144 339 
<< m1 >>
rect 145 338 146 339 
<< m2 >>
rect 146 338 147 339 
<< m1 >>
rect 148 338 149 339 
<< m1 >>
rect 150 338 151 339 
<< m1 >>
rect 154 338 155 339 
<< pdiffusion >>
rect 156 338 157 339 
<< pdiffusion >>
rect 157 338 158 339 
<< pdiffusion >>
rect 158 338 159 339 
<< pdiffusion >>
rect 159 338 160 339 
<< pdiffusion >>
rect 160 338 161 339 
<< pdiffusion >>
rect 161 338 162 339 
<< m1 >>
rect 163 338 164 339 
<< m2 >>
rect 164 338 165 339 
<< pdiffusion >>
rect 174 338 175 339 
<< pdiffusion >>
rect 175 338 176 339 
<< pdiffusion >>
rect 176 338 177 339 
<< pdiffusion >>
rect 177 338 178 339 
<< pdiffusion >>
rect 178 338 179 339 
<< pdiffusion >>
rect 179 338 180 339 
<< m1 >>
rect 181 338 182 339 
<< pdiffusion >>
rect 192 338 193 339 
<< pdiffusion >>
rect 193 338 194 339 
<< pdiffusion >>
rect 194 338 195 339 
<< pdiffusion >>
rect 195 338 196 339 
<< pdiffusion >>
rect 196 338 197 339 
<< pdiffusion >>
rect 197 338 198 339 
<< m1 >>
rect 204 338 205 339 
<< m1 >>
rect 206 338 207 339 
<< pdiffusion >>
rect 210 338 211 339 
<< pdiffusion >>
rect 211 338 212 339 
<< pdiffusion >>
rect 212 338 213 339 
<< pdiffusion >>
rect 213 338 214 339 
<< pdiffusion >>
rect 214 338 215 339 
<< pdiffusion >>
rect 215 338 216 339 
<< m1 >>
rect 217 338 218 339 
<< m1 >>
rect 219 338 220 339 
<< m1 >>
rect 223 338 224 339 
<< m1 >>
rect 225 338 226 339 
<< pdiffusion >>
rect 228 338 229 339 
<< pdiffusion >>
rect 229 338 230 339 
<< pdiffusion >>
rect 230 338 231 339 
<< pdiffusion >>
rect 231 338 232 339 
<< pdiffusion >>
rect 232 338 233 339 
<< pdiffusion >>
rect 233 338 234 339 
<< m1 >>
rect 235 338 236 339 
<< m1 >>
rect 242 338 243 339 
<< m1 >>
rect 244 338 245 339 
<< m2 >>
rect 244 338 245 339 
<< pdiffusion >>
rect 246 338 247 339 
<< pdiffusion >>
rect 247 338 248 339 
<< pdiffusion >>
rect 248 338 249 339 
<< pdiffusion >>
rect 249 338 250 339 
<< pdiffusion >>
rect 250 338 251 339 
<< pdiffusion >>
rect 251 338 252 339 
<< m1 >>
rect 253 338 254 339 
<< pdiffusion >>
rect 264 338 265 339 
<< pdiffusion >>
rect 265 338 266 339 
<< pdiffusion >>
rect 266 338 267 339 
<< pdiffusion >>
rect 267 338 268 339 
<< pdiffusion >>
rect 268 338 269 339 
<< pdiffusion >>
rect 269 338 270 339 
<< m1 >>
rect 276 338 277 339 
<< pdiffusion >>
rect 282 338 283 339 
<< pdiffusion >>
rect 283 338 284 339 
<< pdiffusion >>
rect 284 338 285 339 
<< pdiffusion >>
rect 285 338 286 339 
<< pdiffusion >>
rect 286 338 287 339 
<< pdiffusion >>
rect 287 338 288 339 
<< m1 >>
rect 289 338 290 339 
<< pdiffusion >>
rect 300 338 301 339 
<< pdiffusion >>
rect 301 338 302 339 
<< pdiffusion >>
rect 302 338 303 339 
<< pdiffusion >>
rect 303 338 304 339 
<< pdiffusion >>
rect 304 338 305 339 
<< pdiffusion >>
rect 305 338 306 339 
<< pdiffusion >>
rect 318 338 319 339 
<< pdiffusion >>
rect 319 338 320 339 
<< pdiffusion >>
rect 320 338 321 339 
<< pdiffusion >>
rect 321 338 322 339 
<< pdiffusion >>
rect 322 338 323 339 
<< pdiffusion >>
rect 323 338 324 339 
<< m1 >>
rect 334 338 335 339 
<< pdiffusion >>
rect 336 338 337 339 
<< pdiffusion >>
rect 337 338 338 339 
<< pdiffusion >>
rect 338 338 339 339 
<< pdiffusion >>
rect 339 338 340 339 
<< pdiffusion >>
rect 340 338 341 339 
<< pdiffusion >>
rect 341 338 342 339 
<< m1 >>
rect 347 338 348 339 
<< m2 >>
rect 350 338 351 339 
<< m1 >>
rect 351 338 352 339 
<< pdiffusion >>
rect 354 338 355 339 
<< pdiffusion >>
rect 355 338 356 339 
<< pdiffusion >>
rect 356 338 357 339 
<< pdiffusion >>
rect 357 338 358 339 
<< pdiffusion >>
rect 358 338 359 339 
<< pdiffusion >>
rect 359 338 360 339 
<< m1 >>
rect 361 338 362 339 
<< m1 >>
rect 364 338 365 339 
<< m1 >>
rect 370 338 371 339 
<< pdiffusion >>
rect 372 338 373 339 
<< pdiffusion >>
rect 373 338 374 339 
<< pdiffusion >>
rect 374 338 375 339 
<< pdiffusion >>
rect 375 338 376 339 
<< pdiffusion >>
rect 376 338 377 339 
<< pdiffusion >>
rect 377 338 378 339 
<< m1 >>
rect 379 338 380 339 
<< pdiffusion >>
rect 390 338 391 339 
<< pdiffusion >>
rect 391 338 392 339 
<< pdiffusion >>
rect 392 338 393 339 
<< pdiffusion >>
rect 393 338 394 339 
<< pdiffusion >>
rect 394 338 395 339 
<< pdiffusion >>
rect 395 338 396 339 
<< pdiffusion >>
rect 408 338 409 339 
<< pdiffusion >>
rect 409 338 410 339 
<< pdiffusion >>
rect 410 338 411 339 
<< pdiffusion >>
rect 411 338 412 339 
<< pdiffusion >>
rect 412 338 413 339 
<< pdiffusion >>
rect 413 338 414 339 
<< m1 >>
rect 416 338 417 339 
<< m1 >>
rect 418 338 419 339 
<< m2 >>
rect 421 338 422 339 
<< m1 >>
rect 422 338 423 339 
<< m1 >>
rect 424 338 425 339 
<< m2 >>
rect 424 338 425 339 
<< pdiffusion >>
rect 426 338 427 339 
<< pdiffusion >>
rect 427 338 428 339 
<< pdiffusion >>
rect 428 338 429 339 
<< pdiffusion >>
rect 429 338 430 339 
<< pdiffusion >>
rect 430 338 431 339 
<< pdiffusion >>
rect 431 338 432 339 
<< m1 >>
rect 433 338 434 339 
<< m1 >>
rect 435 338 436 339 
<< m1 >>
rect 439 338 440 339 
<< pdiffusion >>
rect 444 338 445 339 
<< pdiffusion >>
rect 445 338 446 339 
<< pdiffusion >>
rect 446 338 447 339 
<< pdiffusion >>
rect 447 338 448 339 
<< pdiffusion >>
rect 448 338 449 339 
<< pdiffusion >>
rect 449 338 450 339 
<< m1 >>
rect 451 338 452 339 
<< pdiffusion >>
rect 462 338 463 339 
<< pdiffusion >>
rect 463 338 464 339 
<< pdiffusion >>
rect 464 338 465 339 
<< pdiffusion >>
rect 465 338 466 339 
<< pdiffusion >>
rect 466 338 467 339 
<< pdiffusion >>
rect 467 338 468 339 
<< pdiffusion >>
rect 480 338 481 339 
<< pdiffusion >>
rect 481 338 482 339 
<< pdiffusion >>
rect 482 338 483 339 
<< pdiffusion >>
rect 483 338 484 339 
<< pdiffusion >>
rect 484 338 485 339 
<< pdiffusion >>
rect 485 338 486 339 
<< pdiffusion >>
rect 498 338 499 339 
<< pdiffusion >>
rect 499 338 500 339 
<< pdiffusion >>
rect 500 338 501 339 
<< pdiffusion >>
rect 501 338 502 339 
<< pdiffusion >>
rect 502 338 503 339 
<< pdiffusion >>
rect 503 338 504 339 
<< pdiffusion >>
rect 516 338 517 339 
<< pdiffusion >>
rect 517 338 518 339 
<< pdiffusion >>
rect 518 338 519 339 
<< pdiffusion >>
rect 519 338 520 339 
<< pdiffusion >>
rect 520 338 521 339 
<< pdiffusion >>
rect 521 338 522 339 
<< m1 >>
rect 523 338 524 339 
<< pdiffusion >>
rect 12 339 13 340 
<< pdiffusion >>
rect 13 339 14 340 
<< pdiffusion >>
rect 14 339 15 340 
<< pdiffusion >>
rect 15 339 16 340 
<< pdiffusion >>
rect 16 339 17 340 
<< pdiffusion >>
rect 17 339 18 340 
<< m1 >>
rect 19 339 20 340 
<< m2 >>
rect 20 339 21 340 
<< m1 >>
rect 23 339 24 340 
<< pdiffusion >>
rect 30 339 31 340 
<< pdiffusion >>
rect 31 339 32 340 
<< pdiffusion >>
rect 32 339 33 340 
<< pdiffusion >>
rect 33 339 34 340 
<< pdiffusion >>
rect 34 339 35 340 
<< pdiffusion >>
rect 35 339 36 340 
<< m1 >>
rect 44 339 45 340 
<< pdiffusion >>
rect 48 339 49 340 
<< pdiffusion >>
rect 49 339 50 340 
<< pdiffusion >>
rect 50 339 51 340 
<< pdiffusion >>
rect 51 339 52 340 
<< pdiffusion >>
rect 52 339 53 340 
<< pdiffusion >>
rect 53 339 54 340 
<< m2 >>
rect 61 339 62 340 
<< m1 >>
rect 62 339 63 340 
<< m1 >>
rect 64 339 65 340 
<< pdiffusion >>
rect 66 339 67 340 
<< pdiffusion >>
rect 67 339 68 340 
<< pdiffusion >>
rect 68 339 69 340 
<< pdiffusion >>
rect 69 339 70 340 
<< pdiffusion >>
rect 70 339 71 340 
<< pdiffusion >>
rect 71 339 72 340 
<< m1 >>
rect 73 339 74 340 
<< m1 >>
rect 82 339 83 340 
<< pdiffusion >>
rect 84 339 85 340 
<< pdiffusion >>
rect 85 339 86 340 
<< pdiffusion >>
rect 86 339 87 340 
<< pdiffusion >>
rect 87 339 88 340 
<< pdiffusion >>
rect 88 339 89 340 
<< pdiffusion >>
rect 89 339 90 340 
<< m1 >>
rect 91 339 92 340 
<< m1 >>
rect 100 339 101 340 
<< m1 >>
rect 116 339 117 340 
<< m1 >>
rect 118 339 119 340 
<< pdiffusion >>
rect 120 339 121 340 
<< pdiffusion >>
rect 121 339 122 340 
<< pdiffusion >>
rect 122 339 123 340 
<< pdiffusion >>
rect 123 339 124 340 
<< pdiffusion >>
rect 124 339 125 340 
<< pdiffusion >>
rect 125 339 126 340 
<< pdiffusion >>
rect 138 339 139 340 
<< pdiffusion >>
rect 139 339 140 340 
<< pdiffusion >>
rect 140 339 141 340 
<< pdiffusion >>
rect 141 339 142 340 
<< pdiffusion >>
rect 142 339 143 340 
<< pdiffusion >>
rect 143 339 144 340 
<< m1 >>
rect 145 339 146 340 
<< m2 >>
rect 146 339 147 340 
<< m1 >>
rect 148 339 149 340 
<< m1 >>
rect 150 339 151 340 
<< m1 >>
rect 154 339 155 340 
<< pdiffusion >>
rect 156 339 157 340 
<< pdiffusion >>
rect 157 339 158 340 
<< pdiffusion >>
rect 158 339 159 340 
<< pdiffusion >>
rect 159 339 160 340 
<< pdiffusion >>
rect 160 339 161 340 
<< pdiffusion >>
rect 161 339 162 340 
<< m1 >>
rect 163 339 164 340 
<< m2 >>
rect 164 339 165 340 
<< pdiffusion >>
rect 174 339 175 340 
<< pdiffusion >>
rect 175 339 176 340 
<< pdiffusion >>
rect 176 339 177 340 
<< pdiffusion >>
rect 177 339 178 340 
<< pdiffusion >>
rect 178 339 179 340 
<< pdiffusion >>
rect 179 339 180 340 
<< m1 >>
rect 181 339 182 340 
<< pdiffusion >>
rect 192 339 193 340 
<< pdiffusion >>
rect 193 339 194 340 
<< pdiffusion >>
rect 194 339 195 340 
<< pdiffusion >>
rect 195 339 196 340 
<< pdiffusion >>
rect 196 339 197 340 
<< pdiffusion >>
rect 197 339 198 340 
<< m1 >>
rect 204 339 205 340 
<< m1 >>
rect 206 339 207 340 
<< pdiffusion >>
rect 210 339 211 340 
<< pdiffusion >>
rect 211 339 212 340 
<< pdiffusion >>
rect 212 339 213 340 
<< pdiffusion >>
rect 213 339 214 340 
<< pdiffusion >>
rect 214 339 215 340 
<< pdiffusion >>
rect 215 339 216 340 
<< m1 >>
rect 217 339 218 340 
<< m1 >>
rect 219 339 220 340 
<< m1 >>
rect 223 339 224 340 
<< m1 >>
rect 225 339 226 340 
<< pdiffusion >>
rect 228 339 229 340 
<< pdiffusion >>
rect 229 339 230 340 
<< pdiffusion >>
rect 230 339 231 340 
<< pdiffusion >>
rect 231 339 232 340 
<< pdiffusion >>
rect 232 339 233 340 
<< pdiffusion >>
rect 233 339 234 340 
<< m1 >>
rect 235 339 236 340 
<< m1 >>
rect 242 339 243 340 
<< m1 >>
rect 244 339 245 340 
<< m2 >>
rect 244 339 245 340 
<< pdiffusion >>
rect 246 339 247 340 
<< pdiffusion >>
rect 247 339 248 340 
<< pdiffusion >>
rect 248 339 249 340 
<< pdiffusion >>
rect 249 339 250 340 
<< pdiffusion >>
rect 250 339 251 340 
<< pdiffusion >>
rect 251 339 252 340 
<< m1 >>
rect 253 339 254 340 
<< pdiffusion >>
rect 264 339 265 340 
<< pdiffusion >>
rect 265 339 266 340 
<< pdiffusion >>
rect 266 339 267 340 
<< pdiffusion >>
rect 267 339 268 340 
<< pdiffusion >>
rect 268 339 269 340 
<< pdiffusion >>
rect 269 339 270 340 
<< m1 >>
rect 276 339 277 340 
<< pdiffusion >>
rect 282 339 283 340 
<< pdiffusion >>
rect 283 339 284 340 
<< pdiffusion >>
rect 284 339 285 340 
<< pdiffusion >>
rect 285 339 286 340 
<< pdiffusion >>
rect 286 339 287 340 
<< pdiffusion >>
rect 287 339 288 340 
<< m1 >>
rect 289 339 290 340 
<< pdiffusion >>
rect 300 339 301 340 
<< pdiffusion >>
rect 301 339 302 340 
<< pdiffusion >>
rect 302 339 303 340 
<< pdiffusion >>
rect 303 339 304 340 
<< pdiffusion >>
rect 304 339 305 340 
<< pdiffusion >>
rect 305 339 306 340 
<< pdiffusion >>
rect 318 339 319 340 
<< pdiffusion >>
rect 319 339 320 340 
<< pdiffusion >>
rect 320 339 321 340 
<< pdiffusion >>
rect 321 339 322 340 
<< pdiffusion >>
rect 322 339 323 340 
<< pdiffusion >>
rect 323 339 324 340 
<< m1 >>
rect 334 339 335 340 
<< pdiffusion >>
rect 336 339 337 340 
<< pdiffusion >>
rect 337 339 338 340 
<< pdiffusion >>
rect 338 339 339 340 
<< pdiffusion >>
rect 339 339 340 340 
<< pdiffusion >>
rect 340 339 341 340 
<< pdiffusion >>
rect 341 339 342 340 
<< m1 >>
rect 347 339 348 340 
<< m2 >>
rect 350 339 351 340 
<< m1 >>
rect 351 339 352 340 
<< pdiffusion >>
rect 354 339 355 340 
<< pdiffusion >>
rect 355 339 356 340 
<< pdiffusion >>
rect 356 339 357 340 
<< pdiffusion >>
rect 357 339 358 340 
<< pdiffusion >>
rect 358 339 359 340 
<< pdiffusion >>
rect 359 339 360 340 
<< m1 >>
rect 361 339 362 340 
<< m1 >>
rect 364 339 365 340 
<< m1 >>
rect 370 339 371 340 
<< pdiffusion >>
rect 372 339 373 340 
<< pdiffusion >>
rect 373 339 374 340 
<< pdiffusion >>
rect 374 339 375 340 
<< pdiffusion >>
rect 375 339 376 340 
<< pdiffusion >>
rect 376 339 377 340 
<< pdiffusion >>
rect 377 339 378 340 
<< m1 >>
rect 379 339 380 340 
<< pdiffusion >>
rect 390 339 391 340 
<< pdiffusion >>
rect 391 339 392 340 
<< pdiffusion >>
rect 392 339 393 340 
<< pdiffusion >>
rect 393 339 394 340 
<< pdiffusion >>
rect 394 339 395 340 
<< pdiffusion >>
rect 395 339 396 340 
<< pdiffusion >>
rect 408 339 409 340 
<< pdiffusion >>
rect 409 339 410 340 
<< pdiffusion >>
rect 410 339 411 340 
<< pdiffusion >>
rect 411 339 412 340 
<< pdiffusion >>
rect 412 339 413 340 
<< pdiffusion >>
rect 413 339 414 340 
<< m1 >>
rect 416 339 417 340 
<< m1 >>
rect 418 339 419 340 
<< m2 >>
rect 421 339 422 340 
<< m1 >>
rect 422 339 423 340 
<< m1 >>
rect 424 339 425 340 
<< m2 >>
rect 424 339 425 340 
<< pdiffusion >>
rect 426 339 427 340 
<< pdiffusion >>
rect 427 339 428 340 
<< pdiffusion >>
rect 428 339 429 340 
<< pdiffusion >>
rect 429 339 430 340 
<< pdiffusion >>
rect 430 339 431 340 
<< pdiffusion >>
rect 431 339 432 340 
<< m1 >>
rect 433 339 434 340 
<< m1 >>
rect 435 339 436 340 
<< m1 >>
rect 439 339 440 340 
<< pdiffusion >>
rect 444 339 445 340 
<< pdiffusion >>
rect 445 339 446 340 
<< pdiffusion >>
rect 446 339 447 340 
<< pdiffusion >>
rect 447 339 448 340 
<< pdiffusion >>
rect 448 339 449 340 
<< pdiffusion >>
rect 449 339 450 340 
<< m1 >>
rect 451 339 452 340 
<< pdiffusion >>
rect 462 339 463 340 
<< pdiffusion >>
rect 463 339 464 340 
<< pdiffusion >>
rect 464 339 465 340 
<< pdiffusion >>
rect 465 339 466 340 
<< pdiffusion >>
rect 466 339 467 340 
<< pdiffusion >>
rect 467 339 468 340 
<< pdiffusion >>
rect 480 339 481 340 
<< pdiffusion >>
rect 481 339 482 340 
<< pdiffusion >>
rect 482 339 483 340 
<< pdiffusion >>
rect 483 339 484 340 
<< pdiffusion >>
rect 484 339 485 340 
<< pdiffusion >>
rect 485 339 486 340 
<< pdiffusion >>
rect 498 339 499 340 
<< pdiffusion >>
rect 499 339 500 340 
<< pdiffusion >>
rect 500 339 501 340 
<< pdiffusion >>
rect 501 339 502 340 
<< pdiffusion >>
rect 502 339 503 340 
<< pdiffusion >>
rect 503 339 504 340 
<< pdiffusion >>
rect 516 339 517 340 
<< pdiffusion >>
rect 517 339 518 340 
<< pdiffusion >>
rect 518 339 519 340 
<< pdiffusion >>
rect 519 339 520 340 
<< pdiffusion >>
rect 520 339 521 340 
<< pdiffusion >>
rect 521 339 522 340 
<< m1 >>
rect 523 339 524 340 
<< pdiffusion >>
rect 12 340 13 341 
<< pdiffusion >>
rect 13 340 14 341 
<< pdiffusion >>
rect 14 340 15 341 
<< pdiffusion >>
rect 15 340 16 341 
<< pdiffusion >>
rect 16 340 17 341 
<< pdiffusion >>
rect 17 340 18 341 
<< m1 >>
rect 19 340 20 341 
<< m2 >>
rect 20 340 21 341 
<< m1 >>
rect 23 340 24 341 
<< pdiffusion >>
rect 30 340 31 341 
<< pdiffusion >>
rect 31 340 32 341 
<< pdiffusion >>
rect 32 340 33 341 
<< pdiffusion >>
rect 33 340 34 341 
<< pdiffusion >>
rect 34 340 35 341 
<< pdiffusion >>
rect 35 340 36 341 
<< m1 >>
rect 44 340 45 341 
<< pdiffusion >>
rect 48 340 49 341 
<< pdiffusion >>
rect 49 340 50 341 
<< pdiffusion >>
rect 50 340 51 341 
<< pdiffusion >>
rect 51 340 52 341 
<< pdiffusion >>
rect 52 340 53 341 
<< pdiffusion >>
rect 53 340 54 341 
<< m2 >>
rect 61 340 62 341 
<< m1 >>
rect 62 340 63 341 
<< m1 >>
rect 64 340 65 341 
<< pdiffusion >>
rect 66 340 67 341 
<< pdiffusion >>
rect 67 340 68 341 
<< pdiffusion >>
rect 68 340 69 341 
<< pdiffusion >>
rect 69 340 70 341 
<< pdiffusion >>
rect 70 340 71 341 
<< pdiffusion >>
rect 71 340 72 341 
<< m1 >>
rect 73 340 74 341 
<< m1 >>
rect 82 340 83 341 
<< pdiffusion >>
rect 84 340 85 341 
<< pdiffusion >>
rect 85 340 86 341 
<< pdiffusion >>
rect 86 340 87 341 
<< pdiffusion >>
rect 87 340 88 341 
<< pdiffusion >>
rect 88 340 89 341 
<< pdiffusion >>
rect 89 340 90 341 
<< m1 >>
rect 91 340 92 341 
<< m1 >>
rect 100 340 101 341 
<< m1 >>
rect 116 340 117 341 
<< m1 >>
rect 118 340 119 341 
<< pdiffusion >>
rect 120 340 121 341 
<< pdiffusion >>
rect 121 340 122 341 
<< pdiffusion >>
rect 122 340 123 341 
<< pdiffusion >>
rect 123 340 124 341 
<< pdiffusion >>
rect 124 340 125 341 
<< pdiffusion >>
rect 125 340 126 341 
<< pdiffusion >>
rect 138 340 139 341 
<< pdiffusion >>
rect 139 340 140 341 
<< pdiffusion >>
rect 140 340 141 341 
<< pdiffusion >>
rect 141 340 142 341 
<< pdiffusion >>
rect 142 340 143 341 
<< pdiffusion >>
rect 143 340 144 341 
<< m1 >>
rect 145 340 146 341 
<< m2 >>
rect 146 340 147 341 
<< m1 >>
rect 148 340 149 341 
<< m1 >>
rect 150 340 151 341 
<< m1 >>
rect 154 340 155 341 
<< pdiffusion >>
rect 156 340 157 341 
<< pdiffusion >>
rect 157 340 158 341 
<< pdiffusion >>
rect 158 340 159 341 
<< pdiffusion >>
rect 159 340 160 341 
<< pdiffusion >>
rect 160 340 161 341 
<< pdiffusion >>
rect 161 340 162 341 
<< m1 >>
rect 163 340 164 341 
<< m2 >>
rect 164 340 165 341 
<< pdiffusion >>
rect 174 340 175 341 
<< pdiffusion >>
rect 175 340 176 341 
<< pdiffusion >>
rect 176 340 177 341 
<< pdiffusion >>
rect 177 340 178 341 
<< pdiffusion >>
rect 178 340 179 341 
<< pdiffusion >>
rect 179 340 180 341 
<< m1 >>
rect 181 340 182 341 
<< pdiffusion >>
rect 192 340 193 341 
<< pdiffusion >>
rect 193 340 194 341 
<< pdiffusion >>
rect 194 340 195 341 
<< pdiffusion >>
rect 195 340 196 341 
<< pdiffusion >>
rect 196 340 197 341 
<< pdiffusion >>
rect 197 340 198 341 
<< m1 >>
rect 204 340 205 341 
<< m1 >>
rect 206 340 207 341 
<< pdiffusion >>
rect 210 340 211 341 
<< pdiffusion >>
rect 211 340 212 341 
<< pdiffusion >>
rect 212 340 213 341 
<< pdiffusion >>
rect 213 340 214 341 
<< pdiffusion >>
rect 214 340 215 341 
<< pdiffusion >>
rect 215 340 216 341 
<< m1 >>
rect 217 340 218 341 
<< m1 >>
rect 219 340 220 341 
<< m1 >>
rect 223 340 224 341 
<< m1 >>
rect 225 340 226 341 
<< pdiffusion >>
rect 228 340 229 341 
<< pdiffusion >>
rect 229 340 230 341 
<< pdiffusion >>
rect 230 340 231 341 
<< pdiffusion >>
rect 231 340 232 341 
<< pdiffusion >>
rect 232 340 233 341 
<< pdiffusion >>
rect 233 340 234 341 
<< m1 >>
rect 235 340 236 341 
<< m1 >>
rect 242 340 243 341 
<< m1 >>
rect 244 340 245 341 
<< m2 >>
rect 244 340 245 341 
<< pdiffusion >>
rect 246 340 247 341 
<< pdiffusion >>
rect 247 340 248 341 
<< pdiffusion >>
rect 248 340 249 341 
<< pdiffusion >>
rect 249 340 250 341 
<< pdiffusion >>
rect 250 340 251 341 
<< pdiffusion >>
rect 251 340 252 341 
<< m1 >>
rect 253 340 254 341 
<< pdiffusion >>
rect 264 340 265 341 
<< pdiffusion >>
rect 265 340 266 341 
<< pdiffusion >>
rect 266 340 267 341 
<< pdiffusion >>
rect 267 340 268 341 
<< pdiffusion >>
rect 268 340 269 341 
<< pdiffusion >>
rect 269 340 270 341 
<< m1 >>
rect 276 340 277 341 
<< pdiffusion >>
rect 282 340 283 341 
<< pdiffusion >>
rect 283 340 284 341 
<< pdiffusion >>
rect 284 340 285 341 
<< pdiffusion >>
rect 285 340 286 341 
<< pdiffusion >>
rect 286 340 287 341 
<< pdiffusion >>
rect 287 340 288 341 
<< m1 >>
rect 289 340 290 341 
<< pdiffusion >>
rect 300 340 301 341 
<< pdiffusion >>
rect 301 340 302 341 
<< pdiffusion >>
rect 302 340 303 341 
<< pdiffusion >>
rect 303 340 304 341 
<< pdiffusion >>
rect 304 340 305 341 
<< pdiffusion >>
rect 305 340 306 341 
<< pdiffusion >>
rect 318 340 319 341 
<< pdiffusion >>
rect 319 340 320 341 
<< pdiffusion >>
rect 320 340 321 341 
<< pdiffusion >>
rect 321 340 322 341 
<< pdiffusion >>
rect 322 340 323 341 
<< pdiffusion >>
rect 323 340 324 341 
<< m1 >>
rect 334 340 335 341 
<< pdiffusion >>
rect 336 340 337 341 
<< pdiffusion >>
rect 337 340 338 341 
<< pdiffusion >>
rect 338 340 339 341 
<< pdiffusion >>
rect 339 340 340 341 
<< pdiffusion >>
rect 340 340 341 341 
<< pdiffusion >>
rect 341 340 342 341 
<< m1 >>
rect 347 340 348 341 
<< m2 >>
rect 350 340 351 341 
<< m1 >>
rect 351 340 352 341 
<< pdiffusion >>
rect 354 340 355 341 
<< pdiffusion >>
rect 355 340 356 341 
<< pdiffusion >>
rect 356 340 357 341 
<< pdiffusion >>
rect 357 340 358 341 
<< pdiffusion >>
rect 358 340 359 341 
<< pdiffusion >>
rect 359 340 360 341 
<< m1 >>
rect 361 340 362 341 
<< m1 >>
rect 364 340 365 341 
<< m1 >>
rect 370 340 371 341 
<< pdiffusion >>
rect 372 340 373 341 
<< pdiffusion >>
rect 373 340 374 341 
<< pdiffusion >>
rect 374 340 375 341 
<< pdiffusion >>
rect 375 340 376 341 
<< pdiffusion >>
rect 376 340 377 341 
<< pdiffusion >>
rect 377 340 378 341 
<< m1 >>
rect 379 340 380 341 
<< pdiffusion >>
rect 390 340 391 341 
<< pdiffusion >>
rect 391 340 392 341 
<< pdiffusion >>
rect 392 340 393 341 
<< pdiffusion >>
rect 393 340 394 341 
<< pdiffusion >>
rect 394 340 395 341 
<< pdiffusion >>
rect 395 340 396 341 
<< pdiffusion >>
rect 408 340 409 341 
<< pdiffusion >>
rect 409 340 410 341 
<< pdiffusion >>
rect 410 340 411 341 
<< pdiffusion >>
rect 411 340 412 341 
<< pdiffusion >>
rect 412 340 413 341 
<< pdiffusion >>
rect 413 340 414 341 
<< m1 >>
rect 416 340 417 341 
<< m1 >>
rect 418 340 419 341 
<< m2 >>
rect 421 340 422 341 
<< m1 >>
rect 422 340 423 341 
<< m1 >>
rect 424 340 425 341 
<< m2 >>
rect 424 340 425 341 
<< pdiffusion >>
rect 426 340 427 341 
<< pdiffusion >>
rect 427 340 428 341 
<< pdiffusion >>
rect 428 340 429 341 
<< pdiffusion >>
rect 429 340 430 341 
<< pdiffusion >>
rect 430 340 431 341 
<< pdiffusion >>
rect 431 340 432 341 
<< m1 >>
rect 433 340 434 341 
<< m1 >>
rect 435 340 436 341 
<< m1 >>
rect 439 340 440 341 
<< pdiffusion >>
rect 444 340 445 341 
<< pdiffusion >>
rect 445 340 446 341 
<< pdiffusion >>
rect 446 340 447 341 
<< pdiffusion >>
rect 447 340 448 341 
<< pdiffusion >>
rect 448 340 449 341 
<< pdiffusion >>
rect 449 340 450 341 
<< m1 >>
rect 451 340 452 341 
<< pdiffusion >>
rect 462 340 463 341 
<< pdiffusion >>
rect 463 340 464 341 
<< pdiffusion >>
rect 464 340 465 341 
<< pdiffusion >>
rect 465 340 466 341 
<< pdiffusion >>
rect 466 340 467 341 
<< pdiffusion >>
rect 467 340 468 341 
<< pdiffusion >>
rect 480 340 481 341 
<< pdiffusion >>
rect 481 340 482 341 
<< pdiffusion >>
rect 482 340 483 341 
<< pdiffusion >>
rect 483 340 484 341 
<< pdiffusion >>
rect 484 340 485 341 
<< pdiffusion >>
rect 485 340 486 341 
<< pdiffusion >>
rect 498 340 499 341 
<< pdiffusion >>
rect 499 340 500 341 
<< pdiffusion >>
rect 500 340 501 341 
<< pdiffusion >>
rect 501 340 502 341 
<< pdiffusion >>
rect 502 340 503 341 
<< pdiffusion >>
rect 503 340 504 341 
<< pdiffusion >>
rect 516 340 517 341 
<< pdiffusion >>
rect 517 340 518 341 
<< pdiffusion >>
rect 518 340 519 341 
<< pdiffusion >>
rect 519 340 520 341 
<< pdiffusion >>
rect 520 340 521 341 
<< pdiffusion >>
rect 521 340 522 341 
<< m1 >>
rect 523 340 524 341 
<< pdiffusion >>
rect 12 341 13 342 
<< m1 >>
rect 13 341 14 342 
<< pdiffusion >>
rect 13 341 14 342 
<< pdiffusion >>
rect 14 341 15 342 
<< pdiffusion >>
rect 15 341 16 342 
<< pdiffusion >>
rect 16 341 17 342 
<< pdiffusion >>
rect 17 341 18 342 
<< m1 >>
rect 19 341 20 342 
<< m2 >>
rect 20 341 21 342 
<< m1 >>
rect 23 341 24 342 
<< pdiffusion >>
rect 30 341 31 342 
<< pdiffusion >>
rect 31 341 32 342 
<< pdiffusion >>
rect 32 341 33 342 
<< pdiffusion >>
rect 33 341 34 342 
<< pdiffusion >>
rect 34 341 35 342 
<< pdiffusion >>
rect 35 341 36 342 
<< m1 >>
rect 44 341 45 342 
<< pdiffusion >>
rect 48 341 49 342 
<< pdiffusion >>
rect 49 341 50 342 
<< pdiffusion >>
rect 50 341 51 342 
<< pdiffusion >>
rect 51 341 52 342 
<< pdiffusion >>
rect 52 341 53 342 
<< pdiffusion >>
rect 53 341 54 342 
<< m2 >>
rect 61 341 62 342 
<< m1 >>
rect 62 341 63 342 
<< m1 >>
rect 64 341 65 342 
<< pdiffusion >>
rect 66 341 67 342 
<< m1 >>
rect 67 341 68 342 
<< pdiffusion >>
rect 67 341 68 342 
<< pdiffusion >>
rect 68 341 69 342 
<< pdiffusion >>
rect 69 341 70 342 
<< pdiffusion >>
rect 70 341 71 342 
<< pdiffusion >>
rect 71 341 72 342 
<< m1 >>
rect 73 341 74 342 
<< m1 >>
rect 82 341 83 342 
<< pdiffusion >>
rect 84 341 85 342 
<< m1 >>
rect 85 341 86 342 
<< pdiffusion >>
rect 85 341 86 342 
<< pdiffusion >>
rect 86 341 87 342 
<< pdiffusion >>
rect 87 341 88 342 
<< pdiffusion >>
rect 88 341 89 342 
<< pdiffusion >>
rect 89 341 90 342 
<< m1 >>
rect 91 341 92 342 
<< m1 >>
rect 100 341 101 342 
<< m1 >>
rect 116 341 117 342 
<< m1 >>
rect 118 341 119 342 
<< pdiffusion >>
rect 120 341 121 342 
<< pdiffusion >>
rect 121 341 122 342 
<< pdiffusion >>
rect 122 341 123 342 
<< pdiffusion >>
rect 123 341 124 342 
<< pdiffusion >>
rect 124 341 125 342 
<< pdiffusion >>
rect 125 341 126 342 
<< pdiffusion >>
rect 138 341 139 342 
<< pdiffusion >>
rect 139 341 140 342 
<< pdiffusion >>
rect 140 341 141 342 
<< pdiffusion >>
rect 141 341 142 342 
<< pdiffusion >>
rect 142 341 143 342 
<< pdiffusion >>
rect 143 341 144 342 
<< m1 >>
rect 145 341 146 342 
<< m2 >>
rect 146 341 147 342 
<< m1 >>
rect 148 341 149 342 
<< m1 >>
rect 150 341 151 342 
<< m1 >>
rect 154 341 155 342 
<< pdiffusion >>
rect 156 341 157 342 
<< pdiffusion >>
rect 157 341 158 342 
<< pdiffusion >>
rect 158 341 159 342 
<< pdiffusion >>
rect 159 341 160 342 
<< pdiffusion >>
rect 160 341 161 342 
<< pdiffusion >>
rect 161 341 162 342 
<< m1 >>
rect 163 341 164 342 
<< m2 >>
rect 164 341 165 342 
<< pdiffusion >>
rect 174 341 175 342 
<< m1 >>
rect 175 341 176 342 
<< pdiffusion >>
rect 175 341 176 342 
<< pdiffusion >>
rect 176 341 177 342 
<< pdiffusion >>
rect 177 341 178 342 
<< m1 >>
rect 178 341 179 342 
<< pdiffusion >>
rect 178 341 179 342 
<< pdiffusion >>
rect 179 341 180 342 
<< m1 >>
rect 181 341 182 342 
<< pdiffusion >>
rect 192 341 193 342 
<< m1 >>
rect 193 341 194 342 
<< pdiffusion >>
rect 193 341 194 342 
<< pdiffusion >>
rect 194 341 195 342 
<< pdiffusion >>
rect 195 341 196 342 
<< pdiffusion >>
rect 196 341 197 342 
<< pdiffusion >>
rect 197 341 198 342 
<< m1 >>
rect 204 341 205 342 
<< m1 >>
rect 206 341 207 342 
<< pdiffusion >>
rect 210 341 211 342 
<< pdiffusion >>
rect 211 341 212 342 
<< pdiffusion >>
rect 212 341 213 342 
<< pdiffusion >>
rect 213 341 214 342 
<< pdiffusion >>
rect 214 341 215 342 
<< pdiffusion >>
rect 215 341 216 342 
<< m1 >>
rect 217 341 218 342 
<< m1 >>
rect 219 341 220 342 
<< m1 >>
rect 223 341 224 342 
<< m1 >>
rect 225 341 226 342 
<< pdiffusion >>
rect 228 341 229 342 
<< pdiffusion >>
rect 229 341 230 342 
<< pdiffusion >>
rect 230 341 231 342 
<< pdiffusion >>
rect 231 341 232 342 
<< m1 >>
rect 232 341 233 342 
<< pdiffusion >>
rect 232 341 233 342 
<< pdiffusion >>
rect 233 341 234 342 
<< m1 >>
rect 235 341 236 342 
<< m1 >>
rect 242 341 243 342 
<< m1 >>
rect 244 341 245 342 
<< m2 >>
rect 244 341 245 342 
<< pdiffusion >>
rect 246 341 247 342 
<< pdiffusion >>
rect 247 341 248 342 
<< pdiffusion >>
rect 248 341 249 342 
<< pdiffusion >>
rect 249 341 250 342 
<< pdiffusion >>
rect 250 341 251 342 
<< pdiffusion >>
rect 251 341 252 342 
<< m1 >>
rect 253 341 254 342 
<< pdiffusion >>
rect 264 341 265 342 
<< m1 >>
rect 265 341 266 342 
<< pdiffusion >>
rect 265 341 266 342 
<< pdiffusion >>
rect 266 341 267 342 
<< pdiffusion >>
rect 267 341 268 342 
<< pdiffusion >>
rect 268 341 269 342 
<< pdiffusion >>
rect 269 341 270 342 
<< m1 >>
rect 276 341 277 342 
<< pdiffusion >>
rect 282 341 283 342 
<< m1 >>
rect 283 341 284 342 
<< pdiffusion >>
rect 283 341 284 342 
<< pdiffusion >>
rect 284 341 285 342 
<< pdiffusion >>
rect 285 341 286 342 
<< pdiffusion >>
rect 286 341 287 342 
<< pdiffusion >>
rect 287 341 288 342 
<< m1 >>
rect 289 341 290 342 
<< pdiffusion >>
rect 300 341 301 342 
<< pdiffusion >>
rect 301 341 302 342 
<< pdiffusion >>
rect 302 341 303 342 
<< pdiffusion >>
rect 303 341 304 342 
<< pdiffusion >>
rect 304 341 305 342 
<< pdiffusion >>
rect 305 341 306 342 
<< pdiffusion >>
rect 318 341 319 342 
<< pdiffusion >>
rect 319 341 320 342 
<< pdiffusion >>
rect 320 341 321 342 
<< pdiffusion >>
rect 321 341 322 342 
<< m1 >>
rect 322 341 323 342 
<< pdiffusion >>
rect 322 341 323 342 
<< pdiffusion >>
rect 323 341 324 342 
<< m1 >>
rect 334 341 335 342 
<< pdiffusion >>
rect 336 341 337 342 
<< m1 >>
rect 337 341 338 342 
<< pdiffusion >>
rect 337 341 338 342 
<< pdiffusion >>
rect 338 341 339 342 
<< pdiffusion >>
rect 339 341 340 342 
<< pdiffusion >>
rect 340 341 341 342 
<< pdiffusion >>
rect 341 341 342 342 
<< m1 >>
rect 347 341 348 342 
<< m2 >>
rect 350 341 351 342 
<< m1 >>
rect 351 341 352 342 
<< pdiffusion >>
rect 354 341 355 342 
<< m1 >>
rect 355 341 356 342 
<< pdiffusion >>
rect 355 341 356 342 
<< pdiffusion >>
rect 356 341 357 342 
<< pdiffusion >>
rect 357 341 358 342 
<< pdiffusion >>
rect 358 341 359 342 
<< pdiffusion >>
rect 359 341 360 342 
<< m1 >>
rect 361 341 362 342 
<< m1 >>
rect 364 341 365 342 
<< m1 >>
rect 370 341 371 342 
<< pdiffusion >>
rect 372 341 373 342 
<< m1 >>
rect 373 341 374 342 
<< pdiffusion >>
rect 373 341 374 342 
<< pdiffusion >>
rect 374 341 375 342 
<< pdiffusion >>
rect 375 341 376 342 
<< pdiffusion >>
rect 376 341 377 342 
<< pdiffusion >>
rect 377 341 378 342 
<< m1 >>
rect 379 341 380 342 
<< pdiffusion >>
rect 390 341 391 342 
<< pdiffusion >>
rect 391 341 392 342 
<< pdiffusion >>
rect 392 341 393 342 
<< pdiffusion >>
rect 393 341 394 342 
<< pdiffusion >>
rect 394 341 395 342 
<< pdiffusion >>
rect 395 341 396 342 
<< pdiffusion >>
rect 408 341 409 342 
<< pdiffusion >>
rect 409 341 410 342 
<< pdiffusion >>
rect 410 341 411 342 
<< pdiffusion >>
rect 411 341 412 342 
<< pdiffusion >>
rect 412 341 413 342 
<< pdiffusion >>
rect 413 341 414 342 
<< m1 >>
rect 416 341 417 342 
<< m1 >>
rect 418 341 419 342 
<< m2 >>
rect 421 341 422 342 
<< m1 >>
rect 422 341 423 342 
<< m1 >>
rect 424 341 425 342 
<< m2 >>
rect 424 341 425 342 
<< pdiffusion >>
rect 426 341 427 342 
<< pdiffusion >>
rect 427 341 428 342 
<< pdiffusion >>
rect 428 341 429 342 
<< pdiffusion >>
rect 429 341 430 342 
<< pdiffusion >>
rect 430 341 431 342 
<< pdiffusion >>
rect 431 341 432 342 
<< m1 >>
rect 433 341 434 342 
<< m1 >>
rect 435 341 436 342 
<< m1 >>
rect 439 341 440 342 
<< pdiffusion >>
rect 444 341 445 342 
<< pdiffusion >>
rect 445 341 446 342 
<< pdiffusion >>
rect 446 341 447 342 
<< pdiffusion >>
rect 447 341 448 342 
<< pdiffusion >>
rect 448 341 449 342 
<< pdiffusion >>
rect 449 341 450 342 
<< m1 >>
rect 451 341 452 342 
<< pdiffusion >>
rect 462 341 463 342 
<< pdiffusion >>
rect 463 341 464 342 
<< pdiffusion >>
rect 464 341 465 342 
<< pdiffusion >>
rect 465 341 466 342 
<< pdiffusion >>
rect 466 341 467 342 
<< pdiffusion >>
rect 467 341 468 342 
<< pdiffusion >>
rect 480 341 481 342 
<< pdiffusion >>
rect 481 341 482 342 
<< pdiffusion >>
rect 482 341 483 342 
<< pdiffusion >>
rect 483 341 484 342 
<< pdiffusion >>
rect 484 341 485 342 
<< pdiffusion >>
rect 485 341 486 342 
<< pdiffusion >>
rect 498 341 499 342 
<< pdiffusion >>
rect 499 341 500 342 
<< pdiffusion >>
rect 500 341 501 342 
<< pdiffusion >>
rect 501 341 502 342 
<< pdiffusion >>
rect 502 341 503 342 
<< pdiffusion >>
rect 503 341 504 342 
<< pdiffusion >>
rect 516 341 517 342 
<< pdiffusion >>
rect 517 341 518 342 
<< pdiffusion >>
rect 518 341 519 342 
<< pdiffusion >>
rect 519 341 520 342 
<< pdiffusion >>
rect 520 341 521 342 
<< pdiffusion >>
rect 521 341 522 342 
<< m1 >>
rect 523 341 524 342 
<< m1 >>
rect 13 342 14 343 
<< m1 >>
rect 19 342 20 343 
<< m2 >>
rect 20 342 21 343 
<< m1 >>
rect 23 342 24 343 
<< m1 >>
rect 44 342 45 343 
<< m2 >>
rect 61 342 62 343 
<< m1 >>
rect 62 342 63 343 
<< m1 >>
rect 64 342 65 343 
<< m1 >>
rect 67 342 68 343 
<< m1 >>
rect 73 342 74 343 
<< m1 >>
rect 82 342 83 343 
<< m1 >>
rect 85 342 86 343 
<< m1 >>
rect 91 342 92 343 
<< m1 >>
rect 100 342 101 343 
<< m1 >>
rect 116 342 117 343 
<< m1 >>
rect 118 342 119 343 
<< m1 >>
rect 145 342 146 343 
<< m2 >>
rect 146 342 147 343 
<< m1 >>
rect 148 342 149 343 
<< m1 >>
rect 150 342 151 343 
<< m1 >>
rect 154 342 155 343 
<< m1 >>
rect 163 342 164 343 
<< m2 >>
rect 164 342 165 343 
<< m1 >>
rect 175 342 176 343 
<< m1 >>
rect 178 342 179 343 
<< m1 >>
rect 181 342 182 343 
<< m1 >>
rect 193 342 194 343 
<< m1 >>
rect 204 342 205 343 
<< m1 >>
rect 206 342 207 343 
<< m1 >>
rect 217 342 218 343 
<< m1 >>
rect 219 342 220 343 
<< m1 >>
rect 223 342 224 343 
<< m1 >>
rect 225 342 226 343 
<< m1 >>
rect 232 342 233 343 
<< m1 >>
rect 235 342 236 343 
<< m1 >>
rect 242 342 243 343 
<< m1 >>
rect 244 342 245 343 
<< m2 >>
rect 244 342 245 343 
<< m1 >>
rect 253 342 254 343 
<< m1 >>
rect 265 342 266 343 
<< m1 >>
rect 276 342 277 343 
<< m1 >>
rect 283 342 284 343 
<< m1 >>
rect 289 342 290 343 
<< m1 >>
rect 322 342 323 343 
<< m1 >>
rect 334 342 335 343 
<< m1 >>
rect 337 342 338 343 
<< m1 >>
rect 347 342 348 343 
<< m2 >>
rect 350 342 351 343 
<< m1 >>
rect 351 342 352 343 
<< m1 >>
rect 355 342 356 343 
<< m1 >>
rect 361 342 362 343 
<< m2 >>
rect 361 342 362 343 
<< m2c >>
rect 361 342 362 343 
<< m1 >>
rect 361 342 362 343 
<< m2 >>
rect 361 342 362 343 
<< m1 >>
rect 364 342 365 343 
<< m1 >>
rect 365 342 366 343 
<< m1 >>
rect 366 342 367 343 
<< m1 >>
rect 367 342 368 343 
<< m1 >>
rect 368 342 369 343 
<< m2 >>
rect 368 342 369 343 
<< m2c >>
rect 368 342 369 343 
<< m1 >>
rect 368 342 369 343 
<< m2 >>
rect 368 342 369 343 
<< m2 >>
rect 369 342 370 343 
<< m1 >>
rect 370 342 371 343 
<< m2 >>
rect 370 342 371 343 
<< m1 >>
rect 373 342 374 343 
<< m1 >>
rect 379 342 380 343 
<< m1 >>
rect 416 342 417 343 
<< m1 >>
rect 418 342 419 343 
<< m2 >>
rect 421 342 422 343 
<< m1 >>
rect 422 342 423 343 
<< m1 >>
rect 424 342 425 343 
<< m2 >>
rect 424 342 425 343 
<< m1 >>
rect 433 342 434 343 
<< m1 >>
rect 435 342 436 343 
<< m1 >>
rect 439 342 440 343 
<< m1 >>
rect 451 342 452 343 
<< m1 >>
rect 523 342 524 343 
<< m1 >>
rect 13 343 14 344 
<< m1 >>
rect 17 343 18 344 
<< m2 >>
rect 17 343 18 344 
<< m2c >>
rect 17 343 18 344 
<< m1 >>
rect 17 343 18 344 
<< m2 >>
rect 17 343 18 344 
<< m2 >>
rect 18 343 19 344 
<< m1 >>
rect 19 343 20 344 
<< m2 >>
rect 19 343 20 344 
<< m2 >>
rect 20 343 21 344 
<< m1 >>
rect 23 343 24 344 
<< m1 >>
rect 44 343 45 344 
<< m2 >>
rect 61 343 62 344 
<< m1 >>
rect 62 343 63 344 
<< m1 >>
rect 64 343 65 344 
<< m1 >>
rect 67 343 68 344 
<< m1 >>
rect 73 343 74 344 
<< m1 >>
rect 82 343 83 344 
<< m1 >>
rect 85 343 86 344 
<< m1 >>
rect 91 343 92 344 
<< m1 >>
rect 100 343 101 344 
<< m1 >>
rect 116 343 117 344 
<< m1 >>
rect 118 343 119 344 
<< m1 >>
rect 144 343 145 344 
<< m1 >>
rect 145 343 146 344 
<< m2 >>
rect 146 343 147 344 
<< m1 >>
rect 148 343 149 344 
<< m1 >>
rect 150 343 151 344 
<< m1 >>
rect 154 343 155 344 
<< m1 >>
rect 163 343 164 344 
<< m2 >>
rect 164 343 165 344 
<< m1 >>
rect 175 343 176 344 
<< m1 >>
rect 178 343 179 344 
<< m1 >>
rect 179 343 180 344 
<< m1 >>
rect 180 343 181 344 
<< m1 >>
rect 181 343 182 344 
<< m1 >>
rect 193 343 194 344 
<< m1 >>
rect 204 343 205 344 
<< m1 >>
rect 206 343 207 344 
<< m1 >>
rect 217 343 218 344 
<< m1 >>
rect 219 343 220 344 
<< m1 >>
rect 223 343 224 344 
<< m1 >>
rect 225 343 226 344 
<< m1 >>
rect 232 343 233 344 
<< m1 >>
rect 235 343 236 344 
<< m1 >>
rect 242 343 243 344 
<< m1 >>
rect 244 343 245 344 
<< m2 >>
rect 244 343 245 344 
<< m1 >>
rect 253 343 254 344 
<< m1 >>
rect 265 343 266 344 
<< m1 >>
rect 276 343 277 344 
<< m1 >>
rect 283 343 284 344 
<< m1 >>
rect 289 343 290 344 
<< m1 >>
rect 322 343 323 344 
<< m1 >>
rect 334 343 335 344 
<< m1 >>
rect 335 343 336 344 
<< m1 >>
rect 336 343 337 344 
<< m1 >>
rect 337 343 338 344 
<< m1 >>
rect 347 343 348 344 
<< m2 >>
rect 350 343 351 344 
<< m1 >>
rect 351 343 352 344 
<< m1 >>
rect 355 343 356 344 
<< m2 >>
rect 361 343 362 344 
<< m1 >>
rect 370 343 371 344 
<< m2 >>
rect 370 343 371 344 
<< m2 >>
rect 371 343 372 344 
<< m1 >>
rect 372 343 373 344 
<< m2 >>
rect 372 343 373 344 
<< m2c >>
rect 372 343 373 344 
<< m1 >>
rect 372 343 373 344 
<< m2 >>
rect 372 343 373 344 
<< m1 >>
rect 373 343 374 344 
<< m1 >>
rect 379 343 380 344 
<< m1 >>
rect 416 343 417 344 
<< m1 >>
rect 418 343 419 344 
<< m2 >>
rect 421 343 422 344 
<< m1 >>
rect 422 343 423 344 
<< m1 >>
rect 424 343 425 344 
<< m2 >>
rect 424 343 425 344 
<< m2 >>
rect 425 343 426 344 
<< m1 >>
rect 426 343 427 344 
<< m2 >>
rect 426 343 427 344 
<< m2c >>
rect 426 343 427 344 
<< m1 >>
rect 426 343 427 344 
<< m2 >>
rect 426 343 427 344 
<< m1 >>
rect 433 343 434 344 
<< m1 >>
rect 435 343 436 344 
<< m1 >>
rect 439 343 440 344 
<< m1 >>
rect 451 343 452 344 
<< m1 >>
rect 523 343 524 344 
<< m1 >>
rect 13 344 14 345 
<< m1 >>
rect 14 344 15 345 
<< m1 >>
rect 15 344 16 345 
<< m1 >>
rect 16 344 17 345 
<< m1 >>
rect 17 344 18 345 
<< m1 >>
rect 19 344 20 345 
<< m1 >>
rect 23 344 24 345 
<< m1 >>
rect 44 344 45 345 
<< m2 >>
rect 61 344 62 345 
<< m1 >>
rect 62 344 63 345 
<< m1 >>
rect 64 344 65 345 
<< m1 >>
rect 67 344 68 345 
<< m1 >>
rect 73 344 74 345 
<< m1 >>
rect 82 344 83 345 
<< m1 >>
rect 85 344 86 345 
<< m1 >>
rect 86 344 87 345 
<< m1 >>
rect 87 344 88 345 
<< m1 >>
rect 88 344 89 345 
<< m1 >>
rect 89 344 90 345 
<< m1 >>
rect 90 344 91 345 
<< m1 >>
rect 91 344 92 345 
<< m1 >>
rect 100 344 101 345 
<< m1 >>
rect 116 344 117 345 
<< m1 >>
rect 118 344 119 345 
<< m1 >>
rect 142 344 143 345 
<< m2 >>
rect 142 344 143 345 
<< m2c >>
rect 142 344 143 345 
<< m1 >>
rect 142 344 143 345 
<< m2 >>
rect 142 344 143 345 
<< m2 >>
rect 143 344 144 345 
<< m1 >>
rect 144 344 145 345 
<< m2 >>
rect 144 344 145 345 
<< m2 >>
rect 145 344 146 345 
<< m2 >>
rect 146 344 147 345 
<< m1 >>
rect 148 344 149 345 
<< m1 >>
rect 150 344 151 345 
<< m1 >>
rect 154 344 155 345 
<< m1 >>
rect 163 344 164 345 
<< m2 >>
rect 164 344 165 345 
<< m1 >>
rect 175 344 176 345 
<< m1 >>
rect 193 344 194 345 
<< m1 >>
rect 194 344 195 345 
<< m1 >>
rect 195 344 196 345 
<< m1 >>
rect 196 344 197 345 
<< m1 >>
rect 197 344 198 345 
<< m1 >>
rect 198 344 199 345 
<< m1 >>
rect 199 344 200 345 
<< m1 >>
rect 200 344 201 345 
<< m1 >>
rect 201 344 202 345 
<< m1 >>
rect 202 344 203 345 
<< m1 >>
rect 203 344 204 345 
<< m1 >>
rect 204 344 205 345 
<< m1 >>
rect 206 344 207 345 
<< m1 >>
rect 217 344 218 345 
<< m2 >>
rect 217 344 218 345 
<< m2c >>
rect 217 344 218 345 
<< m1 >>
rect 217 344 218 345 
<< m2 >>
rect 217 344 218 345 
<< m1 >>
rect 219 344 220 345 
<< m2 >>
rect 219 344 220 345 
<< m2c >>
rect 219 344 220 345 
<< m1 >>
rect 219 344 220 345 
<< m2 >>
rect 219 344 220 345 
<< m1 >>
rect 221 344 222 345 
<< m2 >>
rect 221 344 222 345 
<< m2c >>
rect 221 344 222 345 
<< m1 >>
rect 221 344 222 345 
<< m2 >>
rect 221 344 222 345 
<< m1 >>
rect 222 344 223 345 
<< m1 >>
rect 223 344 224 345 
<< m2 >>
rect 223 344 224 345 
<< m2 >>
rect 224 344 225 345 
<< m1 >>
rect 225 344 226 345 
<< m2 >>
rect 225 344 226 345 
<< m2c >>
rect 225 344 226 345 
<< m1 >>
rect 225 344 226 345 
<< m2 >>
rect 225 344 226 345 
<< m1 >>
rect 232 344 233 345 
<< m1 >>
rect 235 344 236 345 
<< m1 >>
rect 242 344 243 345 
<< m1 >>
rect 244 344 245 345 
<< m2 >>
rect 244 344 245 345 
<< m1 >>
rect 253 344 254 345 
<< m1 >>
rect 265 344 266 345 
<< m1 >>
rect 276 344 277 345 
<< m1 >>
rect 283 344 284 345 
<< m1 >>
rect 284 344 285 345 
<< m1 >>
rect 285 344 286 345 
<< m1 >>
rect 286 344 287 345 
<< m1 >>
rect 287 344 288 345 
<< m1 >>
rect 288 344 289 345 
<< m1 >>
rect 289 344 290 345 
<< m1 >>
rect 322 344 323 345 
<< m1 >>
rect 347 344 348 345 
<< m2 >>
rect 350 344 351 345 
<< m1 >>
rect 351 344 352 345 
<< m1 >>
rect 355 344 356 345 
<< m1 >>
rect 356 344 357 345 
<< m1 >>
rect 357 344 358 345 
<< m1 >>
rect 358 344 359 345 
<< m1 >>
rect 359 344 360 345 
<< m1 >>
rect 360 344 361 345 
<< m1 >>
rect 361 344 362 345 
<< m2 >>
rect 361 344 362 345 
<< m1 >>
rect 362 344 363 345 
<< m1 >>
rect 363 344 364 345 
<< m1 >>
rect 364 344 365 345 
<< m1 >>
rect 365 344 366 345 
<< m1 >>
rect 366 344 367 345 
<< m1 >>
rect 367 344 368 345 
<< m1 >>
rect 368 344 369 345 
<< m1 >>
rect 369 344 370 345 
<< m1 >>
rect 370 344 371 345 
<< m1 >>
rect 379 344 380 345 
<< m2 >>
rect 379 344 380 345 
<< m2c >>
rect 379 344 380 345 
<< m1 >>
rect 379 344 380 345 
<< m2 >>
rect 379 344 380 345 
<< m1 >>
rect 416 344 417 345 
<< m1 >>
rect 418 344 419 345 
<< m2 >>
rect 421 344 422 345 
<< m1 >>
rect 422 344 423 345 
<< m1 >>
rect 424 344 425 345 
<< m1 >>
rect 426 344 427 345 
<< m1 >>
rect 433 344 434 345 
<< m1 >>
rect 435 344 436 345 
<< m1 >>
rect 439 344 440 345 
<< m1 >>
rect 451 344 452 345 
<< m1 >>
rect 523 344 524 345 
<< m1 >>
rect 19 345 20 346 
<< m1 >>
rect 23 345 24 346 
<< m1 >>
rect 44 345 45 346 
<< m2 >>
rect 61 345 62 346 
<< m1 >>
rect 62 345 63 346 
<< m1 >>
rect 64 345 65 346 
<< m1 >>
rect 67 345 68 346 
<< m1 >>
rect 73 345 74 346 
<< m1 >>
rect 82 345 83 346 
<< m1 >>
rect 100 345 101 346 
<< m1 >>
rect 116 345 117 346 
<< m1 >>
rect 118 345 119 346 
<< m1 >>
rect 142 345 143 346 
<< m1 >>
rect 144 345 145 346 
<< m1 >>
rect 148 345 149 346 
<< m1 >>
rect 150 345 151 346 
<< m1 >>
rect 154 345 155 346 
<< m1 >>
rect 163 345 164 346 
<< m2 >>
rect 164 345 165 346 
<< m1 >>
rect 175 345 176 346 
<< m1 >>
rect 176 345 177 346 
<< m1 >>
rect 177 345 178 346 
<< m1 >>
rect 178 345 179 346 
<< m1 >>
rect 179 345 180 346 
<< m1 >>
rect 180 345 181 346 
<< m1 >>
rect 181 345 182 346 
<< m1 >>
rect 182 345 183 346 
<< m2 >>
rect 182 345 183 346 
<< m2c >>
rect 182 345 183 346 
<< m1 >>
rect 182 345 183 346 
<< m2 >>
rect 182 345 183 346 
<< m1 >>
rect 206 345 207 346 
<< m2 >>
rect 217 345 218 346 
<< m2 >>
rect 219 345 220 346 
<< m2 >>
rect 221 345 222 346 
<< m2 >>
rect 223 345 224 346 
<< m1 >>
rect 232 345 233 346 
<< m1 >>
rect 235 345 236 346 
<< m1 >>
rect 242 345 243 346 
<< m1 >>
rect 244 345 245 346 
<< m2 >>
rect 244 345 245 346 
<< m1 >>
rect 253 345 254 346 
<< m1 >>
rect 265 345 266 346 
<< m1 >>
rect 276 345 277 346 
<< m1 >>
rect 322 345 323 346 
<< m1 >>
rect 347 345 348 346 
<< m2 >>
rect 350 345 351 346 
<< m1 >>
rect 351 345 352 346 
<< m2 >>
rect 361 345 362 346 
<< m2 >>
rect 379 345 380 346 
<< m1 >>
rect 416 345 417 346 
<< m1 >>
rect 418 345 419 346 
<< m2 >>
rect 421 345 422 346 
<< m1 >>
rect 422 345 423 346 
<< m1 >>
rect 424 345 425 346 
<< m1 >>
rect 426 345 427 346 
<< m1 >>
rect 433 345 434 346 
<< m1 >>
rect 435 345 436 346 
<< m1 >>
rect 439 345 440 346 
<< m1 >>
rect 451 345 452 346 
<< m1 >>
rect 523 345 524 346 
<< m1 >>
rect 19 346 20 347 
<< m1 >>
rect 23 346 24 347 
<< m1 >>
rect 44 346 45 347 
<< m2 >>
rect 61 346 62 347 
<< m1 >>
rect 62 346 63 347 
<< m2 >>
rect 62 346 63 347 
<< m2 >>
rect 63 346 64 347 
<< m1 >>
rect 64 346 65 347 
<< m2 >>
rect 64 346 65 347 
<< m2 >>
rect 65 346 66 347 
<< m2 >>
rect 66 346 67 347 
<< m1 >>
rect 67 346 68 347 
<< m2 >>
rect 67 346 68 347 
<< m2 >>
rect 68 346 69 347 
<< m1 >>
rect 69 346 70 347 
<< m2 >>
rect 69 346 70 347 
<< m2c >>
rect 69 346 70 347 
<< m1 >>
rect 69 346 70 347 
<< m2 >>
rect 69 346 70 347 
<< m1 >>
rect 70 346 71 347 
<< m1 >>
rect 71 346 72 347 
<< m2 >>
rect 71 346 72 347 
<< m2c >>
rect 71 346 72 347 
<< m1 >>
rect 71 346 72 347 
<< m2 >>
rect 71 346 72 347 
<< m2 >>
rect 72 346 73 347 
<< m1 >>
rect 73 346 74 347 
<< m2 >>
rect 73 346 74 347 
<< m2 >>
rect 74 346 75 347 
<< m1 >>
rect 75 346 76 347 
<< m2 >>
rect 75 346 76 347 
<< m2c >>
rect 75 346 76 347 
<< m1 >>
rect 75 346 76 347 
<< m2 >>
rect 75 346 76 347 
<< m1 >>
rect 76 346 77 347 
<< m1 >>
rect 77 346 78 347 
<< m1 >>
rect 78 346 79 347 
<< m1 >>
rect 79 346 80 347 
<< m1 >>
rect 80 346 81 347 
<< m2 >>
rect 80 346 81 347 
<< m2c >>
rect 80 346 81 347 
<< m1 >>
rect 80 346 81 347 
<< m2 >>
rect 80 346 81 347 
<< m2 >>
rect 81 346 82 347 
<< m1 >>
rect 82 346 83 347 
<< m2 >>
rect 82 346 83 347 
<< m2 >>
rect 83 346 84 347 
<< m1 >>
rect 84 346 85 347 
<< m2 >>
rect 84 346 85 347 
<< m2c >>
rect 84 346 85 347 
<< m1 >>
rect 84 346 85 347 
<< m2 >>
rect 84 346 85 347 
<< m1 >>
rect 85 346 86 347 
<< m1 >>
rect 86 346 87 347 
<< m1 >>
rect 87 346 88 347 
<< m1 >>
rect 88 346 89 347 
<< m1 >>
rect 89 346 90 347 
<< m1 >>
rect 90 346 91 347 
<< m1 >>
rect 91 346 92 347 
<< m1 >>
rect 100 346 101 347 
<< m1 >>
rect 112 346 113 347 
<< m1 >>
rect 113 346 114 347 
<< m1 >>
rect 114 346 115 347 
<< m2 >>
rect 114 346 115 347 
<< m2c >>
rect 114 346 115 347 
<< m1 >>
rect 114 346 115 347 
<< m2 >>
rect 114 346 115 347 
<< m2 >>
rect 115 346 116 347 
<< m1 >>
rect 116 346 117 347 
<< m2 >>
rect 116 346 117 347 
<< m2 >>
rect 117 346 118 347 
<< m1 >>
rect 118 346 119 347 
<< m2 >>
rect 118 346 119 347 
<< m2 >>
rect 119 346 120 347 
<< m1 >>
rect 120 346 121 347 
<< m2 >>
rect 120 346 121 347 
<< m2c >>
rect 120 346 121 347 
<< m1 >>
rect 120 346 121 347 
<< m2 >>
rect 120 346 121 347 
<< m1 >>
rect 121 346 122 347 
<< m1 >>
rect 122 346 123 347 
<< m1 >>
rect 123 346 124 347 
<< m1 >>
rect 124 346 125 347 
<< m1 >>
rect 125 346 126 347 
<< m1 >>
rect 126 346 127 347 
<< m1 >>
rect 127 346 128 347 
<< m1 >>
rect 128 346 129 347 
<< m1 >>
rect 129 346 130 347 
<< m1 >>
rect 130 346 131 347 
<< m1 >>
rect 131 346 132 347 
<< m1 >>
rect 132 346 133 347 
<< m1 >>
rect 133 346 134 347 
<< m1 >>
rect 134 346 135 347 
<< m1 >>
rect 135 346 136 347 
<< m1 >>
rect 136 346 137 347 
<< m1 >>
rect 137 346 138 347 
<< m1 >>
rect 138 346 139 347 
<< m1 >>
rect 139 346 140 347 
<< m1 >>
rect 140 346 141 347 
<< m1 >>
rect 141 346 142 347 
<< m1 >>
rect 142 346 143 347 
<< m1 >>
rect 144 346 145 347 
<< m1 >>
rect 148 346 149 347 
<< m1 >>
rect 150 346 151 347 
<< m1 >>
rect 154 346 155 347 
<< m1 >>
rect 163 346 164 347 
<< m2 >>
rect 164 346 165 347 
<< m1 >>
rect 165 346 166 347 
<< m2 >>
rect 165 346 166 347 
<< m2c >>
rect 165 346 166 347 
<< m1 >>
rect 165 346 166 347 
<< m2 >>
rect 165 346 166 347 
<< m1 >>
rect 166 346 167 347 
<< m1 >>
rect 167 346 168 347 
<< m1 >>
rect 168 346 169 347 
<< m2 >>
rect 168 346 169 347 
<< m2c >>
rect 168 346 169 347 
<< m1 >>
rect 168 346 169 347 
<< m2 >>
rect 168 346 169 347 
<< m2 >>
rect 182 346 183 347 
<< m1 >>
rect 206 346 207 347 
<< m1 >>
rect 208 346 209 347 
<< m1 >>
rect 209 346 210 347 
<< m1 >>
rect 210 346 211 347 
<< m1 >>
rect 211 346 212 347 
<< m1 >>
rect 212 346 213 347 
<< m1 >>
rect 213 346 214 347 
<< m1 >>
rect 214 346 215 347 
<< m1 >>
rect 215 346 216 347 
<< m1 >>
rect 216 346 217 347 
<< m1 >>
rect 217 346 218 347 
<< m2 >>
rect 217 346 218 347 
<< m1 >>
rect 218 346 219 347 
<< m1 >>
rect 219 346 220 347 
<< m2 >>
rect 219 346 220 347 
<< m1 >>
rect 220 346 221 347 
<< m1 >>
rect 221 346 222 347 
<< m2 >>
rect 221 346 222 347 
<< m1 >>
rect 222 346 223 347 
<< m1 >>
rect 223 346 224 347 
<< m2 >>
rect 223 346 224 347 
<< m1 >>
rect 224 346 225 347 
<< m1 >>
rect 225 346 226 347 
<< m1 >>
rect 226 346 227 347 
<< m1 >>
rect 227 346 228 347 
<< m1 >>
rect 228 346 229 347 
<< m1 >>
rect 229 346 230 347 
<< m1 >>
rect 230 346 231 347 
<< m1 >>
rect 231 346 232 347 
<< m1 >>
rect 232 346 233 347 
<< m1 >>
rect 235 346 236 347 
<< m1 >>
rect 242 346 243 347 
<< m1 >>
rect 244 346 245 347 
<< m2 >>
rect 244 346 245 347 
<< m1 >>
rect 253 346 254 347 
<< m1 >>
rect 265 346 266 347 
<< m1 >>
rect 276 346 277 347 
<< m1 >>
rect 277 346 278 347 
<< m1 >>
rect 278 346 279 347 
<< m1 >>
rect 279 346 280 347 
<< m1 >>
rect 280 346 281 347 
<< m1 >>
rect 281 346 282 347 
<< m1 >>
rect 282 346 283 347 
<< m1 >>
rect 283 346 284 347 
<< m1 >>
rect 284 346 285 347 
<< m1 >>
rect 285 346 286 347 
<< m1 >>
rect 286 346 287 347 
<< m1 >>
rect 287 346 288 347 
<< m1 >>
rect 288 346 289 347 
<< m1 >>
rect 289 346 290 347 
<< m1 >>
rect 290 346 291 347 
<< m1 >>
rect 291 346 292 347 
<< m1 >>
rect 292 346 293 347 
<< m1 >>
rect 293 346 294 347 
<< m1 >>
rect 294 346 295 347 
<< m1 >>
rect 295 346 296 347 
<< m1 >>
rect 296 346 297 347 
<< m1 >>
rect 297 346 298 347 
<< m1 >>
rect 298 346 299 347 
<< m1 >>
rect 299 346 300 347 
<< m1 >>
rect 300 346 301 347 
<< m1 >>
rect 301 346 302 347 
<< m1 >>
rect 302 346 303 347 
<< m1 >>
rect 303 346 304 347 
<< m1 >>
rect 304 346 305 347 
<< m1 >>
rect 305 346 306 347 
<< m1 >>
rect 306 346 307 347 
<< m1 >>
rect 307 346 308 347 
<< m1 >>
rect 308 346 309 347 
<< m1 >>
rect 309 346 310 347 
<< m1 >>
rect 310 346 311 347 
<< m1 >>
rect 311 346 312 347 
<< m1 >>
rect 312 346 313 347 
<< m1 >>
rect 313 346 314 347 
<< m1 >>
rect 314 346 315 347 
<< m2 >>
rect 314 346 315 347 
<< m2c >>
rect 314 346 315 347 
<< m1 >>
rect 314 346 315 347 
<< m2 >>
rect 314 346 315 347 
<< m2 >>
rect 315 346 316 347 
<< m1 >>
rect 316 346 317 347 
<< m2 >>
rect 316 346 317 347 
<< m1 >>
rect 317 346 318 347 
<< m2 >>
rect 317 346 318 347 
<< m1 >>
rect 318 346 319 347 
<< m2 >>
rect 318 346 319 347 
<< m1 >>
rect 319 346 320 347 
<< m2 >>
rect 319 346 320 347 
<< m1 >>
rect 320 346 321 347 
<< m2 >>
rect 320 346 321 347 
<< m1 >>
rect 321 346 322 347 
<< m2 >>
rect 321 346 322 347 
<< m1 >>
rect 322 346 323 347 
<< m1 >>
rect 347 346 348 347 
<< m2 >>
rect 350 346 351 347 
<< m1 >>
rect 351 346 352 347 
<< m1 >>
rect 361 346 362 347 
<< m2 >>
rect 361 346 362 347 
<< m2c >>
rect 361 346 362 347 
<< m1 >>
rect 361 346 362 347 
<< m2 >>
rect 361 346 362 347 
<< m1 >>
rect 362 346 363 347 
<< m1 >>
rect 363 346 364 347 
<< m1 >>
rect 364 346 365 347 
<< m1 >>
rect 365 346 366 347 
<< m1 >>
rect 366 346 367 347 
<< m1 >>
rect 367 346 368 347 
<< m1 >>
rect 368 346 369 347 
<< m1 >>
rect 369 346 370 347 
<< m1 >>
rect 370 346 371 347 
<< m1 >>
rect 371 346 372 347 
<< m1 >>
rect 372 346 373 347 
<< m1 >>
rect 373 346 374 347 
<< m1 >>
rect 374 346 375 347 
<< m1 >>
rect 375 346 376 347 
<< m1 >>
rect 376 346 377 347 
<< m1 >>
rect 377 346 378 347 
<< m1 >>
rect 378 346 379 347 
<< m1 >>
rect 379 346 380 347 
<< m2 >>
rect 379 346 380 347 
<< m1 >>
rect 380 346 381 347 
<< m1 >>
rect 381 346 382 347 
<< m1 >>
rect 382 346 383 347 
<< m1 >>
rect 383 346 384 347 
<< m1 >>
rect 384 346 385 347 
<< m1 >>
rect 385 346 386 347 
<< m1 >>
rect 386 346 387 347 
<< m1 >>
rect 387 346 388 347 
<< m1 >>
rect 388 346 389 347 
<< m1 >>
rect 389 346 390 347 
<< m1 >>
rect 390 346 391 347 
<< m1 >>
rect 391 346 392 347 
<< m1 >>
rect 392 346 393 347 
<< m1 >>
rect 393 346 394 347 
<< m1 >>
rect 416 346 417 347 
<< m1 >>
rect 418 346 419 347 
<< m2 >>
rect 421 346 422 347 
<< m1 >>
rect 422 346 423 347 
<< m1 >>
rect 424 346 425 347 
<< m1 >>
rect 426 346 427 347 
<< m1 >>
rect 427 346 428 347 
<< m1 >>
rect 428 346 429 347 
<< m1 >>
rect 429 346 430 347 
<< m1 >>
rect 430 346 431 347 
<< m1 >>
rect 431 346 432 347 
<< m2 >>
rect 431 346 432 347 
<< m2c >>
rect 431 346 432 347 
<< m1 >>
rect 431 346 432 347 
<< m2 >>
rect 431 346 432 347 
<< m2 >>
rect 432 346 433 347 
<< m1 >>
rect 433 346 434 347 
<< m2 >>
rect 433 346 434 347 
<< m2 >>
rect 434 346 435 347 
<< m1 >>
rect 435 346 436 347 
<< m2 >>
rect 435 346 436 347 
<< m2 >>
rect 436 346 437 347 
<< m1 >>
rect 437 346 438 347 
<< m2 >>
rect 437 346 438 347 
<< m2c >>
rect 437 346 438 347 
<< m1 >>
rect 437 346 438 347 
<< m2 >>
rect 437 346 438 347 
<< m1 >>
rect 439 346 440 347 
<< m1 >>
rect 451 346 452 347 
<< m1 >>
rect 523 346 524 347 
<< m1 >>
rect 19 347 20 348 
<< m1 >>
rect 23 347 24 348 
<< m1 >>
rect 44 347 45 348 
<< m1 >>
rect 62 347 63 348 
<< m1 >>
rect 64 347 65 348 
<< m1 >>
rect 67 347 68 348 
<< m1 >>
rect 73 347 74 348 
<< m1 >>
rect 82 347 83 348 
<< m1 >>
rect 91 347 92 348 
<< m1 >>
rect 100 347 101 348 
<< m1 >>
rect 112 347 113 348 
<< m2 >>
rect 112 347 113 348 
<< m2c >>
rect 112 347 113 348 
<< m1 >>
rect 112 347 113 348 
<< m2 >>
rect 112 347 113 348 
<< m1 >>
rect 116 347 117 348 
<< m1 >>
rect 118 347 119 348 
<< m1 >>
rect 144 347 145 348 
<< m2 >>
rect 144 347 145 348 
<< m2c >>
rect 144 347 145 348 
<< m1 >>
rect 144 347 145 348 
<< m2 >>
rect 144 347 145 348 
<< m1 >>
rect 148 347 149 348 
<< m1 >>
rect 150 347 151 348 
<< m1 >>
rect 154 347 155 348 
<< m1 >>
rect 163 347 164 348 
<< m2 >>
rect 168 347 169 348 
<< m2 >>
rect 174 347 175 348 
<< m2 >>
rect 175 347 176 348 
<< m2 >>
rect 176 347 177 348 
<< m2 >>
rect 177 347 178 348 
<< m2 >>
rect 178 347 179 348 
<< m2 >>
rect 179 347 180 348 
<< m1 >>
rect 180 347 181 348 
<< m2 >>
rect 180 347 181 348 
<< m2c >>
rect 180 347 181 348 
<< m1 >>
rect 180 347 181 348 
<< m2 >>
rect 180 347 181 348 
<< m1 >>
rect 181 347 182 348 
<< m1 >>
rect 182 347 183 348 
<< m2 >>
rect 182 347 183 348 
<< m1 >>
rect 183 347 184 348 
<< m1 >>
rect 184 347 185 348 
<< m1 >>
rect 185 347 186 348 
<< m1 >>
rect 186 347 187 348 
<< m1 >>
rect 187 347 188 348 
<< m1 >>
rect 188 347 189 348 
<< m1 >>
rect 189 347 190 348 
<< m1 >>
rect 190 347 191 348 
<< m1 >>
rect 191 347 192 348 
<< m1 >>
rect 192 347 193 348 
<< m1 >>
rect 193 347 194 348 
<< m1 >>
rect 194 347 195 348 
<< m1 >>
rect 195 347 196 348 
<< m1 >>
rect 196 347 197 348 
<< m1 >>
rect 197 347 198 348 
<< m1 >>
rect 198 347 199 348 
<< m1 >>
rect 199 347 200 348 
<< m1 >>
rect 200 347 201 348 
<< m1 >>
rect 201 347 202 348 
<< m1 >>
rect 202 347 203 348 
<< m1 >>
rect 203 347 204 348 
<< m1 >>
rect 204 347 205 348 
<< m1 >>
rect 205 347 206 348 
<< m1 >>
rect 206 347 207 348 
<< m1 >>
rect 208 347 209 348 
<< m2 >>
rect 217 347 218 348 
<< m2 >>
rect 219 347 220 348 
<< m2 >>
rect 221 347 222 348 
<< m2 >>
rect 223 347 224 348 
<< m1 >>
rect 235 347 236 348 
<< m1 >>
rect 242 347 243 348 
<< m1 >>
rect 244 347 245 348 
<< m2 >>
rect 244 347 245 348 
<< m1 >>
rect 253 347 254 348 
<< m1 >>
rect 265 347 266 348 
<< m1 >>
rect 316 347 317 348 
<< m2 >>
rect 321 347 322 348 
<< m1 >>
rect 347 347 348 348 
<< m2 >>
rect 347 347 348 348 
<< m2c >>
rect 347 347 348 348 
<< m1 >>
rect 347 347 348 348 
<< m2 >>
rect 347 347 348 348 
<< m2 >>
rect 350 347 351 348 
<< m1 >>
rect 351 347 352 348 
<< m2 >>
rect 379 347 380 348 
<< m1 >>
rect 393 347 394 348 
<< m2 >>
rect 393 347 394 348 
<< m2c >>
rect 393 347 394 348 
<< m1 >>
rect 393 347 394 348 
<< m2 >>
rect 393 347 394 348 
<< m1 >>
rect 416 347 417 348 
<< m1 >>
rect 418 347 419 348 
<< m2 >>
rect 421 347 422 348 
<< m1 >>
rect 422 347 423 348 
<< m1 >>
rect 424 347 425 348 
<< m1 >>
rect 433 347 434 348 
<< m1 >>
rect 435 347 436 348 
<< m1 >>
rect 437 347 438 348 
<< m1 >>
rect 439 347 440 348 
<< m1 >>
rect 451 347 452 348 
<< m1 >>
rect 523 347 524 348 
<< m1 >>
rect 19 348 20 349 
<< m1 >>
rect 23 348 24 349 
<< m1 >>
rect 44 348 45 349 
<< m1 >>
rect 62 348 63 349 
<< m1 >>
rect 64 348 65 349 
<< m1 >>
rect 67 348 68 349 
<< m1 >>
rect 73 348 74 349 
<< m1 >>
rect 82 348 83 349 
<< m1 >>
rect 91 348 92 349 
<< m1 >>
rect 100 348 101 349 
<< m2 >>
rect 110 348 111 349 
<< m2 >>
rect 111 348 112 349 
<< m2 >>
rect 112 348 113 349 
<< m1 >>
rect 116 348 117 349 
<< m1 >>
rect 118 348 119 349 
<< m2 >>
rect 144 348 145 349 
<< m1 >>
rect 148 348 149 349 
<< m1 >>
rect 150 348 151 349 
<< m1 >>
rect 154 348 155 349 
<< m1 >>
rect 156 348 157 349 
<< m1 >>
rect 157 348 158 349 
<< m1 >>
rect 158 348 159 349 
<< m1 >>
rect 159 348 160 349 
<< m1 >>
rect 160 348 161 349 
<< m1 >>
rect 161 348 162 349 
<< m2 >>
rect 161 348 162 349 
<< m2c >>
rect 161 348 162 349 
<< m1 >>
rect 161 348 162 349 
<< m2 >>
rect 161 348 162 349 
<< m2 >>
rect 162 348 163 349 
<< m1 >>
rect 163 348 164 349 
<< m2 >>
rect 163 348 164 349 
<< m2 >>
rect 164 348 165 349 
<< m1 >>
rect 165 348 166 349 
<< m2 >>
rect 165 348 166 349 
<< m2c >>
rect 165 348 166 349 
<< m1 >>
rect 165 348 166 349 
<< m2 >>
rect 165 348 166 349 
<< m1 >>
rect 166 348 167 349 
<< m1 >>
rect 167 348 168 349 
<< m1 >>
rect 168 348 169 349 
<< m2 >>
rect 168 348 169 349 
<< m1 >>
rect 169 348 170 349 
<< m1 >>
rect 170 348 171 349 
<< m1 >>
rect 171 348 172 349 
<< m1 >>
rect 172 348 173 349 
<< m1 >>
rect 173 348 174 349 
<< m1 >>
rect 174 348 175 349 
<< m2 >>
rect 174 348 175 349 
<< m1 >>
rect 175 348 176 349 
<< m1 >>
rect 176 348 177 349 
<< m1 >>
rect 177 348 178 349 
<< m1 >>
rect 178 348 179 349 
<< m2 >>
rect 182 348 183 349 
<< m2 >>
rect 183 348 184 349 
<< m2 >>
rect 184 348 185 349 
<< m2 >>
rect 185 348 186 349 
<< m2 >>
rect 186 348 187 349 
<< m2 >>
rect 187 348 188 349 
<< m2 >>
rect 188 348 189 349 
<< m2 >>
rect 189 348 190 349 
<< m2 >>
rect 190 348 191 349 
<< m2 >>
rect 191 348 192 349 
<< m2 >>
rect 192 348 193 349 
<< m2 >>
rect 193 348 194 349 
<< m2 >>
rect 194 348 195 349 
<< m2 >>
rect 195 348 196 349 
<< m2 >>
rect 196 348 197 349 
<< m2 >>
rect 197 348 198 349 
<< m2 >>
rect 198 348 199 349 
<< m2 >>
rect 199 348 200 349 
<< m2 >>
rect 200 348 201 349 
<< m2 >>
rect 201 348 202 349 
<< m2 >>
rect 202 348 203 349 
<< m2 >>
rect 203 348 204 349 
<< m2 >>
rect 204 348 205 349 
<< m2 >>
rect 205 348 206 349 
<< m2 >>
rect 206 348 207 349 
<< m2 >>
rect 207 348 208 349 
<< m1 >>
rect 208 348 209 349 
<< m2 >>
rect 208 348 209 349 
<< m2 >>
rect 209 348 210 349 
<< m1 >>
rect 210 348 211 349 
<< m2 >>
rect 210 348 211 349 
<< m2c >>
rect 210 348 211 349 
<< m1 >>
rect 210 348 211 349 
<< m2 >>
rect 210 348 211 349 
<< m1 >>
rect 211 348 212 349 
<< m1 >>
rect 212 348 213 349 
<< m1 >>
rect 217 348 218 349 
<< m2 >>
rect 217 348 218 349 
<< m2c >>
rect 217 348 218 349 
<< m1 >>
rect 217 348 218 349 
<< m2 >>
rect 217 348 218 349 
<< m1 >>
rect 219 348 220 349 
<< m2 >>
rect 219 348 220 349 
<< m2c >>
rect 219 348 220 349 
<< m1 >>
rect 219 348 220 349 
<< m2 >>
rect 219 348 220 349 
<< m1 >>
rect 221 348 222 349 
<< m2 >>
rect 221 348 222 349 
<< m2c >>
rect 221 348 222 349 
<< m1 >>
rect 221 348 222 349 
<< m2 >>
rect 221 348 222 349 
<< m1 >>
rect 223 348 224 349 
<< m2 >>
rect 223 348 224 349 
<< m2c >>
rect 223 348 224 349 
<< m1 >>
rect 223 348 224 349 
<< m2 >>
rect 223 348 224 349 
<< m1 >>
rect 235 348 236 349 
<< m1 >>
rect 242 348 243 349 
<< m1 >>
rect 244 348 245 349 
<< m2 >>
rect 244 348 245 349 
<< m1 >>
rect 253 348 254 349 
<< m1 >>
rect 265 348 266 349 
<< m1 >>
rect 316 348 317 349 
<< m2 >>
rect 321 348 322 349 
<< m2 >>
rect 336 348 337 349 
<< m2 >>
rect 337 348 338 349 
<< m2 >>
rect 338 348 339 349 
<< m2 >>
rect 339 348 340 349 
<< m2 >>
rect 340 348 341 349 
<< m2 >>
rect 341 348 342 349 
<< m2 >>
rect 342 348 343 349 
<< m2 >>
rect 343 348 344 349 
<< m2 >>
rect 344 348 345 349 
<< m2 >>
rect 345 348 346 349 
<< m2 >>
rect 346 348 347 349 
<< m2 >>
rect 347 348 348 349 
<< m2 >>
rect 350 348 351 349 
<< m1 >>
rect 351 348 352 349 
<< m1 >>
rect 379 348 380 349 
<< m2 >>
rect 379 348 380 349 
<< m2c >>
rect 379 348 380 349 
<< m1 >>
rect 379 348 380 349 
<< m2 >>
rect 379 348 380 349 
<< m2 >>
rect 393 348 394 349 
<< m2 >>
rect 394 348 395 349 
<< m2 >>
rect 395 348 396 349 
<< m2 >>
rect 396 348 397 349 
<< m2 >>
rect 397 348 398 349 
<< m2 >>
rect 398 348 399 349 
<< m2 >>
rect 399 348 400 349 
<< m2 >>
rect 400 348 401 349 
<< m2 >>
rect 401 348 402 349 
<< m2 >>
rect 402 348 403 349 
<< m2 >>
rect 403 348 404 349 
<< m2 >>
rect 404 348 405 349 
<< m2 >>
rect 405 348 406 349 
<< m2 >>
rect 406 348 407 349 
<< m2 >>
rect 407 348 408 349 
<< m2 >>
rect 408 348 409 349 
<< m2 >>
rect 409 348 410 349 
<< m2 >>
rect 410 348 411 349 
<< m1 >>
rect 416 348 417 349 
<< m1 >>
rect 418 348 419 349 
<< m2 >>
rect 421 348 422 349 
<< m1 >>
rect 422 348 423 349 
<< m2 >>
rect 422 348 423 349 
<< m2 >>
rect 423 348 424 349 
<< m1 >>
rect 424 348 425 349 
<< m2 >>
rect 424 348 425 349 
<< m2 >>
rect 425 348 426 349 
<< m1 >>
rect 426 348 427 349 
<< m2 >>
rect 426 348 427 349 
<< m2c >>
rect 426 348 427 349 
<< m1 >>
rect 426 348 427 349 
<< m2 >>
rect 426 348 427 349 
<< m1 >>
rect 427 348 428 349 
<< m1 >>
rect 433 348 434 349 
<< m1 >>
rect 435 348 436 349 
<< m1 >>
rect 437 348 438 349 
<< m2 >>
rect 438 348 439 349 
<< m1 >>
rect 439 348 440 349 
<< m2 >>
rect 439 348 440 349 
<< m2c >>
rect 439 348 440 349 
<< m1 >>
rect 439 348 440 349 
<< m2 >>
rect 439 348 440 349 
<< m1 >>
rect 451 348 452 349 
<< m1 >>
rect 523 348 524 349 
<< m1 >>
rect 19 349 20 350 
<< m1 >>
rect 23 349 24 350 
<< m1 >>
rect 42 349 43 350 
<< m2 >>
rect 42 349 43 350 
<< m2c >>
rect 42 349 43 350 
<< m1 >>
rect 42 349 43 350 
<< m2 >>
rect 42 349 43 350 
<< m2 >>
rect 43 349 44 350 
<< m1 >>
rect 44 349 45 350 
<< m2 >>
rect 44 349 45 350 
<< m2 >>
rect 45 349 46 350 
<< m1 >>
rect 46 349 47 350 
<< m2 >>
rect 46 349 47 350 
<< m2c >>
rect 46 349 47 350 
<< m1 >>
rect 46 349 47 350 
<< m2 >>
rect 46 349 47 350 
<< m1 >>
rect 47 349 48 350 
<< m1 >>
rect 48 349 49 350 
<< m1 >>
rect 49 349 50 350 
<< m1 >>
rect 50 349 51 350 
<< m1 >>
rect 51 349 52 350 
<< m1 >>
rect 52 349 53 350 
<< m1 >>
rect 53 349 54 350 
<< m1 >>
rect 54 349 55 350 
<< m1 >>
rect 55 349 56 350 
<< m1 >>
rect 56 349 57 350 
<< m1 >>
rect 57 349 58 350 
<< m1 >>
rect 58 349 59 350 
<< m1 >>
rect 59 349 60 350 
<< m1 >>
rect 60 349 61 350 
<< m2 >>
rect 60 349 61 350 
<< m2c >>
rect 60 349 61 350 
<< m1 >>
rect 60 349 61 350 
<< m2 >>
rect 60 349 61 350 
<< m2 >>
rect 61 349 62 350 
<< m1 >>
rect 62 349 63 350 
<< m2 >>
rect 62 349 63 350 
<< m2 >>
rect 63 349 64 350 
<< m1 >>
rect 64 349 65 350 
<< m2 >>
rect 64 349 65 350 
<< m2 >>
rect 65 349 66 350 
<< m2 >>
rect 66 349 67 350 
<< m1 >>
rect 67 349 68 350 
<< m2 >>
rect 67 349 68 350 
<< m1 >>
rect 68 349 69 350 
<< m2 >>
rect 68 349 69 350 
<< m1 >>
rect 69 349 70 350 
<< m2 >>
rect 69 349 70 350 
<< m1 >>
rect 70 349 71 350 
<< m2 >>
rect 70 349 71 350 
<< m1 >>
rect 71 349 72 350 
<< m2 >>
rect 71 349 72 350 
<< m2 >>
rect 72 349 73 350 
<< m1 >>
rect 73 349 74 350 
<< m2 >>
rect 73 349 74 350 
<< m2 >>
rect 74 349 75 350 
<< m1 >>
rect 75 349 76 350 
<< m2 >>
rect 75 349 76 350 
<< m2c >>
rect 75 349 76 350 
<< m1 >>
rect 75 349 76 350 
<< m2 >>
rect 75 349 76 350 
<< m1 >>
rect 76 349 77 350 
<< m1 >>
rect 77 349 78 350 
<< m1 >>
rect 78 349 79 350 
<< m1 >>
rect 79 349 80 350 
<< m1 >>
rect 80 349 81 350 
<< m2 >>
rect 80 349 81 350 
<< m2c >>
rect 80 349 81 350 
<< m1 >>
rect 80 349 81 350 
<< m2 >>
rect 80 349 81 350 
<< m2 >>
rect 81 349 82 350 
<< m1 >>
rect 82 349 83 350 
<< m2 >>
rect 82 349 83 350 
<< m2 >>
rect 83 349 84 350 
<< m1 >>
rect 84 349 85 350 
<< m2 >>
rect 84 349 85 350 
<< m2c >>
rect 84 349 85 350 
<< m1 >>
rect 84 349 85 350 
<< m2 >>
rect 84 349 85 350 
<< m1 >>
rect 85 349 86 350 
<< m1 >>
rect 86 349 87 350 
<< m1 >>
rect 87 349 88 350 
<< m1 >>
rect 88 349 89 350 
<< m1 >>
rect 89 349 90 350 
<< m2 >>
rect 89 349 90 350 
<< m2c >>
rect 89 349 90 350 
<< m1 >>
rect 89 349 90 350 
<< m2 >>
rect 89 349 90 350 
<< m2 >>
rect 90 349 91 350 
<< m1 >>
rect 91 349 92 350 
<< m2 >>
rect 91 349 92 350 
<< m2 >>
rect 92 349 93 350 
<< m1 >>
rect 93 349 94 350 
<< m2 >>
rect 93 349 94 350 
<< m2c >>
rect 93 349 94 350 
<< m1 >>
rect 93 349 94 350 
<< m2 >>
rect 93 349 94 350 
<< m1 >>
rect 94 349 95 350 
<< m1 >>
rect 95 349 96 350 
<< m1 >>
rect 96 349 97 350 
<< m1 >>
rect 97 349 98 350 
<< m1 >>
rect 98 349 99 350 
<< m2 >>
rect 98 349 99 350 
<< m2c >>
rect 98 349 99 350 
<< m1 >>
rect 98 349 99 350 
<< m2 >>
rect 98 349 99 350 
<< m2 >>
rect 99 349 100 350 
<< m1 >>
rect 100 349 101 350 
<< m2 >>
rect 100 349 101 350 
<< m2 >>
rect 101 349 102 350 
<< m1 >>
rect 102 349 103 350 
<< m2 >>
rect 102 349 103 350 
<< m2c >>
rect 102 349 103 350 
<< m1 >>
rect 102 349 103 350 
<< m2 >>
rect 102 349 103 350 
<< m1 >>
rect 103 349 104 350 
<< m1 >>
rect 104 349 105 350 
<< m1 >>
rect 105 349 106 350 
<< m1 >>
rect 106 349 107 350 
<< m1 >>
rect 107 349 108 350 
<< m1 >>
rect 108 349 109 350 
<< m1 >>
rect 109 349 110 350 
<< m1 >>
rect 110 349 111 350 
<< m2 >>
rect 110 349 111 350 
<< m1 >>
rect 111 349 112 350 
<< m1 >>
rect 112 349 113 350 
<< m1 >>
rect 113 349 114 350 
<< m1 >>
rect 114 349 115 350 
<< m2 >>
rect 114 349 115 350 
<< m2c >>
rect 114 349 115 350 
<< m1 >>
rect 114 349 115 350 
<< m2 >>
rect 114 349 115 350 
<< m2 >>
rect 115 349 116 350 
<< m1 >>
rect 116 349 117 350 
<< m2 >>
rect 116 349 117 350 
<< m2 >>
rect 117 349 118 350 
<< m1 >>
rect 118 349 119 350 
<< m2 >>
rect 118 349 119 350 
<< m2 >>
rect 119 349 120 350 
<< m1 >>
rect 120 349 121 350 
<< m2 >>
rect 120 349 121 350 
<< m2c >>
rect 120 349 121 350 
<< m1 >>
rect 120 349 121 350 
<< m2 >>
rect 120 349 121 350 
<< m1 >>
rect 121 349 122 350 
<< m1 >>
rect 122 349 123 350 
<< m1 >>
rect 123 349 124 350 
<< m1 >>
rect 124 349 125 350 
<< m1 >>
rect 125 349 126 350 
<< m1 >>
rect 127 349 128 350 
<< m1 >>
rect 128 349 129 350 
<< m1 >>
rect 129 349 130 350 
<< m1 >>
rect 130 349 131 350 
<< m1 >>
rect 131 349 132 350 
<< m1 >>
rect 132 349 133 350 
<< m1 >>
rect 133 349 134 350 
<< m1 >>
rect 134 349 135 350 
<< m1 >>
rect 135 349 136 350 
<< m1 >>
rect 136 349 137 350 
<< m1 >>
rect 137 349 138 350 
<< m1 >>
rect 138 349 139 350 
<< m1 >>
rect 139 349 140 350 
<< m1 >>
rect 140 349 141 350 
<< m1 >>
rect 141 349 142 350 
<< m1 >>
rect 142 349 143 350 
<< m1 >>
rect 143 349 144 350 
<< m1 >>
rect 144 349 145 350 
<< m2 >>
rect 144 349 145 350 
<< m1 >>
rect 145 349 146 350 
<< m1 >>
rect 146 349 147 350 
<< m2 >>
rect 146 349 147 350 
<< m2c >>
rect 146 349 147 350 
<< m1 >>
rect 146 349 147 350 
<< m2 >>
rect 146 349 147 350 
<< m2 >>
rect 147 349 148 350 
<< m1 >>
rect 148 349 149 350 
<< m2 >>
rect 148 349 149 350 
<< m2 >>
rect 149 349 150 350 
<< m1 >>
rect 150 349 151 350 
<< m2 >>
rect 150 349 151 350 
<< m2 >>
rect 151 349 152 350 
<< m1 >>
rect 152 349 153 350 
<< m2 >>
rect 152 349 153 350 
<< m2c >>
rect 152 349 153 350 
<< m1 >>
rect 152 349 153 350 
<< m2 >>
rect 152 349 153 350 
<< m2 >>
rect 153 349 154 350 
<< m1 >>
rect 154 349 155 350 
<< m2 >>
rect 154 349 155 350 
<< m2 >>
rect 155 349 156 350 
<< m1 >>
rect 156 349 157 350 
<< m2 >>
rect 156 349 157 350 
<< m2c >>
rect 156 349 157 350 
<< m1 >>
rect 156 349 157 350 
<< m2 >>
rect 156 349 157 350 
<< m1 >>
rect 163 349 164 350 
<< m2 >>
rect 168 349 169 350 
<< m2 >>
rect 174 349 175 350 
<< m1 >>
rect 178 349 179 350 
<< m1 >>
rect 208 349 209 350 
<< m1 >>
rect 212 349 213 350 
<< m1 >>
rect 217 349 218 350 
<< m1 >>
rect 219 349 220 350 
<< m1 >>
rect 221 349 222 350 
<< m1 >>
rect 223 349 224 350 
<< m1 >>
rect 235 349 236 350 
<< m1 >>
rect 242 349 243 350 
<< m1 >>
rect 244 349 245 350 
<< m2 >>
rect 244 349 245 350 
<< m1 >>
rect 253 349 254 350 
<< m1 >>
rect 255 349 256 350 
<< m1 >>
rect 256 349 257 350 
<< m1 >>
rect 257 349 258 350 
<< m1 >>
rect 258 349 259 350 
<< m1 >>
rect 259 349 260 350 
<< m1 >>
rect 260 349 261 350 
<< m1 >>
rect 261 349 262 350 
<< m1 >>
rect 262 349 263 350 
<< m1 >>
rect 263 349 264 350 
<< m1 >>
rect 264 349 265 350 
<< m1 >>
rect 265 349 266 350 
<< m1 >>
rect 316 349 317 350 
<< m2 >>
rect 321 349 322 350 
<< m1 >>
rect 322 349 323 350 
<< m1 >>
rect 323 349 324 350 
<< m1 >>
rect 324 349 325 350 
<< m1 >>
rect 325 349 326 350 
<< m1 >>
rect 326 349 327 350 
<< m1 >>
rect 327 349 328 350 
<< m1 >>
rect 328 349 329 350 
<< m1 >>
rect 329 349 330 350 
<< m1 >>
rect 330 349 331 350 
<< m1 >>
rect 331 349 332 350 
<< m1 >>
rect 332 349 333 350 
<< m1 >>
rect 333 349 334 350 
<< m1 >>
rect 334 349 335 350 
<< m1 >>
rect 335 349 336 350 
<< m1 >>
rect 336 349 337 350 
<< m2 >>
rect 336 349 337 350 
<< m1 >>
rect 337 349 338 350 
<< m1 >>
rect 338 349 339 350 
<< m1 >>
rect 339 349 340 350 
<< m1 >>
rect 340 349 341 350 
<< m1 >>
rect 341 349 342 350 
<< m1 >>
rect 342 349 343 350 
<< m1 >>
rect 343 349 344 350 
<< m1 >>
rect 344 349 345 350 
<< m1 >>
rect 345 349 346 350 
<< m1 >>
rect 346 349 347 350 
<< m1 >>
rect 347 349 348 350 
<< m1 >>
rect 348 349 349 350 
<< m1 >>
rect 349 349 350 350 
<< m1 >>
rect 350 349 351 350 
<< m2 >>
rect 350 349 351 350 
<< m1 >>
rect 351 349 352 350 
<< m1 >>
rect 379 349 380 350 
<< m1 >>
rect 394 349 395 350 
<< m1 >>
rect 395 349 396 350 
<< m1 >>
rect 396 349 397 350 
<< m1 >>
rect 397 349 398 350 
<< m1 >>
rect 398 349 399 350 
<< m1 >>
rect 399 349 400 350 
<< m1 >>
rect 400 349 401 350 
<< m1 >>
rect 401 349 402 350 
<< m1 >>
rect 402 349 403 350 
<< m1 >>
rect 403 349 404 350 
<< m1 >>
rect 404 349 405 350 
<< m1 >>
rect 405 349 406 350 
<< m1 >>
rect 406 349 407 350 
<< m1 >>
rect 407 349 408 350 
<< m1 >>
rect 408 349 409 350 
<< m1 >>
rect 409 349 410 350 
<< m1 >>
rect 410 349 411 350 
<< m2 >>
rect 410 349 411 350 
<< m1 >>
rect 411 349 412 350 
<< m1 >>
rect 412 349 413 350 
<< m1 >>
rect 413 349 414 350 
<< m1 >>
rect 414 349 415 350 
<< m2 >>
rect 414 349 415 350 
<< m2c >>
rect 414 349 415 350 
<< m1 >>
rect 414 349 415 350 
<< m2 >>
rect 414 349 415 350 
<< m2 >>
rect 415 349 416 350 
<< m1 >>
rect 416 349 417 350 
<< m2 >>
rect 416 349 417 350 
<< m2 >>
rect 417 349 418 350 
<< m1 >>
rect 418 349 419 350 
<< m2 >>
rect 418 349 419 350 
<< m2c >>
rect 418 349 419 350 
<< m1 >>
rect 418 349 419 350 
<< m2 >>
rect 418 349 419 350 
<< m1 >>
rect 422 349 423 350 
<< m1 >>
rect 424 349 425 350 
<< m1 >>
rect 427 349 428 350 
<< m1 >>
rect 433 349 434 350 
<< m1 >>
rect 435 349 436 350 
<< m1 >>
rect 437 349 438 350 
<< m2 >>
rect 438 349 439 350 
<< m1 >>
rect 451 349 452 350 
<< m1 >>
rect 523 349 524 350 
<< m1 >>
rect 19 350 20 351 
<< m1 >>
rect 23 350 24 351 
<< m1 >>
rect 42 350 43 351 
<< m1 >>
rect 44 350 45 351 
<< m1 >>
rect 62 350 63 351 
<< m1 >>
rect 64 350 65 351 
<< m1 >>
rect 71 350 72 351 
<< m1 >>
rect 73 350 74 351 
<< m1 >>
rect 82 350 83 351 
<< m1 >>
rect 91 350 92 351 
<< m1 >>
rect 100 350 101 351 
<< m2 >>
rect 110 350 111 351 
<< m1 >>
rect 116 350 117 351 
<< m1 >>
rect 118 350 119 351 
<< m1 >>
rect 125 350 126 351 
<< m1 >>
rect 127 350 128 351 
<< m2 >>
rect 144 350 145 351 
<< m1 >>
rect 148 350 149 351 
<< m1 >>
rect 150 350 151 351 
<< m1 >>
rect 154 350 155 351 
<< m1 >>
rect 163 350 164 351 
<< m2 >>
rect 163 350 164 351 
<< m2c >>
rect 163 350 164 351 
<< m1 >>
rect 163 350 164 351 
<< m2 >>
rect 163 350 164 351 
<< m1 >>
rect 168 350 169 351 
<< m2 >>
rect 168 350 169 351 
<< m2c >>
rect 168 350 169 351 
<< m1 >>
rect 168 350 169 351 
<< m2 >>
rect 168 350 169 351 
<< m1 >>
rect 174 350 175 351 
<< m2 >>
rect 174 350 175 351 
<< m2c >>
rect 174 350 175 351 
<< m1 >>
rect 174 350 175 351 
<< m2 >>
rect 174 350 175 351 
<< m1 >>
rect 178 350 179 351 
<< m1 >>
rect 208 350 209 351 
<< m1 >>
rect 212 350 213 351 
<< m1 >>
rect 213 350 214 351 
<< m1 >>
rect 214 350 215 351 
<< m1 >>
rect 215 350 216 351 
<< m2 >>
rect 215 350 216 351 
<< m2c >>
rect 215 350 216 351 
<< m1 >>
rect 215 350 216 351 
<< m2 >>
rect 215 350 216 351 
<< m2 >>
rect 216 350 217 351 
<< m1 >>
rect 217 350 218 351 
<< m2 >>
rect 217 350 218 351 
<< m2 >>
rect 218 350 219 351 
<< m1 >>
rect 219 350 220 351 
<< m2 >>
rect 219 350 220 351 
<< m2c >>
rect 219 350 220 351 
<< m1 >>
rect 219 350 220 351 
<< m2 >>
rect 219 350 220 351 
<< m1 >>
rect 221 350 222 351 
<< m1 >>
rect 223 350 224 351 
<< m1 >>
rect 235 350 236 351 
<< m2 >>
rect 235 350 236 351 
<< m2c >>
rect 235 350 236 351 
<< m1 >>
rect 235 350 236 351 
<< m2 >>
rect 235 350 236 351 
<< m1 >>
rect 242 350 243 351 
<< m1 >>
rect 244 350 245 351 
<< m2 >>
rect 244 350 245 351 
<< m1 >>
rect 253 350 254 351 
<< m1 >>
rect 255 350 256 351 
<< m1 >>
rect 316 350 317 351 
<< m2 >>
rect 321 350 322 351 
<< m1 >>
rect 322 350 323 351 
<< m2 >>
rect 336 350 337 351 
<< m2 >>
rect 350 350 351 351 
<< m1 >>
rect 379 350 380 351 
<< m1 >>
rect 394 350 395 351 
<< m2 >>
rect 410 350 411 351 
<< m1 >>
rect 416 350 417 351 
<< m1 >>
rect 422 350 423 351 
<< m1 >>
rect 424 350 425 351 
<< m1 >>
rect 427 350 428 351 
<< m1 >>
rect 433 350 434 351 
<< m1 >>
rect 435 350 436 351 
<< m1 >>
rect 437 350 438 351 
<< m2 >>
rect 438 350 439 351 
<< m1 >>
rect 451 350 452 351 
<< m1 >>
rect 523 350 524 351 
<< m1 >>
rect 19 351 20 352 
<< m1 >>
rect 23 351 24 352 
<< m2 >>
rect 38 351 39 352 
<< m1 >>
rect 39 351 40 352 
<< m2 >>
rect 39 351 40 352 
<< m2c >>
rect 39 351 40 352 
<< m1 >>
rect 39 351 40 352 
<< m2 >>
rect 39 351 40 352 
<< m1 >>
rect 40 351 41 352 
<< m1 >>
rect 41 351 42 352 
<< m1 >>
rect 42 351 43 352 
<< m1 >>
rect 44 351 45 352 
<< m1 >>
rect 62 351 63 352 
<< m1 >>
rect 64 351 65 352 
<< m1 >>
rect 71 351 72 352 
<< m1 >>
rect 73 351 74 352 
<< m1 >>
rect 82 351 83 352 
<< m1 >>
rect 91 351 92 352 
<< m1 >>
rect 100 351 101 352 
<< m1 >>
rect 103 351 104 352 
<< m1 >>
rect 104 351 105 352 
<< m1 >>
rect 105 351 106 352 
<< m1 >>
rect 106 351 107 352 
<< m1 >>
rect 107 351 108 352 
<< m1 >>
rect 108 351 109 352 
<< m1 >>
rect 109 351 110 352 
<< m2 >>
rect 110 351 111 352 
<< m1 >>
rect 116 351 117 352 
<< m1 >>
rect 118 351 119 352 
<< m1 >>
rect 125 351 126 352 
<< m1 >>
rect 127 351 128 352 
<< m1 >>
rect 144 351 145 352 
<< m2 >>
rect 144 351 145 352 
<< m2c >>
rect 144 351 145 352 
<< m1 >>
rect 144 351 145 352 
<< m2 >>
rect 144 351 145 352 
<< m1 >>
rect 145 351 146 352 
<< m1 >>
rect 146 351 147 352 
<< m2 >>
rect 146 351 147 352 
<< m2c >>
rect 146 351 147 352 
<< m1 >>
rect 146 351 147 352 
<< m2 >>
rect 146 351 147 352 
<< m2 >>
rect 147 351 148 352 
<< m1 >>
rect 148 351 149 352 
<< m2 >>
rect 148 351 149 352 
<< m2 >>
rect 149 351 150 352 
<< m1 >>
rect 150 351 151 352 
<< m2 >>
rect 150 351 151 352 
<< m2 >>
rect 151 351 152 352 
<< m1 >>
rect 152 351 153 352 
<< m2 >>
rect 152 351 153 352 
<< m2c >>
rect 152 351 153 352 
<< m1 >>
rect 152 351 153 352 
<< m2 >>
rect 152 351 153 352 
<< m1 >>
rect 154 351 155 352 
<< m2 >>
rect 163 351 164 352 
<< m2 >>
rect 168 351 169 352 
<< m2 >>
rect 172 351 173 352 
<< m2 >>
rect 173 351 174 352 
<< m1 >>
rect 174 351 175 352 
<< m2 >>
rect 174 351 175 352 
<< m1 >>
rect 178 351 179 352 
<< m1 >>
rect 208 351 209 352 
<< m1 >>
rect 217 351 218 352 
<< m1 >>
rect 221 351 222 352 
<< m1 >>
rect 223 351 224 352 
<< m2 >>
rect 235 351 236 352 
<< m1 >>
rect 242 351 243 352 
<< m1 >>
rect 244 351 245 352 
<< m2 >>
rect 244 351 245 352 
<< m1 >>
rect 247 351 248 352 
<< m1 >>
rect 248 351 249 352 
<< m1 >>
rect 249 351 250 352 
<< m1 >>
rect 250 351 251 352 
<< m1 >>
rect 251 351 252 352 
<< m2 >>
rect 251 351 252 352 
<< m2c >>
rect 251 351 252 352 
<< m1 >>
rect 251 351 252 352 
<< m2 >>
rect 251 351 252 352 
<< m2 >>
rect 252 351 253 352 
<< m1 >>
rect 253 351 254 352 
<< m2 >>
rect 253 351 254 352 
<< m1 >>
rect 255 351 256 352 
<< m1 >>
rect 316 351 317 352 
<< m2 >>
rect 321 351 322 352 
<< m1 >>
rect 322 351 323 352 
<< m2 >>
rect 322 351 323 352 
<< m2 >>
rect 323 351 324 352 
<< m1 >>
rect 324 351 325 352 
<< m2 >>
rect 324 351 325 352 
<< m2c >>
rect 324 351 325 352 
<< m1 >>
rect 324 351 325 352 
<< m2 >>
rect 324 351 325 352 
<< m1 >>
rect 325 351 326 352 
<< m1 >>
rect 334 351 335 352 
<< m1 >>
rect 335 351 336 352 
<< m1 >>
rect 336 351 337 352 
<< m2 >>
rect 336 351 337 352 
<< m2c >>
rect 336 351 337 352 
<< m1 >>
rect 336 351 337 352 
<< m2 >>
rect 336 351 337 352 
<< m2 >>
rect 350 351 351 352 
<< m1 >>
rect 379 351 380 352 
<< m1 >>
rect 391 351 392 352 
<< m1 >>
rect 392 351 393 352 
<< m2 >>
rect 392 351 393 352 
<< m2c >>
rect 392 351 393 352 
<< m1 >>
rect 392 351 393 352 
<< m2 >>
rect 392 351 393 352 
<< m2 >>
rect 393 351 394 352 
<< m1 >>
rect 394 351 395 352 
<< m2 >>
rect 394 351 395 352 
<< m2 >>
rect 395 351 396 352 
<< m1 >>
rect 410 351 411 352 
<< m2 >>
rect 410 351 411 352 
<< m2c >>
rect 410 351 411 352 
<< m1 >>
rect 410 351 411 352 
<< m2 >>
rect 410 351 411 352 
<< m1 >>
rect 411 351 412 352 
<< m1 >>
rect 412 351 413 352 
<< m1 >>
rect 416 351 417 352 
<< m2 >>
rect 417 351 418 352 
<< m1 >>
rect 418 351 419 352 
<< m2 >>
rect 418 351 419 352 
<< m2c >>
rect 418 351 419 352 
<< m1 >>
rect 418 351 419 352 
<< m2 >>
rect 418 351 419 352 
<< m1 >>
rect 419 351 420 352 
<< m1 >>
rect 420 351 421 352 
<< m1 >>
rect 421 351 422 352 
<< m1 >>
rect 422 351 423 352 
<< m1 >>
rect 424 351 425 352 
<< m1 >>
rect 427 351 428 352 
<< m1 >>
rect 433 351 434 352 
<< m1 >>
rect 435 351 436 352 
<< m1 >>
rect 437 351 438 352 
<< m2 >>
rect 438 351 439 352 
<< m1 >>
rect 451 351 452 352 
<< m1 >>
rect 523 351 524 352 
<< m1 >>
rect 16 352 17 353 
<< m1 >>
rect 17 352 18 353 
<< m2 >>
rect 17 352 18 353 
<< m2c >>
rect 17 352 18 353 
<< m1 >>
rect 17 352 18 353 
<< m2 >>
rect 17 352 18 353 
<< m2 >>
rect 18 352 19 353 
<< m1 >>
rect 19 352 20 353 
<< m2 >>
rect 19 352 20 353 
<< m2 >>
rect 20 352 21 353 
<< m1 >>
rect 21 352 22 353 
<< m2 >>
rect 21 352 22 353 
<< m2c >>
rect 21 352 22 353 
<< m1 >>
rect 21 352 22 353 
<< m2 >>
rect 21 352 22 353 
<< m2 >>
rect 22 352 23 353 
<< m1 >>
rect 23 352 24 353 
<< m2 >>
rect 23 352 24 353 
<< m1 >>
rect 34 352 35 353 
<< m1 >>
rect 35 352 36 353 
<< m1 >>
rect 36 352 37 353 
<< m1 >>
rect 37 352 38 353 
<< m2 >>
rect 38 352 39 353 
<< m1 >>
rect 44 352 45 353 
<< m1 >>
rect 62 352 63 353 
<< m1 >>
rect 64 352 65 353 
<< m1 >>
rect 71 352 72 353 
<< m2 >>
rect 71 352 72 353 
<< m2c >>
rect 71 352 72 353 
<< m1 >>
rect 71 352 72 353 
<< m2 >>
rect 71 352 72 353 
<< m2 >>
rect 72 352 73 353 
<< m1 >>
rect 73 352 74 353 
<< m2 >>
rect 73 352 74 353 
<< m2 >>
rect 74 352 75 353 
<< m1 >>
rect 82 352 83 353 
<< m1 >>
rect 91 352 92 353 
<< m1 >>
rect 100 352 101 353 
<< m1 >>
rect 103 352 104 353 
<< m1 >>
rect 109 352 110 353 
<< m2 >>
rect 110 352 111 353 
<< m1 >>
rect 116 352 117 353 
<< m1 >>
rect 118 352 119 353 
<< m1 >>
rect 125 352 126 353 
<< m2 >>
rect 125 352 126 353 
<< m2c >>
rect 125 352 126 353 
<< m1 >>
rect 125 352 126 353 
<< m2 >>
rect 125 352 126 353 
<< m2 >>
rect 126 352 127 353 
<< m1 >>
rect 127 352 128 353 
<< m2 >>
rect 127 352 128 353 
<< m2 >>
rect 128 352 129 353 
<< m1 >>
rect 148 352 149 353 
<< m1 >>
rect 150 352 151 353 
<< m1 >>
rect 152 352 153 353 
<< m1 >>
rect 154 352 155 353 
<< m1 >>
rect 160 352 161 353 
<< m1 >>
rect 161 352 162 353 
<< m1 >>
rect 162 352 163 353 
<< m1 >>
rect 163 352 164 353 
<< m2 >>
rect 163 352 164 353 
<< m1 >>
rect 164 352 165 353 
<< m1 >>
rect 165 352 166 353 
<< m1 >>
rect 166 352 167 353 
<< m1 >>
rect 167 352 168 353 
<< m1 >>
rect 168 352 169 353 
<< m2 >>
rect 168 352 169 353 
<< m1 >>
rect 169 352 170 353 
<< m1 >>
rect 170 352 171 353 
<< m1 >>
rect 171 352 172 353 
<< m1 >>
rect 172 352 173 353 
<< m2 >>
rect 172 352 173 353 
<< m1 >>
rect 178 352 179 353 
<< m2 >>
rect 207 352 208 353 
<< m1 >>
rect 208 352 209 353 
<< m2 >>
rect 208 352 209 353 
<< m2 >>
rect 209 352 210 353 
<< m1 >>
rect 210 352 211 353 
<< m2 >>
rect 210 352 211 353 
<< m2c >>
rect 210 352 211 353 
<< m1 >>
rect 210 352 211 353 
<< m2 >>
rect 210 352 211 353 
<< m1 >>
rect 211 352 212 353 
<< m1 >>
rect 217 352 218 353 
<< m1 >>
rect 221 352 222 353 
<< m1 >>
rect 223 352 224 353 
<< m1 >>
rect 232 352 233 353 
<< m1 >>
rect 233 352 234 353 
<< m1 >>
rect 234 352 235 353 
<< m1 >>
rect 235 352 236 353 
<< m2 >>
rect 235 352 236 353 
<< m1 >>
rect 242 352 243 353 
<< m1 >>
rect 244 352 245 353 
<< m2 >>
rect 244 352 245 353 
<< m1 >>
rect 247 352 248 353 
<< m1 >>
rect 253 352 254 353 
<< m2 >>
rect 253 352 254 353 
<< m1 >>
rect 255 352 256 353 
<< m1 >>
rect 316 352 317 353 
<< m1 >>
rect 322 352 323 353 
<< m1 >>
rect 325 352 326 353 
<< m1 >>
rect 334 352 335 353 
<< m1 >>
rect 340 352 341 353 
<< m1 >>
rect 341 352 342 353 
<< m1 >>
rect 342 352 343 353 
<< m1 >>
rect 343 352 344 353 
<< m1 >>
rect 344 352 345 353 
<< m1 >>
rect 345 352 346 353 
<< m1 >>
rect 346 352 347 353 
<< m1 >>
rect 347 352 348 353 
<< m1 >>
rect 348 352 349 353 
<< m1 >>
rect 349 352 350 353 
<< m1 >>
rect 350 352 351 353 
<< m2 >>
rect 350 352 351 353 
<< m1 >>
rect 351 352 352 353 
<< m1 >>
rect 352 352 353 353 
<< m1 >>
rect 379 352 380 353 
<< m1 >>
rect 391 352 392 353 
<< m1 >>
rect 394 352 395 353 
<< m2 >>
rect 395 352 396 353 
<< m1 >>
rect 396 352 397 353 
<< m2 >>
rect 396 352 397 353 
<< m2c >>
rect 396 352 397 353 
<< m1 >>
rect 396 352 397 353 
<< m2 >>
rect 396 352 397 353 
<< m1 >>
rect 397 352 398 353 
<< m1 >>
rect 412 352 413 353 
<< m1 >>
rect 416 352 417 353 
<< m2 >>
rect 417 352 418 353 
<< m1 >>
rect 424 352 425 353 
<< m1 >>
rect 427 352 428 353 
<< m1 >>
rect 433 352 434 353 
<< m1 >>
rect 435 352 436 353 
<< m1 >>
rect 437 352 438 353 
<< m2 >>
rect 438 352 439 353 
<< m1 >>
rect 451 352 452 353 
<< m1 >>
rect 523 352 524 353 
<< m1 >>
rect 16 353 17 354 
<< m1 >>
rect 19 353 20 354 
<< m1 >>
rect 23 353 24 354 
<< m2 >>
rect 23 353 24 354 
<< m1 >>
rect 34 353 35 354 
<< m1 >>
rect 37 353 38 354 
<< m2 >>
rect 38 353 39 354 
<< m1 >>
rect 44 353 45 354 
<< m1 >>
rect 62 353 63 354 
<< m1 >>
rect 64 353 65 354 
<< m1 >>
rect 73 353 74 354 
<< m2 >>
rect 74 353 75 354 
<< m1 >>
rect 82 353 83 354 
<< m1 >>
rect 91 353 92 354 
<< m1 >>
rect 100 353 101 354 
<< m1 >>
rect 103 353 104 354 
<< m1 >>
rect 109 353 110 354 
<< m2 >>
rect 110 353 111 354 
<< m1 >>
rect 116 353 117 354 
<< m1 >>
rect 118 353 119 354 
<< m1 >>
rect 127 353 128 354 
<< m2 >>
rect 128 353 129 354 
<< m1 >>
rect 148 353 149 354 
<< m1 >>
rect 150 353 151 354 
<< m1 >>
rect 152 353 153 354 
<< m1 >>
rect 154 353 155 354 
<< m1 >>
rect 160 353 161 354 
<< m2 >>
rect 163 353 164 354 
<< m2 >>
rect 168 353 169 354 
<< m1 >>
rect 172 353 173 354 
<< m2 >>
rect 172 353 173 354 
<< m1 >>
rect 178 353 179 354 
<< m2 >>
rect 207 353 208 354 
<< m1 >>
rect 208 353 209 354 
<< m1 >>
rect 211 353 212 354 
<< m1 >>
rect 217 353 218 354 
<< m1 >>
rect 221 353 222 354 
<< m1 >>
rect 223 353 224 354 
<< m1 >>
rect 232 353 233 354 
<< m1 >>
rect 235 353 236 354 
<< m2 >>
rect 235 353 236 354 
<< m1 >>
rect 242 353 243 354 
<< m1 >>
rect 244 353 245 354 
<< m2 >>
rect 244 353 245 354 
<< m1 >>
rect 247 353 248 354 
<< m1 >>
rect 253 353 254 354 
<< m2 >>
rect 253 353 254 354 
<< m1 >>
rect 255 353 256 354 
<< m1 >>
rect 316 353 317 354 
<< m1 >>
rect 322 353 323 354 
<< m1 >>
rect 325 353 326 354 
<< m1 >>
rect 334 353 335 354 
<< m1 >>
rect 340 353 341 354 
<< m2 >>
rect 343 353 344 354 
<< m2 >>
rect 344 353 345 354 
<< m2 >>
rect 345 353 346 354 
<< m2 >>
rect 346 353 347 354 
<< m2 >>
rect 347 353 348 354 
<< m2 >>
rect 348 353 349 354 
<< m2 >>
rect 349 353 350 354 
<< m2 >>
rect 350 353 351 354 
<< m1 >>
rect 352 353 353 354 
<< m1 >>
rect 379 353 380 354 
<< m1 >>
rect 391 353 392 354 
<< m1 >>
rect 394 353 395 354 
<< m1 >>
rect 397 353 398 354 
<< m1 >>
rect 412 353 413 354 
<< m1 >>
rect 416 353 417 354 
<< m2 >>
rect 417 353 418 354 
<< m1 >>
rect 424 353 425 354 
<< m1 >>
rect 427 353 428 354 
<< m1 >>
rect 433 353 434 354 
<< m1 >>
rect 435 353 436 354 
<< m1 >>
rect 437 353 438 354 
<< m2 >>
rect 438 353 439 354 
<< m1 >>
rect 451 353 452 354 
<< m1 >>
rect 523 353 524 354 
<< pdiffusion >>
rect 12 354 13 355 
<< pdiffusion >>
rect 13 354 14 355 
<< pdiffusion >>
rect 14 354 15 355 
<< pdiffusion >>
rect 15 354 16 355 
<< m1 >>
rect 16 354 17 355 
<< pdiffusion >>
rect 16 354 17 355 
<< pdiffusion >>
rect 17 354 18 355 
<< m1 >>
rect 19 354 20 355 
<< m1 >>
rect 23 354 24 355 
<< m2 >>
rect 23 354 24 355 
<< pdiffusion >>
rect 30 354 31 355 
<< pdiffusion >>
rect 31 354 32 355 
<< pdiffusion >>
rect 32 354 33 355 
<< pdiffusion >>
rect 33 354 34 355 
<< m1 >>
rect 34 354 35 355 
<< pdiffusion >>
rect 34 354 35 355 
<< pdiffusion >>
rect 35 354 36 355 
<< m1 >>
rect 37 354 38 355 
<< m2 >>
rect 38 354 39 355 
<< m1 >>
rect 44 354 45 355 
<< pdiffusion >>
rect 48 354 49 355 
<< pdiffusion >>
rect 49 354 50 355 
<< pdiffusion >>
rect 50 354 51 355 
<< pdiffusion >>
rect 51 354 52 355 
<< pdiffusion >>
rect 52 354 53 355 
<< pdiffusion >>
rect 53 354 54 355 
<< m1 >>
rect 62 354 63 355 
<< m1 >>
rect 64 354 65 355 
<< pdiffusion >>
rect 66 354 67 355 
<< pdiffusion >>
rect 67 354 68 355 
<< pdiffusion >>
rect 68 354 69 355 
<< pdiffusion >>
rect 69 354 70 355 
<< pdiffusion >>
rect 70 354 71 355 
<< pdiffusion >>
rect 71 354 72 355 
<< m1 >>
rect 73 354 74 355 
<< m2 >>
rect 74 354 75 355 
<< m1 >>
rect 82 354 83 355 
<< pdiffusion >>
rect 84 354 85 355 
<< pdiffusion >>
rect 85 354 86 355 
<< pdiffusion >>
rect 86 354 87 355 
<< pdiffusion >>
rect 87 354 88 355 
<< pdiffusion >>
rect 88 354 89 355 
<< pdiffusion >>
rect 89 354 90 355 
<< m1 >>
rect 91 354 92 355 
<< m1 >>
rect 100 354 101 355 
<< pdiffusion >>
rect 102 354 103 355 
<< m1 >>
rect 103 354 104 355 
<< pdiffusion >>
rect 103 354 104 355 
<< pdiffusion >>
rect 104 354 105 355 
<< pdiffusion >>
rect 105 354 106 355 
<< pdiffusion >>
rect 106 354 107 355 
<< pdiffusion >>
rect 107 354 108 355 
<< m1 >>
rect 109 354 110 355 
<< m2 >>
rect 110 354 111 355 
<< m1 >>
rect 116 354 117 355 
<< m1 >>
rect 118 354 119 355 
<< pdiffusion >>
rect 120 354 121 355 
<< pdiffusion >>
rect 121 354 122 355 
<< pdiffusion >>
rect 122 354 123 355 
<< pdiffusion >>
rect 123 354 124 355 
<< pdiffusion >>
rect 124 354 125 355 
<< pdiffusion >>
rect 125 354 126 355 
<< m1 >>
rect 127 354 128 355 
<< m2 >>
rect 128 354 129 355 
<< pdiffusion >>
rect 138 354 139 355 
<< pdiffusion >>
rect 139 354 140 355 
<< pdiffusion >>
rect 140 354 141 355 
<< pdiffusion >>
rect 141 354 142 355 
<< pdiffusion >>
rect 142 354 143 355 
<< pdiffusion >>
rect 143 354 144 355 
<< m1 >>
rect 148 354 149 355 
<< m1 >>
rect 150 354 151 355 
<< m1 >>
rect 152 354 153 355 
<< m1 >>
rect 154 354 155 355 
<< pdiffusion >>
rect 156 354 157 355 
<< pdiffusion >>
rect 157 354 158 355 
<< pdiffusion >>
rect 158 354 159 355 
<< pdiffusion >>
rect 159 354 160 355 
<< m1 >>
rect 160 354 161 355 
<< pdiffusion >>
rect 160 354 161 355 
<< pdiffusion >>
rect 161 354 162 355 
<< m1 >>
rect 163 354 164 355 
<< m2 >>
rect 163 354 164 355 
<< m2c >>
rect 163 354 164 355 
<< m1 >>
rect 163 354 164 355 
<< m2 >>
rect 163 354 164 355 
<< m2 >>
rect 168 354 169 355 
<< m1 >>
rect 169 354 170 355 
<< m1 >>
rect 170 354 171 355 
<< m2 >>
rect 170 354 171 355 
<< m2c >>
rect 170 354 171 355 
<< m1 >>
rect 170 354 171 355 
<< m2 >>
rect 170 354 171 355 
<< m2 >>
rect 171 354 172 355 
<< m1 >>
rect 172 354 173 355 
<< m2 >>
rect 172 354 173 355 
<< pdiffusion >>
rect 174 354 175 355 
<< pdiffusion >>
rect 175 354 176 355 
<< pdiffusion >>
rect 176 354 177 355 
<< pdiffusion >>
rect 177 354 178 355 
<< m1 >>
rect 178 354 179 355 
<< pdiffusion >>
rect 178 354 179 355 
<< pdiffusion >>
rect 179 354 180 355 
<< pdiffusion >>
rect 192 354 193 355 
<< pdiffusion >>
rect 193 354 194 355 
<< pdiffusion >>
rect 194 354 195 355 
<< pdiffusion >>
rect 195 354 196 355 
<< pdiffusion >>
rect 196 354 197 355 
<< pdiffusion >>
rect 197 354 198 355 
<< m2 >>
rect 207 354 208 355 
<< m1 >>
rect 208 354 209 355 
<< pdiffusion >>
rect 210 354 211 355 
<< m1 >>
rect 211 354 212 355 
<< pdiffusion >>
rect 211 354 212 355 
<< pdiffusion >>
rect 212 354 213 355 
<< pdiffusion >>
rect 213 354 214 355 
<< pdiffusion >>
rect 214 354 215 355 
<< pdiffusion >>
rect 215 354 216 355 
<< m1 >>
rect 217 354 218 355 
<< m1 >>
rect 221 354 222 355 
<< m1 >>
rect 223 354 224 355 
<< pdiffusion >>
rect 228 354 229 355 
<< pdiffusion >>
rect 229 354 230 355 
<< pdiffusion >>
rect 230 354 231 355 
<< pdiffusion >>
rect 231 354 232 355 
<< m1 >>
rect 232 354 233 355 
<< pdiffusion >>
rect 232 354 233 355 
<< pdiffusion >>
rect 233 354 234 355 
<< m1 >>
rect 235 354 236 355 
<< m2 >>
rect 235 354 236 355 
<< m1 >>
rect 242 354 243 355 
<< m1 >>
rect 244 354 245 355 
<< m2 >>
rect 244 354 245 355 
<< pdiffusion >>
rect 246 354 247 355 
<< m1 >>
rect 247 354 248 355 
<< pdiffusion >>
rect 247 354 248 355 
<< pdiffusion >>
rect 248 354 249 355 
<< pdiffusion >>
rect 249 354 250 355 
<< pdiffusion >>
rect 250 354 251 355 
<< pdiffusion >>
rect 251 354 252 355 
<< m1 >>
rect 253 354 254 355 
<< m2 >>
rect 253 354 254 355 
<< m1 >>
rect 255 354 256 355 
<< pdiffusion >>
rect 264 354 265 355 
<< pdiffusion >>
rect 265 354 266 355 
<< pdiffusion >>
rect 266 354 267 355 
<< pdiffusion >>
rect 267 354 268 355 
<< pdiffusion >>
rect 268 354 269 355 
<< pdiffusion >>
rect 269 354 270 355 
<< pdiffusion >>
rect 282 354 283 355 
<< pdiffusion >>
rect 283 354 284 355 
<< pdiffusion >>
rect 284 354 285 355 
<< pdiffusion >>
rect 285 354 286 355 
<< pdiffusion >>
rect 286 354 287 355 
<< pdiffusion >>
rect 287 354 288 355 
<< m1 >>
rect 316 354 317 355 
<< pdiffusion >>
rect 318 354 319 355 
<< pdiffusion >>
rect 319 354 320 355 
<< pdiffusion >>
rect 320 354 321 355 
<< pdiffusion >>
rect 321 354 322 355 
<< m1 >>
rect 322 354 323 355 
<< pdiffusion >>
rect 322 354 323 355 
<< pdiffusion >>
rect 323 354 324 355 
<< m1 >>
rect 325 354 326 355 
<< m1 >>
rect 334 354 335 355 
<< pdiffusion >>
rect 336 354 337 355 
<< pdiffusion >>
rect 337 354 338 355 
<< pdiffusion >>
rect 338 354 339 355 
<< pdiffusion >>
rect 339 354 340 355 
<< m1 >>
rect 340 354 341 355 
<< pdiffusion >>
rect 340 354 341 355 
<< pdiffusion >>
rect 341 354 342 355 
<< m1 >>
rect 343 354 344 355 
<< m2 >>
rect 343 354 344 355 
<< m2c >>
rect 343 354 344 355 
<< m1 >>
rect 343 354 344 355 
<< m2 >>
rect 343 354 344 355 
<< m1 >>
rect 352 354 353 355 
<< pdiffusion >>
rect 354 354 355 355 
<< pdiffusion >>
rect 355 354 356 355 
<< pdiffusion >>
rect 356 354 357 355 
<< pdiffusion >>
rect 357 354 358 355 
<< pdiffusion >>
rect 358 354 359 355 
<< pdiffusion >>
rect 359 354 360 355 
<< pdiffusion >>
rect 372 354 373 355 
<< pdiffusion >>
rect 373 354 374 355 
<< pdiffusion >>
rect 374 354 375 355 
<< pdiffusion >>
rect 375 354 376 355 
<< pdiffusion >>
rect 376 354 377 355 
<< pdiffusion >>
rect 377 354 378 355 
<< m1 >>
rect 379 354 380 355 
<< pdiffusion >>
rect 390 354 391 355 
<< m1 >>
rect 391 354 392 355 
<< pdiffusion >>
rect 391 354 392 355 
<< pdiffusion >>
rect 392 354 393 355 
<< pdiffusion >>
rect 393 354 394 355 
<< m1 >>
rect 394 354 395 355 
<< pdiffusion >>
rect 394 354 395 355 
<< pdiffusion >>
rect 395 354 396 355 
<< m1 >>
rect 397 354 398 355 
<< pdiffusion >>
rect 408 354 409 355 
<< pdiffusion >>
rect 409 354 410 355 
<< pdiffusion >>
rect 410 354 411 355 
<< pdiffusion >>
rect 411 354 412 355 
<< m1 >>
rect 412 354 413 355 
<< pdiffusion >>
rect 412 354 413 355 
<< pdiffusion >>
rect 413 354 414 355 
<< m1 >>
rect 416 354 417 355 
<< m2 >>
rect 417 354 418 355 
<< m1 >>
rect 424 354 425 355 
<< pdiffusion >>
rect 426 354 427 355 
<< m1 >>
rect 427 354 428 355 
<< pdiffusion >>
rect 427 354 428 355 
<< pdiffusion >>
rect 428 354 429 355 
<< pdiffusion >>
rect 429 354 430 355 
<< pdiffusion >>
rect 430 354 431 355 
<< pdiffusion >>
rect 431 354 432 355 
<< m1 >>
rect 433 354 434 355 
<< m1 >>
rect 435 354 436 355 
<< m1 >>
rect 437 354 438 355 
<< m2 >>
rect 438 354 439 355 
<< pdiffusion >>
rect 444 354 445 355 
<< pdiffusion >>
rect 445 354 446 355 
<< pdiffusion >>
rect 446 354 447 355 
<< pdiffusion >>
rect 447 354 448 355 
<< pdiffusion >>
rect 448 354 449 355 
<< pdiffusion >>
rect 449 354 450 355 
<< m1 >>
rect 451 354 452 355 
<< pdiffusion >>
rect 462 354 463 355 
<< pdiffusion >>
rect 463 354 464 355 
<< pdiffusion >>
rect 464 354 465 355 
<< pdiffusion >>
rect 465 354 466 355 
<< pdiffusion >>
rect 466 354 467 355 
<< pdiffusion >>
rect 467 354 468 355 
<< pdiffusion >>
rect 480 354 481 355 
<< pdiffusion >>
rect 481 354 482 355 
<< pdiffusion >>
rect 482 354 483 355 
<< pdiffusion >>
rect 483 354 484 355 
<< pdiffusion >>
rect 484 354 485 355 
<< pdiffusion >>
rect 485 354 486 355 
<< pdiffusion >>
rect 498 354 499 355 
<< pdiffusion >>
rect 499 354 500 355 
<< pdiffusion >>
rect 500 354 501 355 
<< pdiffusion >>
rect 501 354 502 355 
<< pdiffusion >>
rect 502 354 503 355 
<< pdiffusion >>
rect 503 354 504 355 
<< pdiffusion >>
rect 516 354 517 355 
<< pdiffusion >>
rect 517 354 518 355 
<< pdiffusion >>
rect 518 354 519 355 
<< pdiffusion >>
rect 519 354 520 355 
<< pdiffusion >>
rect 520 354 521 355 
<< pdiffusion >>
rect 521 354 522 355 
<< m1 >>
rect 523 354 524 355 
<< pdiffusion >>
rect 12 355 13 356 
<< pdiffusion >>
rect 13 355 14 356 
<< pdiffusion >>
rect 14 355 15 356 
<< pdiffusion >>
rect 15 355 16 356 
<< pdiffusion >>
rect 16 355 17 356 
<< pdiffusion >>
rect 17 355 18 356 
<< m1 >>
rect 19 355 20 356 
<< m1 >>
rect 23 355 24 356 
<< m2 >>
rect 23 355 24 356 
<< pdiffusion >>
rect 30 355 31 356 
<< pdiffusion >>
rect 31 355 32 356 
<< pdiffusion >>
rect 32 355 33 356 
<< pdiffusion >>
rect 33 355 34 356 
<< pdiffusion >>
rect 34 355 35 356 
<< pdiffusion >>
rect 35 355 36 356 
<< m1 >>
rect 37 355 38 356 
<< m2 >>
rect 38 355 39 356 
<< m1 >>
rect 44 355 45 356 
<< pdiffusion >>
rect 48 355 49 356 
<< pdiffusion >>
rect 49 355 50 356 
<< pdiffusion >>
rect 50 355 51 356 
<< pdiffusion >>
rect 51 355 52 356 
<< pdiffusion >>
rect 52 355 53 356 
<< pdiffusion >>
rect 53 355 54 356 
<< m1 >>
rect 62 355 63 356 
<< m1 >>
rect 64 355 65 356 
<< pdiffusion >>
rect 66 355 67 356 
<< pdiffusion >>
rect 67 355 68 356 
<< pdiffusion >>
rect 68 355 69 356 
<< pdiffusion >>
rect 69 355 70 356 
<< pdiffusion >>
rect 70 355 71 356 
<< pdiffusion >>
rect 71 355 72 356 
<< m1 >>
rect 73 355 74 356 
<< m2 >>
rect 74 355 75 356 
<< m1 >>
rect 82 355 83 356 
<< pdiffusion >>
rect 84 355 85 356 
<< pdiffusion >>
rect 85 355 86 356 
<< pdiffusion >>
rect 86 355 87 356 
<< pdiffusion >>
rect 87 355 88 356 
<< pdiffusion >>
rect 88 355 89 356 
<< pdiffusion >>
rect 89 355 90 356 
<< m1 >>
rect 91 355 92 356 
<< m1 >>
rect 100 355 101 356 
<< pdiffusion >>
rect 102 355 103 356 
<< pdiffusion >>
rect 103 355 104 356 
<< pdiffusion >>
rect 104 355 105 356 
<< pdiffusion >>
rect 105 355 106 356 
<< pdiffusion >>
rect 106 355 107 356 
<< pdiffusion >>
rect 107 355 108 356 
<< m1 >>
rect 109 355 110 356 
<< m2 >>
rect 110 355 111 356 
<< m1 >>
rect 116 355 117 356 
<< m1 >>
rect 118 355 119 356 
<< pdiffusion >>
rect 120 355 121 356 
<< pdiffusion >>
rect 121 355 122 356 
<< pdiffusion >>
rect 122 355 123 356 
<< pdiffusion >>
rect 123 355 124 356 
<< pdiffusion >>
rect 124 355 125 356 
<< pdiffusion >>
rect 125 355 126 356 
<< m1 >>
rect 127 355 128 356 
<< m2 >>
rect 128 355 129 356 
<< pdiffusion >>
rect 138 355 139 356 
<< pdiffusion >>
rect 139 355 140 356 
<< pdiffusion >>
rect 140 355 141 356 
<< pdiffusion >>
rect 141 355 142 356 
<< pdiffusion >>
rect 142 355 143 356 
<< pdiffusion >>
rect 143 355 144 356 
<< m1 >>
rect 148 355 149 356 
<< m1 >>
rect 150 355 151 356 
<< m1 >>
rect 152 355 153 356 
<< m1 >>
rect 154 355 155 356 
<< pdiffusion >>
rect 156 355 157 356 
<< pdiffusion >>
rect 157 355 158 356 
<< pdiffusion >>
rect 158 355 159 356 
<< pdiffusion >>
rect 159 355 160 356 
<< pdiffusion >>
rect 160 355 161 356 
<< pdiffusion >>
rect 161 355 162 356 
<< m1 >>
rect 163 355 164 356 
<< m2 >>
rect 168 355 169 356 
<< m1 >>
rect 169 355 170 356 
<< m1 >>
rect 172 355 173 356 
<< pdiffusion >>
rect 174 355 175 356 
<< pdiffusion >>
rect 175 355 176 356 
<< pdiffusion >>
rect 176 355 177 356 
<< pdiffusion >>
rect 177 355 178 356 
<< pdiffusion >>
rect 178 355 179 356 
<< pdiffusion >>
rect 179 355 180 356 
<< pdiffusion >>
rect 192 355 193 356 
<< pdiffusion >>
rect 193 355 194 356 
<< pdiffusion >>
rect 194 355 195 356 
<< pdiffusion >>
rect 195 355 196 356 
<< pdiffusion >>
rect 196 355 197 356 
<< pdiffusion >>
rect 197 355 198 356 
<< m2 >>
rect 207 355 208 356 
<< m1 >>
rect 208 355 209 356 
<< pdiffusion >>
rect 210 355 211 356 
<< pdiffusion >>
rect 211 355 212 356 
<< pdiffusion >>
rect 212 355 213 356 
<< pdiffusion >>
rect 213 355 214 356 
<< pdiffusion >>
rect 214 355 215 356 
<< pdiffusion >>
rect 215 355 216 356 
<< m1 >>
rect 217 355 218 356 
<< m1 >>
rect 221 355 222 356 
<< m1 >>
rect 223 355 224 356 
<< pdiffusion >>
rect 228 355 229 356 
<< pdiffusion >>
rect 229 355 230 356 
<< pdiffusion >>
rect 230 355 231 356 
<< pdiffusion >>
rect 231 355 232 356 
<< pdiffusion >>
rect 232 355 233 356 
<< pdiffusion >>
rect 233 355 234 356 
<< m1 >>
rect 235 355 236 356 
<< m2 >>
rect 235 355 236 356 
<< m1 >>
rect 242 355 243 356 
<< m1 >>
rect 244 355 245 356 
<< m2 >>
rect 244 355 245 356 
<< pdiffusion >>
rect 246 355 247 356 
<< pdiffusion >>
rect 247 355 248 356 
<< pdiffusion >>
rect 248 355 249 356 
<< pdiffusion >>
rect 249 355 250 356 
<< pdiffusion >>
rect 250 355 251 356 
<< pdiffusion >>
rect 251 355 252 356 
<< m1 >>
rect 253 355 254 356 
<< m2 >>
rect 253 355 254 356 
<< m1 >>
rect 255 355 256 356 
<< pdiffusion >>
rect 264 355 265 356 
<< pdiffusion >>
rect 265 355 266 356 
<< pdiffusion >>
rect 266 355 267 356 
<< pdiffusion >>
rect 267 355 268 356 
<< pdiffusion >>
rect 268 355 269 356 
<< pdiffusion >>
rect 269 355 270 356 
<< pdiffusion >>
rect 282 355 283 356 
<< pdiffusion >>
rect 283 355 284 356 
<< pdiffusion >>
rect 284 355 285 356 
<< pdiffusion >>
rect 285 355 286 356 
<< pdiffusion >>
rect 286 355 287 356 
<< pdiffusion >>
rect 287 355 288 356 
<< m1 >>
rect 316 355 317 356 
<< pdiffusion >>
rect 318 355 319 356 
<< pdiffusion >>
rect 319 355 320 356 
<< pdiffusion >>
rect 320 355 321 356 
<< pdiffusion >>
rect 321 355 322 356 
<< pdiffusion >>
rect 322 355 323 356 
<< pdiffusion >>
rect 323 355 324 356 
<< m1 >>
rect 325 355 326 356 
<< m1 >>
rect 334 355 335 356 
<< pdiffusion >>
rect 336 355 337 356 
<< pdiffusion >>
rect 337 355 338 356 
<< pdiffusion >>
rect 338 355 339 356 
<< pdiffusion >>
rect 339 355 340 356 
<< pdiffusion >>
rect 340 355 341 356 
<< pdiffusion >>
rect 341 355 342 356 
<< m1 >>
rect 343 355 344 356 
<< m1 >>
rect 352 355 353 356 
<< pdiffusion >>
rect 354 355 355 356 
<< pdiffusion >>
rect 355 355 356 356 
<< pdiffusion >>
rect 356 355 357 356 
<< pdiffusion >>
rect 357 355 358 356 
<< pdiffusion >>
rect 358 355 359 356 
<< pdiffusion >>
rect 359 355 360 356 
<< pdiffusion >>
rect 372 355 373 356 
<< pdiffusion >>
rect 373 355 374 356 
<< pdiffusion >>
rect 374 355 375 356 
<< pdiffusion >>
rect 375 355 376 356 
<< pdiffusion >>
rect 376 355 377 356 
<< pdiffusion >>
rect 377 355 378 356 
<< m1 >>
rect 379 355 380 356 
<< pdiffusion >>
rect 390 355 391 356 
<< pdiffusion >>
rect 391 355 392 356 
<< pdiffusion >>
rect 392 355 393 356 
<< pdiffusion >>
rect 393 355 394 356 
<< pdiffusion >>
rect 394 355 395 356 
<< pdiffusion >>
rect 395 355 396 356 
<< m1 >>
rect 397 355 398 356 
<< pdiffusion >>
rect 408 355 409 356 
<< pdiffusion >>
rect 409 355 410 356 
<< pdiffusion >>
rect 410 355 411 356 
<< pdiffusion >>
rect 411 355 412 356 
<< pdiffusion >>
rect 412 355 413 356 
<< pdiffusion >>
rect 413 355 414 356 
<< m1 >>
rect 416 355 417 356 
<< m2 >>
rect 417 355 418 356 
<< m1 >>
rect 424 355 425 356 
<< pdiffusion >>
rect 426 355 427 356 
<< pdiffusion >>
rect 427 355 428 356 
<< pdiffusion >>
rect 428 355 429 356 
<< pdiffusion >>
rect 429 355 430 356 
<< pdiffusion >>
rect 430 355 431 356 
<< pdiffusion >>
rect 431 355 432 356 
<< m1 >>
rect 433 355 434 356 
<< m1 >>
rect 435 355 436 356 
<< m1 >>
rect 437 355 438 356 
<< m2 >>
rect 438 355 439 356 
<< pdiffusion >>
rect 444 355 445 356 
<< pdiffusion >>
rect 445 355 446 356 
<< pdiffusion >>
rect 446 355 447 356 
<< pdiffusion >>
rect 447 355 448 356 
<< pdiffusion >>
rect 448 355 449 356 
<< pdiffusion >>
rect 449 355 450 356 
<< m1 >>
rect 451 355 452 356 
<< pdiffusion >>
rect 462 355 463 356 
<< pdiffusion >>
rect 463 355 464 356 
<< pdiffusion >>
rect 464 355 465 356 
<< pdiffusion >>
rect 465 355 466 356 
<< pdiffusion >>
rect 466 355 467 356 
<< pdiffusion >>
rect 467 355 468 356 
<< pdiffusion >>
rect 480 355 481 356 
<< pdiffusion >>
rect 481 355 482 356 
<< pdiffusion >>
rect 482 355 483 356 
<< pdiffusion >>
rect 483 355 484 356 
<< pdiffusion >>
rect 484 355 485 356 
<< pdiffusion >>
rect 485 355 486 356 
<< pdiffusion >>
rect 498 355 499 356 
<< pdiffusion >>
rect 499 355 500 356 
<< pdiffusion >>
rect 500 355 501 356 
<< pdiffusion >>
rect 501 355 502 356 
<< pdiffusion >>
rect 502 355 503 356 
<< pdiffusion >>
rect 503 355 504 356 
<< pdiffusion >>
rect 516 355 517 356 
<< pdiffusion >>
rect 517 355 518 356 
<< pdiffusion >>
rect 518 355 519 356 
<< pdiffusion >>
rect 519 355 520 356 
<< pdiffusion >>
rect 520 355 521 356 
<< pdiffusion >>
rect 521 355 522 356 
<< m1 >>
rect 523 355 524 356 
<< pdiffusion >>
rect 12 356 13 357 
<< pdiffusion >>
rect 13 356 14 357 
<< pdiffusion >>
rect 14 356 15 357 
<< pdiffusion >>
rect 15 356 16 357 
<< pdiffusion >>
rect 16 356 17 357 
<< pdiffusion >>
rect 17 356 18 357 
<< m1 >>
rect 19 356 20 357 
<< m1 >>
rect 23 356 24 357 
<< m2 >>
rect 23 356 24 357 
<< pdiffusion >>
rect 30 356 31 357 
<< pdiffusion >>
rect 31 356 32 357 
<< pdiffusion >>
rect 32 356 33 357 
<< pdiffusion >>
rect 33 356 34 357 
<< pdiffusion >>
rect 34 356 35 357 
<< pdiffusion >>
rect 35 356 36 357 
<< m1 >>
rect 37 356 38 357 
<< m2 >>
rect 38 356 39 357 
<< m1 >>
rect 44 356 45 357 
<< pdiffusion >>
rect 48 356 49 357 
<< pdiffusion >>
rect 49 356 50 357 
<< pdiffusion >>
rect 50 356 51 357 
<< pdiffusion >>
rect 51 356 52 357 
<< pdiffusion >>
rect 52 356 53 357 
<< pdiffusion >>
rect 53 356 54 357 
<< m1 >>
rect 62 356 63 357 
<< m1 >>
rect 64 356 65 357 
<< pdiffusion >>
rect 66 356 67 357 
<< pdiffusion >>
rect 67 356 68 357 
<< pdiffusion >>
rect 68 356 69 357 
<< pdiffusion >>
rect 69 356 70 357 
<< pdiffusion >>
rect 70 356 71 357 
<< pdiffusion >>
rect 71 356 72 357 
<< m1 >>
rect 73 356 74 357 
<< m2 >>
rect 74 356 75 357 
<< m1 >>
rect 82 356 83 357 
<< pdiffusion >>
rect 84 356 85 357 
<< pdiffusion >>
rect 85 356 86 357 
<< pdiffusion >>
rect 86 356 87 357 
<< pdiffusion >>
rect 87 356 88 357 
<< pdiffusion >>
rect 88 356 89 357 
<< pdiffusion >>
rect 89 356 90 357 
<< m1 >>
rect 91 356 92 357 
<< m1 >>
rect 100 356 101 357 
<< pdiffusion >>
rect 102 356 103 357 
<< pdiffusion >>
rect 103 356 104 357 
<< pdiffusion >>
rect 104 356 105 357 
<< pdiffusion >>
rect 105 356 106 357 
<< pdiffusion >>
rect 106 356 107 357 
<< pdiffusion >>
rect 107 356 108 357 
<< m1 >>
rect 109 356 110 357 
<< m2 >>
rect 110 356 111 357 
<< m1 >>
rect 116 356 117 357 
<< m1 >>
rect 118 356 119 357 
<< pdiffusion >>
rect 120 356 121 357 
<< pdiffusion >>
rect 121 356 122 357 
<< pdiffusion >>
rect 122 356 123 357 
<< pdiffusion >>
rect 123 356 124 357 
<< pdiffusion >>
rect 124 356 125 357 
<< pdiffusion >>
rect 125 356 126 357 
<< m1 >>
rect 127 356 128 357 
<< m2 >>
rect 128 356 129 357 
<< pdiffusion >>
rect 138 356 139 357 
<< pdiffusion >>
rect 139 356 140 357 
<< pdiffusion >>
rect 140 356 141 357 
<< pdiffusion >>
rect 141 356 142 357 
<< pdiffusion >>
rect 142 356 143 357 
<< pdiffusion >>
rect 143 356 144 357 
<< m1 >>
rect 148 356 149 357 
<< m1 >>
rect 150 356 151 357 
<< m1 >>
rect 152 356 153 357 
<< m1 >>
rect 154 356 155 357 
<< pdiffusion >>
rect 156 356 157 357 
<< pdiffusion >>
rect 157 356 158 357 
<< pdiffusion >>
rect 158 356 159 357 
<< pdiffusion >>
rect 159 356 160 357 
<< pdiffusion >>
rect 160 356 161 357 
<< pdiffusion >>
rect 161 356 162 357 
<< m1 >>
rect 163 356 164 357 
<< m2 >>
rect 168 356 169 357 
<< m1 >>
rect 169 356 170 357 
<< m1 >>
rect 172 356 173 357 
<< pdiffusion >>
rect 174 356 175 357 
<< pdiffusion >>
rect 175 356 176 357 
<< pdiffusion >>
rect 176 356 177 357 
<< pdiffusion >>
rect 177 356 178 357 
<< pdiffusion >>
rect 178 356 179 357 
<< pdiffusion >>
rect 179 356 180 357 
<< pdiffusion >>
rect 192 356 193 357 
<< pdiffusion >>
rect 193 356 194 357 
<< pdiffusion >>
rect 194 356 195 357 
<< pdiffusion >>
rect 195 356 196 357 
<< pdiffusion >>
rect 196 356 197 357 
<< pdiffusion >>
rect 197 356 198 357 
<< m2 >>
rect 207 356 208 357 
<< m1 >>
rect 208 356 209 357 
<< pdiffusion >>
rect 210 356 211 357 
<< pdiffusion >>
rect 211 356 212 357 
<< pdiffusion >>
rect 212 356 213 357 
<< pdiffusion >>
rect 213 356 214 357 
<< pdiffusion >>
rect 214 356 215 357 
<< pdiffusion >>
rect 215 356 216 357 
<< m1 >>
rect 217 356 218 357 
<< m1 >>
rect 221 356 222 357 
<< m1 >>
rect 223 356 224 357 
<< pdiffusion >>
rect 228 356 229 357 
<< pdiffusion >>
rect 229 356 230 357 
<< pdiffusion >>
rect 230 356 231 357 
<< pdiffusion >>
rect 231 356 232 357 
<< pdiffusion >>
rect 232 356 233 357 
<< pdiffusion >>
rect 233 356 234 357 
<< m1 >>
rect 235 356 236 357 
<< m2 >>
rect 235 356 236 357 
<< m1 >>
rect 242 356 243 357 
<< m1 >>
rect 244 356 245 357 
<< m2 >>
rect 244 356 245 357 
<< pdiffusion >>
rect 246 356 247 357 
<< pdiffusion >>
rect 247 356 248 357 
<< pdiffusion >>
rect 248 356 249 357 
<< pdiffusion >>
rect 249 356 250 357 
<< pdiffusion >>
rect 250 356 251 357 
<< pdiffusion >>
rect 251 356 252 357 
<< m1 >>
rect 253 356 254 357 
<< m2 >>
rect 253 356 254 357 
<< m1 >>
rect 255 356 256 357 
<< pdiffusion >>
rect 264 356 265 357 
<< pdiffusion >>
rect 265 356 266 357 
<< pdiffusion >>
rect 266 356 267 357 
<< pdiffusion >>
rect 267 356 268 357 
<< pdiffusion >>
rect 268 356 269 357 
<< pdiffusion >>
rect 269 356 270 357 
<< pdiffusion >>
rect 282 356 283 357 
<< pdiffusion >>
rect 283 356 284 357 
<< pdiffusion >>
rect 284 356 285 357 
<< pdiffusion >>
rect 285 356 286 357 
<< pdiffusion >>
rect 286 356 287 357 
<< pdiffusion >>
rect 287 356 288 357 
<< m1 >>
rect 316 356 317 357 
<< pdiffusion >>
rect 318 356 319 357 
<< pdiffusion >>
rect 319 356 320 357 
<< pdiffusion >>
rect 320 356 321 357 
<< pdiffusion >>
rect 321 356 322 357 
<< pdiffusion >>
rect 322 356 323 357 
<< pdiffusion >>
rect 323 356 324 357 
<< m1 >>
rect 325 356 326 357 
<< m1 >>
rect 334 356 335 357 
<< pdiffusion >>
rect 336 356 337 357 
<< pdiffusion >>
rect 337 356 338 357 
<< pdiffusion >>
rect 338 356 339 357 
<< pdiffusion >>
rect 339 356 340 357 
<< pdiffusion >>
rect 340 356 341 357 
<< pdiffusion >>
rect 341 356 342 357 
<< m1 >>
rect 343 356 344 357 
<< m1 >>
rect 352 356 353 357 
<< pdiffusion >>
rect 354 356 355 357 
<< pdiffusion >>
rect 355 356 356 357 
<< pdiffusion >>
rect 356 356 357 357 
<< pdiffusion >>
rect 357 356 358 357 
<< pdiffusion >>
rect 358 356 359 357 
<< pdiffusion >>
rect 359 356 360 357 
<< pdiffusion >>
rect 372 356 373 357 
<< pdiffusion >>
rect 373 356 374 357 
<< pdiffusion >>
rect 374 356 375 357 
<< pdiffusion >>
rect 375 356 376 357 
<< pdiffusion >>
rect 376 356 377 357 
<< pdiffusion >>
rect 377 356 378 357 
<< m1 >>
rect 379 356 380 357 
<< pdiffusion >>
rect 390 356 391 357 
<< pdiffusion >>
rect 391 356 392 357 
<< pdiffusion >>
rect 392 356 393 357 
<< pdiffusion >>
rect 393 356 394 357 
<< pdiffusion >>
rect 394 356 395 357 
<< pdiffusion >>
rect 395 356 396 357 
<< m1 >>
rect 397 356 398 357 
<< pdiffusion >>
rect 408 356 409 357 
<< pdiffusion >>
rect 409 356 410 357 
<< pdiffusion >>
rect 410 356 411 357 
<< pdiffusion >>
rect 411 356 412 357 
<< pdiffusion >>
rect 412 356 413 357 
<< pdiffusion >>
rect 413 356 414 357 
<< m1 >>
rect 416 356 417 357 
<< m2 >>
rect 417 356 418 357 
<< m1 >>
rect 424 356 425 357 
<< pdiffusion >>
rect 426 356 427 357 
<< pdiffusion >>
rect 427 356 428 357 
<< pdiffusion >>
rect 428 356 429 357 
<< pdiffusion >>
rect 429 356 430 357 
<< pdiffusion >>
rect 430 356 431 357 
<< pdiffusion >>
rect 431 356 432 357 
<< m1 >>
rect 433 356 434 357 
<< m1 >>
rect 435 356 436 357 
<< m1 >>
rect 437 356 438 357 
<< m2 >>
rect 438 356 439 357 
<< pdiffusion >>
rect 444 356 445 357 
<< pdiffusion >>
rect 445 356 446 357 
<< pdiffusion >>
rect 446 356 447 357 
<< pdiffusion >>
rect 447 356 448 357 
<< pdiffusion >>
rect 448 356 449 357 
<< pdiffusion >>
rect 449 356 450 357 
<< m1 >>
rect 451 356 452 357 
<< pdiffusion >>
rect 462 356 463 357 
<< pdiffusion >>
rect 463 356 464 357 
<< pdiffusion >>
rect 464 356 465 357 
<< pdiffusion >>
rect 465 356 466 357 
<< pdiffusion >>
rect 466 356 467 357 
<< pdiffusion >>
rect 467 356 468 357 
<< pdiffusion >>
rect 480 356 481 357 
<< pdiffusion >>
rect 481 356 482 357 
<< pdiffusion >>
rect 482 356 483 357 
<< pdiffusion >>
rect 483 356 484 357 
<< pdiffusion >>
rect 484 356 485 357 
<< pdiffusion >>
rect 485 356 486 357 
<< pdiffusion >>
rect 498 356 499 357 
<< pdiffusion >>
rect 499 356 500 357 
<< pdiffusion >>
rect 500 356 501 357 
<< pdiffusion >>
rect 501 356 502 357 
<< pdiffusion >>
rect 502 356 503 357 
<< pdiffusion >>
rect 503 356 504 357 
<< pdiffusion >>
rect 516 356 517 357 
<< pdiffusion >>
rect 517 356 518 357 
<< pdiffusion >>
rect 518 356 519 357 
<< pdiffusion >>
rect 519 356 520 357 
<< pdiffusion >>
rect 520 356 521 357 
<< pdiffusion >>
rect 521 356 522 357 
<< m1 >>
rect 523 356 524 357 
<< pdiffusion >>
rect 12 357 13 358 
<< pdiffusion >>
rect 13 357 14 358 
<< pdiffusion >>
rect 14 357 15 358 
<< pdiffusion >>
rect 15 357 16 358 
<< pdiffusion >>
rect 16 357 17 358 
<< pdiffusion >>
rect 17 357 18 358 
<< m1 >>
rect 19 357 20 358 
<< m1 >>
rect 23 357 24 358 
<< m2 >>
rect 23 357 24 358 
<< pdiffusion >>
rect 30 357 31 358 
<< pdiffusion >>
rect 31 357 32 358 
<< pdiffusion >>
rect 32 357 33 358 
<< pdiffusion >>
rect 33 357 34 358 
<< pdiffusion >>
rect 34 357 35 358 
<< pdiffusion >>
rect 35 357 36 358 
<< m1 >>
rect 37 357 38 358 
<< m2 >>
rect 38 357 39 358 
<< m1 >>
rect 44 357 45 358 
<< pdiffusion >>
rect 48 357 49 358 
<< pdiffusion >>
rect 49 357 50 358 
<< pdiffusion >>
rect 50 357 51 358 
<< pdiffusion >>
rect 51 357 52 358 
<< pdiffusion >>
rect 52 357 53 358 
<< pdiffusion >>
rect 53 357 54 358 
<< m1 >>
rect 62 357 63 358 
<< m1 >>
rect 64 357 65 358 
<< pdiffusion >>
rect 66 357 67 358 
<< pdiffusion >>
rect 67 357 68 358 
<< pdiffusion >>
rect 68 357 69 358 
<< pdiffusion >>
rect 69 357 70 358 
<< pdiffusion >>
rect 70 357 71 358 
<< pdiffusion >>
rect 71 357 72 358 
<< m1 >>
rect 73 357 74 358 
<< m2 >>
rect 74 357 75 358 
<< m1 >>
rect 82 357 83 358 
<< pdiffusion >>
rect 84 357 85 358 
<< pdiffusion >>
rect 85 357 86 358 
<< pdiffusion >>
rect 86 357 87 358 
<< pdiffusion >>
rect 87 357 88 358 
<< pdiffusion >>
rect 88 357 89 358 
<< pdiffusion >>
rect 89 357 90 358 
<< m1 >>
rect 91 357 92 358 
<< m1 >>
rect 100 357 101 358 
<< pdiffusion >>
rect 102 357 103 358 
<< pdiffusion >>
rect 103 357 104 358 
<< pdiffusion >>
rect 104 357 105 358 
<< pdiffusion >>
rect 105 357 106 358 
<< pdiffusion >>
rect 106 357 107 358 
<< pdiffusion >>
rect 107 357 108 358 
<< m1 >>
rect 109 357 110 358 
<< m2 >>
rect 110 357 111 358 
<< m1 >>
rect 116 357 117 358 
<< m1 >>
rect 118 357 119 358 
<< pdiffusion >>
rect 120 357 121 358 
<< pdiffusion >>
rect 121 357 122 358 
<< pdiffusion >>
rect 122 357 123 358 
<< pdiffusion >>
rect 123 357 124 358 
<< pdiffusion >>
rect 124 357 125 358 
<< pdiffusion >>
rect 125 357 126 358 
<< m1 >>
rect 127 357 128 358 
<< m2 >>
rect 128 357 129 358 
<< pdiffusion >>
rect 138 357 139 358 
<< pdiffusion >>
rect 139 357 140 358 
<< pdiffusion >>
rect 140 357 141 358 
<< pdiffusion >>
rect 141 357 142 358 
<< pdiffusion >>
rect 142 357 143 358 
<< pdiffusion >>
rect 143 357 144 358 
<< m1 >>
rect 148 357 149 358 
<< m1 >>
rect 150 357 151 358 
<< m1 >>
rect 152 357 153 358 
<< m1 >>
rect 154 357 155 358 
<< pdiffusion >>
rect 156 357 157 358 
<< pdiffusion >>
rect 157 357 158 358 
<< pdiffusion >>
rect 158 357 159 358 
<< pdiffusion >>
rect 159 357 160 358 
<< pdiffusion >>
rect 160 357 161 358 
<< pdiffusion >>
rect 161 357 162 358 
<< m1 >>
rect 163 357 164 358 
<< m2 >>
rect 168 357 169 358 
<< m1 >>
rect 169 357 170 358 
<< m1 >>
rect 172 357 173 358 
<< pdiffusion >>
rect 174 357 175 358 
<< pdiffusion >>
rect 175 357 176 358 
<< pdiffusion >>
rect 176 357 177 358 
<< pdiffusion >>
rect 177 357 178 358 
<< pdiffusion >>
rect 178 357 179 358 
<< pdiffusion >>
rect 179 357 180 358 
<< pdiffusion >>
rect 192 357 193 358 
<< pdiffusion >>
rect 193 357 194 358 
<< pdiffusion >>
rect 194 357 195 358 
<< pdiffusion >>
rect 195 357 196 358 
<< pdiffusion >>
rect 196 357 197 358 
<< pdiffusion >>
rect 197 357 198 358 
<< m2 >>
rect 207 357 208 358 
<< m1 >>
rect 208 357 209 358 
<< pdiffusion >>
rect 210 357 211 358 
<< pdiffusion >>
rect 211 357 212 358 
<< pdiffusion >>
rect 212 357 213 358 
<< pdiffusion >>
rect 213 357 214 358 
<< pdiffusion >>
rect 214 357 215 358 
<< pdiffusion >>
rect 215 357 216 358 
<< m1 >>
rect 217 357 218 358 
<< m1 >>
rect 221 357 222 358 
<< m1 >>
rect 223 357 224 358 
<< pdiffusion >>
rect 228 357 229 358 
<< pdiffusion >>
rect 229 357 230 358 
<< pdiffusion >>
rect 230 357 231 358 
<< pdiffusion >>
rect 231 357 232 358 
<< pdiffusion >>
rect 232 357 233 358 
<< pdiffusion >>
rect 233 357 234 358 
<< m1 >>
rect 235 357 236 358 
<< m2 >>
rect 235 357 236 358 
<< m1 >>
rect 242 357 243 358 
<< m1 >>
rect 244 357 245 358 
<< m2 >>
rect 244 357 245 358 
<< pdiffusion >>
rect 246 357 247 358 
<< pdiffusion >>
rect 247 357 248 358 
<< pdiffusion >>
rect 248 357 249 358 
<< pdiffusion >>
rect 249 357 250 358 
<< pdiffusion >>
rect 250 357 251 358 
<< pdiffusion >>
rect 251 357 252 358 
<< m1 >>
rect 253 357 254 358 
<< m2 >>
rect 253 357 254 358 
<< m1 >>
rect 255 357 256 358 
<< pdiffusion >>
rect 264 357 265 358 
<< pdiffusion >>
rect 265 357 266 358 
<< pdiffusion >>
rect 266 357 267 358 
<< pdiffusion >>
rect 267 357 268 358 
<< pdiffusion >>
rect 268 357 269 358 
<< pdiffusion >>
rect 269 357 270 358 
<< pdiffusion >>
rect 282 357 283 358 
<< pdiffusion >>
rect 283 357 284 358 
<< pdiffusion >>
rect 284 357 285 358 
<< pdiffusion >>
rect 285 357 286 358 
<< pdiffusion >>
rect 286 357 287 358 
<< pdiffusion >>
rect 287 357 288 358 
<< m1 >>
rect 316 357 317 358 
<< pdiffusion >>
rect 318 357 319 358 
<< pdiffusion >>
rect 319 357 320 358 
<< pdiffusion >>
rect 320 357 321 358 
<< pdiffusion >>
rect 321 357 322 358 
<< pdiffusion >>
rect 322 357 323 358 
<< pdiffusion >>
rect 323 357 324 358 
<< m1 >>
rect 325 357 326 358 
<< m1 >>
rect 334 357 335 358 
<< pdiffusion >>
rect 336 357 337 358 
<< pdiffusion >>
rect 337 357 338 358 
<< pdiffusion >>
rect 338 357 339 358 
<< pdiffusion >>
rect 339 357 340 358 
<< pdiffusion >>
rect 340 357 341 358 
<< pdiffusion >>
rect 341 357 342 358 
<< m1 >>
rect 343 357 344 358 
<< m1 >>
rect 352 357 353 358 
<< pdiffusion >>
rect 354 357 355 358 
<< pdiffusion >>
rect 355 357 356 358 
<< pdiffusion >>
rect 356 357 357 358 
<< pdiffusion >>
rect 357 357 358 358 
<< pdiffusion >>
rect 358 357 359 358 
<< pdiffusion >>
rect 359 357 360 358 
<< pdiffusion >>
rect 372 357 373 358 
<< pdiffusion >>
rect 373 357 374 358 
<< pdiffusion >>
rect 374 357 375 358 
<< pdiffusion >>
rect 375 357 376 358 
<< pdiffusion >>
rect 376 357 377 358 
<< pdiffusion >>
rect 377 357 378 358 
<< m1 >>
rect 379 357 380 358 
<< pdiffusion >>
rect 390 357 391 358 
<< pdiffusion >>
rect 391 357 392 358 
<< pdiffusion >>
rect 392 357 393 358 
<< pdiffusion >>
rect 393 357 394 358 
<< pdiffusion >>
rect 394 357 395 358 
<< pdiffusion >>
rect 395 357 396 358 
<< m1 >>
rect 397 357 398 358 
<< pdiffusion >>
rect 408 357 409 358 
<< pdiffusion >>
rect 409 357 410 358 
<< pdiffusion >>
rect 410 357 411 358 
<< pdiffusion >>
rect 411 357 412 358 
<< pdiffusion >>
rect 412 357 413 358 
<< pdiffusion >>
rect 413 357 414 358 
<< m1 >>
rect 416 357 417 358 
<< m2 >>
rect 417 357 418 358 
<< m1 >>
rect 424 357 425 358 
<< pdiffusion >>
rect 426 357 427 358 
<< pdiffusion >>
rect 427 357 428 358 
<< pdiffusion >>
rect 428 357 429 358 
<< pdiffusion >>
rect 429 357 430 358 
<< pdiffusion >>
rect 430 357 431 358 
<< pdiffusion >>
rect 431 357 432 358 
<< m1 >>
rect 433 357 434 358 
<< m1 >>
rect 435 357 436 358 
<< m1 >>
rect 437 357 438 358 
<< m2 >>
rect 438 357 439 358 
<< pdiffusion >>
rect 444 357 445 358 
<< pdiffusion >>
rect 445 357 446 358 
<< pdiffusion >>
rect 446 357 447 358 
<< pdiffusion >>
rect 447 357 448 358 
<< pdiffusion >>
rect 448 357 449 358 
<< pdiffusion >>
rect 449 357 450 358 
<< m1 >>
rect 451 357 452 358 
<< pdiffusion >>
rect 462 357 463 358 
<< pdiffusion >>
rect 463 357 464 358 
<< pdiffusion >>
rect 464 357 465 358 
<< pdiffusion >>
rect 465 357 466 358 
<< pdiffusion >>
rect 466 357 467 358 
<< pdiffusion >>
rect 467 357 468 358 
<< pdiffusion >>
rect 480 357 481 358 
<< pdiffusion >>
rect 481 357 482 358 
<< pdiffusion >>
rect 482 357 483 358 
<< pdiffusion >>
rect 483 357 484 358 
<< pdiffusion >>
rect 484 357 485 358 
<< pdiffusion >>
rect 485 357 486 358 
<< pdiffusion >>
rect 498 357 499 358 
<< pdiffusion >>
rect 499 357 500 358 
<< pdiffusion >>
rect 500 357 501 358 
<< pdiffusion >>
rect 501 357 502 358 
<< pdiffusion >>
rect 502 357 503 358 
<< pdiffusion >>
rect 503 357 504 358 
<< pdiffusion >>
rect 516 357 517 358 
<< pdiffusion >>
rect 517 357 518 358 
<< pdiffusion >>
rect 518 357 519 358 
<< pdiffusion >>
rect 519 357 520 358 
<< pdiffusion >>
rect 520 357 521 358 
<< pdiffusion >>
rect 521 357 522 358 
<< m1 >>
rect 523 357 524 358 
<< pdiffusion >>
rect 12 358 13 359 
<< pdiffusion >>
rect 13 358 14 359 
<< pdiffusion >>
rect 14 358 15 359 
<< pdiffusion >>
rect 15 358 16 359 
<< pdiffusion >>
rect 16 358 17 359 
<< pdiffusion >>
rect 17 358 18 359 
<< m1 >>
rect 19 358 20 359 
<< m1 >>
rect 23 358 24 359 
<< m2 >>
rect 23 358 24 359 
<< pdiffusion >>
rect 30 358 31 359 
<< pdiffusion >>
rect 31 358 32 359 
<< pdiffusion >>
rect 32 358 33 359 
<< pdiffusion >>
rect 33 358 34 359 
<< pdiffusion >>
rect 34 358 35 359 
<< pdiffusion >>
rect 35 358 36 359 
<< m1 >>
rect 37 358 38 359 
<< m2 >>
rect 38 358 39 359 
<< m1 >>
rect 44 358 45 359 
<< pdiffusion >>
rect 48 358 49 359 
<< pdiffusion >>
rect 49 358 50 359 
<< pdiffusion >>
rect 50 358 51 359 
<< pdiffusion >>
rect 51 358 52 359 
<< pdiffusion >>
rect 52 358 53 359 
<< pdiffusion >>
rect 53 358 54 359 
<< m1 >>
rect 62 358 63 359 
<< m1 >>
rect 64 358 65 359 
<< pdiffusion >>
rect 66 358 67 359 
<< pdiffusion >>
rect 67 358 68 359 
<< pdiffusion >>
rect 68 358 69 359 
<< pdiffusion >>
rect 69 358 70 359 
<< pdiffusion >>
rect 70 358 71 359 
<< pdiffusion >>
rect 71 358 72 359 
<< m1 >>
rect 73 358 74 359 
<< m2 >>
rect 74 358 75 359 
<< m1 >>
rect 82 358 83 359 
<< pdiffusion >>
rect 84 358 85 359 
<< pdiffusion >>
rect 85 358 86 359 
<< pdiffusion >>
rect 86 358 87 359 
<< pdiffusion >>
rect 87 358 88 359 
<< pdiffusion >>
rect 88 358 89 359 
<< pdiffusion >>
rect 89 358 90 359 
<< m1 >>
rect 91 358 92 359 
<< m1 >>
rect 100 358 101 359 
<< pdiffusion >>
rect 102 358 103 359 
<< pdiffusion >>
rect 103 358 104 359 
<< pdiffusion >>
rect 104 358 105 359 
<< pdiffusion >>
rect 105 358 106 359 
<< pdiffusion >>
rect 106 358 107 359 
<< pdiffusion >>
rect 107 358 108 359 
<< m1 >>
rect 109 358 110 359 
<< m2 >>
rect 110 358 111 359 
<< m1 >>
rect 116 358 117 359 
<< m1 >>
rect 118 358 119 359 
<< pdiffusion >>
rect 120 358 121 359 
<< pdiffusion >>
rect 121 358 122 359 
<< pdiffusion >>
rect 122 358 123 359 
<< pdiffusion >>
rect 123 358 124 359 
<< pdiffusion >>
rect 124 358 125 359 
<< pdiffusion >>
rect 125 358 126 359 
<< m1 >>
rect 127 358 128 359 
<< m2 >>
rect 128 358 129 359 
<< pdiffusion >>
rect 138 358 139 359 
<< pdiffusion >>
rect 139 358 140 359 
<< pdiffusion >>
rect 140 358 141 359 
<< pdiffusion >>
rect 141 358 142 359 
<< pdiffusion >>
rect 142 358 143 359 
<< pdiffusion >>
rect 143 358 144 359 
<< m1 >>
rect 148 358 149 359 
<< m1 >>
rect 150 358 151 359 
<< m1 >>
rect 152 358 153 359 
<< m1 >>
rect 154 358 155 359 
<< pdiffusion >>
rect 156 358 157 359 
<< pdiffusion >>
rect 157 358 158 359 
<< pdiffusion >>
rect 158 358 159 359 
<< pdiffusion >>
rect 159 358 160 359 
<< pdiffusion >>
rect 160 358 161 359 
<< pdiffusion >>
rect 161 358 162 359 
<< m1 >>
rect 163 358 164 359 
<< m2 >>
rect 168 358 169 359 
<< m1 >>
rect 169 358 170 359 
<< m1 >>
rect 172 358 173 359 
<< pdiffusion >>
rect 174 358 175 359 
<< pdiffusion >>
rect 175 358 176 359 
<< pdiffusion >>
rect 176 358 177 359 
<< pdiffusion >>
rect 177 358 178 359 
<< pdiffusion >>
rect 178 358 179 359 
<< pdiffusion >>
rect 179 358 180 359 
<< pdiffusion >>
rect 192 358 193 359 
<< pdiffusion >>
rect 193 358 194 359 
<< pdiffusion >>
rect 194 358 195 359 
<< pdiffusion >>
rect 195 358 196 359 
<< pdiffusion >>
rect 196 358 197 359 
<< pdiffusion >>
rect 197 358 198 359 
<< m2 >>
rect 207 358 208 359 
<< m1 >>
rect 208 358 209 359 
<< pdiffusion >>
rect 210 358 211 359 
<< pdiffusion >>
rect 211 358 212 359 
<< pdiffusion >>
rect 212 358 213 359 
<< pdiffusion >>
rect 213 358 214 359 
<< pdiffusion >>
rect 214 358 215 359 
<< pdiffusion >>
rect 215 358 216 359 
<< m1 >>
rect 217 358 218 359 
<< m1 >>
rect 221 358 222 359 
<< m1 >>
rect 223 358 224 359 
<< pdiffusion >>
rect 228 358 229 359 
<< pdiffusion >>
rect 229 358 230 359 
<< pdiffusion >>
rect 230 358 231 359 
<< pdiffusion >>
rect 231 358 232 359 
<< pdiffusion >>
rect 232 358 233 359 
<< pdiffusion >>
rect 233 358 234 359 
<< m1 >>
rect 235 358 236 359 
<< m2 >>
rect 235 358 236 359 
<< m1 >>
rect 242 358 243 359 
<< m1 >>
rect 244 358 245 359 
<< m2 >>
rect 244 358 245 359 
<< pdiffusion >>
rect 246 358 247 359 
<< pdiffusion >>
rect 247 358 248 359 
<< pdiffusion >>
rect 248 358 249 359 
<< pdiffusion >>
rect 249 358 250 359 
<< pdiffusion >>
rect 250 358 251 359 
<< pdiffusion >>
rect 251 358 252 359 
<< m1 >>
rect 253 358 254 359 
<< m2 >>
rect 253 358 254 359 
<< m1 >>
rect 255 358 256 359 
<< pdiffusion >>
rect 264 358 265 359 
<< pdiffusion >>
rect 265 358 266 359 
<< pdiffusion >>
rect 266 358 267 359 
<< pdiffusion >>
rect 267 358 268 359 
<< pdiffusion >>
rect 268 358 269 359 
<< pdiffusion >>
rect 269 358 270 359 
<< pdiffusion >>
rect 282 358 283 359 
<< pdiffusion >>
rect 283 358 284 359 
<< pdiffusion >>
rect 284 358 285 359 
<< pdiffusion >>
rect 285 358 286 359 
<< pdiffusion >>
rect 286 358 287 359 
<< pdiffusion >>
rect 287 358 288 359 
<< m1 >>
rect 316 358 317 359 
<< pdiffusion >>
rect 318 358 319 359 
<< pdiffusion >>
rect 319 358 320 359 
<< pdiffusion >>
rect 320 358 321 359 
<< pdiffusion >>
rect 321 358 322 359 
<< pdiffusion >>
rect 322 358 323 359 
<< pdiffusion >>
rect 323 358 324 359 
<< m1 >>
rect 325 358 326 359 
<< m1 >>
rect 334 358 335 359 
<< pdiffusion >>
rect 336 358 337 359 
<< pdiffusion >>
rect 337 358 338 359 
<< pdiffusion >>
rect 338 358 339 359 
<< pdiffusion >>
rect 339 358 340 359 
<< pdiffusion >>
rect 340 358 341 359 
<< pdiffusion >>
rect 341 358 342 359 
<< m1 >>
rect 343 358 344 359 
<< m1 >>
rect 352 358 353 359 
<< pdiffusion >>
rect 354 358 355 359 
<< pdiffusion >>
rect 355 358 356 359 
<< pdiffusion >>
rect 356 358 357 359 
<< pdiffusion >>
rect 357 358 358 359 
<< pdiffusion >>
rect 358 358 359 359 
<< pdiffusion >>
rect 359 358 360 359 
<< pdiffusion >>
rect 372 358 373 359 
<< pdiffusion >>
rect 373 358 374 359 
<< pdiffusion >>
rect 374 358 375 359 
<< pdiffusion >>
rect 375 358 376 359 
<< pdiffusion >>
rect 376 358 377 359 
<< pdiffusion >>
rect 377 358 378 359 
<< m1 >>
rect 379 358 380 359 
<< pdiffusion >>
rect 390 358 391 359 
<< pdiffusion >>
rect 391 358 392 359 
<< pdiffusion >>
rect 392 358 393 359 
<< pdiffusion >>
rect 393 358 394 359 
<< pdiffusion >>
rect 394 358 395 359 
<< pdiffusion >>
rect 395 358 396 359 
<< m1 >>
rect 397 358 398 359 
<< pdiffusion >>
rect 408 358 409 359 
<< pdiffusion >>
rect 409 358 410 359 
<< pdiffusion >>
rect 410 358 411 359 
<< pdiffusion >>
rect 411 358 412 359 
<< pdiffusion >>
rect 412 358 413 359 
<< pdiffusion >>
rect 413 358 414 359 
<< m1 >>
rect 416 358 417 359 
<< m2 >>
rect 417 358 418 359 
<< m1 >>
rect 424 358 425 359 
<< pdiffusion >>
rect 426 358 427 359 
<< pdiffusion >>
rect 427 358 428 359 
<< pdiffusion >>
rect 428 358 429 359 
<< pdiffusion >>
rect 429 358 430 359 
<< pdiffusion >>
rect 430 358 431 359 
<< pdiffusion >>
rect 431 358 432 359 
<< m1 >>
rect 433 358 434 359 
<< m1 >>
rect 435 358 436 359 
<< m1 >>
rect 437 358 438 359 
<< m2 >>
rect 438 358 439 359 
<< pdiffusion >>
rect 444 358 445 359 
<< pdiffusion >>
rect 445 358 446 359 
<< pdiffusion >>
rect 446 358 447 359 
<< pdiffusion >>
rect 447 358 448 359 
<< pdiffusion >>
rect 448 358 449 359 
<< pdiffusion >>
rect 449 358 450 359 
<< m1 >>
rect 451 358 452 359 
<< pdiffusion >>
rect 462 358 463 359 
<< pdiffusion >>
rect 463 358 464 359 
<< pdiffusion >>
rect 464 358 465 359 
<< pdiffusion >>
rect 465 358 466 359 
<< pdiffusion >>
rect 466 358 467 359 
<< pdiffusion >>
rect 467 358 468 359 
<< pdiffusion >>
rect 480 358 481 359 
<< pdiffusion >>
rect 481 358 482 359 
<< pdiffusion >>
rect 482 358 483 359 
<< pdiffusion >>
rect 483 358 484 359 
<< pdiffusion >>
rect 484 358 485 359 
<< pdiffusion >>
rect 485 358 486 359 
<< pdiffusion >>
rect 498 358 499 359 
<< pdiffusion >>
rect 499 358 500 359 
<< pdiffusion >>
rect 500 358 501 359 
<< pdiffusion >>
rect 501 358 502 359 
<< pdiffusion >>
rect 502 358 503 359 
<< pdiffusion >>
rect 503 358 504 359 
<< pdiffusion >>
rect 516 358 517 359 
<< pdiffusion >>
rect 517 358 518 359 
<< pdiffusion >>
rect 518 358 519 359 
<< pdiffusion >>
rect 519 358 520 359 
<< pdiffusion >>
rect 520 358 521 359 
<< pdiffusion >>
rect 521 358 522 359 
<< m1 >>
rect 523 358 524 359 
<< pdiffusion >>
rect 12 359 13 360 
<< pdiffusion >>
rect 13 359 14 360 
<< pdiffusion >>
rect 14 359 15 360 
<< pdiffusion >>
rect 15 359 16 360 
<< m1 >>
rect 16 359 17 360 
<< pdiffusion >>
rect 16 359 17 360 
<< pdiffusion >>
rect 17 359 18 360 
<< m1 >>
rect 19 359 20 360 
<< m1 >>
rect 23 359 24 360 
<< m2 >>
rect 23 359 24 360 
<< pdiffusion >>
rect 30 359 31 360 
<< pdiffusion >>
rect 31 359 32 360 
<< pdiffusion >>
rect 32 359 33 360 
<< pdiffusion >>
rect 33 359 34 360 
<< pdiffusion >>
rect 34 359 35 360 
<< pdiffusion >>
rect 35 359 36 360 
<< m1 >>
rect 37 359 38 360 
<< m2 >>
rect 38 359 39 360 
<< m1 >>
rect 44 359 45 360 
<< pdiffusion >>
rect 48 359 49 360 
<< pdiffusion >>
rect 49 359 50 360 
<< pdiffusion >>
rect 50 359 51 360 
<< pdiffusion >>
rect 51 359 52 360 
<< pdiffusion >>
rect 52 359 53 360 
<< pdiffusion >>
rect 53 359 54 360 
<< m1 >>
rect 62 359 63 360 
<< m1 >>
rect 64 359 65 360 
<< pdiffusion >>
rect 66 359 67 360 
<< pdiffusion >>
rect 67 359 68 360 
<< pdiffusion >>
rect 68 359 69 360 
<< pdiffusion >>
rect 69 359 70 360 
<< m1 >>
rect 70 359 71 360 
<< pdiffusion >>
rect 70 359 71 360 
<< pdiffusion >>
rect 71 359 72 360 
<< m1 >>
rect 73 359 74 360 
<< m2 >>
rect 74 359 75 360 
<< m1 >>
rect 82 359 83 360 
<< pdiffusion >>
rect 84 359 85 360 
<< m1 >>
rect 85 359 86 360 
<< pdiffusion >>
rect 85 359 86 360 
<< pdiffusion >>
rect 86 359 87 360 
<< pdiffusion >>
rect 87 359 88 360 
<< m1 >>
rect 88 359 89 360 
<< pdiffusion >>
rect 88 359 89 360 
<< pdiffusion >>
rect 89 359 90 360 
<< m1 >>
rect 91 359 92 360 
<< m1 >>
rect 100 359 101 360 
<< pdiffusion >>
rect 102 359 103 360 
<< m1 >>
rect 103 359 104 360 
<< pdiffusion >>
rect 103 359 104 360 
<< pdiffusion >>
rect 104 359 105 360 
<< pdiffusion >>
rect 105 359 106 360 
<< pdiffusion >>
rect 106 359 107 360 
<< pdiffusion >>
rect 107 359 108 360 
<< m1 >>
rect 109 359 110 360 
<< m2 >>
rect 110 359 111 360 
<< m1 >>
rect 116 359 117 360 
<< m1 >>
rect 118 359 119 360 
<< pdiffusion >>
rect 120 359 121 360 
<< pdiffusion >>
rect 121 359 122 360 
<< pdiffusion >>
rect 122 359 123 360 
<< pdiffusion >>
rect 123 359 124 360 
<< pdiffusion >>
rect 124 359 125 360 
<< pdiffusion >>
rect 125 359 126 360 
<< m1 >>
rect 127 359 128 360 
<< m2 >>
rect 128 359 129 360 
<< pdiffusion >>
rect 138 359 139 360 
<< pdiffusion >>
rect 139 359 140 360 
<< pdiffusion >>
rect 140 359 141 360 
<< pdiffusion >>
rect 141 359 142 360 
<< pdiffusion >>
rect 142 359 143 360 
<< pdiffusion >>
rect 143 359 144 360 
<< m1 >>
rect 148 359 149 360 
<< m1 >>
rect 150 359 151 360 
<< m1 >>
rect 152 359 153 360 
<< m1 >>
rect 154 359 155 360 
<< pdiffusion >>
rect 156 359 157 360 
<< pdiffusion >>
rect 157 359 158 360 
<< pdiffusion >>
rect 158 359 159 360 
<< pdiffusion >>
rect 159 359 160 360 
<< m1 >>
rect 160 359 161 360 
<< pdiffusion >>
rect 160 359 161 360 
<< pdiffusion >>
rect 161 359 162 360 
<< m1 >>
rect 163 359 164 360 
<< m2 >>
rect 168 359 169 360 
<< m1 >>
rect 169 359 170 360 
<< m1 >>
rect 172 359 173 360 
<< pdiffusion >>
rect 174 359 175 360 
<< m1 >>
rect 175 359 176 360 
<< pdiffusion >>
rect 175 359 176 360 
<< pdiffusion >>
rect 176 359 177 360 
<< pdiffusion >>
rect 177 359 178 360 
<< pdiffusion >>
rect 178 359 179 360 
<< pdiffusion >>
rect 179 359 180 360 
<< pdiffusion >>
rect 192 359 193 360 
<< m1 >>
rect 193 359 194 360 
<< pdiffusion >>
rect 193 359 194 360 
<< pdiffusion >>
rect 194 359 195 360 
<< pdiffusion >>
rect 195 359 196 360 
<< m1 >>
rect 196 359 197 360 
<< pdiffusion >>
rect 196 359 197 360 
<< pdiffusion >>
rect 197 359 198 360 
<< m2 >>
rect 207 359 208 360 
<< m1 >>
rect 208 359 209 360 
<< pdiffusion >>
rect 210 359 211 360 
<< pdiffusion >>
rect 211 359 212 360 
<< pdiffusion >>
rect 212 359 213 360 
<< pdiffusion >>
rect 213 359 214 360 
<< pdiffusion >>
rect 214 359 215 360 
<< pdiffusion >>
rect 215 359 216 360 
<< m1 >>
rect 217 359 218 360 
<< m1 >>
rect 221 359 222 360 
<< m1 >>
rect 223 359 224 360 
<< pdiffusion >>
rect 228 359 229 360 
<< pdiffusion >>
rect 229 359 230 360 
<< pdiffusion >>
rect 230 359 231 360 
<< pdiffusion >>
rect 231 359 232 360 
<< m1 >>
rect 232 359 233 360 
<< pdiffusion >>
rect 232 359 233 360 
<< pdiffusion >>
rect 233 359 234 360 
<< m1 >>
rect 235 359 236 360 
<< m2 >>
rect 235 359 236 360 
<< m1 >>
rect 242 359 243 360 
<< m1 >>
rect 244 359 245 360 
<< m2 >>
rect 244 359 245 360 
<< pdiffusion >>
rect 246 359 247 360 
<< m1 >>
rect 247 359 248 360 
<< pdiffusion >>
rect 247 359 248 360 
<< pdiffusion >>
rect 248 359 249 360 
<< pdiffusion >>
rect 249 359 250 360 
<< pdiffusion >>
rect 250 359 251 360 
<< pdiffusion >>
rect 251 359 252 360 
<< m1 >>
rect 253 359 254 360 
<< m2 >>
rect 253 359 254 360 
<< m1 >>
rect 255 359 256 360 
<< pdiffusion >>
rect 264 359 265 360 
<< pdiffusion >>
rect 265 359 266 360 
<< pdiffusion >>
rect 266 359 267 360 
<< pdiffusion >>
rect 267 359 268 360 
<< pdiffusion >>
rect 268 359 269 360 
<< pdiffusion >>
rect 269 359 270 360 
<< pdiffusion >>
rect 282 359 283 360 
<< pdiffusion >>
rect 283 359 284 360 
<< pdiffusion >>
rect 284 359 285 360 
<< pdiffusion >>
rect 285 359 286 360 
<< pdiffusion >>
rect 286 359 287 360 
<< pdiffusion >>
rect 287 359 288 360 
<< m1 >>
rect 316 359 317 360 
<< pdiffusion >>
rect 318 359 319 360 
<< pdiffusion >>
rect 319 359 320 360 
<< pdiffusion >>
rect 320 359 321 360 
<< pdiffusion >>
rect 321 359 322 360 
<< pdiffusion >>
rect 322 359 323 360 
<< pdiffusion >>
rect 323 359 324 360 
<< m1 >>
rect 325 359 326 360 
<< m1 >>
rect 334 359 335 360 
<< pdiffusion >>
rect 336 359 337 360 
<< pdiffusion >>
rect 337 359 338 360 
<< pdiffusion >>
rect 338 359 339 360 
<< pdiffusion >>
rect 339 359 340 360 
<< pdiffusion >>
rect 340 359 341 360 
<< pdiffusion >>
rect 341 359 342 360 
<< m1 >>
rect 343 359 344 360 
<< m1 >>
rect 352 359 353 360 
<< pdiffusion >>
rect 354 359 355 360 
<< pdiffusion >>
rect 355 359 356 360 
<< pdiffusion >>
rect 356 359 357 360 
<< pdiffusion >>
rect 357 359 358 360 
<< pdiffusion >>
rect 358 359 359 360 
<< pdiffusion >>
rect 359 359 360 360 
<< pdiffusion >>
rect 372 359 373 360 
<< pdiffusion >>
rect 373 359 374 360 
<< pdiffusion >>
rect 374 359 375 360 
<< pdiffusion >>
rect 375 359 376 360 
<< pdiffusion >>
rect 376 359 377 360 
<< pdiffusion >>
rect 377 359 378 360 
<< m1 >>
rect 379 359 380 360 
<< pdiffusion >>
rect 390 359 391 360 
<< pdiffusion >>
rect 391 359 392 360 
<< pdiffusion >>
rect 392 359 393 360 
<< pdiffusion >>
rect 393 359 394 360 
<< pdiffusion >>
rect 394 359 395 360 
<< pdiffusion >>
rect 395 359 396 360 
<< m1 >>
rect 397 359 398 360 
<< pdiffusion >>
rect 408 359 409 360 
<< m1 >>
rect 409 359 410 360 
<< pdiffusion >>
rect 409 359 410 360 
<< pdiffusion >>
rect 410 359 411 360 
<< pdiffusion >>
rect 411 359 412 360 
<< pdiffusion >>
rect 412 359 413 360 
<< pdiffusion >>
rect 413 359 414 360 
<< m1 >>
rect 416 359 417 360 
<< m2 >>
rect 417 359 418 360 
<< m1 >>
rect 424 359 425 360 
<< pdiffusion >>
rect 426 359 427 360 
<< pdiffusion >>
rect 427 359 428 360 
<< pdiffusion >>
rect 428 359 429 360 
<< pdiffusion >>
rect 429 359 430 360 
<< pdiffusion >>
rect 430 359 431 360 
<< pdiffusion >>
rect 431 359 432 360 
<< m1 >>
rect 433 359 434 360 
<< m1 >>
rect 435 359 436 360 
<< m1 >>
rect 437 359 438 360 
<< m2 >>
rect 438 359 439 360 
<< pdiffusion >>
rect 444 359 445 360 
<< pdiffusion >>
rect 445 359 446 360 
<< pdiffusion >>
rect 446 359 447 360 
<< pdiffusion >>
rect 447 359 448 360 
<< pdiffusion >>
rect 448 359 449 360 
<< pdiffusion >>
rect 449 359 450 360 
<< m1 >>
rect 451 359 452 360 
<< pdiffusion >>
rect 462 359 463 360 
<< pdiffusion >>
rect 463 359 464 360 
<< pdiffusion >>
rect 464 359 465 360 
<< pdiffusion >>
rect 465 359 466 360 
<< pdiffusion >>
rect 466 359 467 360 
<< pdiffusion >>
rect 467 359 468 360 
<< pdiffusion >>
rect 480 359 481 360 
<< m1 >>
rect 481 359 482 360 
<< pdiffusion >>
rect 481 359 482 360 
<< pdiffusion >>
rect 482 359 483 360 
<< pdiffusion >>
rect 483 359 484 360 
<< pdiffusion >>
rect 484 359 485 360 
<< pdiffusion >>
rect 485 359 486 360 
<< pdiffusion >>
rect 498 359 499 360 
<< pdiffusion >>
rect 499 359 500 360 
<< pdiffusion >>
rect 500 359 501 360 
<< pdiffusion >>
rect 501 359 502 360 
<< pdiffusion >>
rect 502 359 503 360 
<< pdiffusion >>
rect 503 359 504 360 
<< pdiffusion >>
rect 516 359 517 360 
<< pdiffusion >>
rect 517 359 518 360 
<< pdiffusion >>
rect 518 359 519 360 
<< pdiffusion >>
rect 519 359 520 360 
<< pdiffusion >>
rect 520 359 521 360 
<< pdiffusion >>
rect 521 359 522 360 
<< m1 >>
rect 523 359 524 360 
<< m1 >>
rect 16 360 17 361 
<< m1 >>
rect 19 360 20 361 
<< m1 >>
rect 23 360 24 361 
<< m2 >>
rect 23 360 24 361 
<< m1 >>
rect 37 360 38 361 
<< m2 >>
rect 38 360 39 361 
<< m1 >>
rect 44 360 45 361 
<< m1 >>
rect 62 360 63 361 
<< m1 >>
rect 64 360 65 361 
<< m1 >>
rect 70 360 71 361 
<< m1 >>
rect 73 360 74 361 
<< m2 >>
rect 74 360 75 361 
<< m1 >>
rect 82 360 83 361 
<< m1 >>
rect 85 360 86 361 
<< m1 >>
rect 88 360 89 361 
<< m2 >>
rect 88 360 89 361 
<< m2c >>
rect 88 360 89 361 
<< m1 >>
rect 88 360 89 361 
<< m2 >>
rect 88 360 89 361 
<< m1 >>
rect 91 360 92 361 
<< m2 >>
rect 91 360 92 361 
<< m2c >>
rect 91 360 92 361 
<< m1 >>
rect 91 360 92 361 
<< m2 >>
rect 91 360 92 361 
<< m1 >>
rect 100 360 101 361 
<< m1 >>
rect 103 360 104 361 
<< m1 >>
rect 109 360 110 361 
<< m2 >>
rect 110 360 111 361 
<< m1 >>
rect 116 360 117 361 
<< m1 >>
rect 118 360 119 361 
<< m1 >>
rect 127 360 128 361 
<< m2 >>
rect 128 360 129 361 
<< m1 >>
rect 129 360 130 361 
<< m2 >>
rect 129 360 130 361 
<< m2c >>
rect 129 360 130 361 
<< m1 >>
rect 129 360 130 361 
<< m2 >>
rect 129 360 130 361 
<< m1 >>
rect 148 360 149 361 
<< m2 >>
rect 148 360 149 361 
<< m2c >>
rect 148 360 149 361 
<< m1 >>
rect 148 360 149 361 
<< m2 >>
rect 148 360 149 361 
<< m1 >>
rect 150 360 151 361 
<< m2 >>
rect 150 360 151 361 
<< m2c >>
rect 150 360 151 361 
<< m1 >>
rect 150 360 151 361 
<< m2 >>
rect 150 360 151 361 
<< m1 >>
rect 152 360 153 361 
<< m2 >>
rect 152 360 153 361 
<< m2c >>
rect 152 360 153 361 
<< m1 >>
rect 152 360 153 361 
<< m2 >>
rect 152 360 153 361 
<< m1 >>
rect 154 360 155 361 
<< m1 >>
rect 160 360 161 361 
<< m1 >>
rect 163 360 164 361 
<< m2 >>
rect 168 360 169 361 
<< m1 >>
rect 169 360 170 361 
<< m1 >>
rect 172 360 173 361 
<< m1 >>
rect 175 360 176 361 
<< m1 >>
rect 193 360 194 361 
<< m1 >>
rect 196 360 197 361 
<< m2 >>
rect 207 360 208 361 
<< m1 >>
rect 208 360 209 361 
<< m1 >>
rect 217 360 218 361 
<< m1 >>
rect 221 360 222 361 
<< m1 >>
rect 223 360 224 361 
<< m1 >>
rect 232 360 233 361 
<< m1 >>
rect 235 360 236 361 
<< m2 >>
rect 235 360 236 361 
<< m1 >>
rect 242 360 243 361 
<< m1 >>
rect 244 360 245 361 
<< m2 >>
rect 244 360 245 361 
<< m1 >>
rect 247 360 248 361 
<< m1 >>
rect 253 360 254 361 
<< m2 >>
rect 253 360 254 361 
<< m1 >>
rect 255 360 256 361 
<< m1 >>
rect 316 360 317 361 
<< m1 >>
rect 325 360 326 361 
<< m1 >>
rect 334 360 335 361 
<< m1 >>
rect 343 360 344 361 
<< m1 >>
rect 352 360 353 361 
<< m1 >>
rect 379 360 380 361 
<< m1 >>
rect 397 360 398 361 
<< m1 >>
rect 409 360 410 361 
<< m1 >>
rect 416 360 417 361 
<< m2 >>
rect 417 360 418 361 
<< m1 >>
rect 424 360 425 361 
<< m1 >>
rect 433 360 434 361 
<< m1 >>
rect 435 360 436 361 
<< m1 >>
rect 437 360 438 361 
<< m2 >>
rect 438 360 439 361 
<< m1 >>
rect 451 360 452 361 
<< m1 >>
rect 481 360 482 361 
<< m1 >>
rect 523 360 524 361 
<< m1 >>
rect 16 361 17 362 
<< m1 >>
rect 17 361 18 362 
<< m2 >>
rect 17 361 18 362 
<< m2c >>
rect 17 361 18 362 
<< m1 >>
rect 17 361 18 362 
<< m2 >>
rect 17 361 18 362 
<< m2 >>
rect 18 361 19 362 
<< m1 >>
rect 19 361 20 362 
<< m2 >>
rect 19 361 20 362 
<< m2 >>
rect 20 361 21 362 
<< m1 >>
rect 21 361 22 362 
<< m2 >>
rect 21 361 22 362 
<< m2c >>
rect 21 361 22 362 
<< m1 >>
rect 21 361 22 362 
<< m2 >>
rect 21 361 22 362 
<< m1 >>
rect 22 361 23 362 
<< m1 >>
rect 23 361 24 362 
<< m2 >>
rect 23 361 24 362 
<< m1 >>
rect 35 361 36 362 
<< m2 >>
rect 35 361 36 362 
<< m2c >>
rect 35 361 36 362 
<< m1 >>
rect 35 361 36 362 
<< m2 >>
rect 35 361 36 362 
<< m2 >>
rect 36 361 37 362 
<< m1 >>
rect 37 361 38 362 
<< m2 >>
rect 37 361 38 362 
<< m2 >>
rect 38 361 39 362 
<< m1 >>
rect 44 361 45 362 
<< m1 >>
rect 62 361 63 362 
<< m1 >>
rect 64 361 65 362 
<< m1 >>
rect 70 361 71 362 
<< m1 >>
rect 71 361 72 362 
<< m1 >>
rect 72 361 73 362 
<< m1 >>
rect 73 361 74 362 
<< m2 >>
rect 74 361 75 362 
<< m1 >>
rect 82 361 83 362 
<< m1 >>
rect 85 361 86 362 
<< m2 >>
rect 88 361 89 362 
<< m2 >>
rect 91 361 92 362 
<< m2 >>
rect 92 361 93 362 
<< m2 >>
rect 93 361 94 362 
<< m1 >>
rect 100 361 101 362 
<< m1 >>
rect 103 361 104 362 
<< m1 >>
rect 107 361 108 362 
<< m2 >>
rect 107 361 108 362 
<< m2c >>
rect 107 361 108 362 
<< m1 >>
rect 107 361 108 362 
<< m2 >>
rect 107 361 108 362 
<< m2 >>
rect 108 361 109 362 
<< m1 >>
rect 109 361 110 362 
<< m2 >>
rect 109 361 110 362 
<< m2 >>
rect 110 361 111 362 
<< m1 >>
rect 116 361 117 362 
<< m1 >>
rect 118 361 119 362 
<< m1 >>
rect 127 361 128 362 
<< m1 >>
rect 129 361 130 362 
<< m2 >>
rect 148 361 149 362 
<< m2 >>
rect 150 361 151 362 
<< m2 >>
rect 152 361 153 362 
<< m1 >>
rect 154 361 155 362 
<< m1 >>
rect 160 361 161 362 
<< m1 >>
rect 163 361 164 362 
<< m2 >>
rect 168 361 169 362 
<< m1 >>
rect 169 361 170 362 
<< m1 >>
rect 172 361 173 362 
<< m1 >>
rect 175 361 176 362 
<< m1 >>
rect 193 361 194 362 
<< m1 >>
rect 196 361 197 362 
<< m2 >>
rect 197 361 198 362 
<< m1 >>
rect 198 361 199 362 
<< m2 >>
rect 198 361 199 362 
<< m2c >>
rect 198 361 199 362 
<< m1 >>
rect 198 361 199 362 
<< m2 >>
rect 198 361 199 362 
<< m1 >>
rect 199 361 200 362 
<< m1 >>
rect 200 361 201 362 
<< m1 >>
rect 201 361 202 362 
<< m1 >>
rect 202 361 203 362 
<< m1 >>
rect 203 361 204 362 
<< m1 >>
rect 204 361 205 362 
<< m1 >>
rect 205 361 206 362 
<< m1 >>
rect 206 361 207 362 
<< m1 >>
rect 207 361 208 362 
<< m2 >>
rect 207 361 208 362 
<< m1 >>
rect 208 361 209 362 
<< m1 >>
rect 217 361 218 362 
<< m1 >>
rect 221 361 222 362 
<< m1 >>
rect 223 361 224 362 
<< m1 >>
rect 232 361 233 362 
<< m1 >>
rect 235 361 236 362 
<< m2 >>
rect 235 361 236 362 
<< m1 >>
rect 242 361 243 362 
<< m1 >>
rect 244 361 245 362 
<< m2 >>
rect 244 361 245 362 
<< m2 >>
rect 245 361 246 362 
<< m1 >>
rect 246 361 247 362 
<< m2 >>
rect 246 361 247 362 
<< m2c >>
rect 246 361 247 362 
<< m1 >>
rect 246 361 247 362 
<< m2 >>
rect 246 361 247 362 
<< m1 >>
rect 247 361 248 362 
<< m1 >>
rect 251 361 252 362 
<< m2 >>
rect 251 361 252 362 
<< m2c >>
rect 251 361 252 362 
<< m1 >>
rect 251 361 252 362 
<< m2 >>
rect 251 361 252 362 
<< m2 >>
rect 252 361 253 362 
<< m1 >>
rect 253 361 254 362 
<< m2 >>
rect 253 361 254 362 
<< m1 >>
rect 255 361 256 362 
<< m1 >>
rect 316 361 317 362 
<< m1 >>
rect 325 361 326 362 
<< m1 >>
rect 334 361 335 362 
<< m1 >>
rect 343 361 344 362 
<< m1 >>
rect 352 361 353 362 
<< m1 >>
rect 379 361 380 362 
<< m1 >>
rect 397 361 398 362 
<< m1 >>
rect 409 361 410 362 
<< m1 >>
rect 414 361 415 362 
<< m2 >>
rect 414 361 415 362 
<< m2c >>
rect 414 361 415 362 
<< m1 >>
rect 414 361 415 362 
<< m2 >>
rect 414 361 415 362 
<< m2 >>
rect 415 361 416 362 
<< m1 >>
rect 416 361 417 362 
<< m2 >>
rect 416 361 417 362 
<< m2 >>
rect 417 361 418 362 
<< m1 >>
rect 424 361 425 362 
<< m1 >>
rect 431 361 432 362 
<< m2 >>
rect 431 361 432 362 
<< m2c >>
rect 431 361 432 362 
<< m1 >>
rect 431 361 432 362 
<< m2 >>
rect 431 361 432 362 
<< m2 >>
rect 432 361 433 362 
<< m1 >>
rect 433 361 434 362 
<< m2 >>
rect 433 361 434 362 
<< m2 >>
rect 434 361 435 362 
<< m1 >>
rect 435 361 436 362 
<< m2 >>
rect 435 361 436 362 
<< m2 >>
rect 436 361 437 362 
<< m1 >>
rect 437 361 438 362 
<< m2 >>
rect 437 361 438 362 
<< m2 >>
rect 438 361 439 362 
<< m1 >>
rect 451 361 452 362 
<< m1 >>
rect 481 361 482 362 
<< m1 >>
rect 523 361 524 362 
<< m1 >>
rect 19 362 20 363 
<< m2 >>
rect 23 362 24 363 
<< m1 >>
rect 34 362 35 363 
<< m1 >>
rect 35 362 36 363 
<< m1 >>
rect 37 362 38 363 
<< m1 >>
rect 44 362 45 363 
<< m2 >>
rect 44 362 45 363 
<< m2c >>
rect 44 362 45 363 
<< m1 >>
rect 44 362 45 363 
<< m2 >>
rect 44 362 45 363 
<< m1 >>
rect 62 362 63 363 
<< m2 >>
rect 62 362 63 363 
<< m2c >>
rect 62 362 63 363 
<< m1 >>
rect 62 362 63 363 
<< m2 >>
rect 62 362 63 363 
<< m1 >>
rect 64 362 65 363 
<< m2 >>
rect 64 362 65 363 
<< m2c >>
rect 64 362 65 363 
<< m1 >>
rect 64 362 65 363 
<< m2 >>
rect 64 362 65 363 
<< m2 >>
rect 74 362 75 363 
<< m1 >>
rect 82 362 83 363 
<< m1 >>
rect 85 362 86 363 
<< m1 >>
rect 86 362 87 363 
<< m1 >>
rect 87 362 88 363 
<< m1 >>
rect 88 362 89 363 
<< m2 >>
rect 88 362 89 363 
<< m1 >>
rect 89 362 90 363 
<< m1 >>
rect 90 362 91 363 
<< m1 >>
rect 91 362 92 363 
<< m1 >>
rect 92 362 93 363 
<< m1 >>
rect 93 362 94 363 
<< m2 >>
rect 93 362 94 363 
<< m1 >>
rect 94 362 95 363 
<< m1 >>
rect 95 362 96 363 
<< m1 >>
rect 96 362 97 363 
<< m1 >>
rect 97 362 98 363 
<< m1 >>
rect 98 362 99 363 
<< m1 >>
rect 99 362 100 363 
<< m1 >>
rect 100 362 101 363 
<< m1 >>
rect 103 362 104 363 
<< m2 >>
rect 104 362 105 363 
<< m1 >>
rect 105 362 106 363 
<< m2 >>
rect 105 362 106 363 
<< m2c >>
rect 105 362 106 363 
<< m1 >>
rect 105 362 106 363 
<< m2 >>
rect 105 362 106 363 
<< m1 >>
rect 106 362 107 363 
<< m1 >>
rect 107 362 108 363 
<< m1 >>
rect 109 362 110 363 
<< m1 >>
rect 116 362 117 363 
<< m2 >>
rect 116 362 117 363 
<< m2c >>
rect 116 362 117 363 
<< m1 >>
rect 116 362 117 363 
<< m2 >>
rect 116 362 117 363 
<< m1 >>
rect 118 362 119 363 
<< m2 >>
rect 118 362 119 363 
<< m2c >>
rect 118 362 119 363 
<< m1 >>
rect 118 362 119 363 
<< m2 >>
rect 118 362 119 363 
<< m1 >>
rect 127 362 128 363 
<< m2 >>
rect 127 362 128 363 
<< m2c >>
rect 127 362 128 363 
<< m1 >>
rect 127 362 128 363 
<< m2 >>
rect 127 362 128 363 
<< m1 >>
rect 129 362 130 363 
<< m2 >>
rect 129 362 130 363 
<< m2c >>
rect 129 362 130 363 
<< m1 >>
rect 129 362 130 363 
<< m2 >>
rect 129 362 130 363 
<< m1 >>
rect 142 362 143 363 
<< m1 >>
rect 143 362 144 363 
<< m1 >>
rect 144 362 145 363 
<< m1 >>
rect 145 362 146 363 
<< m1 >>
rect 146 362 147 363 
<< m1 >>
rect 147 362 148 363 
<< m1 >>
rect 148 362 149 363 
<< m2 >>
rect 148 362 149 363 
<< m1 >>
rect 149 362 150 363 
<< m1 >>
rect 150 362 151 363 
<< m2 >>
rect 150 362 151 363 
<< m1 >>
rect 151 362 152 363 
<< m1 >>
rect 152 362 153 363 
<< m2 >>
rect 152 362 153 363 
<< m1 >>
rect 153 362 154 363 
<< m1 >>
rect 154 362 155 363 
<< m1 >>
rect 158 362 159 363 
<< m2 >>
rect 158 362 159 363 
<< m2c >>
rect 158 362 159 363 
<< m1 >>
rect 158 362 159 363 
<< m2 >>
rect 158 362 159 363 
<< m1 >>
rect 159 362 160 363 
<< m1 >>
rect 160 362 161 363 
<< m1 >>
rect 163 362 164 363 
<< m2 >>
rect 163 362 164 363 
<< m2c >>
rect 163 362 164 363 
<< m1 >>
rect 163 362 164 363 
<< m2 >>
rect 163 362 164 363 
<< m2 >>
rect 168 362 169 363 
<< m1 >>
rect 169 362 170 363 
<< m1 >>
rect 172 362 173 363 
<< m1 >>
rect 175 362 176 363 
<< m1 >>
rect 193 362 194 363 
<< m1 >>
rect 194 362 195 363 
<< m2 >>
rect 194 362 195 363 
<< m2c >>
rect 194 362 195 363 
<< m1 >>
rect 194 362 195 363 
<< m2 >>
rect 194 362 195 363 
<< m2 >>
rect 195 362 196 363 
<< m1 >>
rect 196 362 197 363 
<< m2 >>
rect 196 362 197 363 
<< m2 >>
rect 197 362 198 363 
<< m2 >>
rect 200 362 201 363 
<< m2 >>
rect 201 362 202 363 
<< m2 >>
rect 202 362 203 363 
<< m2 >>
rect 203 362 204 363 
<< m2 >>
rect 204 362 205 363 
<< m2 >>
rect 205 362 206 363 
<< m2 >>
rect 206 362 207 363 
<< m2 >>
rect 207 362 208 363 
<< m1 >>
rect 212 362 213 363 
<< m2 >>
rect 212 362 213 363 
<< m2c >>
rect 212 362 213 363 
<< m1 >>
rect 212 362 213 363 
<< m2 >>
rect 212 362 213 363 
<< m1 >>
rect 213 362 214 363 
<< m1 >>
rect 214 362 215 363 
<< m1 >>
rect 215 362 216 363 
<< m2 >>
rect 215 362 216 363 
<< m2c >>
rect 215 362 216 363 
<< m1 >>
rect 215 362 216 363 
<< m2 >>
rect 215 362 216 363 
<< m2 >>
rect 216 362 217 363 
<< m1 >>
rect 217 362 218 363 
<< m2 >>
rect 217 362 218 363 
<< m2 >>
rect 218 362 219 363 
<< m1 >>
rect 219 362 220 363 
<< m2 >>
rect 219 362 220 363 
<< m2c >>
rect 219 362 220 363 
<< m1 >>
rect 219 362 220 363 
<< m2 >>
rect 219 362 220 363 
<< m1 >>
rect 220 362 221 363 
<< m1 >>
rect 221 362 222 363 
<< m2 >>
rect 221 362 222 363 
<< m2 >>
rect 222 362 223 363 
<< m1 >>
rect 223 362 224 363 
<< m2 >>
rect 223 362 224 363 
<< m2c >>
rect 223 362 224 363 
<< m1 >>
rect 223 362 224 363 
<< m2 >>
rect 223 362 224 363 
<< m1 >>
rect 232 362 233 363 
<< m1 >>
rect 235 362 236 363 
<< m2 >>
rect 235 362 236 363 
<< m1 >>
rect 242 362 243 363 
<< m1 >>
rect 244 362 245 363 
<< m1 >>
rect 251 362 252 363 
<< m1 >>
rect 253 362 254 363 
<< m1 >>
rect 255 362 256 363 
<< m1 >>
rect 316 362 317 363 
<< m1 >>
rect 325 362 326 363 
<< m1 >>
rect 334 362 335 363 
<< m2 >>
rect 334 362 335 363 
<< m2c >>
rect 334 362 335 363 
<< m1 >>
rect 334 362 335 363 
<< m2 >>
rect 334 362 335 363 
<< m1 >>
rect 343 362 344 363 
<< m1 >>
rect 352 362 353 363 
<< m1 >>
rect 379 362 380 363 
<< m2 >>
rect 379 362 380 363 
<< m2c >>
rect 379 362 380 363 
<< m1 >>
rect 379 362 380 363 
<< m2 >>
rect 379 362 380 363 
<< m1 >>
rect 397 362 398 363 
<< m2 >>
rect 397 362 398 363 
<< m2c >>
rect 397 362 398 363 
<< m1 >>
rect 397 362 398 363 
<< m2 >>
rect 397 362 398 363 
<< m1 >>
rect 409 362 410 363 
<< m2 >>
rect 409 362 410 363 
<< m2c >>
rect 409 362 410 363 
<< m1 >>
rect 409 362 410 363 
<< m2 >>
rect 409 362 410 363 
<< m1 >>
rect 414 362 415 363 
<< m1 >>
rect 416 362 417 363 
<< m1 >>
rect 424 362 425 363 
<< m1 >>
rect 429 362 430 363 
<< m2 >>
rect 429 362 430 363 
<< m2c >>
rect 429 362 430 363 
<< m1 >>
rect 429 362 430 363 
<< m2 >>
rect 429 362 430 363 
<< m1 >>
rect 430 362 431 363 
<< m1 >>
rect 431 362 432 363 
<< m1 >>
rect 433 362 434 363 
<< m1 >>
rect 435 362 436 363 
<< m1 >>
rect 437 362 438 363 
<< m1 >>
rect 446 362 447 363 
<< m2 >>
rect 446 362 447 363 
<< m2c >>
rect 446 362 447 363 
<< m1 >>
rect 446 362 447 363 
<< m2 >>
rect 446 362 447 363 
<< m1 >>
rect 447 362 448 363 
<< m1 >>
rect 448 362 449 363 
<< m1 >>
rect 449 362 450 363 
<< m2 >>
rect 449 362 450 363 
<< m2c >>
rect 449 362 450 363 
<< m1 >>
rect 449 362 450 363 
<< m2 >>
rect 449 362 450 363 
<< m2 >>
rect 450 362 451 363 
<< m1 >>
rect 451 362 452 363 
<< m2 >>
rect 451 362 452 363 
<< m2 >>
rect 452 362 453 363 
<< m1 >>
rect 481 362 482 363 
<< m1 >>
rect 523 362 524 363 
<< m1 >>
rect 19 363 20 364 
<< m1 >>
rect 23 363 24 364 
<< m2 >>
rect 23 363 24 364 
<< m2c >>
rect 23 363 24 364 
<< m1 >>
rect 23 363 24 364 
<< m2 >>
rect 23 363 24 364 
<< m1 >>
rect 34 363 35 364 
<< m1 >>
rect 37 363 38 364 
<< m2 >>
rect 44 363 45 364 
<< m2 >>
rect 62 363 63 364 
<< m2 >>
rect 64 363 65 364 
<< m2 >>
rect 74 363 75 364 
<< m1 >>
rect 82 363 83 364 
<< m2 >>
rect 88 363 89 364 
<< m2 >>
rect 93 363 94 364 
<< m1 >>
rect 103 363 104 364 
<< m2 >>
rect 104 363 105 364 
<< m1 >>
rect 109 363 110 364 
<< m2 >>
rect 116 363 117 364 
<< m2 >>
rect 118 363 119 364 
<< m2 >>
rect 127 363 128 364 
<< m2 >>
rect 129 363 130 364 
<< m1 >>
rect 142 363 143 364 
<< m2 >>
rect 148 363 149 364 
<< m2 >>
rect 150 363 151 364 
<< m2 >>
rect 152 363 153 364 
<< m2 >>
rect 158 363 159 364 
<< m2 >>
rect 163 363 164 364 
<< m2 >>
rect 168 363 169 364 
<< m1 >>
rect 169 363 170 364 
<< m1 >>
rect 172 363 173 364 
<< m1 >>
rect 175 363 176 364 
<< m1 >>
rect 196 363 197 364 
<< m1 >>
rect 200 363 201 364 
<< m2 >>
rect 200 363 201 364 
<< m2c >>
rect 200 363 201 364 
<< m1 >>
rect 200 363 201 364 
<< m2 >>
rect 200 363 201 364 
<< m2 >>
rect 212 363 213 364 
<< m1 >>
rect 217 363 218 364 
<< m2 >>
rect 221 363 222 364 
<< m1 >>
rect 232 363 233 364 
<< m1 >>
rect 235 363 236 364 
<< m2 >>
rect 235 363 236 364 
<< m1 >>
rect 242 363 243 364 
<< m1 >>
rect 244 363 245 364 
<< m1 >>
rect 251 363 252 364 
<< m1 >>
rect 253 363 254 364 
<< m1 >>
rect 255 363 256 364 
<< m1 >>
rect 316 363 317 364 
<< m1 >>
rect 325 363 326 364 
<< m2 >>
rect 334 363 335 364 
<< m1 >>
rect 343 363 344 364 
<< m1 >>
rect 352 363 353 364 
<< m2 >>
rect 379 363 380 364 
<< m2 >>
rect 397 363 398 364 
<< m2 >>
rect 409 363 410 364 
<< m2 >>
rect 410 363 411 364 
<< m2 >>
rect 411 363 412 364 
<< m2 >>
rect 412 363 413 364 
<< m2 >>
rect 413 363 414 364 
<< m1 >>
rect 414 363 415 364 
<< m2 >>
rect 414 363 415 364 
<< m2 >>
rect 415 363 416 364 
<< m1 >>
rect 416 363 417 364 
<< m2 >>
rect 416 363 417 364 
<< m2 >>
rect 417 363 418 364 
<< m1 >>
rect 418 363 419 364 
<< m2 >>
rect 418 363 419 364 
<< m2c >>
rect 418 363 419 364 
<< m1 >>
rect 418 363 419 364 
<< m2 >>
rect 418 363 419 364 
<< m1 >>
rect 419 363 420 364 
<< m1 >>
rect 420 363 421 364 
<< m1 >>
rect 421 363 422 364 
<< m1 >>
rect 422 363 423 364 
<< m2 >>
rect 422 363 423 364 
<< m2c >>
rect 422 363 423 364 
<< m1 >>
rect 422 363 423 364 
<< m2 >>
rect 422 363 423 364 
<< m2 >>
rect 423 363 424 364 
<< m1 >>
rect 424 363 425 364 
<< m2 >>
rect 424 363 425 364 
<< m2 >>
rect 425 363 426 364 
<< m1 >>
rect 426 363 427 364 
<< m2 >>
rect 426 363 427 364 
<< m2c >>
rect 426 363 427 364 
<< m1 >>
rect 426 363 427 364 
<< m2 >>
rect 426 363 427 364 
<< m2 >>
rect 429 363 430 364 
<< m1 >>
rect 433 363 434 364 
<< m1 >>
rect 435 363 436 364 
<< m1 >>
rect 437 363 438 364 
<< m2 >>
rect 446 363 447 364 
<< m1 >>
rect 451 363 452 364 
<< m2 >>
rect 452 363 453 364 
<< m1 >>
rect 481 363 482 364 
<< m1 >>
rect 523 363 524 364 
<< m1 >>
rect 19 364 20 365 
<< m1 >>
rect 23 364 24 365 
<< m1 >>
rect 34 364 35 365 
<< m1 >>
rect 37 364 38 365 
<< m1 >>
rect 38 364 39 365 
<< m1 >>
rect 39 364 40 365 
<< m1 >>
rect 40 364 41 365 
<< m1 >>
rect 41 364 42 365 
<< m1 >>
rect 42 364 43 365 
<< m1 >>
rect 43 364 44 365 
<< m1 >>
rect 44 364 45 365 
<< m2 >>
rect 44 364 45 365 
<< m1 >>
rect 45 364 46 365 
<< m1 >>
rect 46 364 47 365 
<< m1 >>
rect 47 364 48 365 
<< m1 >>
rect 48 364 49 365 
<< m1 >>
rect 49 364 50 365 
<< m1 >>
rect 50 364 51 365 
<< m1 >>
rect 51 364 52 365 
<< m1 >>
rect 52 364 53 365 
<< m1 >>
rect 53 364 54 365 
<< m1 >>
rect 54 364 55 365 
<< m1 >>
rect 55 364 56 365 
<< m1 >>
rect 56 364 57 365 
<< m1 >>
rect 57 364 58 365 
<< m1 >>
rect 58 364 59 365 
<< m1 >>
rect 59 364 60 365 
<< m1 >>
rect 60 364 61 365 
<< m1 >>
rect 61 364 62 365 
<< m1 >>
rect 62 364 63 365 
<< m2 >>
rect 62 364 63 365 
<< m1 >>
rect 63 364 64 365 
<< m1 >>
rect 64 364 65 365 
<< m2 >>
rect 64 364 65 365 
<< m1 >>
rect 65 364 66 365 
<< m1 >>
rect 66 364 67 365 
<< m1 >>
rect 67 364 68 365 
<< m1 >>
rect 68 364 69 365 
<< m1 >>
rect 69 364 70 365 
<< m1 >>
rect 70 364 71 365 
<< m1 >>
rect 71 364 72 365 
<< m1 >>
rect 72 364 73 365 
<< m1 >>
rect 73 364 74 365 
<< m1 >>
rect 74 364 75 365 
<< m2 >>
rect 74 364 75 365 
<< m1 >>
rect 75 364 76 365 
<< m1 >>
rect 76 364 77 365 
<< m1 >>
rect 77 364 78 365 
<< m1 >>
rect 78 364 79 365 
<< m1 >>
rect 79 364 80 365 
<< m1 >>
rect 80 364 81 365 
<< m2 >>
rect 80 364 81 365 
<< m2c >>
rect 80 364 81 365 
<< m1 >>
rect 80 364 81 365 
<< m2 >>
rect 80 364 81 365 
<< m2 >>
rect 81 364 82 365 
<< m1 >>
rect 82 364 83 365 
<< m2 >>
rect 82 364 83 365 
<< m2 >>
rect 83 364 84 365 
<< m1 >>
rect 84 364 85 365 
<< m2 >>
rect 84 364 85 365 
<< m2c >>
rect 84 364 85 365 
<< m1 >>
rect 84 364 85 365 
<< m2 >>
rect 84 364 85 365 
<< m1 >>
rect 85 364 86 365 
<< m1 >>
rect 86 364 87 365 
<< m1 >>
rect 87 364 88 365 
<< m1 >>
rect 88 364 89 365 
<< m2 >>
rect 88 364 89 365 
<< m1 >>
rect 89 364 90 365 
<< m1 >>
rect 90 364 91 365 
<< m1 >>
rect 91 364 92 365 
<< m1 >>
rect 92 364 93 365 
<< m1 >>
rect 93 364 94 365 
<< m2 >>
rect 93 364 94 365 
<< m1 >>
rect 94 364 95 365 
<< m1 >>
rect 95 364 96 365 
<< m1 >>
rect 96 364 97 365 
<< m1 >>
rect 97 364 98 365 
<< m1 >>
rect 98 364 99 365 
<< m1 >>
rect 99 364 100 365 
<< m1 >>
rect 100 364 101 365 
<< m1 >>
rect 101 364 102 365 
<< m1 >>
rect 102 364 103 365 
<< m2 >>
rect 102 364 103 365 
<< m1 >>
rect 103 364 104 365 
<< m2 >>
rect 103 364 104 365 
<< m2 >>
rect 104 364 105 365 
<< m1 >>
rect 109 364 110 365 
<< m1 >>
rect 110 364 111 365 
<< m1 >>
rect 111 364 112 365 
<< m1 >>
rect 112 364 113 365 
<< m1 >>
rect 113 364 114 365 
<< m1 >>
rect 114 364 115 365 
<< m1 >>
rect 115 364 116 365 
<< m1 >>
rect 116 364 117 365 
<< m2 >>
rect 116 364 117 365 
<< m1 >>
rect 117 364 118 365 
<< m1 >>
rect 118 364 119 365 
<< m2 >>
rect 118 364 119 365 
<< m1 >>
rect 119 364 120 365 
<< m1 >>
rect 120 364 121 365 
<< m1 >>
rect 121 364 122 365 
<< m1 >>
rect 122 364 123 365 
<< m1 >>
rect 123 364 124 365 
<< m1 >>
rect 124 364 125 365 
<< m1 >>
rect 125 364 126 365 
<< m1 >>
rect 126 364 127 365 
<< m1 >>
rect 127 364 128 365 
<< m2 >>
rect 127 364 128 365 
<< m1 >>
rect 128 364 129 365 
<< m1 >>
rect 129 364 130 365 
<< m2 >>
rect 129 364 130 365 
<< m1 >>
rect 130 364 131 365 
<< m1 >>
rect 131 364 132 365 
<< m1 >>
rect 132 364 133 365 
<< m1 >>
rect 133 364 134 365 
<< m1 >>
rect 134 364 135 365 
<< m1 >>
rect 135 364 136 365 
<< m1 >>
rect 136 364 137 365 
<< m1 >>
rect 137 364 138 365 
<< m1 >>
rect 138 364 139 365 
<< m1 >>
rect 139 364 140 365 
<< m1 >>
rect 140 364 141 365 
<< m2 >>
rect 140 364 141 365 
<< m2c >>
rect 140 364 141 365 
<< m1 >>
rect 140 364 141 365 
<< m2 >>
rect 140 364 141 365 
<< m2 >>
rect 141 364 142 365 
<< m1 >>
rect 142 364 143 365 
<< m2 >>
rect 142 364 143 365 
<< m2 >>
rect 143 364 144 365 
<< m1 >>
rect 144 364 145 365 
<< m2 >>
rect 144 364 145 365 
<< m2c >>
rect 144 364 145 365 
<< m1 >>
rect 144 364 145 365 
<< m2 >>
rect 144 364 145 365 
<< m1 >>
rect 145 364 146 365 
<< m1 >>
rect 146 364 147 365 
<< m1 >>
rect 147 364 148 365 
<< m1 >>
rect 148 364 149 365 
<< m2 >>
rect 148 364 149 365 
<< m1 >>
rect 149 364 150 365 
<< m1 >>
rect 150 364 151 365 
<< m2 >>
rect 150 364 151 365 
<< m1 >>
rect 151 364 152 365 
<< m1 >>
rect 152 364 153 365 
<< m2 >>
rect 152 364 153 365 
<< m1 >>
rect 153 364 154 365 
<< m2 >>
rect 153 364 154 365 
<< m1 >>
rect 154 364 155 365 
<< m2 >>
rect 154 364 155 365 
<< m1 >>
rect 155 364 156 365 
<< m2 >>
rect 155 364 156 365 
<< m1 >>
rect 156 364 157 365 
<< m2 >>
rect 156 364 157 365 
<< m1 >>
rect 157 364 158 365 
<< m2 >>
rect 157 364 158 365 
<< m1 >>
rect 158 364 159 365 
<< m2 >>
rect 158 364 159 365 
<< m1 >>
rect 159 364 160 365 
<< m1 >>
rect 160 364 161 365 
<< m1 >>
rect 161 364 162 365 
<< m1 >>
rect 162 364 163 365 
<< m1 >>
rect 163 364 164 365 
<< m2 >>
rect 163 364 164 365 
<< m2 >>
rect 168 364 169 365 
<< m1 >>
rect 169 364 170 365 
<< m2 >>
rect 169 364 170 365 
<< m2 >>
rect 170 364 171 365 
<< m2 >>
rect 171 364 172 365 
<< m1 >>
rect 172 364 173 365 
<< m2 >>
rect 172 364 173 365 
<< m2 >>
rect 173 364 174 365 
<< m2 >>
rect 174 364 175 365 
<< m1 >>
rect 175 364 176 365 
<< m2 >>
rect 175 364 176 365 
<< m2 >>
rect 176 364 177 365 
<< m2 >>
rect 177 364 178 365 
<< m1 >>
rect 178 364 179 365 
<< m2 >>
rect 178 364 179 365 
<< m1 >>
rect 179 364 180 365 
<< m2 >>
rect 179 364 180 365 
<< m1 >>
rect 180 364 181 365 
<< m2 >>
rect 180 364 181 365 
<< m1 >>
rect 181 364 182 365 
<< m2 >>
rect 181 364 182 365 
<< m1 >>
rect 182 364 183 365 
<< m2 >>
rect 182 364 183 365 
<< m1 >>
rect 183 364 184 365 
<< m2 >>
rect 183 364 184 365 
<< m1 >>
rect 184 364 185 365 
<< m2 >>
rect 184 364 185 365 
<< m1 >>
rect 185 364 186 365 
<< m2 >>
rect 185 364 186 365 
<< m1 >>
rect 186 364 187 365 
<< m2 >>
rect 186 364 187 365 
<< m1 >>
rect 187 364 188 365 
<< m2 >>
rect 187 364 188 365 
<< m1 >>
rect 188 364 189 365 
<< m2 >>
rect 188 364 189 365 
<< m1 >>
rect 189 364 190 365 
<< m2 >>
rect 189 364 190 365 
<< m1 >>
rect 190 364 191 365 
<< m2 >>
rect 190 364 191 365 
<< m1 >>
rect 191 364 192 365 
<< m2 >>
rect 191 364 192 365 
<< m1 >>
rect 192 364 193 365 
<< m2 >>
rect 192 364 193 365 
<< m1 >>
rect 193 364 194 365 
<< m2 >>
rect 193 364 194 365 
<< m1 >>
rect 194 364 195 365 
<< m2 >>
rect 194 364 195 365 
<< m1 >>
rect 195 364 196 365 
<< m2 >>
rect 195 364 196 365 
<< m1 >>
rect 196 364 197 365 
<< m2 >>
rect 196 364 197 365 
<< m1 >>
rect 200 364 201 365 
<< m1 >>
rect 204 364 205 365 
<< m2 >>
rect 204 364 205 365 
<< m2c >>
rect 204 364 205 365 
<< m1 >>
rect 204 364 205 365 
<< m2 >>
rect 204 364 205 365 
<< m1 >>
rect 205 364 206 365 
<< m1 >>
rect 206 364 207 365 
<< m1 >>
rect 207 364 208 365 
<< m1 >>
rect 208 364 209 365 
<< m1 >>
rect 209 364 210 365 
<< m1 >>
rect 210 364 211 365 
<< m1 >>
rect 211 364 212 365 
<< m1 >>
rect 212 364 213 365 
<< m2 >>
rect 212 364 213 365 
<< m1 >>
rect 213 364 214 365 
<< m1 >>
rect 214 364 215 365 
<< m1 >>
rect 215 364 216 365 
<< m2 >>
rect 215 364 216 365 
<< m2c >>
rect 215 364 216 365 
<< m1 >>
rect 215 364 216 365 
<< m2 >>
rect 215 364 216 365 
<< m2 >>
rect 216 364 217 365 
<< m1 >>
rect 217 364 218 365 
<< m2 >>
rect 217 364 218 365 
<< m2 >>
rect 218 364 219 365 
<< m1 >>
rect 219 364 220 365 
<< m2 >>
rect 219 364 220 365 
<< m2c >>
rect 219 364 220 365 
<< m1 >>
rect 219 364 220 365 
<< m2 >>
rect 219 364 220 365 
<< m1 >>
rect 220 364 221 365 
<< m1 >>
rect 221 364 222 365 
<< m2 >>
rect 221 364 222 365 
<< m1 >>
rect 222 364 223 365 
<< m1 >>
rect 223 364 224 365 
<< m2 >>
rect 223 364 224 365 
<< m1 >>
rect 224 364 225 365 
<< m2 >>
rect 224 364 225 365 
<< m1 >>
rect 225 364 226 365 
<< m2 >>
rect 225 364 226 365 
<< m1 >>
rect 226 364 227 365 
<< m2 >>
rect 226 364 227 365 
<< m1 >>
rect 227 364 228 365 
<< m2 >>
rect 227 364 228 365 
<< m1 >>
rect 228 364 229 365 
<< m2 >>
rect 228 364 229 365 
<< m1 >>
rect 229 364 230 365 
<< m2 >>
rect 229 364 230 365 
<< m1 >>
rect 230 364 231 365 
<< m2 >>
rect 230 364 231 365 
<< m1 >>
rect 231 364 232 365 
<< m2 >>
rect 231 364 232 365 
<< m1 >>
rect 232 364 233 365 
<< m2 >>
rect 232 364 233 365 
<< m2 >>
rect 233 364 234 365 
<< m2 >>
rect 234 364 235 365 
<< m1 >>
rect 235 364 236 365 
<< m2 >>
rect 235 364 236 365 
<< m1 >>
rect 242 364 243 365 
<< m2 >>
rect 242 364 243 365 
<< m2c >>
rect 242 364 243 365 
<< m1 >>
rect 242 364 243 365 
<< m2 >>
rect 242 364 243 365 
<< m2 >>
rect 243 364 244 365 
<< m1 >>
rect 244 364 245 365 
<< m2 >>
rect 244 364 245 365 
<< m2 >>
rect 245 364 246 365 
<< m1 >>
rect 246 364 247 365 
<< m2 >>
rect 246 364 247 365 
<< m2c >>
rect 246 364 247 365 
<< m1 >>
rect 246 364 247 365 
<< m2 >>
rect 246 364 247 365 
<< m1 >>
rect 247 364 248 365 
<< m1 >>
rect 248 364 249 365 
<< m1 >>
rect 249 364 250 365 
<< m1 >>
rect 250 364 251 365 
<< m1 >>
rect 251 364 252 365 
<< m1 >>
rect 253 364 254 365 
<< m1 >>
rect 255 364 256 365 
<< m1 >>
rect 316 364 317 365 
<< m1 >>
rect 325 364 326 365 
<< m1 >>
rect 334 364 335 365 
<< m2 >>
rect 334 364 335 365 
<< m1 >>
rect 335 364 336 365 
<< m1 >>
rect 336 364 337 365 
<< m1 >>
rect 337 364 338 365 
<< m1 >>
rect 338 364 339 365 
<< m1 >>
rect 339 364 340 365 
<< m1 >>
rect 340 364 341 365 
<< m1 >>
rect 341 364 342 365 
<< m2 >>
rect 341 364 342 365 
<< m2c >>
rect 341 364 342 365 
<< m1 >>
rect 341 364 342 365 
<< m2 >>
rect 341 364 342 365 
<< m2 >>
rect 342 364 343 365 
<< m1 >>
rect 343 364 344 365 
<< m2 >>
rect 343 364 344 365 
<< m2 >>
rect 344 364 345 365 
<< m1 >>
rect 345 364 346 365 
<< m2 >>
rect 345 364 346 365 
<< m2c >>
rect 345 364 346 365 
<< m1 >>
rect 345 364 346 365 
<< m2 >>
rect 345 364 346 365 
<< m1 >>
rect 346 364 347 365 
<< m1 >>
rect 347 364 348 365 
<< m1 >>
rect 348 364 349 365 
<< m1 >>
rect 349 364 350 365 
<< m1 >>
rect 350 364 351 365 
<< m2 >>
rect 350 364 351 365 
<< m2c >>
rect 350 364 351 365 
<< m1 >>
rect 350 364 351 365 
<< m2 >>
rect 350 364 351 365 
<< m2 >>
rect 351 364 352 365 
<< m1 >>
rect 352 364 353 365 
<< m2 >>
rect 352 364 353 365 
<< m2 >>
rect 353 364 354 365 
<< m1 >>
rect 354 364 355 365 
<< m2 >>
rect 354 364 355 365 
<< m2c >>
rect 354 364 355 365 
<< m1 >>
rect 354 364 355 365 
<< m2 >>
rect 354 364 355 365 
<< m1 >>
rect 355 364 356 365 
<< m1 >>
rect 356 364 357 365 
<< m1 >>
rect 357 364 358 365 
<< m1 >>
rect 358 364 359 365 
<< m1 >>
rect 359 364 360 365 
<< m1 >>
rect 360 364 361 365 
<< m1 >>
rect 361 364 362 365 
<< m1 >>
rect 362 364 363 365 
<< m1 >>
rect 363 364 364 365 
<< m1 >>
rect 364 364 365 365 
<< m1 >>
rect 365 364 366 365 
<< m1 >>
rect 366 364 367 365 
<< m1 >>
rect 367 364 368 365 
<< m1 >>
rect 368 364 369 365 
<< m1 >>
rect 369 364 370 365 
<< m1 >>
rect 370 364 371 365 
<< m1 >>
rect 371 364 372 365 
<< m1 >>
rect 372 364 373 365 
<< m1 >>
rect 373 364 374 365 
<< m1 >>
rect 374 364 375 365 
<< m1 >>
rect 375 364 376 365 
<< m1 >>
rect 376 364 377 365 
<< m1 >>
rect 377 364 378 365 
<< m1 >>
rect 378 364 379 365 
<< m1 >>
rect 379 364 380 365 
<< m2 >>
rect 379 364 380 365 
<< m1 >>
rect 380 364 381 365 
<< m2 >>
rect 380 364 381 365 
<< m1 >>
rect 381 364 382 365 
<< m2 >>
rect 381 364 382 365 
<< m1 >>
rect 382 364 383 365 
<< m2 >>
rect 382 364 383 365 
<< m1 >>
rect 383 364 384 365 
<< m2 >>
rect 383 364 384 365 
<< m1 >>
rect 384 364 385 365 
<< m2 >>
rect 384 364 385 365 
<< m1 >>
rect 385 364 386 365 
<< m2 >>
rect 385 364 386 365 
<< m1 >>
rect 386 364 387 365 
<< m2 >>
rect 386 364 387 365 
<< m1 >>
rect 387 364 388 365 
<< m2 >>
rect 387 364 388 365 
<< m1 >>
rect 388 364 389 365 
<< m2 >>
rect 388 364 389 365 
<< m1 >>
rect 389 364 390 365 
<< m2 >>
rect 389 364 390 365 
<< m1 >>
rect 390 364 391 365 
<< m2 >>
rect 390 364 391 365 
<< m1 >>
rect 391 364 392 365 
<< m2 >>
rect 391 364 392 365 
<< m1 >>
rect 392 364 393 365 
<< m2 >>
rect 392 364 393 365 
<< m1 >>
rect 393 364 394 365 
<< m1 >>
rect 394 364 395 365 
<< m1 >>
rect 395 364 396 365 
<< m1 >>
rect 396 364 397 365 
<< m1 >>
rect 397 364 398 365 
<< m2 >>
rect 397 364 398 365 
<< m1 >>
rect 398 364 399 365 
<< m1 >>
rect 399 364 400 365 
<< m1 >>
rect 400 364 401 365 
<< m1 >>
rect 401 364 402 365 
<< m1 >>
rect 402 364 403 365 
<< m1 >>
rect 403 364 404 365 
<< m1 >>
rect 404 364 405 365 
<< m1 >>
rect 405 364 406 365 
<< m1 >>
rect 406 364 407 365 
<< m1 >>
rect 407 364 408 365 
<< m1 >>
rect 408 364 409 365 
<< m1 >>
rect 409 364 410 365 
<< m1 >>
rect 410 364 411 365 
<< m1 >>
rect 411 364 412 365 
<< m1 >>
rect 412 364 413 365 
<< m1 >>
rect 413 364 414 365 
<< m1 >>
rect 414 364 415 365 
<< m1 >>
rect 416 364 417 365 
<< m1 >>
rect 424 364 425 365 
<< m1 >>
rect 426 364 427 365 
<< m1 >>
rect 427 364 428 365 
<< m1 >>
rect 428 364 429 365 
<< m1 >>
rect 429 364 430 365 
<< m2 >>
rect 429 364 430 365 
<< m1 >>
rect 430 364 431 365 
<< m1 >>
rect 431 364 432 365 
<< m2 >>
rect 431 364 432 365 
<< m2c >>
rect 431 364 432 365 
<< m1 >>
rect 431 364 432 365 
<< m2 >>
rect 431 364 432 365 
<< m2 >>
rect 432 364 433 365 
<< m1 >>
rect 433 364 434 365 
<< m2 >>
rect 433 364 434 365 
<< m2 >>
rect 434 364 435 365 
<< m1 >>
rect 435 364 436 365 
<< m2 >>
rect 435 364 436 365 
<< m2 >>
rect 436 364 437 365 
<< m1 >>
rect 437 364 438 365 
<< m2 >>
rect 437 364 438 365 
<< m1 >>
rect 438 364 439 365 
<< m2 >>
rect 438 364 439 365 
<< m1 >>
rect 439 364 440 365 
<< m2 >>
rect 439 364 440 365 
<< m1 >>
rect 440 364 441 365 
<< m2 >>
rect 440 364 441 365 
<< m1 >>
rect 441 364 442 365 
<< m2 >>
rect 441 364 442 365 
<< m1 >>
rect 442 364 443 365 
<< m2 >>
rect 442 364 443 365 
<< m1 >>
rect 443 364 444 365 
<< m2 >>
rect 443 364 444 365 
<< m1 >>
rect 444 364 445 365 
<< m2 >>
rect 444 364 445 365 
<< m1 >>
rect 445 364 446 365 
<< m2 >>
rect 445 364 446 365 
<< m1 >>
rect 446 364 447 365 
<< m2 >>
rect 446 364 447 365 
<< m1 >>
rect 447 364 448 365 
<< m1 >>
rect 448 364 449 365 
<< m1 >>
rect 449 364 450 365 
<< m2 >>
rect 449 364 450 365 
<< m2c >>
rect 449 364 450 365 
<< m1 >>
rect 449 364 450 365 
<< m2 >>
rect 449 364 450 365 
<< m2 >>
rect 450 364 451 365 
<< m1 >>
rect 451 364 452 365 
<< m2 >>
rect 452 364 453 365 
<< m1 >>
rect 481 364 482 365 
<< m1 >>
rect 482 364 483 365 
<< m1 >>
rect 483 364 484 365 
<< m1 >>
rect 484 364 485 365 
<< m1 >>
rect 485 364 486 365 
<< m1 >>
rect 486 364 487 365 
<< m1 >>
rect 487 364 488 365 
<< m1 >>
rect 488 364 489 365 
<< m1 >>
rect 489 364 490 365 
<< m1 >>
rect 490 364 491 365 
<< m1 >>
rect 491 364 492 365 
<< m1 >>
rect 492 364 493 365 
<< m1 >>
rect 493 364 494 365 
<< m1 >>
rect 494 364 495 365 
<< m1 >>
rect 495 364 496 365 
<< m1 >>
rect 496 364 497 365 
<< m1 >>
rect 497 364 498 365 
<< m1 >>
rect 498 364 499 365 
<< m1 >>
rect 499 364 500 365 
<< m1 >>
rect 523 364 524 365 
<< m1 >>
rect 19 365 20 366 
<< m1 >>
rect 23 365 24 366 
<< m1 >>
rect 34 365 35 366 
<< m2 >>
rect 44 365 45 366 
<< m2 >>
rect 62 365 63 366 
<< m2 >>
rect 64 365 65 366 
<< m2 >>
rect 74 365 75 366 
<< m2 >>
rect 75 365 76 366 
<< m2 >>
rect 76 365 77 366 
<< m2 >>
rect 77 365 78 366 
<< m2 >>
rect 78 365 79 366 
<< m1 >>
rect 82 365 83 366 
<< m2 >>
rect 88 365 89 366 
<< m2 >>
rect 93 365 94 366 
<< m2 >>
rect 102 365 103 366 
<< m2 >>
rect 116 365 117 366 
<< m2 >>
rect 118 365 119 366 
<< m2 >>
rect 127 365 128 366 
<< m2 >>
rect 129 365 130 366 
<< m1 >>
rect 142 365 143 366 
<< m2 >>
rect 148 365 149 366 
<< m2 >>
rect 150 365 151 366 
<< m1 >>
rect 163 365 164 366 
<< m2 >>
rect 163 365 164 366 
<< m1 >>
rect 169 365 170 366 
<< m1 >>
rect 172 365 173 366 
<< m1 >>
rect 175 365 176 366 
<< m1 >>
rect 178 365 179 366 
<< m2 >>
rect 196 365 197 366 
<< m1 >>
rect 200 365 201 366 
<< m2 >>
rect 204 365 205 366 
<< m2 >>
rect 212 365 213 366 
<< m1 >>
rect 217 365 218 366 
<< m2 >>
rect 221 365 222 366 
<< m2 >>
rect 223 365 224 366 
<< m1 >>
rect 235 365 236 366 
<< m1 >>
rect 244 365 245 366 
<< m1 >>
rect 253 365 254 366 
<< m1 >>
rect 255 365 256 366 
<< m1 >>
rect 316 365 317 366 
<< m1 >>
rect 325 365 326 366 
<< m1 >>
rect 334 365 335 366 
<< m2 >>
rect 334 365 335 366 
<< m1 >>
rect 343 365 344 366 
<< m1 >>
rect 352 365 353 366 
<< m2 >>
rect 392 365 393 366 
<< m2 >>
rect 397 365 398 366 
<< m2 >>
rect 406 365 407 366 
<< m2 >>
rect 407 365 408 366 
<< m2 >>
rect 408 365 409 366 
<< m2 >>
rect 409 365 410 366 
<< m2 >>
rect 410 365 411 366 
<< m2 >>
rect 411 365 412 366 
<< m2 >>
rect 412 365 413 366 
<< m2 >>
rect 413 365 414 366 
<< m2 >>
rect 414 365 415 366 
<< m2 >>
rect 415 365 416 366 
<< m1 >>
rect 416 365 417 366 
<< m2 >>
rect 416 365 417 366 
<< m2 >>
rect 417 365 418 366 
<< m1 >>
rect 418 365 419 366 
<< m2 >>
rect 418 365 419 366 
<< m2c >>
rect 418 365 419 366 
<< m1 >>
rect 418 365 419 366 
<< m2 >>
rect 418 365 419 366 
<< m1 >>
rect 419 365 420 366 
<< m1 >>
rect 420 365 421 366 
<< m1 >>
rect 421 365 422 366 
<< m1 >>
rect 422 365 423 366 
<< m2 >>
rect 422 365 423 366 
<< m2c >>
rect 422 365 423 366 
<< m1 >>
rect 422 365 423 366 
<< m2 >>
rect 422 365 423 366 
<< m2 >>
rect 423 365 424 366 
<< m1 >>
rect 424 365 425 366 
<< m2 >>
rect 424 365 425 366 
<< m2 >>
rect 425 365 426 366 
<< m2 >>
rect 426 365 427 366 
<< m2 >>
rect 427 365 428 366 
<< m2 >>
rect 428 365 429 366 
<< m2 >>
rect 429 365 430 366 
<< m1 >>
rect 433 365 434 366 
<< m1 >>
rect 435 365 436 366 
<< m2 >>
rect 450 365 451 366 
<< m1 >>
rect 451 365 452 366 
<< m2 >>
rect 452 365 453 366 
<< m1 >>
rect 499 365 500 366 
<< m1 >>
rect 523 365 524 366 
<< m1 >>
rect 19 366 20 367 
<< m1 >>
rect 23 366 24 367 
<< m1 >>
rect 34 366 35 367 
<< m1 >>
rect 44 366 45 367 
<< m2 >>
rect 44 366 45 367 
<< m2c >>
rect 44 366 45 367 
<< m1 >>
rect 44 366 45 367 
<< m2 >>
rect 44 366 45 367 
<< m1 >>
rect 62 366 63 367 
<< m2 >>
rect 62 366 63 367 
<< m2c >>
rect 62 366 63 367 
<< m1 >>
rect 62 366 63 367 
<< m2 >>
rect 62 366 63 367 
<< m1 >>
rect 64 366 65 367 
<< m2 >>
rect 64 366 65 367 
<< m2c >>
rect 64 366 65 367 
<< m1 >>
rect 64 366 65 367 
<< m2 >>
rect 64 366 65 367 
<< m1 >>
rect 65 366 66 367 
<< m1 >>
rect 66 366 67 367 
<< m1 >>
rect 67 366 68 367 
<< m1 >>
rect 68 366 69 367 
<< m1 >>
rect 69 366 70 367 
<< m1 >>
rect 70 366 71 367 
<< m1 >>
rect 78 366 79 367 
<< m2 >>
rect 78 366 79 367 
<< m2c >>
rect 78 366 79 367 
<< m1 >>
rect 78 366 79 367 
<< m2 >>
rect 78 366 79 367 
<< m1 >>
rect 80 366 81 367 
<< m2 >>
rect 80 366 81 367 
<< m2c >>
rect 80 366 81 367 
<< m1 >>
rect 80 366 81 367 
<< m2 >>
rect 80 366 81 367 
<< m2 >>
rect 81 366 82 367 
<< m1 >>
rect 82 366 83 367 
<< m2 >>
rect 82 366 83 367 
<< m2 >>
rect 83 366 84 367 
<< m1 >>
rect 84 366 85 367 
<< m2 >>
rect 84 366 85 367 
<< m2c >>
rect 84 366 85 367 
<< m1 >>
rect 84 366 85 367 
<< m2 >>
rect 84 366 85 367 
<< m1 >>
rect 85 366 86 367 
<< m1 >>
rect 86 366 87 367 
<< m1 >>
rect 87 366 88 367 
<< m1 >>
rect 88 366 89 367 
<< m2 >>
rect 88 366 89 367 
<< m1 >>
rect 89 366 90 367 
<< m1 >>
rect 90 366 91 367 
<< m1 >>
rect 91 366 92 367 
<< m1 >>
rect 92 366 93 367 
<< m1 >>
rect 93 366 94 367 
<< m2 >>
rect 93 366 94 367 
<< m1 >>
rect 94 366 95 367 
<< m1 >>
rect 95 366 96 367 
<< m1 >>
rect 96 366 97 367 
<< m1 >>
rect 97 366 98 367 
<< m1 >>
rect 98 366 99 367 
<< m1 >>
rect 99 366 100 367 
<< m1 >>
rect 100 366 101 367 
<< m1 >>
rect 101 366 102 367 
<< m1 >>
rect 102 366 103 367 
<< m2 >>
rect 102 366 103 367 
<< m1 >>
rect 103 366 104 367 
<< m1 >>
rect 104 366 105 367 
<< m1 >>
rect 105 366 106 367 
<< m1 >>
rect 106 366 107 367 
<< m1 >>
rect 107 366 108 367 
<< m1 >>
rect 108 366 109 367 
<< m1 >>
rect 109 366 110 367 
<< m1 >>
rect 110 366 111 367 
<< m1 >>
rect 111 366 112 367 
<< m1 >>
rect 112 366 113 367 
<< m1 >>
rect 113 366 114 367 
<< m1 >>
rect 114 366 115 367 
<< m1 >>
rect 115 366 116 367 
<< m1 >>
rect 116 366 117 367 
<< m2 >>
rect 116 366 117 367 
<< m1 >>
rect 117 366 118 367 
<< m1 >>
rect 118 366 119 367 
<< m2 >>
rect 118 366 119 367 
<< m1 >>
rect 119 366 120 367 
<< m1 >>
rect 120 366 121 367 
<< m1 >>
rect 121 366 122 367 
<< m1 >>
rect 122 366 123 367 
<< m1 >>
rect 123 366 124 367 
<< m1 >>
rect 124 366 125 367 
<< m1 >>
rect 125 366 126 367 
<< m1 >>
rect 126 366 127 367 
<< m1 >>
rect 127 366 128 367 
<< m2 >>
rect 127 366 128 367 
<< m1 >>
rect 128 366 129 367 
<< m1 >>
rect 129 366 130 367 
<< m2 >>
rect 129 366 130 367 
<< m1 >>
rect 130 366 131 367 
<< m1 >>
rect 131 366 132 367 
<< m1 >>
rect 132 366 133 367 
<< m1 >>
rect 133 366 134 367 
<< m1 >>
rect 134 366 135 367 
<< m1 >>
rect 135 366 136 367 
<< m1 >>
rect 136 366 137 367 
<< m1 >>
rect 137 366 138 367 
<< m1 >>
rect 138 366 139 367 
<< m1 >>
rect 139 366 140 367 
<< m1 >>
rect 140 366 141 367 
<< m2 >>
rect 140 366 141 367 
<< m2c >>
rect 140 366 141 367 
<< m1 >>
rect 140 366 141 367 
<< m2 >>
rect 140 366 141 367 
<< m2 >>
rect 141 366 142 367 
<< m1 >>
rect 142 366 143 367 
<< m2 >>
rect 142 366 143 367 
<< m2 >>
rect 143 366 144 367 
<< m1 >>
rect 144 366 145 367 
<< m2 >>
rect 144 366 145 367 
<< m2c >>
rect 144 366 145 367 
<< m1 >>
rect 144 366 145 367 
<< m2 >>
rect 144 366 145 367 
<< m1 >>
rect 145 366 146 367 
<< m1 >>
rect 146 366 147 367 
<< m1 >>
rect 147 366 148 367 
<< m1 >>
rect 148 366 149 367 
<< m2 >>
rect 148 366 149 367 
<< m2c >>
rect 148 366 149 367 
<< m1 >>
rect 148 366 149 367 
<< m2 >>
rect 148 366 149 367 
<< m1 >>
rect 150 366 151 367 
<< m2 >>
rect 150 366 151 367 
<< m2c >>
rect 150 366 151 367 
<< m1 >>
rect 150 366 151 367 
<< m2 >>
rect 150 366 151 367 
<< m1 >>
rect 163 366 164 367 
<< m2 >>
rect 163 366 164 367 
<< m1 >>
rect 169 366 170 367 
<< m1 >>
rect 172 366 173 367 
<< m1 >>
rect 175 366 176 367 
<< m1 >>
rect 176 366 177 367 
<< m2 >>
rect 176 366 177 367 
<< m2c >>
rect 176 366 177 367 
<< m1 >>
rect 176 366 177 367 
<< m2 >>
rect 176 366 177 367 
<< m2 >>
rect 177 366 178 367 
<< m1 >>
rect 178 366 179 367 
<< m2 >>
rect 178 366 179 367 
<< m2 >>
rect 179 366 180 367 
<< m1 >>
rect 180 366 181 367 
<< m2 >>
rect 180 366 181 367 
<< m2c >>
rect 180 366 181 367 
<< m1 >>
rect 180 366 181 367 
<< m2 >>
rect 180 366 181 367 
<< m1 >>
rect 181 366 182 367 
<< m1 >>
rect 182 366 183 367 
<< m1 >>
rect 183 366 184 367 
<< m1 >>
rect 184 366 185 367 
<< m1 >>
rect 185 366 186 367 
<< m1 >>
rect 186 366 187 367 
<< m1 >>
rect 187 366 188 367 
<< m1 >>
rect 188 366 189 367 
<< m1 >>
rect 189 366 190 367 
<< m1 >>
rect 190 366 191 367 
<< m1 >>
rect 191 366 192 367 
<< m1 >>
rect 192 366 193 367 
<< m1 >>
rect 193 366 194 367 
<< m1 >>
rect 194 366 195 367 
<< m1 >>
rect 195 366 196 367 
<< m1 >>
rect 196 366 197 367 
<< m2 >>
rect 196 366 197 367 
<< m1 >>
rect 197 366 198 367 
<< m1 >>
rect 198 366 199 367 
<< m2 >>
rect 198 366 199 367 
<< m2c >>
rect 198 366 199 367 
<< m1 >>
rect 198 366 199 367 
<< m2 >>
rect 198 366 199 367 
<< m2 >>
rect 199 366 200 367 
<< m1 >>
rect 200 366 201 367 
<< m2 >>
rect 200 366 201 367 
<< m2 >>
rect 201 366 202 367 
<< m1 >>
rect 202 366 203 367 
<< m2 >>
rect 202 366 203 367 
<< m2c >>
rect 202 366 203 367 
<< m1 >>
rect 202 366 203 367 
<< m2 >>
rect 202 366 203 367 
<< m1 >>
rect 203 366 204 367 
<< m1 >>
rect 204 366 205 367 
<< m2 >>
rect 204 366 205 367 
<< m1 >>
rect 205 366 206 367 
<< m1 >>
rect 206 366 207 367 
<< m1 >>
rect 207 366 208 367 
<< m1 >>
rect 208 366 209 367 
<< m1 >>
rect 209 366 210 367 
<< m1 >>
rect 210 366 211 367 
<< m1 >>
rect 211 366 212 367 
<< m1 >>
rect 212 366 213 367 
<< m2 >>
rect 212 366 213 367 
<< m1 >>
rect 213 366 214 367 
<< m1 >>
rect 214 366 215 367 
<< m1 >>
rect 215 366 216 367 
<< m2 >>
rect 215 366 216 367 
<< m2c >>
rect 215 366 216 367 
<< m1 >>
rect 215 366 216 367 
<< m2 >>
rect 215 366 216 367 
<< m2 >>
rect 216 366 217 367 
<< m1 >>
rect 217 366 218 367 
<< m2 >>
rect 217 366 218 367 
<< m2 >>
rect 218 366 219 367 
<< m1 >>
rect 219 366 220 367 
<< m2 >>
rect 219 366 220 367 
<< m2c >>
rect 219 366 220 367 
<< m1 >>
rect 219 366 220 367 
<< m2 >>
rect 219 366 220 367 
<< m1 >>
rect 220 366 221 367 
<< m1 >>
rect 221 366 222 367 
<< m2 >>
rect 221 366 222 367 
<< m1 >>
rect 222 366 223 367 
<< m1 >>
rect 223 366 224 367 
<< m2 >>
rect 223 366 224 367 
<< m1 >>
rect 224 366 225 367 
<< m1 >>
rect 225 366 226 367 
<< m1 >>
rect 226 366 227 367 
<< m1 >>
rect 227 366 228 367 
<< m1 >>
rect 228 366 229 367 
<< m1 >>
rect 229 366 230 367 
<< m1 >>
rect 230 366 231 367 
<< m1 >>
rect 231 366 232 367 
<< m1 >>
rect 232 366 233 367 
<< m1 >>
rect 233 366 234 367 
<< m2 >>
rect 233 366 234 367 
<< m2c >>
rect 233 366 234 367 
<< m1 >>
rect 233 366 234 367 
<< m2 >>
rect 233 366 234 367 
<< m2 >>
rect 234 366 235 367 
<< m1 >>
rect 235 366 236 367 
<< m2 >>
rect 235 366 236 367 
<< m2 >>
rect 236 366 237 367 
<< m1 >>
rect 237 366 238 367 
<< m2 >>
rect 237 366 238 367 
<< m2c >>
rect 237 366 238 367 
<< m1 >>
rect 237 366 238 367 
<< m2 >>
rect 237 366 238 367 
<< m1 >>
rect 238 366 239 367 
<< m1 >>
rect 239 366 240 367 
<< m1 >>
rect 240 366 241 367 
<< m1 >>
rect 241 366 242 367 
<< m1 >>
rect 242 366 243 367 
<< m1 >>
rect 244 366 245 367 
<< m1 >>
rect 253 366 254 367 
<< m1 >>
rect 255 366 256 367 
<< m1 >>
rect 316 366 317 367 
<< m1 >>
rect 325 366 326 367 
<< m1 >>
rect 334 366 335 367 
<< m2 >>
rect 334 366 335 367 
<< m2 >>
rect 335 366 336 367 
<< m1 >>
rect 336 366 337 367 
<< m2 >>
rect 336 366 337 367 
<< m2c >>
rect 336 366 337 367 
<< m1 >>
rect 336 366 337 367 
<< m2 >>
rect 336 366 337 367 
<< m1 >>
rect 337 366 338 367 
<< m1 >>
rect 338 366 339 367 
<< m1 >>
rect 339 366 340 367 
<< m1 >>
rect 340 366 341 367 
<< m1 >>
rect 341 366 342 367 
<< m2 >>
rect 341 366 342 367 
<< m2c >>
rect 341 366 342 367 
<< m1 >>
rect 341 366 342 367 
<< m2 >>
rect 341 366 342 367 
<< m2 >>
rect 342 366 343 367 
<< m1 >>
rect 343 366 344 367 
<< m2 >>
rect 343 366 344 367 
<< m2 >>
rect 344 366 345 367 
<< m1 >>
rect 345 366 346 367 
<< m2 >>
rect 345 366 346 367 
<< m2c >>
rect 345 366 346 367 
<< m1 >>
rect 345 366 346 367 
<< m2 >>
rect 345 366 346 367 
<< m1 >>
rect 346 366 347 367 
<< m1 >>
rect 347 366 348 367 
<< m1 >>
rect 348 366 349 367 
<< m1 >>
rect 349 366 350 367 
<< m1 >>
rect 350 366 351 367 
<< m2 >>
rect 350 366 351 367 
<< m2c >>
rect 350 366 351 367 
<< m1 >>
rect 350 366 351 367 
<< m2 >>
rect 350 366 351 367 
<< m2 >>
rect 351 366 352 367 
<< m1 >>
rect 352 366 353 367 
<< m2 >>
rect 352 366 353 367 
<< m2 >>
rect 353 366 354 367 
<< m2 >>
rect 354 366 355 367 
<< m2 >>
rect 355 366 356 367 
<< m2 >>
rect 356 366 357 367 
<< m2 >>
rect 392 366 393 367 
<< m2 >>
rect 397 366 398 367 
<< m2 >>
rect 406 366 407 367 
<< m1 >>
rect 416 366 417 367 
<< m1 >>
rect 424 366 425 367 
<< m1 >>
rect 433 366 434 367 
<< m1 >>
rect 435 366 436 367 
<< m2 >>
rect 450 366 451 367 
<< m1 >>
rect 451 366 452 367 
<< m2 >>
rect 452 366 453 367 
<< m2 >>
rect 453 366 454 367 
<< m2 >>
rect 454 366 455 367 
<< m2 >>
rect 455 366 456 367 
<< m2 >>
rect 456 366 457 367 
<< m2 >>
rect 457 366 458 367 
<< m1 >>
rect 499 366 500 367 
<< m1 >>
rect 523 366 524 367 
<< m1 >>
rect 19 367 20 368 
<< m1 >>
rect 23 367 24 368 
<< m1 >>
rect 34 367 35 368 
<< m1 >>
rect 44 367 45 368 
<< m1 >>
rect 62 367 63 368 
<< m1 >>
rect 70 367 71 368 
<< m1 >>
rect 78 367 79 368 
<< m1 >>
rect 80 367 81 368 
<< m1 >>
rect 82 367 83 368 
<< m2 >>
rect 88 367 89 368 
<< m2 >>
rect 89 367 90 368 
<< m2 >>
rect 90 367 91 368 
<< m2 >>
rect 91 367 92 368 
<< m2 >>
rect 93 367 94 368 
<< m2 >>
rect 102 367 103 368 
<< m2 >>
rect 116 367 117 368 
<< m2 >>
rect 118 367 119 368 
<< m2 >>
rect 127 367 128 368 
<< m2 >>
rect 129 367 130 368 
<< m1 >>
rect 142 367 143 368 
<< m1 >>
rect 150 367 151 368 
<< m1 >>
rect 156 367 157 368 
<< m1 >>
rect 157 367 158 368 
<< m1 >>
rect 158 367 159 368 
<< m1 >>
rect 159 367 160 368 
<< m1 >>
rect 160 367 161 368 
<< m1 >>
rect 163 367 164 368 
<< m2 >>
rect 163 367 164 368 
<< m1 >>
rect 169 367 170 368 
<< m1 >>
rect 172 367 173 368 
<< m1 >>
rect 178 367 179 368 
<< m2 >>
rect 196 367 197 368 
<< m1 >>
rect 200 367 201 368 
<< m2 >>
rect 204 367 205 368 
<< m2 >>
rect 208 367 209 368 
<< m2 >>
rect 209 367 210 368 
<< m2 >>
rect 210 367 211 368 
<< m2 >>
rect 211 367 212 368 
<< m2 >>
rect 212 367 213 368 
<< m1 >>
rect 217 367 218 368 
<< m2 >>
rect 221 367 222 368 
<< m2 >>
rect 223 367 224 368 
<< m1 >>
rect 235 367 236 368 
<< m1 >>
rect 242 367 243 368 
<< m2 >>
rect 242 367 243 368 
<< m2c >>
rect 242 367 243 368 
<< m1 >>
rect 242 367 243 368 
<< m2 >>
rect 242 367 243 368 
<< m2 >>
rect 243 367 244 368 
<< m1 >>
rect 244 367 245 368 
<< m2 >>
rect 244 367 245 368 
<< m2 >>
rect 245 367 246 368 
<< m1 >>
rect 246 367 247 368 
<< m2 >>
rect 246 367 247 368 
<< m2c >>
rect 246 367 247 368 
<< m1 >>
rect 246 367 247 368 
<< m2 >>
rect 246 367 247 368 
<< m1 >>
rect 247 367 248 368 
<< m1 >>
rect 248 367 249 368 
<< m1 >>
rect 249 367 250 368 
<< m1 >>
rect 250 367 251 368 
<< m1 >>
rect 251 367 252 368 
<< m2 >>
rect 251 367 252 368 
<< m2c >>
rect 251 367 252 368 
<< m1 >>
rect 251 367 252 368 
<< m2 >>
rect 251 367 252 368 
<< m2 >>
rect 252 367 253 368 
<< m1 >>
rect 253 367 254 368 
<< m2 >>
rect 253 367 254 368 
<< m2 >>
rect 254 367 255 368 
<< m1 >>
rect 255 367 256 368 
<< m2 >>
rect 255 367 256 368 
<< m2 >>
rect 256 367 257 368 
<< m1 >>
rect 257 367 258 368 
<< m2 >>
rect 257 367 258 368 
<< m2c >>
rect 257 367 258 368 
<< m1 >>
rect 257 367 258 368 
<< m2 >>
rect 257 367 258 368 
<< m1 >>
rect 258 367 259 368 
<< m1 >>
rect 259 367 260 368 
<< m1 >>
rect 260 367 261 368 
<< m1 >>
rect 261 367 262 368 
<< m1 >>
rect 262 367 263 368 
<< m1 >>
rect 263 367 264 368 
<< m1 >>
rect 264 367 265 368 
<< m1 >>
rect 265 367 266 368 
<< m1 >>
rect 266 367 267 368 
<< m1 >>
rect 267 367 268 368 
<< m1 >>
rect 268 367 269 368 
<< m1 >>
rect 316 367 317 368 
<< m1 >>
rect 325 367 326 368 
<< m1 >>
rect 334 367 335 368 
<< m1 >>
rect 343 367 344 368 
<< m1 >>
rect 352 367 353 368 
<< m1 >>
rect 353 367 354 368 
<< m1 >>
rect 354 367 355 368 
<< m1 >>
rect 355 367 356 368 
<< m1 >>
rect 356 367 357 368 
<< m2 >>
rect 356 367 357 368 
<< m1 >>
rect 357 367 358 368 
<< m1 >>
rect 358 367 359 368 
<< m1 >>
rect 359 367 360 368 
<< m1 >>
rect 360 367 361 368 
<< m1 >>
rect 361 367 362 368 
<< m1 >>
rect 362 367 363 368 
<< m1 >>
rect 363 367 364 368 
<< m1 >>
rect 364 367 365 368 
<< m1 >>
rect 365 367 366 368 
<< m1 >>
rect 366 367 367 368 
<< m1 >>
rect 367 367 368 368 
<< m1 >>
rect 368 367 369 368 
<< m1 >>
rect 369 367 370 368 
<< m1 >>
rect 370 367 371 368 
<< m1 >>
rect 371 367 372 368 
<< m1 >>
rect 372 367 373 368 
<< m1 >>
rect 373 367 374 368 
<< m1 >>
rect 374 367 375 368 
<< m1 >>
rect 375 367 376 368 
<< m1 >>
rect 376 367 377 368 
<< m1 >>
rect 377 367 378 368 
<< m1 >>
rect 378 367 379 368 
<< m1 >>
rect 379 367 380 368 
<< m1 >>
rect 380 367 381 368 
<< m1 >>
rect 381 367 382 368 
<< m1 >>
rect 382 367 383 368 
<< m1 >>
rect 383 367 384 368 
<< m1 >>
rect 384 367 385 368 
<< m1 >>
rect 385 367 386 368 
<< m1 >>
rect 386 367 387 368 
<< m1 >>
rect 387 367 388 368 
<< m1 >>
rect 388 367 389 368 
<< m1 >>
rect 389 367 390 368 
<< m1 >>
rect 390 367 391 368 
<< m1 >>
rect 391 367 392 368 
<< m1 >>
rect 392 367 393 368 
<< m2 >>
rect 392 367 393 368 
<< m1 >>
rect 393 367 394 368 
<< m1 >>
rect 394 367 395 368 
<< m1 >>
rect 395 367 396 368 
<< m1 >>
rect 396 367 397 368 
<< m1 >>
rect 397 367 398 368 
<< m2 >>
rect 397 367 398 368 
<< m1 >>
rect 398 367 399 368 
<< m1 >>
rect 399 367 400 368 
<< m1 >>
rect 400 367 401 368 
<< m1 >>
rect 401 367 402 368 
<< m1 >>
rect 402 367 403 368 
<< m1 >>
rect 403 367 404 368 
<< m1 >>
rect 404 367 405 368 
<< m1 >>
rect 405 367 406 368 
<< m1 >>
rect 406 367 407 368 
<< m2 >>
rect 406 367 407 368 
<< m1 >>
rect 407 367 408 368 
<< m1 >>
rect 408 367 409 368 
<< m1 >>
rect 409 367 410 368 
<< m1 >>
rect 410 367 411 368 
<< m1 >>
rect 411 367 412 368 
<< m1 >>
rect 412 367 413 368 
<< m1 >>
rect 416 367 417 368 
<< m1 >>
rect 424 367 425 368 
<< m1 >>
rect 425 367 426 368 
<< m1 >>
rect 426 367 427 368 
<< m1 >>
rect 427 367 428 368 
<< m1 >>
rect 428 367 429 368 
<< m1 >>
rect 429 367 430 368 
<< m1 >>
rect 430 367 431 368 
<< m1 >>
rect 433 367 434 368 
<< m1 >>
rect 435 367 436 368 
<< m2 >>
rect 450 367 451 368 
<< m1 >>
rect 451 367 452 368 
<< m1 >>
rect 453 367 454 368 
<< m1 >>
rect 454 367 455 368 
<< m1 >>
rect 455 367 456 368 
<< m1 >>
rect 456 367 457 368 
<< m1 >>
rect 457 367 458 368 
<< m2 >>
rect 457 367 458 368 
<< m1 >>
rect 458 367 459 368 
<< m1 >>
rect 459 367 460 368 
<< m1 >>
rect 460 367 461 368 
<< m1 >>
rect 461 367 462 368 
<< m1 >>
rect 462 367 463 368 
<< m1 >>
rect 463 367 464 368 
<< m1 >>
rect 464 367 465 368 
<< m1 >>
rect 465 367 466 368 
<< m1 >>
rect 466 367 467 368 
<< m1 >>
rect 499 367 500 368 
<< m1 >>
rect 523 367 524 368 
<< m1 >>
rect 19 368 20 369 
<< m1 >>
rect 23 368 24 369 
<< m1 >>
rect 34 368 35 369 
<< m1 >>
rect 44 368 45 369 
<< m1 >>
rect 62 368 63 369 
<< m1 >>
rect 70 368 71 369 
<< m1 >>
rect 76 368 77 369 
<< m2 >>
rect 76 368 77 369 
<< m2c >>
rect 76 368 77 369 
<< m1 >>
rect 76 368 77 369 
<< m2 >>
rect 76 368 77 369 
<< m2 >>
rect 77 368 78 369 
<< m1 >>
rect 78 368 79 369 
<< m2 >>
rect 78 368 79 369 
<< m2 >>
rect 79 368 80 369 
<< m1 >>
rect 80 368 81 369 
<< m2 >>
rect 80 368 81 369 
<< m2c >>
rect 80 368 81 369 
<< m1 >>
rect 80 368 81 369 
<< m2 >>
rect 80 368 81 369 
<< m1 >>
rect 82 368 83 369 
<< m1 >>
rect 91 368 92 369 
<< m2 >>
rect 91 368 92 369 
<< m2c >>
rect 91 368 92 369 
<< m1 >>
rect 91 368 92 369 
<< m2 >>
rect 91 368 92 369 
<< m1 >>
rect 93 368 94 369 
<< m2 >>
rect 93 368 94 369 
<< m2c >>
rect 93 368 94 369 
<< m1 >>
rect 93 368 94 369 
<< m2 >>
rect 93 368 94 369 
<< m1 >>
rect 100 368 101 369 
<< m1 >>
rect 101 368 102 369 
<< m1 >>
rect 102 368 103 369 
<< m2 >>
rect 102 368 103 369 
<< m2c >>
rect 102 368 103 369 
<< m1 >>
rect 102 368 103 369 
<< m2 >>
rect 102 368 103 369 
<< m1 >>
rect 110 368 111 369 
<< m2 >>
rect 110 368 111 369 
<< m2c >>
rect 110 368 111 369 
<< m1 >>
rect 110 368 111 369 
<< m2 >>
rect 110 368 111 369 
<< m2 >>
rect 111 368 112 369 
<< m1 >>
rect 112 368 113 369 
<< m2 >>
rect 112 368 113 369 
<< m1 >>
rect 113 368 114 369 
<< m2 >>
rect 113 368 114 369 
<< m1 >>
rect 114 368 115 369 
<< m2 >>
rect 114 368 115 369 
<< m1 >>
rect 115 368 116 369 
<< m2 >>
rect 115 368 116 369 
<< m1 >>
rect 116 368 117 369 
<< m2 >>
rect 116 368 117 369 
<< m1 >>
rect 117 368 118 369 
<< m1 >>
rect 118 368 119 369 
<< m2 >>
rect 118 368 119 369 
<< m2c >>
rect 118 368 119 369 
<< m1 >>
rect 118 368 119 369 
<< m2 >>
rect 118 368 119 369 
<< m1 >>
rect 127 368 128 369 
<< m2 >>
rect 127 368 128 369 
<< m2c >>
rect 127 368 128 369 
<< m1 >>
rect 127 368 128 369 
<< m2 >>
rect 127 368 128 369 
<< m1 >>
rect 129 368 130 369 
<< m2 >>
rect 129 368 130 369 
<< m2c >>
rect 129 368 130 369 
<< m1 >>
rect 129 368 130 369 
<< m2 >>
rect 129 368 130 369 
<< m1 >>
rect 142 368 143 369 
<< m1 >>
rect 148 368 149 369 
<< m2 >>
rect 148 368 149 369 
<< m2c >>
rect 148 368 149 369 
<< m1 >>
rect 148 368 149 369 
<< m2 >>
rect 148 368 149 369 
<< m2 >>
rect 149 368 150 369 
<< m1 >>
rect 150 368 151 369 
<< m2 >>
rect 150 368 151 369 
<< m2 >>
rect 151 368 152 369 
<< m1 >>
rect 152 368 153 369 
<< m2 >>
rect 152 368 153 369 
<< m2c >>
rect 152 368 153 369 
<< m1 >>
rect 152 368 153 369 
<< m2 >>
rect 152 368 153 369 
<< m1 >>
rect 153 368 154 369 
<< m1 >>
rect 154 368 155 369 
<< m1 >>
rect 155 368 156 369 
<< m1 >>
rect 156 368 157 369 
<< m1 >>
rect 160 368 161 369 
<< m1 >>
rect 163 368 164 369 
<< m2 >>
rect 163 368 164 369 
<< m1 >>
rect 169 368 170 369 
<< m1 >>
rect 172 368 173 369 
<< m1 >>
rect 178 368 179 369 
<< m1 >>
rect 196 368 197 369 
<< m2 >>
rect 196 368 197 369 
<< m2c >>
rect 196 368 197 369 
<< m1 >>
rect 196 368 197 369 
<< m2 >>
rect 196 368 197 369 
<< m1 >>
rect 200 368 201 369 
<< m1 >>
rect 204 368 205 369 
<< m2 >>
rect 204 368 205 369 
<< m2c >>
rect 204 368 205 369 
<< m1 >>
rect 204 368 205 369 
<< m2 >>
rect 204 368 205 369 
<< m1 >>
rect 208 368 209 369 
<< m2 >>
rect 208 368 209 369 
<< m2c >>
rect 208 368 209 369 
<< m1 >>
rect 208 368 209 369 
<< m2 >>
rect 208 368 209 369 
<< m1 >>
rect 217 368 218 369 
<< m1 >>
rect 221 368 222 369 
<< m2 >>
rect 221 368 222 369 
<< m2c >>
rect 221 368 222 369 
<< m1 >>
rect 221 368 222 369 
<< m2 >>
rect 221 368 222 369 
<< m1 >>
rect 223 368 224 369 
<< m2 >>
rect 223 368 224 369 
<< m2c >>
rect 223 368 224 369 
<< m1 >>
rect 223 368 224 369 
<< m2 >>
rect 223 368 224 369 
<< m1 >>
rect 235 368 236 369 
<< m2 >>
rect 235 368 236 369 
<< m2c >>
rect 235 368 236 369 
<< m1 >>
rect 235 368 236 369 
<< m2 >>
rect 235 368 236 369 
<< m1 >>
rect 244 368 245 369 
<< m1 >>
rect 253 368 254 369 
<< m1 >>
rect 255 368 256 369 
<< m1 >>
rect 268 368 269 369 
<< m1 >>
rect 316 368 317 369 
<< m1 >>
rect 325 368 326 369 
<< m1 >>
rect 334 368 335 369 
<< m1 >>
rect 343 368 344 369 
<< m2 >>
rect 356 368 357 369 
<< m2 >>
rect 392 368 393 369 
<< m2 >>
rect 397 368 398 369 
<< m2 >>
rect 406 368 407 369 
<< m1 >>
rect 412 368 413 369 
<< m1 >>
rect 416 368 417 369 
<< m1 >>
rect 430 368 431 369 
<< m1 >>
rect 433 368 434 369 
<< m1 >>
rect 435 368 436 369 
<< m2 >>
rect 450 368 451 369 
<< m1 >>
rect 451 368 452 369 
<< m1 >>
rect 453 368 454 369 
<< m2 >>
rect 457 368 458 369 
<< m1 >>
rect 466 368 467 369 
<< m1 >>
rect 499 368 500 369 
<< m1 >>
rect 523 368 524 369 
<< m1 >>
rect 19 369 20 370 
<< m1 >>
rect 23 369 24 370 
<< m1 >>
rect 34 369 35 370 
<< m1 >>
rect 44 369 45 370 
<< m1 >>
rect 62 369 63 370 
<< m1 >>
rect 70 369 71 370 
<< m1 >>
rect 76 369 77 370 
<< m1 >>
rect 78 369 79 370 
<< m1 >>
rect 82 369 83 370 
<< m1 >>
rect 91 369 92 370 
<< m1 >>
rect 93 369 94 370 
<< m1 >>
rect 100 369 101 370 
<< m1 >>
rect 110 369 111 370 
<< m1 >>
rect 112 369 113 370 
<< m1 >>
rect 127 369 128 370 
<< m1 >>
rect 129 369 130 370 
<< m1 >>
rect 142 369 143 370 
<< m1 >>
rect 148 369 149 370 
<< m1 >>
rect 150 369 151 370 
<< m1 >>
rect 160 369 161 370 
<< m1 >>
rect 163 369 164 370 
<< m2 >>
rect 163 369 164 370 
<< m1 >>
rect 169 369 170 370 
<< m1 >>
rect 172 369 173 370 
<< m1 >>
rect 178 369 179 370 
<< m1 >>
rect 196 369 197 370 
<< m1 >>
rect 200 369 201 370 
<< m1 >>
rect 204 369 205 370 
<< m1 >>
rect 208 369 209 370 
<< m1 >>
rect 217 369 218 370 
<< m1 >>
rect 221 369 222 370 
<< m1 >>
rect 223 369 224 370 
<< m2 >>
rect 235 369 236 370 
<< m1 >>
rect 244 369 245 370 
<< m1 >>
rect 253 369 254 370 
<< m1 >>
rect 255 369 256 370 
<< m1 >>
rect 268 369 269 370 
<< m1 >>
rect 316 369 317 370 
<< m1 >>
rect 325 369 326 370 
<< m1 >>
rect 334 369 335 370 
<< m1 >>
rect 343 369 344 370 
<< m1 >>
rect 356 369 357 370 
<< m2 >>
rect 356 369 357 370 
<< m2c >>
rect 356 369 357 370 
<< m1 >>
rect 356 369 357 370 
<< m2 >>
rect 356 369 357 370 
<< m1 >>
rect 357 369 358 370 
<< m1 >>
rect 358 369 359 370 
<< m1 >>
rect 359 369 360 370 
<< m1 >>
rect 360 369 361 370 
<< m1 >>
rect 361 369 362 370 
<< m1 >>
rect 362 369 363 370 
<< m1 >>
rect 363 369 364 370 
<< m1 >>
rect 364 369 365 370 
<< m1 >>
rect 365 369 366 370 
<< m1 >>
rect 392 369 393 370 
<< m2 >>
rect 392 369 393 370 
<< m2c >>
rect 392 369 393 370 
<< m1 >>
rect 392 369 393 370 
<< m2 >>
rect 392 369 393 370 
<< m1 >>
rect 393 369 394 370 
<< m1 >>
rect 394 369 395 370 
<< m1 >>
rect 395 369 396 370 
<< m1 >>
rect 396 369 397 370 
<< m1 >>
rect 397 369 398 370 
<< m2 >>
rect 397 369 398 370 
<< m1 >>
rect 398 369 399 370 
<< m1 >>
rect 399 369 400 370 
<< m1 >>
rect 400 369 401 370 
<< m1 >>
rect 401 369 402 370 
<< m1 >>
rect 402 369 403 370 
<< m1 >>
rect 403 369 404 370 
<< m1 >>
rect 404 369 405 370 
<< m1 >>
rect 405 369 406 370 
<< m2 >>
rect 406 369 407 370 
<< m1 >>
rect 412 369 413 370 
<< m1 >>
rect 416 369 417 370 
<< m1 >>
rect 430 369 431 370 
<< m1 >>
rect 433 369 434 370 
<< m1 >>
rect 435 369 436 370 
<< m2 >>
rect 450 369 451 370 
<< m1 >>
rect 451 369 452 370 
<< m2 >>
rect 451 369 452 370 
<< m2 >>
rect 452 369 453 370 
<< m1 >>
rect 453 369 454 370 
<< m2 >>
rect 453 369 454 370 
<< m2 >>
rect 454 369 455 370 
<< m1 >>
rect 455 369 456 370 
<< m2 >>
rect 455 369 456 370 
<< m2c >>
rect 455 369 456 370 
<< m1 >>
rect 455 369 456 370 
<< m2 >>
rect 455 369 456 370 
<< m1 >>
rect 457 369 458 370 
<< m2 >>
rect 457 369 458 370 
<< m2c >>
rect 457 369 458 370 
<< m1 >>
rect 457 369 458 370 
<< m2 >>
rect 457 369 458 370 
<< m1 >>
rect 466 369 467 370 
<< m1 >>
rect 499 369 500 370 
<< m1 >>
rect 523 369 524 370 
<< m1 >>
rect 19 370 20 371 
<< m1 >>
rect 23 370 24 371 
<< m1 >>
rect 34 370 35 371 
<< m1 >>
rect 44 370 45 371 
<< m1 >>
rect 62 370 63 371 
<< m1 >>
rect 70 370 71 371 
<< m1 >>
rect 76 370 77 371 
<< m1 >>
rect 78 370 79 371 
<< m1 >>
rect 82 370 83 371 
<< m1 >>
rect 91 370 92 371 
<< m1 >>
rect 93 370 94 371 
<< m1 >>
rect 100 370 101 371 
<< m1 >>
rect 110 370 111 371 
<< m1 >>
rect 112 370 113 371 
<< m1 >>
rect 127 370 128 371 
<< m1 >>
rect 129 370 130 371 
<< m1 >>
rect 142 370 143 371 
<< m1 >>
rect 148 370 149 371 
<< m1 >>
rect 150 370 151 371 
<< m1 >>
rect 160 370 161 371 
<< m1 >>
rect 163 370 164 371 
<< m2 >>
rect 163 370 164 371 
<< m1 >>
rect 169 370 170 371 
<< m1 >>
rect 172 370 173 371 
<< m1 >>
rect 178 370 179 371 
<< m1 >>
rect 190 370 191 371 
<< m1 >>
rect 191 370 192 371 
<< m1 >>
rect 192 370 193 371 
<< m1 >>
rect 193 370 194 371 
<< m1 >>
rect 196 370 197 371 
<< m1 >>
rect 200 370 201 371 
<< m1 >>
rect 204 370 205 371 
<< m1 >>
rect 208 370 209 371 
<< m1 >>
rect 217 370 218 371 
<< m1 >>
rect 221 370 222 371 
<< m1 >>
rect 223 370 224 371 
<< m1 >>
rect 232 370 233 371 
<< m1 >>
rect 233 370 234 371 
<< m1 >>
rect 234 370 235 371 
<< m1 >>
rect 235 370 236 371 
<< m2 >>
rect 235 370 236 371 
<< m1 >>
rect 244 370 245 371 
<< m1 >>
rect 253 370 254 371 
<< m1 >>
rect 255 370 256 371 
<< m1 >>
rect 268 370 269 371 
<< m1 >>
rect 271 370 272 371 
<< m1 >>
rect 272 370 273 371 
<< m1 >>
rect 273 370 274 371 
<< m1 >>
rect 274 370 275 371 
<< m1 >>
rect 275 370 276 371 
<< m1 >>
rect 276 370 277 371 
<< m1 >>
rect 277 370 278 371 
<< m1 >>
rect 278 370 279 371 
<< m1 >>
rect 279 370 280 371 
<< m1 >>
rect 280 370 281 371 
<< m1 >>
rect 281 370 282 371 
<< m1 >>
rect 282 370 283 371 
<< m1 >>
rect 283 370 284 371 
<< m1 >>
rect 304 370 305 371 
<< m1 >>
rect 305 370 306 371 
<< m1 >>
rect 306 370 307 371 
<< m1 >>
rect 307 370 308 371 
<< m1 >>
rect 316 370 317 371 
<< m1 >>
rect 325 370 326 371 
<< m1 >>
rect 334 370 335 371 
<< m1 >>
rect 343 370 344 371 
<< m1 >>
rect 365 370 366 371 
<< m2 >>
rect 397 370 398 371 
<< m1 >>
rect 405 370 406 371 
<< m2 >>
rect 406 370 407 371 
<< m1 >>
rect 412 370 413 371 
<< m1 >>
rect 416 370 417 371 
<< m1 >>
rect 430 370 431 371 
<< m1 >>
rect 433 370 434 371 
<< m1 >>
rect 435 370 436 371 
<< m1 >>
rect 451 370 452 371 
<< m1 >>
rect 453 370 454 371 
<< m1 >>
rect 455 370 456 371 
<< m1 >>
rect 457 370 458 371 
<< m1 >>
rect 466 370 467 371 
<< m1 >>
rect 499 370 500 371 
<< m1 >>
rect 523 370 524 371 
<< m1 >>
rect 19 371 20 372 
<< m1 >>
rect 23 371 24 372 
<< m1 >>
rect 34 371 35 372 
<< m1 >>
rect 44 371 45 372 
<< m1 >>
rect 62 371 63 372 
<< m1 >>
rect 70 371 71 372 
<< m1 >>
rect 76 371 77 372 
<< m1 >>
rect 78 371 79 372 
<< m1 >>
rect 82 371 83 372 
<< m1 >>
rect 91 371 92 372 
<< m1 >>
rect 93 371 94 372 
<< m1 >>
rect 100 371 101 372 
<< m1 >>
rect 110 371 111 372 
<< m1 >>
rect 112 371 113 372 
<< m1 >>
rect 127 371 128 372 
<< m1 >>
rect 129 371 130 372 
<< m1 >>
rect 142 371 143 372 
<< m1 >>
rect 148 371 149 372 
<< m1 >>
rect 150 371 151 372 
<< m1 >>
rect 160 371 161 372 
<< m1 >>
rect 163 371 164 372 
<< m2 >>
rect 163 371 164 372 
<< m1 >>
rect 169 371 170 372 
<< m1 >>
rect 172 371 173 372 
<< m1 >>
rect 178 371 179 372 
<< m1 >>
rect 190 371 191 372 
<< m1 >>
rect 193 371 194 372 
<< m1 >>
rect 196 371 197 372 
<< m1 >>
rect 200 371 201 372 
<< m1 >>
rect 204 371 205 372 
<< m1 >>
rect 208 371 209 372 
<< m1 >>
rect 217 371 218 372 
<< m1 >>
rect 221 371 222 372 
<< m1 >>
rect 223 371 224 372 
<< m1 >>
rect 232 371 233 372 
<< m1 >>
rect 235 371 236 372 
<< m2 >>
rect 235 371 236 372 
<< m1 >>
rect 244 371 245 372 
<< m1 >>
rect 253 371 254 372 
<< m1 >>
rect 255 371 256 372 
<< m1 >>
rect 268 371 269 372 
<< m1 >>
rect 271 371 272 372 
<< m1 >>
rect 283 371 284 372 
<< m1 >>
rect 304 371 305 372 
<< m1 >>
rect 307 371 308 372 
<< m1 >>
rect 316 371 317 372 
<< m1 >>
rect 325 371 326 372 
<< m1 >>
rect 334 371 335 372 
<< m1 >>
rect 343 371 344 372 
<< m1 >>
rect 365 371 366 372 
<< m1 >>
rect 397 371 398 372 
<< m2 >>
rect 397 371 398 372 
<< m2c >>
rect 397 371 398 372 
<< m1 >>
rect 397 371 398 372 
<< m2 >>
rect 397 371 398 372 
<< m1 >>
rect 402 371 403 372 
<< m1 >>
rect 403 371 404 372 
<< m2 >>
rect 403 371 404 372 
<< m2c >>
rect 403 371 404 372 
<< m1 >>
rect 403 371 404 372 
<< m2 >>
rect 403 371 404 372 
<< m2 >>
rect 404 371 405 372 
<< m1 >>
rect 405 371 406 372 
<< m2 >>
rect 405 371 406 372 
<< m2 >>
rect 406 371 407 372 
<< m1 >>
rect 412 371 413 372 
<< m1 >>
rect 416 371 417 372 
<< m1 >>
rect 430 371 431 372 
<< m1 >>
rect 433 371 434 372 
<< m1 >>
rect 435 371 436 372 
<< m1 >>
rect 451 371 452 372 
<< m1 >>
rect 453 371 454 372 
<< m1 >>
rect 455 371 456 372 
<< m1 >>
rect 457 371 458 372 
<< m1 >>
rect 466 371 467 372 
<< m1 >>
rect 499 371 500 372 
<< m1 >>
rect 523 371 524 372 
<< pdiffusion >>
rect 12 372 13 373 
<< pdiffusion >>
rect 13 372 14 373 
<< pdiffusion >>
rect 14 372 15 373 
<< pdiffusion >>
rect 15 372 16 373 
<< pdiffusion >>
rect 16 372 17 373 
<< pdiffusion >>
rect 17 372 18 373 
<< m1 >>
rect 19 372 20 373 
<< m1 >>
rect 23 372 24 373 
<< pdiffusion >>
rect 30 372 31 373 
<< pdiffusion >>
rect 31 372 32 373 
<< pdiffusion >>
rect 32 372 33 373 
<< pdiffusion >>
rect 33 372 34 373 
<< m1 >>
rect 34 372 35 373 
<< pdiffusion >>
rect 34 372 35 373 
<< pdiffusion >>
rect 35 372 36 373 
<< m1 >>
rect 44 372 45 373 
<< pdiffusion >>
rect 48 372 49 373 
<< pdiffusion >>
rect 49 372 50 373 
<< pdiffusion >>
rect 50 372 51 373 
<< pdiffusion >>
rect 51 372 52 373 
<< pdiffusion >>
rect 52 372 53 373 
<< pdiffusion >>
rect 53 372 54 373 
<< m1 >>
rect 62 372 63 373 
<< pdiffusion >>
rect 66 372 67 373 
<< pdiffusion >>
rect 67 372 68 373 
<< pdiffusion >>
rect 68 372 69 373 
<< pdiffusion >>
rect 69 372 70 373 
<< m1 >>
rect 70 372 71 373 
<< pdiffusion >>
rect 70 372 71 373 
<< pdiffusion >>
rect 71 372 72 373 
<< m1 >>
rect 76 372 77 373 
<< m1 >>
rect 78 372 79 373 
<< m1 >>
rect 82 372 83 373 
<< pdiffusion >>
rect 84 372 85 373 
<< pdiffusion >>
rect 85 372 86 373 
<< pdiffusion >>
rect 86 372 87 373 
<< pdiffusion >>
rect 87 372 88 373 
<< pdiffusion >>
rect 88 372 89 373 
<< pdiffusion >>
rect 89 372 90 373 
<< m1 >>
rect 91 372 92 373 
<< m1 >>
rect 93 372 94 373 
<< m1 >>
rect 100 372 101 373 
<< pdiffusion >>
rect 102 372 103 373 
<< pdiffusion >>
rect 103 372 104 373 
<< pdiffusion >>
rect 104 372 105 373 
<< pdiffusion >>
rect 105 372 106 373 
<< pdiffusion >>
rect 106 372 107 373 
<< pdiffusion >>
rect 107 372 108 373 
<< m1 >>
rect 110 372 111 373 
<< m1 >>
rect 112 372 113 373 
<< pdiffusion >>
rect 120 372 121 373 
<< pdiffusion >>
rect 121 372 122 373 
<< pdiffusion >>
rect 122 372 123 373 
<< pdiffusion >>
rect 123 372 124 373 
<< pdiffusion >>
rect 124 372 125 373 
<< pdiffusion >>
rect 125 372 126 373 
<< m1 >>
rect 127 372 128 373 
<< m1 >>
rect 129 372 130 373 
<< pdiffusion >>
rect 138 372 139 373 
<< pdiffusion >>
rect 139 372 140 373 
<< pdiffusion >>
rect 140 372 141 373 
<< pdiffusion >>
rect 141 372 142 373 
<< m1 >>
rect 142 372 143 373 
<< pdiffusion >>
rect 142 372 143 373 
<< pdiffusion >>
rect 143 372 144 373 
<< m1 >>
rect 148 372 149 373 
<< m1 >>
rect 150 372 151 373 
<< pdiffusion >>
rect 156 372 157 373 
<< pdiffusion >>
rect 157 372 158 373 
<< pdiffusion >>
rect 158 372 159 373 
<< pdiffusion >>
rect 159 372 160 373 
<< m1 >>
rect 160 372 161 373 
<< pdiffusion >>
rect 160 372 161 373 
<< pdiffusion >>
rect 161 372 162 373 
<< m1 >>
rect 163 372 164 373 
<< m2 >>
rect 163 372 164 373 
<< m1 >>
rect 169 372 170 373 
<< m1 >>
rect 172 372 173 373 
<< pdiffusion >>
rect 174 372 175 373 
<< pdiffusion >>
rect 175 372 176 373 
<< pdiffusion >>
rect 176 372 177 373 
<< pdiffusion >>
rect 177 372 178 373 
<< m1 >>
rect 178 372 179 373 
<< pdiffusion >>
rect 178 372 179 373 
<< pdiffusion >>
rect 179 372 180 373 
<< m1 >>
rect 190 372 191 373 
<< pdiffusion >>
rect 192 372 193 373 
<< m1 >>
rect 193 372 194 373 
<< pdiffusion >>
rect 193 372 194 373 
<< pdiffusion >>
rect 194 372 195 373 
<< pdiffusion >>
rect 195 372 196 373 
<< m1 >>
rect 196 372 197 373 
<< pdiffusion >>
rect 196 372 197 373 
<< pdiffusion >>
rect 197 372 198 373 
<< m1 >>
rect 200 372 201 373 
<< m1 >>
rect 204 372 205 373 
<< m1 >>
rect 208 372 209 373 
<< pdiffusion >>
rect 210 372 211 373 
<< pdiffusion >>
rect 211 372 212 373 
<< pdiffusion >>
rect 212 372 213 373 
<< pdiffusion >>
rect 213 372 214 373 
<< pdiffusion >>
rect 214 372 215 373 
<< pdiffusion >>
rect 215 372 216 373 
<< m1 >>
rect 217 372 218 373 
<< m1 >>
rect 221 372 222 373 
<< m1 >>
rect 223 372 224 373 
<< pdiffusion >>
rect 228 372 229 373 
<< pdiffusion >>
rect 229 372 230 373 
<< pdiffusion >>
rect 230 372 231 373 
<< pdiffusion >>
rect 231 372 232 373 
<< m1 >>
rect 232 372 233 373 
<< pdiffusion >>
rect 232 372 233 373 
<< pdiffusion >>
rect 233 372 234 373 
<< m1 >>
rect 235 372 236 373 
<< m2 >>
rect 235 372 236 373 
<< m1 >>
rect 244 372 245 373 
<< pdiffusion >>
rect 246 372 247 373 
<< pdiffusion >>
rect 247 372 248 373 
<< pdiffusion >>
rect 248 372 249 373 
<< pdiffusion >>
rect 249 372 250 373 
<< pdiffusion >>
rect 250 372 251 373 
<< pdiffusion >>
rect 251 372 252 373 
<< m1 >>
rect 253 372 254 373 
<< m1 >>
rect 255 372 256 373 
<< pdiffusion >>
rect 264 372 265 373 
<< pdiffusion >>
rect 265 372 266 373 
<< pdiffusion >>
rect 266 372 267 373 
<< pdiffusion >>
rect 267 372 268 373 
<< m1 >>
rect 268 372 269 373 
<< pdiffusion >>
rect 268 372 269 373 
<< pdiffusion >>
rect 269 372 270 373 
<< m1 >>
rect 271 372 272 373 
<< pdiffusion >>
rect 282 372 283 373 
<< m1 >>
rect 283 372 284 373 
<< pdiffusion >>
rect 283 372 284 373 
<< pdiffusion >>
rect 284 372 285 373 
<< pdiffusion >>
rect 285 372 286 373 
<< pdiffusion >>
rect 286 372 287 373 
<< pdiffusion >>
rect 287 372 288 373 
<< pdiffusion >>
rect 300 372 301 373 
<< pdiffusion >>
rect 301 372 302 373 
<< pdiffusion >>
rect 302 372 303 373 
<< pdiffusion >>
rect 303 372 304 373 
<< m1 >>
rect 304 372 305 373 
<< pdiffusion >>
rect 304 372 305 373 
<< pdiffusion >>
rect 305 372 306 373 
<< m1 >>
rect 307 372 308 373 
<< m1 >>
rect 316 372 317 373 
<< pdiffusion >>
rect 318 372 319 373 
<< pdiffusion >>
rect 319 372 320 373 
<< pdiffusion >>
rect 320 372 321 373 
<< pdiffusion >>
rect 321 372 322 373 
<< pdiffusion >>
rect 322 372 323 373 
<< pdiffusion >>
rect 323 372 324 373 
<< m1 >>
rect 325 372 326 373 
<< m1 >>
rect 334 372 335 373 
<< pdiffusion >>
rect 336 372 337 373 
<< pdiffusion >>
rect 337 372 338 373 
<< pdiffusion >>
rect 338 372 339 373 
<< pdiffusion >>
rect 339 372 340 373 
<< pdiffusion >>
rect 340 372 341 373 
<< pdiffusion >>
rect 341 372 342 373 
<< m1 >>
rect 343 372 344 373 
<< pdiffusion >>
rect 354 372 355 373 
<< pdiffusion >>
rect 355 372 356 373 
<< pdiffusion >>
rect 356 372 357 373 
<< pdiffusion >>
rect 357 372 358 373 
<< pdiffusion >>
rect 358 372 359 373 
<< pdiffusion >>
rect 359 372 360 373 
<< m1 >>
rect 365 372 366 373 
<< pdiffusion >>
rect 372 372 373 373 
<< pdiffusion >>
rect 373 372 374 373 
<< pdiffusion >>
rect 374 372 375 373 
<< pdiffusion >>
rect 375 372 376 373 
<< pdiffusion >>
rect 376 372 377 373 
<< pdiffusion >>
rect 377 372 378 373 
<< pdiffusion >>
rect 390 372 391 373 
<< pdiffusion >>
rect 391 372 392 373 
<< pdiffusion >>
rect 392 372 393 373 
<< pdiffusion >>
rect 393 372 394 373 
<< pdiffusion >>
rect 394 372 395 373 
<< pdiffusion >>
rect 395 372 396 373 
<< m1 >>
rect 397 372 398 373 
<< m1 >>
rect 402 372 403 373 
<< m1 >>
rect 405 372 406 373 
<< pdiffusion >>
rect 408 372 409 373 
<< pdiffusion >>
rect 409 372 410 373 
<< pdiffusion >>
rect 410 372 411 373 
<< pdiffusion >>
rect 411 372 412 373 
<< m1 >>
rect 412 372 413 373 
<< pdiffusion >>
rect 412 372 413 373 
<< pdiffusion >>
rect 413 372 414 373 
<< m1 >>
rect 416 372 417 373 
<< pdiffusion >>
rect 426 372 427 373 
<< pdiffusion >>
rect 427 372 428 373 
<< pdiffusion >>
rect 428 372 429 373 
<< pdiffusion >>
rect 429 372 430 373 
<< m1 >>
rect 430 372 431 373 
<< pdiffusion >>
rect 430 372 431 373 
<< pdiffusion >>
rect 431 372 432 373 
<< m1 >>
rect 433 372 434 373 
<< m1 >>
rect 435 372 436 373 
<< pdiffusion >>
rect 444 372 445 373 
<< pdiffusion >>
rect 445 372 446 373 
<< pdiffusion >>
rect 446 372 447 373 
<< pdiffusion >>
rect 447 372 448 373 
<< pdiffusion >>
rect 448 372 449 373 
<< pdiffusion >>
rect 449 372 450 373 
<< m1 >>
rect 451 372 452 373 
<< m1 >>
rect 453 372 454 373 
<< m1 >>
rect 455 372 456 373 
<< m1 >>
rect 457 372 458 373 
<< pdiffusion >>
rect 462 372 463 373 
<< pdiffusion >>
rect 463 372 464 373 
<< pdiffusion >>
rect 464 372 465 373 
<< pdiffusion >>
rect 465 372 466 373 
<< m1 >>
rect 466 372 467 373 
<< pdiffusion >>
rect 466 372 467 373 
<< pdiffusion >>
rect 467 372 468 373 
<< pdiffusion >>
rect 498 372 499 373 
<< m1 >>
rect 499 372 500 373 
<< pdiffusion >>
rect 499 372 500 373 
<< pdiffusion >>
rect 500 372 501 373 
<< pdiffusion >>
rect 501 372 502 373 
<< pdiffusion >>
rect 502 372 503 373 
<< pdiffusion >>
rect 503 372 504 373 
<< pdiffusion >>
rect 516 372 517 373 
<< pdiffusion >>
rect 517 372 518 373 
<< pdiffusion >>
rect 518 372 519 373 
<< pdiffusion >>
rect 519 372 520 373 
<< pdiffusion >>
rect 520 372 521 373 
<< pdiffusion >>
rect 521 372 522 373 
<< m1 >>
rect 523 372 524 373 
<< pdiffusion >>
rect 12 373 13 374 
<< pdiffusion >>
rect 13 373 14 374 
<< pdiffusion >>
rect 14 373 15 374 
<< pdiffusion >>
rect 15 373 16 374 
<< pdiffusion >>
rect 16 373 17 374 
<< pdiffusion >>
rect 17 373 18 374 
<< m1 >>
rect 19 373 20 374 
<< m1 >>
rect 23 373 24 374 
<< pdiffusion >>
rect 30 373 31 374 
<< pdiffusion >>
rect 31 373 32 374 
<< pdiffusion >>
rect 32 373 33 374 
<< pdiffusion >>
rect 33 373 34 374 
<< pdiffusion >>
rect 34 373 35 374 
<< pdiffusion >>
rect 35 373 36 374 
<< m1 >>
rect 44 373 45 374 
<< pdiffusion >>
rect 48 373 49 374 
<< pdiffusion >>
rect 49 373 50 374 
<< pdiffusion >>
rect 50 373 51 374 
<< pdiffusion >>
rect 51 373 52 374 
<< pdiffusion >>
rect 52 373 53 374 
<< pdiffusion >>
rect 53 373 54 374 
<< m1 >>
rect 62 373 63 374 
<< pdiffusion >>
rect 66 373 67 374 
<< pdiffusion >>
rect 67 373 68 374 
<< pdiffusion >>
rect 68 373 69 374 
<< pdiffusion >>
rect 69 373 70 374 
<< pdiffusion >>
rect 70 373 71 374 
<< pdiffusion >>
rect 71 373 72 374 
<< m1 >>
rect 76 373 77 374 
<< m1 >>
rect 78 373 79 374 
<< m1 >>
rect 82 373 83 374 
<< pdiffusion >>
rect 84 373 85 374 
<< pdiffusion >>
rect 85 373 86 374 
<< pdiffusion >>
rect 86 373 87 374 
<< pdiffusion >>
rect 87 373 88 374 
<< pdiffusion >>
rect 88 373 89 374 
<< pdiffusion >>
rect 89 373 90 374 
<< m1 >>
rect 91 373 92 374 
<< m1 >>
rect 93 373 94 374 
<< m1 >>
rect 100 373 101 374 
<< pdiffusion >>
rect 102 373 103 374 
<< pdiffusion >>
rect 103 373 104 374 
<< pdiffusion >>
rect 104 373 105 374 
<< pdiffusion >>
rect 105 373 106 374 
<< pdiffusion >>
rect 106 373 107 374 
<< pdiffusion >>
rect 107 373 108 374 
<< m1 >>
rect 110 373 111 374 
<< m1 >>
rect 112 373 113 374 
<< pdiffusion >>
rect 120 373 121 374 
<< pdiffusion >>
rect 121 373 122 374 
<< pdiffusion >>
rect 122 373 123 374 
<< pdiffusion >>
rect 123 373 124 374 
<< pdiffusion >>
rect 124 373 125 374 
<< pdiffusion >>
rect 125 373 126 374 
<< m1 >>
rect 127 373 128 374 
<< m1 >>
rect 129 373 130 374 
<< pdiffusion >>
rect 138 373 139 374 
<< pdiffusion >>
rect 139 373 140 374 
<< pdiffusion >>
rect 140 373 141 374 
<< pdiffusion >>
rect 141 373 142 374 
<< pdiffusion >>
rect 142 373 143 374 
<< pdiffusion >>
rect 143 373 144 374 
<< m1 >>
rect 148 373 149 374 
<< m1 >>
rect 150 373 151 374 
<< pdiffusion >>
rect 156 373 157 374 
<< pdiffusion >>
rect 157 373 158 374 
<< pdiffusion >>
rect 158 373 159 374 
<< pdiffusion >>
rect 159 373 160 374 
<< pdiffusion >>
rect 160 373 161 374 
<< pdiffusion >>
rect 161 373 162 374 
<< m1 >>
rect 163 373 164 374 
<< m2 >>
rect 163 373 164 374 
<< m1 >>
rect 169 373 170 374 
<< m1 >>
rect 172 373 173 374 
<< pdiffusion >>
rect 174 373 175 374 
<< pdiffusion >>
rect 175 373 176 374 
<< pdiffusion >>
rect 176 373 177 374 
<< pdiffusion >>
rect 177 373 178 374 
<< pdiffusion >>
rect 178 373 179 374 
<< pdiffusion >>
rect 179 373 180 374 
<< m1 >>
rect 190 373 191 374 
<< pdiffusion >>
rect 192 373 193 374 
<< pdiffusion >>
rect 193 373 194 374 
<< pdiffusion >>
rect 194 373 195 374 
<< pdiffusion >>
rect 195 373 196 374 
<< pdiffusion >>
rect 196 373 197 374 
<< pdiffusion >>
rect 197 373 198 374 
<< m1 >>
rect 200 373 201 374 
<< m1 >>
rect 204 373 205 374 
<< m1 >>
rect 208 373 209 374 
<< pdiffusion >>
rect 210 373 211 374 
<< pdiffusion >>
rect 211 373 212 374 
<< pdiffusion >>
rect 212 373 213 374 
<< pdiffusion >>
rect 213 373 214 374 
<< pdiffusion >>
rect 214 373 215 374 
<< pdiffusion >>
rect 215 373 216 374 
<< m1 >>
rect 217 373 218 374 
<< m1 >>
rect 221 373 222 374 
<< m1 >>
rect 223 373 224 374 
<< pdiffusion >>
rect 228 373 229 374 
<< pdiffusion >>
rect 229 373 230 374 
<< pdiffusion >>
rect 230 373 231 374 
<< pdiffusion >>
rect 231 373 232 374 
<< pdiffusion >>
rect 232 373 233 374 
<< pdiffusion >>
rect 233 373 234 374 
<< m1 >>
rect 235 373 236 374 
<< m2 >>
rect 235 373 236 374 
<< m1 >>
rect 244 373 245 374 
<< pdiffusion >>
rect 246 373 247 374 
<< pdiffusion >>
rect 247 373 248 374 
<< pdiffusion >>
rect 248 373 249 374 
<< pdiffusion >>
rect 249 373 250 374 
<< pdiffusion >>
rect 250 373 251 374 
<< pdiffusion >>
rect 251 373 252 374 
<< m1 >>
rect 253 373 254 374 
<< m1 >>
rect 255 373 256 374 
<< pdiffusion >>
rect 264 373 265 374 
<< pdiffusion >>
rect 265 373 266 374 
<< pdiffusion >>
rect 266 373 267 374 
<< pdiffusion >>
rect 267 373 268 374 
<< pdiffusion >>
rect 268 373 269 374 
<< pdiffusion >>
rect 269 373 270 374 
<< m1 >>
rect 271 373 272 374 
<< pdiffusion >>
rect 282 373 283 374 
<< pdiffusion >>
rect 283 373 284 374 
<< pdiffusion >>
rect 284 373 285 374 
<< pdiffusion >>
rect 285 373 286 374 
<< pdiffusion >>
rect 286 373 287 374 
<< pdiffusion >>
rect 287 373 288 374 
<< pdiffusion >>
rect 300 373 301 374 
<< pdiffusion >>
rect 301 373 302 374 
<< pdiffusion >>
rect 302 373 303 374 
<< pdiffusion >>
rect 303 373 304 374 
<< pdiffusion >>
rect 304 373 305 374 
<< pdiffusion >>
rect 305 373 306 374 
<< m1 >>
rect 307 373 308 374 
<< m1 >>
rect 316 373 317 374 
<< pdiffusion >>
rect 318 373 319 374 
<< pdiffusion >>
rect 319 373 320 374 
<< pdiffusion >>
rect 320 373 321 374 
<< pdiffusion >>
rect 321 373 322 374 
<< pdiffusion >>
rect 322 373 323 374 
<< pdiffusion >>
rect 323 373 324 374 
<< m1 >>
rect 325 373 326 374 
<< m1 >>
rect 334 373 335 374 
<< pdiffusion >>
rect 336 373 337 374 
<< pdiffusion >>
rect 337 373 338 374 
<< pdiffusion >>
rect 338 373 339 374 
<< pdiffusion >>
rect 339 373 340 374 
<< pdiffusion >>
rect 340 373 341 374 
<< pdiffusion >>
rect 341 373 342 374 
<< m1 >>
rect 343 373 344 374 
<< pdiffusion >>
rect 354 373 355 374 
<< pdiffusion >>
rect 355 373 356 374 
<< pdiffusion >>
rect 356 373 357 374 
<< pdiffusion >>
rect 357 373 358 374 
<< pdiffusion >>
rect 358 373 359 374 
<< pdiffusion >>
rect 359 373 360 374 
<< m1 >>
rect 365 373 366 374 
<< pdiffusion >>
rect 372 373 373 374 
<< pdiffusion >>
rect 373 373 374 374 
<< pdiffusion >>
rect 374 373 375 374 
<< pdiffusion >>
rect 375 373 376 374 
<< pdiffusion >>
rect 376 373 377 374 
<< pdiffusion >>
rect 377 373 378 374 
<< pdiffusion >>
rect 390 373 391 374 
<< pdiffusion >>
rect 391 373 392 374 
<< pdiffusion >>
rect 392 373 393 374 
<< pdiffusion >>
rect 393 373 394 374 
<< pdiffusion >>
rect 394 373 395 374 
<< pdiffusion >>
rect 395 373 396 374 
<< m1 >>
rect 397 373 398 374 
<< m1 >>
rect 402 373 403 374 
<< m1 >>
rect 405 373 406 374 
<< pdiffusion >>
rect 408 373 409 374 
<< pdiffusion >>
rect 409 373 410 374 
<< pdiffusion >>
rect 410 373 411 374 
<< pdiffusion >>
rect 411 373 412 374 
<< pdiffusion >>
rect 412 373 413 374 
<< pdiffusion >>
rect 413 373 414 374 
<< m1 >>
rect 416 373 417 374 
<< pdiffusion >>
rect 426 373 427 374 
<< pdiffusion >>
rect 427 373 428 374 
<< pdiffusion >>
rect 428 373 429 374 
<< pdiffusion >>
rect 429 373 430 374 
<< pdiffusion >>
rect 430 373 431 374 
<< pdiffusion >>
rect 431 373 432 374 
<< m1 >>
rect 433 373 434 374 
<< m1 >>
rect 435 373 436 374 
<< pdiffusion >>
rect 444 373 445 374 
<< pdiffusion >>
rect 445 373 446 374 
<< pdiffusion >>
rect 446 373 447 374 
<< pdiffusion >>
rect 447 373 448 374 
<< pdiffusion >>
rect 448 373 449 374 
<< pdiffusion >>
rect 449 373 450 374 
<< m1 >>
rect 451 373 452 374 
<< m1 >>
rect 453 373 454 374 
<< m1 >>
rect 455 373 456 374 
<< m1 >>
rect 457 373 458 374 
<< pdiffusion >>
rect 462 373 463 374 
<< pdiffusion >>
rect 463 373 464 374 
<< pdiffusion >>
rect 464 373 465 374 
<< pdiffusion >>
rect 465 373 466 374 
<< pdiffusion >>
rect 466 373 467 374 
<< pdiffusion >>
rect 467 373 468 374 
<< pdiffusion >>
rect 498 373 499 374 
<< pdiffusion >>
rect 499 373 500 374 
<< pdiffusion >>
rect 500 373 501 374 
<< pdiffusion >>
rect 501 373 502 374 
<< pdiffusion >>
rect 502 373 503 374 
<< pdiffusion >>
rect 503 373 504 374 
<< pdiffusion >>
rect 516 373 517 374 
<< pdiffusion >>
rect 517 373 518 374 
<< pdiffusion >>
rect 518 373 519 374 
<< pdiffusion >>
rect 519 373 520 374 
<< pdiffusion >>
rect 520 373 521 374 
<< pdiffusion >>
rect 521 373 522 374 
<< m1 >>
rect 523 373 524 374 
<< pdiffusion >>
rect 12 374 13 375 
<< pdiffusion >>
rect 13 374 14 375 
<< pdiffusion >>
rect 14 374 15 375 
<< pdiffusion >>
rect 15 374 16 375 
<< pdiffusion >>
rect 16 374 17 375 
<< pdiffusion >>
rect 17 374 18 375 
<< m1 >>
rect 19 374 20 375 
<< m1 >>
rect 23 374 24 375 
<< pdiffusion >>
rect 30 374 31 375 
<< pdiffusion >>
rect 31 374 32 375 
<< pdiffusion >>
rect 32 374 33 375 
<< pdiffusion >>
rect 33 374 34 375 
<< pdiffusion >>
rect 34 374 35 375 
<< pdiffusion >>
rect 35 374 36 375 
<< m1 >>
rect 44 374 45 375 
<< pdiffusion >>
rect 48 374 49 375 
<< pdiffusion >>
rect 49 374 50 375 
<< pdiffusion >>
rect 50 374 51 375 
<< pdiffusion >>
rect 51 374 52 375 
<< pdiffusion >>
rect 52 374 53 375 
<< pdiffusion >>
rect 53 374 54 375 
<< m1 >>
rect 62 374 63 375 
<< pdiffusion >>
rect 66 374 67 375 
<< pdiffusion >>
rect 67 374 68 375 
<< pdiffusion >>
rect 68 374 69 375 
<< pdiffusion >>
rect 69 374 70 375 
<< pdiffusion >>
rect 70 374 71 375 
<< pdiffusion >>
rect 71 374 72 375 
<< m1 >>
rect 76 374 77 375 
<< m1 >>
rect 78 374 79 375 
<< m1 >>
rect 82 374 83 375 
<< pdiffusion >>
rect 84 374 85 375 
<< pdiffusion >>
rect 85 374 86 375 
<< pdiffusion >>
rect 86 374 87 375 
<< pdiffusion >>
rect 87 374 88 375 
<< pdiffusion >>
rect 88 374 89 375 
<< pdiffusion >>
rect 89 374 90 375 
<< m1 >>
rect 91 374 92 375 
<< m1 >>
rect 93 374 94 375 
<< m1 >>
rect 100 374 101 375 
<< pdiffusion >>
rect 102 374 103 375 
<< pdiffusion >>
rect 103 374 104 375 
<< pdiffusion >>
rect 104 374 105 375 
<< pdiffusion >>
rect 105 374 106 375 
<< pdiffusion >>
rect 106 374 107 375 
<< pdiffusion >>
rect 107 374 108 375 
<< m1 >>
rect 110 374 111 375 
<< m1 >>
rect 112 374 113 375 
<< pdiffusion >>
rect 120 374 121 375 
<< pdiffusion >>
rect 121 374 122 375 
<< pdiffusion >>
rect 122 374 123 375 
<< pdiffusion >>
rect 123 374 124 375 
<< pdiffusion >>
rect 124 374 125 375 
<< pdiffusion >>
rect 125 374 126 375 
<< m1 >>
rect 127 374 128 375 
<< m1 >>
rect 129 374 130 375 
<< pdiffusion >>
rect 138 374 139 375 
<< pdiffusion >>
rect 139 374 140 375 
<< pdiffusion >>
rect 140 374 141 375 
<< pdiffusion >>
rect 141 374 142 375 
<< pdiffusion >>
rect 142 374 143 375 
<< pdiffusion >>
rect 143 374 144 375 
<< m1 >>
rect 148 374 149 375 
<< m1 >>
rect 150 374 151 375 
<< pdiffusion >>
rect 156 374 157 375 
<< pdiffusion >>
rect 157 374 158 375 
<< pdiffusion >>
rect 158 374 159 375 
<< pdiffusion >>
rect 159 374 160 375 
<< pdiffusion >>
rect 160 374 161 375 
<< pdiffusion >>
rect 161 374 162 375 
<< m1 >>
rect 163 374 164 375 
<< m2 >>
rect 163 374 164 375 
<< m1 >>
rect 169 374 170 375 
<< m1 >>
rect 172 374 173 375 
<< pdiffusion >>
rect 174 374 175 375 
<< pdiffusion >>
rect 175 374 176 375 
<< pdiffusion >>
rect 176 374 177 375 
<< pdiffusion >>
rect 177 374 178 375 
<< pdiffusion >>
rect 178 374 179 375 
<< pdiffusion >>
rect 179 374 180 375 
<< m1 >>
rect 190 374 191 375 
<< pdiffusion >>
rect 192 374 193 375 
<< pdiffusion >>
rect 193 374 194 375 
<< pdiffusion >>
rect 194 374 195 375 
<< pdiffusion >>
rect 195 374 196 375 
<< pdiffusion >>
rect 196 374 197 375 
<< pdiffusion >>
rect 197 374 198 375 
<< m1 >>
rect 200 374 201 375 
<< m1 >>
rect 204 374 205 375 
<< m1 >>
rect 208 374 209 375 
<< pdiffusion >>
rect 210 374 211 375 
<< pdiffusion >>
rect 211 374 212 375 
<< pdiffusion >>
rect 212 374 213 375 
<< pdiffusion >>
rect 213 374 214 375 
<< pdiffusion >>
rect 214 374 215 375 
<< pdiffusion >>
rect 215 374 216 375 
<< m1 >>
rect 217 374 218 375 
<< m1 >>
rect 221 374 222 375 
<< m1 >>
rect 223 374 224 375 
<< pdiffusion >>
rect 228 374 229 375 
<< pdiffusion >>
rect 229 374 230 375 
<< pdiffusion >>
rect 230 374 231 375 
<< pdiffusion >>
rect 231 374 232 375 
<< pdiffusion >>
rect 232 374 233 375 
<< pdiffusion >>
rect 233 374 234 375 
<< m1 >>
rect 235 374 236 375 
<< m2 >>
rect 235 374 236 375 
<< m1 >>
rect 244 374 245 375 
<< pdiffusion >>
rect 246 374 247 375 
<< pdiffusion >>
rect 247 374 248 375 
<< pdiffusion >>
rect 248 374 249 375 
<< pdiffusion >>
rect 249 374 250 375 
<< pdiffusion >>
rect 250 374 251 375 
<< pdiffusion >>
rect 251 374 252 375 
<< m1 >>
rect 253 374 254 375 
<< m1 >>
rect 255 374 256 375 
<< pdiffusion >>
rect 264 374 265 375 
<< pdiffusion >>
rect 265 374 266 375 
<< pdiffusion >>
rect 266 374 267 375 
<< pdiffusion >>
rect 267 374 268 375 
<< pdiffusion >>
rect 268 374 269 375 
<< pdiffusion >>
rect 269 374 270 375 
<< m1 >>
rect 271 374 272 375 
<< pdiffusion >>
rect 282 374 283 375 
<< pdiffusion >>
rect 283 374 284 375 
<< pdiffusion >>
rect 284 374 285 375 
<< pdiffusion >>
rect 285 374 286 375 
<< pdiffusion >>
rect 286 374 287 375 
<< pdiffusion >>
rect 287 374 288 375 
<< pdiffusion >>
rect 300 374 301 375 
<< pdiffusion >>
rect 301 374 302 375 
<< pdiffusion >>
rect 302 374 303 375 
<< pdiffusion >>
rect 303 374 304 375 
<< pdiffusion >>
rect 304 374 305 375 
<< pdiffusion >>
rect 305 374 306 375 
<< m1 >>
rect 307 374 308 375 
<< m1 >>
rect 316 374 317 375 
<< pdiffusion >>
rect 318 374 319 375 
<< pdiffusion >>
rect 319 374 320 375 
<< pdiffusion >>
rect 320 374 321 375 
<< pdiffusion >>
rect 321 374 322 375 
<< pdiffusion >>
rect 322 374 323 375 
<< pdiffusion >>
rect 323 374 324 375 
<< m1 >>
rect 325 374 326 375 
<< m1 >>
rect 334 374 335 375 
<< pdiffusion >>
rect 336 374 337 375 
<< pdiffusion >>
rect 337 374 338 375 
<< pdiffusion >>
rect 338 374 339 375 
<< pdiffusion >>
rect 339 374 340 375 
<< pdiffusion >>
rect 340 374 341 375 
<< pdiffusion >>
rect 341 374 342 375 
<< m1 >>
rect 343 374 344 375 
<< pdiffusion >>
rect 354 374 355 375 
<< pdiffusion >>
rect 355 374 356 375 
<< pdiffusion >>
rect 356 374 357 375 
<< pdiffusion >>
rect 357 374 358 375 
<< pdiffusion >>
rect 358 374 359 375 
<< pdiffusion >>
rect 359 374 360 375 
<< m1 >>
rect 365 374 366 375 
<< pdiffusion >>
rect 372 374 373 375 
<< pdiffusion >>
rect 373 374 374 375 
<< pdiffusion >>
rect 374 374 375 375 
<< pdiffusion >>
rect 375 374 376 375 
<< pdiffusion >>
rect 376 374 377 375 
<< pdiffusion >>
rect 377 374 378 375 
<< pdiffusion >>
rect 390 374 391 375 
<< pdiffusion >>
rect 391 374 392 375 
<< pdiffusion >>
rect 392 374 393 375 
<< pdiffusion >>
rect 393 374 394 375 
<< pdiffusion >>
rect 394 374 395 375 
<< pdiffusion >>
rect 395 374 396 375 
<< m1 >>
rect 397 374 398 375 
<< m1 >>
rect 402 374 403 375 
<< m1 >>
rect 405 374 406 375 
<< pdiffusion >>
rect 408 374 409 375 
<< pdiffusion >>
rect 409 374 410 375 
<< pdiffusion >>
rect 410 374 411 375 
<< pdiffusion >>
rect 411 374 412 375 
<< pdiffusion >>
rect 412 374 413 375 
<< pdiffusion >>
rect 413 374 414 375 
<< m1 >>
rect 416 374 417 375 
<< pdiffusion >>
rect 426 374 427 375 
<< pdiffusion >>
rect 427 374 428 375 
<< pdiffusion >>
rect 428 374 429 375 
<< pdiffusion >>
rect 429 374 430 375 
<< pdiffusion >>
rect 430 374 431 375 
<< pdiffusion >>
rect 431 374 432 375 
<< m1 >>
rect 433 374 434 375 
<< m1 >>
rect 435 374 436 375 
<< pdiffusion >>
rect 444 374 445 375 
<< pdiffusion >>
rect 445 374 446 375 
<< pdiffusion >>
rect 446 374 447 375 
<< pdiffusion >>
rect 447 374 448 375 
<< pdiffusion >>
rect 448 374 449 375 
<< pdiffusion >>
rect 449 374 450 375 
<< m1 >>
rect 451 374 452 375 
<< m1 >>
rect 453 374 454 375 
<< m1 >>
rect 455 374 456 375 
<< m1 >>
rect 457 374 458 375 
<< pdiffusion >>
rect 462 374 463 375 
<< pdiffusion >>
rect 463 374 464 375 
<< pdiffusion >>
rect 464 374 465 375 
<< pdiffusion >>
rect 465 374 466 375 
<< pdiffusion >>
rect 466 374 467 375 
<< pdiffusion >>
rect 467 374 468 375 
<< pdiffusion >>
rect 498 374 499 375 
<< pdiffusion >>
rect 499 374 500 375 
<< pdiffusion >>
rect 500 374 501 375 
<< pdiffusion >>
rect 501 374 502 375 
<< pdiffusion >>
rect 502 374 503 375 
<< pdiffusion >>
rect 503 374 504 375 
<< pdiffusion >>
rect 516 374 517 375 
<< pdiffusion >>
rect 517 374 518 375 
<< pdiffusion >>
rect 518 374 519 375 
<< pdiffusion >>
rect 519 374 520 375 
<< pdiffusion >>
rect 520 374 521 375 
<< pdiffusion >>
rect 521 374 522 375 
<< m1 >>
rect 523 374 524 375 
<< pdiffusion >>
rect 12 375 13 376 
<< pdiffusion >>
rect 13 375 14 376 
<< pdiffusion >>
rect 14 375 15 376 
<< pdiffusion >>
rect 15 375 16 376 
<< pdiffusion >>
rect 16 375 17 376 
<< pdiffusion >>
rect 17 375 18 376 
<< m1 >>
rect 19 375 20 376 
<< m1 >>
rect 23 375 24 376 
<< pdiffusion >>
rect 30 375 31 376 
<< pdiffusion >>
rect 31 375 32 376 
<< pdiffusion >>
rect 32 375 33 376 
<< pdiffusion >>
rect 33 375 34 376 
<< pdiffusion >>
rect 34 375 35 376 
<< pdiffusion >>
rect 35 375 36 376 
<< m1 >>
rect 44 375 45 376 
<< pdiffusion >>
rect 48 375 49 376 
<< pdiffusion >>
rect 49 375 50 376 
<< pdiffusion >>
rect 50 375 51 376 
<< pdiffusion >>
rect 51 375 52 376 
<< pdiffusion >>
rect 52 375 53 376 
<< pdiffusion >>
rect 53 375 54 376 
<< m1 >>
rect 62 375 63 376 
<< pdiffusion >>
rect 66 375 67 376 
<< pdiffusion >>
rect 67 375 68 376 
<< pdiffusion >>
rect 68 375 69 376 
<< pdiffusion >>
rect 69 375 70 376 
<< pdiffusion >>
rect 70 375 71 376 
<< pdiffusion >>
rect 71 375 72 376 
<< m1 >>
rect 76 375 77 376 
<< m1 >>
rect 78 375 79 376 
<< m1 >>
rect 82 375 83 376 
<< pdiffusion >>
rect 84 375 85 376 
<< pdiffusion >>
rect 85 375 86 376 
<< pdiffusion >>
rect 86 375 87 376 
<< pdiffusion >>
rect 87 375 88 376 
<< pdiffusion >>
rect 88 375 89 376 
<< pdiffusion >>
rect 89 375 90 376 
<< m1 >>
rect 91 375 92 376 
<< m1 >>
rect 93 375 94 376 
<< m1 >>
rect 100 375 101 376 
<< pdiffusion >>
rect 102 375 103 376 
<< pdiffusion >>
rect 103 375 104 376 
<< pdiffusion >>
rect 104 375 105 376 
<< pdiffusion >>
rect 105 375 106 376 
<< pdiffusion >>
rect 106 375 107 376 
<< pdiffusion >>
rect 107 375 108 376 
<< m1 >>
rect 110 375 111 376 
<< m1 >>
rect 112 375 113 376 
<< pdiffusion >>
rect 120 375 121 376 
<< pdiffusion >>
rect 121 375 122 376 
<< pdiffusion >>
rect 122 375 123 376 
<< pdiffusion >>
rect 123 375 124 376 
<< pdiffusion >>
rect 124 375 125 376 
<< pdiffusion >>
rect 125 375 126 376 
<< m1 >>
rect 127 375 128 376 
<< m1 >>
rect 129 375 130 376 
<< pdiffusion >>
rect 138 375 139 376 
<< pdiffusion >>
rect 139 375 140 376 
<< pdiffusion >>
rect 140 375 141 376 
<< pdiffusion >>
rect 141 375 142 376 
<< pdiffusion >>
rect 142 375 143 376 
<< pdiffusion >>
rect 143 375 144 376 
<< m1 >>
rect 148 375 149 376 
<< m1 >>
rect 150 375 151 376 
<< pdiffusion >>
rect 156 375 157 376 
<< pdiffusion >>
rect 157 375 158 376 
<< pdiffusion >>
rect 158 375 159 376 
<< pdiffusion >>
rect 159 375 160 376 
<< pdiffusion >>
rect 160 375 161 376 
<< pdiffusion >>
rect 161 375 162 376 
<< m1 >>
rect 163 375 164 376 
<< m2 >>
rect 163 375 164 376 
<< m1 >>
rect 169 375 170 376 
<< m1 >>
rect 172 375 173 376 
<< pdiffusion >>
rect 174 375 175 376 
<< pdiffusion >>
rect 175 375 176 376 
<< pdiffusion >>
rect 176 375 177 376 
<< pdiffusion >>
rect 177 375 178 376 
<< pdiffusion >>
rect 178 375 179 376 
<< pdiffusion >>
rect 179 375 180 376 
<< m1 >>
rect 190 375 191 376 
<< pdiffusion >>
rect 192 375 193 376 
<< pdiffusion >>
rect 193 375 194 376 
<< pdiffusion >>
rect 194 375 195 376 
<< pdiffusion >>
rect 195 375 196 376 
<< pdiffusion >>
rect 196 375 197 376 
<< pdiffusion >>
rect 197 375 198 376 
<< m1 >>
rect 200 375 201 376 
<< m1 >>
rect 204 375 205 376 
<< m1 >>
rect 208 375 209 376 
<< pdiffusion >>
rect 210 375 211 376 
<< pdiffusion >>
rect 211 375 212 376 
<< pdiffusion >>
rect 212 375 213 376 
<< pdiffusion >>
rect 213 375 214 376 
<< pdiffusion >>
rect 214 375 215 376 
<< pdiffusion >>
rect 215 375 216 376 
<< m1 >>
rect 217 375 218 376 
<< m1 >>
rect 221 375 222 376 
<< m1 >>
rect 223 375 224 376 
<< pdiffusion >>
rect 228 375 229 376 
<< pdiffusion >>
rect 229 375 230 376 
<< pdiffusion >>
rect 230 375 231 376 
<< pdiffusion >>
rect 231 375 232 376 
<< pdiffusion >>
rect 232 375 233 376 
<< pdiffusion >>
rect 233 375 234 376 
<< m1 >>
rect 235 375 236 376 
<< m2 >>
rect 235 375 236 376 
<< m1 >>
rect 244 375 245 376 
<< pdiffusion >>
rect 246 375 247 376 
<< pdiffusion >>
rect 247 375 248 376 
<< pdiffusion >>
rect 248 375 249 376 
<< pdiffusion >>
rect 249 375 250 376 
<< pdiffusion >>
rect 250 375 251 376 
<< pdiffusion >>
rect 251 375 252 376 
<< m1 >>
rect 253 375 254 376 
<< m1 >>
rect 255 375 256 376 
<< pdiffusion >>
rect 264 375 265 376 
<< pdiffusion >>
rect 265 375 266 376 
<< pdiffusion >>
rect 266 375 267 376 
<< pdiffusion >>
rect 267 375 268 376 
<< pdiffusion >>
rect 268 375 269 376 
<< pdiffusion >>
rect 269 375 270 376 
<< m1 >>
rect 271 375 272 376 
<< pdiffusion >>
rect 282 375 283 376 
<< pdiffusion >>
rect 283 375 284 376 
<< pdiffusion >>
rect 284 375 285 376 
<< pdiffusion >>
rect 285 375 286 376 
<< pdiffusion >>
rect 286 375 287 376 
<< pdiffusion >>
rect 287 375 288 376 
<< pdiffusion >>
rect 300 375 301 376 
<< pdiffusion >>
rect 301 375 302 376 
<< pdiffusion >>
rect 302 375 303 376 
<< pdiffusion >>
rect 303 375 304 376 
<< pdiffusion >>
rect 304 375 305 376 
<< pdiffusion >>
rect 305 375 306 376 
<< m1 >>
rect 307 375 308 376 
<< m1 >>
rect 316 375 317 376 
<< pdiffusion >>
rect 318 375 319 376 
<< pdiffusion >>
rect 319 375 320 376 
<< pdiffusion >>
rect 320 375 321 376 
<< pdiffusion >>
rect 321 375 322 376 
<< pdiffusion >>
rect 322 375 323 376 
<< pdiffusion >>
rect 323 375 324 376 
<< m1 >>
rect 325 375 326 376 
<< m1 >>
rect 334 375 335 376 
<< pdiffusion >>
rect 336 375 337 376 
<< pdiffusion >>
rect 337 375 338 376 
<< pdiffusion >>
rect 338 375 339 376 
<< pdiffusion >>
rect 339 375 340 376 
<< pdiffusion >>
rect 340 375 341 376 
<< pdiffusion >>
rect 341 375 342 376 
<< m1 >>
rect 343 375 344 376 
<< pdiffusion >>
rect 354 375 355 376 
<< pdiffusion >>
rect 355 375 356 376 
<< pdiffusion >>
rect 356 375 357 376 
<< pdiffusion >>
rect 357 375 358 376 
<< pdiffusion >>
rect 358 375 359 376 
<< pdiffusion >>
rect 359 375 360 376 
<< m1 >>
rect 365 375 366 376 
<< pdiffusion >>
rect 372 375 373 376 
<< pdiffusion >>
rect 373 375 374 376 
<< pdiffusion >>
rect 374 375 375 376 
<< pdiffusion >>
rect 375 375 376 376 
<< pdiffusion >>
rect 376 375 377 376 
<< pdiffusion >>
rect 377 375 378 376 
<< pdiffusion >>
rect 390 375 391 376 
<< pdiffusion >>
rect 391 375 392 376 
<< pdiffusion >>
rect 392 375 393 376 
<< pdiffusion >>
rect 393 375 394 376 
<< pdiffusion >>
rect 394 375 395 376 
<< pdiffusion >>
rect 395 375 396 376 
<< m1 >>
rect 397 375 398 376 
<< m1 >>
rect 402 375 403 376 
<< m1 >>
rect 405 375 406 376 
<< pdiffusion >>
rect 408 375 409 376 
<< pdiffusion >>
rect 409 375 410 376 
<< pdiffusion >>
rect 410 375 411 376 
<< pdiffusion >>
rect 411 375 412 376 
<< pdiffusion >>
rect 412 375 413 376 
<< pdiffusion >>
rect 413 375 414 376 
<< m1 >>
rect 416 375 417 376 
<< pdiffusion >>
rect 426 375 427 376 
<< pdiffusion >>
rect 427 375 428 376 
<< pdiffusion >>
rect 428 375 429 376 
<< pdiffusion >>
rect 429 375 430 376 
<< pdiffusion >>
rect 430 375 431 376 
<< pdiffusion >>
rect 431 375 432 376 
<< m1 >>
rect 433 375 434 376 
<< m1 >>
rect 435 375 436 376 
<< pdiffusion >>
rect 444 375 445 376 
<< pdiffusion >>
rect 445 375 446 376 
<< pdiffusion >>
rect 446 375 447 376 
<< pdiffusion >>
rect 447 375 448 376 
<< pdiffusion >>
rect 448 375 449 376 
<< pdiffusion >>
rect 449 375 450 376 
<< m1 >>
rect 451 375 452 376 
<< m1 >>
rect 453 375 454 376 
<< m1 >>
rect 455 375 456 376 
<< m1 >>
rect 457 375 458 376 
<< pdiffusion >>
rect 462 375 463 376 
<< pdiffusion >>
rect 463 375 464 376 
<< pdiffusion >>
rect 464 375 465 376 
<< pdiffusion >>
rect 465 375 466 376 
<< pdiffusion >>
rect 466 375 467 376 
<< pdiffusion >>
rect 467 375 468 376 
<< pdiffusion >>
rect 498 375 499 376 
<< pdiffusion >>
rect 499 375 500 376 
<< pdiffusion >>
rect 500 375 501 376 
<< pdiffusion >>
rect 501 375 502 376 
<< pdiffusion >>
rect 502 375 503 376 
<< pdiffusion >>
rect 503 375 504 376 
<< pdiffusion >>
rect 516 375 517 376 
<< pdiffusion >>
rect 517 375 518 376 
<< pdiffusion >>
rect 518 375 519 376 
<< pdiffusion >>
rect 519 375 520 376 
<< pdiffusion >>
rect 520 375 521 376 
<< pdiffusion >>
rect 521 375 522 376 
<< m1 >>
rect 523 375 524 376 
<< pdiffusion >>
rect 12 376 13 377 
<< pdiffusion >>
rect 13 376 14 377 
<< pdiffusion >>
rect 14 376 15 377 
<< pdiffusion >>
rect 15 376 16 377 
<< pdiffusion >>
rect 16 376 17 377 
<< pdiffusion >>
rect 17 376 18 377 
<< m1 >>
rect 19 376 20 377 
<< m1 >>
rect 23 376 24 377 
<< pdiffusion >>
rect 30 376 31 377 
<< pdiffusion >>
rect 31 376 32 377 
<< pdiffusion >>
rect 32 376 33 377 
<< pdiffusion >>
rect 33 376 34 377 
<< pdiffusion >>
rect 34 376 35 377 
<< pdiffusion >>
rect 35 376 36 377 
<< m1 >>
rect 44 376 45 377 
<< pdiffusion >>
rect 48 376 49 377 
<< pdiffusion >>
rect 49 376 50 377 
<< pdiffusion >>
rect 50 376 51 377 
<< pdiffusion >>
rect 51 376 52 377 
<< pdiffusion >>
rect 52 376 53 377 
<< pdiffusion >>
rect 53 376 54 377 
<< m1 >>
rect 62 376 63 377 
<< pdiffusion >>
rect 66 376 67 377 
<< pdiffusion >>
rect 67 376 68 377 
<< pdiffusion >>
rect 68 376 69 377 
<< pdiffusion >>
rect 69 376 70 377 
<< pdiffusion >>
rect 70 376 71 377 
<< pdiffusion >>
rect 71 376 72 377 
<< m1 >>
rect 76 376 77 377 
<< m1 >>
rect 78 376 79 377 
<< m1 >>
rect 82 376 83 377 
<< pdiffusion >>
rect 84 376 85 377 
<< pdiffusion >>
rect 85 376 86 377 
<< pdiffusion >>
rect 86 376 87 377 
<< pdiffusion >>
rect 87 376 88 377 
<< pdiffusion >>
rect 88 376 89 377 
<< pdiffusion >>
rect 89 376 90 377 
<< m1 >>
rect 91 376 92 377 
<< m1 >>
rect 93 376 94 377 
<< m1 >>
rect 100 376 101 377 
<< pdiffusion >>
rect 102 376 103 377 
<< pdiffusion >>
rect 103 376 104 377 
<< pdiffusion >>
rect 104 376 105 377 
<< pdiffusion >>
rect 105 376 106 377 
<< pdiffusion >>
rect 106 376 107 377 
<< pdiffusion >>
rect 107 376 108 377 
<< m1 >>
rect 110 376 111 377 
<< m1 >>
rect 112 376 113 377 
<< pdiffusion >>
rect 120 376 121 377 
<< pdiffusion >>
rect 121 376 122 377 
<< pdiffusion >>
rect 122 376 123 377 
<< pdiffusion >>
rect 123 376 124 377 
<< pdiffusion >>
rect 124 376 125 377 
<< pdiffusion >>
rect 125 376 126 377 
<< m1 >>
rect 127 376 128 377 
<< m1 >>
rect 129 376 130 377 
<< pdiffusion >>
rect 138 376 139 377 
<< pdiffusion >>
rect 139 376 140 377 
<< pdiffusion >>
rect 140 376 141 377 
<< pdiffusion >>
rect 141 376 142 377 
<< pdiffusion >>
rect 142 376 143 377 
<< pdiffusion >>
rect 143 376 144 377 
<< m1 >>
rect 148 376 149 377 
<< m1 >>
rect 150 376 151 377 
<< pdiffusion >>
rect 156 376 157 377 
<< pdiffusion >>
rect 157 376 158 377 
<< pdiffusion >>
rect 158 376 159 377 
<< pdiffusion >>
rect 159 376 160 377 
<< pdiffusion >>
rect 160 376 161 377 
<< pdiffusion >>
rect 161 376 162 377 
<< m1 >>
rect 163 376 164 377 
<< m2 >>
rect 163 376 164 377 
<< m1 >>
rect 169 376 170 377 
<< m1 >>
rect 172 376 173 377 
<< pdiffusion >>
rect 174 376 175 377 
<< pdiffusion >>
rect 175 376 176 377 
<< pdiffusion >>
rect 176 376 177 377 
<< pdiffusion >>
rect 177 376 178 377 
<< pdiffusion >>
rect 178 376 179 377 
<< pdiffusion >>
rect 179 376 180 377 
<< m1 >>
rect 190 376 191 377 
<< pdiffusion >>
rect 192 376 193 377 
<< pdiffusion >>
rect 193 376 194 377 
<< pdiffusion >>
rect 194 376 195 377 
<< pdiffusion >>
rect 195 376 196 377 
<< pdiffusion >>
rect 196 376 197 377 
<< pdiffusion >>
rect 197 376 198 377 
<< m1 >>
rect 200 376 201 377 
<< m1 >>
rect 204 376 205 377 
<< m1 >>
rect 208 376 209 377 
<< pdiffusion >>
rect 210 376 211 377 
<< pdiffusion >>
rect 211 376 212 377 
<< pdiffusion >>
rect 212 376 213 377 
<< pdiffusion >>
rect 213 376 214 377 
<< pdiffusion >>
rect 214 376 215 377 
<< pdiffusion >>
rect 215 376 216 377 
<< m1 >>
rect 217 376 218 377 
<< m1 >>
rect 221 376 222 377 
<< m1 >>
rect 223 376 224 377 
<< pdiffusion >>
rect 228 376 229 377 
<< pdiffusion >>
rect 229 376 230 377 
<< pdiffusion >>
rect 230 376 231 377 
<< pdiffusion >>
rect 231 376 232 377 
<< pdiffusion >>
rect 232 376 233 377 
<< pdiffusion >>
rect 233 376 234 377 
<< m1 >>
rect 235 376 236 377 
<< m2 >>
rect 235 376 236 377 
<< m1 >>
rect 244 376 245 377 
<< pdiffusion >>
rect 246 376 247 377 
<< pdiffusion >>
rect 247 376 248 377 
<< pdiffusion >>
rect 248 376 249 377 
<< pdiffusion >>
rect 249 376 250 377 
<< pdiffusion >>
rect 250 376 251 377 
<< pdiffusion >>
rect 251 376 252 377 
<< m1 >>
rect 253 376 254 377 
<< m1 >>
rect 255 376 256 377 
<< pdiffusion >>
rect 264 376 265 377 
<< pdiffusion >>
rect 265 376 266 377 
<< pdiffusion >>
rect 266 376 267 377 
<< pdiffusion >>
rect 267 376 268 377 
<< pdiffusion >>
rect 268 376 269 377 
<< pdiffusion >>
rect 269 376 270 377 
<< m1 >>
rect 271 376 272 377 
<< pdiffusion >>
rect 282 376 283 377 
<< pdiffusion >>
rect 283 376 284 377 
<< pdiffusion >>
rect 284 376 285 377 
<< pdiffusion >>
rect 285 376 286 377 
<< pdiffusion >>
rect 286 376 287 377 
<< pdiffusion >>
rect 287 376 288 377 
<< pdiffusion >>
rect 300 376 301 377 
<< pdiffusion >>
rect 301 376 302 377 
<< pdiffusion >>
rect 302 376 303 377 
<< pdiffusion >>
rect 303 376 304 377 
<< pdiffusion >>
rect 304 376 305 377 
<< pdiffusion >>
rect 305 376 306 377 
<< m1 >>
rect 307 376 308 377 
<< m1 >>
rect 316 376 317 377 
<< pdiffusion >>
rect 318 376 319 377 
<< pdiffusion >>
rect 319 376 320 377 
<< pdiffusion >>
rect 320 376 321 377 
<< pdiffusion >>
rect 321 376 322 377 
<< pdiffusion >>
rect 322 376 323 377 
<< pdiffusion >>
rect 323 376 324 377 
<< m1 >>
rect 325 376 326 377 
<< m1 >>
rect 334 376 335 377 
<< pdiffusion >>
rect 336 376 337 377 
<< pdiffusion >>
rect 337 376 338 377 
<< pdiffusion >>
rect 338 376 339 377 
<< pdiffusion >>
rect 339 376 340 377 
<< pdiffusion >>
rect 340 376 341 377 
<< pdiffusion >>
rect 341 376 342 377 
<< m1 >>
rect 343 376 344 377 
<< pdiffusion >>
rect 354 376 355 377 
<< pdiffusion >>
rect 355 376 356 377 
<< pdiffusion >>
rect 356 376 357 377 
<< pdiffusion >>
rect 357 376 358 377 
<< pdiffusion >>
rect 358 376 359 377 
<< pdiffusion >>
rect 359 376 360 377 
<< m1 >>
rect 365 376 366 377 
<< pdiffusion >>
rect 372 376 373 377 
<< pdiffusion >>
rect 373 376 374 377 
<< pdiffusion >>
rect 374 376 375 377 
<< pdiffusion >>
rect 375 376 376 377 
<< pdiffusion >>
rect 376 376 377 377 
<< pdiffusion >>
rect 377 376 378 377 
<< pdiffusion >>
rect 390 376 391 377 
<< pdiffusion >>
rect 391 376 392 377 
<< pdiffusion >>
rect 392 376 393 377 
<< pdiffusion >>
rect 393 376 394 377 
<< pdiffusion >>
rect 394 376 395 377 
<< pdiffusion >>
rect 395 376 396 377 
<< m1 >>
rect 397 376 398 377 
<< m1 >>
rect 402 376 403 377 
<< m1 >>
rect 405 376 406 377 
<< pdiffusion >>
rect 408 376 409 377 
<< pdiffusion >>
rect 409 376 410 377 
<< pdiffusion >>
rect 410 376 411 377 
<< pdiffusion >>
rect 411 376 412 377 
<< pdiffusion >>
rect 412 376 413 377 
<< pdiffusion >>
rect 413 376 414 377 
<< m1 >>
rect 416 376 417 377 
<< pdiffusion >>
rect 426 376 427 377 
<< pdiffusion >>
rect 427 376 428 377 
<< pdiffusion >>
rect 428 376 429 377 
<< pdiffusion >>
rect 429 376 430 377 
<< pdiffusion >>
rect 430 376 431 377 
<< pdiffusion >>
rect 431 376 432 377 
<< m1 >>
rect 433 376 434 377 
<< m1 >>
rect 435 376 436 377 
<< pdiffusion >>
rect 444 376 445 377 
<< pdiffusion >>
rect 445 376 446 377 
<< pdiffusion >>
rect 446 376 447 377 
<< pdiffusion >>
rect 447 376 448 377 
<< pdiffusion >>
rect 448 376 449 377 
<< pdiffusion >>
rect 449 376 450 377 
<< m1 >>
rect 451 376 452 377 
<< m1 >>
rect 453 376 454 377 
<< m1 >>
rect 455 376 456 377 
<< m1 >>
rect 457 376 458 377 
<< pdiffusion >>
rect 462 376 463 377 
<< pdiffusion >>
rect 463 376 464 377 
<< pdiffusion >>
rect 464 376 465 377 
<< pdiffusion >>
rect 465 376 466 377 
<< pdiffusion >>
rect 466 376 467 377 
<< pdiffusion >>
rect 467 376 468 377 
<< pdiffusion >>
rect 498 376 499 377 
<< pdiffusion >>
rect 499 376 500 377 
<< pdiffusion >>
rect 500 376 501 377 
<< pdiffusion >>
rect 501 376 502 377 
<< pdiffusion >>
rect 502 376 503 377 
<< pdiffusion >>
rect 503 376 504 377 
<< pdiffusion >>
rect 516 376 517 377 
<< pdiffusion >>
rect 517 376 518 377 
<< pdiffusion >>
rect 518 376 519 377 
<< pdiffusion >>
rect 519 376 520 377 
<< pdiffusion >>
rect 520 376 521 377 
<< pdiffusion >>
rect 521 376 522 377 
<< m1 >>
rect 523 376 524 377 
<< pdiffusion >>
rect 12 377 13 378 
<< pdiffusion >>
rect 13 377 14 378 
<< pdiffusion >>
rect 14 377 15 378 
<< pdiffusion >>
rect 15 377 16 378 
<< m1 >>
rect 16 377 17 378 
<< pdiffusion >>
rect 16 377 17 378 
<< pdiffusion >>
rect 17 377 18 378 
<< m1 >>
rect 19 377 20 378 
<< m1 >>
rect 23 377 24 378 
<< pdiffusion >>
rect 30 377 31 378 
<< pdiffusion >>
rect 31 377 32 378 
<< pdiffusion >>
rect 32 377 33 378 
<< pdiffusion >>
rect 33 377 34 378 
<< pdiffusion >>
rect 34 377 35 378 
<< pdiffusion >>
rect 35 377 36 378 
<< m1 >>
rect 44 377 45 378 
<< pdiffusion >>
rect 48 377 49 378 
<< pdiffusion >>
rect 49 377 50 378 
<< pdiffusion >>
rect 50 377 51 378 
<< pdiffusion >>
rect 51 377 52 378 
<< pdiffusion >>
rect 52 377 53 378 
<< pdiffusion >>
rect 53 377 54 378 
<< m1 >>
rect 62 377 63 378 
<< pdiffusion >>
rect 66 377 67 378 
<< m1 >>
rect 67 377 68 378 
<< pdiffusion >>
rect 67 377 68 378 
<< pdiffusion >>
rect 68 377 69 378 
<< pdiffusion >>
rect 69 377 70 378 
<< pdiffusion >>
rect 70 377 71 378 
<< pdiffusion >>
rect 71 377 72 378 
<< m1 >>
rect 76 377 77 378 
<< m1 >>
rect 78 377 79 378 
<< m1 >>
rect 82 377 83 378 
<< pdiffusion >>
rect 84 377 85 378 
<< pdiffusion >>
rect 85 377 86 378 
<< pdiffusion >>
rect 86 377 87 378 
<< pdiffusion >>
rect 87 377 88 378 
<< m1 >>
rect 88 377 89 378 
<< pdiffusion >>
rect 88 377 89 378 
<< pdiffusion >>
rect 89 377 90 378 
<< m1 >>
rect 91 377 92 378 
<< m1 >>
rect 93 377 94 378 
<< m1 >>
rect 100 377 101 378 
<< m2 >>
rect 100 377 101 378 
<< m2c >>
rect 100 377 101 378 
<< m1 >>
rect 100 377 101 378 
<< m2 >>
rect 100 377 101 378 
<< pdiffusion >>
rect 102 377 103 378 
<< m1 >>
rect 103 377 104 378 
<< pdiffusion >>
rect 103 377 104 378 
<< pdiffusion >>
rect 104 377 105 378 
<< pdiffusion >>
rect 105 377 106 378 
<< pdiffusion >>
rect 106 377 107 378 
<< pdiffusion >>
rect 107 377 108 378 
<< m1 >>
rect 110 377 111 378 
<< m1 >>
rect 112 377 113 378 
<< pdiffusion >>
rect 120 377 121 378 
<< m1 >>
rect 121 377 122 378 
<< pdiffusion >>
rect 121 377 122 378 
<< pdiffusion >>
rect 122 377 123 378 
<< m1 >>
rect 123 377 124 378 
<< m2 >>
rect 123 377 124 378 
<< m2c >>
rect 123 377 124 378 
<< m1 >>
rect 123 377 124 378 
<< m2 >>
rect 123 377 124 378 
<< pdiffusion >>
rect 123 377 124 378 
<< m1 >>
rect 124 377 125 378 
<< pdiffusion >>
rect 124 377 125 378 
<< pdiffusion >>
rect 125 377 126 378 
<< m1 >>
rect 127 377 128 378 
<< m1 >>
rect 129 377 130 378 
<< pdiffusion >>
rect 138 377 139 378 
<< m1 >>
rect 139 377 140 378 
<< pdiffusion >>
rect 139 377 140 378 
<< pdiffusion >>
rect 140 377 141 378 
<< pdiffusion >>
rect 141 377 142 378 
<< pdiffusion >>
rect 142 377 143 378 
<< pdiffusion >>
rect 143 377 144 378 
<< m1 >>
rect 148 377 149 378 
<< m1 >>
rect 150 377 151 378 
<< pdiffusion >>
rect 156 377 157 378 
<< m1 >>
rect 157 377 158 378 
<< pdiffusion >>
rect 157 377 158 378 
<< pdiffusion >>
rect 158 377 159 378 
<< pdiffusion >>
rect 159 377 160 378 
<< pdiffusion >>
rect 160 377 161 378 
<< pdiffusion >>
rect 161 377 162 378 
<< m1 >>
rect 163 377 164 378 
<< m2 >>
rect 163 377 164 378 
<< m1 >>
rect 169 377 170 378 
<< m1 >>
rect 172 377 173 378 
<< pdiffusion >>
rect 174 377 175 378 
<< pdiffusion >>
rect 175 377 176 378 
<< pdiffusion >>
rect 176 377 177 378 
<< pdiffusion >>
rect 177 377 178 378 
<< pdiffusion >>
rect 178 377 179 378 
<< pdiffusion >>
rect 179 377 180 378 
<< m1 >>
rect 190 377 191 378 
<< pdiffusion >>
rect 192 377 193 378 
<< m1 >>
rect 193 377 194 378 
<< pdiffusion >>
rect 193 377 194 378 
<< pdiffusion >>
rect 194 377 195 378 
<< pdiffusion >>
rect 195 377 196 378 
<< pdiffusion >>
rect 196 377 197 378 
<< pdiffusion >>
rect 197 377 198 378 
<< m1 >>
rect 200 377 201 378 
<< m1 >>
rect 204 377 205 378 
<< m1 >>
rect 208 377 209 378 
<< pdiffusion >>
rect 210 377 211 378 
<< pdiffusion >>
rect 211 377 212 378 
<< pdiffusion >>
rect 212 377 213 378 
<< pdiffusion >>
rect 213 377 214 378 
<< pdiffusion >>
rect 214 377 215 378 
<< pdiffusion >>
rect 215 377 216 378 
<< m1 >>
rect 217 377 218 378 
<< m1 >>
rect 221 377 222 378 
<< m1 >>
rect 223 377 224 378 
<< pdiffusion >>
rect 228 377 229 378 
<< pdiffusion >>
rect 229 377 230 378 
<< pdiffusion >>
rect 230 377 231 378 
<< pdiffusion >>
rect 231 377 232 378 
<< m1 >>
rect 232 377 233 378 
<< pdiffusion >>
rect 232 377 233 378 
<< pdiffusion >>
rect 233 377 234 378 
<< m1 >>
rect 235 377 236 378 
<< m2 >>
rect 235 377 236 378 
<< m1 >>
rect 244 377 245 378 
<< pdiffusion >>
rect 246 377 247 378 
<< pdiffusion >>
rect 247 377 248 378 
<< pdiffusion >>
rect 248 377 249 378 
<< pdiffusion >>
rect 249 377 250 378 
<< pdiffusion >>
rect 250 377 251 378 
<< pdiffusion >>
rect 251 377 252 378 
<< m1 >>
rect 253 377 254 378 
<< m1 >>
rect 255 377 256 378 
<< pdiffusion >>
rect 264 377 265 378 
<< m1 >>
rect 265 377 266 378 
<< pdiffusion >>
rect 265 377 266 378 
<< pdiffusion >>
rect 266 377 267 378 
<< pdiffusion >>
rect 267 377 268 378 
<< pdiffusion >>
rect 268 377 269 378 
<< pdiffusion >>
rect 269 377 270 378 
<< m1 >>
rect 271 377 272 378 
<< pdiffusion >>
rect 282 377 283 378 
<< pdiffusion >>
rect 283 377 284 378 
<< pdiffusion >>
rect 284 377 285 378 
<< pdiffusion >>
rect 285 377 286 378 
<< pdiffusion >>
rect 286 377 287 378 
<< pdiffusion >>
rect 287 377 288 378 
<< pdiffusion >>
rect 300 377 301 378 
<< pdiffusion >>
rect 301 377 302 378 
<< pdiffusion >>
rect 302 377 303 378 
<< pdiffusion >>
rect 303 377 304 378 
<< pdiffusion >>
rect 304 377 305 378 
<< pdiffusion >>
rect 305 377 306 378 
<< m1 >>
rect 307 377 308 378 
<< m1 >>
rect 316 377 317 378 
<< pdiffusion >>
rect 318 377 319 378 
<< pdiffusion >>
rect 319 377 320 378 
<< pdiffusion >>
rect 320 377 321 378 
<< pdiffusion >>
rect 321 377 322 378 
<< pdiffusion >>
rect 322 377 323 378 
<< pdiffusion >>
rect 323 377 324 378 
<< m1 >>
rect 325 377 326 378 
<< m1 >>
rect 334 377 335 378 
<< pdiffusion >>
rect 336 377 337 378 
<< pdiffusion >>
rect 337 377 338 378 
<< pdiffusion >>
rect 338 377 339 378 
<< pdiffusion >>
rect 339 377 340 378 
<< pdiffusion >>
rect 340 377 341 378 
<< pdiffusion >>
rect 341 377 342 378 
<< m1 >>
rect 343 377 344 378 
<< pdiffusion >>
rect 354 377 355 378 
<< m1 >>
rect 355 377 356 378 
<< pdiffusion >>
rect 355 377 356 378 
<< pdiffusion >>
rect 356 377 357 378 
<< pdiffusion >>
rect 357 377 358 378 
<< pdiffusion >>
rect 358 377 359 378 
<< pdiffusion >>
rect 359 377 360 378 
<< m1 >>
rect 365 377 366 378 
<< pdiffusion >>
rect 372 377 373 378 
<< pdiffusion >>
rect 373 377 374 378 
<< pdiffusion >>
rect 374 377 375 378 
<< pdiffusion >>
rect 375 377 376 378 
<< m1 >>
rect 376 377 377 378 
<< pdiffusion >>
rect 376 377 377 378 
<< pdiffusion >>
rect 377 377 378 378 
<< pdiffusion >>
rect 390 377 391 378 
<< pdiffusion >>
rect 391 377 392 378 
<< pdiffusion >>
rect 392 377 393 378 
<< pdiffusion >>
rect 393 377 394 378 
<< m1 >>
rect 394 377 395 378 
<< pdiffusion >>
rect 394 377 395 378 
<< pdiffusion >>
rect 395 377 396 378 
<< m1 >>
rect 397 377 398 378 
<< m1 >>
rect 402 377 403 378 
<< m1 >>
rect 405 377 406 378 
<< pdiffusion >>
rect 408 377 409 378 
<< pdiffusion >>
rect 409 377 410 378 
<< pdiffusion >>
rect 410 377 411 378 
<< pdiffusion >>
rect 411 377 412 378 
<< pdiffusion >>
rect 412 377 413 378 
<< pdiffusion >>
rect 413 377 414 378 
<< m1 >>
rect 416 377 417 378 
<< pdiffusion >>
rect 426 377 427 378 
<< pdiffusion >>
rect 427 377 428 378 
<< pdiffusion >>
rect 428 377 429 378 
<< pdiffusion >>
rect 429 377 430 378 
<< m1 >>
rect 430 377 431 378 
<< pdiffusion >>
rect 430 377 431 378 
<< pdiffusion >>
rect 431 377 432 378 
<< m1 >>
rect 433 377 434 378 
<< m1 >>
rect 435 377 436 378 
<< pdiffusion >>
rect 444 377 445 378 
<< pdiffusion >>
rect 445 377 446 378 
<< pdiffusion >>
rect 446 377 447 378 
<< pdiffusion >>
rect 447 377 448 378 
<< pdiffusion >>
rect 448 377 449 378 
<< pdiffusion >>
rect 449 377 450 378 
<< m1 >>
rect 451 377 452 378 
<< m1 >>
rect 453 377 454 378 
<< m1 >>
rect 455 377 456 378 
<< m1 >>
rect 457 377 458 378 
<< pdiffusion >>
rect 462 377 463 378 
<< pdiffusion >>
rect 463 377 464 378 
<< pdiffusion >>
rect 464 377 465 378 
<< pdiffusion >>
rect 465 377 466 378 
<< pdiffusion >>
rect 466 377 467 378 
<< pdiffusion >>
rect 467 377 468 378 
<< pdiffusion >>
rect 498 377 499 378 
<< pdiffusion >>
rect 499 377 500 378 
<< pdiffusion >>
rect 500 377 501 378 
<< pdiffusion >>
rect 501 377 502 378 
<< pdiffusion >>
rect 502 377 503 378 
<< pdiffusion >>
rect 503 377 504 378 
<< pdiffusion >>
rect 516 377 517 378 
<< pdiffusion >>
rect 517 377 518 378 
<< pdiffusion >>
rect 518 377 519 378 
<< pdiffusion >>
rect 519 377 520 378 
<< m1 >>
rect 520 377 521 378 
<< pdiffusion >>
rect 520 377 521 378 
<< pdiffusion >>
rect 521 377 522 378 
<< m1 >>
rect 523 377 524 378 
<< m1 >>
rect 16 378 17 379 
<< m1 >>
rect 19 378 20 379 
<< m1 >>
rect 23 378 24 379 
<< m1 >>
rect 44 378 45 379 
<< m1 >>
rect 60 378 61 379 
<< m2 >>
rect 60 378 61 379 
<< m2c >>
rect 60 378 61 379 
<< m1 >>
rect 60 378 61 379 
<< m2 >>
rect 60 378 61 379 
<< m2 >>
rect 61 378 62 379 
<< m1 >>
rect 62 378 63 379 
<< m2 >>
rect 62 378 63 379 
<< m2 >>
rect 63 378 64 379 
<< m1 >>
rect 64 378 65 379 
<< m2 >>
rect 64 378 65 379 
<< m2c >>
rect 64 378 65 379 
<< m1 >>
rect 64 378 65 379 
<< m2 >>
rect 64 378 65 379 
<< m1 >>
rect 67 378 68 379 
<< m1 >>
rect 76 378 77 379 
<< m1 >>
rect 78 378 79 379 
<< m1 >>
rect 82 378 83 379 
<< m1 >>
rect 88 378 89 379 
<< m1 >>
rect 91 378 92 379 
<< m1 >>
rect 93 378 94 379 
<< m2 >>
rect 100 378 101 379 
<< m1 >>
rect 103 378 104 379 
<< m1 >>
rect 110 378 111 379 
<< m1 >>
rect 112 378 113 379 
<< m1 >>
rect 121 378 122 379 
<< m1 >>
rect 124 378 125 379 
<< m2 >>
rect 124 378 125 379 
<< m1 >>
rect 127 378 128 379 
<< m1 >>
rect 129 378 130 379 
<< m1 >>
rect 139 378 140 379 
<< m1 >>
rect 148 378 149 379 
<< m1 >>
rect 150 378 151 379 
<< m1 >>
rect 157 378 158 379 
<< m1 >>
rect 163 378 164 379 
<< m2 >>
rect 163 378 164 379 
<< m1 >>
rect 169 378 170 379 
<< m1 >>
rect 172 378 173 379 
<< m1 >>
rect 190 378 191 379 
<< m1 >>
rect 193 378 194 379 
<< m1 >>
rect 200 378 201 379 
<< m1 >>
rect 204 378 205 379 
<< m1 >>
rect 208 378 209 379 
<< m1 >>
rect 217 378 218 379 
<< m1 >>
rect 221 378 222 379 
<< m1 >>
rect 223 378 224 379 
<< m1 >>
rect 232 378 233 379 
<< m1 >>
rect 235 378 236 379 
<< m2 >>
rect 235 378 236 379 
<< m1 >>
rect 244 378 245 379 
<< m1 >>
rect 253 378 254 379 
<< m1 >>
rect 255 378 256 379 
<< m1 >>
rect 265 378 266 379 
<< m1 >>
rect 271 378 272 379 
<< m1 >>
rect 307 378 308 379 
<< m1 >>
rect 316 378 317 379 
<< m1 >>
rect 325 378 326 379 
<< m1 >>
rect 334 378 335 379 
<< m1 >>
rect 343 378 344 379 
<< m1 >>
rect 355 378 356 379 
<< m1 >>
rect 365 378 366 379 
<< m1 >>
rect 376 378 377 379 
<< m1 >>
rect 394 378 395 379 
<< m1 >>
rect 397 378 398 379 
<< m1 >>
rect 402 378 403 379 
<< m1 >>
rect 405 378 406 379 
<< m1 >>
rect 416 378 417 379 
<< m1 >>
rect 430 378 431 379 
<< m1 >>
rect 433 378 434 379 
<< m1 >>
rect 435 378 436 379 
<< m1 >>
rect 451 378 452 379 
<< m1 >>
rect 453 378 454 379 
<< m1 >>
rect 455 378 456 379 
<< m1 >>
rect 457 378 458 379 
<< m1 >>
rect 520 378 521 379 
<< m1 >>
rect 523 378 524 379 
<< m1 >>
rect 16 379 17 380 
<< m1 >>
rect 19 379 20 380 
<< m1 >>
rect 23 379 24 380 
<< m1 >>
rect 44 379 45 380 
<< m1 >>
rect 60 379 61 380 
<< m1 >>
rect 62 379 63 380 
<< m1 >>
rect 64 379 65 380 
<< m1 >>
rect 65 379 66 380 
<< m1 >>
rect 66 379 67 380 
<< m1 >>
rect 67 379 68 380 
<< m1 >>
rect 76 379 77 380 
<< m1 >>
rect 78 379 79 380 
<< m1 >>
rect 82 379 83 380 
<< m1 >>
rect 88 379 89 380 
<< m1 >>
rect 89 379 90 380 
<< m2 >>
rect 89 379 90 380 
<< m2c >>
rect 89 379 90 380 
<< m1 >>
rect 89 379 90 380 
<< m2 >>
rect 89 379 90 380 
<< m2 >>
rect 90 379 91 380 
<< m1 >>
rect 91 379 92 380 
<< m2 >>
rect 91 379 92 380 
<< m2 >>
rect 92 379 93 380 
<< m1 >>
rect 93 379 94 380 
<< m2 >>
rect 93 379 94 380 
<< m2 >>
rect 94 379 95 380 
<< m1 >>
rect 95 379 96 380 
<< m2 >>
rect 95 379 96 380 
<< m2c >>
rect 95 379 96 380 
<< m1 >>
rect 95 379 96 380 
<< m2 >>
rect 95 379 96 380 
<< m1 >>
rect 96 379 97 380 
<< m1 >>
rect 97 379 98 380 
<< m1 >>
rect 98 379 99 380 
<< m1 >>
rect 99 379 100 380 
<< m1 >>
rect 100 379 101 380 
<< m2 >>
rect 100 379 101 380 
<< m1 >>
rect 101 379 102 380 
<< m1 >>
rect 102 379 103 380 
<< m1 >>
rect 103 379 104 380 
<< m1 >>
rect 110 379 111 380 
<< m1 >>
rect 112 379 113 380 
<< m1 >>
rect 121 379 122 380 
<< m2 >>
rect 124 379 125 380 
<< m2 >>
rect 125 379 126 380 
<< m2 >>
rect 126 379 127 380 
<< m1 >>
rect 127 379 128 380 
<< m2 >>
rect 127 379 128 380 
<< m2 >>
rect 128 379 129 380 
<< m1 >>
rect 129 379 130 380 
<< m2 >>
rect 129 379 130 380 
<< m2c >>
rect 129 379 130 380 
<< m1 >>
rect 129 379 130 380 
<< m2 >>
rect 129 379 130 380 
<< m1 >>
rect 139 379 140 380 
<< m1 >>
rect 148 379 149 380 
<< m1 >>
rect 150 379 151 380 
<< m2 >>
rect 151 379 152 380 
<< m1 >>
rect 152 379 153 380 
<< m2 >>
rect 152 379 153 380 
<< m2c >>
rect 152 379 153 380 
<< m1 >>
rect 152 379 153 380 
<< m2 >>
rect 152 379 153 380 
<< m1 >>
rect 153 379 154 380 
<< m1 >>
rect 154 379 155 380 
<< m1 >>
rect 155 379 156 380 
<< m1 >>
rect 156 379 157 380 
<< m1 >>
rect 157 379 158 380 
<< m1 >>
rect 163 379 164 380 
<< m2 >>
rect 163 379 164 380 
<< m1 >>
rect 169 379 170 380 
<< m1 >>
rect 172 379 173 380 
<< m1 >>
rect 190 379 191 380 
<< m1 >>
rect 193 379 194 380 
<< m1 >>
rect 200 379 201 380 
<< m1 >>
rect 204 379 205 380 
<< m1 >>
rect 208 379 209 380 
<< m1 >>
rect 217 379 218 380 
<< m1 >>
rect 221 379 222 380 
<< m1 >>
rect 223 379 224 380 
<< m1 >>
rect 232 379 233 380 
<< m1 >>
rect 233 379 234 380 
<< m2 >>
rect 233 379 234 380 
<< m2c >>
rect 233 379 234 380 
<< m1 >>
rect 233 379 234 380 
<< m2 >>
rect 233 379 234 380 
<< m2 >>
rect 234 379 235 380 
<< m1 >>
rect 235 379 236 380 
<< m2 >>
rect 235 379 236 380 
<< m1 >>
rect 244 379 245 380 
<< m1 >>
rect 253 379 254 380 
<< m1 >>
rect 255 379 256 380 
<< m1 >>
rect 265 379 266 380 
<< m1 >>
rect 271 379 272 380 
<< m1 >>
rect 307 379 308 380 
<< m1 >>
rect 316 379 317 380 
<< m1 >>
rect 325 379 326 380 
<< m1 >>
rect 334 379 335 380 
<< m1 >>
rect 343 379 344 380 
<< m1 >>
rect 355 379 356 380 
<< m1 >>
rect 365 379 366 380 
<< m1 >>
rect 376 379 377 380 
<< m1 >>
rect 394 379 395 380 
<< m1 >>
rect 397 379 398 380 
<< m1 >>
rect 402 379 403 380 
<< m1 >>
rect 405 379 406 380 
<< m1 >>
rect 416 379 417 380 
<< m1 >>
rect 429 379 430 380 
<< m1 >>
rect 430 379 431 380 
<< m1 >>
rect 433 379 434 380 
<< m1 >>
rect 435 379 436 380 
<< m1 >>
rect 451 379 452 380 
<< m1 >>
rect 453 379 454 380 
<< m1 >>
rect 455 379 456 380 
<< m1 >>
rect 457 379 458 380 
<< m1 >>
rect 520 379 521 380 
<< m1 >>
rect 523 379 524 380 
<< m1 >>
rect 16 380 17 381 
<< m1 >>
rect 19 380 20 381 
<< m1 >>
rect 23 380 24 381 
<< m1 >>
rect 44 380 45 381 
<< m2 >>
rect 44 380 45 381 
<< m2c >>
rect 44 380 45 381 
<< m1 >>
rect 44 380 45 381 
<< m2 >>
rect 44 380 45 381 
<< m1 >>
rect 60 380 61 381 
<< m2 >>
rect 60 380 61 381 
<< m2c >>
rect 60 380 61 381 
<< m1 >>
rect 60 380 61 381 
<< m2 >>
rect 60 380 61 381 
<< m1 >>
rect 62 380 63 381 
<< m2 >>
rect 62 380 63 381 
<< m2c >>
rect 62 380 63 381 
<< m1 >>
rect 62 380 63 381 
<< m2 >>
rect 62 380 63 381 
<< m1 >>
rect 76 380 77 381 
<< m1 >>
rect 78 380 79 381 
<< m1 >>
rect 82 380 83 381 
<< m1 >>
rect 91 380 92 381 
<< m1 >>
rect 93 380 94 381 
<< m2 >>
rect 100 380 101 381 
<< m1 >>
rect 110 380 111 381 
<< m1 >>
rect 112 380 113 381 
<< m1 >>
rect 121 380 122 381 
<< m1 >>
rect 122 380 123 381 
<< m1 >>
rect 123 380 124 381 
<< m1 >>
rect 124 380 125 381 
<< m1 >>
rect 125 380 126 381 
<< m1 >>
rect 126 380 127 381 
<< m1 >>
rect 127 380 128 381 
<< m1 >>
rect 139 380 140 381 
<< m2 >>
rect 140 380 141 381 
<< m1 >>
rect 141 380 142 381 
<< m2 >>
rect 141 380 142 381 
<< m2c >>
rect 141 380 142 381 
<< m1 >>
rect 141 380 142 381 
<< m2 >>
rect 141 380 142 381 
<< m1 >>
rect 142 380 143 381 
<< m1 >>
rect 143 380 144 381 
<< m1 >>
rect 144 380 145 381 
<< m1 >>
rect 145 380 146 381 
<< m1 >>
rect 146 380 147 381 
<< m1 >>
rect 147 380 148 381 
<< m1 >>
rect 148 380 149 381 
<< m1 >>
rect 150 380 151 381 
<< m2 >>
rect 151 380 152 381 
<< m1 >>
rect 163 380 164 381 
<< m2 >>
rect 163 380 164 381 
<< m1 >>
rect 169 380 170 381 
<< m1 >>
rect 172 380 173 381 
<< m1 >>
rect 190 380 191 381 
<< m1 >>
rect 193 380 194 381 
<< m1 >>
rect 194 380 195 381 
<< m1 >>
rect 195 380 196 381 
<< m1 >>
rect 196 380 197 381 
<< m1 >>
rect 197 380 198 381 
<< m1 >>
rect 198 380 199 381 
<< m2 >>
rect 198 380 199 381 
<< m2c >>
rect 198 380 199 381 
<< m1 >>
rect 198 380 199 381 
<< m2 >>
rect 198 380 199 381 
<< m2 >>
rect 199 380 200 381 
<< m1 >>
rect 200 380 201 381 
<< m2 >>
rect 200 380 201 381 
<< m2 >>
rect 201 380 202 381 
<< m1 >>
rect 202 380 203 381 
<< m2 >>
rect 202 380 203 381 
<< m2c >>
rect 202 380 203 381 
<< m1 >>
rect 202 380 203 381 
<< m2 >>
rect 202 380 203 381 
<< m2 >>
rect 203 380 204 381 
<< m1 >>
rect 204 380 205 381 
<< m2 >>
rect 204 380 205 381 
<< m2 >>
rect 205 380 206 381 
<< m1 >>
rect 206 380 207 381 
<< m2 >>
rect 206 380 207 381 
<< m2c >>
rect 206 380 207 381 
<< m1 >>
rect 206 380 207 381 
<< m2 >>
rect 206 380 207 381 
<< m1 >>
rect 208 380 209 381 
<< m2 >>
rect 208 380 209 381 
<< m2c >>
rect 208 380 209 381 
<< m1 >>
rect 208 380 209 381 
<< m2 >>
rect 208 380 209 381 
<< m1 >>
rect 217 380 218 381 
<< m1 >>
rect 221 380 222 381 
<< m2 >>
rect 221 380 222 381 
<< m2c >>
rect 221 380 222 381 
<< m1 >>
rect 221 380 222 381 
<< m2 >>
rect 221 380 222 381 
<< m1 >>
rect 223 380 224 381 
<< m2 >>
rect 223 380 224 381 
<< m2c >>
rect 223 380 224 381 
<< m1 >>
rect 223 380 224 381 
<< m2 >>
rect 223 380 224 381 
<< m1 >>
rect 235 380 236 381 
<< m1 >>
rect 244 380 245 381 
<< m1 >>
rect 253 380 254 381 
<< m1 >>
rect 255 380 256 381 
<< m1 >>
rect 265 380 266 381 
<< m2 >>
rect 266 380 267 381 
<< m1 >>
rect 267 380 268 381 
<< m2 >>
rect 267 380 268 381 
<< m2c >>
rect 267 380 268 381 
<< m1 >>
rect 267 380 268 381 
<< m2 >>
rect 267 380 268 381 
<< m1 >>
rect 268 380 269 381 
<< m1 >>
rect 269 380 270 381 
<< m1 >>
rect 270 380 271 381 
<< m1 >>
rect 271 380 272 381 
<< m1 >>
rect 307 380 308 381 
<< m2 >>
rect 307 380 308 381 
<< m2c >>
rect 307 380 308 381 
<< m1 >>
rect 307 380 308 381 
<< m2 >>
rect 307 380 308 381 
<< m1 >>
rect 316 380 317 381 
<< m1 >>
rect 321 380 322 381 
<< m2 >>
rect 321 380 322 381 
<< m2c >>
rect 321 380 322 381 
<< m1 >>
rect 321 380 322 381 
<< m2 >>
rect 321 380 322 381 
<< m1 >>
rect 322 380 323 381 
<< m1 >>
rect 323 380 324 381 
<< m1 >>
rect 324 380 325 381 
<< m1 >>
rect 325 380 326 381 
<< m1 >>
rect 334 380 335 381 
<< m2 >>
rect 334 380 335 381 
<< m2c >>
rect 334 380 335 381 
<< m1 >>
rect 334 380 335 381 
<< m2 >>
rect 334 380 335 381 
<< m1 >>
rect 338 380 339 381 
<< m2 >>
rect 338 380 339 381 
<< m2c >>
rect 338 380 339 381 
<< m1 >>
rect 338 380 339 381 
<< m2 >>
rect 338 380 339 381 
<< m1 >>
rect 339 380 340 381 
<< m1 >>
rect 340 380 341 381 
<< m1 >>
rect 341 380 342 381 
<< m1 >>
rect 342 380 343 381 
<< m1 >>
rect 343 380 344 381 
<< m1 >>
rect 355 380 356 381 
<< m1 >>
rect 356 380 357 381 
<< m1 >>
rect 357 380 358 381 
<< m1 >>
rect 358 380 359 381 
<< m1 >>
rect 359 380 360 381 
<< m2 >>
rect 359 380 360 381 
<< m2c >>
rect 359 380 360 381 
<< m1 >>
rect 359 380 360 381 
<< m2 >>
rect 359 380 360 381 
<< m1 >>
rect 365 380 366 381 
<< m1 >>
rect 376 380 377 381 
<< m1 >>
rect 394 380 395 381 
<< m1 >>
rect 397 380 398 381 
<< m1 >>
rect 402 380 403 381 
<< m1 >>
rect 405 380 406 381 
<< m2 >>
rect 405 380 406 381 
<< m2c >>
rect 405 380 406 381 
<< m1 >>
rect 405 380 406 381 
<< m2 >>
rect 405 380 406 381 
<< m1 >>
rect 416 380 417 381 
<< m1 >>
rect 429 380 430 381 
<< m2 >>
rect 429 380 430 381 
<< m2c >>
rect 429 380 430 381 
<< m1 >>
rect 429 380 430 381 
<< m2 >>
rect 429 380 430 381 
<< m1 >>
rect 433 380 434 381 
<< m1 >>
rect 435 380 436 381 
<< m1 >>
rect 446 380 447 381 
<< m2 >>
rect 446 380 447 381 
<< m2c >>
rect 446 380 447 381 
<< m1 >>
rect 446 380 447 381 
<< m2 >>
rect 446 380 447 381 
<< m1 >>
rect 447 380 448 381 
<< m1 >>
rect 448 380 449 381 
<< m1 >>
rect 449 380 450 381 
<< m2 >>
rect 449 380 450 381 
<< m2c >>
rect 449 380 450 381 
<< m1 >>
rect 449 380 450 381 
<< m2 >>
rect 449 380 450 381 
<< m2 >>
rect 450 380 451 381 
<< m1 >>
rect 451 380 452 381 
<< m2 >>
rect 451 380 452 381 
<< m2 >>
rect 452 380 453 381 
<< m1 >>
rect 453 380 454 381 
<< m2 >>
rect 453 380 454 381 
<< m2c >>
rect 453 380 454 381 
<< m1 >>
rect 453 380 454 381 
<< m2 >>
rect 453 380 454 381 
<< m1 >>
rect 455 380 456 381 
<< m2 >>
rect 455 380 456 381 
<< m2c >>
rect 455 380 456 381 
<< m1 >>
rect 455 380 456 381 
<< m2 >>
rect 455 380 456 381 
<< m1 >>
rect 457 380 458 381 
<< m2 >>
rect 457 380 458 381 
<< m2c >>
rect 457 380 458 381 
<< m1 >>
rect 457 380 458 381 
<< m2 >>
rect 457 380 458 381 
<< m1 >>
rect 520 380 521 381 
<< m1 >>
rect 523 380 524 381 
<< m1 >>
rect 16 381 17 382 
<< m1 >>
rect 19 381 20 382 
<< m1 >>
rect 23 381 24 382 
<< m2 >>
rect 44 381 45 382 
<< m2 >>
rect 60 381 61 382 
<< m2 >>
rect 62 381 63 382 
<< m2 >>
rect 63 381 64 382 
<< m1 >>
rect 76 381 77 382 
<< m1 >>
rect 78 381 79 382 
<< m1 >>
rect 82 381 83 382 
<< m1 >>
rect 91 381 92 382 
<< m1 >>
rect 93 381 94 382 
<< m1 >>
rect 100 381 101 382 
<< m2 >>
rect 100 381 101 382 
<< m2c >>
rect 100 381 101 382 
<< m1 >>
rect 100 381 101 382 
<< m2 >>
rect 100 381 101 382 
<< m1 >>
rect 110 381 111 382 
<< m1 >>
rect 112 381 113 382 
<< m1 >>
rect 139 381 140 382 
<< m2 >>
rect 140 381 141 382 
<< m1 >>
rect 150 381 151 382 
<< m2 >>
rect 151 381 152 382 
<< m1 >>
rect 163 381 164 382 
<< m2 >>
rect 163 381 164 382 
<< m1 >>
rect 169 381 170 382 
<< m1 >>
rect 172 381 173 382 
<< m1 >>
rect 190 381 191 382 
<< m1 >>
rect 200 381 201 382 
<< m1 >>
rect 204 381 205 382 
<< m1 >>
rect 206 381 207 382 
<< m2 >>
rect 208 381 209 382 
<< m1 >>
rect 212 381 213 382 
<< m1 >>
rect 213 381 214 382 
<< m1 >>
rect 214 381 215 382 
<< m1 >>
rect 215 381 216 382 
<< m2 >>
rect 215 381 216 382 
<< m2c >>
rect 215 381 216 382 
<< m1 >>
rect 215 381 216 382 
<< m2 >>
rect 215 381 216 382 
<< m2 >>
rect 216 381 217 382 
<< m1 >>
rect 217 381 218 382 
<< m2 >>
rect 217 381 218 382 
<< m2 >>
rect 218 381 219 382 
<< m1 >>
rect 219 381 220 382 
<< m2 >>
rect 219 381 220 382 
<< m2c >>
rect 219 381 220 382 
<< m1 >>
rect 219 381 220 382 
<< m2 >>
rect 219 381 220 382 
<< m2 >>
rect 221 381 222 382 
<< m2 >>
rect 223 381 224 382 
<< m1 >>
rect 235 381 236 382 
<< m1 >>
rect 237 381 238 382 
<< m1 >>
rect 238 381 239 382 
<< m1 >>
rect 239 381 240 382 
<< m1 >>
rect 240 381 241 382 
<< m1 >>
rect 241 381 242 382 
<< m1 >>
rect 242 381 243 382 
<< m2 >>
rect 242 381 243 382 
<< m2c >>
rect 242 381 243 382 
<< m1 >>
rect 242 381 243 382 
<< m2 >>
rect 242 381 243 382 
<< m2 >>
rect 243 381 244 382 
<< m1 >>
rect 244 381 245 382 
<< m2 >>
rect 244 381 245 382 
<< m2 >>
rect 245 381 246 382 
<< m1 >>
rect 246 381 247 382 
<< m2 >>
rect 246 381 247 382 
<< m2c >>
rect 246 381 247 382 
<< m1 >>
rect 246 381 247 382 
<< m2 >>
rect 246 381 247 382 
<< m1 >>
rect 248 381 249 382 
<< m1 >>
rect 249 381 250 382 
<< m1 >>
rect 250 381 251 382 
<< m1 >>
rect 251 381 252 382 
<< m2 >>
rect 251 381 252 382 
<< m2c >>
rect 251 381 252 382 
<< m1 >>
rect 251 381 252 382 
<< m2 >>
rect 251 381 252 382 
<< m2 >>
rect 252 381 253 382 
<< m1 >>
rect 253 381 254 382 
<< m2 >>
rect 253 381 254 382 
<< m2 >>
rect 254 381 255 382 
<< m1 >>
rect 255 381 256 382 
<< m2 >>
rect 255 381 256 382 
<< m2 >>
rect 256 381 257 382 
<< m1 >>
rect 257 381 258 382 
<< m2 >>
rect 257 381 258 382 
<< m2c >>
rect 257 381 258 382 
<< m1 >>
rect 257 381 258 382 
<< m2 >>
rect 257 381 258 382 
<< m1 >>
rect 265 381 266 382 
<< m2 >>
rect 266 381 267 382 
<< m2 >>
rect 307 381 308 382 
<< m1 >>
rect 316 381 317 382 
<< m2 >>
rect 321 381 322 382 
<< m2 >>
rect 323 381 324 382 
<< m2 >>
rect 324 381 325 382 
<< m2 >>
rect 325 381 326 382 
<< m2 >>
rect 326 381 327 382 
<< m2 >>
rect 327 381 328 382 
<< m2 >>
rect 328 381 329 382 
<< m2 >>
rect 329 381 330 382 
<< m2 >>
rect 330 381 331 382 
<< m2 >>
rect 331 381 332 382 
<< m2 >>
rect 332 381 333 382 
<< m2 >>
rect 333 381 334 382 
<< m2 >>
rect 334 381 335 382 
<< m2 >>
rect 338 381 339 382 
<< m2 >>
rect 359 381 360 382 
<< m1 >>
rect 365 381 366 382 
<< m1 >>
rect 376 381 377 382 
<< m1 >>
rect 394 381 395 382 
<< m1 >>
rect 397 381 398 382 
<< m1 >>
rect 402 381 403 382 
<< m2 >>
rect 405 381 406 382 
<< m1 >>
rect 416 381 417 382 
<< m2 >>
rect 429 381 430 382 
<< m1 >>
rect 433 381 434 382 
<< m1 >>
rect 435 381 436 382 
<< m2 >>
rect 446 381 447 382 
<< m1 >>
rect 451 381 452 382 
<< m2 >>
rect 455 381 456 382 
<< m2 >>
rect 457 381 458 382 
<< m1 >>
rect 520 381 521 382 
<< m1 >>
rect 523 381 524 382 
<< m1 >>
rect 13 382 14 383 
<< m1 >>
rect 14 382 15 383 
<< m1 >>
rect 15 382 16 383 
<< m1 >>
rect 16 382 17 383 
<< m1 >>
rect 19 382 20 383 
<< m1 >>
rect 23 382 24 383 
<< m1 >>
rect 31 382 32 383 
<< m1 >>
rect 32 382 33 383 
<< m1 >>
rect 33 382 34 383 
<< m1 >>
rect 34 382 35 383 
<< m1 >>
rect 35 382 36 383 
<< m1 >>
rect 36 382 37 383 
<< m1 >>
rect 37 382 38 383 
<< m1 >>
rect 38 382 39 383 
<< m1 >>
rect 39 382 40 383 
<< m1 >>
rect 40 382 41 383 
<< m1 >>
rect 41 382 42 383 
<< m1 >>
rect 42 382 43 383 
<< m1 >>
rect 43 382 44 383 
<< m1 >>
rect 44 382 45 383 
<< m2 >>
rect 44 382 45 383 
<< m1 >>
rect 45 382 46 383 
<< m1 >>
rect 46 382 47 383 
<< m1 >>
rect 47 382 48 383 
<< m1 >>
rect 48 382 49 383 
<< m2 >>
rect 48 382 49 383 
<< m1 >>
rect 49 382 50 383 
<< m2 >>
rect 49 382 50 383 
<< m1 >>
rect 50 382 51 383 
<< m2 >>
rect 50 382 51 383 
<< m1 >>
rect 51 382 52 383 
<< m2 >>
rect 51 382 52 383 
<< m1 >>
rect 52 382 53 383 
<< m2 >>
rect 52 382 53 383 
<< m1 >>
rect 53 382 54 383 
<< m2 >>
rect 53 382 54 383 
<< m1 >>
rect 54 382 55 383 
<< m2 >>
rect 54 382 55 383 
<< m1 >>
rect 55 382 56 383 
<< m2 >>
rect 55 382 56 383 
<< m1 >>
rect 56 382 57 383 
<< m2 >>
rect 56 382 57 383 
<< m1 >>
rect 57 382 58 383 
<< m2 >>
rect 57 382 58 383 
<< m1 >>
rect 58 382 59 383 
<< m2 >>
rect 58 382 59 383 
<< m1 >>
rect 59 382 60 383 
<< m2 >>
rect 59 382 60 383 
<< m1 >>
rect 60 382 61 383 
<< m2 >>
rect 60 382 61 383 
<< m1 >>
rect 61 382 62 383 
<< m1 >>
rect 62 382 63 383 
<< m1 >>
rect 63 382 64 383 
<< m2 >>
rect 63 382 64 383 
<< m1 >>
rect 64 382 65 383 
<< m1 >>
rect 65 382 66 383 
<< m1 >>
rect 66 382 67 383 
<< m1 >>
rect 67 382 68 383 
<< m1 >>
rect 68 382 69 383 
<< m1 >>
rect 69 382 70 383 
<< m1 >>
rect 70 382 71 383 
<< m1 >>
rect 71 382 72 383 
<< m1 >>
rect 72 382 73 383 
<< m1 >>
rect 73 382 74 383 
<< m1 >>
rect 74 382 75 383 
<< m1 >>
rect 75 382 76 383 
<< m1 >>
rect 76 382 77 383 
<< m1 >>
rect 78 382 79 383 
<< m1 >>
rect 82 382 83 383 
<< m1 >>
rect 91 382 92 383 
<< m1 >>
rect 93 382 94 383 
<< m1 >>
rect 100 382 101 383 
<< m1 >>
rect 110 382 111 383 
<< m1 >>
rect 112 382 113 383 
<< m1 >>
rect 118 382 119 383 
<< m1 >>
rect 119 382 120 383 
<< m1 >>
rect 120 382 121 383 
<< m1 >>
rect 121 382 122 383 
<< m1 >>
rect 122 382 123 383 
<< m1 >>
rect 123 382 124 383 
<< m1 >>
rect 124 382 125 383 
<< m1 >>
rect 125 382 126 383 
<< m1 >>
rect 126 382 127 383 
<< m1 >>
rect 127 382 128 383 
<< m1 >>
rect 128 382 129 383 
<< m1 >>
rect 129 382 130 383 
<< m1 >>
rect 130 382 131 383 
<< m1 >>
rect 131 382 132 383 
<< m1 >>
rect 132 382 133 383 
<< m1 >>
rect 133 382 134 383 
<< m1 >>
rect 134 382 135 383 
<< m1 >>
rect 135 382 136 383 
<< m1 >>
rect 136 382 137 383 
<< m1 >>
rect 137 382 138 383 
<< m2 >>
rect 137 382 138 383 
<< m2c >>
rect 137 382 138 383 
<< m1 >>
rect 137 382 138 383 
<< m2 >>
rect 137 382 138 383 
<< m2 >>
rect 138 382 139 383 
<< m1 >>
rect 139 382 140 383 
<< m2 >>
rect 139 382 140 383 
<< m2 >>
rect 140 382 141 383 
<< m1 >>
rect 148 382 149 383 
<< m2 >>
rect 148 382 149 383 
<< m2c >>
rect 148 382 149 383 
<< m1 >>
rect 148 382 149 383 
<< m2 >>
rect 148 382 149 383 
<< m2 >>
rect 149 382 150 383 
<< m1 >>
rect 150 382 151 383 
<< m2 >>
rect 150 382 151 383 
<< m2 >>
rect 151 382 152 383 
<< m1 >>
rect 163 382 164 383 
<< m2 >>
rect 163 382 164 383 
<< m1 >>
rect 167 382 168 383 
<< m2 >>
rect 167 382 168 383 
<< m2c >>
rect 167 382 168 383 
<< m1 >>
rect 167 382 168 383 
<< m2 >>
rect 167 382 168 383 
<< m2 >>
rect 168 382 169 383 
<< m1 >>
rect 169 382 170 383 
<< m2 >>
rect 169 382 170 383 
<< m2 >>
rect 170 382 171 383 
<< m2 >>
rect 171 382 172 383 
<< m1 >>
rect 172 382 173 383 
<< m2 >>
rect 172 382 173 383 
<< m2 >>
rect 173 382 174 383 
<< m1 >>
rect 174 382 175 383 
<< m2 >>
rect 174 382 175 383 
<< m2c >>
rect 174 382 175 383 
<< m1 >>
rect 174 382 175 383 
<< m2 >>
rect 174 382 175 383 
<< m1 >>
rect 175 382 176 383 
<< m1 >>
rect 176 382 177 383 
<< m1 >>
rect 177 382 178 383 
<< m1 >>
rect 178 382 179 383 
<< m1 >>
rect 179 382 180 383 
<< m1 >>
rect 180 382 181 383 
<< m1 >>
rect 181 382 182 383 
<< m1 >>
rect 182 382 183 383 
<< m1 >>
rect 183 382 184 383 
<< m1 >>
rect 184 382 185 383 
<< m1 >>
rect 185 382 186 383 
<< m1 >>
rect 186 382 187 383 
<< m1 >>
rect 187 382 188 383 
<< m1 >>
rect 188 382 189 383 
<< m1 >>
rect 189 382 190 383 
<< m1 >>
rect 190 382 191 383 
<< m1 >>
rect 200 382 201 383 
<< m1 >>
rect 204 382 205 383 
<< m1 >>
rect 206 382 207 383 
<< m1 >>
rect 207 382 208 383 
<< m1 >>
rect 208 382 209 383 
<< m2 >>
rect 208 382 209 383 
<< m1 >>
rect 209 382 210 383 
<< m1 >>
rect 210 382 211 383 
<< m1 >>
rect 211 382 212 383 
<< m1 >>
rect 212 382 213 383 
<< m1 >>
rect 217 382 218 383 
<< m1 >>
rect 219 382 220 383 
<< m1 >>
rect 220 382 221 383 
<< m1 >>
rect 221 382 222 383 
<< m2 >>
rect 221 382 222 383 
<< m1 >>
rect 222 382 223 383 
<< m1 >>
rect 223 382 224 383 
<< m2 >>
rect 223 382 224 383 
<< m1 >>
rect 224 382 225 383 
<< m1 >>
rect 225 382 226 383 
<< m1 >>
rect 226 382 227 383 
<< m1 >>
rect 227 382 228 383 
<< m1 >>
rect 228 382 229 383 
<< m1 >>
rect 229 382 230 383 
<< m1 >>
rect 230 382 231 383 
<< m1 >>
rect 231 382 232 383 
<< m1 >>
rect 232 382 233 383 
<< m1 >>
rect 233 382 234 383 
<< m2 >>
rect 233 382 234 383 
<< m2c >>
rect 233 382 234 383 
<< m1 >>
rect 233 382 234 383 
<< m2 >>
rect 233 382 234 383 
<< m2 >>
rect 234 382 235 383 
<< m1 >>
rect 235 382 236 383 
<< m2 >>
rect 235 382 236 383 
<< m2 >>
rect 236 382 237 383 
<< m1 >>
rect 237 382 238 383 
<< m2 >>
rect 237 382 238 383 
<< m2c >>
rect 237 382 238 383 
<< m1 >>
rect 237 382 238 383 
<< m2 >>
rect 237 382 238 383 
<< m1 >>
rect 244 382 245 383 
<< m1 >>
rect 246 382 247 383 
<< m1 >>
rect 247 382 248 383 
<< m1 >>
rect 248 382 249 383 
<< m1 >>
rect 253 382 254 383 
<< m1 >>
rect 255 382 256 383 
<< m1 >>
rect 257 382 258 383 
<< m1 >>
rect 265 382 266 383 
<< m1 >>
rect 266 382 267 383 
<< m2 >>
rect 266 382 267 383 
<< m1 >>
rect 267 382 268 383 
<< m1 >>
rect 268 382 269 383 
<< m1 >>
rect 269 382 270 383 
<< m1 >>
rect 270 382 271 383 
<< m1 >>
rect 271 382 272 383 
<< m1 >>
rect 272 382 273 383 
<< m1 >>
rect 273 382 274 383 
<< m1 >>
rect 274 382 275 383 
<< m1 >>
rect 275 382 276 383 
<< m1 >>
rect 276 382 277 383 
<< m1 >>
rect 277 382 278 383 
<< m1 >>
rect 278 382 279 383 
<< m1 >>
rect 279 382 280 383 
<< m1 >>
rect 280 382 281 383 
<< m1 >>
rect 281 382 282 383 
<< m1 >>
rect 282 382 283 383 
<< m1 >>
rect 283 382 284 383 
<< m1 >>
rect 284 382 285 383 
<< m1 >>
rect 285 382 286 383 
<< m1 >>
rect 286 382 287 383 
<< m1 >>
rect 287 382 288 383 
<< m1 >>
rect 288 382 289 383 
<< m1 >>
rect 289 382 290 383 
<< m1 >>
rect 290 382 291 383 
<< m1 >>
rect 291 382 292 383 
<< m1 >>
rect 292 382 293 383 
<< m1 >>
rect 293 382 294 383 
<< m1 >>
rect 294 382 295 383 
<< m1 >>
rect 295 382 296 383 
<< m1 >>
rect 296 382 297 383 
<< m1 >>
rect 297 382 298 383 
<< m1 >>
rect 298 382 299 383 
<< m1 >>
rect 299 382 300 383 
<< m1 >>
rect 300 382 301 383 
<< m1 >>
rect 301 382 302 383 
<< m1 >>
rect 302 382 303 383 
<< m1 >>
rect 303 382 304 383 
<< m1 >>
rect 304 382 305 383 
<< m1 >>
rect 305 382 306 383 
<< m1 >>
rect 306 382 307 383 
<< m1 >>
rect 307 382 308 383 
<< m2 >>
rect 307 382 308 383 
<< m1 >>
rect 308 382 309 383 
<< m1 >>
rect 309 382 310 383 
<< m1 >>
rect 310 382 311 383 
<< m1 >>
rect 311 382 312 383 
<< m1 >>
rect 312 382 313 383 
<< m1 >>
rect 313 382 314 383 
<< m1 >>
rect 314 382 315 383 
<< m2 >>
rect 314 382 315 383 
<< m2c >>
rect 314 382 315 383 
<< m1 >>
rect 314 382 315 383 
<< m2 >>
rect 314 382 315 383 
<< m2 >>
rect 315 382 316 383 
<< m1 >>
rect 316 382 317 383 
<< m2 >>
rect 316 382 317 383 
<< m2 >>
rect 317 382 318 383 
<< m1 >>
rect 318 382 319 383 
<< m2 >>
rect 318 382 319 383 
<< m2c >>
rect 318 382 319 383 
<< m1 >>
rect 318 382 319 383 
<< m2 >>
rect 318 382 319 383 
<< m1 >>
rect 319 382 320 383 
<< m1 >>
rect 320 382 321 383 
<< m1 >>
rect 321 382 322 383 
<< m2 >>
rect 321 382 322 383 
<< m1 >>
rect 322 382 323 383 
<< m1 >>
rect 323 382 324 383 
<< m2 >>
rect 323 382 324 383 
<< m1 >>
rect 324 382 325 383 
<< m1 >>
rect 325 382 326 383 
<< m1 >>
rect 326 382 327 383 
<< m1 >>
rect 327 382 328 383 
<< m1 >>
rect 328 382 329 383 
<< m1 >>
rect 329 382 330 383 
<< m1 >>
rect 330 382 331 383 
<< m1 >>
rect 331 382 332 383 
<< m1 >>
rect 332 382 333 383 
<< m1 >>
rect 333 382 334 383 
<< m1 >>
rect 334 382 335 383 
<< m1 >>
rect 335 382 336 383 
<< m1 >>
rect 336 382 337 383 
<< m1 >>
rect 337 382 338 383 
<< m1 >>
rect 338 382 339 383 
<< m2 >>
rect 338 382 339 383 
<< m1 >>
rect 339 382 340 383 
<< m1 >>
rect 340 382 341 383 
<< m1 >>
rect 341 382 342 383 
<< m1 >>
rect 342 382 343 383 
<< m1 >>
rect 343 382 344 383 
<< m1 >>
rect 344 382 345 383 
<< m1 >>
rect 345 382 346 383 
<< m1 >>
rect 346 382 347 383 
<< m1 >>
rect 347 382 348 383 
<< m1 >>
rect 348 382 349 383 
<< m1 >>
rect 349 382 350 383 
<< m1 >>
rect 350 382 351 383 
<< m1 >>
rect 351 382 352 383 
<< m1 >>
rect 352 382 353 383 
<< m1 >>
rect 353 382 354 383 
<< m1 >>
rect 354 382 355 383 
<< m1 >>
rect 355 382 356 383 
<< m1 >>
rect 356 382 357 383 
<< m1 >>
rect 357 382 358 383 
<< m1 >>
rect 358 382 359 383 
<< m1 >>
rect 359 382 360 383 
<< m2 >>
rect 359 382 360 383 
<< m1 >>
rect 360 382 361 383 
<< m1 >>
rect 361 382 362 383 
<< m1 >>
rect 362 382 363 383 
<< m1 >>
rect 363 382 364 383 
<< m1 >>
rect 365 382 366 383 
<< m1 >>
rect 366 382 367 383 
<< m1 >>
rect 367 382 368 383 
<< m1 >>
rect 368 382 369 383 
<< m1 >>
rect 369 382 370 383 
<< m1 >>
rect 370 382 371 383 
<< m1 >>
rect 371 382 372 383 
<< m1 >>
rect 372 382 373 383 
<< m1 >>
rect 373 382 374 383 
<< m1 >>
rect 374 382 375 383 
<< m1 >>
rect 375 382 376 383 
<< m1 >>
rect 376 382 377 383 
<< m1 >>
rect 394 382 395 383 
<< m1 >>
rect 397 382 398 383 
<< m1 >>
rect 402 382 403 383 
<< m2 >>
rect 405 382 406 383 
<< m1 >>
rect 406 382 407 383 
<< m2 >>
rect 406 382 407 383 
<< m1 >>
rect 407 382 408 383 
<< m2 >>
rect 407 382 408 383 
<< m1 >>
rect 408 382 409 383 
<< m2 >>
rect 408 382 409 383 
<< m1 >>
rect 409 382 410 383 
<< m2 >>
rect 409 382 410 383 
<< m1 >>
rect 410 382 411 383 
<< m2 >>
rect 410 382 411 383 
<< m1 >>
rect 411 382 412 383 
<< m1 >>
rect 412 382 413 383 
<< m1 >>
rect 413 382 414 383 
<< m1 >>
rect 414 382 415 383 
<< m2 >>
rect 414 382 415 383 
<< m2c >>
rect 414 382 415 383 
<< m1 >>
rect 414 382 415 383 
<< m2 >>
rect 414 382 415 383 
<< m2 >>
rect 415 382 416 383 
<< m1 >>
rect 416 382 417 383 
<< m2 >>
rect 416 382 417 383 
<< m2 >>
rect 417 382 418 383 
<< m1 >>
rect 418 382 419 383 
<< m2 >>
rect 418 382 419 383 
<< m2c >>
rect 418 382 419 383 
<< m1 >>
rect 418 382 419 383 
<< m2 >>
rect 418 382 419 383 
<< m1 >>
rect 419 382 420 383 
<< m1 >>
rect 420 382 421 383 
<< m1 >>
rect 421 382 422 383 
<< m1 >>
rect 422 382 423 383 
<< m1 >>
rect 423 382 424 383 
<< m1 >>
rect 424 382 425 383 
<< m1 >>
rect 425 382 426 383 
<< m1 >>
rect 426 382 427 383 
<< m1 >>
rect 427 382 428 383 
<< m1 >>
rect 428 382 429 383 
<< m1 >>
rect 429 382 430 383 
<< m2 >>
rect 429 382 430 383 
<< m1 >>
rect 430 382 431 383 
<< m1 >>
rect 431 382 432 383 
<< m2 >>
rect 431 382 432 383 
<< m2c >>
rect 431 382 432 383 
<< m1 >>
rect 431 382 432 383 
<< m2 >>
rect 431 382 432 383 
<< m2 >>
rect 432 382 433 383 
<< m1 >>
rect 433 382 434 383 
<< m2 >>
rect 433 382 434 383 
<< m2 >>
rect 434 382 435 383 
<< m1 >>
rect 435 382 436 383 
<< m2 >>
rect 435 382 436 383 
<< m2 >>
rect 436 382 437 383 
<< m1 >>
rect 437 382 438 383 
<< m2 >>
rect 437 382 438 383 
<< m2c >>
rect 437 382 438 383 
<< m1 >>
rect 437 382 438 383 
<< m2 >>
rect 437 382 438 383 
<< m1 >>
rect 438 382 439 383 
<< m1 >>
rect 439 382 440 383 
<< m1 >>
rect 440 382 441 383 
<< m1 >>
rect 441 382 442 383 
<< m1 >>
rect 442 382 443 383 
<< m1 >>
rect 443 382 444 383 
<< m1 >>
rect 444 382 445 383 
<< m1 >>
rect 445 382 446 383 
<< m1 >>
rect 446 382 447 383 
<< m2 >>
rect 446 382 447 383 
<< m1 >>
rect 447 382 448 383 
<< m1 >>
rect 448 382 449 383 
<< m1 >>
rect 449 382 450 383 
<< m2 >>
rect 449 382 450 383 
<< m2c >>
rect 449 382 450 383 
<< m1 >>
rect 449 382 450 383 
<< m2 >>
rect 449 382 450 383 
<< m2 >>
rect 450 382 451 383 
<< m1 >>
rect 451 382 452 383 
<< m2 >>
rect 451 382 452 383 
<< m2 >>
rect 452 382 453 383 
<< m1 >>
rect 453 382 454 383 
<< m2 >>
rect 453 382 454 383 
<< m2c >>
rect 453 382 454 383 
<< m1 >>
rect 453 382 454 383 
<< m2 >>
rect 453 382 454 383 
<< m1 >>
rect 454 382 455 383 
<< m1 >>
rect 455 382 456 383 
<< m2 >>
rect 455 382 456 383 
<< m1 >>
rect 456 382 457 383 
<< m1 >>
rect 457 382 458 383 
<< m2 >>
rect 457 382 458 383 
<< m1 >>
rect 458 382 459 383 
<< m1 >>
rect 459 382 460 383 
<< m1 >>
rect 460 382 461 383 
<< m1 >>
rect 461 382 462 383 
<< m1 >>
rect 462 382 463 383 
<< m1 >>
rect 463 382 464 383 
<< m1 >>
rect 464 382 465 383 
<< m1 >>
rect 465 382 466 383 
<< m1 >>
rect 466 382 467 383 
<< m1 >>
rect 467 382 468 383 
<< m1 >>
rect 468 382 469 383 
<< m1 >>
rect 469 382 470 383 
<< m1 >>
rect 470 382 471 383 
<< m1 >>
rect 471 382 472 383 
<< m1 >>
rect 472 382 473 383 
<< m1 >>
rect 473 382 474 383 
<< m1 >>
rect 474 382 475 383 
<< m1 >>
rect 475 382 476 383 
<< m1 >>
rect 476 382 477 383 
<< m1 >>
rect 477 382 478 383 
<< m1 >>
rect 478 382 479 383 
<< m1 >>
rect 479 382 480 383 
<< m1 >>
rect 480 382 481 383 
<< m1 >>
rect 481 382 482 383 
<< m1 >>
rect 482 382 483 383 
<< m1 >>
rect 483 382 484 383 
<< m1 >>
rect 484 382 485 383 
<< m1 >>
rect 485 382 486 383 
<< m1 >>
rect 486 382 487 383 
<< m1 >>
rect 487 382 488 383 
<< m1 >>
rect 488 382 489 383 
<< m1 >>
rect 489 382 490 383 
<< m1 >>
rect 490 382 491 383 
<< m1 >>
rect 491 382 492 383 
<< m1 >>
rect 492 382 493 383 
<< m1 >>
rect 493 382 494 383 
<< m1 >>
rect 494 382 495 383 
<< m1 >>
rect 495 382 496 383 
<< m1 >>
rect 496 382 497 383 
<< m1 >>
rect 497 382 498 383 
<< m1 >>
rect 498 382 499 383 
<< m1 >>
rect 499 382 500 383 
<< m1 >>
rect 500 382 501 383 
<< m1 >>
rect 501 382 502 383 
<< m1 >>
rect 502 382 503 383 
<< m1 >>
rect 503 382 504 383 
<< m1 >>
rect 504 382 505 383 
<< m1 >>
rect 505 382 506 383 
<< m1 >>
rect 506 382 507 383 
<< m1 >>
rect 507 382 508 383 
<< m1 >>
rect 508 382 509 383 
<< m1 >>
rect 509 382 510 383 
<< m1 >>
rect 510 382 511 383 
<< m1 >>
rect 511 382 512 383 
<< m1 >>
rect 512 382 513 383 
<< m1 >>
rect 513 382 514 383 
<< m1 >>
rect 514 382 515 383 
<< m1 >>
rect 515 382 516 383 
<< m1 >>
rect 516 382 517 383 
<< m1 >>
rect 517 382 518 383 
<< m1 >>
rect 518 382 519 383 
<< m1 >>
rect 519 382 520 383 
<< m1 >>
rect 520 382 521 383 
<< m1 >>
rect 523 382 524 383 
<< m1 >>
rect 13 383 14 384 
<< m1 >>
rect 19 383 20 384 
<< m1 >>
rect 23 383 24 384 
<< m2 >>
rect 23 383 24 384 
<< m2c >>
rect 23 383 24 384 
<< m1 >>
rect 23 383 24 384 
<< m2 >>
rect 23 383 24 384 
<< m1 >>
rect 31 383 32 384 
<< m2 >>
rect 44 383 45 384 
<< m2 >>
rect 48 383 49 384 
<< m2 >>
rect 63 383 64 384 
<< m2 >>
rect 73 383 74 384 
<< m2 >>
rect 74 383 75 384 
<< m2 >>
rect 75 383 76 384 
<< m2 >>
rect 76 383 77 384 
<< m2 >>
rect 77 383 78 384 
<< m1 >>
rect 78 383 79 384 
<< m2 >>
rect 78 383 79 384 
<< m2 >>
rect 79 383 80 384 
<< m1 >>
rect 80 383 81 384 
<< m2 >>
rect 80 383 81 384 
<< m2c >>
rect 80 383 81 384 
<< m1 >>
rect 80 383 81 384 
<< m2 >>
rect 80 383 81 384 
<< m2 >>
rect 81 383 82 384 
<< m1 >>
rect 82 383 83 384 
<< m2 >>
rect 82 383 83 384 
<< m2 >>
rect 83 383 84 384 
<< m1 >>
rect 84 383 85 384 
<< m2 >>
rect 84 383 85 384 
<< m2c >>
rect 84 383 85 384 
<< m1 >>
rect 84 383 85 384 
<< m2 >>
rect 84 383 85 384 
<< m1 >>
rect 85 383 86 384 
<< m1 >>
rect 86 383 87 384 
<< m1 >>
rect 87 383 88 384 
<< m1 >>
rect 88 383 89 384 
<< m1 >>
rect 89 383 90 384 
<< m1 >>
rect 90 383 91 384 
<< m1 >>
rect 91 383 92 384 
<< m1 >>
rect 93 383 94 384 
<< m2 >>
rect 93 383 94 384 
<< m2c >>
rect 93 383 94 384 
<< m1 >>
rect 93 383 94 384 
<< m2 >>
rect 93 383 94 384 
<< m1 >>
rect 100 383 101 384 
<< m2 >>
rect 100 383 101 384 
<< m2c >>
rect 100 383 101 384 
<< m1 >>
rect 100 383 101 384 
<< m2 >>
rect 100 383 101 384 
<< m1 >>
rect 110 383 111 384 
<< m2 >>
rect 110 383 111 384 
<< m2c >>
rect 110 383 111 384 
<< m1 >>
rect 110 383 111 384 
<< m2 >>
rect 110 383 111 384 
<< m1 >>
rect 112 383 113 384 
<< m2 >>
rect 112 383 113 384 
<< m2c >>
rect 112 383 113 384 
<< m1 >>
rect 112 383 113 384 
<< m2 >>
rect 112 383 113 384 
<< m1 >>
rect 114 383 115 384 
<< m2 >>
rect 114 383 115 384 
<< m2c >>
rect 114 383 115 384 
<< m1 >>
rect 114 383 115 384 
<< m2 >>
rect 114 383 115 384 
<< m1 >>
rect 115 383 116 384 
<< m1 >>
rect 116 383 117 384 
<< m2 >>
rect 116 383 117 384 
<< m2c >>
rect 116 383 117 384 
<< m1 >>
rect 116 383 117 384 
<< m2 >>
rect 116 383 117 384 
<< m2 >>
rect 117 383 118 384 
<< m1 >>
rect 118 383 119 384 
<< m2 >>
rect 118 383 119 384 
<< m2 >>
rect 119 383 120 384 
<< m2 >>
rect 120 383 121 384 
<< m2 >>
rect 121 383 122 384 
<< m2 >>
rect 122 383 123 384 
<< m2 >>
rect 123 383 124 384 
<< m2 >>
rect 124 383 125 384 
<< m2 >>
rect 125 383 126 384 
<< m2 >>
rect 126 383 127 384 
<< m2 >>
rect 127 383 128 384 
<< m2 >>
rect 128 383 129 384 
<< m2 >>
rect 129 383 130 384 
<< m2 >>
rect 130 383 131 384 
<< m2 >>
rect 131 383 132 384 
<< m2 >>
rect 132 383 133 384 
<< m2 >>
rect 133 383 134 384 
<< m2 >>
rect 134 383 135 384 
<< m2 >>
rect 135 383 136 384 
<< m1 >>
rect 139 383 140 384 
<< m1 >>
rect 148 383 149 384 
<< m1 >>
rect 150 383 151 384 
<< m1 >>
rect 163 383 164 384 
<< m2 >>
rect 163 383 164 384 
<< m1 >>
rect 167 383 168 384 
<< m1 >>
rect 169 383 170 384 
<< m1 >>
rect 172 383 173 384 
<< m1 >>
rect 196 383 197 384 
<< m2 >>
rect 196 383 197 384 
<< m2c >>
rect 196 383 197 384 
<< m1 >>
rect 196 383 197 384 
<< m2 >>
rect 196 383 197 384 
<< m1 >>
rect 197 383 198 384 
<< m1 >>
rect 198 383 199 384 
<< m1 >>
rect 199 383 200 384 
<< m2 >>
rect 199 383 200 384 
<< m1 >>
rect 200 383 201 384 
<< m2 >>
rect 200 383 201 384 
<< m2 >>
rect 201 383 202 384 
<< m1 >>
rect 202 383 203 384 
<< m2 >>
rect 202 383 203 384 
<< m2c >>
rect 202 383 203 384 
<< m1 >>
rect 202 383 203 384 
<< m2 >>
rect 202 383 203 384 
<< m1 >>
rect 203 383 204 384 
<< m1 >>
rect 204 383 205 384 
<< m2 >>
rect 208 383 209 384 
<< m1 >>
rect 217 383 218 384 
<< m2 >>
rect 217 383 218 384 
<< m2c >>
rect 217 383 218 384 
<< m1 >>
rect 217 383 218 384 
<< m2 >>
rect 217 383 218 384 
<< m2 >>
rect 221 383 222 384 
<< m2 >>
rect 223 383 224 384 
<< m1 >>
rect 235 383 236 384 
<< m1 >>
rect 244 383 245 384 
<< m2 >>
rect 244 383 245 384 
<< m2c >>
rect 244 383 245 384 
<< m1 >>
rect 244 383 245 384 
<< m2 >>
rect 244 383 245 384 
<< m1 >>
rect 253 383 254 384 
<< m2 >>
rect 253 383 254 384 
<< m2c >>
rect 253 383 254 384 
<< m1 >>
rect 253 383 254 384 
<< m2 >>
rect 253 383 254 384 
<< m1 >>
rect 255 383 256 384 
<< m2 >>
rect 255 383 256 384 
<< m2c >>
rect 255 383 256 384 
<< m1 >>
rect 255 383 256 384 
<< m2 >>
rect 255 383 256 384 
<< m1 >>
rect 257 383 258 384 
<< m2 >>
rect 257 383 258 384 
<< m2c >>
rect 257 383 258 384 
<< m1 >>
rect 257 383 258 384 
<< m2 >>
rect 257 383 258 384 
<< m2 >>
rect 264 383 265 384 
<< m2 >>
rect 265 383 266 384 
<< m2 >>
rect 266 383 267 384 
<< m2 >>
rect 307 383 308 384 
<< m1 >>
rect 316 383 317 384 
<< m2 >>
rect 321 383 322 384 
<< m2 >>
rect 323 383 324 384 
<< m2 >>
rect 325 383 326 384 
<< m2 >>
rect 326 383 327 384 
<< m2 >>
rect 327 383 328 384 
<< m2 >>
rect 328 383 329 384 
<< m2 >>
rect 329 383 330 384 
<< m2 >>
rect 330 383 331 384 
<< m2 >>
rect 331 383 332 384 
<< m2 >>
rect 332 383 333 384 
<< m2 >>
rect 333 383 334 384 
<< m2 >>
rect 334 383 335 384 
<< m2 >>
rect 335 383 336 384 
<< m2 >>
rect 336 383 337 384 
<< m2 >>
rect 337 383 338 384 
<< m2 >>
rect 338 383 339 384 
<< m2 >>
rect 359 383 360 384 
<< m1 >>
rect 363 383 364 384 
<< m2 >>
rect 367 383 368 384 
<< m2 >>
rect 368 383 369 384 
<< m2 >>
rect 369 383 370 384 
<< m2 >>
rect 370 383 371 384 
<< m2 >>
rect 371 383 372 384 
<< m2 >>
rect 372 383 373 384 
<< m2 >>
rect 373 383 374 384 
<< m2 >>
rect 374 383 375 384 
<< m2 >>
rect 375 383 376 384 
<< m2 >>
rect 376 383 377 384 
<< m2 >>
rect 377 383 378 384 
<< m1 >>
rect 378 383 379 384 
<< m2 >>
rect 378 383 379 384 
<< m2c >>
rect 378 383 379 384 
<< m1 >>
rect 378 383 379 384 
<< m2 >>
rect 378 383 379 384 
<< m1 >>
rect 379 383 380 384 
<< m1 >>
rect 380 383 381 384 
<< m1 >>
rect 381 383 382 384 
<< m1 >>
rect 382 383 383 384 
<< m1 >>
rect 383 383 384 384 
<< m1 >>
rect 384 383 385 384 
<< m1 >>
rect 385 383 386 384 
<< m2 >>
rect 385 383 386 384 
<< m1 >>
rect 386 383 387 384 
<< m2 >>
rect 386 383 387 384 
<< m1 >>
rect 387 383 388 384 
<< m2 >>
rect 387 383 388 384 
<< m1 >>
rect 388 383 389 384 
<< m2 >>
rect 388 383 389 384 
<< m1 >>
rect 389 383 390 384 
<< m2 >>
rect 389 383 390 384 
<< m1 >>
rect 390 383 391 384 
<< m2 >>
rect 390 383 391 384 
<< m1 >>
rect 391 383 392 384 
<< m2 >>
rect 391 383 392 384 
<< m1 >>
rect 392 383 393 384 
<< m2 >>
rect 392 383 393 384 
<< m1 >>
rect 393 383 394 384 
<< m2 >>
rect 393 383 394 384 
<< m1 >>
rect 394 383 395 384 
<< m2 >>
rect 394 383 395 384 
<< m2 >>
rect 395 383 396 384 
<< m1 >>
rect 396 383 397 384 
<< m2 >>
rect 396 383 397 384 
<< m2c >>
rect 396 383 397 384 
<< m1 >>
rect 396 383 397 384 
<< m2 >>
rect 396 383 397 384 
<< m1 >>
rect 397 383 398 384 
<< m1 >>
rect 402 383 403 384 
<< m2 >>
rect 402 383 403 384 
<< m2c >>
rect 402 383 403 384 
<< m1 >>
rect 402 383 403 384 
<< m2 >>
rect 402 383 403 384 
<< m1 >>
rect 406 383 407 384 
<< m2 >>
rect 410 383 411 384 
<< m1 >>
rect 416 383 417 384 
<< m2 >>
rect 429 383 430 384 
<< m1 >>
rect 433 383 434 384 
<< m1 >>
rect 435 383 436 384 
<< m2 >>
rect 439 383 440 384 
<< m2 >>
rect 440 383 441 384 
<< m2 >>
rect 441 383 442 384 
<< m2 >>
rect 442 383 443 384 
<< m2 >>
rect 443 383 444 384 
<< m2 >>
rect 444 383 445 384 
<< m2 >>
rect 445 383 446 384 
<< m2 >>
rect 446 383 447 384 
<< m1 >>
rect 451 383 452 384 
<< m2 >>
rect 455 383 456 384 
<< m2 >>
rect 457 383 458 384 
<< m1 >>
rect 523 383 524 384 
<< m1 >>
rect 13 384 14 385 
<< m1 >>
rect 19 384 20 385 
<< m2 >>
rect 23 384 24 385 
<< m1 >>
rect 31 384 32 385 
<< m2 >>
rect 44 384 45 385 
<< m2 >>
rect 48 384 49 385 
<< m2 >>
rect 63 384 64 385 
<< m2 >>
rect 73 384 74 385 
<< m1 >>
rect 78 384 79 385 
<< m1 >>
rect 82 384 83 385 
<< m2 >>
rect 93 384 94 385 
<< m2 >>
rect 100 384 101 385 
<< m2 >>
rect 110 384 111 385 
<< m2 >>
rect 112 384 113 385 
<< m2 >>
rect 114 384 115 385 
<< m1 >>
rect 118 384 119 385 
<< m2 >>
rect 135 384 136 385 
<< m2 >>
rect 136 384 137 385 
<< m2 >>
rect 137 384 138 385 
<< m2 >>
rect 138 384 139 385 
<< m1 >>
rect 139 384 140 385 
<< m2 >>
rect 139 384 140 385 
<< m2 >>
rect 140 384 141 385 
<< m1 >>
rect 141 384 142 385 
<< m2 >>
rect 141 384 142 385 
<< m2c >>
rect 141 384 142 385 
<< m1 >>
rect 141 384 142 385 
<< m2 >>
rect 141 384 142 385 
<< m1 >>
rect 142 384 143 385 
<< m1 >>
rect 143 384 144 385 
<< m1 >>
rect 144 384 145 385 
<< m1 >>
rect 145 384 146 385 
<< m1 >>
rect 146 384 147 385 
<< m1 >>
rect 147 384 148 385 
<< m1 >>
rect 148 384 149 385 
<< m1 >>
rect 150 384 151 385 
<< m1 >>
rect 163 384 164 385 
<< m2 >>
rect 163 384 164 385 
<< m1 >>
rect 167 384 168 385 
<< m1 >>
rect 169 384 170 385 
<< m1 >>
rect 172 384 173 385 
<< m2 >>
rect 196 384 197 385 
<< m2 >>
rect 199 384 200 385 
<< m2 >>
rect 208 384 209 385 
<< m2 >>
rect 210 384 211 385 
<< m2 >>
rect 211 384 212 385 
<< m2 >>
rect 212 384 213 385 
<< m2 >>
rect 213 384 214 385 
<< m2 >>
rect 214 384 215 385 
<< m2 >>
rect 215 384 216 385 
<< m2 >>
rect 216 384 217 385 
<< m2 >>
rect 217 384 218 385 
<< m2 >>
rect 221 384 222 385 
<< m2 >>
rect 223 384 224 385 
<< m1 >>
rect 235 384 236 385 
<< m2 >>
rect 244 384 245 385 
<< m2 >>
rect 253 384 254 385 
<< m2 >>
rect 255 384 256 385 
<< m2 >>
rect 257 384 258 385 
<< m1 >>
rect 264 384 265 385 
<< m2 >>
rect 264 384 265 385 
<< m2c >>
rect 264 384 265 385 
<< m1 >>
rect 264 384 265 385 
<< m2 >>
rect 264 384 265 385 
<< m1 >>
rect 280 384 281 385 
<< m1 >>
rect 281 384 282 385 
<< m1 >>
rect 282 384 283 385 
<< m1 >>
rect 283 384 284 385 
<< m1 >>
rect 284 384 285 385 
<< m1 >>
rect 285 384 286 385 
<< m1 >>
rect 286 384 287 385 
<< m1 >>
rect 287 384 288 385 
<< m1 >>
rect 288 384 289 385 
<< m1 >>
rect 289 384 290 385 
<< m1 >>
rect 290 384 291 385 
<< m1 >>
rect 291 384 292 385 
<< m1 >>
rect 292 384 293 385 
<< m1 >>
rect 293 384 294 385 
<< m1 >>
rect 294 384 295 385 
<< m1 >>
rect 295 384 296 385 
<< m1 >>
rect 296 384 297 385 
<< m1 >>
rect 297 384 298 385 
<< m1 >>
rect 298 384 299 385 
<< m1 >>
rect 299 384 300 385 
<< m1 >>
rect 300 384 301 385 
<< m1 >>
rect 301 384 302 385 
<< m1 >>
rect 302 384 303 385 
<< m1 >>
rect 303 384 304 385 
<< m1 >>
rect 304 384 305 385 
<< m1 >>
rect 305 384 306 385 
<< m1 >>
rect 306 384 307 385 
<< m1 >>
rect 307 384 308 385 
<< m2 >>
rect 307 384 308 385 
<< m1 >>
rect 308 384 309 385 
<< m1 >>
rect 309 384 310 385 
<< m1 >>
rect 310 384 311 385 
<< m1 >>
rect 311 384 312 385 
<< m1 >>
rect 312 384 313 385 
<< m1 >>
rect 313 384 314 385 
<< m1 >>
rect 314 384 315 385 
<< m2 >>
rect 314 384 315 385 
<< m2c >>
rect 314 384 315 385 
<< m1 >>
rect 314 384 315 385 
<< m2 >>
rect 314 384 315 385 
<< m2 >>
rect 315 384 316 385 
<< m1 >>
rect 316 384 317 385 
<< m2 >>
rect 316 384 317 385 
<< m2 >>
rect 317 384 318 385 
<< m1 >>
rect 318 384 319 385 
<< m2 >>
rect 318 384 319 385 
<< m2c >>
rect 318 384 319 385 
<< m1 >>
rect 318 384 319 385 
<< m2 >>
rect 318 384 319 385 
<< m1 >>
rect 319 384 320 385 
<< m1 >>
rect 320 384 321 385 
<< m1 >>
rect 321 384 322 385 
<< m2 >>
rect 321 384 322 385 
<< m1 >>
rect 322 384 323 385 
<< m1 >>
rect 323 384 324 385 
<< m2 >>
rect 323 384 324 385 
<< m2c >>
rect 323 384 324 385 
<< m1 >>
rect 323 384 324 385 
<< m2 >>
rect 323 384 324 385 
<< m1 >>
rect 325 384 326 385 
<< m2 >>
rect 325 384 326 385 
<< m2c >>
rect 325 384 326 385 
<< m1 >>
rect 325 384 326 385 
<< m2 >>
rect 325 384 326 385 
<< m2 >>
rect 359 384 360 385 
<< m1 >>
rect 363 384 364 385 
<< m2 >>
rect 367 384 368 385 
<< m2 >>
rect 385 384 386 385 
<< m2 >>
rect 402 384 403 385 
<< m1 >>
rect 406 384 407 385 
<< m2 >>
rect 410 384 411 385 
<< m1 >>
rect 416 384 417 385 
<< m2 >>
rect 429 384 430 385 
<< m1 >>
rect 433 384 434 385 
<< m1 >>
rect 435 384 436 385 
<< m1 >>
rect 439 384 440 385 
<< m2 >>
rect 439 384 440 385 
<< m2c >>
rect 439 384 440 385 
<< m1 >>
rect 439 384 440 385 
<< m2 >>
rect 439 384 440 385 
<< m1 >>
rect 451 384 452 385 
<< m1 >>
rect 455 384 456 385 
<< m2 >>
rect 455 384 456 385 
<< m2c >>
rect 455 384 456 385 
<< m1 >>
rect 455 384 456 385 
<< m2 >>
rect 455 384 456 385 
<< m1 >>
rect 456 384 457 385 
<< m1 >>
rect 457 384 458 385 
<< m2 >>
rect 457 384 458 385 
<< m1 >>
rect 458 384 459 385 
<< m1 >>
rect 459 384 460 385 
<< m1 >>
rect 460 384 461 385 
<< m1 >>
rect 461 384 462 385 
<< m1 >>
rect 462 384 463 385 
<< m1 >>
rect 463 384 464 385 
<< m1 >>
rect 464 384 465 385 
<< m1 >>
rect 465 384 466 385 
<< m1 >>
rect 466 384 467 385 
<< m1 >>
rect 467 384 468 385 
<< m1 >>
rect 468 384 469 385 
<< m1 >>
rect 469 384 470 385 
<< m1 >>
rect 470 384 471 385 
<< m1 >>
rect 471 384 472 385 
<< m1 >>
rect 472 384 473 385 
<< m1 >>
rect 523 384 524 385 
<< m1 >>
rect 13 385 14 386 
<< m1 >>
rect 19 385 20 386 
<< m2 >>
rect 20 385 21 386 
<< m1 >>
rect 21 385 22 386 
<< m2 >>
rect 21 385 22 386 
<< m2c >>
rect 21 385 22 386 
<< m1 >>
rect 21 385 22 386 
<< m2 >>
rect 21 385 22 386 
<< m1 >>
rect 22 385 23 386 
<< m1 >>
rect 23 385 24 386 
<< m2 >>
rect 23 385 24 386 
<< m1 >>
rect 24 385 25 386 
<< m1 >>
rect 25 385 26 386 
<< m1 >>
rect 26 385 27 386 
<< m1 >>
rect 27 385 28 386 
<< m1 >>
rect 28 385 29 386 
<< m1 >>
rect 29 385 30 386 
<< m2 >>
rect 29 385 30 386 
<< m2c >>
rect 29 385 30 386 
<< m1 >>
rect 29 385 30 386 
<< m2 >>
rect 29 385 30 386 
<< m2 >>
rect 30 385 31 386 
<< m1 >>
rect 31 385 32 386 
<< m2 >>
rect 31 385 32 386 
<< m2 >>
rect 32 385 33 386 
<< m1 >>
rect 33 385 34 386 
<< m2 >>
rect 33 385 34 386 
<< m2c >>
rect 33 385 34 386 
<< m1 >>
rect 33 385 34 386 
<< m2 >>
rect 33 385 34 386 
<< m1 >>
rect 34 385 35 386 
<< m1 >>
rect 35 385 36 386 
<< m1 >>
rect 36 385 37 386 
<< m1 >>
rect 37 385 38 386 
<< m1 >>
rect 38 385 39 386 
<< m1 >>
rect 39 385 40 386 
<< m1 >>
rect 40 385 41 386 
<< m1 >>
rect 41 385 42 386 
<< m1 >>
rect 42 385 43 386 
<< m1 >>
rect 43 385 44 386 
<< m1 >>
rect 44 385 45 386 
<< m2 >>
rect 44 385 45 386 
<< m1 >>
rect 45 385 46 386 
<< m1 >>
rect 46 385 47 386 
<< m1 >>
rect 47 385 48 386 
<< m1 >>
rect 48 385 49 386 
<< m2 >>
rect 48 385 49 386 
<< m1 >>
rect 49 385 50 386 
<< m1 >>
rect 50 385 51 386 
<< m1 >>
rect 51 385 52 386 
<< m1 >>
rect 52 385 53 386 
<< m1 >>
rect 53 385 54 386 
<< m1 >>
rect 54 385 55 386 
<< m1 >>
rect 55 385 56 386 
<< m1 >>
rect 56 385 57 386 
<< m1 >>
rect 57 385 58 386 
<< m1 >>
rect 58 385 59 386 
<< m1 >>
rect 59 385 60 386 
<< m1 >>
rect 60 385 61 386 
<< m1 >>
rect 61 385 62 386 
<< m1 >>
rect 62 385 63 386 
<< m1 >>
rect 63 385 64 386 
<< m2 >>
rect 63 385 64 386 
<< m1 >>
rect 64 385 65 386 
<< m1 >>
rect 65 385 66 386 
<< m1 >>
rect 66 385 67 386 
<< m1 >>
rect 67 385 68 386 
<< m1 >>
rect 68 385 69 386 
<< m1 >>
rect 69 385 70 386 
<< m1 >>
rect 70 385 71 386 
<< m1 >>
rect 71 385 72 386 
<< m1 >>
rect 72 385 73 386 
<< m1 >>
rect 73 385 74 386 
<< m2 >>
rect 73 385 74 386 
<< m1 >>
rect 74 385 75 386 
<< m1 >>
rect 75 385 76 386 
<< m1 >>
rect 76 385 77 386 
<< m2 >>
rect 76 385 77 386 
<< m2c >>
rect 76 385 77 386 
<< m1 >>
rect 76 385 77 386 
<< m2 >>
rect 76 385 77 386 
<< m2 >>
rect 77 385 78 386 
<< m1 >>
rect 78 385 79 386 
<< m2 >>
rect 78 385 79 386 
<< m2 >>
rect 79 385 80 386 
<< m1 >>
rect 80 385 81 386 
<< m2 >>
rect 80 385 81 386 
<< m2c >>
rect 80 385 81 386 
<< m1 >>
rect 80 385 81 386 
<< m2 >>
rect 80 385 81 386 
<< m2 >>
rect 81 385 82 386 
<< m1 >>
rect 82 385 83 386 
<< m2 >>
rect 82 385 83 386 
<< m2 >>
rect 83 385 84 386 
<< m1 >>
rect 84 385 85 386 
<< m2 >>
rect 84 385 85 386 
<< m2c >>
rect 84 385 85 386 
<< m1 >>
rect 84 385 85 386 
<< m2 >>
rect 84 385 85 386 
<< m1 >>
rect 85 385 86 386 
<< m1 >>
rect 86 385 87 386 
<< m1 >>
rect 87 385 88 386 
<< m1 >>
rect 88 385 89 386 
<< m1 >>
rect 89 385 90 386 
<< m1 >>
rect 90 385 91 386 
<< m1 >>
rect 91 385 92 386 
<< m1 >>
rect 92 385 93 386 
<< m1 >>
rect 93 385 94 386 
<< m2 >>
rect 93 385 94 386 
<< m1 >>
rect 94 385 95 386 
<< m1 >>
rect 95 385 96 386 
<< m1 >>
rect 96 385 97 386 
<< m1 >>
rect 97 385 98 386 
<< m1 >>
rect 98 385 99 386 
<< m1 >>
rect 99 385 100 386 
<< m1 >>
rect 100 385 101 386 
<< m2 >>
rect 100 385 101 386 
<< m1 >>
rect 101 385 102 386 
<< m1 >>
rect 102 385 103 386 
<< m1 >>
rect 103 385 104 386 
<< m1 >>
rect 104 385 105 386 
<< m1 >>
rect 105 385 106 386 
<< m1 >>
rect 106 385 107 386 
<< m1 >>
rect 107 385 108 386 
<< m1 >>
rect 108 385 109 386 
<< m1 >>
rect 109 385 110 386 
<< m1 >>
rect 110 385 111 386 
<< m2 >>
rect 110 385 111 386 
<< m1 >>
rect 111 385 112 386 
<< m1 >>
rect 112 385 113 386 
<< m2 >>
rect 112 385 113 386 
<< m1 >>
rect 113 385 114 386 
<< m1 >>
rect 114 385 115 386 
<< m2 >>
rect 114 385 115 386 
<< m1 >>
rect 115 385 116 386 
<< m1 >>
rect 116 385 117 386 
<< m2 >>
rect 116 385 117 386 
<< m2c >>
rect 116 385 117 386 
<< m1 >>
rect 116 385 117 386 
<< m2 >>
rect 116 385 117 386 
<< m2 >>
rect 117 385 118 386 
<< m1 >>
rect 118 385 119 386 
<< m2 >>
rect 118 385 119 386 
<< m2 >>
rect 119 385 120 386 
<< m1 >>
rect 120 385 121 386 
<< m2 >>
rect 120 385 121 386 
<< m2c >>
rect 120 385 121 386 
<< m1 >>
rect 120 385 121 386 
<< m2 >>
rect 120 385 121 386 
<< m1 >>
rect 121 385 122 386 
<< m1 >>
rect 122 385 123 386 
<< m1 >>
rect 123 385 124 386 
<< m1 >>
rect 124 385 125 386 
<< m1 >>
rect 125 385 126 386 
<< m1 >>
rect 127 385 128 386 
<< m1 >>
rect 128 385 129 386 
<< m1 >>
rect 129 385 130 386 
<< m1 >>
rect 130 385 131 386 
<< m1 >>
rect 131 385 132 386 
<< m1 >>
rect 132 385 133 386 
<< m1 >>
rect 133 385 134 386 
<< m1 >>
rect 134 385 135 386 
<< m1 >>
rect 135 385 136 386 
<< m1 >>
rect 136 385 137 386 
<< m1 >>
rect 137 385 138 386 
<< m1 >>
rect 138 385 139 386 
<< m1 >>
rect 139 385 140 386 
<< m1 >>
rect 150 385 151 386 
<< m1 >>
rect 163 385 164 386 
<< m2 >>
rect 163 385 164 386 
<< m1 >>
rect 167 385 168 386 
<< m1 >>
rect 169 385 170 386 
<< m2 >>
rect 171 385 172 386 
<< m1 >>
rect 172 385 173 386 
<< m2 >>
rect 172 385 173 386 
<< m1 >>
rect 173 385 174 386 
<< m2 >>
rect 173 385 174 386 
<< m1 >>
rect 174 385 175 386 
<< m2 >>
rect 174 385 175 386 
<< m1 >>
rect 175 385 176 386 
<< m2 >>
rect 175 385 176 386 
<< m1 >>
rect 176 385 177 386 
<< m2 >>
rect 176 385 177 386 
<< m1 >>
rect 177 385 178 386 
<< m2 >>
rect 177 385 178 386 
<< m1 >>
rect 178 385 179 386 
<< m2 >>
rect 178 385 179 386 
<< m1 >>
rect 179 385 180 386 
<< m2 >>
rect 179 385 180 386 
<< m1 >>
rect 180 385 181 386 
<< m2 >>
rect 180 385 181 386 
<< m1 >>
rect 181 385 182 386 
<< m2 >>
rect 181 385 182 386 
<< m1 >>
rect 182 385 183 386 
<< m2 >>
rect 182 385 183 386 
<< m1 >>
rect 183 385 184 386 
<< m2 >>
rect 183 385 184 386 
<< m1 >>
rect 184 385 185 386 
<< m2 >>
rect 184 385 185 386 
<< m1 >>
rect 185 385 186 386 
<< m2 >>
rect 185 385 186 386 
<< m1 >>
rect 186 385 187 386 
<< m2 >>
rect 186 385 187 386 
<< m1 >>
rect 187 385 188 386 
<< m2 >>
rect 187 385 188 386 
<< m1 >>
rect 188 385 189 386 
<< m2 >>
rect 188 385 189 386 
<< m1 >>
rect 189 385 190 386 
<< m2 >>
rect 189 385 190 386 
<< m1 >>
rect 190 385 191 386 
<< m2 >>
rect 190 385 191 386 
<< m2 >>
rect 191 385 192 386 
<< m1 >>
rect 192 385 193 386 
<< m2 >>
rect 192 385 193 386 
<< m2c >>
rect 192 385 193 386 
<< m1 >>
rect 192 385 193 386 
<< m2 >>
rect 192 385 193 386 
<< m1 >>
rect 193 385 194 386 
<< m1 >>
rect 194 385 195 386 
<< m1 >>
rect 195 385 196 386 
<< m1 >>
rect 196 385 197 386 
<< m2 >>
rect 196 385 197 386 
<< m1 >>
rect 197 385 198 386 
<< m1 >>
rect 198 385 199 386 
<< m1 >>
rect 199 385 200 386 
<< m2 >>
rect 199 385 200 386 
<< m1 >>
rect 200 385 201 386 
<< m1 >>
rect 201 385 202 386 
<< m1 >>
rect 202 385 203 386 
<< m1 >>
rect 203 385 204 386 
<< m1 >>
rect 204 385 205 386 
<< m1 >>
rect 205 385 206 386 
<< m1 >>
rect 206 385 207 386 
<< m1 >>
rect 207 385 208 386 
<< m1 >>
rect 208 385 209 386 
<< m2 >>
rect 208 385 209 386 
<< m1 >>
rect 209 385 210 386 
<< m1 >>
rect 210 385 211 386 
<< m2 >>
rect 210 385 211 386 
<< m1 >>
rect 211 385 212 386 
<< m1 >>
rect 212 385 213 386 
<< m1 >>
rect 213 385 214 386 
<< m1 >>
rect 214 385 215 386 
<< m1 >>
rect 215 385 216 386 
<< m1 >>
rect 216 385 217 386 
<< m1 >>
rect 217 385 218 386 
<< m1 >>
rect 218 385 219 386 
<< m1 >>
rect 219 385 220 386 
<< m1 >>
rect 220 385 221 386 
<< m1 >>
rect 221 385 222 386 
<< m2 >>
rect 221 385 222 386 
<< m1 >>
rect 222 385 223 386 
<< m1 >>
rect 223 385 224 386 
<< m2 >>
rect 223 385 224 386 
<< m1 >>
rect 224 385 225 386 
<< m1 >>
rect 225 385 226 386 
<< m1 >>
rect 226 385 227 386 
<< m1 >>
rect 227 385 228 386 
<< m1 >>
rect 228 385 229 386 
<< m1 >>
rect 229 385 230 386 
<< m1 >>
rect 230 385 231 386 
<< m1 >>
rect 231 385 232 386 
<< m1 >>
rect 232 385 233 386 
<< m1 >>
rect 233 385 234 386 
<< m2 >>
rect 233 385 234 386 
<< m2c >>
rect 233 385 234 386 
<< m1 >>
rect 233 385 234 386 
<< m2 >>
rect 233 385 234 386 
<< m2 >>
rect 234 385 235 386 
<< m1 >>
rect 235 385 236 386 
<< m2 >>
rect 235 385 236 386 
<< m2 >>
rect 236 385 237 386 
<< m1 >>
rect 237 385 238 386 
<< m2 >>
rect 237 385 238 386 
<< m2c >>
rect 237 385 238 386 
<< m1 >>
rect 237 385 238 386 
<< m2 >>
rect 237 385 238 386 
<< m1 >>
rect 238 385 239 386 
<< m1 >>
rect 239 385 240 386 
<< m1 >>
rect 240 385 241 386 
<< m1 >>
rect 241 385 242 386 
<< m1 >>
rect 242 385 243 386 
<< m1 >>
rect 243 385 244 386 
<< m1 >>
rect 244 385 245 386 
<< m2 >>
rect 244 385 245 386 
<< m1 >>
rect 245 385 246 386 
<< m1 >>
rect 246 385 247 386 
<< m1 >>
rect 247 385 248 386 
<< m1 >>
rect 248 385 249 386 
<< m1 >>
rect 249 385 250 386 
<< m1 >>
rect 250 385 251 386 
<< m1 >>
rect 251 385 252 386 
<< m1 >>
rect 252 385 253 386 
<< m1 >>
rect 253 385 254 386 
<< m2 >>
rect 253 385 254 386 
<< m1 >>
rect 254 385 255 386 
<< m1 >>
rect 255 385 256 386 
<< m2 >>
rect 255 385 256 386 
<< m1 >>
rect 256 385 257 386 
<< m1 >>
rect 257 385 258 386 
<< m2 >>
rect 257 385 258 386 
<< m1 >>
rect 258 385 259 386 
<< m1 >>
rect 259 385 260 386 
<< m1 >>
rect 260 385 261 386 
<< m1 >>
rect 261 385 262 386 
<< m1 >>
rect 262 385 263 386 
<< m1 >>
rect 263 385 264 386 
<< m1 >>
rect 264 385 265 386 
<< m1 >>
rect 280 385 281 386 
<< m2 >>
rect 307 385 308 386 
<< m1 >>
rect 316 385 317 386 
<< m2 >>
rect 321 385 322 386 
<< m1 >>
rect 325 385 326 386 
<< m1 >>
rect 327 385 328 386 
<< m1 >>
rect 328 385 329 386 
<< m1 >>
rect 329 385 330 386 
<< m1 >>
rect 330 385 331 386 
<< m1 >>
rect 331 385 332 386 
<< m1 >>
rect 332 385 333 386 
<< m1 >>
rect 333 385 334 386 
<< m1 >>
rect 334 385 335 386 
<< m1 >>
rect 335 385 336 386 
<< m1 >>
rect 336 385 337 386 
<< m1 >>
rect 337 385 338 386 
<< m1 >>
rect 338 385 339 386 
<< m1 >>
rect 339 385 340 386 
<< m1 >>
rect 340 385 341 386 
<< m1 >>
rect 341 385 342 386 
<< m1 >>
rect 342 385 343 386 
<< m1 >>
rect 343 385 344 386 
<< m1 >>
rect 344 385 345 386 
<< m1 >>
rect 345 385 346 386 
<< m1 >>
rect 346 385 347 386 
<< m1 >>
rect 347 385 348 386 
<< m1 >>
rect 348 385 349 386 
<< m1 >>
rect 349 385 350 386 
<< m1 >>
rect 350 385 351 386 
<< m1 >>
rect 351 385 352 386 
<< m1 >>
rect 352 385 353 386 
<< m1 >>
rect 353 385 354 386 
<< m1 >>
rect 354 385 355 386 
<< m1 >>
rect 355 385 356 386 
<< m1 >>
rect 356 385 357 386 
<< m1 >>
rect 357 385 358 386 
<< m1 >>
rect 358 385 359 386 
<< m1 >>
rect 359 385 360 386 
<< m2 >>
rect 359 385 360 386 
<< m1 >>
rect 360 385 361 386 
<< m1 >>
rect 361 385 362 386 
<< m2 >>
rect 361 385 362 386 
<< m2c >>
rect 361 385 362 386 
<< m1 >>
rect 361 385 362 386 
<< m2 >>
rect 361 385 362 386 
<< m2 >>
rect 362 385 363 386 
<< m1 >>
rect 363 385 364 386 
<< m2 >>
rect 363 385 364 386 
<< m2 >>
rect 364 385 365 386 
<< m1 >>
rect 365 385 366 386 
<< m2 >>
rect 365 385 366 386 
<< m2c >>
rect 365 385 366 386 
<< m1 >>
rect 365 385 366 386 
<< m2 >>
rect 365 385 366 386 
<< m1 >>
rect 366 385 367 386 
<< m1 >>
rect 367 385 368 386 
<< m2 >>
rect 367 385 368 386 
<< m1 >>
rect 368 385 369 386 
<< m1 >>
rect 369 385 370 386 
<< m1 >>
rect 370 385 371 386 
<< m1 >>
rect 371 385 372 386 
<< m1 >>
rect 372 385 373 386 
<< m1 >>
rect 373 385 374 386 
<< m1 >>
rect 374 385 375 386 
<< m1 >>
rect 375 385 376 386 
<< m1 >>
rect 376 385 377 386 
<< m1 >>
rect 377 385 378 386 
<< m1 >>
rect 378 385 379 386 
<< m1 >>
rect 379 385 380 386 
<< m1 >>
rect 380 385 381 386 
<< m1 >>
rect 381 385 382 386 
<< m1 >>
rect 382 385 383 386 
<< m1 >>
rect 383 385 384 386 
<< m1 >>
rect 384 385 385 386 
<< m1 >>
rect 385 385 386 386 
<< m2 >>
rect 385 385 386 386 
<< m1 >>
rect 386 385 387 386 
<< m1 >>
rect 387 385 388 386 
<< m1 >>
rect 388 385 389 386 
<< m1 >>
rect 389 385 390 386 
<< m1 >>
rect 390 385 391 386 
<< m1 >>
rect 391 385 392 386 
<< m1 >>
rect 392 385 393 386 
<< m1 >>
rect 393 385 394 386 
<< m1 >>
rect 394 385 395 386 
<< m1 >>
rect 395 385 396 386 
<< m1 >>
rect 396 385 397 386 
<< m1 >>
rect 397 385 398 386 
<< m1 >>
rect 398 385 399 386 
<< m1 >>
rect 399 385 400 386 
<< m1 >>
rect 400 385 401 386 
<< m1 >>
rect 401 385 402 386 
<< m1 >>
rect 402 385 403 386 
<< m2 >>
rect 402 385 403 386 
<< m1 >>
rect 403 385 404 386 
<< m1 >>
rect 404 385 405 386 
<< m2 >>
rect 404 385 405 386 
<< m2c >>
rect 404 385 405 386 
<< m1 >>
rect 404 385 405 386 
<< m2 >>
rect 404 385 405 386 
<< m2 >>
rect 405 385 406 386 
<< m1 >>
rect 406 385 407 386 
<< m2 >>
rect 406 385 407 386 
<< m2 >>
rect 407 385 408 386 
<< m1 >>
rect 408 385 409 386 
<< m2 >>
rect 408 385 409 386 
<< m2c >>
rect 408 385 409 386 
<< m1 >>
rect 408 385 409 386 
<< m2 >>
rect 408 385 409 386 
<< m1 >>
rect 409 385 410 386 
<< m1 >>
rect 410 385 411 386 
<< m2 >>
rect 410 385 411 386 
<< m1 >>
rect 411 385 412 386 
<< m1 >>
rect 412 385 413 386 
<< m1 >>
rect 413 385 414 386 
<< m1 >>
rect 414 385 415 386 
<< m2 >>
rect 414 385 415 386 
<< m2c >>
rect 414 385 415 386 
<< m1 >>
rect 414 385 415 386 
<< m2 >>
rect 414 385 415 386 
<< m2 >>
rect 415 385 416 386 
<< m1 >>
rect 416 385 417 386 
<< m2 >>
rect 416 385 417 386 
<< m2 >>
rect 417 385 418 386 
<< m1 >>
rect 418 385 419 386 
<< m2 >>
rect 418 385 419 386 
<< m2c >>
rect 418 385 419 386 
<< m1 >>
rect 418 385 419 386 
<< m2 >>
rect 418 385 419 386 
<< m1 >>
rect 419 385 420 386 
<< m1 >>
rect 420 385 421 386 
<< m1 >>
rect 421 385 422 386 
<< m1 >>
rect 422 385 423 386 
<< m1 >>
rect 423 385 424 386 
<< m1 >>
rect 424 385 425 386 
<< m1 >>
rect 425 385 426 386 
<< m1 >>
rect 426 385 427 386 
<< m1 >>
rect 427 385 428 386 
<< m1 >>
rect 428 385 429 386 
<< m1 >>
rect 429 385 430 386 
<< m2 >>
rect 429 385 430 386 
<< m1 >>
rect 430 385 431 386 
<< m1 >>
rect 431 385 432 386 
<< m2 >>
rect 431 385 432 386 
<< m2c >>
rect 431 385 432 386 
<< m1 >>
rect 431 385 432 386 
<< m2 >>
rect 431 385 432 386 
<< m2 >>
rect 432 385 433 386 
<< m1 >>
rect 433 385 434 386 
<< m2 >>
rect 433 385 434 386 
<< m2 >>
rect 434 385 435 386 
<< m1 >>
rect 435 385 436 386 
<< m2 >>
rect 435 385 436 386 
<< m2 >>
rect 436 385 437 386 
<< m1 >>
rect 437 385 438 386 
<< m2 >>
rect 437 385 438 386 
<< m2c >>
rect 437 385 438 386 
<< m1 >>
rect 437 385 438 386 
<< m2 >>
rect 437 385 438 386 
<< m1 >>
rect 438 385 439 386 
<< m1 >>
rect 439 385 440 386 
<< m1 >>
rect 451 385 452 386 
<< m2 >>
rect 457 385 458 386 
<< m2 >>
rect 459 385 460 386 
<< m2 >>
rect 460 385 461 386 
<< m2 >>
rect 461 385 462 386 
<< m2 >>
rect 462 385 463 386 
<< m2 >>
rect 463 385 464 386 
<< m2 >>
rect 464 385 465 386 
<< m2 >>
rect 465 385 466 386 
<< m2 >>
rect 466 385 467 386 
<< m2 >>
rect 467 385 468 386 
<< m2 >>
rect 468 385 469 386 
<< m2 >>
rect 469 385 470 386 
<< m2 >>
rect 470 385 471 386 
<< m2 >>
rect 471 385 472 386 
<< m1 >>
rect 472 385 473 386 
<< m2 >>
rect 472 385 473 386 
<< m2 >>
rect 473 385 474 386 
<< m1 >>
rect 474 385 475 386 
<< m2 >>
rect 474 385 475 386 
<< m2c >>
rect 474 385 475 386 
<< m1 >>
rect 474 385 475 386 
<< m2 >>
rect 474 385 475 386 
<< m1 >>
rect 475 385 476 386 
<< m1 >>
rect 476 385 477 386 
<< m1 >>
rect 523 385 524 386 
<< m1 >>
rect 13 386 14 387 
<< m1 >>
rect 19 386 20 387 
<< m2 >>
rect 20 386 21 387 
<< m2 >>
rect 23 386 24 387 
<< m1 >>
rect 31 386 32 387 
<< m2 >>
rect 44 386 45 387 
<< m2 >>
rect 48 386 49 387 
<< m2 >>
rect 63 386 64 387 
<< m2 >>
rect 73 386 74 387 
<< m1 >>
rect 78 386 79 387 
<< m1 >>
rect 82 386 83 387 
<< m2 >>
rect 93 386 94 387 
<< m2 >>
rect 100 386 101 387 
<< m2 >>
rect 110 386 111 387 
<< m2 >>
rect 112 386 113 387 
<< m2 >>
rect 114 386 115 387 
<< m1 >>
rect 118 386 119 387 
<< m1 >>
rect 125 386 126 387 
<< m1 >>
rect 127 386 128 387 
<< m1 >>
rect 150 386 151 387 
<< m1 >>
rect 163 386 164 387 
<< m2 >>
rect 163 386 164 387 
<< m1 >>
rect 167 386 168 387 
<< m1 >>
rect 169 386 170 387 
<< m2 >>
rect 171 386 172 387 
<< m1 >>
rect 190 386 191 387 
<< m2 >>
rect 196 386 197 387 
<< m2 >>
rect 199 386 200 387 
<< m2 >>
rect 208 386 209 387 
<< m2 >>
rect 210 386 211 387 
<< m2 >>
rect 217 386 218 387 
<< m2 >>
rect 218 386 219 387 
<< m2 >>
rect 219 386 220 387 
<< m2 >>
rect 220 386 221 387 
<< m2 >>
rect 221 386 222 387 
<< m2 >>
rect 223 386 224 387 
<< m1 >>
rect 235 386 236 387 
<< m2 >>
rect 244 386 245 387 
<< m2 >>
rect 253 386 254 387 
<< m2 >>
rect 255 386 256 387 
<< m2 >>
rect 257 386 258 387 
<< m1 >>
rect 280 386 281 387 
<< m1 >>
rect 307 386 308 387 
<< m2 >>
rect 307 386 308 387 
<< m2c >>
rect 307 386 308 387 
<< m1 >>
rect 307 386 308 387 
<< m2 >>
rect 307 386 308 387 
<< m1 >>
rect 316 386 317 387 
<< m1 >>
rect 321 386 322 387 
<< m2 >>
rect 321 386 322 387 
<< m2c >>
rect 321 386 322 387 
<< m1 >>
rect 321 386 322 387 
<< m2 >>
rect 321 386 322 387 
<< m1 >>
rect 322 386 323 387 
<< m1 >>
rect 323 386 324 387 
<< m2 >>
rect 323 386 324 387 
<< m2c >>
rect 323 386 324 387 
<< m1 >>
rect 323 386 324 387 
<< m2 >>
rect 323 386 324 387 
<< m2 >>
rect 324 386 325 387 
<< m1 >>
rect 325 386 326 387 
<< m2 >>
rect 325 386 326 387 
<< m2 >>
rect 326 386 327 387 
<< m1 >>
rect 327 386 328 387 
<< m2 >>
rect 327 386 328 387 
<< m2c >>
rect 327 386 328 387 
<< m1 >>
rect 327 386 328 387 
<< m2 >>
rect 327 386 328 387 
<< m2 >>
rect 359 386 360 387 
<< m1 >>
rect 363 386 364 387 
<< m2 >>
rect 367 386 368 387 
<< m2 >>
rect 385 386 386 387 
<< m2 >>
rect 402 386 403 387 
<< m1 >>
rect 406 386 407 387 
<< m2 >>
rect 410 386 411 387 
<< m1 >>
rect 416 386 417 387 
<< m2 >>
rect 429 386 430 387 
<< m1 >>
rect 433 386 434 387 
<< m1 >>
rect 435 386 436 387 
<< m1 >>
rect 451 386 452 387 
<< m1 >>
rect 457 386 458 387 
<< m2 >>
rect 457 386 458 387 
<< m2c >>
rect 457 386 458 387 
<< m1 >>
rect 457 386 458 387 
<< m2 >>
rect 457 386 458 387 
<< m1 >>
rect 459 386 460 387 
<< m2 >>
rect 459 386 460 387 
<< m2c >>
rect 459 386 460 387 
<< m1 >>
rect 459 386 460 387 
<< m2 >>
rect 459 386 460 387 
<< m1 >>
rect 472 386 473 387 
<< m1 >>
rect 476 386 477 387 
<< m1 >>
rect 523 386 524 387 
<< m1 >>
rect 13 387 14 388 
<< m1 >>
rect 19 387 20 388 
<< m2 >>
rect 20 387 21 388 
<< m1 >>
rect 23 387 24 388 
<< m2 >>
rect 23 387 24 388 
<< m2c >>
rect 23 387 24 388 
<< m1 >>
rect 23 387 24 388 
<< m2 >>
rect 23 387 24 388 
<< m1 >>
rect 31 387 32 388 
<< m1 >>
rect 44 387 45 388 
<< m2 >>
rect 44 387 45 388 
<< m2c >>
rect 44 387 45 388 
<< m1 >>
rect 44 387 45 388 
<< m2 >>
rect 44 387 45 388 
<< m1 >>
rect 46 387 47 388 
<< m1 >>
rect 47 387 48 388 
<< m1 >>
rect 48 387 49 388 
<< m2 >>
rect 48 387 49 388 
<< m2c >>
rect 48 387 49 388 
<< m1 >>
rect 48 387 49 388 
<< m2 >>
rect 48 387 49 388 
<< m2 >>
rect 63 387 64 388 
<< m1 >>
rect 73 387 74 388 
<< m2 >>
rect 73 387 74 388 
<< m2c >>
rect 73 387 74 388 
<< m1 >>
rect 73 387 74 388 
<< m2 >>
rect 73 387 74 388 
<< m1 >>
rect 78 387 79 388 
<< m1 >>
rect 82 387 83 388 
<< m1 >>
rect 93 387 94 388 
<< m2 >>
rect 93 387 94 388 
<< m2c >>
rect 93 387 94 388 
<< m1 >>
rect 93 387 94 388 
<< m2 >>
rect 93 387 94 388 
<< m1 >>
rect 100 387 101 388 
<< m2 >>
rect 100 387 101 388 
<< m2c >>
rect 100 387 101 388 
<< m1 >>
rect 100 387 101 388 
<< m2 >>
rect 100 387 101 388 
<< m1 >>
rect 110 387 111 388 
<< m2 >>
rect 110 387 111 388 
<< m2c >>
rect 110 387 111 388 
<< m1 >>
rect 110 387 111 388 
<< m2 >>
rect 110 387 111 388 
<< m1 >>
rect 112 387 113 388 
<< m2 >>
rect 112 387 113 388 
<< m2c >>
rect 112 387 113 388 
<< m1 >>
rect 112 387 113 388 
<< m2 >>
rect 112 387 113 388 
<< m1 >>
rect 114 387 115 388 
<< m2 >>
rect 114 387 115 388 
<< m2c >>
rect 114 387 115 388 
<< m1 >>
rect 114 387 115 388 
<< m2 >>
rect 114 387 115 388 
<< m1 >>
rect 118 387 119 388 
<< m1 >>
rect 125 387 126 388 
<< m1 >>
rect 127 387 128 388 
<< m1 >>
rect 150 387 151 388 
<< m1 >>
rect 163 387 164 388 
<< m2 >>
rect 163 387 164 388 
<< m1 >>
rect 167 387 168 388 
<< m1 >>
rect 169 387 170 388 
<< m1 >>
rect 171 387 172 388 
<< m2 >>
rect 171 387 172 388 
<< m2c >>
rect 171 387 172 388 
<< m1 >>
rect 171 387 172 388 
<< m2 >>
rect 171 387 172 388 
<< m1 >>
rect 190 387 191 388 
<< m1 >>
rect 196 387 197 388 
<< m2 >>
rect 196 387 197 388 
<< m2c >>
rect 196 387 197 388 
<< m1 >>
rect 196 387 197 388 
<< m2 >>
rect 196 387 197 388 
<< m1 >>
rect 199 387 200 388 
<< m2 >>
rect 199 387 200 388 
<< m2c >>
rect 199 387 200 388 
<< m1 >>
rect 199 387 200 388 
<< m2 >>
rect 199 387 200 388 
<< m1 >>
rect 206 387 207 388 
<< m1 >>
rect 207 387 208 388 
<< m1 >>
rect 208 387 209 388 
<< m2 >>
rect 208 387 209 388 
<< m1 >>
rect 209 387 210 388 
<< m1 >>
rect 210 387 211 388 
<< m2 >>
rect 210 387 211 388 
<< m2c >>
rect 210 387 211 388 
<< m1 >>
rect 210 387 211 388 
<< m2 >>
rect 210 387 211 388 
<< m1 >>
rect 217 387 218 388 
<< m2 >>
rect 217 387 218 388 
<< m2c >>
rect 217 387 218 388 
<< m1 >>
rect 217 387 218 388 
<< m2 >>
rect 217 387 218 388 
<< m1 >>
rect 223 387 224 388 
<< m2 >>
rect 223 387 224 388 
<< m2c >>
rect 223 387 224 388 
<< m1 >>
rect 223 387 224 388 
<< m2 >>
rect 223 387 224 388 
<< m1 >>
rect 235 387 236 388 
<< m1 >>
rect 244 387 245 388 
<< m2 >>
rect 244 387 245 388 
<< m2c >>
rect 244 387 245 388 
<< m1 >>
rect 244 387 245 388 
<< m2 >>
rect 244 387 245 388 
<< m1 >>
rect 253 387 254 388 
<< m2 >>
rect 253 387 254 388 
<< m2c >>
rect 253 387 254 388 
<< m1 >>
rect 253 387 254 388 
<< m2 >>
rect 253 387 254 388 
<< m1 >>
rect 255 387 256 388 
<< m2 >>
rect 255 387 256 388 
<< m2c >>
rect 255 387 256 388 
<< m1 >>
rect 255 387 256 388 
<< m2 >>
rect 255 387 256 388 
<< m1 >>
rect 257 387 258 388 
<< m2 >>
rect 257 387 258 388 
<< m2c >>
rect 257 387 258 388 
<< m1 >>
rect 257 387 258 388 
<< m2 >>
rect 257 387 258 388 
<< m1 >>
rect 258 387 259 388 
<< m1 >>
rect 259 387 260 388 
<< m1 >>
rect 280 387 281 388 
<< m1 >>
rect 307 387 308 388 
<< m1 >>
rect 316 387 317 388 
<< m1 >>
rect 325 387 326 388 
<< m1 >>
rect 337 387 338 388 
<< m1 >>
rect 338 387 339 388 
<< m1 >>
rect 339 387 340 388 
<< m1 >>
rect 340 387 341 388 
<< m1 >>
rect 341 387 342 388 
<< m1 >>
rect 342 387 343 388 
<< m1 >>
rect 343 387 344 388 
<< m1 >>
rect 355 387 356 388 
<< m1 >>
rect 356 387 357 388 
<< m1 >>
rect 357 387 358 388 
<< m1 >>
rect 358 387 359 388 
<< m1 >>
rect 359 387 360 388 
<< m2 >>
rect 359 387 360 388 
<< m1 >>
rect 360 387 361 388 
<< m1 >>
rect 361 387 362 388 
<< m1 >>
rect 363 387 364 388 
<< m1 >>
rect 367 387 368 388 
<< m2 >>
rect 367 387 368 388 
<< m2c >>
rect 367 387 368 388 
<< m1 >>
rect 367 387 368 388 
<< m2 >>
rect 367 387 368 388 
<< m1 >>
rect 385 387 386 388 
<< m2 >>
rect 385 387 386 388 
<< m2c >>
rect 385 387 386 388 
<< m1 >>
rect 385 387 386 388 
<< m2 >>
rect 385 387 386 388 
<< m1 >>
rect 402 387 403 388 
<< m2 >>
rect 402 387 403 388 
<< m2c >>
rect 402 387 403 388 
<< m1 >>
rect 402 387 403 388 
<< m2 >>
rect 402 387 403 388 
<< m1 >>
rect 406 387 407 388 
<< m1 >>
rect 410 387 411 388 
<< m2 >>
rect 410 387 411 388 
<< m2c >>
rect 410 387 411 388 
<< m1 >>
rect 410 387 411 388 
<< m2 >>
rect 410 387 411 388 
<< m1 >>
rect 411 387 412 388 
<< m1 >>
rect 412 387 413 388 
<< m1 >>
rect 413 387 414 388 
<< m1 >>
rect 414 387 415 388 
<< m2 >>
rect 414 387 415 388 
<< m2c >>
rect 414 387 415 388 
<< m1 >>
rect 414 387 415 388 
<< m2 >>
rect 414 387 415 388 
<< m2 >>
rect 415 387 416 388 
<< m1 >>
rect 416 387 417 388 
<< m2 >>
rect 416 387 417 388 
<< m2 >>
rect 417 387 418 388 
<< m1 >>
rect 418 387 419 388 
<< m2 >>
rect 418 387 419 388 
<< m2c >>
rect 418 387 419 388 
<< m1 >>
rect 418 387 419 388 
<< m2 >>
rect 418 387 419 388 
<< m1 >>
rect 429 387 430 388 
<< m2 >>
rect 429 387 430 388 
<< m2c >>
rect 429 387 430 388 
<< m1 >>
rect 429 387 430 388 
<< m2 >>
rect 429 387 430 388 
<< m1 >>
rect 430 387 431 388 
<< m1 >>
rect 431 387 432 388 
<< m2 >>
rect 431 387 432 388 
<< m2c >>
rect 431 387 432 388 
<< m1 >>
rect 431 387 432 388 
<< m2 >>
rect 431 387 432 388 
<< m2 >>
rect 432 387 433 388 
<< m1 >>
rect 433 387 434 388 
<< m2 >>
rect 433 387 434 388 
<< m2 >>
rect 434 387 435 388 
<< m1 >>
rect 435 387 436 388 
<< m2 >>
rect 435 387 436 388 
<< m2 >>
rect 436 387 437 388 
<< m1 >>
rect 437 387 438 388 
<< m2 >>
rect 437 387 438 388 
<< m2c >>
rect 437 387 438 388 
<< m1 >>
rect 437 387 438 388 
<< m2 >>
rect 437 387 438 388 
<< m1 >>
rect 451 387 452 388 
<< m1 >>
rect 457 387 458 388 
<< m1 >>
rect 459 387 460 388 
<< m1 >>
rect 472 387 473 388 
<< m1 >>
rect 476 387 477 388 
<< m1 >>
rect 523 387 524 388 
<< m1 >>
rect 13 388 14 389 
<< m1 >>
rect 19 388 20 389 
<< m2 >>
rect 20 388 21 389 
<< m1 >>
rect 23 388 24 389 
<< m1 >>
rect 31 388 32 389 
<< m1 >>
rect 44 388 45 389 
<< m1 >>
rect 46 388 47 389 
<< m2 >>
rect 63 388 64 389 
<< m1 >>
rect 64 388 65 389 
<< m1 >>
rect 65 388 66 389 
<< m1 >>
rect 66 388 67 389 
<< m1 >>
rect 67 388 68 389 
<< m1 >>
rect 73 388 74 389 
<< m1 >>
rect 78 388 79 389 
<< m1 >>
rect 82 388 83 389 
<< m1 >>
rect 93 388 94 389 
<< m1 >>
rect 100 388 101 389 
<< m1 >>
rect 110 388 111 389 
<< m1 >>
rect 112 388 113 389 
<< m1 >>
rect 114 388 115 389 
<< m1 >>
rect 118 388 119 389 
<< m1 >>
rect 125 388 126 389 
<< m2 >>
rect 125 388 126 389 
<< m2c >>
rect 125 388 126 389 
<< m1 >>
rect 125 388 126 389 
<< m2 >>
rect 125 388 126 389 
<< m2 >>
rect 126 388 127 389 
<< m1 >>
rect 127 388 128 389 
<< m2 >>
rect 127 388 128 389 
<< m2 >>
rect 128 388 129 389 
<< m1 >>
rect 136 388 137 389 
<< m1 >>
rect 137 388 138 389 
<< m1 >>
rect 138 388 139 389 
<< m1 >>
rect 139 388 140 389 
<< m1 >>
rect 150 388 151 389 
<< m1 >>
rect 160 388 161 389 
<< m1 >>
rect 161 388 162 389 
<< m2 >>
rect 161 388 162 389 
<< m2c >>
rect 161 388 162 389 
<< m1 >>
rect 161 388 162 389 
<< m2 >>
rect 161 388 162 389 
<< m2 >>
rect 162 388 163 389 
<< m1 >>
rect 163 388 164 389 
<< m2 >>
rect 163 388 164 389 
<< m1 >>
rect 167 388 168 389 
<< m1 >>
rect 169 388 170 389 
<< m1 >>
rect 171 388 172 389 
<< m1 >>
rect 190 388 191 389 
<< m1 >>
rect 196 388 197 389 
<< m1 >>
rect 199 388 200 389 
<< m2 >>
rect 205 388 206 389 
<< m1 >>
rect 206 388 207 389 
<< m2 >>
rect 206 388 207 389 
<< m2 >>
rect 207 388 208 389 
<< m2 >>
rect 208 388 209 389 
<< m1 >>
rect 217 388 218 389 
<< m1 >>
rect 223 388 224 389 
<< m1 >>
rect 235 388 236 389 
<< m1 >>
rect 244 388 245 389 
<< m1 >>
rect 253 388 254 389 
<< m1 >>
rect 255 388 256 389 
<< m1 >>
rect 259 388 260 389 
<< m1 >>
rect 280 388 281 389 
<< m1 >>
rect 307 388 308 389 
<< m1 >>
rect 310 388 311 389 
<< m1 >>
rect 311 388 312 389 
<< m1 >>
rect 312 388 313 389 
<< m1 >>
rect 313 388 314 389 
<< m1 >>
rect 314 388 315 389 
<< m2 >>
rect 314 388 315 389 
<< m2c >>
rect 314 388 315 389 
<< m1 >>
rect 314 388 315 389 
<< m2 >>
rect 314 388 315 389 
<< m2 >>
rect 315 388 316 389 
<< m1 >>
rect 316 388 317 389 
<< m2 >>
rect 316 388 317 389 
<< m2 >>
rect 317 388 318 389 
<< m1 >>
rect 318 388 319 389 
<< m2 >>
rect 318 388 319 389 
<< m2c >>
rect 318 388 319 389 
<< m1 >>
rect 318 388 319 389 
<< m2 >>
rect 318 388 319 389 
<< m1 >>
rect 319 388 320 389 
<< m1 >>
rect 325 388 326 389 
<< m1 >>
rect 337 388 338 389 
<< m1 >>
rect 343 388 344 389 
<< m1 >>
rect 355 388 356 389 
<< m2 >>
rect 359 388 360 389 
<< m2 >>
rect 360 388 361 389 
<< m1 >>
rect 361 388 362 389 
<< m2 >>
rect 361 388 362 389 
<< m2 >>
rect 362 388 363 389 
<< m1 >>
rect 363 388 364 389 
<< m2 >>
rect 363 388 364 389 
<< m2 >>
rect 364 388 365 389 
<< m1 >>
rect 367 388 368 389 
<< m1 >>
rect 385 388 386 389 
<< m1 >>
rect 402 388 403 389 
<< m1 >>
rect 406 388 407 389 
<< m1 >>
rect 416 388 417 389 
<< m1 >>
rect 418 388 419 389 
<< m1 >>
rect 433 388 434 389 
<< m1 >>
rect 435 388 436 389 
<< m1 >>
rect 437 388 438 389 
<< m1 >>
rect 451 388 452 389 
<< m1 >>
rect 457 388 458 389 
<< m1 >>
rect 459 388 460 389 
<< m1 >>
rect 472 388 473 389 
<< m1 >>
rect 476 388 477 389 
<< m1 >>
rect 478 388 479 389 
<< m1 >>
rect 479 388 480 389 
<< m1 >>
rect 480 388 481 389 
<< m1 >>
rect 481 388 482 389 
<< m1 >>
rect 523 388 524 389 
<< m1 >>
rect 13 389 14 390 
<< m1 >>
rect 19 389 20 390 
<< m2 >>
rect 20 389 21 390 
<< m1 >>
rect 23 389 24 390 
<< m1 >>
rect 31 389 32 390 
<< m1 >>
rect 42 389 43 390 
<< m2 >>
rect 42 389 43 390 
<< m2c >>
rect 42 389 43 390 
<< m1 >>
rect 42 389 43 390 
<< m2 >>
rect 42 389 43 390 
<< m2 >>
rect 43 389 44 390 
<< m1 >>
rect 44 389 45 390 
<< m2 >>
rect 44 389 45 390 
<< m2 >>
rect 45 389 46 390 
<< m1 >>
rect 46 389 47 390 
<< m2 >>
rect 46 389 47 390 
<< m2c >>
rect 46 389 47 390 
<< m1 >>
rect 46 389 47 390 
<< m2 >>
rect 46 389 47 390 
<< m2 >>
rect 63 389 64 390 
<< m1 >>
rect 64 389 65 390 
<< m1 >>
rect 67 389 68 390 
<< m1 >>
rect 73 389 74 390 
<< m1 >>
rect 78 389 79 390 
<< m1 >>
rect 82 389 83 390 
<< m1 >>
rect 93 389 94 390 
<< m1 >>
rect 100 389 101 390 
<< m1 >>
rect 110 389 111 390 
<< m1 >>
rect 112 389 113 390 
<< m1 >>
rect 114 389 115 390 
<< m1 >>
rect 118 389 119 390 
<< m1 >>
rect 127 389 128 390 
<< m2 >>
rect 128 389 129 390 
<< m1 >>
rect 136 389 137 390 
<< m1 >>
rect 139 389 140 390 
<< m1 >>
rect 150 389 151 390 
<< m1 >>
rect 160 389 161 390 
<< m1 >>
rect 163 389 164 390 
<< m1 >>
rect 167 389 168 390 
<< m1 >>
rect 169 389 170 390 
<< m1 >>
rect 171 389 172 390 
<< m1 >>
rect 190 389 191 390 
<< m1 >>
rect 196 389 197 390 
<< m1 >>
rect 199 389 200 390 
<< m2 >>
rect 205 389 206 390 
<< m1 >>
rect 206 389 207 390 
<< m1 >>
rect 217 389 218 390 
<< m1 >>
rect 223 389 224 390 
<< m1 >>
rect 235 389 236 390 
<< m1 >>
rect 244 389 245 390 
<< m1 >>
rect 253 389 254 390 
<< m1 >>
rect 255 389 256 390 
<< m1 >>
rect 259 389 260 390 
<< m1 >>
rect 280 389 281 390 
<< m1 >>
rect 307 389 308 390 
<< m1 >>
rect 310 389 311 390 
<< m1 >>
rect 316 389 317 390 
<< m1 >>
rect 319 389 320 390 
<< m1 >>
rect 325 389 326 390 
<< m1 >>
rect 337 389 338 390 
<< m1 >>
rect 343 389 344 390 
<< m1 >>
rect 355 389 356 390 
<< m1 >>
rect 361 389 362 390 
<< m1 >>
rect 363 389 364 390 
<< m2 >>
rect 364 389 365 390 
<< m1 >>
rect 367 389 368 390 
<< m1 >>
rect 385 389 386 390 
<< m1 >>
rect 402 389 403 390 
<< m1 >>
rect 406 389 407 390 
<< m1 >>
rect 416 389 417 390 
<< m1 >>
rect 418 389 419 390 
<< m1 >>
rect 433 389 434 390 
<< m1 >>
rect 435 389 436 390 
<< m1 >>
rect 437 389 438 390 
<< m1 >>
rect 451 389 452 390 
<< m1 >>
rect 457 389 458 390 
<< m1 >>
rect 459 389 460 390 
<< m1 >>
rect 472 389 473 390 
<< m1 >>
rect 476 389 477 390 
<< m1 >>
rect 478 389 479 390 
<< m1 >>
rect 481 389 482 390 
<< m1 >>
rect 523 389 524 390 
<< pdiffusion >>
rect 12 390 13 391 
<< m1 >>
rect 13 390 14 391 
<< pdiffusion >>
rect 13 390 14 391 
<< pdiffusion >>
rect 14 390 15 391 
<< pdiffusion >>
rect 15 390 16 391 
<< pdiffusion >>
rect 16 390 17 391 
<< pdiffusion >>
rect 17 390 18 391 
<< m1 >>
rect 19 390 20 391 
<< m2 >>
rect 20 390 21 391 
<< m1 >>
rect 23 390 24 391 
<< pdiffusion >>
rect 30 390 31 391 
<< m1 >>
rect 31 390 32 391 
<< pdiffusion >>
rect 31 390 32 391 
<< pdiffusion >>
rect 32 390 33 391 
<< pdiffusion >>
rect 33 390 34 391 
<< pdiffusion >>
rect 34 390 35 391 
<< pdiffusion >>
rect 35 390 36 391 
<< m1 >>
rect 42 390 43 391 
<< m1 >>
rect 44 390 45 391 
<< pdiffusion >>
rect 48 390 49 391 
<< pdiffusion >>
rect 49 390 50 391 
<< pdiffusion >>
rect 50 390 51 391 
<< pdiffusion >>
rect 51 390 52 391 
<< pdiffusion >>
rect 52 390 53 391 
<< pdiffusion >>
rect 53 390 54 391 
<< m2 >>
rect 63 390 64 391 
<< m1 >>
rect 64 390 65 391 
<< pdiffusion >>
rect 66 390 67 391 
<< m1 >>
rect 67 390 68 391 
<< pdiffusion >>
rect 67 390 68 391 
<< pdiffusion >>
rect 68 390 69 391 
<< pdiffusion >>
rect 69 390 70 391 
<< pdiffusion >>
rect 70 390 71 391 
<< pdiffusion >>
rect 71 390 72 391 
<< m1 >>
rect 73 390 74 391 
<< m1 >>
rect 78 390 79 391 
<< m1 >>
rect 82 390 83 391 
<< pdiffusion >>
rect 84 390 85 391 
<< pdiffusion >>
rect 85 390 86 391 
<< pdiffusion >>
rect 86 390 87 391 
<< pdiffusion >>
rect 87 390 88 391 
<< pdiffusion >>
rect 88 390 89 391 
<< pdiffusion >>
rect 89 390 90 391 
<< m1 >>
rect 93 390 94 391 
<< m1 >>
rect 100 390 101 391 
<< pdiffusion >>
rect 102 390 103 391 
<< pdiffusion >>
rect 103 390 104 391 
<< pdiffusion >>
rect 104 390 105 391 
<< pdiffusion >>
rect 105 390 106 391 
<< pdiffusion >>
rect 106 390 107 391 
<< pdiffusion >>
rect 107 390 108 391 
<< m1 >>
rect 110 390 111 391 
<< m1 >>
rect 112 390 113 391 
<< m1 >>
rect 114 390 115 391 
<< m1 >>
rect 118 390 119 391 
<< pdiffusion >>
rect 120 390 121 391 
<< pdiffusion >>
rect 121 390 122 391 
<< pdiffusion >>
rect 122 390 123 391 
<< pdiffusion >>
rect 123 390 124 391 
<< pdiffusion >>
rect 124 390 125 391 
<< pdiffusion >>
rect 125 390 126 391 
<< m1 >>
rect 127 390 128 391 
<< m2 >>
rect 128 390 129 391 
<< m1 >>
rect 136 390 137 391 
<< pdiffusion >>
rect 138 390 139 391 
<< m1 >>
rect 139 390 140 391 
<< pdiffusion >>
rect 139 390 140 391 
<< pdiffusion >>
rect 140 390 141 391 
<< pdiffusion >>
rect 141 390 142 391 
<< pdiffusion >>
rect 142 390 143 391 
<< pdiffusion >>
rect 143 390 144 391 
<< m1 >>
rect 150 390 151 391 
<< pdiffusion >>
rect 156 390 157 391 
<< pdiffusion >>
rect 157 390 158 391 
<< pdiffusion >>
rect 158 390 159 391 
<< pdiffusion >>
rect 159 390 160 391 
<< m1 >>
rect 160 390 161 391 
<< pdiffusion >>
rect 160 390 161 391 
<< pdiffusion >>
rect 161 390 162 391 
<< m1 >>
rect 163 390 164 391 
<< m1 >>
rect 167 390 168 391 
<< m1 >>
rect 169 390 170 391 
<< m1 >>
rect 171 390 172 391 
<< pdiffusion >>
rect 174 390 175 391 
<< pdiffusion >>
rect 175 390 176 391 
<< pdiffusion >>
rect 176 390 177 391 
<< pdiffusion >>
rect 177 390 178 391 
<< pdiffusion >>
rect 178 390 179 391 
<< pdiffusion >>
rect 179 390 180 391 
<< m1 >>
rect 190 390 191 391 
<< pdiffusion >>
rect 192 390 193 391 
<< pdiffusion >>
rect 193 390 194 391 
<< pdiffusion >>
rect 194 390 195 391 
<< pdiffusion >>
rect 195 390 196 391 
<< m1 >>
rect 196 390 197 391 
<< pdiffusion >>
rect 196 390 197 391 
<< pdiffusion >>
rect 197 390 198 391 
<< m1 >>
rect 199 390 200 391 
<< m2 >>
rect 205 390 206 391 
<< m1 >>
rect 206 390 207 391 
<< pdiffusion >>
rect 210 390 211 391 
<< pdiffusion >>
rect 211 390 212 391 
<< pdiffusion >>
rect 212 390 213 391 
<< pdiffusion >>
rect 213 390 214 391 
<< pdiffusion >>
rect 214 390 215 391 
<< pdiffusion >>
rect 215 390 216 391 
<< m1 >>
rect 217 390 218 391 
<< m1 >>
rect 223 390 224 391 
<< pdiffusion >>
rect 228 390 229 391 
<< pdiffusion >>
rect 229 390 230 391 
<< pdiffusion >>
rect 230 390 231 391 
<< pdiffusion >>
rect 231 390 232 391 
<< pdiffusion >>
rect 232 390 233 391 
<< pdiffusion >>
rect 233 390 234 391 
<< m1 >>
rect 235 390 236 391 
<< m1 >>
rect 244 390 245 391 
<< pdiffusion >>
rect 246 390 247 391 
<< pdiffusion >>
rect 247 390 248 391 
<< pdiffusion >>
rect 248 390 249 391 
<< pdiffusion >>
rect 249 390 250 391 
<< pdiffusion >>
rect 250 390 251 391 
<< pdiffusion >>
rect 251 390 252 391 
<< m1 >>
rect 253 390 254 391 
<< m1 >>
rect 255 390 256 391 
<< m1 >>
rect 259 390 260 391 
<< pdiffusion >>
rect 264 390 265 391 
<< pdiffusion >>
rect 265 390 266 391 
<< pdiffusion >>
rect 266 390 267 391 
<< pdiffusion >>
rect 267 390 268 391 
<< pdiffusion >>
rect 268 390 269 391 
<< pdiffusion >>
rect 269 390 270 391 
<< m1 >>
rect 280 390 281 391 
<< pdiffusion >>
rect 282 390 283 391 
<< pdiffusion >>
rect 283 390 284 391 
<< pdiffusion >>
rect 284 390 285 391 
<< pdiffusion >>
rect 285 390 286 391 
<< pdiffusion >>
rect 286 390 287 391 
<< pdiffusion >>
rect 287 390 288 391 
<< pdiffusion >>
rect 300 390 301 391 
<< pdiffusion >>
rect 301 390 302 391 
<< pdiffusion >>
rect 302 390 303 391 
<< pdiffusion >>
rect 303 390 304 391 
<< pdiffusion >>
rect 304 390 305 391 
<< pdiffusion >>
rect 305 390 306 391 
<< m1 >>
rect 307 390 308 391 
<< m1 >>
rect 310 390 311 391 
<< m1 >>
rect 316 390 317 391 
<< pdiffusion >>
rect 318 390 319 391 
<< m1 >>
rect 319 390 320 391 
<< pdiffusion >>
rect 319 390 320 391 
<< pdiffusion >>
rect 320 390 321 391 
<< pdiffusion >>
rect 321 390 322 391 
<< pdiffusion >>
rect 322 390 323 391 
<< pdiffusion >>
rect 323 390 324 391 
<< m1 >>
rect 325 390 326 391 
<< pdiffusion >>
rect 336 390 337 391 
<< m1 >>
rect 337 390 338 391 
<< pdiffusion >>
rect 337 390 338 391 
<< pdiffusion >>
rect 338 390 339 391 
<< pdiffusion >>
rect 339 390 340 391 
<< pdiffusion >>
rect 340 390 341 391 
<< pdiffusion >>
rect 341 390 342 391 
<< m1 >>
rect 343 390 344 391 
<< pdiffusion >>
rect 354 390 355 391 
<< m1 >>
rect 355 390 356 391 
<< pdiffusion >>
rect 355 390 356 391 
<< pdiffusion >>
rect 356 390 357 391 
<< pdiffusion >>
rect 357 390 358 391 
<< pdiffusion >>
rect 358 390 359 391 
<< pdiffusion >>
rect 359 390 360 391 
<< m1 >>
rect 361 390 362 391 
<< m1 >>
rect 363 390 364 391 
<< m2 >>
rect 364 390 365 391 
<< m1 >>
rect 367 390 368 391 
<< pdiffusion >>
rect 372 390 373 391 
<< pdiffusion >>
rect 373 390 374 391 
<< pdiffusion >>
rect 374 390 375 391 
<< pdiffusion >>
rect 375 390 376 391 
<< pdiffusion >>
rect 376 390 377 391 
<< pdiffusion >>
rect 377 390 378 391 
<< m1 >>
rect 385 390 386 391 
<< m1 >>
rect 402 390 403 391 
<< m1 >>
rect 406 390 407 391 
<< pdiffusion >>
rect 408 390 409 391 
<< pdiffusion >>
rect 409 390 410 391 
<< pdiffusion >>
rect 410 390 411 391 
<< pdiffusion >>
rect 411 390 412 391 
<< pdiffusion >>
rect 412 390 413 391 
<< pdiffusion >>
rect 413 390 414 391 
<< m1 >>
rect 416 390 417 391 
<< m1 >>
rect 418 390 419 391 
<< pdiffusion >>
rect 426 390 427 391 
<< pdiffusion >>
rect 427 390 428 391 
<< pdiffusion >>
rect 428 390 429 391 
<< pdiffusion >>
rect 429 390 430 391 
<< pdiffusion >>
rect 430 390 431 391 
<< pdiffusion >>
rect 431 390 432 391 
<< m1 >>
rect 433 390 434 391 
<< m1 >>
rect 435 390 436 391 
<< m1 >>
rect 437 390 438 391 
<< pdiffusion >>
rect 444 390 445 391 
<< pdiffusion >>
rect 445 390 446 391 
<< pdiffusion >>
rect 446 390 447 391 
<< pdiffusion >>
rect 447 390 448 391 
<< pdiffusion >>
rect 448 390 449 391 
<< pdiffusion >>
rect 449 390 450 391 
<< m1 >>
rect 451 390 452 391 
<< m1 >>
rect 457 390 458 391 
<< m1 >>
rect 459 390 460 391 
<< pdiffusion >>
rect 462 390 463 391 
<< pdiffusion >>
rect 463 390 464 391 
<< pdiffusion >>
rect 464 390 465 391 
<< pdiffusion >>
rect 465 390 466 391 
<< pdiffusion >>
rect 466 390 467 391 
<< pdiffusion >>
rect 467 390 468 391 
<< m1 >>
rect 472 390 473 391 
<< m1 >>
rect 476 390 477 391 
<< m1 >>
rect 478 390 479 391 
<< pdiffusion >>
rect 480 390 481 391 
<< m1 >>
rect 481 390 482 391 
<< pdiffusion >>
rect 481 390 482 391 
<< pdiffusion >>
rect 482 390 483 391 
<< pdiffusion >>
rect 483 390 484 391 
<< pdiffusion >>
rect 484 390 485 391 
<< pdiffusion >>
rect 485 390 486 391 
<< pdiffusion >>
rect 498 390 499 391 
<< pdiffusion >>
rect 499 390 500 391 
<< pdiffusion >>
rect 500 390 501 391 
<< pdiffusion >>
rect 501 390 502 391 
<< pdiffusion >>
rect 502 390 503 391 
<< pdiffusion >>
rect 503 390 504 391 
<< pdiffusion >>
rect 516 390 517 391 
<< pdiffusion >>
rect 517 390 518 391 
<< pdiffusion >>
rect 518 390 519 391 
<< pdiffusion >>
rect 519 390 520 391 
<< pdiffusion >>
rect 520 390 521 391 
<< pdiffusion >>
rect 521 390 522 391 
<< m1 >>
rect 523 390 524 391 
<< pdiffusion >>
rect 12 391 13 392 
<< pdiffusion >>
rect 13 391 14 392 
<< pdiffusion >>
rect 14 391 15 392 
<< pdiffusion >>
rect 15 391 16 392 
<< pdiffusion >>
rect 16 391 17 392 
<< pdiffusion >>
rect 17 391 18 392 
<< m1 >>
rect 19 391 20 392 
<< m2 >>
rect 20 391 21 392 
<< m1 >>
rect 23 391 24 392 
<< pdiffusion >>
rect 30 391 31 392 
<< pdiffusion >>
rect 31 391 32 392 
<< pdiffusion >>
rect 32 391 33 392 
<< pdiffusion >>
rect 33 391 34 392 
<< pdiffusion >>
rect 34 391 35 392 
<< pdiffusion >>
rect 35 391 36 392 
<< m1 >>
rect 42 391 43 392 
<< m1 >>
rect 44 391 45 392 
<< pdiffusion >>
rect 48 391 49 392 
<< pdiffusion >>
rect 49 391 50 392 
<< pdiffusion >>
rect 50 391 51 392 
<< pdiffusion >>
rect 51 391 52 392 
<< pdiffusion >>
rect 52 391 53 392 
<< pdiffusion >>
rect 53 391 54 392 
<< m2 >>
rect 63 391 64 392 
<< m1 >>
rect 64 391 65 392 
<< pdiffusion >>
rect 66 391 67 392 
<< pdiffusion >>
rect 67 391 68 392 
<< pdiffusion >>
rect 68 391 69 392 
<< pdiffusion >>
rect 69 391 70 392 
<< pdiffusion >>
rect 70 391 71 392 
<< pdiffusion >>
rect 71 391 72 392 
<< m1 >>
rect 73 391 74 392 
<< m1 >>
rect 78 391 79 392 
<< m1 >>
rect 82 391 83 392 
<< pdiffusion >>
rect 84 391 85 392 
<< pdiffusion >>
rect 85 391 86 392 
<< pdiffusion >>
rect 86 391 87 392 
<< pdiffusion >>
rect 87 391 88 392 
<< pdiffusion >>
rect 88 391 89 392 
<< pdiffusion >>
rect 89 391 90 392 
<< m1 >>
rect 93 391 94 392 
<< m1 >>
rect 100 391 101 392 
<< pdiffusion >>
rect 102 391 103 392 
<< pdiffusion >>
rect 103 391 104 392 
<< pdiffusion >>
rect 104 391 105 392 
<< pdiffusion >>
rect 105 391 106 392 
<< pdiffusion >>
rect 106 391 107 392 
<< pdiffusion >>
rect 107 391 108 392 
<< m1 >>
rect 110 391 111 392 
<< m1 >>
rect 112 391 113 392 
<< m1 >>
rect 114 391 115 392 
<< m1 >>
rect 118 391 119 392 
<< pdiffusion >>
rect 120 391 121 392 
<< pdiffusion >>
rect 121 391 122 392 
<< pdiffusion >>
rect 122 391 123 392 
<< pdiffusion >>
rect 123 391 124 392 
<< pdiffusion >>
rect 124 391 125 392 
<< pdiffusion >>
rect 125 391 126 392 
<< m1 >>
rect 127 391 128 392 
<< m2 >>
rect 128 391 129 392 
<< m1 >>
rect 136 391 137 392 
<< pdiffusion >>
rect 138 391 139 392 
<< pdiffusion >>
rect 139 391 140 392 
<< pdiffusion >>
rect 140 391 141 392 
<< pdiffusion >>
rect 141 391 142 392 
<< pdiffusion >>
rect 142 391 143 392 
<< pdiffusion >>
rect 143 391 144 392 
<< m1 >>
rect 150 391 151 392 
<< pdiffusion >>
rect 156 391 157 392 
<< pdiffusion >>
rect 157 391 158 392 
<< pdiffusion >>
rect 158 391 159 392 
<< pdiffusion >>
rect 159 391 160 392 
<< pdiffusion >>
rect 160 391 161 392 
<< pdiffusion >>
rect 161 391 162 392 
<< m1 >>
rect 163 391 164 392 
<< m1 >>
rect 167 391 168 392 
<< m1 >>
rect 169 391 170 392 
<< m1 >>
rect 171 391 172 392 
<< pdiffusion >>
rect 174 391 175 392 
<< pdiffusion >>
rect 175 391 176 392 
<< pdiffusion >>
rect 176 391 177 392 
<< pdiffusion >>
rect 177 391 178 392 
<< pdiffusion >>
rect 178 391 179 392 
<< pdiffusion >>
rect 179 391 180 392 
<< m1 >>
rect 190 391 191 392 
<< pdiffusion >>
rect 192 391 193 392 
<< pdiffusion >>
rect 193 391 194 392 
<< pdiffusion >>
rect 194 391 195 392 
<< pdiffusion >>
rect 195 391 196 392 
<< pdiffusion >>
rect 196 391 197 392 
<< pdiffusion >>
rect 197 391 198 392 
<< m1 >>
rect 199 391 200 392 
<< m2 >>
rect 205 391 206 392 
<< m1 >>
rect 206 391 207 392 
<< pdiffusion >>
rect 210 391 211 392 
<< pdiffusion >>
rect 211 391 212 392 
<< pdiffusion >>
rect 212 391 213 392 
<< pdiffusion >>
rect 213 391 214 392 
<< pdiffusion >>
rect 214 391 215 392 
<< pdiffusion >>
rect 215 391 216 392 
<< m1 >>
rect 217 391 218 392 
<< m1 >>
rect 223 391 224 392 
<< pdiffusion >>
rect 228 391 229 392 
<< pdiffusion >>
rect 229 391 230 392 
<< pdiffusion >>
rect 230 391 231 392 
<< pdiffusion >>
rect 231 391 232 392 
<< pdiffusion >>
rect 232 391 233 392 
<< pdiffusion >>
rect 233 391 234 392 
<< m1 >>
rect 235 391 236 392 
<< m1 >>
rect 244 391 245 392 
<< pdiffusion >>
rect 246 391 247 392 
<< pdiffusion >>
rect 247 391 248 392 
<< pdiffusion >>
rect 248 391 249 392 
<< pdiffusion >>
rect 249 391 250 392 
<< pdiffusion >>
rect 250 391 251 392 
<< pdiffusion >>
rect 251 391 252 392 
<< m1 >>
rect 253 391 254 392 
<< m1 >>
rect 255 391 256 392 
<< m1 >>
rect 259 391 260 392 
<< pdiffusion >>
rect 264 391 265 392 
<< pdiffusion >>
rect 265 391 266 392 
<< pdiffusion >>
rect 266 391 267 392 
<< pdiffusion >>
rect 267 391 268 392 
<< pdiffusion >>
rect 268 391 269 392 
<< pdiffusion >>
rect 269 391 270 392 
<< m1 >>
rect 280 391 281 392 
<< pdiffusion >>
rect 282 391 283 392 
<< pdiffusion >>
rect 283 391 284 392 
<< pdiffusion >>
rect 284 391 285 392 
<< pdiffusion >>
rect 285 391 286 392 
<< pdiffusion >>
rect 286 391 287 392 
<< pdiffusion >>
rect 287 391 288 392 
<< pdiffusion >>
rect 300 391 301 392 
<< pdiffusion >>
rect 301 391 302 392 
<< pdiffusion >>
rect 302 391 303 392 
<< pdiffusion >>
rect 303 391 304 392 
<< pdiffusion >>
rect 304 391 305 392 
<< pdiffusion >>
rect 305 391 306 392 
<< m1 >>
rect 307 391 308 392 
<< m1 >>
rect 310 391 311 392 
<< m1 >>
rect 316 391 317 392 
<< pdiffusion >>
rect 318 391 319 392 
<< pdiffusion >>
rect 319 391 320 392 
<< pdiffusion >>
rect 320 391 321 392 
<< pdiffusion >>
rect 321 391 322 392 
<< pdiffusion >>
rect 322 391 323 392 
<< pdiffusion >>
rect 323 391 324 392 
<< m1 >>
rect 325 391 326 392 
<< pdiffusion >>
rect 336 391 337 392 
<< pdiffusion >>
rect 337 391 338 392 
<< pdiffusion >>
rect 338 391 339 392 
<< pdiffusion >>
rect 339 391 340 392 
<< pdiffusion >>
rect 340 391 341 392 
<< pdiffusion >>
rect 341 391 342 392 
<< m1 >>
rect 343 391 344 392 
<< pdiffusion >>
rect 354 391 355 392 
<< pdiffusion >>
rect 355 391 356 392 
<< pdiffusion >>
rect 356 391 357 392 
<< pdiffusion >>
rect 357 391 358 392 
<< pdiffusion >>
rect 358 391 359 392 
<< pdiffusion >>
rect 359 391 360 392 
<< m1 >>
rect 361 391 362 392 
<< m1 >>
rect 363 391 364 392 
<< m2 >>
rect 364 391 365 392 
<< m1 >>
rect 367 391 368 392 
<< pdiffusion >>
rect 372 391 373 392 
<< pdiffusion >>
rect 373 391 374 392 
<< pdiffusion >>
rect 374 391 375 392 
<< pdiffusion >>
rect 375 391 376 392 
<< pdiffusion >>
rect 376 391 377 392 
<< pdiffusion >>
rect 377 391 378 392 
<< m1 >>
rect 385 391 386 392 
<< m1 >>
rect 402 391 403 392 
<< m1 >>
rect 406 391 407 392 
<< pdiffusion >>
rect 408 391 409 392 
<< pdiffusion >>
rect 409 391 410 392 
<< pdiffusion >>
rect 410 391 411 392 
<< pdiffusion >>
rect 411 391 412 392 
<< pdiffusion >>
rect 412 391 413 392 
<< pdiffusion >>
rect 413 391 414 392 
<< m1 >>
rect 416 391 417 392 
<< m1 >>
rect 418 391 419 392 
<< pdiffusion >>
rect 426 391 427 392 
<< pdiffusion >>
rect 427 391 428 392 
<< pdiffusion >>
rect 428 391 429 392 
<< pdiffusion >>
rect 429 391 430 392 
<< pdiffusion >>
rect 430 391 431 392 
<< pdiffusion >>
rect 431 391 432 392 
<< m1 >>
rect 433 391 434 392 
<< m1 >>
rect 435 391 436 392 
<< m1 >>
rect 437 391 438 392 
<< pdiffusion >>
rect 444 391 445 392 
<< pdiffusion >>
rect 445 391 446 392 
<< pdiffusion >>
rect 446 391 447 392 
<< pdiffusion >>
rect 447 391 448 392 
<< pdiffusion >>
rect 448 391 449 392 
<< pdiffusion >>
rect 449 391 450 392 
<< m1 >>
rect 451 391 452 392 
<< m1 >>
rect 457 391 458 392 
<< m1 >>
rect 459 391 460 392 
<< pdiffusion >>
rect 462 391 463 392 
<< pdiffusion >>
rect 463 391 464 392 
<< pdiffusion >>
rect 464 391 465 392 
<< pdiffusion >>
rect 465 391 466 392 
<< pdiffusion >>
rect 466 391 467 392 
<< pdiffusion >>
rect 467 391 468 392 
<< m1 >>
rect 472 391 473 392 
<< m1 >>
rect 476 391 477 392 
<< m1 >>
rect 478 391 479 392 
<< pdiffusion >>
rect 480 391 481 392 
<< pdiffusion >>
rect 481 391 482 392 
<< pdiffusion >>
rect 482 391 483 392 
<< pdiffusion >>
rect 483 391 484 392 
<< pdiffusion >>
rect 484 391 485 392 
<< pdiffusion >>
rect 485 391 486 392 
<< pdiffusion >>
rect 498 391 499 392 
<< pdiffusion >>
rect 499 391 500 392 
<< pdiffusion >>
rect 500 391 501 392 
<< pdiffusion >>
rect 501 391 502 392 
<< pdiffusion >>
rect 502 391 503 392 
<< pdiffusion >>
rect 503 391 504 392 
<< pdiffusion >>
rect 516 391 517 392 
<< pdiffusion >>
rect 517 391 518 392 
<< pdiffusion >>
rect 518 391 519 392 
<< pdiffusion >>
rect 519 391 520 392 
<< pdiffusion >>
rect 520 391 521 392 
<< pdiffusion >>
rect 521 391 522 392 
<< m1 >>
rect 523 391 524 392 
<< pdiffusion >>
rect 12 392 13 393 
<< pdiffusion >>
rect 13 392 14 393 
<< pdiffusion >>
rect 14 392 15 393 
<< pdiffusion >>
rect 15 392 16 393 
<< pdiffusion >>
rect 16 392 17 393 
<< pdiffusion >>
rect 17 392 18 393 
<< m1 >>
rect 19 392 20 393 
<< m2 >>
rect 20 392 21 393 
<< m1 >>
rect 23 392 24 393 
<< pdiffusion >>
rect 30 392 31 393 
<< pdiffusion >>
rect 31 392 32 393 
<< pdiffusion >>
rect 32 392 33 393 
<< pdiffusion >>
rect 33 392 34 393 
<< pdiffusion >>
rect 34 392 35 393 
<< pdiffusion >>
rect 35 392 36 393 
<< m1 >>
rect 42 392 43 393 
<< m1 >>
rect 44 392 45 393 
<< pdiffusion >>
rect 48 392 49 393 
<< pdiffusion >>
rect 49 392 50 393 
<< pdiffusion >>
rect 50 392 51 393 
<< pdiffusion >>
rect 51 392 52 393 
<< pdiffusion >>
rect 52 392 53 393 
<< pdiffusion >>
rect 53 392 54 393 
<< m2 >>
rect 63 392 64 393 
<< m1 >>
rect 64 392 65 393 
<< pdiffusion >>
rect 66 392 67 393 
<< pdiffusion >>
rect 67 392 68 393 
<< pdiffusion >>
rect 68 392 69 393 
<< pdiffusion >>
rect 69 392 70 393 
<< pdiffusion >>
rect 70 392 71 393 
<< pdiffusion >>
rect 71 392 72 393 
<< m1 >>
rect 73 392 74 393 
<< m1 >>
rect 78 392 79 393 
<< m1 >>
rect 82 392 83 393 
<< pdiffusion >>
rect 84 392 85 393 
<< pdiffusion >>
rect 85 392 86 393 
<< pdiffusion >>
rect 86 392 87 393 
<< pdiffusion >>
rect 87 392 88 393 
<< pdiffusion >>
rect 88 392 89 393 
<< pdiffusion >>
rect 89 392 90 393 
<< m1 >>
rect 93 392 94 393 
<< m1 >>
rect 100 392 101 393 
<< pdiffusion >>
rect 102 392 103 393 
<< pdiffusion >>
rect 103 392 104 393 
<< pdiffusion >>
rect 104 392 105 393 
<< pdiffusion >>
rect 105 392 106 393 
<< pdiffusion >>
rect 106 392 107 393 
<< pdiffusion >>
rect 107 392 108 393 
<< m1 >>
rect 110 392 111 393 
<< m1 >>
rect 112 392 113 393 
<< m1 >>
rect 114 392 115 393 
<< m1 >>
rect 118 392 119 393 
<< pdiffusion >>
rect 120 392 121 393 
<< pdiffusion >>
rect 121 392 122 393 
<< pdiffusion >>
rect 122 392 123 393 
<< pdiffusion >>
rect 123 392 124 393 
<< pdiffusion >>
rect 124 392 125 393 
<< pdiffusion >>
rect 125 392 126 393 
<< m1 >>
rect 127 392 128 393 
<< m2 >>
rect 128 392 129 393 
<< m1 >>
rect 136 392 137 393 
<< pdiffusion >>
rect 138 392 139 393 
<< pdiffusion >>
rect 139 392 140 393 
<< pdiffusion >>
rect 140 392 141 393 
<< pdiffusion >>
rect 141 392 142 393 
<< pdiffusion >>
rect 142 392 143 393 
<< pdiffusion >>
rect 143 392 144 393 
<< m1 >>
rect 150 392 151 393 
<< pdiffusion >>
rect 156 392 157 393 
<< pdiffusion >>
rect 157 392 158 393 
<< pdiffusion >>
rect 158 392 159 393 
<< pdiffusion >>
rect 159 392 160 393 
<< pdiffusion >>
rect 160 392 161 393 
<< pdiffusion >>
rect 161 392 162 393 
<< m1 >>
rect 163 392 164 393 
<< m1 >>
rect 167 392 168 393 
<< m1 >>
rect 169 392 170 393 
<< m1 >>
rect 171 392 172 393 
<< pdiffusion >>
rect 174 392 175 393 
<< pdiffusion >>
rect 175 392 176 393 
<< pdiffusion >>
rect 176 392 177 393 
<< pdiffusion >>
rect 177 392 178 393 
<< pdiffusion >>
rect 178 392 179 393 
<< pdiffusion >>
rect 179 392 180 393 
<< m1 >>
rect 190 392 191 393 
<< pdiffusion >>
rect 192 392 193 393 
<< pdiffusion >>
rect 193 392 194 393 
<< pdiffusion >>
rect 194 392 195 393 
<< pdiffusion >>
rect 195 392 196 393 
<< pdiffusion >>
rect 196 392 197 393 
<< pdiffusion >>
rect 197 392 198 393 
<< m1 >>
rect 199 392 200 393 
<< m2 >>
rect 205 392 206 393 
<< m1 >>
rect 206 392 207 393 
<< pdiffusion >>
rect 210 392 211 393 
<< pdiffusion >>
rect 211 392 212 393 
<< pdiffusion >>
rect 212 392 213 393 
<< pdiffusion >>
rect 213 392 214 393 
<< pdiffusion >>
rect 214 392 215 393 
<< pdiffusion >>
rect 215 392 216 393 
<< m1 >>
rect 217 392 218 393 
<< m1 >>
rect 223 392 224 393 
<< pdiffusion >>
rect 228 392 229 393 
<< pdiffusion >>
rect 229 392 230 393 
<< pdiffusion >>
rect 230 392 231 393 
<< pdiffusion >>
rect 231 392 232 393 
<< pdiffusion >>
rect 232 392 233 393 
<< pdiffusion >>
rect 233 392 234 393 
<< m1 >>
rect 235 392 236 393 
<< m1 >>
rect 244 392 245 393 
<< pdiffusion >>
rect 246 392 247 393 
<< pdiffusion >>
rect 247 392 248 393 
<< pdiffusion >>
rect 248 392 249 393 
<< pdiffusion >>
rect 249 392 250 393 
<< pdiffusion >>
rect 250 392 251 393 
<< pdiffusion >>
rect 251 392 252 393 
<< m1 >>
rect 253 392 254 393 
<< m1 >>
rect 255 392 256 393 
<< m1 >>
rect 259 392 260 393 
<< pdiffusion >>
rect 264 392 265 393 
<< pdiffusion >>
rect 265 392 266 393 
<< pdiffusion >>
rect 266 392 267 393 
<< pdiffusion >>
rect 267 392 268 393 
<< pdiffusion >>
rect 268 392 269 393 
<< pdiffusion >>
rect 269 392 270 393 
<< m1 >>
rect 280 392 281 393 
<< pdiffusion >>
rect 282 392 283 393 
<< pdiffusion >>
rect 283 392 284 393 
<< pdiffusion >>
rect 284 392 285 393 
<< pdiffusion >>
rect 285 392 286 393 
<< pdiffusion >>
rect 286 392 287 393 
<< pdiffusion >>
rect 287 392 288 393 
<< pdiffusion >>
rect 300 392 301 393 
<< pdiffusion >>
rect 301 392 302 393 
<< pdiffusion >>
rect 302 392 303 393 
<< pdiffusion >>
rect 303 392 304 393 
<< pdiffusion >>
rect 304 392 305 393 
<< pdiffusion >>
rect 305 392 306 393 
<< m1 >>
rect 307 392 308 393 
<< m1 >>
rect 310 392 311 393 
<< m1 >>
rect 316 392 317 393 
<< pdiffusion >>
rect 318 392 319 393 
<< pdiffusion >>
rect 319 392 320 393 
<< pdiffusion >>
rect 320 392 321 393 
<< pdiffusion >>
rect 321 392 322 393 
<< pdiffusion >>
rect 322 392 323 393 
<< pdiffusion >>
rect 323 392 324 393 
<< m1 >>
rect 325 392 326 393 
<< pdiffusion >>
rect 336 392 337 393 
<< pdiffusion >>
rect 337 392 338 393 
<< pdiffusion >>
rect 338 392 339 393 
<< pdiffusion >>
rect 339 392 340 393 
<< pdiffusion >>
rect 340 392 341 393 
<< pdiffusion >>
rect 341 392 342 393 
<< m1 >>
rect 343 392 344 393 
<< pdiffusion >>
rect 354 392 355 393 
<< pdiffusion >>
rect 355 392 356 393 
<< pdiffusion >>
rect 356 392 357 393 
<< pdiffusion >>
rect 357 392 358 393 
<< pdiffusion >>
rect 358 392 359 393 
<< pdiffusion >>
rect 359 392 360 393 
<< m1 >>
rect 361 392 362 393 
<< m1 >>
rect 363 392 364 393 
<< m2 >>
rect 364 392 365 393 
<< m1 >>
rect 367 392 368 393 
<< pdiffusion >>
rect 372 392 373 393 
<< pdiffusion >>
rect 373 392 374 393 
<< pdiffusion >>
rect 374 392 375 393 
<< pdiffusion >>
rect 375 392 376 393 
<< pdiffusion >>
rect 376 392 377 393 
<< pdiffusion >>
rect 377 392 378 393 
<< m1 >>
rect 385 392 386 393 
<< m1 >>
rect 402 392 403 393 
<< m1 >>
rect 406 392 407 393 
<< pdiffusion >>
rect 408 392 409 393 
<< pdiffusion >>
rect 409 392 410 393 
<< pdiffusion >>
rect 410 392 411 393 
<< pdiffusion >>
rect 411 392 412 393 
<< pdiffusion >>
rect 412 392 413 393 
<< pdiffusion >>
rect 413 392 414 393 
<< m1 >>
rect 416 392 417 393 
<< m1 >>
rect 418 392 419 393 
<< pdiffusion >>
rect 426 392 427 393 
<< pdiffusion >>
rect 427 392 428 393 
<< pdiffusion >>
rect 428 392 429 393 
<< pdiffusion >>
rect 429 392 430 393 
<< pdiffusion >>
rect 430 392 431 393 
<< pdiffusion >>
rect 431 392 432 393 
<< m1 >>
rect 433 392 434 393 
<< m1 >>
rect 435 392 436 393 
<< m1 >>
rect 437 392 438 393 
<< pdiffusion >>
rect 444 392 445 393 
<< pdiffusion >>
rect 445 392 446 393 
<< pdiffusion >>
rect 446 392 447 393 
<< pdiffusion >>
rect 447 392 448 393 
<< pdiffusion >>
rect 448 392 449 393 
<< pdiffusion >>
rect 449 392 450 393 
<< m1 >>
rect 451 392 452 393 
<< m1 >>
rect 457 392 458 393 
<< m1 >>
rect 459 392 460 393 
<< pdiffusion >>
rect 462 392 463 393 
<< pdiffusion >>
rect 463 392 464 393 
<< pdiffusion >>
rect 464 392 465 393 
<< pdiffusion >>
rect 465 392 466 393 
<< pdiffusion >>
rect 466 392 467 393 
<< pdiffusion >>
rect 467 392 468 393 
<< m1 >>
rect 472 392 473 393 
<< m1 >>
rect 476 392 477 393 
<< m1 >>
rect 478 392 479 393 
<< pdiffusion >>
rect 480 392 481 393 
<< pdiffusion >>
rect 481 392 482 393 
<< pdiffusion >>
rect 482 392 483 393 
<< pdiffusion >>
rect 483 392 484 393 
<< pdiffusion >>
rect 484 392 485 393 
<< pdiffusion >>
rect 485 392 486 393 
<< pdiffusion >>
rect 498 392 499 393 
<< pdiffusion >>
rect 499 392 500 393 
<< pdiffusion >>
rect 500 392 501 393 
<< pdiffusion >>
rect 501 392 502 393 
<< pdiffusion >>
rect 502 392 503 393 
<< pdiffusion >>
rect 503 392 504 393 
<< pdiffusion >>
rect 516 392 517 393 
<< pdiffusion >>
rect 517 392 518 393 
<< pdiffusion >>
rect 518 392 519 393 
<< pdiffusion >>
rect 519 392 520 393 
<< pdiffusion >>
rect 520 392 521 393 
<< pdiffusion >>
rect 521 392 522 393 
<< m1 >>
rect 523 392 524 393 
<< pdiffusion >>
rect 12 393 13 394 
<< pdiffusion >>
rect 13 393 14 394 
<< pdiffusion >>
rect 14 393 15 394 
<< pdiffusion >>
rect 15 393 16 394 
<< pdiffusion >>
rect 16 393 17 394 
<< pdiffusion >>
rect 17 393 18 394 
<< m1 >>
rect 19 393 20 394 
<< m2 >>
rect 20 393 21 394 
<< m1 >>
rect 23 393 24 394 
<< pdiffusion >>
rect 30 393 31 394 
<< pdiffusion >>
rect 31 393 32 394 
<< pdiffusion >>
rect 32 393 33 394 
<< pdiffusion >>
rect 33 393 34 394 
<< pdiffusion >>
rect 34 393 35 394 
<< pdiffusion >>
rect 35 393 36 394 
<< m1 >>
rect 42 393 43 394 
<< m1 >>
rect 44 393 45 394 
<< pdiffusion >>
rect 48 393 49 394 
<< pdiffusion >>
rect 49 393 50 394 
<< pdiffusion >>
rect 50 393 51 394 
<< pdiffusion >>
rect 51 393 52 394 
<< pdiffusion >>
rect 52 393 53 394 
<< pdiffusion >>
rect 53 393 54 394 
<< m2 >>
rect 63 393 64 394 
<< m1 >>
rect 64 393 65 394 
<< pdiffusion >>
rect 66 393 67 394 
<< pdiffusion >>
rect 67 393 68 394 
<< pdiffusion >>
rect 68 393 69 394 
<< pdiffusion >>
rect 69 393 70 394 
<< pdiffusion >>
rect 70 393 71 394 
<< pdiffusion >>
rect 71 393 72 394 
<< m1 >>
rect 73 393 74 394 
<< m1 >>
rect 78 393 79 394 
<< m1 >>
rect 82 393 83 394 
<< pdiffusion >>
rect 84 393 85 394 
<< pdiffusion >>
rect 85 393 86 394 
<< pdiffusion >>
rect 86 393 87 394 
<< pdiffusion >>
rect 87 393 88 394 
<< pdiffusion >>
rect 88 393 89 394 
<< pdiffusion >>
rect 89 393 90 394 
<< m1 >>
rect 93 393 94 394 
<< m1 >>
rect 100 393 101 394 
<< pdiffusion >>
rect 102 393 103 394 
<< pdiffusion >>
rect 103 393 104 394 
<< pdiffusion >>
rect 104 393 105 394 
<< pdiffusion >>
rect 105 393 106 394 
<< pdiffusion >>
rect 106 393 107 394 
<< pdiffusion >>
rect 107 393 108 394 
<< m1 >>
rect 110 393 111 394 
<< m1 >>
rect 112 393 113 394 
<< m1 >>
rect 114 393 115 394 
<< m1 >>
rect 118 393 119 394 
<< pdiffusion >>
rect 120 393 121 394 
<< pdiffusion >>
rect 121 393 122 394 
<< pdiffusion >>
rect 122 393 123 394 
<< pdiffusion >>
rect 123 393 124 394 
<< pdiffusion >>
rect 124 393 125 394 
<< pdiffusion >>
rect 125 393 126 394 
<< m1 >>
rect 127 393 128 394 
<< m2 >>
rect 128 393 129 394 
<< m1 >>
rect 136 393 137 394 
<< pdiffusion >>
rect 138 393 139 394 
<< pdiffusion >>
rect 139 393 140 394 
<< pdiffusion >>
rect 140 393 141 394 
<< pdiffusion >>
rect 141 393 142 394 
<< pdiffusion >>
rect 142 393 143 394 
<< pdiffusion >>
rect 143 393 144 394 
<< m1 >>
rect 150 393 151 394 
<< pdiffusion >>
rect 156 393 157 394 
<< pdiffusion >>
rect 157 393 158 394 
<< pdiffusion >>
rect 158 393 159 394 
<< pdiffusion >>
rect 159 393 160 394 
<< pdiffusion >>
rect 160 393 161 394 
<< pdiffusion >>
rect 161 393 162 394 
<< m1 >>
rect 163 393 164 394 
<< m1 >>
rect 167 393 168 394 
<< m2 >>
rect 167 393 168 394 
<< m2c >>
rect 167 393 168 394 
<< m1 >>
rect 167 393 168 394 
<< m2 >>
rect 167 393 168 394 
<< m1 >>
rect 169 393 170 394 
<< m2 >>
rect 169 393 170 394 
<< m2c >>
rect 169 393 170 394 
<< m1 >>
rect 169 393 170 394 
<< m2 >>
rect 169 393 170 394 
<< m1 >>
rect 171 393 172 394 
<< pdiffusion >>
rect 174 393 175 394 
<< pdiffusion >>
rect 175 393 176 394 
<< pdiffusion >>
rect 176 393 177 394 
<< pdiffusion >>
rect 177 393 178 394 
<< pdiffusion >>
rect 178 393 179 394 
<< pdiffusion >>
rect 179 393 180 394 
<< m1 >>
rect 190 393 191 394 
<< pdiffusion >>
rect 192 393 193 394 
<< pdiffusion >>
rect 193 393 194 394 
<< pdiffusion >>
rect 194 393 195 394 
<< pdiffusion >>
rect 195 393 196 394 
<< pdiffusion >>
rect 196 393 197 394 
<< pdiffusion >>
rect 197 393 198 394 
<< m1 >>
rect 199 393 200 394 
<< m2 >>
rect 205 393 206 394 
<< m1 >>
rect 206 393 207 394 
<< pdiffusion >>
rect 210 393 211 394 
<< pdiffusion >>
rect 211 393 212 394 
<< pdiffusion >>
rect 212 393 213 394 
<< pdiffusion >>
rect 213 393 214 394 
<< pdiffusion >>
rect 214 393 215 394 
<< pdiffusion >>
rect 215 393 216 394 
<< m1 >>
rect 217 393 218 394 
<< m1 >>
rect 223 393 224 394 
<< pdiffusion >>
rect 228 393 229 394 
<< pdiffusion >>
rect 229 393 230 394 
<< pdiffusion >>
rect 230 393 231 394 
<< pdiffusion >>
rect 231 393 232 394 
<< pdiffusion >>
rect 232 393 233 394 
<< pdiffusion >>
rect 233 393 234 394 
<< m1 >>
rect 235 393 236 394 
<< m1 >>
rect 244 393 245 394 
<< pdiffusion >>
rect 246 393 247 394 
<< pdiffusion >>
rect 247 393 248 394 
<< pdiffusion >>
rect 248 393 249 394 
<< pdiffusion >>
rect 249 393 250 394 
<< pdiffusion >>
rect 250 393 251 394 
<< pdiffusion >>
rect 251 393 252 394 
<< m1 >>
rect 253 393 254 394 
<< m1 >>
rect 255 393 256 394 
<< m1 >>
rect 259 393 260 394 
<< pdiffusion >>
rect 264 393 265 394 
<< pdiffusion >>
rect 265 393 266 394 
<< pdiffusion >>
rect 266 393 267 394 
<< pdiffusion >>
rect 267 393 268 394 
<< pdiffusion >>
rect 268 393 269 394 
<< pdiffusion >>
rect 269 393 270 394 
<< m1 >>
rect 280 393 281 394 
<< pdiffusion >>
rect 282 393 283 394 
<< pdiffusion >>
rect 283 393 284 394 
<< pdiffusion >>
rect 284 393 285 394 
<< pdiffusion >>
rect 285 393 286 394 
<< pdiffusion >>
rect 286 393 287 394 
<< pdiffusion >>
rect 287 393 288 394 
<< pdiffusion >>
rect 300 393 301 394 
<< pdiffusion >>
rect 301 393 302 394 
<< pdiffusion >>
rect 302 393 303 394 
<< pdiffusion >>
rect 303 393 304 394 
<< pdiffusion >>
rect 304 393 305 394 
<< pdiffusion >>
rect 305 393 306 394 
<< m1 >>
rect 307 393 308 394 
<< m1 >>
rect 310 393 311 394 
<< m1 >>
rect 316 393 317 394 
<< pdiffusion >>
rect 318 393 319 394 
<< pdiffusion >>
rect 319 393 320 394 
<< pdiffusion >>
rect 320 393 321 394 
<< pdiffusion >>
rect 321 393 322 394 
<< pdiffusion >>
rect 322 393 323 394 
<< pdiffusion >>
rect 323 393 324 394 
<< m1 >>
rect 325 393 326 394 
<< pdiffusion >>
rect 336 393 337 394 
<< pdiffusion >>
rect 337 393 338 394 
<< pdiffusion >>
rect 338 393 339 394 
<< pdiffusion >>
rect 339 393 340 394 
<< pdiffusion >>
rect 340 393 341 394 
<< pdiffusion >>
rect 341 393 342 394 
<< m1 >>
rect 343 393 344 394 
<< pdiffusion >>
rect 354 393 355 394 
<< pdiffusion >>
rect 355 393 356 394 
<< pdiffusion >>
rect 356 393 357 394 
<< pdiffusion >>
rect 357 393 358 394 
<< pdiffusion >>
rect 358 393 359 394 
<< pdiffusion >>
rect 359 393 360 394 
<< m1 >>
rect 361 393 362 394 
<< m1 >>
rect 363 393 364 394 
<< m2 >>
rect 364 393 365 394 
<< m1 >>
rect 367 393 368 394 
<< pdiffusion >>
rect 372 393 373 394 
<< pdiffusion >>
rect 373 393 374 394 
<< pdiffusion >>
rect 374 393 375 394 
<< pdiffusion >>
rect 375 393 376 394 
<< pdiffusion >>
rect 376 393 377 394 
<< pdiffusion >>
rect 377 393 378 394 
<< m1 >>
rect 385 393 386 394 
<< m1 >>
rect 402 393 403 394 
<< m1 >>
rect 406 393 407 394 
<< pdiffusion >>
rect 408 393 409 394 
<< pdiffusion >>
rect 409 393 410 394 
<< pdiffusion >>
rect 410 393 411 394 
<< pdiffusion >>
rect 411 393 412 394 
<< pdiffusion >>
rect 412 393 413 394 
<< pdiffusion >>
rect 413 393 414 394 
<< m1 >>
rect 416 393 417 394 
<< m1 >>
rect 418 393 419 394 
<< pdiffusion >>
rect 426 393 427 394 
<< pdiffusion >>
rect 427 393 428 394 
<< pdiffusion >>
rect 428 393 429 394 
<< pdiffusion >>
rect 429 393 430 394 
<< pdiffusion >>
rect 430 393 431 394 
<< pdiffusion >>
rect 431 393 432 394 
<< m1 >>
rect 433 393 434 394 
<< m1 >>
rect 435 393 436 394 
<< m1 >>
rect 437 393 438 394 
<< pdiffusion >>
rect 444 393 445 394 
<< pdiffusion >>
rect 445 393 446 394 
<< pdiffusion >>
rect 446 393 447 394 
<< pdiffusion >>
rect 447 393 448 394 
<< pdiffusion >>
rect 448 393 449 394 
<< pdiffusion >>
rect 449 393 450 394 
<< m1 >>
rect 451 393 452 394 
<< m1 >>
rect 455 393 456 394 
<< m2 >>
rect 455 393 456 394 
<< m2c >>
rect 455 393 456 394 
<< m1 >>
rect 455 393 456 394 
<< m2 >>
rect 455 393 456 394 
<< m2 >>
rect 456 393 457 394 
<< m1 >>
rect 457 393 458 394 
<< m2 >>
rect 457 393 458 394 
<< m2 >>
rect 458 393 459 394 
<< m1 >>
rect 459 393 460 394 
<< m2 >>
rect 459 393 460 394 
<< m2c >>
rect 459 393 460 394 
<< m1 >>
rect 459 393 460 394 
<< m2 >>
rect 459 393 460 394 
<< pdiffusion >>
rect 462 393 463 394 
<< pdiffusion >>
rect 463 393 464 394 
<< pdiffusion >>
rect 464 393 465 394 
<< pdiffusion >>
rect 465 393 466 394 
<< pdiffusion >>
rect 466 393 467 394 
<< pdiffusion >>
rect 467 393 468 394 
<< m1 >>
rect 472 393 473 394 
<< m1 >>
rect 476 393 477 394 
<< m1 >>
rect 478 393 479 394 
<< pdiffusion >>
rect 480 393 481 394 
<< pdiffusion >>
rect 481 393 482 394 
<< pdiffusion >>
rect 482 393 483 394 
<< pdiffusion >>
rect 483 393 484 394 
<< pdiffusion >>
rect 484 393 485 394 
<< pdiffusion >>
rect 485 393 486 394 
<< pdiffusion >>
rect 498 393 499 394 
<< pdiffusion >>
rect 499 393 500 394 
<< pdiffusion >>
rect 500 393 501 394 
<< pdiffusion >>
rect 501 393 502 394 
<< pdiffusion >>
rect 502 393 503 394 
<< pdiffusion >>
rect 503 393 504 394 
<< pdiffusion >>
rect 516 393 517 394 
<< pdiffusion >>
rect 517 393 518 394 
<< pdiffusion >>
rect 518 393 519 394 
<< pdiffusion >>
rect 519 393 520 394 
<< pdiffusion >>
rect 520 393 521 394 
<< pdiffusion >>
rect 521 393 522 394 
<< m1 >>
rect 523 393 524 394 
<< pdiffusion >>
rect 12 394 13 395 
<< pdiffusion >>
rect 13 394 14 395 
<< pdiffusion >>
rect 14 394 15 395 
<< pdiffusion >>
rect 15 394 16 395 
<< pdiffusion >>
rect 16 394 17 395 
<< pdiffusion >>
rect 17 394 18 395 
<< m1 >>
rect 19 394 20 395 
<< m2 >>
rect 20 394 21 395 
<< m1 >>
rect 23 394 24 395 
<< pdiffusion >>
rect 30 394 31 395 
<< pdiffusion >>
rect 31 394 32 395 
<< pdiffusion >>
rect 32 394 33 395 
<< pdiffusion >>
rect 33 394 34 395 
<< pdiffusion >>
rect 34 394 35 395 
<< pdiffusion >>
rect 35 394 36 395 
<< m1 >>
rect 42 394 43 395 
<< m1 >>
rect 44 394 45 395 
<< pdiffusion >>
rect 48 394 49 395 
<< pdiffusion >>
rect 49 394 50 395 
<< pdiffusion >>
rect 50 394 51 395 
<< pdiffusion >>
rect 51 394 52 395 
<< pdiffusion >>
rect 52 394 53 395 
<< pdiffusion >>
rect 53 394 54 395 
<< m2 >>
rect 63 394 64 395 
<< m1 >>
rect 64 394 65 395 
<< pdiffusion >>
rect 66 394 67 395 
<< pdiffusion >>
rect 67 394 68 395 
<< pdiffusion >>
rect 68 394 69 395 
<< pdiffusion >>
rect 69 394 70 395 
<< pdiffusion >>
rect 70 394 71 395 
<< pdiffusion >>
rect 71 394 72 395 
<< m1 >>
rect 73 394 74 395 
<< m1 >>
rect 78 394 79 395 
<< m1 >>
rect 82 394 83 395 
<< pdiffusion >>
rect 84 394 85 395 
<< pdiffusion >>
rect 85 394 86 395 
<< pdiffusion >>
rect 86 394 87 395 
<< pdiffusion >>
rect 87 394 88 395 
<< pdiffusion >>
rect 88 394 89 395 
<< pdiffusion >>
rect 89 394 90 395 
<< m1 >>
rect 93 394 94 395 
<< m1 >>
rect 100 394 101 395 
<< pdiffusion >>
rect 102 394 103 395 
<< pdiffusion >>
rect 103 394 104 395 
<< pdiffusion >>
rect 104 394 105 395 
<< pdiffusion >>
rect 105 394 106 395 
<< pdiffusion >>
rect 106 394 107 395 
<< pdiffusion >>
rect 107 394 108 395 
<< m1 >>
rect 110 394 111 395 
<< m1 >>
rect 112 394 113 395 
<< m1 >>
rect 114 394 115 395 
<< m1 >>
rect 118 394 119 395 
<< pdiffusion >>
rect 120 394 121 395 
<< pdiffusion >>
rect 121 394 122 395 
<< pdiffusion >>
rect 122 394 123 395 
<< pdiffusion >>
rect 123 394 124 395 
<< pdiffusion >>
rect 124 394 125 395 
<< pdiffusion >>
rect 125 394 126 395 
<< m1 >>
rect 127 394 128 395 
<< m2 >>
rect 128 394 129 395 
<< m1 >>
rect 136 394 137 395 
<< pdiffusion >>
rect 138 394 139 395 
<< pdiffusion >>
rect 139 394 140 395 
<< pdiffusion >>
rect 140 394 141 395 
<< pdiffusion >>
rect 141 394 142 395 
<< pdiffusion >>
rect 142 394 143 395 
<< pdiffusion >>
rect 143 394 144 395 
<< m1 >>
rect 150 394 151 395 
<< pdiffusion >>
rect 156 394 157 395 
<< pdiffusion >>
rect 157 394 158 395 
<< pdiffusion >>
rect 158 394 159 395 
<< pdiffusion >>
rect 159 394 160 395 
<< pdiffusion >>
rect 160 394 161 395 
<< pdiffusion >>
rect 161 394 162 395 
<< m1 >>
rect 163 394 164 395 
<< m2 >>
rect 167 394 168 395 
<< m2 >>
rect 169 394 170 395 
<< m1 >>
rect 171 394 172 395 
<< pdiffusion >>
rect 174 394 175 395 
<< pdiffusion >>
rect 175 394 176 395 
<< pdiffusion >>
rect 176 394 177 395 
<< pdiffusion >>
rect 177 394 178 395 
<< pdiffusion >>
rect 178 394 179 395 
<< pdiffusion >>
rect 179 394 180 395 
<< m1 >>
rect 190 394 191 395 
<< pdiffusion >>
rect 192 394 193 395 
<< pdiffusion >>
rect 193 394 194 395 
<< pdiffusion >>
rect 194 394 195 395 
<< pdiffusion >>
rect 195 394 196 395 
<< pdiffusion >>
rect 196 394 197 395 
<< pdiffusion >>
rect 197 394 198 395 
<< m1 >>
rect 199 394 200 395 
<< m2 >>
rect 205 394 206 395 
<< m1 >>
rect 206 394 207 395 
<< pdiffusion >>
rect 210 394 211 395 
<< pdiffusion >>
rect 211 394 212 395 
<< pdiffusion >>
rect 212 394 213 395 
<< pdiffusion >>
rect 213 394 214 395 
<< pdiffusion >>
rect 214 394 215 395 
<< pdiffusion >>
rect 215 394 216 395 
<< m1 >>
rect 217 394 218 395 
<< m1 >>
rect 223 394 224 395 
<< pdiffusion >>
rect 228 394 229 395 
<< pdiffusion >>
rect 229 394 230 395 
<< pdiffusion >>
rect 230 394 231 395 
<< pdiffusion >>
rect 231 394 232 395 
<< pdiffusion >>
rect 232 394 233 395 
<< pdiffusion >>
rect 233 394 234 395 
<< m1 >>
rect 235 394 236 395 
<< m1 >>
rect 244 394 245 395 
<< pdiffusion >>
rect 246 394 247 395 
<< pdiffusion >>
rect 247 394 248 395 
<< pdiffusion >>
rect 248 394 249 395 
<< pdiffusion >>
rect 249 394 250 395 
<< pdiffusion >>
rect 250 394 251 395 
<< pdiffusion >>
rect 251 394 252 395 
<< m1 >>
rect 253 394 254 395 
<< m1 >>
rect 255 394 256 395 
<< m1 >>
rect 259 394 260 395 
<< pdiffusion >>
rect 264 394 265 395 
<< pdiffusion >>
rect 265 394 266 395 
<< pdiffusion >>
rect 266 394 267 395 
<< pdiffusion >>
rect 267 394 268 395 
<< pdiffusion >>
rect 268 394 269 395 
<< pdiffusion >>
rect 269 394 270 395 
<< m1 >>
rect 280 394 281 395 
<< pdiffusion >>
rect 282 394 283 395 
<< pdiffusion >>
rect 283 394 284 395 
<< pdiffusion >>
rect 284 394 285 395 
<< pdiffusion >>
rect 285 394 286 395 
<< pdiffusion >>
rect 286 394 287 395 
<< pdiffusion >>
rect 287 394 288 395 
<< pdiffusion >>
rect 300 394 301 395 
<< pdiffusion >>
rect 301 394 302 395 
<< pdiffusion >>
rect 302 394 303 395 
<< pdiffusion >>
rect 303 394 304 395 
<< pdiffusion >>
rect 304 394 305 395 
<< pdiffusion >>
rect 305 394 306 395 
<< m1 >>
rect 307 394 308 395 
<< m1 >>
rect 310 394 311 395 
<< m1 >>
rect 316 394 317 395 
<< pdiffusion >>
rect 318 394 319 395 
<< pdiffusion >>
rect 319 394 320 395 
<< pdiffusion >>
rect 320 394 321 395 
<< pdiffusion >>
rect 321 394 322 395 
<< pdiffusion >>
rect 322 394 323 395 
<< pdiffusion >>
rect 323 394 324 395 
<< m1 >>
rect 325 394 326 395 
<< pdiffusion >>
rect 336 394 337 395 
<< pdiffusion >>
rect 337 394 338 395 
<< pdiffusion >>
rect 338 394 339 395 
<< pdiffusion >>
rect 339 394 340 395 
<< pdiffusion >>
rect 340 394 341 395 
<< pdiffusion >>
rect 341 394 342 395 
<< m1 >>
rect 343 394 344 395 
<< pdiffusion >>
rect 354 394 355 395 
<< pdiffusion >>
rect 355 394 356 395 
<< pdiffusion >>
rect 356 394 357 395 
<< pdiffusion >>
rect 357 394 358 395 
<< pdiffusion >>
rect 358 394 359 395 
<< pdiffusion >>
rect 359 394 360 395 
<< m1 >>
rect 361 394 362 395 
<< m1 >>
rect 363 394 364 395 
<< m2 >>
rect 364 394 365 395 
<< m1 >>
rect 367 394 368 395 
<< pdiffusion >>
rect 372 394 373 395 
<< pdiffusion >>
rect 373 394 374 395 
<< pdiffusion >>
rect 374 394 375 395 
<< pdiffusion >>
rect 375 394 376 395 
<< pdiffusion >>
rect 376 394 377 395 
<< pdiffusion >>
rect 377 394 378 395 
<< m1 >>
rect 385 394 386 395 
<< m1 >>
rect 402 394 403 395 
<< m1 >>
rect 406 394 407 395 
<< pdiffusion >>
rect 408 394 409 395 
<< pdiffusion >>
rect 409 394 410 395 
<< pdiffusion >>
rect 410 394 411 395 
<< pdiffusion >>
rect 411 394 412 395 
<< pdiffusion >>
rect 412 394 413 395 
<< pdiffusion >>
rect 413 394 414 395 
<< m1 >>
rect 416 394 417 395 
<< m1 >>
rect 418 394 419 395 
<< pdiffusion >>
rect 426 394 427 395 
<< pdiffusion >>
rect 427 394 428 395 
<< pdiffusion >>
rect 428 394 429 395 
<< pdiffusion >>
rect 429 394 430 395 
<< pdiffusion >>
rect 430 394 431 395 
<< pdiffusion >>
rect 431 394 432 395 
<< m1 >>
rect 433 394 434 395 
<< m1 >>
rect 435 394 436 395 
<< m1 >>
rect 437 394 438 395 
<< pdiffusion >>
rect 444 394 445 395 
<< pdiffusion >>
rect 445 394 446 395 
<< pdiffusion >>
rect 446 394 447 395 
<< pdiffusion >>
rect 447 394 448 395 
<< pdiffusion >>
rect 448 394 449 395 
<< pdiffusion >>
rect 449 394 450 395 
<< m1 >>
rect 451 394 452 395 
<< m1 >>
rect 455 394 456 395 
<< m1 >>
rect 457 394 458 395 
<< pdiffusion >>
rect 462 394 463 395 
<< pdiffusion >>
rect 463 394 464 395 
<< pdiffusion >>
rect 464 394 465 395 
<< pdiffusion >>
rect 465 394 466 395 
<< pdiffusion >>
rect 466 394 467 395 
<< pdiffusion >>
rect 467 394 468 395 
<< m1 >>
rect 472 394 473 395 
<< m1 >>
rect 476 394 477 395 
<< m1 >>
rect 478 394 479 395 
<< pdiffusion >>
rect 480 394 481 395 
<< pdiffusion >>
rect 481 394 482 395 
<< pdiffusion >>
rect 482 394 483 395 
<< pdiffusion >>
rect 483 394 484 395 
<< pdiffusion >>
rect 484 394 485 395 
<< pdiffusion >>
rect 485 394 486 395 
<< pdiffusion >>
rect 498 394 499 395 
<< pdiffusion >>
rect 499 394 500 395 
<< pdiffusion >>
rect 500 394 501 395 
<< pdiffusion >>
rect 501 394 502 395 
<< pdiffusion >>
rect 502 394 503 395 
<< pdiffusion >>
rect 503 394 504 395 
<< pdiffusion >>
rect 516 394 517 395 
<< pdiffusion >>
rect 517 394 518 395 
<< pdiffusion >>
rect 518 394 519 395 
<< pdiffusion >>
rect 519 394 520 395 
<< pdiffusion >>
rect 520 394 521 395 
<< pdiffusion >>
rect 521 394 522 395 
<< m1 >>
rect 523 394 524 395 
<< pdiffusion >>
rect 12 395 13 396 
<< pdiffusion >>
rect 13 395 14 396 
<< pdiffusion >>
rect 14 395 15 396 
<< pdiffusion >>
rect 15 395 16 396 
<< pdiffusion >>
rect 16 395 17 396 
<< pdiffusion >>
rect 17 395 18 396 
<< m1 >>
rect 19 395 20 396 
<< m2 >>
rect 20 395 21 396 
<< m1 >>
rect 23 395 24 396 
<< pdiffusion >>
rect 30 395 31 396 
<< pdiffusion >>
rect 31 395 32 396 
<< pdiffusion >>
rect 32 395 33 396 
<< pdiffusion >>
rect 33 395 34 396 
<< pdiffusion >>
rect 34 395 35 396 
<< pdiffusion >>
rect 35 395 36 396 
<< m1 >>
rect 42 395 43 396 
<< m1 >>
rect 44 395 45 396 
<< pdiffusion >>
rect 48 395 49 396 
<< pdiffusion >>
rect 49 395 50 396 
<< pdiffusion >>
rect 50 395 51 396 
<< pdiffusion >>
rect 51 395 52 396 
<< m1 >>
rect 52 395 53 396 
<< pdiffusion >>
rect 52 395 53 396 
<< pdiffusion >>
rect 53 395 54 396 
<< m2 >>
rect 63 395 64 396 
<< m1 >>
rect 64 395 65 396 
<< pdiffusion >>
rect 66 395 67 396 
<< m1 >>
rect 67 395 68 396 
<< pdiffusion >>
rect 67 395 68 396 
<< pdiffusion >>
rect 68 395 69 396 
<< pdiffusion >>
rect 69 395 70 396 
<< pdiffusion >>
rect 70 395 71 396 
<< pdiffusion >>
rect 71 395 72 396 
<< m1 >>
rect 73 395 74 396 
<< m1 >>
rect 78 395 79 396 
<< m1 >>
rect 82 395 83 396 
<< pdiffusion >>
rect 84 395 85 396 
<< pdiffusion >>
rect 85 395 86 396 
<< pdiffusion >>
rect 86 395 87 396 
<< pdiffusion >>
rect 87 395 88 396 
<< pdiffusion >>
rect 88 395 89 396 
<< pdiffusion >>
rect 89 395 90 396 
<< m1 >>
rect 93 395 94 396 
<< m1 >>
rect 100 395 101 396 
<< pdiffusion >>
rect 102 395 103 396 
<< pdiffusion >>
rect 103 395 104 396 
<< pdiffusion >>
rect 104 395 105 396 
<< pdiffusion >>
rect 105 395 106 396 
<< m1 >>
rect 106 395 107 396 
<< pdiffusion >>
rect 106 395 107 396 
<< pdiffusion >>
rect 107 395 108 396 
<< m1 >>
rect 110 395 111 396 
<< m2 >>
rect 110 395 111 396 
<< m2c >>
rect 110 395 111 396 
<< m1 >>
rect 110 395 111 396 
<< m2 >>
rect 110 395 111 396 
<< m1 >>
rect 112 395 113 396 
<< m1 >>
rect 114 395 115 396 
<< m1 >>
rect 118 395 119 396 
<< pdiffusion >>
rect 120 395 121 396 
<< pdiffusion >>
rect 121 395 122 396 
<< pdiffusion >>
rect 122 395 123 396 
<< pdiffusion >>
rect 123 395 124 396 
<< pdiffusion >>
rect 124 395 125 396 
<< pdiffusion >>
rect 125 395 126 396 
<< m1 >>
rect 127 395 128 396 
<< m2 >>
rect 128 395 129 396 
<< m1 >>
rect 136 395 137 396 
<< pdiffusion >>
rect 138 395 139 396 
<< pdiffusion >>
rect 139 395 140 396 
<< pdiffusion >>
rect 140 395 141 396 
<< pdiffusion >>
rect 141 395 142 396 
<< pdiffusion >>
rect 142 395 143 396 
<< pdiffusion >>
rect 143 395 144 396 
<< m1 >>
rect 150 395 151 396 
<< pdiffusion >>
rect 156 395 157 396 
<< m1 >>
rect 157 395 158 396 
<< pdiffusion >>
rect 157 395 158 396 
<< pdiffusion >>
rect 158 395 159 396 
<< pdiffusion >>
rect 159 395 160 396 
<< m1 >>
rect 160 395 161 396 
<< pdiffusion >>
rect 160 395 161 396 
<< pdiffusion >>
rect 161 395 162 396 
<< m1 >>
rect 163 395 164 396 
<< m2 >>
rect 163 395 164 396 
<< m2 >>
rect 164 395 165 396 
<< m1 >>
rect 165 395 166 396 
<< m2 >>
rect 165 395 166 396 
<< m2c >>
rect 165 395 166 396 
<< m1 >>
rect 165 395 166 396 
<< m2 >>
rect 165 395 166 396 
<< m1 >>
rect 166 395 167 396 
<< m1 >>
rect 167 395 168 396 
<< m2 >>
rect 167 395 168 396 
<< m1 >>
rect 168 395 169 396 
<< m1 >>
rect 169 395 170 396 
<< m2 >>
rect 169 395 170 396 
<< m1 >>
rect 170 395 171 396 
<< m1 >>
rect 171 395 172 396 
<< pdiffusion >>
rect 174 395 175 396 
<< m1 >>
rect 175 395 176 396 
<< pdiffusion >>
rect 175 395 176 396 
<< pdiffusion >>
rect 176 395 177 396 
<< pdiffusion >>
rect 177 395 178 396 
<< pdiffusion >>
rect 178 395 179 396 
<< pdiffusion >>
rect 179 395 180 396 
<< m1 >>
rect 190 395 191 396 
<< pdiffusion >>
rect 192 395 193 396 
<< m1 >>
rect 193 395 194 396 
<< pdiffusion >>
rect 193 395 194 396 
<< pdiffusion >>
rect 194 395 195 396 
<< pdiffusion >>
rect 195 395 196 396 
<< pdiffusion >>
rect 196 395 197 396 
<< pdiffusion >>
rect 197 395 198 396 
<< m1 >>
rect 199 395 200 396 
<< m2 >>
rect 205 395 206 396 
<< m1 >>
rect 206 395 207 396 
<< pdiffusion >>
rect 210 395 211 396 
<< pdiffusion >>
rect 211 395 212 396 
<< pdiffusion >>
rect 212 395 213 396 
<< pdiffusion >>
rect 213 395 214 396 
<< m1 >>
rect 214 395 215 396 
<< pdiffusion >>
rect 214 395 215 396 
<< pdiffusion >>
rect 215 395 216 396 
<< m1 >>
rect 217 395 218 396 
<< m1 >>
rect 223 395 224 396 
<< pdiffusion >>
rect 228 395 229 396 
<< pdiffusion >>
rect 229 395 230 396 
<< pdiffusion >>
rect 230 395 231 396 
<< pdiffusion >>
rect 231 395 232 396 
<< pdiffusion >>
rect 232 395 233 396 
<< pdiffusion >>
rect 233 395 234 396 
<< m1 >>
rect 235 395 236 396 
<< m1 >>
rect 244 395 245 396 
<< pdiffusion >>
rect 246 395 247 396 
<< m1 >>
rect 247 395 248 396 
<< pdiffusion >>
rect 247 395 248 396 
<< pdiffusion >>
rect 248 395 249 396 
<< pdiffusion >>
rect 249 395 250 396 
<< pdiffusion >>
rect 250 395 251 396 
<< pdiffusion >>
rect 251 395 252 396 
<< m1 >>
rect 253 395 254 396 
<< m1 >>
rect 255 395 256 396 
<< m1 >>
rect 259 395 260 396 
<< pdiffusion >>
rect 264 395 265 396 
<< pdiffusion >>
rect 265 395 266 396 
<< pdiffusion >>
rect 266 395 267 396 
<< pdiffusion >>
rect 267 395 268 396 
<< pdiffusion >>
rect 268 395 269 396 
<< pdiffusion >>
rect 269 395 270 396 
<< m1 >>
rect 280 395 281 396 
<< pdiffusion >>
rect 282 395 283 396 
<< pdiffusion >>
rect 283 395 284 396 
<< pdiffusion >>
rect 284 395 285 396 
<< pdiffusion >>
rect 285 395 286 396 
<< pdiffusion >>
rect 286 395 287 396 
<< pdiffusion >>
rect 287 395 288 396 
<< pdiffusion >>
rect 300 395 301 396 
<< m1 >>
rect 301 395 302 396 
<< pdiffusion >>
rect 301 395 302 396 
<< pdiffusion >>
rect 302 395 303 396 
<< pdiffusion >>
rect 303 395 304 396 
<< pdiffusion >>
rect 304 395 305 396 
<< pdiffusion >>
rect 305 395 306 396 
<< m1 >>
rect 307 395 308 396 
<< m1 >>
rect 310 395 311 396 
<< m1 >>
rect 316 395 317 396 
<< pdiffusion >>
rect 318 395 319 396 
<< pdiffusion >>
rect 319 395 320 396 
<< pdiffusion >>
rect 320 395 321 396 
<< pdiffusion >>
rect 321 395 322 396 
<< m1 >>
rect 322 395 323 396 
<< pdiffusion >>
rect 322 395 323 396 
<< pdiffusion >>
rect 323 395 324 396 
<< m1 >>
rect 325 395 326 396 
<< pdiffusion >>
rect 336 395 337 396 
<< pdiffusion >>
rect 337 395 338 396 
<< pdiffusion >>
rect 338 395 339 396 
<< pdiffusion >>
rect 339 395 340 396 
<< pdiffusion >>
rect 340 395 341 396 
<< pdiffusion >>
rect 341 395 342 396 
<< m1 >>
rect 343 395 344 396 
<< pdiffusion >>
rect 354 395 355 396 
<< pdiffusion >>
rect 355 395 356 396 
<< pdiffusion >>
rect 356 395 357 396 
<< pdiffusion >>
rect 357 395 358 396 
<< pdiffusion >>
rect 358 395 359 396 
<< pdiffusion >>
rect 359 395 360 396 
<< m1 >>
rect 361 395 362 396 
<< m1 >>
rect 363 395 364 396 
<< m2 >>
rect 364 395 365 396 
<< m1 >>
rect 367 395 368 396 
<< pdiffusion >>
rect 372 395 373 396 
<< pdiffusion >>
rect 373 395 374 396 
<< pdiffusion >>
rect 374 395 375 396 
<< pdiffusion >>
rect 375 395 376 396 
<< pdiffusion >>
rect 376 395 377 396 
<< pdiffusion >>
rect 377 395 378 396 
<< m1 >>
rect 385 395 386 396 
<< m1 >>
rect 402 395 403 396 
<< m1 >>
rect 406 395 407 396 
<< pdiffusion >>
rect 408 395 409 396 
<< pdiffusion >>
rect 409 395 410 396 
<< pdiffusion >>
rect 410 395 411 396 
<< pdiffusion >>
rect 411 395 412 396 
<< pdiffusion >>
rect 412 395 413 396 
<< pdiffusion >>
rect 413 395 414 396 
<< m1 >>
rect 416 395 417 396 
<< m1 >>
rect 418 395 419 396 
<< pdiffusion >>
rect 426 395 427 396 
<< m1 >>
rect 427 395 428 396 
<< pdiffusion >>
rect 427 395 428 396 
<< pdiffusion >>
rect 428 395 429 396 
<< pdiffusion >>
rect 429 395 430 396 
<< pdiffusion >>
rect 430 395 431 396 
<< pdiffusion >>
rect 431 395 432 396 
<< m1 >>
rect 433 395 434 396 
<< m1 >>
rect 435 395 436 396 
<< m1 >>
rect 437 395 438 396 
<< pdiffusion >>
rect 444 395 445 396 
<< m1 >>
rect 445 395 446 396 
<< pdiffusion >>
rect 445 395 446 396 
<< pdiffusion >>
rect 446 395 447 396 
<< pdiffusion >>
rect 447 395 448 396 
<< m1 >>
rect 448 395 449 396 
<< pdiffusion >>
rect 448 395 449 396 
<< pdiffusion >>
rect 449 395 450 396 
<< m1 >>
rect 451 395 452 396 
<< m1 >>
rect 455 395 456 396 
<< m2 >>
rect 455 395 456 396 
<< m2c >>
rect 455 395 456 396 
<< m1 >>
rect 455 395 456 396 
<< m2 >>
rect 455 395 456 396 
<< m1 >>
rect 457 395 458 396 
<< m2 >>
rect 457 395 458 396 
<< m2c >>
rect 457 395 458 396 
<< m1 >>
rect 457 395 458 396 
<< m2 >>
rect 457 395 458 396 
<< pdiffusion >>
rect 462 395 463 396 
<< m1 >>
rect 463 395 464 396 
<< pdiffusion >>
rect 463 395 464 396 
<< pdiffusion >>
rect 464 395 465 396 
<< pdiffusion >>
rect 465 395 466 396 
<< pdiffusion >>
rect 466 395 467 396 
<< pdiffusion >>
rect 467 395 468 396 
<< m1 >>
rect 472 395 473 396 
<< m1 >>
rect 476 395 477 396 
<< m1 >>
rect 478 395 479 396 
<< pdiffusion >>
rect 480 395 481 396 
<< pdiffusion >>
rect 481 395 482 396 
<< pdiffusion >>
rect 482 395 483 396 
<< pdiffusion >>
rect 483 395 484 396 
<< pdiffusion >>
rect 484 395 485 396 
<< pdiffusion >>
rect 485 395 486 396 
<< pdiffusion >>
rect 498 395 499 396 
<< pdiffusion >>
rect 499 395 500 396 
<< pdiffusion >>
rect 500 395 501 396 
<< pdiffusion >>
rect 501 395 502 396 
<< pdiffusion >>
rect 502 395 503 396 
<< pdiffusion >>
rect 503 395 504 396 
<< pdiffusion >>
rect 516 395 517 396 
<< pdiffusion >>
rect 517 395 518 396 
<< pdiffusion >>
rect 518 395 519 396 
<< pdiffusion >>
rect 519 395 520 396 
<< pdiffusion >>
rect 520 395 521 396 
<< pdiffusion >>
rect 521 395 522 396 
<< m1 >>
rect 523 395 524 396 
<< m1 >>
rect 19 396 20 397 
<< m2 >>
rect 20 396 21 397 
<< m1 >>
rect 23 396 24 397 
<< m1 >>
rect 42 396 43 397 
<< m1 >>
rect 44 396 45 397 
<< m1 >>
rect 52 396 53 397 
<< m2 >>
rect 63 396 64 397 
<< m1 >>
rect 64 396 65 397 
<< m1 >>
rect 67 396 68 397 
<< m1 >>
rect 73 396 74 397 
<< m1 >>
rect 78 396 79 397 
<< m1 >>
rect 82 396 83 397 
<< m1 >>
rect 93 396 94 397 
<< m1 >>
rect 100 396 101 397 
<< m1 >>
rect 106 396 107 397 
<< m2 >>
rect 110 396 111 397 
<< m1 >>
rect 112 396 113 397 
<< m1 >>
rect 114 396 115 397 
<< m1 >>
rect 118 396 119 397 
<< m1 >>
rect 127 396 128 397 
<< m2 >>
rect 128 396 129 397 
<< m1 >>
rect 136 396 137 397 
<< m1 >>
rect 150 396 151 397 
<< m1 >>
rect 157 396 158 397 
<< m1 >>
rect 160 396 161 397 
<< m1 >>
rect 163 396 164 397 
<< m2 >>
rect 163 396 164 397 
<< m2 >>
rect 167 396 168 397 
<< m2 >>
rect 169 396 170 397 
<< m1 >>
rect 175 396 176 397 
<< m1 >>
rect 190 396 191 397 
<< m1 >>
rect 193 396 194 397 
<< m1 >>
rect 199 396 200 397 
<< m2 >>
rect 205 396 206 397 
<< m1 >>
rect 206 396 207 397 
<< m1 >>
rect 214 396 215 397 
<< m1 >>
rect 217 396 218 397 
<< m1 >>
rect 223 396 224 397 
<< m1 >>
rect 235 396 236 397 
<< m1 >>
rect 244 396 245 397 
<< m1 >>
rect 247 396 248 397 
<< m1 >>
rect 253 396 254 397 
<< m1 >>
rect 255 396 256 397 
<< m1 >>
rect 259 396 260 397 
<< m1 >>
rect 280 396 281 397 
<< m1 >>
rect 301 396 302 397 
<< m1 >>
rect 307 396 308 397 
<< m1 >>
rect 310 396 311 397 
<< m1 >>
rect 316 396 317 397 
<< m1 >>
rect 322 396 323 397 
<< m1 >>
rect 325 396 326 397 
<< m1 >>
rect 343 396 344 397 
<< m1 >>
rect 361 396 362 397 
<< m1 >>
rect 363 396 364 397 
<< m2 >>
rect 364 396 365 397 
<< m1 >>
rect 365 396 366 397 
<< m2 >>
rect 365 396 366 397 
<< m2c >>
rect 365 396 366 397 
<< m1 >>
rect 365 396 366 397 
<< m2 >>
rect 365 396 366 397 
<< m2 >>
rect 366 396 367 397 
<< m1 >>
rect 367 396 368 397 
<< m2 >>
rect 367 396 368 397 
<< m2 >>
rect 368 396 369 397 
<< m1 >>
rect 385 396 386 397 
<< m1 >>
rect 402 396 403 397 
<< m1 >>
rect 406 396 407 397 
<< m1 >>
rect 416 396 417 397 
<< m1 >>
rect 418 396 419 397 
<< m1 >>
rect 427 396 428 397 
<< m1 >>
rect 433 396 434 397 
<< m1 >>
rect 435 396 436 397 
<< m1 >>
rect 437 396 438 397 
<< m1 >>
rect 445 396 446 397 
<< m1 >>
rect 448 396 449 397 
<< m1 >>
rect 451 396 452 397 
<< m2 >>
rect 455 396 456 397 
<< m2 >>
rect 457 396 458 397 
<< m1 >>
rect 463 396 464 397 
<< m1 >>
rect 472 396 473 397 
<< m1 >>
rect 476 396 477 397 
<< m1 >>
rect 478 396 479 397 
<< m1 >>
rect 523 396 524 397 
<< m1 >>
rect 19 397 20 398 
<< m2 >>
rect 20 397 21 398 
<< m1 >>
rect 23 397 24 398 
<< m1 >>
rect 42 397 43 398 
<< m1 >>
rect 44 397 45 398 
<< m1 >>
rect 52 397 53 398 
<< m2 >>
rect 63 397 64 398 
<< m1 >>
rect 64 397 65 398 
<< m1 >>
rect 67 397 68 398 
<< m1 >>
rect 73 397 74 398 
<< m1 >>
rect 78 397 79 398 
<< m1 >>
rect 82 397 83 398 
<< m1 >>
rect 93 397 94 398 
<< m1 >>
rect 100 397 101 398 
<< m1 >>
rect 106 397 107 398 
<< m2 >>
rect 107 397 108 398 
<< m1 >>
rect 108 397 109 398 
<< m2 >>
rect 108 397 109 398 
<< m2c >>
rect 108 397 109 398 
<< m1 >>
rect 108 397 109 398 
<< m2 >>
rect 108 397 109 398 
<< m1 >>
rect 109 397 110 398 
<< m1 >>
rect 110 397 111 398 
<< m2 >>
rect 110 397 111 398 
<< m1 >>
rect 111 397 112 398 
<< m1 >>
rect 112 397 113 398 
<< m1 >>
rect 114 397 115 398 
<< m1 >>
rect 118 397 119 398 
<< m1 >>
rect 127 397 128 398 
<< m2 >>
rect 128 397 129 398 
<< m1 >>
rect 136 397 137 398 
<< m1 >>
rect 150 397 151 398 
<< m1 >>
rect 157 397 158 398 
<< m1 >>
rect 160 397 161 398 
<< m1 >>
rect 161 397 162 398 
<< m2 >>
rect 161 397 162 398 
<< m2c >>
rect 161 397 162 398 
<< m1 >>
rect 161 397 162 398 
<< m2 >>
rect 161 397 162 398 
<< m2 >>
rect 162 397 163 398 
<< m1 >>
rect 163 397 164 398 
<< m2 >>
rect 163 397 164 398 
<< m1 >>
rect 164 397 165 398 
<< m1 >>
rect 165 397 166 398 
<< m1 >>
rect 166 397 167 398 
<< m1 >>
rect 167 397 168 398 
<< m2 >>
rect 167 397 168 398 
<< m1 >>
rect 168 397 169 398 
<< m1 >>
rect 169 397 170 398 
<< m2 >>
rect 169 397 170 398 
<< m1 >>
rect 170 397 171 398 
<< m1 >>
rect 171 397 172 398 
<< m1 >>
rect 172 397 173 398 
<< m1 >>
rect 173 397 174 398 
<< m1 >>
rect 174 397 175 398 
<< m1 >>
rect 175 397 176 398 
<< m1 >>
rect 190 397 191 398 
<< m1 >>
rect 191 397 192 398 
<< m1 >>
rect 192 397 193 398 
<< m1 >>
rect 193 397 194 398 
<< m1 >>
rect 199 397 200 398 
<< m2 >>
rect 205 397 206 398 
<< m1 >>
rect 206 397 207 398 
<< m1 >>
rect 214 397 215 398 
<< m1 >>
rect 217 397 218 398 
<< m1 >>
rect 223 397 224 398 
<< m1 >>
rect 235 397 236 398 
<< m1 >>
rect 244 397 245 398 
<< m1 >>
rect 247 397 248 398 
<< m1 >>
rect 253 397 254 398 
<< m1 >>
rect 255 397 256 398 
<< m1 >>
rect 259 397 260 398 
<< m1 >>
rect 280 397 281 398 
<< m1 >>
rect 301 397 302 398 
<< m1 >>
rect 307 397 308 398 
<< m1 >>
rect 310 397 311 398 
<< m1 >>
rect 316 397 317 398 
<< m1 >>
rect 322 397 323 398 
<< m1 >>
rect 325 397 326 398 
<< m1 >>
rect 343 397 344 398 
<< m1 >>
rect 361 397 362 398 
<< m1 >>
rect 363 397 364 398 
<< m1 >>
rect 367 397 368 398 
<< m2 >>
rect 368 397 369 398 
<< m1 >>
rect 385 397 386 398 
<< m1 >>
rect 402 397 403 398 
<< m1 >>
rect 406 397 407 398 
<< m1 >>
rect 416 397 417 398 
<< m1 >>
rect 418 397 419 398 
<< m1 >>
rect 419 397 420 398 
<< m1 >>
rect 420 397 421 398 
<< m1 >>
rect 421 397 422 398 
<< m1 >>
rect 422 397 423 398 
<< m1 >>
rect 423 397 424 398 
<< m1 >>
rect 424 397 425 398 
<< m1 >>
rect 425 397 426 398 
<< m2 >>
rect 425 397 426 398 
<< m2c >>
rect 425 397 426 398 
<< m1 >>
rect 425 397 426 398 
<< m2 >>
rect 425 397 426 398 
<< m2 >>
rect 426 397 427 398 
<< m1 >>
rect 427 397 428 398 
<< m1 >>
rect 433 397 434 398 
<< m1 >>
rect 435 397 436 398 
<< m1 >>
rect 437 397 438 398 
<< m1 >>
rect 438 397 439 398 
<< m1 >>
rect 439 397 440 398 
<< m1 >>
rect 440 397 441 398 
<< m1 >>
rect 441 397 442 398 
<< m1 >>
rect 442 397 443 398 
<< m1 >>
rect 443 397 444 398 
<< m2 >>
rect 443 397 444 398 
<< m2c >>
rect 443 397 444 398 
<< m1 >>
rect 443 397 444 398 
<< m2 >>
rect 443 397 444 398 
<< m2 >>
rect 444 397 445 398 
<< m1 >>
rect 445 397 446 398 
<< m1 >>
rect 448 397 449 398 
<< m1 >>
rect 451 397 452 398 
<< m1 >>
rect 452 397 453 398 
<< m1 >>
rect 453 397 454 398 
<< m1 >>
rect 454 397 455 398 
<< m1 >>
rect 455 397 456 398 
<< m2 >>
rect 455 397 456 398 
<< m1 >>
rect 456 397 457 398 
<< m1 >>
rect 457 397 458 398 
<< m2 >>
rect 457 397 458 398 
<< m1 >>
rect 458 397 459 398 
<< m1 >>
rect 459 397 460 398 
<< m1 >>
rect 460 397 461 398 
<< m1 >>
rect 461 397 462 398 
<< m1 >>
rect 462 397 463 398 
<< m1 >>
rect 463 397 464 398 
<< m1 >>
rect 472 397 473 398 
<< m1 >>
rect 476 397 477 398 
<< m1 >>
rect 478 397 479 398 
<< m1 >>
rect 523 397 524 398 
<< m1 >>
rect 19 398 20 399 
<< m2 >>
rect 20 398 21 399 
<< m1 >>
rect 23 398 24 399 
<< m1 >>
rect 42 398 43 399 
<< m1 >>
rect 44 398 45 399 
<< m1 >>
rect 52 398 53 399 
<< m2 >>
rect 63 398 64 399 
<< m1 >>
rect 64 398 65 399 
<< m1 >>
rect 67 398 68 399 
<< m1 >>
rect 73 398 74 399 
<< m1 >>
rect 78 398 79 399 
<< m1 >>
rect 82 398 83 399 
<< m1 >>
rect 93 398 94 399 
<< m2 >>
rect 93 398 94 399 
<< m2c >>
rect 93 398 94 399 
<< m1 >>
rect 93 398 94 399 
<< m2 >>
rect 93 398 94 399 
<< m1 >>
rect 100 398 101 399 
<< m2 >>
rect 100 398 101 399 
<< m2c >>
rect 100 398 101 399 
<< m1 >>
rect 100 398 101 399 
<< m2 >>
rect 100 398 101 399 
<< m1 >>
rect 104 398 105 399 
<< m2 >>
rect 104 398 105 399 
<< m2c >>
rect 104 398 105 399 
<< m1 >>
rect 104 398 105 399 
<< m2 >>
rect 104 398 105 399 
<< m2 >>
rect 105 398 106 399 
<< m1 >>
rect 106 398 107 399 
<< m2 >>
rect 106 398 107 399 
<< m2 >>
rect 107 398 108 399 
<< m2 >>
rect 110 398 111 399 
<< m1 >>
rect 114 398 115 399 
<< m2 >>
rect 114 398 115 399 
<< m2c >>
rect 114 398 115 399 
<< m1 >>
rect 114 398 115 399 
<< m2 >>
rect 114 398 115 399 
<< m1 >>
rect 118 398 119 399 
<< m2 >>
rect 118 398 119 399 
<< m2c >>
rect 118 398 119 399 
<< m1 >>
rect 118 398 119 399 
<< m2 >>
rect 118 398 119 399 
<< m1 >>
rect 122 398 123 399 
<< m2 >>
rect 122 398 123 399 
<< m2c >>
rect 122 398 123 399 
<< m1 >>
rect 122 398 123 399 
<< m2 >>
rect 122 398 123 399 
<< m1 >>
rect 123 398 124 399 
<< m1 >>
rect 124 398 125 399 
<< m1 >>
rect 125 398 126 399 
<< m1 >>
rect 126 398 127 399 
<< m1 >>
rect 127 398 128 399 
<< m2 >>
rect 128 398 129 399 
<< m1 >>
rect 136 398 137 399 
<< m1 >>
rect 150 398 151 399 
<< m1 >>
rect 157 398 158 399 
<< m2 >>
rect 167 398 168 399 
<< m2 >>
rect 169 398 170 399 
<< m2 >>
rect 194 398 195 399 
<< m1 >>
rect 195 398 196 399 
<< m2 >>
rect 195 398 196 399 
<< m2c >>
rect 195 398 196 399 
<< m1 >>
rect 195 398 196 399 
<< m2 >>
rect 195 398 196 399 
<< m1 >>
rect 196 398 197 399 
<< m1 >>
rect 197 398 198 399 
<< m1 >>
rect 198 398 199 399 
<< m1 >>
rect 199 398 200 399 
<< m2 >>
rect 205 398 206 399 
<< m1 >>
rect 206 398 207 399 
<< m1 >>
rect 214 398 215 399 
<< m1 >>
rect 217 398 218 399 
<< m1 >>
rect 223 398 224 399 
<< m1 >>
rect 235 398 236 399 
<< m1 >>
rect 244 398 245 399 
<< m1 >>
rect 247 398 248 399 
<< m1 >>
rect 253 398 254 399 
<< m1 >>
rect 255 398 256 399 
<< m1 >>
rect 259 398 260 399 
<< m1 >>
rect 280 398 281 399 
<< m1 >>
rect 301 398 302 399 
<< m1 >>
rect 302 398 303 399 
<< m1 >>
rect 303 398 304 399 
<< m1 >>
rect 304 398 305 399 
<< m1 >>
rect 305 398 306 399 
<< m1 >>
rect 306 398 307 399 
<< m1 >>
rect 307 398 308 399 
<< m1 >>
rect 310 398 311 399 
<< m1 >>
rect 316 398 317 399 
<< m1 >>
rect 322 398 323 399 
<< m1 >>
rect 325 398 326 399 
<< m1 >>
rect 343 398 344 399 
<< m1 >>
rect 357 398 358 399 
<< m2 >>
rect 357 398 358 399 
<< m2c >>
rect 357 398 358 399 
<< m1 >>
rect 357 398 358 399 
<< m2 >>
rect 357 398 358 399 
<< m1 >>
rect 358 398 359 399 
<< m1 >>
rect 359 398 360 399 
<< m2 >>
rect 359 398 360 399 
<< m2c >>
rect 359 398 360 399 
<< m1 >>
rect 359 398 360 399 
<< m2 >>
rect 359 398 360 399 
<< m2 >>
rect 360 398 361 399 
<< m1 >>
rect 361 398 362 399 
<< m2 >>
rect 361 398 362 399 
<< m2 >>
rect 362 398 363 399 
<< m1 >>
rect 363 398 364 399 
<< m2 >>
rect 363 398 364 399 
<< m2 >>
rect 364 398 365 399 
<< m1 >>
rect 365 398 366 399 
<< m2 >>
rect 365 398 366 399 
<< m2c >>
rect 365 398 366 399 
<< m1 >>
rect 365 398 366 399 
<< m2 >>
rect 365 398 366 399 
<< m1 >>
rect 366 398 367 399 
<< m1 >>
rect 367 398 368 399 
<< m2 >>
rect 368 398 369 399 
<< m1 >>
rect 385 398 386 399 
<< m1 >>
rect 402 398 403 399 
<< m1 >>
rect 406 398 407 399 
<< m1 >>
rect 416 398 417 399 
<< m2 >>
rect 426 398 427 399 
<< m1 >>
rect 427 398 428 399 
<< m1 >>
rect 433 398 434 399 
<< m1 >>
rect 435 398 436 399 
<< m2 >>
rect 444 398 445 399 
<< m1 >>
rect 445 398 446 399 
<< m2 >>
rect 446 398 447 399 
<< m1 >>
rect 447 398 448 399 
<< m2 >>
rect 447 398 448 399 
<< m2c >>
rect 447 398 448 399 
<< m1 >>
rect 447 398 448 399 
<< m2 >>
rect 447 398 448 399 
<< m1 >>
rect 448 398 449 399 
<< m2 >>
rect 455 398 456 399 
<< m2 >>
rect 457 398 458 399 
<< m1 >>
rect 472 398 473 399 
<< m1 >>
rect 476 398 477 399 
<< m1 >>
rect 478 398 479 399 
<< m1 >>
rect 523 398 524 399 
<< m1 >>
rect 19 399 20 400 
<< m2 >>
rect 20 399 21 400 
<< m1 >>
rect 23 399 24 400 
<< m1 >>
rect 42 399 43 400 
<< m1 >>
rect 44 399 45 400 
<< m1 >>
rect 52 399 53 400 
<< m2 >>
rect 63 399 64 400 
<< m1 >>
rect 64 399 65 400 
<< m1 >>
rect 67 399 68 400 
<< m1 >>
rect 73 399 74 400 
<< m1 >>
rect 78 399 79 400 
<< m1 >>
rect 82 399 83 400 
<< m2 >>
rect 93 399 94 400 
<< m2 >>
rect 99 399 100 400 
<< m2 >>
rect 100 399 101 400 
<< m1 >>
rect 104 399 105 400 
<< m1 >>
rect 106 399 107 400 
<< m2 >>
rect 110 399 111 400 
<< m2 >>
rect 114 399 115 400 
<< m2 >>
rect 118 399 119 400 
<< m2 >>
rect 122 399 123 400 
<< m2 >>
rect 128 399 129 400 
<< m1 >>
rect 136 399 137 400 
<< m1 >>
rect 150 399 151 400 
<< m1 >>
rect 157 399 158 400 
<< m2 >>
rect 158 399 159 400 
<< m1 >>
rect 159 399 160 400 
<< m2 >>
rect 159 399 160 400 
<< m2c >>
rect 159 399 160 400 
<< m1 >>
rect 159 399 160 400 
<< m2 >>
rect 159 399 160 400 
<< m1 >>
rect 160 399 161 400 
<< m1 >>
rect 161 399 162 400 
<< m1 >>
rect 162 399 163 400 
<< m1 >>
rect 163 399 164 400 
<< m1 >>
rect 164 399 165 400 
<< m1 >>
rect 165 399 166 400 
<< m1 >>
rect 166 399 167 400 
<< m1 >>
rect 167 399 168 400 
<< m2 >>
rect 167 399 168 400 
<< m1 >>
rect 168 399 169 400 
<< m1 >>
rect 169 399 170 400 
<< m2 >>
rect 169 399 170 400 
<< m2c >>
rect 169 399 170 400 
<< m1 >>
rect 169 399 170 400 
<< m2 >>
rect 169 399 170 400 
<< m2 >>
rect 194 399 195 400 
<< m2 >>
rect 205 399 206 400 
<< m1 >>
rect 206 399 207 400 
<< m1 >>
rect 214 399 215 400 
<< m1 >>
rect 217 399 218 400 
<< m1 >>
rect 223 399 224 400 
<< m1 >>
rect 235 399 236 400 
<< m1 >>
rect 244 399 245 400 
<< m1 >>
rect 245 399 246 400 
<< m2 >>
rect 245 399 246 400 
<< m2c >>
rect 245 399 246 400 
<< m1 >>
rect 245 399 246 400 
<< m2 >>
rect 245 399 246 400 
<< m2 >>
rect 246 399 247 400 
<< m1 >>
rect 247 399 248 400 
<< m1 >>
rect 253 399 254 400 
<< m1 >>
rect 255 399 256 400 
<< m1 >>
rect 259 399 260 400 
<< m2 >>
rect 259 399 260 400 
<< m2c >>
rect 259 399 260 400 
<< m1 >>
rect 259 399 260 400 
<< m2 >>
rect 259 399 260 400 
<< m1 >>
rect 280 399 281 400 
<< m1 >>
rect 310 399 311 400 
<< m1 >>
rect 316 399 317 400 
<< m1 >>
rect 322 399 323 400 
<< m1 >>
rect 325 399 326 400 
<< m1 >>
rect 343 399 344 400 
<< m2 >>
rect 357 399 358 400 
<< m1 >>
rect 361 399 362 400 
<< m1 >>
rect 363 399 364 400 
<< m2 >>
rect 368 399 369 400 
<< m1 >>
rect 385 399 386 400 
<< m1 >>
rect 402 399 403 400 
<< m1 >>
rect 406 399 407 400 
<< m1 >>
rect 416 399 417 400 
<< m2 >>
rect 426 399 427 400 
<< m1 >>
rect 427 399 428 400 
<< m1 >>
rect 433 399 434 400 
<< m1 >>
rect 435 399 436 400 
<< m2 >>
rect 444 399 445 400 
<< m1 >>
rect 445 399 446 400 
<< m2 >>
rect 446 399 447 400 
<< m2 >>
rect 455 399 456 400 
<< m2 >>
rect 457 399 458 400 
<< m1 >>
rect 472 399 473 400 
<< m1 >>
rect 476 399 477 400 
<< m1 >>
rect 478 399 479 400 
<< m1 >>
rect 523 399 524 400 
<< m1 >>
rect 19 400 20 401 
<< m2 >>
rect 20 400 21 401 
<< m1 >>
rect 23 400 24 401 
<< m1 >>
rect 26 400 27 401 
<< m1 >>
rect 27 400 28 401 
<< m1 >>
rect 28 400 29 401 
<< m1 >>
rect 29 400 30 401 
<< m1 >>
rect 30 400 31 401 
<< m1 >>
rect 31 400 32 401 
<< m1 >>
rect 32 400 33 401 
<< m1 >>
rect 33 400 34 401 
<< m1 >>
rect 34 400 35 401 
<< m1 >>
rect 35 400 36 401 
<< m1 >>
rect 36 400 37 401 
<< m1 >>
rect 37 400 38 401 
<< m1 >>
rect 38 400 39 401 
<< m1 >>
rect 39 400 40 401 
<< m1 >>
rect 40 400 41 401 
<< m1 >>
rect 41 400 42 401 
<< m1 >>
rect 42 400 43 401 
<< m1 >>
rect 44 400 45 401 
<< m1 >>
rect 52 400 53 401 
<< m2 >>
rect 63 400 64 401 
<< m1 >>
rect 64 400 65 401 
<< m1 >>
rect 67 400 68 401 
<< m1 >>
rect 68 400 69 401 
<< m1 >>
rect 69 400 70 401 
<< m1 >>
rect 70 400 71 401 
<< m1 >>
rect 71 400 72 401 
<< m2 >>
rect 71 400 72 401 
<< m2c >>
rect 71 400 72 401 
<< m1 >>
rect 71 400 72 401 
<< m2 >>
rect 71 400 72 401 
<< m2 >>
rect 72 400 73 401 
<< m1 >>
rect 73 400 74 401 
<< m2 >>
rect 73 400 74 401 
<< m2 >>
rect 74 400 75 401 
<< m1 >>
rect 75 400 76 401 
<< m2 >>
rect 75 400 76 401 
<< m1 >>
rect 76 400 77 401 
<< m2 >>
rect 76 400 77 401 
<< m2c >>
rect 76 400 77 401 
<< m1 >>
rect 76 400 77 401 
<< m2 >>
rect 76 400 77 401 
<< m2 >>
rect 77 400 78 401 
<< m1 >>
rect 78 400 79 401 
<< m2 >>
rect 78 400 79 401 
<< m2 >>
rect 79 400 80 401 
<< m1 >>
rect 80 400 81 401 
<< m2 >>
rect 80 400 81 401 
<< m2c >>
rect 80 400 81 401 
<< m1 >>
rect 80 400 81 401 
<< m2 >>
rect 80 400 81 401 
<< m2 >>
rect 81 400 82 401 
<< m1 >>
rect 82 400 83 401 
<< m2 >>
rect 82 400 83 401 
<< m2 >>
rect 83 400 84 401 
<< m1 >>
rect 84 400 85 401 
<< m2 >>
rect 84 400 85 401 
<< m2c >>
rect 84 400 85 401 
<< m1 >>
rect 84 400 85 401 
<< m2 >>
rect 84 400 85 401 
<< m1 >>
rect 85 400 86 401 
<< m1 >>
rect 86 400 87 401 
<< m1 >>
rect 87 400 88 401 
<< m1 >>
rect 88 400 89 401 
<< m1 >>
rect 89 400 90 401 
<< m1 >>
rect 90 400 91 401 
<< m1 >>
rect 91 400 92 401 
<< m1 >>
rect 92 400 93 401 
<< m1 >>
rect 93 400 94 401 
<< m2 >>
rect 93 400 94 401 
<< m1 >>
rect 94 400 95 401 
<< m1 >>
rect 95 400 96 401 
<< m1 >>
rect 96 400 97 401 
<< m1 >>
rect 97 400 98 401 
<< m1 >>
rect 98 400 99 401 
<< m1 >>
rect 99 400 100 401 
<< m2 >>
rect 99 400 100 401 
<< m1 >>
rect 100 400 101 401 
<< m1 >>
rect 101 400 102 401 
<< m1 >>
rect 102 400 103 401 
<< m1 >>
rect 103 400 104 401 
<< m1 >>
rect 104 400 105 401 
<< m1 >>
rect 106 400 107 401 
<< m1 >>
rect 107 400 108 401 
<< m1 >>
rect 108 400 109 401 
<< m1 >>
rect 109 400 110 401 
<< m1 >>
rect 110 400 111 401 
<< m2 >>
rect 110 400 111 401 
<< m1 >>
rect 111 400 112 401 
<< m1 >>
rect 112 400 113 401 
<< m1 >>
rect 113 400 114 401 
<< m1 >>
rect 114 400 115 401 
<< m2 >>
rect 114 400 115 401 
<< m1 >>
rect 115 400 116 401 
<< m1 >>
rect 116 400 117 401 
<< m1 >>
rect 117 400 118 401 
<< m1 >>
rect 118 400 119 401 
<< m2 >>
rect 118 400 119 401 
<< m1 >>
rect 119 400 120 401 
<< m1 >>
rect 120 400 121 401 
<< m1 >>
rect 121 400 122 401 
<< m1 >>
rect 122 400 123 401 
<< m2 >>
rect 122 400 123 401 
<< m1 >>
rect 123 400 124 401 
<< m1 >>
rect 124 400 125 401 
<< m1 >>
rect 125 400 126 401 
<< m1 >>
rect 126 400 127 401 
<< m1 >>
rect 127 400 128 401 
<< m1 >>
rect 128 400 129 401 
<< m2 >>
rect 128 400 129 401 
<< m1 >>
rect 129 400 130 401 
<< m1 >>
rect 130 400 131 401 
<< m1 >>
rect 131 400 132 401 
<< m1 >>
rect 132 400 133 401 
<< m1 >>
rect 133 400 134 401 
<< m1 >>
rect 134 400 135 401 
<< m1 >>
rect 135 400 136 401 
<< m1 >>
rect 136 400 137 401 
<< m1 >>
rect 148 400 149 401 
<< m2 >>
rect 148 400 149 401 
<< m2c >>
rect 148 400 149 401 
<< m1 >>
rect 148 400 149 401 
<< m2 >>
rect 148 400 149 401 
<< m2 >>
rect 149 400 150 401 
<< m1 >>
rect 150 400 151 401 
<< m2 >>
rect 150 400 151 401 
<< m2 >>
rect 151 400 152 401 
<< m1 >>
rect 152 400 153 401 
<< m2 >>
rect 152 400 153 401 
<< m2c >>
rect 152 400 153 401 
<< m1 >>
rect 152 400 153 401 
<< m2 >>
rect 152 400 153 401 
<< m1 >>
rect 153 400 154 401 
<< m1 >>
rect 154 400 155 401 
<< m1 >>
rect 155 400 156 401 
<< m2 >>
rect 155 400 156 401 
<< m2c >>
rect 155 400 156 401 
<< m1 >>
rect 155 400 156 401 
<< m2 >>
rect 155 400 156 401 
<< m2 >>
rect 156 400 157 401 
<< m1 >>
rect 157 400 158 401 
<< m2 >>
rect 157 400 158 401 
<< m2 >>
rect 158 400 159 401 
<< m2 >>
rect 167 400 168 401 
<< m1 >>
rect 178 400 179 401 
<< m1 >>
rect 179 400 180 401 
<< m1 >>
rect 180 400 181 401 
<< m1 >>
rect 181 400 182 401 
<< m1 >>
rect 182 400 183 401 
<< m1 >>
rect 183 400 184 401 
<< m1 >>
rect 184 400 185 401 
<< m1 >>
rect 185 400 186 401 
<< m1 >>
rect 186 400 187 401 
<< m1 >>
rect 187 400 188 401 
<< m1 >>
rect 188 400 189 401 
<< m1 >>
rect 189 400 190 401 
<< m1 >>
rect 190 400 191 401 
<< m1 >>
rect 191 400 192 401 
<< m1 >>
rect 192 400 193 401 
<< m1 >>
rect 193 400 194 401 
<< m1 >>
rect 194 400 195 401 
<< m2 >>
rect 194 400 195 401 
<< m1 >>
rect 195 400 196 401 
<< m1 >>
rect 196 400 197 401 
<< m1 >>
rect 197 400 198 401 
<< m1 >>
rect 198 400 199 401 
<< m1 >>
rect 199 400 200 401 
<< m1 >>
rect 200 400 201 401 
<< m1 >>
rect 201 400 202 401 
<< m1 >>
rect 202 400 203 401 
<< m1 >>
rect 203 400 204 401 
<< m1 >>
rect 204 400 205 401 
<< m1 >>
rect 205 400 206 401 
<< m2 >>
rect 205 400 206 401 
<< m1 >>
rect 206 400 207 401 
<< m1 >>
rect 208 400 209 401 
<< m1 >>
rect 209 400 210 401 
<< m1 >>
rect 210 400 211 401 
<< m1 >>
rect 211 400 212 401 
<< m1 >>
rect 212 400 213 401 
<< m1 >>
rect 213 400 214 401 
<< m1 >>
rect 214 400 215 401 
<< m1 >>
rect 217 400 218 401 
<< m1 >>
rect 223 400 224 401 
<< m1 >>
rect 235 400 236 401 
<< m2 >>
rect 246 400 247 401 
<< m1 >>
rect 247 400 248 401 
<< m1 >>
rect 253 400 254 401 
<< m1 >>
rect 255 400 256 401 
<< m2 >>
rect 259 400 260 401 
<< m2 >>
rect 260 400 261 401 
<< m2 >>
rect 261 400 262 401 
<< m2 >>
rect 262 400 263 401 
<< m2 >>
rect 263 400 264 401 
<< m2 >>
rect 264 400 265 401 
<< m2 >>
rect 265 400 266 401 
<< m2 >>
rect 266 400 267 401 
<< m2 >>
rect 267 400 268 401 
<< m2 >>
rect 268 400 269 401 
<< m2 >>
rect 269 400 270 401 
<< m2 >>
rect 270 400 271 401 
<< m2 >>
rect 271 400 272 401 
<< m2 >>
rect 272 400 273 401 
<< m2 >>
rect 273 400 274 401 
<< m2 >>
rect 274 400 275 401 
<< m2 >>
rect 275 400 276 401 
<< m2 >>
rect 276 400 277 401 
<< m2 >>
rect 277 400 278 401 
<< m2 >>
rect 278 400 279 401 
<< m2 >>
rect 279 400 280 401 
<< m1 >>
rect 280 400 281 401 
<< m2 >>
rect 280 400 281 401 
<< m2 >>
rect 281 400 282 401 
<< m1 >>
rect 282 400 283 401 
<< m2 >>
rect 282 400 283 401 
<< m2c >>
rect 282 400 283 401 
<< m1 >>
rect 282 400 283 401 
<< m2 >>
rect 282 400 283 401 
<< m1 >>
rect 283 400 284 401 
<< m1 >>
rect 284 400 285 401 
<< m1 >>
rect 310 400 311 401 
<< m1 >>
rect 314 400 315 401 
<< m2 >>
rect 314 400 315 401 
<< m2c >>
rect 314 400 315 401 
<< m1 >>
rect 314 400 315 401 
<< m2 >>
rect 314 400 315 401 
<< m2 >>
rect 315 400 316 401 
<< m1 >>
rect 316 400 317 401 
<< m2 >>
rect 316 400 317 401 
<< m2 >>
rect 317 400 318 401 
<< m1 >>
rect 318 400 319 401 
<< m2 >>
rect 318 400 319 401 
<< m2c >>
rect 318 400 319 401 
<< m1 >>
rect 318 400 319 401 
<< m2 >>
rect 318 400 319 401 
<< m1 >>
rect 319 400 320 401 
<< m1 >>
rect 320 400 321 401 
<< m1 >>
rect 321 400 322 401 
<< m1 >>
rect 322 400 323 401 
<< m1 >>
rect 325 400 326 401 
<< m1 >>
rect 343 400 344 401 
<< m1 >>
rect 344 400 345 401 
<< m1 >>
rect 345 400 346 401 
<< m1 >>
rect 346 400 347 401 
<< m1 >>
rect 347 400 348 401 
<< m1 >>
rect 348 400 349 401 
<< m1 >>
rect 349 400 350 401 
<< m1 >>
rect 350 400 351 401 
<< m1 >>
rect 351 400 352 401 
<< m1 >>
rect 352 400 353 401 
<< m1 >>
rect 353 400 354 401 
<< m1 >>
rect 354 400 355 401 
<< m1 >>
rect 355 400 356 401 
<< m1 >>
rect 356 400 357 401 
<< m1 >>
rect 357 400 358 401 
<< m2 >>
rect 357 400 358 401 
<< m1 >>
rect 358 400 359 401 
<< m1 >>
rect 359 400 360 401 
<< m2 >>
rect 359 400 360 401 
<< m2c >>
rect 359 400 360 401 
<< m1 >>
rect 359 400 360 401 
<< m2 >>
rect 359 400 360 401 
<< m2 >>
rect 360 400 361 401 
<< m1 >>
rect 361 400 362 401 
<< m2 >>
rect 361 400 362 401 
<< m2 >>
rect 362 400 363 401 
<< m1 >>
rect 363 400 364 401 
<< m2 >>
rect 363 400 364 401 
<< m2 >>
rect 364 400 365 401 
<< m1 >>
rect 365 400 366 401 
<< m2 >>
rect 365 400 366 401 
<< m2c >>
rect 365 400 366 401 
<< m1 >>
rect 365 400 366 401 
<< m2 >>
rect 365 400 366 401 
<< m1 >>
rect 366 400 367 401 
<< m1 >>
rect 367 400 368 401 
<< m1 >>
rect 368 400 369 401 
<< m2 >>
rect 368 400 369 401 
<< m1 >>
rect 369 400 370 401 
<< m1 >>
rect 370 400 371 401 
<< m1 >>
rect 371 400 372 401 
<< m1 >>
rect 372 400 373 401 
<< m1 >>
rect 373 400 374 401 
<< m1 >>
rect 374 400 375 401 
<< m1 >>
rect 375 400 376 401 
<< m1 >>
rect 376 400 377 401 
<< m1 >>
rect 377 400 378 401 
<< m1 >>
rect 378 400 379 401 
<< m1 >>
rect 379 400 380 401 
<< m1 >>
rect 385 400 386 401 
<< m1 >>
rect 402 400 403 401 
<< m1 >>
rect 406 400 407 401 
<< m1 >>
rect 416 400 417 401 
<< m2 >>
rect 426 400 427 401 
<< m1 >>
rect 427 400 428 401 
<< m2 >>
rect 427 400 428 401 
<< m2 >>
rect 428 400 429 401 
<< m1 >>
rect 429 400 430 401 
<< m2 >>
rect 429 400 430 401 
<< m2c >>
rect 429 400 430 401 
<< m1 >>
rect 429 400 430 401 
<< m2 >>
rect 429 400 430 401 
<< m1 >>
rect 430 400 431 401 
<< m1 >>
rect 431 400 432 401 
<< m2 >>
rect 431 400 432 401 
<< m2c >>
rect 431 400 432 401 
<< m1 >>
rect 431 400 432 401 
<< m2 >>
rect 431 400 432 401 
<< m2 >>
rect 432 400 433 401 
<< m1 >>
rect 433 400 434 401 
<< m2 >>
rect 433 400 434 401 
<< m2 >>
rect 434 400 435 401 
<< m1 >>
rect 435 400 436 401 
<< m2 >>
rect 435 400 436 401 
<< m2 >>
rect 436 400 437 401 
<< m1 >>
rect 437 400 438 401 
<< m2 >>
rect 437 400 438 401 
<< m2c >>
rect 437 400 438 401 
<< m1 >>
rect 437 400 438 401 
<< m2 >>
rect 437 400 438 401 
<< m1 >>
rect 438 400 439 401 
<< m1 >>
rect 439 400 440 401 
<< m2 >>
rect 444 400 445 401 
<< m1 >>
rect 445 400 446 401 
<< m2 >>
rect 445 400 446 401 
<< m1 >>
rect 446 400 447 401 
<< m2 >>
rect 446 400 447 401 
<< m1 >>
rect 447 400 448 401 
<< m1 >>
rect 448 400 449 401 
<< m1 >>
rect 449 400 450 401 
<< m1 >>
rect 450 400 451 401 
<< m1 >>
rect 451 400 452 401 
<< m1 >>
rect 452 400 453 401 
<< m1 >>
rect 453 400 454 401 
<< m1 >>
rect 454 400 455 401 
<< m1 >>
rect 455 400 456 401 
<< m2 >>
rect 455 400 456 401 
<< m1 >>
rect 456 400 457 401 
<< m1 >>
rect 457 400 458 401 
<< m2 >>
rect 457 400 458 401 
<< m1 >>
rect 458 400 459 401 
<< m2 >>
rect 458 400 459 401 
<< m1 >>
rect 459 400 460 401 
<< m2 >>
rect 459 400 460 401 
<< m1 >>
rect 460 400 461 401 
<< m2 >>
rect 460 400 461 401 
<< m1 >>
rect 461 400 462 401 
<< m2 >>
rect 461 400 462 401 
<< m1 >>
rect 462 400 463 401 
<< m2 >>
rect 462 400 463 401 
<< m1 >>
rect 463 400 464 401 
<< m2 >>
rect 463 400 464 401 
<< m1 >>
rect 464 400 465 401 
<< m2 >>
rect 464 400 465 401 
<< m1 >>
rect 465 400 466 401 
<< m1 >>
rect 466 400 467 401 
<< m1 >>
rect 467 400 468 401 
<< m1 >>
rect 468 400 469 401 
<< m1 >>
rect 469 400 470 401 
<< m1 >>
rect 470 400 471 401 
<< m1 >>
rect 472 400 473 401 
<< m1 >>
rect 476 400 477 401 
<< m2 >>
rect 476 400 477 401 
<< m2c >>
rect 476 400 477 401 
<< m1 >>
rect 476 400 477 401 
<< m2 >>
rect 476 400 477 401 
<< m1 >>
rect 478 400 479 401 
<< m1 >>
rect 479 400 480 401 
<< m1 >>
rect 480 400 481 401 
<< m1 >>
rect 481 400 482 401 
<< m2 >>
rect 481 400 482 401 
<< m2c >>
rect 481 400 482 401 
<< m1 >>
rect 481 400 482 401 
<< m2 >>
rect 481 400 482 401 
<< m1 >>
rect 523 400 524 401 
<< m1 >>
rect 19 401 20 402 
<< m2 >>
rect 20 401 21 402 
<< m1 >>
rect 23 401 24 402 
<< m1 >>
rect 26 401 27 402 
<< m1 >>
rect 44 401 45 402 
<< m2 >>
rect 44 401 45 402 
<< m2c >>
rect 44 401 45 402 
<< m1 >>
rect 44 401 45 402 
<< m2 >>
rect 44 401 45 402 
<< m1 >>
rect 52 401 53 402 
<< m2 >>
rect 63 401 64 402 
<< m1 >>
rect 64 401 65 402 
<< m1 >>
rect 73 401 74 402 
<< m1 >>
rect 78 401 79 402 
<< m1 >>
rect 82 401 83 402 
<< m2 >>
rect 93 401 94 402 
<< m2 >>
rect 99 401 100 402 
<< m2 >>
rect 110 401 111 402 
<< m2 >>
rect 114 401 115 402 
<< m2 >>
rect 118 401 119 402 
<< m2 >>
rect 121 401 122 402 
<< m2 >>
rect 122 401 123 402 
<< m2 >>
rect 128 401 129 402 
<< m2 >>
rect 129 401 130 402 
<< m2 >>
rect 130 401 131 402 
<< m2 >>
rect 131 401 132 402 
<< m2 >>
rect 132 401 133 402 
<< m2 >>
rect 133 401 134 402 
<< m2 >>
rect 134 401 135 402 
<< m2 >>
rect 135 401 136 402 
<< m2 >>
rect 136 401 137 402 
<< m2 >>
rect 137 401 138 402 
<< m2 >>
rect 138 401 139 402 
<< m2 >>
rect 139 401 140 402 
<< m2 >>
rect 140 401 141 402 
<< m2 >>
rect 141 401 142 402 
<< m2 >>
rect 142 401 143 402 
<< m2 >>
rect 143 401 144 402 
<< m2 >>
rect 144 401 145 402 
<< m2 >>
rect 145 401 146 402 
<< m2 >>
rect 146 401 147 402 
<< m1 >>
rect 148 401 149 402 
<< m1 >>
rect 150 401 151 402 
<< m1 >>
rect 157 401 158 402 
<< m1 >>
rect 167 401 168 402 
<< m2 >>
rect 167 401 168 402 
<< m2c >>
rect 167 401 168 402 
<< m1 >>
rect 167 401 168 402 
<< m2 >>
rect 167 401 168 402 
<< m2 >>
rect 177 401 178 402 
<< m1 >>
rect 178 401 179 402 
<< m2 >>
rect 178 401 179 402 
<< m2 >>
rect 179 401 180 402 
<< m2 >>
rect 180 401 181 402 
<< m2 >>
rect 181 401 182 402 
<< m2 >>
rect 182 401 183 402 
<< m2 >>
rect 183 401 184 402 
<< m2 >>
rect 184 401 185 402 
<< m2 >>
rect 185 401 186 402 
<< m2 >>
rect 186 401 187 402 
<< m2 >>
rect 187 401 188 402 
<< m2 >>
rect 188 401 189 402 
<< m2 >>
rect 189 401 190 402 
<< m2 >>
rect 190 401 191 402 
<< m2 >>
rect 191 401 192 402 
<< m2 >>
rect 192 401 193 402 
<< m2 >>
rect 193 401 194 402 
<< m2 >>
rect 194 401 195 402 
<< m2 >>
rect 196 401 197 402 
<< m2 >>
rect 197 401 198 402 
<< m2 >>
rect 198 401 199 402 
<< m2 >>
rect 199 401 200 402 
<< m2 >>
rect 200 401 201 402 
<< m2 >>
rect 201 401 202 402 
<< m2 >>
rect 202 401 203 402 
<< m2 >>
rect 203 401 204 402 
<< m2 >>
rect 204 401 205 402 
<< m2 >>
rect 205 401 206 402 
<< m2 >>
rect 207 401 208 402 
<< m1 >>
rect 208 401 209 402 
<< m2 >>
rect 208 401 209 402 
<< m2 >>
rect 209 401 210 402 
<< m2 >>
rect 210 401 211 402 
<< m2 >>
rect 211 401 212 402 
<< m2 >>
rect 212 401 213 402 
<< m2 >>
rect 213 401 214 402 
<< m2 >>
rect 214 401 215 402 
<< m2 >>
rect 215 401 216 402 
<< m1 >>
rect 216 401 217 402 
<< m2 >>
rect 216 401 217 402 
<< m2c >>
rect 216 401 217 402 
<< m1 >>
rect 216 401 217 402 
<< m2 >>
rect 216 401 217 402 
<< m1 >>
rect 217 401 218 402 
<< m2 >>
rect 218 401 219 402 
<< m1 >>
rect 219 401 220 402 
<< m2 >>
rect 219 401 220 402 
<< m2c >>
rect 219 401 220 402 
<< m1 >>
rect 219 401 220 402 
<< m2 >>
rect 219 401 220 402 
<< m1 >>
rect 220 401 221 402 
<< m1 >>
rect 221 401 222 402 
<< m1 >>
rect 222 401 223 402 
<< m1 >>
rect 223 401 224 402 
<< m2 >>
rect 234 401 235 402 
<< m1 >>
rect 235 401 236 402 
<< m2 >>
rect 235 401 236 402 
<< m2 >>
rect 236 401 237 402 
<< m1 >>
rect 237 401 238 402 
<< m2 >>
rect 237 401 238 402 
<< m2c >>
rect 237 401 238 402 
<< m1 >>
rect 237 401 238 402 
<< m2 >>
rect 237 401 238 402 
<< m1 >>
rect 238 401 239 402 
<< m1 >>
rect 239 401 240 402 
<< m1 >>
rect 240 401 241 402 
<< m1 >>
rect 241 401 242 402 
<< m1 >>
rect 242 401 243 402 
<< m1 >>
rect 243 401 244 402 
<< m1 >>
rect 244 401 245 402 
<< m1 >>
rect 245 401 246 402 
<< m1 >>
rect 246 401 247 402 
<< m2 >>
rect 246 401 247 402 
<< m1 >>
rect 247 401 248 402 
<< m2 >>
rect 247 401 248 402 
<< m2 >>
rect 248 401 249 402 
<< m1 >>
rect 249 401 250 402 
<< m2 >>
rect 249 401 250 402 
<< m2c >>
rect 249 401 250 402 
<< m1 >>
rect 249 401 250 402 
<< m2 >>
rect 249 401 250 402 
<< m1 >>
rect 250 401 251 402 
<< m1 >>
rect 251 401 252 402 
<< m2 >>
rect 251 401 252 402 
<< m2c >>
rect 251 401 252 402 
<< m1 >>
rect 251 401 252 402 
<< m2 >>
rect 251 401 252 402 
<< m2 >>
rect 252 401 253 402 
<< m1 >>
rect 253 401 254 402 
<< m2 >>
rect 253 401 254 402 
<< m2 >>
rect 254 401 255 402 
<< m1 >>
rect 255 401 256 402 
<< m2 >>
rect 255 401 256 402 
<< m2 >>
rect 256 401 257 402 
<< m1 >>
rect 257 401 258 402 
<< m2 >>
rect 257 401 258 402 
<< m2c >>
rect 257 401 258 402 
<< m1 >>
rect 257 401 258 402 
<< m2 >>
rect 257 401 258 402 
<< m1 >>
rect 258 401 259 402 
<< m1 >>
rect 259 401 260 402 
<< m1 >>
rect 260 401 261 402 
<< m1 >>
rect 261 401 262 402 
<< m1 >>
rect 262 401 263 402 
<< m1 >>
rect 263 401 264 402 
<< m1 >>
rect 264 401 265 402 
<< m1 >>
rect 265 401 266 402 
<< m1 >>
rect 266 401 267 402 
<< m1 >>
rect 267 401 268 402 
<< m1 >>
rect 268 401 269 402 
<< m1 >>
rect 269 401 270 402 
<< m1 >>
rect 270 401 271 402 
<< m1 >>
rect 271 401 272 402 
<< m1 >>
rect 272 401 273 402 
<< m1 >>
rect 273 401 274 402 
<< m1 >>
rect 274 401 275 402 
<< m1 >>
rect 275 401 276 402 
<< m1 >>
rect 276 401 277 402 
<< m1 >>
rect 277 401 278 402 
<< m1 >>
rect 278 401 279 402 
<< m1 >>
rect 280 401 281 402 
<< m1 >>
rect 284 401 285 402 
<< m2 >>
rect 284 401 285 402 
<< m2c >>
rect 284 401 285 402 
<< m1 >>
rect 284 401 285 402 
<< m2 >>
rect 284 401 285 402 
<< m1 >>
rect 310 401 311 402 
<< m2 >>
rect 310 401 311 402 
<< m2c >>
rect 310 401 311 402 
<< m1 >>
rect 310 401 311 402 
<< m2 >>
rect 310 401 311 402 
<< m1 >>
rect 314 401 315 402 
<< m1 >>
rect 316 401 317 402 
<< m1 >>
rect 325 401 326 402 
<< m2 >>
rect 357 401 358 402 
<< m1 >>
rect 361 401 362 402 
<< m1 >>
rect 363 401 364 402 
<< m2 >>
rect 368 401 369 402 
<< m2 >>
rect 369 401 370 402 
<< m2 >>
rect 370 401 371 402 
<< m2 >>
rect 371 401 372 402 
<< m2 >>
rect 372 401 373 402 
<< m2 >>
rect 373 401 374 402 
<< m2 >>
rect 374 401 375 402 
<< m2 >>
rect 375 401 376 402 
<< m2 >>
rect 376 401 377 402 
<< m2 >>
rect 377 401 378 402 
<< m2 >>
rect 378 401 379 402 
<< m1 >>
rect 379 401 380 402 
<< m2 >>
rect 379 401 380 402 
<< m2 >>
rect 380 401 381 402 
<< m1 >>
rect 381 401 382 402 
<< m2 >>
rect 381 401 382 402 
<< m2c >>
rect 381 401 382 402 
<< m1 >>
rect 381 401 382 402 
<< m2 >>
rect 381 401 382 402 
<< m1 >>
rect 382 401 383 402 
<< m1 >>
rect 383 401 384 402 
<< m2 >>
rect 383 401 384 402 
<< m2c >>
rect 383 401 384 402 
<< m1 >>
rect 383 401 384 402 
<< m2 >>
rect 383 401 384 402 
<< m1 >>
rect 385 401 386 402 
<< m2 >>
rect 385 401 386 402 
<< m2c >>
rect 385 401 386 402 
<< m1 >>
rect 385 401 386 402 
<< m2 >>
rect 385 401 386 402 
<< m1 >>
rect 402 401 403 402 
<< m2 >>
rect 402 401 403 402 
<< m2c >>
rect 402 401 403 402 
<< m1 >>
rect 402 401 403 402 
<< m2 >>
rect 402 401 403 402 
<< m1 >>
rect 406 401 407 402 
<< m1 >>
rect 416 401 417 402 
<< m1 >>
rect 427 401 428 402 
<< m1 >>
rect 433 401 434 402 
<< m1 >>
rect 435 401 436 402 
<< m1 >>
rect 439 401 440 402 
<< m2 >>
rect 439 401 440 402 
<< m2c >>
rect 439 401 440 402 
<< m1 >>
rect 439 401 440 402 
<< m2 >>
rect 439 401 440 402 
<< m2 >>
rect 455 401 456 402 
<< m2 >>
rect 464 401 465 402 
<< m1 >>
rect 470 401 471 402 
<< m1 >>
rect 472 401 473 402 
<< m2 >>
rect 476 401 477 402 
<< m2 >>
rect 481 401 482 402 
<< m2 >>
rect 490 401 491 402 
<< m1 >>
rect 491 401 492 402 
<< m2 >>
rect 491 401 492 402 
<< m2c >>
rect 491 401 492 402 
<< m1 >>
rect 491 401 492 402 
<< m2 >>
rect 491 401 492 402 
<< m1 >>
rect 492 401 493 402 
<< m1 >>
rect 493 401 494 402 
<< m1 >>
rect 494 401 495 402 
<< m1 >>
rect 495 401 496 402 
<< m1 >>
rect 496 401 497 402 
<< m1 >>
rect 497 401 498 402 
<< m1 >>
rect 498 401 499 402 
<< m1 >>
rect 499 401 500 402 
<< m1 >>
rect 500 401 501 402 
<< m1 >>
rect 501 401 502 402 
<< m1 >>
rect 502 401 503 402 
<< m1 >>
rect 503 401 504 402 
<< m1 >>
rect 504 401 505 402 
<< m1 >>
rect 505 401 506 402 
<< m1 >>
rect 506 401 507 402 
<< m1 >>
rect 507 401 508 402 
<< m1 >>
rect 508 401 509 402 
<< m1 >>
rect 509 401 510 402 
<< m1 >>
rect 510 401 511 402 
<< m1 >>
rect 511 401 512 402 
<< m1 >>
rect 512 401 513 402 
<< m1 >>
rect 513 401 514 402 
<< m1 >>
rect 514 401 515 402 
<< m1 >>
rect 515 401 516 402 
<< m1 >>
rect 516 401 517 402 
<< m1 >>
rect 517 401 518 402 
<< m1 >>
rect 518 401 519 402 
<< m1 >>
rect 519 401 520 402 
<< m1 >>
rect 520 401 521 402 
<< m1 >>
rect 521 401 522 402 
<< m1 >>
rect 522 401 523 402 
<< m1 >>
rect 523 401 524 402 
<< m1 >>
rect 19 402 20 403 
<< m2 >>
rect 20 402 21 403 
<< m1 >>
rect 23 402 24 403 
<< m1 >>
rect 26 402 27 403 
<< m2 >>
rect 44 402 45 403 
<< m1 >>
rect 52 402 53 403 
<< m2 >>
rect 63 402 64 403 
<< m1 >>
rect 64 402 65 403 
<< m2 >>
rect 64 402 65 403 
<< m2 >>
rect 65 402 66 403 
<< m1 >>
rect 66 402 67 403 
<< m2 >>
rect 66 402 67 403 
<< m2c >>
rect 66 402 67 403 
<< m1 >>
rect 66 402 67 403 
<< m2 >>
rect 66 402 67 403 
<< m1 >>
rect 67 402 68 403 
<< m1 >>
rect 68 402 69 403 
<< m1 >>
rect 69 402 70 403 
<< m1 >>
rect 70 402 71 403 
<< m1 >>
rect 71 402 72 403 
<< m2 >>
rect 71 402 72 403 
<< m2c >>
rect 71 402 72 403 
<< m1 >>
rect 71 402 72 403 
<< m2 >>
rect 71 402 72 403 
<< m2 >>
rect 72 402 73 403 
<< m1 >>
rect 73 402 74 403 
<< m2 >>
rect 73 402 74 403 
<< m1 >>
rect 78 402 79 403 
<< m1 >>
rect 82 402 83 403 
<< m2 >>
rect 93 402 94 403 
<< m2 >>
rect 99 402 100 403 
<< m2 >>
rect 102 402 103 403 
<< m2 >>
rect 103 402 104 403 
<< m2 >>
rect 104 402 105 403 
<< m1 >>
rect 105 402 106 403 
<< m2 >>
rect 105 402 106 403 
<< m2c >>
rect 105 402 106 403 
<< m1 >>
rect 105 402 106 403 
<< m2 >>
rect 105 402 106 403 
<< m1 >>
rect 106 402 107 403 
<< m1 >>
rect 107 402 108 403 
<< m1 >>
rect 108 402 109 403 
<< m1 >>
rect 109 402 110 403 
<< m1 >>
rect 110 402 111 403 
<< m2 >>
rect 110 402 111 403 
<< m1 >>
rect 111 402 112 403 
<< m1 >>
rect 112 402 113 403 
<< m1 >>
rect 113 402 114 403 
<< m1 >>
rect 114 402 115 403 
<< m2 >>
rect 114 402 115 403 
<< m1 >>
rect 115 402 116 403 
<< m1 >>
rect 116 402 117 403 
<< m1 >>
rect 117 402 118 403 
<< m1 >>
rect 118 402 119 403 
<< m2 >>
rect 118 402 119 403 
<< m2c >>
rect 118 402 119 403 
<< m1 >>
rect 118 402 119 403 
<< m2 >>
rect 118 402 119 403 
<< m1 >>
rect 121 402 122 403 
<< m2 >>
rect 121 402 122 403 
<< m2c >>
rect 121 402 122 403 
<< m1 >>
rect 121 402 122 403 
<< m2 >>
rect 121 402 122 403 
<< m1 >>
rect 136 402 137 403 
<< m1 >>
rect 137 402 138 403 
<< m1 >>
rect 138 402 139 403 
<< m1 >>
rect 139 402 140 403 
<< m1 >>
rect 140 402 141 403 
<< m1 >>
rect 141 402 142 403 
<< m1 >>
rect 142 402 143 403 
<< m1 >>
rect 143 402 144 403 
<< m1 >>
rect 144 402 145 403 
<< m1 >>
rect 145 402 146 403 
<< m1 >>
rect 146 402 147 403 
<< m2 >>
rect 146 402 147 403 
<< m1 >>
rect 147 402 148 403 
<< m2 >>
rect 147 402 148 403 
<< m1 >>
rect 148 402 149 403 
<< m2 >>
rect 148 402 149 403 
<< m2 >>
rect 149 402 150 403 
<< m1 >>
rect 150 402 151 403 
<< m2 >>
rect 150 402 151 403 
<< m2 >>
rect 151 402 152 403 
<< m1 >>
rect 152 402 153 403 
<< m2 >>
rect 152 402 153 403 
<< m2c >>
rect 152 402 153 403 
<< m1 >>
rect 152 402 153 403 
<< m2 >>
rect 152 402 153 403 
<< m1 >>
rect 153 402 154 403 
<< m1 >>
rect 154 402 155 403 
<< m1 >>
rect 155 402 156 403 
<< m2 >>
rect 155 402 156 403 
<< m2c >>
rect 155 402 156 403 
<< m1 >>
rect 155 402 156 403 
<< m2 >>
rect 155 402 156 403 
<< m2 >>
rect 156 402 157 403 
<< m1 >>
rect 157 402 158 403 
<< m2 >>
rect 157 402 158 403 
<< m2 >>
rect 158 402 159 403 
<< m1 >>
rect 159 402 160 403 
<< m2 >>
rect 159 402 160 403 
<< m2c >>
rect 159 402 160 403 
<< m1 >>
rect 159 402 160 403 
<< m2 >>
rect 159 402 160 403 
<< m1 >>
rect 160 402 161 403 
<< m1 >>
rect 161 402 162 403 
<< m1 >>
rect 162 402 163 403 
<< m1 >>
rect 163 402 164 403 
<< m1 >>
rect 164 402 165 403 
<< m1 >>
rect 165 402 166 403 
<< m1 >>
rect 166 402 167 403 
<< m1 >>
rect 167 402 168 403 
<< m2 >>
rect 177 402 178 403 
<< m1 >>
rect 178 402 179 403 
<< m1 >>
rect 196 402 197 403 
<< m2 >>
rect 196 402 197 403 
<< m2c >>
rect 196 402 197 403 
<< m1 >>
rect 196 402 197 403 
<< m2 >>
rect 196 402 197 403 
<< m2 >>
rect 207 402 208 403 
<< m1 >>
rect 208 402 209 403 
<< m2 >>
rect 218 402 219 403 
<< m2 >>
rect 234 402 235 403 
<< m1 >>
rect 235 402 236 403 
<< m1 >>
rect 253 402 254 403 
<< m1 >>
rect 255 402 256 403 
<< m1 >>
rect 278 402 279 403 
<< m1 >>
rect 280 402 281 403 
<< m2 >>
rect 284 402 285 403 
<< m2 >>
rect 285 402 286 403 
<< m2 >>
rect 286 402 287 403 
<< m2 >>
rect 287 402 288 403 
<< m2 >>
rect 288 402 289 403 
<< m2 >>
rect 289 402 290 403 
<< m2 >>
rect 290 402 291 403 
<< m2 >>
rect 291 402 292 403 
<< m2 >>
rect 292 402 293 403 
<< m2 >>
rect 293 402 294 403 
<< m2 >>
rect 294 402 295 403 
<< m2 >>
rect 295 402 296 403 
<< m2 >>
rect 296 402 297 403 
<< m2 >>
rect 297 402 298 403 
<< m2 >>
rect 298 402 299 403 
<< m2 >>
rect 299 402 300 403 
<< m2 >>
rect 300 402 301 403 
<< m2 >>
rect 301 402 302 403 
<< m2 >>
rect 302 402 303 403 
<< m2 >>
rect 304 402 305 403 
<< m2 >>
rect 305 402 306 403 
<< m2 >>
rect 306 402 307 403 
<< m2 >>
rect 307 402 308 403 
<< m2 >>
rect 308 402 309 403 
<< m2 >>
rect 309 402 310 403 
<< m2 >>
rect 310 402 311 403 
<< m1 >>
rect 314 402 315 403 
<< m1 >>
rect 316 402 317 403 
<< m1 >>
rect 325 402 326 403 
<< m2 >>
rect 357 402 358 403 
<< m1 >>
rect 361 402 362 403 
<< m1 >>
rect 363 402 364 403 
<< m1 >>
rect 379 402 380 403 
<< m2 >>
rect 383 402 384 403 
<< m2 >>
rect 385 402 386 403 
<< m2 >>
rect 402 402 403 403 
<< m1 >>
rect 406 402 407 403 
<< m1 >>
rect 416 402 417 403 
<< m1 >>
rect 427 402 428 403 
<< m1 >>
rect 433 402 434 403 
<< m1 >>
rect 435 402 436 403 
<< m2 >>
rect 439 402 440 403 
<< m2 >>
rect 440 402 441 403 
<< m2 >>
rect 441 402 442 403 
<< m2 >>
rect 442 402 443 403 
<< m2 >>
rect 443 402 444 403 
<< m2 >>
rect 444 402 445 403 
<< m2 >>
rect 445 402 446 403 
<< m2 >>
rect 446 402 447 403 
<< m2 >>
rect 447 402 448 403 
<< m2 >>
rect 448 402 449 403 
<< m2 >>
rect 449 402 450 403 
<< m1 >>
rect 450 402 451 403 
<< m2 >>
rect 450 402 451 403 
<< m2c >>
rect 450 402 451 403 
<< m1 >>
rect 450 402 451 403 
<< m2 >>
rect 450 402 451 403 
<< m1 >>
rect 451 402 452 403 
<< m1 >>
rect 452 402 453 403 
<< m1 >>
rect 453 402 454 403 
<< m1 >>
rect 454 402 455 403 
<< m1 >>
rect 455 402 456 403 
<< m2 >>
rect 455 402 456 403 
<< m1 >>
rect 456 402 457 403 
<< m1 >>
rect 457 402 458 403 
<< m1 >>
rect 458 402 459 403 
<< m1 >>
rect 459 402 460 403 
<< m1 >>
rect 460 402 461 403 
<< m1 >>
rect 461 402 462 403 
<< m1 >>
rect 462 402 463 403 
<< m1 >>
rect 463 402 464 403 
<< m1 >>
rect 464 402 465 403 
<< m2 >>
rect 464 402 465 403 
<< m1 >>
rect 465 402 466 403 
<< m1 >>
rect 466 402 467 403 
<< m1 >>
rect 467 402 468 403 
<< m1 >>
rect 468 402 469 403 
<< m2 >>
rect 468 402 469 403 
<< m2c >>
rect 468 402 469 403 
<< m1 >>
rect 468 402 469 403 
<< m2 >>
rect 468 402 469 403 
<< m2 >>
rect 469 402 470 403 
<< m1 >>
rect 470 402 471 403 
<< m2 >>
rect 470 402 471 403 
<< m2 >>
rect 471 402 472 403 
<< m1 >>
rect 472 402 473 403 
<< m2 >>
rect 472 402 473 403 
<< m2 >>
rect 473 402 474 403 
<< m1 >>
rect 474 402 475 403 
<< m2 >>
rect 474 402 475 403 
<< m2c >>
rect 474 402 475 403 
<< m1 >>
rect 474 402 475 403 
<< m2 >>
rect 474 402 475 403 
<< m1 >>
rect 475 402 476 403 
<< m1 >>
rect 476 402 477 403 
<< m2 >>
rect 476 402 477 403 
<< m1 >>
rect 477 402 478 403 
<< m1 >>
rect 478 402 479 403 
<< m1 >>
rect 479 402 480 403 
<< m1 >>
rect 480 402 481 403 
<< m1 >>
rect 481 402 482 403 
<< m2 >>
rect 481 402 482 403 
<< m1 >>
rect 482 402 483 403 
<< m1 >>
rect 483 402 484 403 
<< m1 >>
rect 484 402 485 403 
<< m1 >>
rect 485 402 486 403 
<< m1 >>
rect 486 402 487 403 
<< m1 >>
rect 487 402 488 403 
<< m1 >>
rect 488 402 489 403 
<< m1 >>
rect 489 402 490 403 
<< m2 >>
rect 490 402 491 403 
<< m1 >>
rect 19 403 20 404 
<< m2 >>
rect 20 403 21 404 
<< m1 >>
rect 23 403 24 404 
<< m1 >>
rect 26 403 27 404 
<< m1 >>
rect 37 403 38 404 
<< m1 >>
rect 38 403 39 404 
<< m1 >>
rect 39 403 40 404 
<< m1 >>
rect 40 403 41 404 
<< m1 >>
rect 41 403 42 404 
<< m1 >>
rect 42 403 43 404 
<< m1 >>
rect 43 403 44 404 
<< m1 >>
rect 44 403 45 404 
<< m2 >>
rect 44 403 45 404 
<< m1 >>
rect 45 403 46 404 
<< m1 >>
rect 46 403 47 404 
<< m1 >>
rect 47 403 48 404 
<< m1 >>
rect 48 403 49 404 
<< m1 >>
rect 49 403 50 404 
<< m1 >>
rect 50 403 51 404 
<< m1 >>
rect 51 403 52 404 
<< m1 >>
rect 52 403 53 404 
<< m1 >>
rect 64 403 65 404 
<< m1 >>
rect 73 403 74 404 
<< m2 >>
rect 73 403 74 404 
<< m1 >>
rect 78 403 79 404 
<< m1 >>
rect 79 403 80 404 
<< m1 >>
rect 80 403 81 404 
<< m2 >>
rect 80 403 81 404 
<< m2c >>
rect 80 403 81 404 
<< m1 >>
rect 80 403 81 404 
<< m2 >>
rect 80 403 81 404 
<< m2 >>
rect 81 403 82 404 
<< m1 >>
rect 82 403 83 404 
<< m2 >>
rect 82 403 83 404 
<< m2 >>
rect 83 403 84 404 
<< m1 >>
rect 84 403 85 404 
<< m2 >>
rect 84 403 85 404 
<< m2c >>
rect 84 403 85 404 
<< m1 >>
rect 84 403 85 404 
<< m2 >>
rect 84 403 85 404 
<< m1 >>
rect 85 403 86 404 
<< m1 >>
rect 86 403 87 404 
<< m1 >>
rect 87 403 88 404 
<< m1 >>
rect 88 403 89 404 
<< m1 >>
rect 89 403 90 404 
<< m1 >>
rect 90 403 91 404 
<< m1 >>
rect 91 403 92 404 
<< m1 >>
rect 92 403 93 404 
<< m1 >>
rect 93 403 94 404 
<< m2 >>
rect 93 403 94 404 
<< m1 >>
rect 94 403 95 404 
<< m1 >>
rect 95 403 96 404 
<< m1 >>
rect 96 403 97 404 
<< m1 >>
rect 97 403 98 404 
<< m1 >>
rect 98 403 99 404 
<< m1 >>
rect 99 403 100 404 
<< m2 >>
rect 99 403 100 404 
<< m1 >>
rect 100 403 101 404 
<< m1 >>
rect 101 403 102 404 
<< m1 >>
rect 102 403 103 404 
<< m2 >>
rect 102 403 103 404 
<< m1 >>
rect 103 403 104 404 
<< m2 >>
rect 110 403 111 404 
<< m2 >>
rect 114 403 115 404 
<< m1 >>
rect 121 403 122 404 
<< m1 >>
rect 136 403 137 404 
<< m1 >>
rect 150 403 151 404 
<< m1 >>
rect 157 403 158 404 
<< m1 >>
rect 169 403 170 404 
<< m1 >>
rect 170 403 171 404 
<< m1 >>
rect 171 403 172 404 
<< m1 >>
rect 172 403 173 404 
<< m1 >>
rect 173 403 174 404 
<< m1 >>
rect 174 403 175 404 
<< m1 >>
rect 175 403 176 404 
<< m1 >>
rect 176 403 177 404 
<< m2 >>
rect 176 403 177 404 
<< m2c >>
rect 176 403 177 404 
<< m1 >>
rect 176 403 177 404 
<< m2 >>
rect 176 403 177 404 
<< m2 >>
rect 177 403 178 404 
<< m1 >>
rect 178 403 179 404 
<< m1 >>
rect 181 403 182 404 
<< m1 >>
rect 182 403 183 404 
<< m1 >>
rect 183 403 184 404 
<< m1 >>
rect 184 403 185 404 
<< m1 >>
rect 185 403 186 404 
<< m1 >>
rect 186 403 187 404 
<< m1 >>
rect 187 403 188 404 
<< m1 >>
rect 188 403 189 404 
<< m1 >>
rect 189 403 190 404 
<< m1 >>
rect 190 403 191 404 
<< m1 >>
rect 191 403 192 404 
<< m1 >>
rect 192 403 193 404 
<< m1 >>
rect 193 403 194 404 
<< m1 >>
rect 194 403 195 404 
<< m1 >>
rect 195 403 196 404 
<< m1 >>
rect 196 403 197 404 
<< m2 >>
rect 207 403 208 404 
<< m1 >>
rect 208 403 209 404 
<< m1 >>
rect 210 403 211 404 
<< m1 >>
rect 211 403 212 404 
<< m1 >>
rect 212 403 213 404 
<< m1 >>
rect 213 403 214 404 
<< m1 >>
rect 214 403 215 404 
<< m1 >>
rect 215 403 216 404 
<< m1 >>
rect 216 403 217 404 
<< m1 >>
rect 217 403 218 404 
<< m1 >>
rect 218 403 219 404 
<< m2 >>
rect 218 403 219 404 
<< m1 >>
rect 219 403 220 404 
<< m1 >>
rect 220 403 221 404 
<< m1 >>
rect 221 403 222 404 
<< m1 >>
rect 222 403 223 404 
<< m1 >>
rect 223 403 224 404 
<< m1 >>
rect 224 403 225 404 
<< m1 >>
rect 225 403 226 404 
<< m1 >>
rect 226 403 227 404 
<< m1 >>
rect 227 403 228 404 
<< m1 >>
rect 228 403 229 404 
<< m1 >>
rect 229 403 230 404 
<< m1 >>
rect 230 403 231 404 
<< m1 >>
rect 231 403 232 404 
<< m1 >>
rect 232 403 233 404 
<< m1 >>
rect 233 403 234 404 
<< m2 >>
rect 233 403 234 404 
<< m2c >>
rect 233 403 234 404 
<< m1 >>
rect 233 403 234 404 
<< m2 >>
rect 233 403 234 404 
<< m2 >>
rect 234 403 235 404 
<< m1 >>
rect 235 403 236 404 
<< m1 >>
rect 237 403 238 404 
<< m1 >>
rect 238 403 239 404 
<< m1 >>
rect 239 403 240 404 
<< m1 >>
rect 240 403 241 404 
<< m1 >>
rect 241 403 242 404 
<< m1 >>
rect 242 403 243 404 
<< m1 >>
rect 243 403 244 404 
<< m1 >>
rect 244 403 245 404 
<< m1 >>
rect 245 403 246 404 
<< m1 >>
rect 246 403 247 404 
<< m1 >>
rect 247 403 248 404 
<< m1 >>
rect 248 403 249 404 
<< m1 >>
rect 249 403 250 404 
<< m1 >>
rect 250 403 251 404 
<< m1 >>
rect 251 403 252 404 
<< m2 >>
rect 251 403 252 404 
<< m2c >>
rect 251 403 252 404 
<< m1 >>
rect 251 403 252 404 
<< m2 >>
rect 251 403 252 404 
<< m2 >>
rect 252 403 253 404 
<< m1 >>
rect 253 403 254 404 
<< m2 >>
rect 253 403 254 404 
<< m2 >>
rect 254 403 255 404 
<< m1 >>
rect 255 403 256 404 
<< m2 >>
rect 255 403 256 404 
<< m2c >>
rect 255 403 256 404 
<< m1 >>
rect 255 403 256 404 
<< m2 >>
rect 255 403 256 404 
<< m1 >>
rect 278 403 279 404 
<< m2 >>
rect 278 403 279 404 
<< m2c >>
rect 278 403 279 404 
<< m1 >>
rect 278 403 279 404 
<< m2 >>
rect 278 403 279 404 
<< m2 >>
rect 279 403 280 404 
<< m1 >>
rect 280 403 281 404 
<< m2 >>
rect 280 403 281 404 
<< m2 >>
rect 281 403 282 404 
<< m1 >>
rect 282 403 283 404 
<< m2 >>
rect 282 403 283 404 
<< m2c >>
rect 282 403 283 404 
<< m1 >>
rect 282 403 283 404 
<< m2 >>
rect 282 403 283 404 
<< m1 >>
rect 283 403 284 404 
<< m1 >>
rect 284 403 285 404 
<< m1 >>
rect 285 403 286 404 
<< m1 >>
rect 286 403 287 404 
<< m1 >>
rect 287 403 288 404 
<< m1 >>
rect 288 403 289 404 
<< m1 >>
rect 289 403 290 404 
<< m1 >>
rect 290 403 291 404 
<< m1 >>
rect 291 403 292 404 
<< m1 >>
rect 292 403 293 404 
<< m1 >>
rect 293 403 294 404 
<< m1 >>
rect 294 403 295 404 
<< m1 >>
rect 295 403 296 404 
<< m1 >>
rect 296 403 297 404 
<< m1 >>
rect 297 403 298 404 
<< m1 >>
rect 298 403 299 404 
<< m1 >>
rect 299 403 300 404 
<< m1 >>
rect 300 403 301 404 
<< m1 >>
rect 301 403 302 404 
<< m1 >>
rect 302 403 303 404 
<< m2 >>
rect 302 403 303 404 
<< m1 >>
rect 303 403 304 404 
<< m1 >>
rect 304 403 305 404 
<< m2 >>
rect 304 403 305 404 
<< m1 >>
rect 305 403 306 404 
<< m1 >>
rect 306 403 307 404 
<< m1 >>
rect 307 403 308 404 
<< m1 >>
rect 308 403 309 404 
<< m1 >>
rect 309 403 310 404 
<< m1 >>
rect 310 403 311 404 
<< m1 >>
rect 311 403 312 404 
<< m1 >>
rect 312 403 313 404 
<< m2 >>
rect 312 403 313 404 
<< m2c >>
rect 312 403 313 404 
<< m1 >>
rect 312 403 313 404 
<< m2 >>
rect 312 403 313 404 
<< m2 >>
rect 313 403 314 404 
<< m1 >>
rect 314 403 315 404 
<< m2 >>
rect 314 403 315 404 
<< m2 >>
rect 315 403 316 404 
<< m1 >>
rect 316 403 317 404 
<< m2 >>
rect 316 403 317 404 
<< m2 >>
rect 317 403 318 404 
<< m1 >>
rect 318 403 319 404 
<< m2 >>
rect 318 403 319 404 
<< m2c >>
rect 318 403 319 404 
<< m1 >>
rect 318 403 319 404 
<< m2 >>
rect 318 403 319 404 
<< m1 >>
rect 319 403 320 404 
<< m1 >>
rect 320 403 321 404 
<< m1 >>
rect 321 403 322 404 
<< m1 >>
rect 322 403 323 404 
<< m1 >>
rect 323 403 324 404 
<< m2 >>
rect 323 403 324 404 
<< m2c >>
rect 323 403 324 404 
<< m1 >>
rect 323 403 324 404 
<< m2 >>
rect 323 403 324 404 
<< m2 >>
rect 324 403 325 404 
<< m1 >>
rect 325 403 326 404 
<< m2 >>
rect 325 403 326 404 
<< m2 >>
rect 326 403 327 404 
<< m1 >>
rect 327 403 328 404 
<< m2 >>
rect 327 403 328 404 
<< m2c >>
rect 327 403 328 404 
<< m1 >>
rect 327 403 328 404 
<< m2 >>
rect 327 403 328 404 
<< m1 >>
rect 328 403 329 404 
<< m1 >>
rect 329 403 330 404 
<< m2 >>
rect 329 403 330 404 
<< m1 >>
rect 330 403 331 404 
<< m2 >>
rect 330 403 331 404 
<< m1 >>
rect 331 403 332 404 
<< m2 >>
rect 331 403 332 404 
<< m1 >>
rect 332 403 333 404 
<< m2 >>
rect 332 403 333 404 
<< m1 >>
rect 333 403 334 404 
<< m2 >>
rect 333 403 334 404 
<< m1 >>
rect 334 403 335 404 
<< m2 >>
rect 334 403 335 404 
<< m1 >>
rect 335 403 336 404 
<< m2 >>
rect 335 403 336 404 
<< m1 >>
rect 336 403 337 404 
<< m2 >>
rect 336 403 337 404 
<< m1 >>
rect 337 403 338 404 
<< m2 >>
rect 337 403 338 404 
<< m1 >>
rect 338 403 339 404 
<< m2 >>
rect 338 403 339 404 
<< m1 >>
rect 339 403 340 404 
<< m1 >>
rect 340 403 341 404 
<< m1 >>
rect 341 403 342 404 
<< m1 >>
rect 342 403 343 404 
<< m1 >>
rect 343 403 344 404 
<< m1 >>
rect 344 403 345 404 
<< m1 >>
rect 345 403 346 404 
<< m1 >>
rect 346 403 347 404 
<< m1 >>
rect 347 403 348 404 
<< m1 >>
rect 348 403 349 404 
<< m1 >>
rect 349 403 350 404 
<< m1 >>
rect 350 403 351 404 
<< m1 >>
rect 351 403 352 404 
<< m1 >>
rect 352 403 353 404 
<< m1 >>
rect 353 403 354 404 
<< m1 >>
rect 354 403 355 404 
<< m1 >>
rect 355 403 356 404 
<< m1 >>
rect 356 403 357 404 
<< m1 >>
rect 357 403 358 404 
<< m2 >>
rect 357 403 358 404 
<< m1 >>
rect 358 403 359 404 
<< m1 >>
rect 359 403 360 404 
<< m2 >>
rect 359 403 360 404 
<< m2c >>
rect 359 403 360 404 
<< m1 >>
rect 359 403 360 404 
<< m2 >>
rect 359 403 360 404 
<< m2 >>
rect 360 403 361 404 
<< m1 >>
rect 361 403 362 404 
<< m2 >>
rect 361 403 362 404 
<< m2 >>
rect 362 403 363 404 
<< m1 >>
rect 363 403 364 404 
<< m2 >>
rect 363 403 364 404 
<< m2 >>
rect 364 403 365 404 
<< m1 >>
rect 365 403 366 404 
<< m2 >>
rect 365 403 366 404 
<< m2c >>
rect 365 403 366 404 
<< m1 >>
rect 365 403 366 404 
<< m2 >>
rect 365 403 366 404 
<< m1 >>
rect 366 403 367 404 
<< m1 >>
rect 367 403 368 404 
<< m2 >>
rect 367 403 368 404 
<< m1 >>
rect 368 403 369 404 
<< m2 >>
rect 368 403 369 404 
<< m1 >>
rect 369 403 370 404 
<< m2 >>
rect 369 403 370 404 
<< m1 >>
rect 370 403 371 404 
<< m2 >>
rect 370 403 371 404 
<< m1 >>
rect 371 403 372 404 
<< m2 >>
rect 371 403 372 404 
<< m1 >>
rect 372 403 373 404 
<< m2 >>
rect 372 403 373 404 
<< m1 >>
rect 373 403 374 404 
<< m2 >>
rect 373 403 374 404 
<< m1 >>
rect 374 403 375 404 
<< m2 >>
rect 374 403 375 404 
<< m1 >>
rect 375 403 376 404 
<< m1 >>
rect 376 403 377 404 
<< m1 >>
rect 377 403 378 404 
<< m2 >>
rect 377 403 378 404 
<< m2c >>
rect 377 403 378 404 
<< m1 >>
rect 377 403 378 404 
<< m2 >>
rect 377 403 378 404 
<< m2 >>
rect 378 403 379 404 
<< m1 >>
rect 379 403 380 404 
<< m2 >>
rect 379 403 380 404 
<< m2 >>
rect 380 403 381 404 
<< m1 >>
rect 381 403 382 404 
<< m2 >>
rect 381 403 382 404 
<< m2c >>
rect 381 403 382 404 
<< m1 >>
rect 381 403 382 404 
<< m2 >>
rect 381 403 382 404 
<< m1 >>
rect 382 403 383 404 
<< m1 >>
rect 383 403 384 404 
<< m2 >>
rect 383 403 384 404 
<< m1 >>
rect 384 403 385 404 
<< m1 >>
rect 385 403 386 404 
<< m2 >>
rect 385 403 386 404 
<< m1 >>
rect 386 403 387 404 
<< m1 >>
rect 387 403 388 404 
<< m1 >>
rect 388 403 389 404 
<< m1 >>
rect 389 403 390 404 
<< m1 >>
rect 390 403 391 404 
<< m1 >>
rect 391 403 392 404 
<< m1 >>
rect 392 403 393 404 
<< m1 >>
rect 393 403 394 404 
<< m1 >>
rect 394 403 395 404 
<< m1 >>
rect 395 403 396 404 
<< m1 >>
rect 396 403 397 404 
<< m1 >>
rect 397 403 398 404 
<< m1 >>
rect 398 403 399 404 
<< m1 >>
rect 399 403 400 404 
<< m1 >>
rect 400 403 401 404 
<< m1 >>
rect 401 403 402 404 
<< m1 >>
rect 402 403 403 404 
<< m2 >>
rect 402 403 403 404 
<< m1 >>
rect 403 403 404 404 
<< m1 >>
rect 404 403 405 404 
<< m2 >>
rect 404 403 405 404 
<< m2c >>
rect 404 403 405 404 
<< m1 >>
rect 404 403 405 404 
<< m2 >>
rect 404 403 405 404 
<< m2 >>
rect 405 403 406 404 
<< m1 >>
rect 406 403 407 404 
<< m2 >>
rect 406 403 407 404 
<< m2 >>
rect 407 403 408 404 
<< m1 >>
rect 408 403 409 404 
<< m2 >>
rect 408 403 409 404 
<< m2c >>
rect 408 403 409 404 
<< m1 >>
rect 408 403 409 404 
<< m2 >>
rect 408 403 409 404 
<< m1 >>
rect 409 403 410 404 
<< m1 >>
rect 410 403 411 404 
<< m1 >>
rect 411 403 412 404 
<< m1 >>
rect 412 403 413 404 
<< m1 >>
rect 413 403 414 404 
<< m1 >>
rect 414 403 415 404 
<< m2 >>
rect 414 403 415 404 
<< m2c >>
rect 414 403 415 404 
<< m1 >>
rect 414 403 415 404 
<< m2 >>
rect 414 403 415 404 
<< m2 >>
rect 415 403 416 404 
<< m1 >>
rect 416 403 417 404 
<< m2 >>
rect 416 403 417 404 
<< m2 >>
rect 417 403 418 404 
<< m1 >>
rect 418 403 419 404 
<< m2 >>
rect 418 403 419 404 
<< m2c >>
rect 418 403 419 404 
<< m1 >>
rect 418 403 419 404 
<< m2 >>
rect 418 403 419 404 
<< m1 >>
rect 419 403 420 404 
<< m1 >>
rect 420 403 421 404 
<< m1 >>
rect 421 403 422 404 
<< m1 >>
rect 422 403 423 404 
<< m2 >>
rect 422 403 423 404 
<< m2c >>
rect 422 403 423 404 
<< m1 >>
rect 422 403 423 404 
<< m2 >>
rect 422 403 423 404 
<< m2 >>
rect 423 403 424 404 
<< m1 >>
rect 424 403 425 404 
<< m2 >>
rect 424 403 425 404 
<< m1 >>
rect 425 403 426 404 
<< m2 >>
rect 425 403 426 404 
<< m1 >>
rect 426 403 427 404 
<< m2 >>
rect 426 403 427 404 
<< m1 >>
rect 427 403 428 404 
<< m2 >>
rect 427 403 428 404 
<< m2 >>
rect 428 403 429 404 
<< m1 >>
rect 429 403 430 404 
<< m2 >>
rect 429 403 430 404 
<< m2c >>
rect 429 403 430 404 
<< m1 >>
rect 429 403 430 404 
<< m2 >>
rect 429 403 430 404 
<< m1 >>
rect 430 403 431 404 
<< m1 >>
rect 431 403 432 404 
<< m2 >>
rect 431 403 432 404 
<< m2c >>
rect 431 403 432 404 
<< m1 >>
rect 431 403 432 404 
<< m2 >>
rect 431 403 432 404 
<< m2 >>
rect 432 403 433 404 
<< m1 >>
rect 433 403 434 404 
<< m2 >>
rect 433 403 434 404 
<< m2 >>
rect 434 403 435 404 
<< m1 >>
rect 435 403 436 404 
<< m2 >>
rect 435 403 436 404 
<< m2 >>
rect 436 403 437 404 
<< m1 >>
rect 437 403 438 404 
<< m2 >>
rect 437 403 438 404 
<< m2c >>
rect 437 403 438 404 
<< m1 >>
rect 437 403 438 404 
<< m2 >>
rect 437 403 438 404 
<< m1 >>
rect 438 403 439 404 
<< m1 >>
rect 439 403 440 404 
<< m1 >>
rect 440 403 441 404 
<< m1 >>
rect 441 403 442 404 
<< m1 >>
rect 442 403 443 404 
<< m1 >>
rect 443 403 444 404 
<< m1 >>
rect 444 403 445 404 
<< m1 >>
rect 445 403 446 404 
<< m1 >>
rect 446 403 447 404 
<< m1 >>
rect 447 403 448 404 
<< m1 >>
rect 448 403 449 404 
<< m2 >>
rect 455 403 456 404 
<< m2 >>
rect 456 403 457 404 
<< m2 >>
rect 457 403 458 404 
<< m2 >>
rect 458 403 459 404 
<< m2 >>
rect 459 403 460 404 
<< m2 >>
rect 460 403 461 404 
<< m2 >>
rect 461 403 462 404 
<< m2 >>
rect 462 403 463 404 
<< m2 >>
rect 464 403 465 404 
<< m1 >>
rect 470 403 471 404 
<< m1 >>
rect 472 403 473 404 
<< m2 >>
rect 476 403 477 404 
<< m2 >>
rect 481 403 482 404 
<< m1 >>
rect 489 403 490 404 
<< m2 >>
rect 490 403 491 404 
<< m1 >>
rect 19 404 20 405 
<< m2 >>
rect 20 404 21 405 
<< m1 >>
rect 23 404 24 405 
<< m1 >>
rect 26 404 27 405 
<< m1 >>
rect 37 404 38 405 
<< m2 >>
rect 44 404 45 405 
<< m1 >>
rect 64 404 65 405 
<< m1 >>
rect 73 404 74 405 
<< m2 >>
rect 73 404 74 405 
<< m1 >>
rect 82 404 83 405 
<< m2 >>
rect 93 404 94 405 
<< m2 >>
rect 99 404 100 405 
<< m2 >>
rect 102 404 103 405 
<< m1 >>
rect 103 404 104 405 
<< m1 >>
rect 110 404 111 405 
<< m2 >>
rect 110 404 111 405 
<< m2c >>
rect 110 404 111 405 
<< m1 >>
rect 110 404 111 405 
<< m2 >>
rect 110 404 111 405 
<< m1 >>
rect 114 404 115 405 
<< m2 >>
rect 114 404 115 405 
<< m2c >>
rect 114 404 115 405 
<< m1 >>
rect 114 404 115 405 
<< m2 >>
rect 114 404 115 405 
<< m1 >>
rect 121 404 122 405 
<< m1 >>
rect 136 404 137 405 
<< m1 >>
rect 150 404 151 405 
<< m1 >>
rect 157 404 158 405 
<< m1 >>
rect 169 404 170 405 
<< m1 >>
rect 178 404 179 405 
<< m1 >>
rect 181 404 182 405 
<< m1 >>
rect 199 404 200 405 
<< m2 >>
rect 199 404 200 405 
<< m2c >>
rect 199 404 200 405 
<< m1 >>
rect 199 404 200 405 
<< m2 >>
rect 199 404 200 405 
<< m1 >>
rect 200 404 201 405 
<< m1 >>
rect 201 404 202 405 
<< m1 >>
rect 202 404 203 405 
<< m1 >>
rect 203 404 204 405 
<< m1 >>
rect 204 404 205 405 
<< m1 >>
rect 205 404 206 405 
<< m1 >>
rect 206 404 207 405 
<< m2 >>
rect 206 404 207 405 
<< m2c >>
rect 206 404 207 405 
<< m1 >>
rect 206 404 207 405 
<< m2 >>
rect 206 404 207 405 
<< m2 >>
rect 207 404 208 405 
<< m1 >>
rect 208 404 209 405 
<< m1 >>
rect 210 404 211 405 
<< m2 >>
rect 217 404 218 405 
<< m2 >>
rect 218 404 219 405 
<< m1 >>
rect 235 404 236 405 
<< m1 >>
rect 237 404 238 405 
<< m1 >>
rect 253 404 254 405 
<< m1 >>
rect 280 404 281 405 
<< m2 >>
rect 302 404 303 405 
<< m2 >>
rect 304 404 305 405 
<< m1 >>
rect 314 404 315 405 
<< m1 >>
rect 316 404 317 405 
<< m1 >>
rect 325 404 326 405 
<< m2 >>
rect 329 404 330 405 
<< m2 >>
rect 338 404 339 405 
<< m2 >>
rect 357 404 358 405 
<< m1 >>
rect 361 404 362 405 
<< m1 >>
rect 363 404 364 405 
<< m2 >>
rect 367 404 368 405 
<< m2 >>
rect 374 404 375 405 
<< m1 >>
rect 379 404 380 405 
<< m2 >>
rect 383 404 384 405 
<< m2 >>
rect 385 404 386 405 
<< m2 >>
rect 402 404 403 405 
<< m1 >>
rect 406 404 407 405 
<< m1 >>
rect 416 404 417 405 
<< m1 >>
rect 424 404 425 405 
<< m1 >>
rect 433 404 434 405 
<< m1 >>
rect 435 404 436 405 
<< m1 >>
rect 448 404 449 405 
<< m1 >>
rect 462 404 463 405 
<< m2 >>
rect 462 404 463 405 
<< m2c >>
rect 462 404 463 405 
<< m1 >>
rect 462 404 463 405 
<< m2 >>
rect 462 404 463 405 
<< m1 >>
rect 464 404 465 405 
<< m2 >>
rect 464 404 465 405 
<< m2c >>
rect 464 404 465 405 
<< m1 >>
rect 464 404 465 405 
<< m2 >>
rect 464 404 465 405 
<< m1 >>
rect 465 404 466 405 
<< m1 >>
rect 466 404 467 405 
<< m1 >>
rect 467 404 468 405 
<< m1 >>
rect 468 404 469 405 
<< m2 >>
rect 468 404 469 405 
<< m2c >>
rect 468 404 469 405 
<< m1 >>
rect 468 404 469 405 
<< m2 >>
rect 468 404 469 405 
<< m2 >>
rect 469 404 470 405 
<< m1 >>
rect 470 404 471 405 
<< m2 >>
rect 470 404 471 405 
<< m2 >>
rect 471 404 472 405 
<< m1 >>
rect 472 404 473 405 
<< m2 >>
rect 472 404 473 405 
<< m2 >>
rect 473 404 474 405 
<< m1 >>
rect 474 404 475 405 
<< m2 >>
rect 474 404 475 405 
<< m2c >>
rect 474 404 475 405 
<< m1 >>
rect 474 404 475 405 
<< m2 >>
rect 474 404 475 405 
<< m1 >>
rect 476 404 477 405 
<< m2 >>
rect 476 404 477 405 
<< m2c >>
rect 476 404 477 405 
<< m1 >>
rect 476 404 477 405 
<< m2 >>
rect 476 404 477 405 
<< m1 >>
rect 481 404 482 405 
<< m2 >>
rect 481 404 482 405 
<< m2c >>
rect 481 404 482 405 
<< m1 >>
rect 481 404 482 405 
<< m2 >>
rect 481 404 482 405 
<< m1 >>
rect 489 404 490 405 
<< m2 >>
rect 490 404 491 405 
<< m1 >>
rect 19 405 20 406 
<< m2 >>
rect 20 405 21 406 
<< m1 >>
rect 23 405 24 406 
<< m1 >>
rect 26 405 27 406 
<< m1 >>
rect 37 405 38 406 
<< m1 >>
rect 44 405 45 406 
<< m2 >>
rect 44 405 45 406 
<< m2c >>
rect 44 405 45 406 
<< m1 >>
rect 44 405 45 406 
<< m2 >>
rect 44 405 45 406 
<< m1 >>
rect 64 405 65 406 
<< m1 >>
rect 73 405 74 406 
<< m2 >>
rect 73 405 74 406 
<< m1 >>
rect 82 405 83 406 
<< m1 >>
rect 88 405 89 406 
<< m1 >>
rect 89 405 90 406 
<< m1 >>
rect 90 405 91 406 
<< m1 >>
rect 91 405 92 406 
<< m1 >>
rect 92 405 93 406 
<< m1 >>
rect 93 405 94 406 
<< m2 >>
rect 93 405 94 406 
<< m1 >>
rect 94 405 95 406 
<< m1 >>
rect 95 405 96 406 
<< m1 >>
rect 96 405 97 406 
<< m1 >>
rect 97 405 98 406 
<< m1 >>
rect 98 405 99 406 
<< m1 >>
rect 99 405 100 406 
<< m2 >>
rect 99 405 100 406 
<< m1 >>
rect 100 405 101 406 
<< m1 >>
rect 101 405 102 406 
<< m2 >>
rect 101 405 102 406 
<< m2c >>
rect 101 405 102 406 
<< m1 >>
rect 101 405 102 406 
<< m2 >>
rect 101 405 102 406 
<< m2 >>
rect 102 405 103 406 
<< m1 >>
rect 103 405 104 406 
<< m1 >>
rect 110 405 111 406 
<< m1 >>
rect 114 405 115 406 
<< m1 >>
rect 121 405 122 406 
<< m1 >>
rect 136 405 137 406 
<< m1 >>
rect 150 405 151 406 
<< m1 >>
rect 157 405 158 406 
<< m1 >>
rect 169 405 170 406 
<< m1 >>
rect 178 405 179 406 
<< m1 >>
rect 181 405 182 406 
<< m2 >>
rect 199 405 200 406 
<< m1 >>
rect 208 405 209 406 
<< m1 >>
rect 210 405 211 406 
<< m1 >>
rect 217 405 218 406 
<< m2 >>
rect 217 405 218 406 
<< m2c >>
rect 217 405 218 406 
<< m1 >>
rect 217 405 218 406 
<< m2 >>
rect 217 405 218 406 
<< m1 >>
rect 229 405 230 406 
<< m1 >>
rect 230 405 231 406 
<< m1 >>
rect 231 405 232 406 
<< m1 >>
rect 232 405 233 406 
<< m1 >>
rect 233 405 234 406 
<< m2 >>
rect 233 405 234 406 
<< m2c >>
rect 233 405 234 406 
<< m1 >>
rect 233 405 234 406 
<< m2 >>
rect 233 405 234 406 
<< m2 >>
rect 234 405 235 406 
<< m1 >>
rect 235 405 236 406 
<< m2 >>
rect 235 405 236 406 
<< m2 >>
rect 236 405 237 406 
<< m1 >>
rect 237 405 238 406 
<< m2 >>
rect 237 405 238 406 
<< m2c >>
rect 237 405 238 406 
<< m1 >>
rect 237 405 238 406 
<< m2 >>
rect 237 405 238 406 
<< m1 >>
rect 253 405 254 406 
<< m1 >>
rect 280 405 281 406 
<< m1 >>
rect 302 405 303 406 
<< m2 >>
rect 302 405 303 406 
<< m2c >>
rect 302 405 303 406 
<< m1 >>
rect 302 405 303 406 
<< m2 >>
rect 302 405 303 406 
<< m1 >>
rect 303 405 304 406 
<< m1 >>
rect 304 405 305 406 
<< m2 >>
rect 304 405 305 406 
<< m1 >>
rect 305 405 306 406 
<< m1 >>
rect 306 405 307 406 
<< m1 >>
rect 307 405 308 406 
<< m1 >>
rect 314 405 315 406 
<< m1 >>
rect 316 405 317 406 
<< m1 >>
rect 325 405 326 406 
<< m1 >>
rect 329 405 330 406 
<< m2 >>
rect 329 405 330 406 
<< m2c >>
rect 329 405 330 406 
<< m1 >>
rect 329 405 330 406 
<< m2 >>
rect 329 405 330 406 
<< m1 >>
rect 338 405 339 406 
<< m2 >>
rect 338 405 339 406 
<< m2c >>
rect 338 405 339 406 
<< m1 >>
rect 338 405 339 406 
<< m2 >>
rect 338 405 339 406 
<< m1 >>
rect 339 405 340 406 
<< m1 >>
rect 340 405 341 406 
<< m1 >>
rect 357 405 358 406 
<< m2 >>
rect 357 405 358 406 
<< m2c >>
rect 357 405 358 406 
<< m1 >>
rect 357 405 358 406 
<< m2 >>
rect 357 405 358 406 
<< m1 >>
rect 361 405 362 406 
<< m1 >>
rect 363 405 364 406 
<< m1 >>
rect 367 405 368 406 
<< m2 >>
rect 367 405 368 406 
<< m2c >>
rect 367 405 368 406 
<< m1 >>
rect 367 405 368 406 
<< m2 >>
rect 367 405 368 406 
<< m1 >>
rect 374 405 375 406 
<< m2 >>
rect 374 405 375 406 
<< m2c >>
rect 374 405 375 406 
<< m1 >>
rect 374 405 375 406 
<< m2 >>
rect 374 405 375 406 
<< m1 >>
rect 375 405 376 406 
<< m1 >>
rect 376 405 377 406 
<< m1 >>
rect 377 405 378 406 
<< m2 >>
rect 377 405 378 406 
<< m2c >>
rect 377 405 378 406 
<< m1 >>
rect 377 405 378 406 
<< m2 >>
rect 377 405 378 406 
<< m2 >>
rect 378 405 379 406 
<< m1 >>
rect 379 405 380 406 
<< m2 >>
rect 379 405 380 406 
<< m2 >>
rect 380 405 381 406 
<< m1 >>
rect 381 405 382 406 
<< m2 >>
rect 381 405 382 406 
<< m2c >>
rect 381 405 382 406 
<< m1 >>
rect 381 405 382 406 
<< m2 >>
rect 381 405 382 406 
<< m1 >>
rect 382 405 383 406 
<< m1 >>
rect 383 405 384 406 
<< m2 >>
rect 383 405 384 406 
<< m1 >>
rect 384 405 385 406 
<< m1 >>
rect 385 405 386 406 
<< m2 >>
rect 385 405 386 406 
<< m1 >>
rect 386 405 387 406 
<< m1 >>
rect 387 405 388 406 
<< m1 >>
rect 388 405 389 406 
<< m1 >>
rect 389 405 390 406 
<< m1 >>
rect 390 405 391 406 
<< m1 >>
rect 391 405 392 406 
<< m1 >>
rect 402 405 403 406 
<< m2 >>
rect 402 405 403 406 
<< m2c >>
rect 402 405 403 406 
<< m1 >>
rect 402 405 403 406 
<< m2 >>
rect 402 405 403 406 
<< m1 >>
rect 406 405 407 406 
<< m1 >>
rect 409 405 410 406 
<< m1 >>
rect 410 405 411 406 
<< m1 >>
rect 411 405 412 406 
<< m1 >>
rect 412 405 413 406 
<< m1 >>
rect 413 405 414 406 
<< m1 >>
rect 414 405 415 406 
<< m1 >>
rect 416 405 417 406 
<< m1 >>
rect 424 405 425 406 
<< m1 >>
rect 433 405 434 406 
<< m1 >>
rect 435 405 436 406 
<< m1 >>
rect 448 405 449 406 
<< m1 >>
rect 462 405 463 406 
<< m1 >>
rect 470 405 471 406 
<< m1 >>
rect 472 405 473 406 
<< m1 >>
rect 474 405 475 406 
<< m1 >>
rect 476 405 477 406 
<< m1 >>
rect 481 405 482 406 
<< m1 >>
rect 489 405 490 406 
<< m2 >>
rect 490 405 491 406 
<< m1 >>
rect 19 406 20 407 
<< m2 >>
rect 20 406 21 407 
<< m1 >>
rect 23 406 24 407 
<< m1 >>
rect 26 406 27 407 
<< m1 >>
rect 37 406 38 407 
<< m1 >>
rect 44 406 45 407 
<< m1 >>
rect 64 406 65 407 
<< m1 >>
rect 73 406 74 407 
<< m2 >>
rect 73 406 74 407 
<< m1 >>
rect 82 406 83 407 
<< m1 >>
rect 88 406 89 407 
<< m2 >>
rect 93 406 94 407 
<< m2 >>
rect 99 406 100 407 
<< m1 >>
rect 103 406 104 407 
<< m1 >>
rect 110 406 111 407 
<< m1 >>
rect 114 406 115 407 
<< m1 >>
rect 121 406 122 407 
<< m1 >>
rect 136 406 137 407 
<< m1 >>
rect 150 406 151 407 
<< m1 >>
rect 157 406 158 407 
<< m1 >>
rect 169 406 170 407 
<< m1 >>
rect 178 406 179 407 
<< m1 >>
rect 181 406 182 407 
<< m1 >>
rect 196 406 197 407 
<< m1 >>
rect 197 406 198 407 
<< m1 >>
rect 198 406 199 407 
<< m1 >>
rect 199 406 200 407 
<< m2 >>
rect 199 406 200 407 
<< m1 >>
rect 200 406 201 407 
<< m1 >>
rect 201 406 202 407 
<< m1 >>
rect 202 406 203 407 
<< m1 >>
rect 203 406 204 407 
<< m1 >>
rect 204 406 205 407 
<< m1 >>
rect 205 406 206 407 
<< m1 >>
rect 206 406 207 407 
<< m2 >>
rect 206 406 207 407 
<< m2c >>
rect 206 406 207 407 
<< m1 >>
rect 206 406 207 407 
<< m2 >>
rect 206 406 207 407 
<< m2 >>
rect 207 406 208 407 
<< m1 >>
rect 208 406 209 407 
<< m2 >>
rect 208 406 209 407 
<< m2 >>
rect 209 406 210 407 
<< m1 >>
rect 210 406 211 407 
<< m2 >>
rect 210 406 211 407 
<< m2c >>
rect 210 406 211 407 
<< m1 >>
rect 210 406 211 407 
<< m2 >>
rect 210 406 211 407 
<< m1 >>
rect 217 406 218 407 
<< m1 >>
rect 229 406 230 407 
<< m1 >>
rect 235 406 236 407 
<< m1 >>
rect 253 406 254 407 
<< m1 >>
rect 280 406 281 407 
<< m2 >>
rect 304 406 305 407 
<< m1 >>
rect 307 406 308 407 
<< m1 >>
rect 314 406 315 407 
<< m1 >>
rect 316 406 317 407 
<< m1 >>
rect 325 406 326 407 
<< m1 >>
rect 329 406 330 407 
<< m1 >>
rect 340 406 341 407 
<< m1 >>
rect 357 406 358 407 
<< m1 >>
rect 361 406 362 407 
<< m1 >>
rect 363 406 364 407 
<< m1 >>
rect 367 406 368 407 
<< m1 >>
rect 379 406 380 407 
<< m2 >>
rect 383 406 384 407 
<< m2 >>
rect 385 406 386 407 
<< m1 >>
rect 391 406 392 407 
<< m1 >>
rect 394 406 395 407 
<< m1 >>
rect 395 406 396 407 
<< m1 >>
rect 396 406 397 407 
<< m1 >>
rect 397 406 398 407 
<< m1 >>
rect 398 406 399 407 
<< m1 >>
rect 399 406 400 407 
<< m1 >>
rect 400 406 401 407 
<< m1 >>
rect 402 406 403 407 
<< m1 >>
rect 406 406 407 407 
<< m1 >>
rect 409 406 410 407 
<< m1 >>
rect 414 406 415 407 
<< m2 >>
rect 414 406 415 407 
<< m2c >>
rect 414 406 415 407 
<< m1 >>
rect 414 406 415 407 
<< m2 >>
rect 414 406 415 407 
<< m2 >>
rect 415 406 416 407 
<< m1 >>
rect 416 406 417 407 
<< m2 >>
rect 416 406 417 407 
<< m2 >>
rect 417 406 418 407 
<< m1 >>
rect 424 406 425 407 
<< m1 >>
rect 433 406 434 407 
<< m1 >>
rect 435 406 436 407 
<< m1 >>
rect 448 406 449 407 
<< m1 >>
rect 462 406 463 407 
<< m1 >>
rect 463 406 464 407 
<< m1 >>
rect 470 406 471 407 
<< m1 >>
rect 472 406 473 407 
<< m1 >>
rect 474 406 475 407 
<< m1 >>
rect 476 406 477 407 
<< m1 >>
rect 481 406 482 407 
<< m1 >>
rect 489 406 490 407 
<< m2 >>
rect 490 406 491 407 
<< m1 >>
rect 19 407 20 408 
<< m2 >>
rect 20 407 21 408 
<< m1 >>
rect 23 407 24 408 
<< m1 >>
rect 26 407 27 408 
<< m1 >>
rect 37 407 38 408 
<< m1 >>
rect 44 407 45 408 
<< m1 >>
rect 64 407 65 408 
<< m1 >>
rect 73 407 74 408 
<< m2 >>
rect 73 407 74 408 
<< m1 >>
rect 82 407 83 408 
<< m1 >>
rect 88 407 89 408 
<< m1 >>
rect 93 407 94 408 
<< m2 >>
rect 93 407 94 408 
<< m2c >>
rect 93 407 94 408 
<< m1 >>
rect 93 407 94 408 
<< m2 >>
rect 93 407 94 408 
<< m1 >>
rect 96 407 97 408 
<< m1 >>
rect 97 407 98 408 
<< m1 >>
rect 98 407 99 408 
<< m1 >>
rect 99 407 100 408 
<< m2 >>
rect 99 407 100 408 
<< m2c >>
rect 99 407 100 408 
<< m1 >>
rect 99 407 100 408 
<< m2 >>
rect 99 407 100 408 
<< m1 >>
rect 103 407 104 408 
<< m1 >>
rect 110 407 111 408 
<< m1 >>
rect 114 407 115 408 
<< m1 >>
rect 121 407 122 408 
<< m1 >>
rect 136 407 137 408 
<< m1 >>
rect 150 407 151 408 
<< m1 >>
rect 157 407 158 408 
<< m1 >>
rect 169 407 170 408 
<< m1 >>
rect 178 407 179 408 
<< m1 >>
rect 181 407 182 408 
<< m1 >>
rect 196 407 197 408 
<< m2 >>
rect 199 407 200 408 
<< m1 >>
rect 208 407 209 408 
<< m1 >>
rect 217 407 218 408 
<< m1 >>
rect 229 407 230 408 
<< m1 >>
rect 235 407 236 408 
<< m1 >>
rect 253 407 254 408 
<< m1 >>
rect 280 407 281 408 
<< m1 >>
rect 304 407 305 408 
<< m2 >>
rect 304 407 305 408 
<< m2c >>
rect 304 407 305 408 
<< m1 >>
rect 304 407 305 408 
<< m2 >>
rect 304 407 305 408 
<< m1 >>
rect 307 407 308 408 
<< m1 >>
rect 314 407 315 408 
<< m1 >>
rect 316 407 317 408 
<< m1 >>
rect 325 407 326 408 
<< m1 >>
rect 329 407 330 408 
<< m1 >>
rect 340 407 341 408 
<< m1 >>
rect 357 407 358 408 
<< m1 >>
rect 361 407 362 408 
<< m1 >>
rect 363 407 364 408 
<< m1 >>
rect 367 407 368 408 
<< m1 >>
rect 379 407 380 408 
<< m1 >>
rect 383 407 384 408 
<< m2 >>
rect 383 407 384 408 
<< m2c >>
rect 383 407 384 408 
<< m1 >>
rect 383 407 384 408 
<< m2 >>
rect 383 407 384 408 
<< m1 >>
rect 385 407 386 408 
<< m2 >>
rect 385 407 386 408 
<< m2c >>
rect 385 407 386 408 
<< m1 >>
rect 385 407 386 408 
<< m2 >>
rect 385 407 386 408 
<< m1 >>
rect 391 407 392 408 
<< m1 >>
rect 394 407 395 408 
<< m1 >>
rect 400 407 401 408 
<< m1 >>
rect 402 407 403 408 
<< m1 >>
rect 406 407 407 408 
<< m1 >>
rect 409 407 410 408 
<< m1 >>
rect 416 407 417 408 
<< m2 >>
rect 417 407 418 408 
<< m1 >>
rect 424 407 425 408 
<< m1 >>
rect 433 407 434 408 
<< m1 >>
rect 435 407 436 408 
<< m1 >>
rect 448 407 449 408 
<< m1 >>
rect 463 407 464 408 
<< m1 >>
rect 470 407 471 408 
<< m1 >>
rect 472 407 473 408 
<< m1 >>
rect 474 407 475 408 
<< m1 >>
rect 476 407 477 408 
<< m1 >>
rect 481 407 482 408 
<< m1 >>
rect 489 407 490 408 
<< m2 >>
rect 490 407 491 408 
<< pdiffusion >>
rect 12 408 13 409 
<< pdiffusion >>
rect 13 408 14 409 
<< pdiffusion >>
rect 14 408 15 409 
<< pdiffusion >>
rect 15 408 16 409 
<< pdiffusion >>
rect 16 408 17 409 
<< pdiffusion >>
rect 17 408 18 409 
<< m1 >>
rect 19 408 20 409 
<< m2 >>
rect 20 408 21 409 
<< m1 >>
rect 23 408 24 409 
<< m1 >>
rect 26 408 27 409 
<< pdiffusion >>
rect 30 408 31 409 
<< pdiffusion >>
rect 31 408 32 409 
<< pdiffusion >>
rect 32 408 33 409 
<< pdiffusion >>
rect 33 408 34 409 
<< pdiffusion >>
rect 34 408 35 409 
<< pdiffusion >>
rect 35 408 36 409 
<< m1 >>
rect 37 408 38 409 
<< m1 >>
rect 44 408 45 409 
<< pdiffusion >>
rect 48 408 49 409 
<< pdiffusion >>
rect 49 408 50 409 
<< pdiffusion >>
rect 50 408 51 409 
<< pdiffusion >>
rect 51 408 52 409 
<< pdiffusion >>
rect 52 408 53 409 
<< pdiffusion >>
rect 53 408 54 409 
<< m1 >>
rect 64 408 65 409 
<< pdiffusion >>
rect 66 408 67 409 
<< pdiffusion >>
rect 67 408 68 409 
<< pdiffusion >>
rect 68 408 69 409 
<< pdiffusion >>
rect 69 408 70 409 
<< pdiffusion >>
rect 70 408 71 409 
<< pdiffusion >>
rect 71 408 72 409 
<< m1 >>
rect 73 408 74 409 
<< m2 >>
rect 73 408 74 409 
<< m1 >>
rect 82 408 83 409 
<< pdiffusion >>
rect 84 408 85 409 
<< pdiffusion >>
rect 85 408 86 409 
<< pdiffusion >>
rect 86 408 87 409 
<< pdiffusion >>
rect 87 408 88 409 
<< m1 >>
rect 88 408 89 409 
<< pdiffusion >>
rect 88 408 89 409 
<< pdiffusion >>
rect 89 408 90 409 
<< m1 >>
rect 93 408 94 409 
<< m1 >>
rect 96 408 97 409 
<< pdiffusion >>
rect 102 408 103 409 
<< m1 >>
rect 103 408 104 409 
<< pdiffusion >>
rect 103 408 104 409 
<< pdiffusion >>
rect 104 408 105 409 
<< pdiffusion >>
rect 105 408 106 409 
<< pdiffusion >>
rect 106 408 107 409 
<< pdiffusion >>
rect 107 408 108 409 
<< m1 >>
rect 110 408 111 409 
<< m1 >>
rect 114 408 115 409 
<< pdiffusion >>
rect 120 408 121 409 
<< m1 >>
rect 121 408 122 409 
<< pdiffusion >>
rect 121 408 122 409 
<< pdiffusion >>
rect 122 408 123 409 
<< pdiffusion >>
rect 123 408 124 409 
<< pdiffusion >>
rect 124 408 125 409 
<< pdiffusion >>
rect 125 408 126 409 
<< m1 >>
rect 136 408 137 409 
<< pdiffusion >>
rect 138 408 139 409 
<< pdiffusion >>
rect 139 408 140 409 
<< pdiffusion >>
rect 140 408 141 409 
<< pdiffusion >>
rect 141 408 142 409 
<< pdiffusion >>
rect 142 408 143 409 
<< pdiffusion >>
rect 143 408 144 409 
<< m1 >>
rect 150 408 151 409 
<< m1 >>
rect 157 408 158 409 
<< m1 >>
rect 169 408 170 409 
<< pdiffusion >>
rect 174 408 175 409 
<< pdiffusion >>
rect 175 408 176 409 
<< pdiffusion >>
rect 176 408 177 409 
<< pdiffusion >>
rect 177 408 178 409 
<< m1 >>
rect 178 408 179 409 
<< pdiffusion >>
rect 178 408 179 409 
<< pdiffusion >>
rect 179 408 180 409 
<< m1 >>
rect 181 408 182 409 
<< pdiffusion >>
rect 192 408 193 409 
<< pdiffusion >>
rect 193 408 194 409 
<< pdiffusion >>
rect 194 408 195 409 
<< pdiffusion >>
rect 195 408 196 409 
<< m1 >>
rect 196 408 197 409 
<< pdiffusion >>
rect 196 408 197 409 
<< pdiffusion >>
rect 197 408 198 409 
<< m1 >>
rect 199 408 200 409 
<< m2 >>
rect 199 408 200 409 
<< m2c >>
rect 199 408 200 409 
<< m1 >>
rect 199 408 200 409 
<< m2 >>
rect 199 408 200 409 
<< m1 >>
rect 208 408 209 409 
<< pdiffusion >>
rect 210 408 211 409 
<< pdiffusion >>
rect 211 408 212 409 
<< pdiffusion >>
rect 212 408 213 409 
<< pdiffusion >>
rect 213 408 214 409 
<< pdiffusion >>
rect 214 408 215 409 
<< pdiffusion >>
rect 215 408 216 409 
<< m1 >>
rect 217 408 218 409 
<< pdiffusion >>
rect 228 408 229 409 
<< m1 >>
rect 229 408 230 409 
<< pdiffusion >>
rect 229 408 230 409 
<< pdiffusion >>
rect 230 408 231 409 
<< pdiffusion >>
rect 231 408 232 409 
<< pdiffusion >>
rect 232 408 233 409 
<< pdiffusion >>
rect 233 408 234 409 
<< m1 >>
rect 235 408 236 409 
<< pdiffusion >>
rect 246 408 247 409 
<< pdiffusion >>
rect 247 408 248 409 
<< pdiffusion >>
rect 248 408 249 409 
<< pdiffusion >>
rect 249 408 250 409 
<< pdiffusion >>
rect 250 408 251 409 
<< pdiffusion >>
rect 251 408 252 409 
<< m1 >>
rect 253 408 254 409 
<< pdiffusion >>
rect 264 408 265 409 
<< pdiffusion >>
rect 265 408 266 409 
<< pdiffusion >>
rect 266 408 267 409 
<< pdiffusion >>
rect 267 408 268 409 
<< pdiffusion >>
rect 268 408 269 409 
<< pdiffusion >>
rect 269 408 270 409 
<< m1 >>
rect 280 408 281 409 
<< pdiffusion >>
rect 282 408 283 409 
<< pdiffusion >>
rect 283 408 284 409 
<< pdiffusion >>
rect 284 408 285 409 
<< pdiffusion >>
rect 285 408 286 409 
<< pdiffusion >>
rect 286 408 287 409 
<< pdiffusion >>
rect 287 408 288 409 
<< pdiffusion >>
rect 300 408 301 409 
<< pdiffusion >>
rect 301 408 302 409 
<< pdiffusion >>
rect 302 408 303 409 
<< pdiffusion >>
rect 303 408 304 409 
<< m1 >>
rect 304 408 305 409 
<< pdiffusion >>
rect 304 408 305 409 
<< pdiffusion >>
rect 305 408 306 409 
<< m1 >>
rect 307 408 308 409 
<< m1 >>
rect 314 408 315 409 
<< m1 >>
rect 316 408 317 409 
<< pdiffusion >>
rect 318 408 319 409 
<< pdiffusion >>
rect 319 408 320 409 
<< pdiffusion >>
rect 320 408 321 409 
<< pdiffusion >>
rect 321 408 322 409 
<< pdiffusion >>
rect 322 408 323 409 
<< pdiffusion >>
rect 323 408 324 409 
<< m1 >>
rect 325 408 326 409 
<< m1 >>
rect 329 408 330 409 
<< pdiffusion >>
rect 336 408 337 409 
<< pdiffusion >>
rect 337 408 338 409 
<< pdiffusion >>
rect 338 408 339 409 
<< pdiffusion >>
rect 339 408 340 409 
<< m1 >>
rect 340 408 341 409 
<< pdiffusion >>
rect 340 408 341 409 
<< pdiffusion >>
rect 341 408 342 409 
<< m1 >>
rect 357 408 358 409 
<< m1 >>
rect 361 408 362 409 
<< m1 >>
rect 363 408 364 409 
<< m1 >>
rect 367 408 368 409 
<< pdiffusion >>
rect 372 408 373 409 
<< pdiffusion >>
rect 373 408 374 409 
<< pdiffusion >>
rect 374 408 375 409 
<< pdiffusion >>
rect 375 408 376 409 
<< pdiffusion >>
rect 376 408 377 409 
<< pdiffusion >>
rect 377 408 378 409 
<< m1 >>
rect 379 408 380 409 
<< m1 >>
rect 383 408 384 409 
<< m1 >>
rect 385 408 386 409 
<< pdiffusion >>
rect 390 408 391 409 
<< m1 >>
rect 391 408 392 409 
<< pdiffusion >>
rect 391 408 392 409 
<< pdiffusion >>
rect 392 408 393 409 
<< pdiffusion >>
rect 393 408 394 409 
<< m1 >>
rect 394 408 395 409 
<< pdiffusion >>
rect 394 408 395 409 
<< pdiffusion >>
rect 395 408 396 409 
<< m1 >>
rect 400 408 401 409 
<< m1 >>
rect 402 408 403 409 
<< m1 >>
rect 406 408 407 409 
<< pdiffusion >>
rect 408 408 409 409 
<< m1 >>
rect 409 408 410 409 
<< pdiffusion >>
rect 409 408 410 409 
<< pdiffusion >>
rect 410 408 411 409 
<< pdiffusion >>
rect 411 408 412 409 
<< pdiffusion >>
rect 412 408 413 409 
<< pdiffusion >>
rect 413 408 414 409 
<< m1 >>
rect 416 408 417 409 
<< m2 >>
rect 417 408 418 409 
<< m1 >>
rect 424 408 425 409 
<< pdiffusion >>
rect 426 408 427 409 
<< pdiffusion >>
rect 427 408 428 409 
<< pdiffusion >>
rect 428 408 429 409 
<< pdiffusion >>
rect 429 408 430 409 
<< pdiffusion >>
rect 430 408 431 409 
<< pdiffusion >>
rect 431 408 432 409 
<< m1 >>
rect 433 408 434 409 
<< m1 >>
rect 435 408 436 409 
<< pdiffusion >>
rect 444 408 445 409 
<< pdiffusion >>
rect 445 408 446 409 
<< pdiffusion >>
rect 446 408 447 409 
<< pdiffusion >>
rect 447 408 448 409 
<< m1 >>
rect 448 408 449 409 
<< pdiffusion >>
rect 448 408 449 409 
<< pdiffusion >>
rect 449 408 450 409 
<< pdiffusion >>
rect 462 408 463 409 
<< m1 >>
rect 463 408 464 409 
<< pdiffusion >>
rect 463 408 464 409 
<< pdiffusion >>
rect 464 408 465 409 
<< pdiffusion >>
rect 465 408 466 409 
<< pdiffusion >>
rect 466 408 467 409 
<< pdiffusion >>
rect 467 408 468 409 
<< m1 >>
rect 470 408 471 409 
<< m1 >>
rect 472 408 473 409 
<< m1 >>
rect 474 408 475 409 
<< m1 >>
rect 476 408 477 409 
<< pdiffusion >>
rect 480 408 481 409 
<< m1 >>
rect 481 408 482 409 
<< pdiffusion >>
rect 481 408 482 409 
<< pdiffusion >>
rect 482 408 483 409 
<< pdiffusion >>
rect 483 408 484 409 
<< pdiffusion >>
rect 484 408 485 409 
<< pdiffusion >>
rect 485 408 486 409 
<< m1 >>
rect 489 408 490 409 
<< m2 >>
rect 490 408 491 409 
<< pdiffusion >>
rect 498 408 499 409 
<< pdiffusion >>
rect 499 408 500 409 
<< pdiffusion >>
rect 500 408 501 409 
<< pdiffusion >>
rect 501 408 502 409 
<< pdiffusion >>
rect 502 408 503 409 
<< pdiffusion >>
rect 503 408 504 409 
<< pdiffusion >>
rect 516 408 517 409 
<< pdiffusion >>
rect 517 408 518 409 
<< pdiffusion >>
rect 518 408 519 409 
<< pdiffusion >>
rect 519 408 520 409 
<< pdiffusion >>
rect 520 408 521 409 
<< pdiffusion >>
rect 521 408 522 409 
<< pdiffusion >>
rect 12 409 13 410 
<< pdiffusion >>
rect 13 409 14 410 
<< pdiffusion >>
rect 14 409 15 410 
<< pdiffusion >>
rect 15 409 16 410 
<< pdiffusion >>
rect 16 409 17 410 
<< pdiffusion >>
rect 17 409 18 410 
<< m1 >>
rect 19 409 20 410 
<< m2 >>
rect 20 409 21 410 
<< m1 >>
rect 23 409 24 410 
<< m1 >>
rect 26 409 27 410 
<< pdiffusion >>
rect 30 409 31 410 
<< pdiffusion >>
rect 31 409 32 410 
<< pdiffusion >>
rect 32 409 33 410 
<< pdiffusion >>
rect 33 409 34 410 
<< pdiffusion >>
rect 34 409 35 410 
<< pdiffusion >>
rect 35 409 36 410 
<< m1 >>
rect 37 409 38 410 
<< m1 >>
rect 44 409 45 410 
<< pdiffusion >>
rect 48 409 49 410 
<< pdiffusion >>
rect 49 409 50 410 
<< pdiffusion >>
rect 50 409 51 410 
<< pdiffusion >>
rect 51 409 52 410 
<< pdiffusion >>
rect 52 409 53 410 
<< pdiffusion >>
rect 53 409 54 410 
<< m1 >>
rect 64 409 65 410 
<< pdiffusion >>
rect 66 409 67 410 
<< pdiffusion >>
rect 67 409 68 410 
<< pdiffusion >>
rect 68 409 69 410 
<< pdiffusion >>
rect 69 409 70 410 
<< pdiffusion >>
rect 70 409 71 410 
<< pdiffusion >>
rect 71 409 72 410 
<< m1 >>
rect 73 409 74 410 
<< m2 >>
rect 73 409 74 410 
<< m1 >>
rect 82 409 83 410 
<< pdiffusion >>
rect 84 409 85 410 
<< pdiffusion >>
rect 85 409 86 410 
<< pdiffusion >>
rect 86 409 87 410 
<< pdiffusion >>
rect 87 409 88 410 
<< pdiffusion >>
rect 88 409 89 410 
<< pdiffusion >>
rect 89 409 90 410 
<< m1 >>
rect 93 409 94 410 
<< m1 >>
rect 96 409 97 410 
<< pdiffusion >>
rect 102 409 103 410 
<< pdiffusion >>
rect 103 409 104 410 
<< pdiffusion >>
rect 104 409 105 410 
<< pdiffusion >>
rect 105 409 106 410 
<< pdiffusion >>
rect 106 409 107 410 
<< pdiffusion >>
rect 107 409 108 410 
<< m1 >>
rect 110 409 111 410 
<< m1 >>
rect 114 409 115 410 
<< pdiffusion >>
rect 120 409 121 410 
<< pdiffusion >>
rect 121 409 122 410 
<< pdiffusion >>
rect 122 409 123 410 
<< pdiffusion >>
rect 123 409 124 410 
<< pdiffusion >>
rect 124 409 125 410 
<< pdiffusion >>
rect 125 409 126 410 
<< m1 >>
rect 136 409 137 410 
<< pdiffusion >>
rect 138 409 139 410 
<< pdiffusion >>
rect 139 409 140 410 
<< pdiffusion >>
rect 140 409 141 410 
<< pdiffusion >>
rect 141 409 142 410 
<< pdiffusion >>
rect 142 409 143 410 
<< pdiffusion >>
rect 143 409 144 410 
<< m1 >>
rect 150 409 151 410 
<< m1 >>
rect 157 409 158 410 
<< m1 >>
rect 169 409 170 410 
<< pdiffusion >>
rect 174 409 175 410 
<< pdiffusion >>
rect 175 409 176 410 
<< pdiffusion >>
rect 176 409 177 410 
<< pdiffusion >>
rect 177 409 178 410 
<< pdiffusion >>
rect 178 409 179 410 
<< pdiffusion >>
rect 179 409 180 410 
<< m1 >>
rect 181 409 182 410 
<< pdiffusion >>
rect 192 409 193 410 
<< pdiffusion >>
rect 193 409 194 410 
<< pdiffusion >>
rect 194 409 195 410 
<< pdiffusion >>
rect 195 409 196 410 
<< pdiffusion >>
rect 196 409 197 410 
<< pdiffusion >>
rect 197 409 198 410 
<< m1 >>
rect 199 409 200 410 
<< m1 >>
rect 208 409 209 410 
<< pdiffusion >>
rect 210 409 211 410 
<< pdiffusion >>
rect 211 409 212 410 
<< pdiffusion >>
rect 212 409 213 410 
<< pdiffusion >>
rect 213 409 214 410 
<< pdiffusion >>
rect 214 409 215 410 
<< pdiffusion >>
rect 215 409 216 410 
<< m1 >>
rect 217 409 218 410 
<< pdiffusion >>
rect 228 409 229 410 
<< pdiffusion >>
rect 229 409 230 410 
<< pdiffusion >>
rect 230 409 231 410 
<< pdiffusion >>
rect 231 409 232 410 
<< pdiffusion >>
rect 232 409 233 410 
<< pdiffusion >>
rect 233 409 234 410 
<< m1 >>
rect 235 409 236 410 
<< pdiffusion >>
rect 246 409 247 410 
<< pdiffusion >>
rect 247 409 248 410 
<< pdiffusion >>
rect 248 409 249 410 
<< pdiffusion >>
rect 249 409 250 410 
<< pdiffusion >>
rect 250 409 251 410 
<< pdiffusion >>
rect 251 409 252 410 
<< m1 >>
rect 253 409 254 410 
<< pdiffusion >>
rect 264 409 265 410 
<< pdiffusion >>
rect 265 409 266 410 
<< pdiffusion >>
rect 266 409 267 410 
<< pdiffusion >>
rect 267 409 268 410 
<< pdiffusion >>
rect 268 409 269 410 
<< pdiffusion >>
rect 269 409 270 410 
<< m1 >>
rect 280 409 281 410 
<< pdiffusion >>
rect 282 409 283 410 
<< pdiffusion >>
rect 283 409 284 410 
<< pdiffusion >>
rect 284 409 285 410 
<< pdiffusion >>
rect 285 409 286 410 
<< pdiffusion >>
rect 286 409 287 410 
<< pdiffusion >>
rect 287 409 288 410 
<< pdiffusion >>
rect 300 409 301 410 
<< pdiffusion >>
rect 301 409 302 410 
<< pdiffusion >>
rect 302 409 303 410 
<< pdiffusion >>
rect 303 409 304 410 
<< pdiffusion >>
rect 304 409 305 410 
<< pdiffusion >>
rect 305 409 306 410 
<< m1 >>
rect 307 409 308 410 
<< m1 >>
rect 314 409 315 410 
<< m1 >>
rect 316 409 317 410 
<< pdiffusion >>
rect 318 409 319 410 
<< pdiffusion >>
rect 319 409 320 410 
<< pdiffusion >>
rect 320 409 321 410 
<< pdiffusion >>
rect 321 409 322 410 
<< pdiffusion >>
rect 322 409 323 410 
<< pdiffusion >>
rect 323 409 324 410 
<< m1 >>
rect 325 409 326 410 
<< m1 >>
rect 329 409 330 410 
<< pdiffusion >>
rect 336 409 337 410 
<< pdiffusion >>
rect 337 409 338 410 
<< pdiffusion >>
rect 338 409 339 410 
<< pdiffusion >>
rect 339 409 340 410 
<< pdiffusion >>
rect 340 409 341 410 
<< pdiffusion >>
rect 341 409 342 410 
<< m1 >>
rect 357 409 358 410 
<< m1 >>
rect 361 409 362 410 
<< m1 >>
rect 363 409 364 410 
<< m1 >>
rect 367 409 368 410 
<< pdiffusion >>
rect 372 409 373 410 
<< pdiffusion >>
rect 373 409 374 410 
<< pdiffusion >>
rect 374 409 375 410 
<< pdiffusion >>
rect 375 409 376 410 
<< pdiffusion >>
rect 376 409 377 410 
<< pdiffusion >>
rect 377 409 378 410 
<< m1 >>
rect 379 409 380 410 
<< m1 >>
rect 383 409 384 410 
<< m1 >>
rect 385 409 386 410 
<< pdiffusion >>
rect 390 409 391 410 
<< pdiffusion >>
rect 391 409 392 410 
<< pdiffusion >>
rect 392 409 393 410 
<< pdiffusion >>
rect 393 409 394 410 
<< pdiffusion >>
rect 394 409 395 410 
<< pdiffusion >>
rect 395 409 396 410 
<< m1 >>
rect 400 409 401 410 
<< m1 >>
rect 402 409 403 410 
<< m1 >>
rect 406 409 407 410 
<< pdiffusion >>
rect 408 409 409 410 
<< pdiffusion >>
rect 409 409 410 410 
<< pdiffusion >>
rect 410 409 411 410 
<< pdiffusion >>
rect 411 409 412 410 
<< pdiffusion >>
rect 412 409 413 410 
<< pdiffusion >>
rect 413 409 414 410 
<< m1 >>
rect 416 409 417 410 
<< m2 >>
rect 417 409 418 410 
<< m1 >>
rect 424 409 425 410 
<< pdiffusion >>
rect 426 409 427 410 
<< pdiffusion >>
rect 427 409 428 410 
<< pdiffusion >>
rect 428 409 429 410 
<< pdiffusion >>
rect 429 409 430 410 
<< pdiffusion >>
rect 430 409 431 410 
<< pdiffusion >>
rect 431 409 432 410 
<< m1 >>
rect 433 409 434 410 
<< m1 >>
rect 435 409 436 410 
<< pdiffusion >>
rect 444 409 445 410 
<< pdiffusion >>
rect 445 409 446 410 
<< pdiffusion >>
rect 446 409 447 410 
<< pdiffusion >>
rect 447 409 448 410 
<< pdiffusion >>
rect 448 409 449 410 
<< pdiffusion >>
rect 449 409 450 410 
<< pdiffusion >>
rect 462 409 463 410 
<< pdiffusion >>
rect 463 409 464 410 
<< pdiffusion >>
rect 464 409 465 410 
<< pdiffusion >>
rect 465 409 466 410 
<< pdiffusion >>
rect 466 409 467 410 
<< pdiffusion >>
rect 467 409 468 410 
<< m1 >>
rect 470 409 471 410 
<< m1 >>
rect 472 409 473 410 
<< m1 >>
rect 474 409 475 410 
<< m1 >>
rect 476 409 477 410 
<< pdiffusion >>
rect 480 409 481 410 
<< pdiffusion >>
rect 481 409 482 410 
<< pdiffusion >>
rect 482 409 483 410 
<< pdiffusion >>
rect 483 409 484 410 
<< pdiffusion >>
rect 484 409 485 410 
<< pdiffusion >>
rect 485 409 486 410 
<< m1 >>
rect 489 409 490 410 
<< m2 >>
rect 490 409 491 410 
<< pdiffusion >>
rect 498 409 499 410 
<< pdiffusion >>
rect 499 409 500 410 
<< pdiffusion >>
rect 500 409 501 410 
<< pdiffusion >>
rect 501 409 502 410 
<< pdiffusion >>
rect 502 409 503 410 
<< pdiffusion >>
rect 503 409 504 410 
<< pdiffusion >>
rect 516 409 517 410 
<< pdiffusion >>
rect 517 409 518 410 
<< pdiffusion >>
rect 518 409 519 410 
<< pdiffusion >>
rect 519 409 520 410 
<< pdiffusion >>
rect 520 409 521 410 
<< pdiffusion >>
rect 521 409 522 410 
<< pdiffusion >>
rect 12 410 13 411 
<< pdiffusion >>
rect 13 410 14 411 
<< pdiffusion >>
rect 14 410 15 411 
<< pdiffusion >>
rect 15 410 16 411 
<< pdiffusion >>
rect 16 410 17 411 
<< pdiffusion >>
rect 17 410 18 411 
<< m1 >>
rect 19 410 20 411 
<< m2 >>
rect 20 410 21 411 
<< m1 >>
rect 23 410 24 411 
<< m1 >>
rect 26 410 27 411 
<< pdiffusion >>
rect 30 410 31 411 
<< pdiffusion >>
rect 31 410 32 411 
<< pdiffusion >>
rect 32 410 33 411 
<< pdiffusion >>
rect 33 410 34 411 
<< pdiffusion >>
rect 34 410 35 411 
<< pdiffusion >>
rect 35 410 36 411 
<< m1 >>
rect 37 410 38 411 
<< m1 >>
rect 44 410 45 411 
<< pdiffusion >>
rect 48 410 49 411 
<< pdiffusion >>
rect 49 410 50 411 
<< pdiffusion >>
rect 50 410 51 411 
<< pdiffusion >>
rect 51 410 52 411 
<< pdiffusion >>
rect 52 410 53 411 
<< pdiffusion >>
rect 53 410 54 411 
<< m1 >>
rect 64 410 65 411 
<< pdiffusion >>
rect 66 410 67 411 
<< pdiffusion >>
rect 67 410 68 411 
<< pdiffusion >>
rect 68 410 69 411 
<< pdiffusion >>
rect 69 410 70 411 
<< pdiffusion >>
rect 70 410 71 411 
<< pdiffusion >>
rect 71 410 72 411 
<< m1 >>
rect 73 410 74 411 
<< m2 >>
rect 73 410 74 411 
<< m1 >>
rect 82 410 83 411 
<< pdiffusion >>
rect 84 410 85 411 
<< pdiffusion >>
rect 85 410 86 411 
<< pdiffusion >>
rect 86 410 87 411 
<< pdiffusion >>
rect 87 410 88 411 
<< pdiffusion >>
rect 88 410 89 411 
<< pdiffusion >>
rect 89 410 90 411 
<< m1 >>
rect 93 410 94 411 
<< m1 >>
rect 96 410 97 411 
<< pdiffusion >>
rect 102 410 103 411 
<< pdiffusion >>
rect 103 410 104 411 
<< pdiffusion >>
rect 104 410 105 411 
<< pdiffusion >>
rect 105 410 106 411 
<< pdiffusion >>
rect 106 410 107 411 
<< pdiffusion >>
rect 107 410 108 411 
<< m1 >>
rect 110 410 111 411 
<< m1 >>
rect 114 410 115 411 
<< pdiffusion >>
rect 120 410 121 411 
<< pdiffusion >>
rect 121 410 122 411 
<< pdiffusion >>
rect 122 410 123 411 
<< pdiffusion >>
rect 123 410 124 411 
<< pdiffusion >>
rect 124 410 125 411 
<< pdiffusion >>
rect 125 410 126 411 
<< m1 >>
rect 136 410 137 411 
<< pdiffusion >>
rect 138 410 139 411 
<< pdiffusion >>
rect 139 410 140 411 
<< pdiffusion >>
rect 140 410 141 411 
<< pdiffusion >>
rect 141 410 142 411 
<< pdiffusion >>
rect 142 410 143 411 
<< pdiffusion >>
rect 143 410 144 411 
<< m1 >>
rect 150 410 151 411 
<< m1 >>
rect 157 410 158 411 
<< m1 >>
rect 169 410 170 411 
<< pdiffusion >>
rect 174 410 175 411 
<< pdiffusion >>
rect 175 410 176 411 
<< pdiffusion >>
rect 176 410 177 411 
<< pdiffusion >>
rect 177 410 178 411 
<< pdiffusion >>
rect 178 410 179 411 
<< pdiffusion >>
rect 179 410 180 411 
<< m1 >>
rect 181 410 182 411 
<< pdiffusion >>
rect 192 410 193 411 
<< pdiffusion >>
rect 193 410 194 411 
<< pdiffusion >>
rect 194 410 195 411 
<< pdiffusion >>
rect 195 410 196 411 
<< pdiffusion >>
rect 196 410 197 411 
<< pdiffusion >>
rect 197 410 198 411 
<< m1 >>
rect 199 410 200 411 
<< m1 >>
rect 208 410 209 411 
<< pdiffusion >>
rect 210 410 211 411 
<< pdiffusion >>
rect 211 410 212 411 
<< pdiffusion >>
rect 212 410 213 411 
<< pdiffusion >>
rect 213 410 214 411 
<< pdiffusion >>
rect 214 410 215 411 
<< pdiffusion >>
rect 215 410 216 411 
<< m1 >>
rect 217 410 218 411 
<< pdiffusion >>
rect 228 410 229 411 
<< pdiffusion >>
rect 229 410 230 411 
<< pdiffusion >>
rect 230 410 231 411 
<< pdiffusion >>
rect 231 410 232 411 
<< pdiffusion >>
rect 232 410 233 411 
<< pdiffusion >>
rect 233 410 234 411 
<< m1 >>
rect 235 410 236 411 
<< pdiffusion >>
rect 246 410 247 411 
<< pdiffusion >>
rect 247 410 248 411 
<< pdiffusion >>
rect 248 410 249 411 
<< pdiffusion >>
rect 249 410 250 411 
<< pdiffusion >>
rect 250 410 251 411 
<< pdiffusion >>
rect 251 410 252 411 
<< m1 >>
rect 253 410 254 411 
<< pdiffusion >>
rect 264 410 265 411 
<< pdiffusion >>
rect 265 410 266 411 
<< pdiffusion >>
rect 266 410 267 411 
<< pdiffusion >>
rect 267 410 268 411 
<< pdiffusion >>
rect 268 410 269 411 
<< pdiffusion >>
rect 269 410 270 411 
<< m1 >>
rect 280 410 281 411 
<< pdiffusion >>
rect 282 410 283 411 
<< pdiffusion >>
rect 283 410 284 411 
<< pdiffusion >>
rect 284 410 285 411 
<< pdiffusion >>
rect 285 410 286 411 
<< pdiffusion >>
rect 286 410 287 411 
<< pdiffusion >>
rect 287 410 288 411 
<< pdiffusion >>
rect 300 410 301 411 
<< pdiffusion >>
rect 301 410 302 411 
<< pdiffusion >>
rect 302 410 303 411 
<< pdiffusion >>
rect 303 410 304 411 
<< pdiffusion >>
rect 304 410 305 411 
<< pdiffusion >>
rect 305 410 306 411 
<< m1 >>
rect 307 410 308 411 
<< m1 >>
rect 314 410 315 411 
<< m1 >>
rect 316 410 317 411 
<< pdiffusion >>
rect 318 410 319 411 
<< pdiffusion >>
rect 319 410 320 411 
<< pdiffusion >>
rect 320 410 321 411 
<< pdiffusion >>
rect 321 410 322 411 
<< pdiffusion >>
rect 322 410 323 411 
<< pdiffusion >>
rect 323 410 324 411 
<< m1 >>
rect 325 410 326 411 
<< m1 >>
rect 329 410 330 411 
<< pdiffusion >>
rect 336 410 337 411 
<< pdiffusion >>
rect 337 410 338 411 
<< pdiffusion >>
rect 338 410 339 411 
<< pdiffusion >>
rect 339 410 340 411 
<< pdiffusion >>
rect 340 410 341 411 
<< pdiffusion >>
rect 341 410 342 411 
<< m1 >>
rect 357 410 358 411 
<< m1 >>
rect 361 410 362 411 
<< m1 >>
rect 363 410 364 411 
<< m1 >>
rect 367 410 368 411 
<< pdiffusion >>
rect 372 410 373 411 
<< pdiffusion >>
rect 373 410 374 411 
<< pdiffusion >>
rect 374 410 375 411 
<< pdiffusion >>
rect 375 410 376 411 
<< pdiffusion >>
rect 376 410 377 411 
<< pdiffusion >>
rect 377 410 378 411 
<< m1 >>
rect 379 410 380 411 
<< m1 >>
rect 383 410 384 411 
<< m1 >>
rect 385 410 386 411 
<< pdiffusion >>
rect 390 410 391 411 
<< pdiffusion >>
rect 391 410 392 411 
<< pdiffusion >>
rect 392 410 393 411 
<< pdiffusion >>
rect 393 410 394 411 
<< pdiffusion >>
rect 394 410 395 411 
<< pdiffusion >>
rect 395 410 396 411 
<< m1 >>
rect 400 410 401 411 
<< m1 >>
rect 402 410 403 411 
<< m1 >>
rect 406 410 407 411 
<< pdiffusion >>
rect 408 410 409 411 
<< pdiffusion >>
rect 409 410 410 411 
<< pdiffusion >>
rect 410 410 411 411 
<< pdiffusion >>
rect 411 410 412 411 
<< pdiffusion >>
rect 412 410 413 411 
<< pdiffusion >>
rect 413 410 414 411 
<< m1 >>
rect 416 410 417 411 
<< m2 >>
rect 417 410 418 411 
<< m1 >>
rect 424 410 425 411 
<< pdiffusion >>
rect 426 410 427 411 
<< pdiffusion >>
rect 427 410 428 411 
<< pdiffusion >>
rect 428 410 429 411 
<< pdiffusion >>
rect 429 410 430 411 
<< pdiffusion >>
rect 430 410 431 411 
<< pdiffusion >>
rect 431 410 432 411 
<< m1 >>
rect 433 410 434 411 
<< m1 >>
rect 435 410 436 411 
<< pdiffusion >>
rect 444 410 445 411 
<< pdiffusion >>
rect 445 410 446 411 
<< pdiffusion >>
rect 446 410 447 411 
<< pdiffusion >>
rect 447 410 448 411 
<< pdiffusion >>
rect 448 410 449 411 
<< pdiffusion >>
rect 449 410 450 411 
<< pdiffusion >>
rect 462 410 463 411 
<< pdiffusion >>
rect 463 410 464 411 
<< pdiffusion >>
rect 464 410 465 411 
<< pdiffusion >>
rect 465 410 466 411 
<< pdiffusion >>
rect 466 410 467 411 
<< pdiffusion >>
rect 467 410 468 411 
<< m1 >>
rect 470 410 471 411 
<< m1 >>
rect 472 410 473 411 
<< m1 >>
rect 474 410 475 411 
<< m1 >>
rect 476 410 477 411 
<< pdiffusion >>
rect 480 410 481 411 
<< pdiffusion >>
rect 481 410 482 411 
<< pdiffusion >>
rect 482 410 483 411 
<< pdiffusion >>
rect 483 410 484 411 
<< pdiffusion >>
rect 484 410 485 411 
<< pdiffusion >>
rect 485 410 486 411 
<< m1 >>
rect 489 410 490 411 
<< m2 >>
rect 490 410 491 411 
<< pdiffusion >>
rect 498 410 499 411 
<< pdiffusion >>
rect 499 410 500 411 
<< pdiffusion >>
rect 500 410 501 411 
<< pdiffusion >>
rect 501 410 502 411 
<< pdiffusion >>
rect 502 410 503 411 
<< pdiffusion >>
rect 503 410 504 411 
<< pdiffusion >>
rect 516 410 517 411 
<< pdiffusion >>
rect 517 410 518 411 
<< pdiffusion >>
rect 518 410 519 411 
<< pdiffusion >>
rect 519 410 520 411 
<< pdiffusion >>
rect 520 410 521 411 
<< pdiffusion >>
rect 521 410 522 411 
<< pdiffusion >>
rect 12 411 13 412 
<< pdiffusion >>
rect 13 411 14 412 
<< pdiffusion >>
rect 14 411 15 412 
<< pdiffusion >>
rect 15 411 16 412 
<< pdiffusion >>
rect 16 411 17 412 
<< pdiffusion >>
rect 17 411 18 412 
<< m1 >>
rect 19 411 20 412 
<< m2 >>
rect 20 411 21 412 
<< m1 >>
rect 23 411 24 412 
<< m1 >>
rect 26 411 27 412 
<< pdiffusion >>
rect 30 411 31 412 
<< pdiffusion >>
rect 31 411 32 412 
<< pdiffusion >>
rect 32 411 33 412 
<< pdiffusion >>
rect 33 411 34 412 
<< pdiffusion >>
rect 34 411 35 412 
<< pdiffusion >>
rect 35 411 36 412 
<< m1 >>
rect 37 411 38 412 
<< m1 >>
rect 44 411 45 412 
<< pdiffusion >>
rect 48 411 49 412 
<< pdiffusion >>
rect 49 411 50 412 
<< pdiffusion >>
rect 50 411 51 412 
<< pdiffusion >>
rect 51 411 52 412 
<< pdiffusion >>
rect 52 411 53 412 
<< pdiffusion >>
rect 53 411 54 412 
<< m1 >>
rect 64 411 65 412 
<< pdiffusion >>
rect 66 411 67 412 
<< pdiffusion >>
rect 67 411 68 412 
<< pdiffusion >>
rect 68 411 69 412 
<< pdiffusion >>
rect 69 411 70 412 
<< pdiffusion >>
rect 70 411 71 412 
<< pdiffusion >>
rect 71 411 72 412 
<< m1 >>
rect 73 411 74 412 
<< m2 >>
rect 73 411 74 412 
<< m1 >>
rect 82 411 83 412 
<< pdiffusion >>
rect 84 411 85 412 
<< pdiffusion >>
rect 85 411 86 412 
<< pdiffusion >>
rect 86 411 87 412 
<< pdiffusion >>
rect 87 411 88 412 
<< pdiffusion >>
rect 88 411 89 412 
<< pdiffusion >>
rect 89 411 90 412 
<< m1 >>
rect 93 411 94 412 
<< m1 >>
rect 96 411 97 412 
<< pdiffusion >>
rect 102 411 103 412 
<< pdiffusion >>
rect 103 411 104 412 
<< pdiffusion >>
rect 104 411 105 412 
<< pdiffusion >>
rect 105 411 106 412 
<< pdiffusion >>
rect 106 411 107 412 
<< pdiffusion >>
rect 107 411 108 412 
<< m1 >>
rect 110 411 111 412 
<< m1 >>
rect 114 411 115 412 
<< pdiffusion >>
rect 120 411 121 412 
<< pdiffusion >>
rect 121 411 122 412 
<< pdiffusion >>
rect 122 411 123 412 
<< pdiffusion >>
rect 123 411 124 412 
<< pdiffusion >>
rect 124 411 125 412 
<< pdiffusion >>
rect 125 411 126 412 
<< m1 >>
rect 136 411 137 412 
<< pdiffusion >>
rect 138 411 139 412 
<< pdiffusion >>
rect 139 411 140 412 
<< pdiffusion >>
rect 140 411 141 412 
<< pdiffusion >>
rect 141 411 142 412 
<< pdiffusion >>
rect 142 411 143 412 
<< pdiffusion >>
rect 143 411 144 412 
<< m1 >>
rect 150 411 151 412 
<< m1 >>
rect 157 411 158 412 
<< m1 >>
rect 169 411 170 412 
<< pdiffusion >>
rect 174 411 175 412 
<< pdiffusion >>
rect 175 411 176 412 
<< pdiffusion >>
rect 176 411 177 412 
<< pdiffusion >>
rect 177 411 178 412 
<< pdiffusion >>
rect 178 411 179 412 
<< pdiffusion >>
rect 179 411 180 412 
<< m1 >>
rect 181 411 182 412 
<< pdiffusion >>
rect 192 411 193 412 
<< pdiffusion >>
rect 193 411 194 412 
<< pdiffusion >>
rect 194 411 195 412 
<< pdiffusion >>
rect 195 411 196 412 
<< pdiffusion >>
rect 196 411 197 412 
<< pdiffusion >>
rect 197 411 198 412 
<< m1 >>
rect 199 411 200 412 
<< m1 >>
rect 208 411 209 412 
<< pdiffusion >>
rect 210 411 211 412 
<< pdiffusion >>
rect 211 411 212 412 
<< pdiffusion >>
rect 212 411 213 412 
<< pdiffusion >>
rect 213 411 214 412 
<< pdiffusion >>
rect 214 411 215 412 
<< pdiffusion >>
rect 215 411 216 412 
<< m1 >>
rect 217 411 218 412 
<< pdiffusion >>
rect 228 411 229 412 
<< pdiffusion >>
rect 229 411 230 412 
<< pdiffusion >>
rect 230 411 231 412 
<< pdiffusion >>
rect 231 411 232 412 
<< pdiffusion >>
rect 232 411 233 412 
<< pdiffusion >>
rect 233 411 234 412 
<< m1 >>
rect 235 411 236 412 
<< pdiffusion >>
rect 246 411 247 412 
<< pdiffusion >>
rect 247 411 248 412 
<< pdiffusion >>
rect 248 411 249 412 
<< pdiffusion >>
rect 249 411 250 412 
<< pdiffusion >>
rect 250 411 251 412 
<< pdiffusion >>
rect 251 411 252 412 
<< m1 >>
rect 253 411 254 412 
<< pdiffusion >>
rect 264 411 265 412 
<< pdiffusion >>
rect 265 411 266 412 
<< pdiffusion >>
rect 266 411 267 412 
<< pdiffusion >>
rect 267 411 268 412 
<< pdiffusion >>
rect 268 411 269 412 
<< pdiffusion >>
rect 269 411 270 412 
<< m1 >>
rect 280 411 281 412 
<< pdiffusion >>
rect 282 411 283 412 
<< pdiffusion >>
rect 283 411 284 412 
<< pdiffusion >>
rect 284 411 285 412 
<< pdiffusion >>
rect 285 411 286 412 
<< pdiffusion >>
rect 286 411 287 412 
<< pdiffusion >>
rect 287 411 288 412 
<< pdiffusion >>
rect 300 411 301 412 
<< pdiffusion >>
rect 301 411 302 412 
<< pdiffusion >>
rect 302 411 303 412 
<< pdiffusion >>
rect 303 411 304 412 
<< pdiffusion >>
rect 304 411 305 412 
<< pdiffusion >>
rect 305 411 306 412 
<< m1 >>
rect 307 411 308 412 
<< m1 >>
rect 314 411 315 412 
<< m1 >>
rect 316 411 317 412 
<< pdiffusion >>
rect 318 411 319 412 
<< pdiffusion >>
rect 319 411 320 412 
<< pdiffusion >>
rect 320 411 321 412 
<< pdiffusion >>
rect 321 411 322 412 
<< pdiffusion >>
rect 322 411 323 412 
<< pdiffusion >>
rect 323 411 324 412 
<< m1 >>
rect 325 411 326 412 
<< m1 >>
rect 329 411 330 412 
<< pdiffusion >>
rect 336 411 337 412 
<< pdiffusion >>
rect 337 411 338 412 
<< pdiffusion >>
rect 338 411 339 412 
<< pdiffusion >>
rect 339 411 340 412 
<< pdiffusion >>
rect 340 411 341 412 
<< pdiffusion >>
rect 341 411 342 412 
<< m1 >>
rect 357 411 358 412 
<< m1 >>
rect 361 411 362 412 
<< m1 >>
rect 363 411 364 412 
<< m1 >>
rect 367 411 368 412 
<< pdiffusion >>
rect 372 411 373 412 
<< pdiffusion >>
rect 373 411 374 412 
<< pdiffusion >>
rect 374 411 375 412 
<< pdiffusion >>
rect 375 411 376 412 
<< pdiffusion >>
rect 376 411 377 412 
<< pdiffusion >>
rect 377 411 378 412 
<< m1 >>
rect 379 411 380 412 
<< m1 >>
rect 383 411 384 412 
<< m1 >>
rect 385 411 386 412 
<< pdiffusion >>
rect 390 411 391 412 
<< pdiffusion >>
rect 391 411 392 412 
<< pdiffusion >>
rect 392 411 393 412 
<< pdiffusion >>
rect 393 411 394 412 
<< pdiffusion >>
rect 394 411 395 412 
<< pdiffusion >>
rect 395 411 396 412 
<< m1 >>
rect 400 411 401 412 
<< m1 >>
rect 402 411 403 412 
<< m1 >>
rect 406 411 407 412 
<< pdiffusion >>
rect 408 411 409 412 
<< pdiffusion >>
rect 409 411 410 412 
<< pdiffusion >>
rect 410 411 411 412 
<< pdiffusion >>
rect 411 411 412 412 
<< pdiffusion >>
rect 412 411 413 412 
<< pdiffusion >>
rect 413 411 414 412 
<< m1 >>
rect 416 411 417 412 
<< m2 >>
rect 417 411 418 412 
<< m1 >>
rect 424 411 425 412 
<< pdiffusion >>
rect 426 411 427 412 
<< pdiffusion >>
rect 427 411 428 412 
<< pdiffusion >>
rect 428 411 429 412 
<< pdiffusion >>
rect 429 411 430 412 
<< pdiffusion >>
rect 430 411 431 412 
<< pdiffusion >>
rect 431 411 432 412 
<< m1 >>
rect 433 411 434 412 
<< m1 >>
rect 435 411 436 412 
<< pdiffusion >>
rect 444 411 445 412 
<< pdiffusion >>
rect 445 411 446 412 
<< pdiffusion >>
rect 446 411 447 412 
<< pdiffusion >>
rect 447 411 448 412 
<< pdiffusion >>
rect 448 411 449 412 
<< pdiffusion >>
rect 449 411 450 412 
<< pdiffusion >>
rect 462 411 463 412 
<< pdiffusion >>
rect 463 411 464 412 
<< pdiffusion >>
rect 464 411 465 412 
<< pdiffusion >>
rect 465 411 466 412 
<< pdiffusion >>
rect 466 411 467 412 
<< pdiffusion >>
rect 467 411 468 412 
<< m1 >>
rect 470 411 471 412 
<< m1 >>
rect 472 411 473 412 
<< m1 >>
rect 474 411 475 412 
<< m1 >>
rect 476 411 477 412 
<< pdiffusion >>
rect 480 411 481 412 
<< pdiffusion >>
rect 481 411 482 412 
<< pdiffusion >>
rect 482 411 483 412 
<< pdiffusion >>
rect 483 411 484 412 
<< pdiffusion >>
rect 484 411 485 412 
<< pdiffusion >>
rect 485 411 486 412 
<< m1 >>
rect 489 411 490 412 
<< m2 >>
rect 490 411 491 412 
<< pdiffusion >>
rect 498 411 499 412 
<< pdiffusion >>
rect 499 411 500 412 
<< pdiffusion >>
rect 500 411 501 412 
<< pdiffusion >>
rect 501 411 502 412 
<< pdiffusion >>
rect 502 411 503 412 
<< pdiffusion >>
rect 503 411 504 412 
<< pdiffusion >>
rect 516 411 517 412 
<< pdiffusion >>
rect 517 411 518 412 
<< pdiffusion >>
rect 518 411 519 412 
<< pdiffusion >>
rect 519 411 520 412 
<< pdiffusion >>
rect 520 411 521 412 
<< pdiffusion >>
rect 521 411 522 412 
<< pdiffusion >>
rect 12 412 13 413 
<< pdiffusion >>
rect 13 412 14 413 
<< pdiffusion >>
rect 14 412 15 413 
<< pdiffusion >>
rect 15 412 16 413 
<< pdiffusion >>
rect 16 412 17 413 
<< pdiffusion >>
rect 17 412 18 413 
<< m1 >>
rect 19 412 20 413 
<< m2 >>
rect 20 412 21 413 
<< m1 >>
rect 23 412 24 413 
<< m1 >>
rect 26 412 27 413 
<< pdiffusion >>
rect 30 412 31 413 
<< pdiffusion >>
rect 31 412 32 413 
<< pdiffusion >>
rect 32 412 33 413 
<< pdiffusion >>
rect 33 412 34 413 
<< pdiffusion >>
rect 34 412 35 413 
<< pdiffusion >>
rect 35 412 36 413 
<< m1 >>
rect 37 412 38 413 
<< m1 >>
rect 44 412 45 413 
<< pdiffusion >>
rect 48 412 49 413 
<< pdiffusion >>
rect 49 412 50 413 
<< pdiffusion >>
rect 50 412 51 413 
<< pdiffusion >>
rect 51 412 52 413 
<< pdiffusion >>
rect 52 412 53 413 
<< pdiffusion >>
rect 53 412 54 413 
<< m1 >>
rect 64 412 65 413 
<< pdiffusion >>
rect 66 412 67 413 
<< pdiffusion >>
rect 67 412 68 413 
<< pdiffusion >>
rect 68 412 69 413 
<< pdiffusion >>
rect 69 412 70 413 
<< pdiffusion >>
rect 70 412 71 413 
<< pdiffusion >>
rect 71 412 72 413 
<< m1 >>
rect 73 412 74 413 
<< m2 >>
rect 73 412 74 413 
<< m1 >>
rect 82 412 83 413 
<< pdiffusion >>
rect 84 412 85 413 
<< pdiffusion >>
rect 85 412 86 413 
<< pdiffusion >>
rect 86 412 87 413 
<< pdiffusion >>
rect 87 412 88 413 
<< pdiffusion >>
rect 88 412 89 413 
<< pdiffusion >>
rect 89 412 90 413 
<< m1 >>
rect 93 412 94 413 
<< m1 >>
rect 96 412 97 413 
<< pdiffusion >>
rect 102 412 103 413 
<< pdiffusion >>
rect 103 412 104 413 
<< pdiffusion >>
rect 104 412 105 413 
<< pdiffusion >>
rect 105 412 106 413 
<< pdiffusion >>
rect 106 412 107 413 
<< pdiffusion >>
rect 107 412 108 413 
<< m1 >>
rect 110 412 111 413 
<< m1 >>
rect 114 412 115 413 
<< pdiffusion >>
rect 120 412 121 413 
<< pdiffusion >>
rect 121 412 122 413 
<< pdiffusion >>
rect 122 412 123 413 
<< pdiffusion >>
rect 123 412 124 413 
<< pdiffusion >>
rect 124 412 125 413 
<< pdiffusion >>
rect 125 412 126 413 
<< m1 >>
rect 136 412 137 413 
<< pdiffusion >>
rect 138 412 139 413 
<< pdiffusion >>
rect 139 412 140 413 
<< pdiffusion >>
rect 140 412 141 413 
<< pdiffusion >>
rect 141 412 142 413 
<< pdiffusion >>
rect 142 412 143 413 
<< pdiffusion >>
rect 143 412 144 413 
<< m1 >>
rect 150 412 151 413 
<< m1 >>
rect 157 412 158 413 
<< m1 >>
rect 169 412 170 413 
<< pdiffusion >>
rect 174 412 175 413 
<< pdiffusion >>
rect 175 412 176 413 
<< pdiffusion >>
rect 176 412 177 413 
<< pdiffusion >>
rect 177 412 178 413 
<< pdiffusion >>
rect 178 412 179 413 
<< pdiffusion >>
rect 179 412 180 413 
<< m1 >>
rect 181 412 182 413 
<< pdiffusion >>
rect 192 412 193 413 
<< pdiffusion >>
rect 193 412 194 413 
<< pdiffusion >>
rect 194 412 195 413 
<< pdiffusion >>
rect 195 412 196 413 
<< pdiffusion >>
rect 196 412 197 413 
<< pdiffusion >>
rect 197 412 198 413 
<< m1 >>
rect 199 412 200 413 
<< m1 >>
rect 208 412 209 413 
<< pdiffusion >>
rect 210 412 211 413 
<< pdiffusion >>
rect 211 412 212 413 
<< pdiffusion >>
rect 212 412 213 413 
<< pdiffusion >>
rect 213 412 214 413 
<< pdiffusion >>
rect 214 412 215 413 
<< pdiffusion >>
rect 215 412 216 413 
<< m1 >>
rect 217 412 218 413 
<< pdiffusion >>
rect 228 412 229 413 
<< pdiffusion >>
rect 229 412 230 413 
<< pdiffusion >>
rect 230 412 231 413 
<< pdiffusion >>
rect 231 412 232 413 
<< pdiffusion >>
rect 232 412 233 413 
<< pdiffusion >>
rect 233 412 234 413 
<< m1 >>
rect 235 412 236 413 
<< pdiffusion >>
rect 246 412 247 413 
<< pdiffusion >>
rect 247 412 248 413 
<< pdiffusion >>
rect 248 412 249 413 
<< pdiffusion >>
rect 249 412 250 413 
<< pdiffusion >>
rect 250 412 251 413 
<< pdiffusion >>
rect 251 412 252 413 
<< m1 >>
rect 253 412 254 413 
<< pdiffusion >>
rect 264 412 265 413 
<< pdiffusion >>
rect 265 412 266 413 
<< pdiffusion >>
rect 266 412 267 413 
<< pdiffusion >>
rect 267 412 268 413 
<< pdiffusion >>
rect 268 412 269 413 
<< pdiffusion >>
rect 269 412 270 413 
<< m1 >>
rect 280 412 281 413 
<< pdiffusion >>
rect 282 412 283 413 
<< pdiffusion >>
rect 283 412 284 413 
<< pdiffusion >>
rect 284 412 285 413 
<< pdiffusion >>
rect 285 412 286 413 
<< pdiffusion >>
rect 286 412 287 413 
<< pdiffusion >>
rect 287 412 288 413 
<< pdiffusion >>
rect 300 412 301 413 
<< pdiffusion >>
rect 301 412 302 413 
<< pdiffusion >>
rect 302 412 303 413 
<< pdiffusion >>
rect 303 412 304 413 
<< pdiffusion >>
rect 304 412 305 413 
<< pdiffusion >>
rect 305 412 306 413 
<< m1 >>
rect 307 412 308 413 
<< m1 >>
rect 314 412 315 413 
<< m1 >>
rect 316 412 317 413 
<< pdiffusion >>
rect 318 412 319 413 
<< pdiffusion >>
rect 319 412 320 413 
<< pdiffusion >>
rect 320 412 321 413 
<< pdiffusion >>
rect 321 412 322 413 
<< pdiffusion >>
rect 322 412 323 413 
<< pdiffusion >>
rect 323 412 324 413 
<< m1 >>
rect 325 412 326 413 
<< m1 >>
rect 329 412 330 413 
<< pdiffusion >>
rect 336 412 337 413 
<< pdiffusion >>
rect 337 412 338 413 
<< pdiffusion >>
rect 338 412 339 413 
<< pdiffusion >>
rect 339 412 340 413 
<< pdiffusion >>
rect 340 412 341 413 
<< pdiffusion >>
rect 341 412 342 413 
<< m1 >>
rect 357 412 358 413 
<< m1 >>
rect 361 412 362 413 
<< m1 >>
rect 363 412 364 413 
<< m1 >>
rect 367 412 368 413 
<< pdiffusion >>
rect 372 412 373 413 
<< pdiffusion >>
rect 373 412 374 413 
<< pdiffusion >>
rect 374 412 375 413 
<< pdiffusion >>
rect 375 412 376 413 
<< pdiffusion >>
rect 376 412 377 413 
<< pdiffusion >>
rect 377 412 378 413 
<< m1 >>
rect 379 412 380 413 
<< m1 >>
rect 383 412 384 413 
<< m1 >>
rect 385 412 386 413 
<< pdiffusion >>
rect 390 412 391 413 
<< pdiffusion >>
rect 391 412 392 413 
<< pdiffusion >>
rect 392 412 393 413 
<< pdiffusion >>
rect 393 412 394 413 
<< pdiffusion >>
rect 394 412 395 413 
<< pdiffusion >>
rect 395 412 396 413 
<< m1 >>
rect 400 412 401 413 
<< m1 >>
rect 402 412 403 413 
<< m1 >>
rect 406 412 407 413 
<< pdiffusion >>
rect 408 412 409 413 
<< pdiffusion >>
rect 409 412 410 413 
<< pdiffusion >>
rect 410 412 411 413 
<< pdiffusion >>
rect 411 412 412 413 
<< pdiffusion >>
rect 412 412 413 413 
<< pdiffusion >>
rect 413 412 414 413 
<< m1 >>
rect 416 412 417 413 
<< m2 >>
rect 417 412 418 413 
<< m1 >>
rect 424 412 425 413 
<< pdiffusion >>
rect 426 412 427 413 
<< pdiffusion >>
rect 427 412 428 413 
<< pdiffusion >>
rect 428 412 429 413 
<< pdiffusion >>
rect 429 412 430 413 
<< pdiffusion >>
rect 430 412 431 413 
<< pdiffusion >>
rect 431 412 432 413 
<< m1 >>
rect 433 412 434 413 
<< m1 >>
rect 435 412 436 413 
<< pdiffusion >>
rect 444 412 445 413 
<< pdiffusion >>
rect 445 412 446 413 
<< pdiffusion >>
rect 446 412 447 413 
<< pdiffusion >>
rect 447 412 448 413 
<< pdiffusion >>
rect 448 412 449 413 
<< pdiffusion >>
rect 449 412 450 413 
<< pdiffusion >>
rect 462 412 463 413 
<< pdiffusion >>
rect 463 412 464 413 
<< pdiffusion >>
rect 464 412 465 413 
<< pdiffusion >>
rect 465 412 466 413 
<< pdiffusion >>
rect 466 412 467 413 
<< pdiffusion >>
rect 467 412 468 413 
<< m1 >>
rect 470 412 471 413 
<< m1 >>
rect 472 412 473 413 
<< m1 >>
rect 474 412 475 413 
<< m1 >>
rect 476 412 477 413 
<< pdiffusion >>
rect 480 412 481 413 
<< pdiffusion >>
rect 481 412 482 413 
<< pdiffusion >>
rect 482 412 483 413 
<< pdiffusion >>
rect 483 412 484 413 
<< pdiffusion >>
rect 484 412 485 413 
<< pdiffusion >>
rect 485 412 486 413 
<< m1 >>
rect 489 412 490 413 
<< m2 >>
rect 490 412 491 413 
<< pdiffusion >>
rect 498 412 499 413 
<< pdiffusion >>
rect 499 412 500 413 
<< pdiffusion >>
rect 500 412 501 413 
<< pdiffusion >>
rect 501 412 502 413 
<< pdiffusion >>
rect 502 412 503 413 
<< pdiffusion >>
rect 503 412 504 413 
<< pdiffusion >>
rect 516 412 517 413 
<< pdiffusion >>
rect 517 412 518 413 
<< pdiffusion >>
rect 518 412 519 413 
<< pdiffusion >>
rect 519 412 520 413 
<< pdiffusion >>
rect 520 412 521 413 
<< pdiffusion >>
rect 521 412 522 413 
<< pdiffusion >>
rect 12 413 13 414 
<< m1 >>
rect 13 413 14 414 
<< pdiffusion >>
rect 13 413 14 414 
<< pdiffusion >>
rect 14 413 15 414 
<< pdiffusion >>
rect 15 413 16 414 
<< pdiffusion >>
rect 16 413 17 414 
<< pdiffusion >>
rect 17 413 18 414 
<< m1 >>
rect 19 413 20 414 
<< m2 >>
rect 20 413 21 414 
<< m1 >>
rect 23 413 24 414 
<< m1 >>
rect 26 413 27 414 
<< pdiffusion >>
rect 30 413 31 414 
<< m1 >>
rect 31 413 32 414 
<< pdiffusion >>
rect 31 413 32 414 
<< pdiffusion >>
rect 32 413 33 414 
<< pdiffusion >>
rect 33 413 34 414 
<< pdiffusion >>
rect 34 413 35 414 
<< pdiffusion >>
rect 35 413 36 414 
<< m1 >>
rect 37 413 38 414 
<< m1 >>
rect 44 413 45 414 
<< pdiffusion >>
rect 48 413 49 414 
<< pdiffusion >>
rect 49 413 50 414 
<< pdiffusion >>
rect 50 413 51 414 
<< pdiffusion >>
rect 51 413 52 414 
<< pdiffusion >>
rect 52 413 53 414 
<< pdiffusion >>
rect 53 413 54 414 
<< m1 >>
rect 64 413 65 414 
<< pdiffusion >>
rect 66 413 67 414 
<< pdiffusion >>
rect 67 413 68 414 
<< pdiffusion >>
rect 68 413 69 414 
<< pdiffusion >>
rect 69 413 70 414 
<< pdiffusion >>
rect 70 413 71 414 
<< pdiffusion >>
rect 71 413 72 414 
<< m1 >>
rect 73 413 74 414 
<< m2 >>
rect 73 413 74 414 
<< m1 >>
rect 82 413 83 414 
<< pdiffusion >>
rect 84 413 85 414 
<< m1 >>
rect 85 413 86 414 
<< pdiffusion >>
rect 85 413 86 414 
<< pdiffusion >>
rect 86 413 87 414 
<< pdiffusion >>
rect 87 413 88 414 
<< pdiffusion >>
rect 88 413 89 414 
<< pdiffusion >>
rect 89 413 90 414 
<< m1 >>
rect 93 413 94 414 
<< m1 >>
rect 96 413 97 414 
<< pdiffusion >>
rect 102 413 103 414 
<< pdiffusion >>
rect 103 413 104 414 
<< pdiffusion >>
rect 104 413 105 414 
<< pdiffusion >>
rect 105 413 106 414 
<< m1 >>
rect 106 413 107 414 
<< pdiffusion >>
rect 106 413 107 414 
<< pdiffusion >>
rect 107 413 108 414 
<< m1 >>
rect 110 413 111 414 
<< m1 >>
rect 114 413 115 414 
<< pdiffusion >>
rect 120 413 121 414 
<< pdiffusion >>
rect 121 413 122 414 
<< pdiffusion >>
rect 122 413 123 414 
<< pdiffusion >>
rect 123 413 124 414 
<< m1 >>
rect 124 413 125 414 
<< pdiffusion >>
rect 124 413 125 414 
<< pdiffusion >>
rect 125 413 126 414 
<< m1 >>
rect 136 413 137 414 
<< pdiffusion >>
rect 138 413 139 414 
<< m1 >>
rect 139 413 140 414 
<< pdiffusion >>
rect 139 413 140 414 
<< pdiffusion >>
rect 140 413 141 414 
<< pdiffusion >>
rect 141 413 142 414 
<< pdiffusion >>
rect 142 413 143 414 
<< pdiffusion >>
rect 143 413 144 414 
<< m1 >>
rect 150 413 151 414 
<< m1 >>
rect 157 413 158 414 
<< m1 >>
rect 169 413 170 414 
<< pdiffusion >>
rect 174 413 175 414 
<< pdiffusion >>
rect 175 413 176 414 
<< pdiffusion >>
rect 176 413 177 414 
<< pdiffusion >>
rect 177 413 178 414 
<< pdiffusion >>
rect 178 413 179 414 
<< pdiffusion >>
rect 179 413 180 414 
<< m1 >>
rect 181 413 182 414 
<< pdiffusion >>
rect 192 413 193 414 
<< pdiffusion >>
rect 193 413 194 414 
<< pdiffusion >>
rect 194 413 195 414 
<< pdiffusion >>
rect 195 413 196 414 
<< pdiffusion >>
rect 196 413 197 414 
<< pdiffusion >>
rect 197 413 198 414 
<< m1 >>
rect 199 413 200 414 
<< m1 >>
rect 208 413 209 414 
<< pdiffusion >>
rect 210 413 211 414 
<< pdiffusion >>
rect 211 413 212 414 
<< pdiffusion >>
rect 212 413 213 414 
<< pdiffusion >>
rect 213 413 214 414 
<< pdiffusion >>
rect 214 413 215 414 
<< pdiffusion >>
rect 215 413 216 414 
<< m1 >>
rect 217 413 218 414 
<< pdiffusion >>
rect 228 413 229 414 
<< m1 >>
rect 229 413 230 414 
<< pdiffusion >>
rect 229 413 230 414 
<< pdiffusion >>
rect 230 413 231 414 
<< pdiffusion >>
rect 231 413 232 414 
<< pdiffusion >>
rect 232 413 233 414 
<< pdiffusion >>
rect 233 413 234 414 
<< m1 >>
rect 235 413 236 414 
<< pdiffusion >>
rect 246 413 247 414 
<< pdiffusion >>
rect 247 413 248 414 
<< pdiffusion >>
rect 248 413 249 414 
<< pdiffusion >>
rect 249 413 250 414 
<< pdiffusion >>
rect 250 413 251 414 
<< pdiffusion >>
rect 251 413 252 414 
<< m1 >>
rect 253 413 254 414 
<< pdiffusion >>
rect 264 413 265 414 
<< pdiffusion >>
rect 265 413 266 414 
<< pdiffusion >>
rect 266 413 267 414 
<< pdiffusion >>
rect 267 413 268 414 
<< m1 >>
rect 268 413 269 414 
<< pdiffusion >>
rect 268 413 269 414 
<< pdiffusion >>
rect 269 413 270 414 
<< m1 >>
rect 280 413 281 414 
<< pdiffusion >>
rect 282 413 283 414 
<< pdiffusion >>
rect 283 413 284 414 
<< pdiffusion >>
rect 284 413 285 414 
<< pdiffusion >>
rect 285 413 286 414 
<< pdiffusion >>
rect 286 413 287 414 
<< pdiffusion >>
rect 287 413 288 414 
<< pdiffusion >>
rect 300 413 301 414 
<< m1 >>
rect 301 413 302 414 
<< pdiffusion >>
rect 301 413 302 414 
<< pdiffusion >>
rect 302 413 303 414 
<< pdiffusion >>
rect 303 413 304 414 
<< pdiffusion >>
rect 304 413 305 414 
<< pdiffusion >>
rect 305 413 306 414 
<< m1 >>
rect 307 413 308 414 
<< m1 >>
rect 314 413 315 414 
<< m1 >>
rect 316 413 317 414 
<< pdiffusion >>
rect 318 413 319 414 
<< pdiffusion >>
rect 319 413 320 414 
<< pdiffusion >>
rect 320 413 321 414 
<< pdiffusion >>
rect 321 413 322 414 
<< m1 >>
rect 322 413 323 414 
<< pdiffusion >>
rect 322 413 323 414 
<< pdiffusion >>
rect 323 413 324 414 
<< m1 >>
rect 325 413 326 414 
<< m1 >>
rect 329 413 330 414 
<< pdiffusion >>
rect 336 413 337 414 
<< pdiffusion >>
rect 337 413 338 414 
<< pdiffusion >>
rect 338 413 339 414 
<< pdiffusion >>
rect 339 413 340 414 
<< pdiffusion >>
rect 340 413 341 414 
<< pdiffusion >>
rect 341 413 342 414 
<< m1 >>
rect 357 413 358 414 
<< m1 >>
rect 361 413 362 414 
<< m1 >>
rect 363 413 364 414 
<< m1 >>
rect 367 413 368 414 
<< pdiffusion >>
rect 372 413 373 414 
<< m1 >>
rect 373 413 374 414 
<< pdiffusion >>
rect 373 413 374 414 
<< pdiffusion >>
rect 374 413 375 414 
<< pdiffusion >>
rect 375 413 376 414 
<< m1 >>
rect 376 413 377 414 
<< pdiffusion >>
rect 376 413 377 414 
<< pdiffusion >>
rect 377 413 378 414 
<< m1 >>
rect 379 413 380 414 
<< m1 >>
rect 383 413 384 414 
<< m1 >>
rect 385 413 386 414 
<< pdiffusion >>
rect 390 413 391 414 
<< pdiffusion >>
rect 391 413 392 414 
<< pdiffusion >>
rect 392 413 393 414 
<< pdiffusion >>
rect 393 413 394 414 
<< m1 >>
rect 394 413 395 414 
<< pdiffusion >>
rect 394 413 395 414 
<< pdiffusion >>
rect 395 413 396 414 
<< m1 >>
rect 400 413 401 414 
<< m1 >>
rect 402 413 403 414 
<< m1 >>
rect 406 413 407 414 
<< pdiffusion >>
rect 408 413 409 414 
<< pdiffusion >>
rect 409 413 410 414 
<< pdiffusion >>
rect 410 413 411 414 
<< pdiffusion >>
rect 411 413 412 414 
<< pdiffusion >>
rect 412 413 413 414 
<< pdiffusion >>
rect 413 413 414 414 
<< m1 >>
rect 416 413 417 414 
<< m2 >>
rect 417 413 418 414 
<< m1 >>
rect 424 413 425 414 
<< pdiffusion >>
rect 426 413 427 414 
<< pdiffusion >>
rect 427 413 428 414 
<< pdiffusion >>
rect 428 413 429 414 
<< pdiffusion >>
rect 429 413 430 414 
<< pdiffusion >>
rect 430 413 431 414 
<< pdiffusion >>
rect 431 413 432 414 
<< m1 >>
rect 433 413 434 414 
<< m1 >>
rect 435 413 436 414 
<< pdiffusion >>
rect 444 413 445 414 
<< pdiffusion >>
rect 445 413 446 414 
<< pdiffusion >>
rect 446 413 447 414 
<< pdiffusion >>
rect 447 413 448 414 
<< pdiffusion >>
rect 448 413 449 414 
<< pdiffusion >>
rect 449 413 450 414 
<< pdiffusion >>
rect 462 413 463 414 
<< pdiffusion >>
rect 463 413 464 414 
<< pdiffusion >>
rect 464 413 465 414 
<< pdiffusion >>
rect 465 413 466 414 
<< pdiffusion >>
rect 466 413 467 414 
<< pdiffusion >>
rect 467 413 468 414 
<< m1 >>
rect 470 413 471 414 
<< m1 >>
rect 472 413 473 414 
<< m1 >>
rect 474 413 475 414 
<< m1 >>
rect 476 413 477 414 
<< pdiffusion >>
rect 480 413 481 414 
<< pdiffusion >>
rect 481 413 482 414 
<< pdiffusion >>
rect 482 413 483 414 
<< pdiffusion >>
rect 483 413 484 414 
<< pdiffusion >>
rect 484 413 485 414 
<< pdiffusion >>
rect 485 413 486 414 
<< m1 >>
rect 489 413 490 414 
<< m2 >>
rect 490 413 491 414 
<< pdiffusion >>
rect 498 413 499 414 
<< pdiffusion >>
rect 499 413 500 414 
<< pdiffusion >>
rect 500 413 501 414 
<< pdiffusion >>
rect 501 413 502 414 
<< pdiffusion >>
rect 502 413 503 414 
<< pdiffusion >>
rect 503 413 504 414 
<< pdiffusion >>
rect 516 413 517 414 
<< pdiffusion >>
rect 517 413 518 414 
<< pdiffusion >>
rect 518 413 519 414 
<< pdiffusion >>
rect 519 413 520 414 
<< pdiffusion >>
rect 520 413 521 414 
<< pdiffusion >>
rect 521 413 522 414 
<< m1 >>
rect 13 414 14 415 
<< m1 >>
rect 19 414 20 415 
<< m2 >>
rect 20 414 21 415 
<< m1 >>
rect 23 414 24 415 
<< m1 >>
rect 26 414 27 415 
<< m1 >>
rect 31 414 32 415 
<< m1 >>
rect 37 414 38 415 
<< m1 >>
rect 44 414 45 415 
<< m1 >>
rect 64 414 65 415 
<< m1 >>
rect 73 414 74 415 
<< m2 >>
rect 73 414 74 415 
<< m1 >>
rect 82 414 83 415 
<< m1 >>
rect 85 414 86 415 
<< m1 >>
rect 93 414 94 415 
<< m1 >>
rect 96 414 97 415 
<< m1 >>
rect 106 414 107 415 
<< m1 >>
rect 110 414 111 415 
<< m1 >>
rect 114 414 115 415 
<< m1 >>
rect 124 414 125 415 
<< m1 >>
rect 136 414 137 415 
<< m1 >>
rect 139 414 140 415 
<< m1 >>
rect 150 414 151 415 
<< m1 >>
rect 157 414 158 415 
<< m1 >>
rect 169 414 170 415 
<< m1 >>
rect 181 414 182 415 
<< m1 >>
rect 199 414 200 415 
<< m1 >>
rect 208 414 209 415 
<< m1 >>
rect 217 414 218 415 
<< m1 >>
rect 229 414 230 415 
<< m1 >>
rect 235 414 236 415 
<< m1 >>
rect 253 414 254 415 
<< m1 >>
rect 268 414 269 415 
<< m1 >>
rect 280 414 281 415 
<< m1 >>
rect 301 414 302 415 
<< m1 >>
rect 307 414 308 415 
<< m2 >>
rect 307 414 308 415 
<< m2c >>
rect 307 414 308 415 
<< m1 >>
rect 307 414 308 415 
<< m2 >>
rect 307 414 308 415 
<< m1 >>
rect 314 414 315 415 
<< m1 >>
rect 316 414 317 415 
<< m1 >>
rect 322 414 323 415 
<< m1 >>
rect 325 414 326 415 
<< m1 >>
rect 329 414 330 415 
<< m1 >>
rect 357 414 358 415 
<< m1 >>
rect 361 414 362 415 
<< m1 >>
rect 363 414 364 415 
<< m1 >>
rect 367 414 368 415 
<< m1 >>
rect 373 414 374 415 
<< m1 >>
rect 376 414 377 415 
<< m1 >>
rect 379 414 380 415 
<< m1 >>
rect 383 414 384 415 
<< m1 >>
rect 385 414 386 415 
<< m1 >>
rect 394 414 395 415 
<< m1 >>
rect 400 414 401 415 
<< m1 >>
rect 402 414 403 415 
<< m1 >>
rect 406 414 407 415 
<< m1 >>
rect 416 414 417 415 
<< m2 >>
rect 417 414 418 415 
<< m1 >>
rect 424 414 425 415 
<< m1 >>
rect 433 414 434 415 
<< m1 >>
rect 435 414 436 415 
<< m1 >>
rect 470 414 471 415 
<< m1 >>
rect 472 414 473 415 
<< m1 >>
rect 474 414 475 415 
<< m1 >>
rect 476 414 477 415 
<< m1 >>
rect 489 414 490 415 
<< m2 >>
rect 490 414 491 415 
<< m1 >>
rect 13 415 14 416 
<< m1 >>
rect 17 415 18 416 
<< m2 >>
rect 17 415 18 416 
<< m2c >>
rect 17 415 18 416 
<< m1 >>
rect 17 415 18 416 
<< m2 >>
rect 17 415 18 416 
<< m2 >>
rect 18 415 19 416 
<< m1 >>
rect 19 415 20 416 
<< m2 >>
rect 19 415 20 416 
<< m2 >>
rect 20 415 21 416 
<< m1 >>
rect 23 415 24 416 
<< m1 >>
rect 26 415 27 416 
<< m1 >>
rect 31 415 32 416 
<< m1 >>
rect 37 415 38 416 
<< m1 >>
rect 44 415 45 416 
<< m1 >>
rect 64 415 65 416 
<< m1 >>
rect 73 415 74 416 
<< m2 >>
rect 73 415 74 416 
<< m1 >>
rect 82 415 83 416 
<< m1 >>
rect 85 415 86 416 
<< m1 >>
rect 93 415 94 416 
<< m1 >>
rect 96 415 97 416 
<< m1 >>
rect 106 415 107 416 
<< m1 >>
rect 110 415 111 416 
<< m1 >>
rect 114 415 115 416 
<< m1 >>
rect 124 415 125 416 
<< m2 >>
rect 125 415 126 416 
<< m1 >>
rect 126 415 127 416 
<< m2 >>
rect 126 415 127 416 
<< m2c >>
rect 126 415 127 416 
<< m1 >>
rect 126 415 127 416 
<< m2 >>
rect 126 415 127 416 
<< m1 >>
rect 127 415 128 416 
<< m1 >>
rect 128 415 129 416 
<< m1 >>
rect 129 415 130 416 
<< m1 >>
rect 130 415 131 416 
<< m1 >>
rect 131 415 132 416 
<< m1 >>
rect 132 415 133 416 
<< m1 >>
rect 133 415 134 416 
<< m1 >>
rect 134 415 135 416 
<< m1 >>
rect 135 415 136 416 
<< m1 >>
rect 136 415 137 416 
<< m1 >>
rect 139 415 140 416 
<< m1 >>
rect 150 415 151 416 
<< m1 >>
rect 157 415 158 416 
<< m1 >>
rect 169 415 170 416 
<< m1 >>
rect 181 415 182 416 
<< m1 >>
rect 199 415 200 416 
<< m1 >>
rect 208 415 209 416 
<< m1 >>
rect 217 415 218 416 
<< m1 >>
rect 229 415 230 416 
<< m1 >>
rect 235 415 236 416 
<< m1 >>
rect 253 415 254 416 
<< m1 >>
rect 268 415 269 416 
<< m2 >>
rect 269 415 270 416 
<< m1 >>
rect 270 415 271 416 
<< m2 >>
rect 270 415 271 416 
<< m2c >>
rect 270 415 271 416 
<< m1 >>
rect 270 415 271 416 
<< m2 >>
rect 270 415 271 416 
<< m1 >>
rect 271 415 272 416 
<< m1 >>
rect 272 415 273 416 
<< m1 >>
rect 273 415 274 416 
<< m1 >>
rect 274 415 275 416 
<< m1 >>
rect 275 415 276 416 
<< m1 >>
rect 276 415 277 416 
<< m1 >>
rect 277 415 278 416 
<< m1 >>
rect 278 415 279 416 
<< m1 >>
rect 279 415 280 416 
<< m1 >>
rect 280 415 281 416 
<< m1 >>
rect 301 415 302 416 
<< m2 >>
rect 307 415 308 416 
<< m2 >>
rect 308 415 309 416 
<< m2 >>
rect 309 415 310 416 
<< m2 >>
rect 310 415 311 416 
<< m2 >>
rect 311 415 312 416 
<< m2 >>
rect 312 415 313 416 
<< m2 >>
rect 313 415 314 416 
<< m1 >>
rect 314 415 315 416 
<< m2 >>
rect 314 415 315 416 
<< m2 >>
rect 315 415 316 416 
<< m1 >>
rect 316 415 317 416 
<< m2 >>
rect 316 415 317 416 
<< m2 >>
rect 317 415 318 416 
<< m1 >>
rect 318 415 319 416 
<< m2 >>
rect 318 415 319 416 
<< m2c >>
rect 318 415 319 416 
<< m1 >>
rect 318 415 319 416 
<< m2 >>
rect 318 415 319 416 
<< m1 >>
rect 322 415 323 416 
<< m1 >>
rect 325 415 326 416 
<< m1 >>
rect 329 415 330 416 
<< m1 >>
rect 357 415 358 416 
<< m1 >>
rect 361 415 362 416 
<< m1 >>
rect 363 415 364 416 
<< m1 >>
rect 367 415 368 416 
<< m1 >>
rect 373 415 374 416 
<< m1 >>
rect 374 415 375 416 
<< m2 >>
rect 374 415 375 416 
<< m2c >>
rect 374 415 375 416 
<< m1 >>
rect 374 415 375 416 
<< m2 >>
rect 374 415 375 416 
<< m2 >>
rect 375 415 376 416 
<< m1 >>
rect 376 415 377 416 
<< m1 >>
rect 379 415 380 416 
<< m1 >>
rect 383 415 384 416 
<< m1 >>
rect 385 415 386 416 
<< m1 >>
rect 394 415 395 416 
<< m1 >>
rect 395 415 396 416 
<< m1 >>
rect 396 415 397 416 
<< m1 >>
rect 397 415 398 416 
<< m1 >>
rect 400 415 401 416 
<< m1 >>
rect 402 415 403 416 
<< m1 >>
rect 406 415 407 416 
<< m1 >>
rect 416 415 417 416 
<< m2 >>
rect 417 415 418 416 
<< m1 >>
rect 424 415 425 416 
<< m1 >>
rect 433 415 434 416 
<< m1 >>
rect 435 415 436 416 
<< m1 >>
rect 470 415 471 416 
<< m1 >>
rect 472 415 473 416 
<< m1 >>
rect 474 415 475 416 
<< m1 >>
rect 476 415 477 416 
<< m1 >>
rect 489 415 490 416 
<< m2 >>
rect 490 415 491 416 
<< m1 >>
rect 13 416 14 417 
<< m1 >>
rect 14 416 15 417 
<< m1 >>
rect 15 416 16 417 
<< m1 >>
rect 16 416 17 417 
<< m1 >>
rect 17 416 18 417 
<< m1 >>
rect 19 416 20 417 
<< m1 >>
rect 23 416 24 417 
<< m1 >>
rect 26 416 27 417 
<< m1 >>
rect 31 416 32 417 
<< m1 >>
rect 32 416 33 417 
<< m1 >>
rect 33 416 34 417 
<< m1 >>
rect 34 416 35 417 
<< m1 >>
rect 35 416 36 417 
<< m1 >>
rect 36 416 37 417 
<< m1 >>
rect 37 416 38 417 
<< m1 >>
rect 44 416 45 417 
<< m1 >>
rect 64 416 65 417 
<< m1 >>
rect 73 416 74 417 
<< m2 >>
rect 73 416 74 417 
<< m1 >>
rect 82 416 83 417 
<< m1 >>
rect 85 416 86 417 
<< m1 >>
rect 93 416 94 417 
<< m1 >>
rect 96 416 97 417 
<< m1 >>
rect 106 416 107 417 
<< m1 >>
rect 110 416 111 417 
<< m1 >>
rect 114 416 115 417 
<< m1 >>
rect 122 416 123 417 
<< m2 >>
rect 122 416 123 417 
<< m2c >>
rect 122 416 123 417 
<< m1 >>
rect 122 416 123 417 
<< m2 >>
rect 122 416 123 417 
<< m2 >>
rect 123 416 124 417 
<< m1 >>
rect 124 416 125 417 
<< m2 >>
rect 124 416 125 417 
<< m2 >>
rect 125 416 126 417 
<< m1 >>
rect 139 416 140 417 
<< m1 >>
rect 150 416 151 417 
<< m1 >>
rect 157 416 158 417 
<< m1 >>
rect 169 416 170 417 
<< m1 >>
rect 181 416 182 417 
<< m1 >>
rect 199 416 200 417 
<< m1 >>
rect 208 416 209 417 
<< m1 >>
rect 217 416 218 417 
<< m1 >>
rect 229 416 230 417 
<< m1 >>
rect 235 416 236 417 
<< m1 >>
rect 253 416 254 417 
<< m2 >>
rect 253 416 254 417 
<< m2c >>
rect 253 416 254 417 
<< m1 >>
rect 253 416 254 417 
<< m2 >>
rect 253 416 254 417 
<< m1 >>
rect 268 416 269 417 
<< m2 >>
rect 269 416 270 417 
<< m1 >>
rect 301 416 302 417 
<< m1 >>
rect 302 416 303 417 
<< m1 >>
rect 303 416 304 417 
<< m1 >>
rect 304 416 305 417 
<< m1 >>
rect 305 416 306 417 
<< m1 >>
rect 306 416 307 417 
<< m1 >>
rect 307 416 308 417 
<< m1 >>
rect 308 416 309 417 
<< m1 >>
rect 309 416 310 417 
<< m1 >>
rect 310 416 311 417 
<< m1 >>
rect 311 416 312 417 
<< m1 >>
rect 312 416 313 417 
<< m1 >>
rect 313 416 314 417 
<< m1 >>
rect 314 416 315 417 
<< m1 >>
rect 316 416 317 417 
<< m1 >>
rect 318 416 319 417 
<< m1 >>
rect 322 416 323 417 
<< m1 >>
rect 325 416 326 417 
<< m1 >>
rect 329 416 330 417 
<< m1 >>
rect 357 416 358 417 
<< m2 >>
rect 360 416 361 417 
<< m1 >>
rect 361 416 362 417 
<< m2 >>
rect 361 416 362 417 
<< m2 >>
rect 362 416 363 417 
<< m1 >>
rect 363 416 364 417 
<< m2 >>
rect 363 416 364 417 
<< m2 >>
rect 364 416 365 417 
<< m1 >>
rect 365 416 366 417 
<< m2 >>
rect 365 416 366 417 
<< m2c >>
rect 365 416 366 417 
<< m1 >>
rect 365 416 366 417 
<< m2 >>
rect 365 416 366 417 
<< m1 >>
rect 366 416 367 417 
<< m1 >>
rect 367 416 368 417 
<< m2 >>
rect 375 416 376 417 
<< m1 >>
rect 376 416 377 417 
<< m2 >>
rect 376 416 377 417 
<< m2 >>
rect 377 416 378 417 
<< m2 >>
rect 378 416 379 417 
<< m1 >>
rect 379 416 380 417 
<< m2 >>
rect 379 416 380 417 
<< m1 >>
rect 383 416 384 417 
<< m1 >>
rect 385 416 386 417 
<< m1 >>
rect 397 416 398 417 
<< m1 >>
rect 400 416 401 417 
<< m1 >>
rect 402 416 403 417 
<< m1 >>
rect 406 416 407 417 
<< m1 >>
rect 416 416 417 417 
<< m2 >>
rect 417 416 418 417 
<< m1 >>
rect 424 416 425 417 
<< m1 >>
rect 425 416 426 417 
<< m1 >>
rect 426 416 427 417 
<< m2 >>
rect 426 416 427 417 
<< m2c >>
rect 426 416 427 417 
<< m1 >>
rect 426 416 427 417 
<< m2 >>
rect 426 416 427 417 
<< m1 >>
rect 433 416 434 417 
<< m2 >>
rect 433 416 434 417 
<< m2c >>
rect 433 416 434 417 
<< m1 >>
rect 433 416 434 417 
<< m2 >>
rect 433 416 434 417 
<< m1 >>
rect 435 416 436 417 
<< m2 >>
rect 435 416 436 417 
<< m2c >>
rect 435 416 436 417 
<< m1 >>
rect 435 416 436 417 
<< m2 >>
rect 435 416 436 417 
<< m1 >>
rect 470 416 471 417 
<< m2 >>
rect 470 416 471 417 
<< m2c >>
rect 470 416 471 417 
<< m1 >>
rect 470 416 471 417 
<< m2 >>
rect 470 416 471 417 
<< m1 >>
rect 472 416 473 417 
<< m2 >>
rect 472 416 473 417 
<< m2c >>
rect 472 416 473 417 
<< m1 >>
rect 472 416 473 417 
<< m2 >>
rect 472 416 473 417 
<< m1 >>
rect 474 416 475 417 
<< m2 >>
rect 474 416 475 417 
<< m2c >>
rect 474 416 475 417 
<< m1 >>
rect 474 416 475 417 
<< m2 >>
rect 474 416 475 417 
<< m1 >>
rect 476 416 477 417 
<< m2 >>
rect 476 416 477 417 
<< m2c >>
rect 476 416 477 417 
<< m1 >>
rect 476 416 477 417 
<< m2 >>
rect 476 416 477 417 
<< m1 >>
rect 489 416 490 417 
<< m2 >>
rect 490 416 491 417 
<< m1 >>
rect 19 417 20 418 
<< m1 >>
rect 23 417 24 418 
<< m2 >>
rect 23 417 24 418 
<< m2c >>
rect 23 417 24 418 
<< m1 >>
rect 23 417 24 418 
<< m2 >>
rect 23 417 24 418 
<< m1 >>
rect 26 417 27 418 
<< m2 >>
rect 26 417 27 418 
<< m2c >>
rect 26 417 27 418 
<< m1 >>
rect 26 417 27 418 
<< m2 >>
rect 26 417 27 418 
<< m1 >>
rect 44 417 45 418 
<< m2 >>
rect 44 417 45 418 
<< m2c >>
rect 44 417 45 418 
<< m1 >>
rect 44 417 45 418 
<< m2 >>
rect 44 417 45 418 
<< m1 >>
rect 64 417 65 418 
<< m2 >>
rect 64 417 65 418 
<< m2c >>
rect 64 417 65 418 
<< m1 >>
rect 64 417 65 418 
<< m2 >>
rect 64 417 65 418 
<< m1 >>
rect 68 417 69 418 
<< m2 >>
rect 68 417 69 418 
<< m2c >>
rect 68 417 69 418 
<< m1 >>
rect 68 417 69 418 
<< m2 >>
rect 68 417 69 418 
<< m1 >>
rect 69 417 70 418 
<< m1 >>
rect 70 417 71 418 
<< m1 >>
rect 71 417 72 418 
<< m1 >>
rect 72 417 73 418 
<< m1 >>
rect 73 417 74 418 
<< m2 >>
rect 73 417 74 418 
<< m1 >>
rect 82 417 83 418 
<< m1 >>
rect 85 417 86 418 
<< m1 >>
rect 93 417 94 418 
<< m1 >>
rect 96 417 97 418 
<< m1 >>
rect 106 417 107 418 
<< m1 >>
rect 110 417 111 418 
<< m1 >>
rect 114 417 115 418 
<< m1 >>
rect 122 417 123 418 
<< m1 >>
rect 124 417 125 418 
<< m1 >>
rect 139 417 140 418 
<< m1 >>
rect 150 417 151 418 
<< m1 >>
rect 157 417 158 418 
<< m1 >>
rect 169 417 170 418 
<< m1 >>
rect 181 417 182 418 
<< m1 >>
rect 199 417 200 418 
<< m1 >>
rect 208 417 209 418 
<< m1 >>
rect 217 417 218 418 
<< m1 >>
rect 229 417 230 418 
<< m1 >>
rect 235 417 236 418 
<< m2 >>
rect 253 417 254 418 
<< m1 >>
rect 268 417 269 418 
<< m2 >>
rect 269 417 270 418 
<< m1 >>
rect 316 417 317 418 
<< m1 >>
rect 318 417 319 418 
<< m1 >>
rect 322 417 323 418 
<< m1 >>
rect 325 417 326 418 
<< m1 >>
rect 329 417 330 418 
<< m1 >>
rect 357 417 358 418 
<< m2 >>
rect 360 417 361 418 
<< m1 >>
rect 361 417 362 418 
<< m1 >>
rect 363 417 364 418 
<< m1 >>
rect 376 417 377 418 
<< m1 >>
rect 379 417 380 418 
<< m2 >>
rect 379 417 380 418 
<< m1 >>
rect 383 417 384 418 
<< m1 >>
rect 385 417 386 418 
<< m1 >>
rect 397 417 398 418 
<< m1 >>
rect 400 417 401 418 
<< m1 >>
rect 402 417 403 418 
<< m1 >>
rect 406 417 407 418 
<< m1 >>
rect 416 417 417 418 
<< m2 >>
rect 417 417 418 418 
<< m2 >>
rect 426 417 427 418 
<< m2 >>
rect 433 417 434 418 
<< m2 >>
rect 435 417 436 418 
<< m2 >>
rect 470 417 471 418 
<< m2 >>
rect 472 417 473 418 
<< m2 >>
rect 474 417 475 418 
<< m2 >>
rect 476 417 477 418 
<< m1 >>
rect 489 417 490 418 
<< m2 >>
rect 490 417 491 418 
<< m1 >>
rect 16 418 17 419 
<< m1 >>
rect 17 418 18 419 
<< m2 >>
rect 17 418 18 419 
<< m2c >>
rect 17 418 18 419 
<< m1 >>
rect 17 418 18 419 
<< m2 >>
rect 17 418 18 419 
<< m2 >>
rect 18 418 19 419 
<< m1 >>
rect 19 418 20 419 
<< m2 >>
rect 19 418 20 419 
<< m2 >>
rect 20 418 21 419 
<< m2 >>
rect 21 418 22 419 
<< m2 >>
rect 22 418 23 419 
<< m2 >>
rect 23 418 24 419 
<< m2 >>
rect 26 418 27 419 
<< m2 >>
rect 28 418 29 419 
<< m2 >>
rect 29 418 30 419 
<< m2 >>
rect 30 418 31 419 
<< m2 >>
rect 31 418 32 419 
<< m2 >>
rect 32 418 33 419 
<< m2 >>
rect 33 418 34 419 
<< m2 >>
rect 34 418 35 419 
<< m2 >>
rect 35 418 36 419 
<< m2 >>
rect 36 418 37 419 
<< m2 >>
rect 37 418 38 419 
<< m2 >>
rect 38 418 39 419 
<< m2 >>
rect 39 418 40 419 
<< m2 >>
rect 40 418 41 419 
<< m2 >>
rect 41 418 42 419 
<< m2 >>
rect 42 418 43 419 
<< m2 >>
rect 43 418 44 419 
<< m2 >>
rect 44 418 45 419 
<< m2 >>
rect 64 418 65 419 
<< m2 >>
rect 68 418 69 419 
<< m2 >>
rect 73 418 74 419 
<< m1 >>
rect 82 418 83 419 
<< m1 >>
rect 85 418 86 419 
<< m1 >>
rect 93 418 94 419 
<< m1 >>
rect 96 418 97 419 
<< m1 >>
rect 100 418 101 419 
<< m1 >>
rect 101 418 102 419 
<< m1 >>
rect 102 418 103 419 
<< m1 >>
rect 103 418 104 419 
<< m1 >>
rect 104 418 105 419 
<< m1 >>
rect 105 418 106 419 
<< m1 >>
rect 106 418 107 419 
<< m1 >>
rect 110 418 111 419 
<< m1 >>
rect 114 418 115 419 
<< m1 >>
rect 122 418 123 419 
<< m1 >>
rect 124 418 125 419 
<< m1 >>
rect 139 418 140 419 
<< m1 >>
rect 150 418 151 419 
<< m1 >>
rect 157 418 158 419 
<< m1 >>
rect 169 418 170 419 
<< m1 >>
rect 181 418 182 419 
<< m1 >>
rect 199 418 200 419 
<< m1 >>
rect 208 418 209 419 
<< m1 >>
rect 217 418 218 419 
<< m1 >>
rect 229 418 230 419 
<< m1 >>
rect 235 418 236 419 
<< m1 >>
rect 236 418 237 419 
<< m1 >>
rect 237 418 238 419 
<< m1 >>
rect 238 418 239 419 
<< m1 >>
rect 239 418 240 419 
<< m1 >>
rect 240 418 241 419 
<< m1 >>
rect 241 418 242 419 
<< m1 >>
rect 242 418 243 419 
<< m1 >>
rect 243 418 244 419 
<< m1 >>
rect 244 418 245 419 
<< m1 >>
rect 245 418 246 419 
<< m1 >>
rect 246 418 247 419 
<< m1 >>
rect 247 418 248 419 
<< m1 >>
rect 248 418 249 419 
<< m1 >>
rect 249 418 250 419 
<< m1 >>
rect 250 418 251 419 
<< m1 >>
rect 251 418 252 419 
<< m1 >>
rect 252 418 253 419 
<< m1 >>
rect 253 418 254 419 
<< m2 >>
rect 253 418 254 419 
<< m1 >>
rect 254 418 255 419 
<< m1 >>
rect 255 418 256 419 
<< m1 >>
rect 256 418 257 419 
<< m1 >>
rect 257 418 258 419 
<< m1 >>
rect 258 418 259 419 
<< m1 >>
rect 259 418 260 419 
<< m1 >>
rect 260 418 261 419 
<< m1 >>
rect 261 418 262 419 
<< m1 >>
rect 262 418 263 419 
<< m1 >>
rect 263 418 264 419 
<< m1 >>
rect 264 418 265 419 
<< m2 >>
rect 264 418 265 419 
<< m1 >>
rect 265 418 266 419 
<< m2 >>
rect 265 418 266 419 
<< m1 >>
rect 266 418 267 419 
<< m2 >>
rect 266 418 267 419 
<< m1 >>
rect 267 418 268 419 
<< m2 >>
rect 267 418 268 419 
<< m1 >>
rect 268 418 269 419 
<< m2 >>
rect 268 418 269 419 
<< m2 >>
rect 269 418 270 419 
<< m1 >>
rect 316 418 317 419 
<< m1 >>
rect 318 418 319 419 
<< m1 >>
rect 319 418 320 419 
<< m1 >>
rect 320 418 321 419 
<< m2 >>
rect 320 418 321 419 
<< m2c >>
rect 320 418 321 419 
<< m1 >>
rect 320 418 321 419 
<< m2 >>
rect 320 418 321 419 
<< m2 >>
rect 321 418 322 419 
<< m1 >>
rect 322 418 323 419 
<< m2 >>
rect 322 418 323 419 
<< m2 >>
rect 323 418 324 419 
<< m2 >>
rect 324 418 325 419 
<< m1 >>
rect 325 418 326 419 
<< m2 >>
rect 325 418 326 419 
<< m2 >>
rect 326 418 327 419 
<< m1 >>
rect 327 418 328 419 
<< m2 >>
rect 327 418 328 419 
<< m2c >>
rect 327 418 328 419 
<< m1 >>
rect 327 418 328 419 
<< m2 >>
rect 327 418 328 419 
<< m1 >>
rect 328 418 329 419 
<< m1 >>
rect 329 418 330 419 
<< m1 >>
rect 357 418 358 419 
<< m2 >>
rect 360 418 361 419 
<< m1 >>
rect 361 418 362 419 
<< m1 >>
rect 363 418 364 419 
<< m1 >>
rect 364 418 365 419 
<< m1 >>
rect 365 418 366 419 
<< m1 >>
rect 366 418 367 419 
<< m1 >>
rect 367 418 368 419 
<< m1 >>
rect 368 418 369 419 
<< m1 >>
rect 369 418 370 419 
<< m1 >>
rect 370 418 371 419 
<< m1 >>
rect 371 418 372 419 
<< m1 >>
rect 372 418 373 419 
<< m1 >>
rect 373 418 374 419 
<< m1 >>
rect 374 418 375 419 
<< m1 >>
rect 375 418 376 419 
<< m1 >>
rect 376 418 377 419 
<< m1 >>
rect 379 418 380 419 
<< m2 >>
rect 379 418 380 419 
<< m1 >>
rect 383 418 384 419 
<< m1 >>
rect 385 418 386 419 
<< m1 >>
rect 397 418 398 419 
<< m1 >>
rect 400 418 401 419 
<< m1 >>
rect 402 418 403 419 
<< m1 >>
rect 406 418 407 419 
<< m1 >>
rect 416 418 417 419 
<< m1 >>
rect 417 418 418 419 
<< m2 >>
rect 417 418 418 419 
<< m1 >>
rect 418 418 419 419 
<< m1 >>
rect 419 418 420 419 
<< m1 >>
rect 420 418 421 419 
<< m1 >>
rect 421 418 422 419 
<< m1 >>
rect 422 418 423 419 
<< m1 >>
rect 423 418 424 419 
<< m1 >>
rect 424 418 425 419 
<< m1 >>
rect 425 418 426 419 
<< m1 >>
rect 426 418 427 419 
<< m2 >>
rect 426 418 427 419 
<< m1 >>
rect 427 418 428 419 
<< m1 >>
rect 428 418 429 419 
<< m1 >>
rect 429 418 430 419 
<< m1 >>
rect 430 418 431 419 
<< m1 >>
rect 431 418 432 419 
<< m1 >>
rect 432 418 433 419 
<< m1 >>
rect 433 418 434 419 
<< m2 >>
rect 433 418 434 419 
<< m1 >>
rect 434 418 435 419 
<< m1 >>
rect 435 418 436 419 
<< m2 >>
rect 435 418 436 419 
<< m1 >>
rect 436 418 437 419 
<< m2 >>
rect 436 418 437 419 
<< m1 >>
rect 437 418 438 419 
<< m2 >>
rect 437 418 438 419 
<< m1 >>
rect 438 418 439 419 
<< m2 >>
rect 438 418 439 419 
<< m1 >>
rect 439 418 440 419 
<< m2 >>
rect 439 418 440 419 
<< m1 >>
rect 440 418 441 419 
<< m2 >>
rect 440 418 441 419 
<< m1 >>
rect 441 418 442 419 
<< m2 >>
rect 441 418 442 419 
<< m1 >>
rect 442 418 443 419 
<< m2 >>
rect 442 418 443 419 
<< m1 >>
rect 443 418 444 419 
<< m2 >>
rect 443 418 444 419 
<< m1 >>
rect 444 418 445 419 
<< m2 >>
rect 444 418 445 419 
<< m1 >>
rect 445 418 446 419 
<< m2 >>
rect 445 418 446 419 
<< m1 >>
rect 446 418 447 419 
<< m2 >>
rect 446 418 447 419 
<< m1 >>
rect 447 418 448 419 
<< m2 >>
rect 447 418 448 419 
<< m1 >>
rect 448 418 449 419 
<< m2 >>
rect 448 418 449 419 
<< m1 >>
rect 449 418 450 419 
<< m2 >>
rect 449 418 450 419 
<< m1 >>
rect 450 418 451 419 
<< m2 >>
rect 450 418 451 419 
<< m1 >>
rect 451 418 452 419 
<< m2 >>
rect 451 418 452 419 
<< m1 >>
rect 452 418 453 419 
<< m2 >>
rect 452 418 453 419 
<< m1 >>
rect 453 418 454 419 
<< m2 >>
rect 453 418 454 419 
<< m1 >>
rect 454 418 455 419 
<< m2 >>
rect 454 418 455 419 
<< m1 >>
rect 455 418 456 419 
<< m2 >>
rect 455 418 456 419 
<< m1 >>
rect 456 418 457 419 
<< m2 >>
rect 456 418 457 419 
<< m1 >>
rect 457 418 458 419 
<< m2 >>
rect 457 418 458 419 
<< m1 >>
rect 458 418 459 419 
<< m2 >>
rect 458 418 459 419 
<< m1 >>
rect 459 418 460 419 
<< m2 >>
rect 459 418 460 419 
<< m1 >>
rect 460 418 461 419 
<< m2 >>
rect 460 418 461 419 
<< m1 >>
rect 461 418 462 419 
<< m2 >>
rect 461 418 462 419 
<< m1 >>
rect 462 418 463 419 
<< m2 >>
rect 462 418 463 419 
<< m1 >>
rect 463 418 464 419 
<< m2 >>
rect 463 418 464 419 
<< m1 >>
rect 464 418 465 419 
<< m2 >>
rect 464 418 465 419 
<< m1 >>
rect 465 418 466 419 
<< m2 >>
rect 465 418 466 419 
<< m1 >>
rect 466 418 467 419 
<< m2 >>
rect 466 418 467 419 
<< m2 >>
rect 467 418 468 419 
<< m1 >>
rect 468 418 469 419 
<< m2 >>
rect 468 418 469 419 
<< m2c >>
rect 468 418 469 419 
<< m1 >>
rect 468 418 469 419 
<< m2 >>
rect 468 418 469 419 
<< m1 >>
rect 469 418 470 419 
<< m1 >>
rect 470 418 471 419 
<< m2 >>
rect 470 418 471 419 
<< m1 >>
rect 471 418 472 419 
<< m1 >>
rect 472 418 473 419 
<< m2 >>
rect 472 418 473 419 
<< m1 >>
rect 473 418 474 419 
<< m1 >>
rect 474 418 475 419 
<< m2 >>
rect 474 418 475 419 
<< m1 >>
rect 475 418 476 419 
<< m1 >>
rect 476 418 477 419 
<< m2 >>
rect 476 418 477 419 
<< m1 >>
rect 477 418 478 419 
<< m1 >>
rect 478 418 479 419 
<< m1 >>
rect 479 418 480 419 
<< m1 >>
rect 480 418 481 419 
<< m2 >>
rect 480 418 481 419 
<< m1 >>
rect 481 418 482 419 
<< m2 >>
rect 481 418 482 419 
<< m1 >>
rect 482 418 483 419 
<< m2 >>
rect 482 418 483 419 
<< m1 >>
rect 483 418 484 419 
<< m2 >>
rect 483 418 484 419 
<< m1 >>
rect 484 418 485 419 
<< m2 >>
rect 484 418 485 419 
<< m1 >>
rect 485 418 486 419 
<< m2 >>
rect 485 418 486 419 
<< m1 >>
rect 486 418 487 419 
<< m2 >>
rect 486 418 487 419 
<< m2 >>
rect 487 418 488 419 
<< m2 >>
rect 488 418 489 419 
<< m1 >>
rect 489 418 490 419 
<< m2 >>
rect 489 418 490 419 
<< m2 >>
rect 490 418 491 419 
<< m1 >>
rect 16 419 17 420 
<< m1 >>
rect 19 419 20 420 
<< m1 >>
rect 21 419 22 420 
<< m1 >>
rect 22 419 23 420 
<< m1 >>
rect 23 419 24 420 
<< m1 >>
rect 24 419 25 420 
<< m1 >>
rect 25 419 26 420 
<< m1 >>
rect 26 419 27 420 
<< m2 >>
rect 26 419 27 420 
<< m1 >>
rect 27 419 28 420 
<< m1 >>
rect 28 419 29 420 
<< m2 >>
rect 28 419 29 420 
<< m1 >>
rect 29 419 30 420 
<< m1 >>
rect 30 419 31 420 
<< m1 >>
rect 31 419 32 420 
<< m1 >>
rect 32 419 33 420 
<< m1 >>
rect 33 419 34 420 
<< m1 >>
rect 34 419 35 420 
<< m1 >>
rect 35 419 36 420 
<< m1 >>
rect 36 419 37 420 
<< m1 >>
rect 37 419 38 420 
<< m1 >>
rect 38 419 39 420 
<< m1 >>
rect 39 419 40 420 
<< m1 >>
rect 40 419 41 420 
<< m1 >>
rect 41 419 42 420 
<< m1 >>
rect 42 419 43 420 
<< m1 >>
rect 43 419 44 420 
<< m1 >>
rect 44 419 45 420 
<< m1 >>
rect 45 419 46 420 
<< m1 >>
rect 46 419 47 420 
<< m1 >>
rect 47 419 48 420 
<< m1 >>
rect 48 419 49 420 
<< m1 >>
rect 49 419 50 420 
<< m1 >>
rect 50 419 51 420 
<< m1 >>
rect 51 419 52 420 
<< m1 >>
rect 52 419 53 420 
<< m1 >>
rect 53 419 54 420 
<< m1 >>
rect 54 419 55 420 
<< m1 >>
rect 55 419 56 420 
<< m1 >>
rect 56 419 57 420 
<< m1 >>
rect 57 419 58 420 
<< m1 >>
rect 58 419 59 420 
<< m1 >>
rect 59 419 60 420 
<< m1 >>
rect 60 419 61 420 
<< m1 >>
rect 61 419 62 420 
<< m1 >>
rect 62 419 63 420 
<< m1 >>
rect 63 419 64 420 
<< m1 >>
rect 64 419 65 420 
<< m2 >>
rect 64 419 65 420 
<< m1 >>
rect 65 419 66 420 
<< m1 >>
rect 66 419 67 420 
<< m1 >>
rect 67 419 68 420 
<< m1 >>
rect 68 419 69 420 
<< m2 >>
rect 68 419 69 420 
<< m1 >>
rect 69 419 70 420 
<< m1 >>
rect 70 419 71 420 
<< m1 >>
rect 71 419 72 420 
<< m1 >>
rect 72 419 73 420 
<< m1 >>
rect 73 419 74 420 
<< m2 >>
rect 73 419 74 420 
<< m1 >>
rect 74 419 75 420 
<< m1 >>
rect 75 419 76 420 
<< m1 >>
rect 76 419 77 420 
<< m1 >>
rect 77 419 78 420 
<< m1 >>
rect 78 419 79 420 
<< m1 >>
rect 79 419 80 420 
<< m1 >>
rect 80 419 81 420 
<< m2 >>
rect 80 419 81 420 
<< m2c >>
rect 80 419 81 420 
<< m1 >>
rect 80 419 81 420 
<< m2 >>
rect 80 419 81 420 
<< m2 >>
rect 81 419 82 420 
<< m1 >>
rect 82 419 83 420 
<< m2 >>
rect 82 419 83 420 
<< m2 >>
rect 83 419 84 420 
<< m1 >>
rect 84 419 85 420 
<< m2 >>
rect 84 419 85 420 
<< m2c >>
rect 84 419 85 420 
<< m1 >>
rect 84 419 85 420 
<< m2 >>
rect 84 419 85 420 
<< m1 >>
rect 85 419 86 420 
<< m1 >>
rect 93 419 94 420 
<< m2 >>
rect 93 419 94 420 
<< m2c >>
rect 93 419 94 420 
<< m1 >>
rect 93 419 94 420 
<< m2 >>
rect 93 419 94 420 
<< m1 >>
rect 96 419 97 420 
<< m2 >>
rect 96 419 97 420 
<< m2c >>
rect 96 419 97 420 
<< m1 >>
rect 96 419 97 420 
<< m2 >>
rect 96 419 97 420 
<< m1 >>
rect 100 419 101 420 
<< m1 >>
rect 110 419 111 420 
<< m2 >>
rect 110 419 111 420 
<< m2c >>
rect 110 419 111 420 
<< m1 >>
rect 110 419 111 420 
<< m2 >>
rect 110 419 111 420 
<< m1 >>
rect 114 419 115 420 
<< m2 >>
rect 114 419 115 420 
<< m2c >>
rect 114 419 115 420 
<< m1 >>
rect 114 419 115 420 
<< m2 >>
rect 114 419 115 420 
<< m1 >>
rect 122 419 123 420 
<< m2 >>
rect 122 419 123 420 
<< m2c >>
rect 122 419 123 420 
<< m1 >>
rect 122 419 123 420 
<< m2 >>
rect 122 419 123 420 
<< m1 >>
rect 124 419 125 420 
<< m2 >>
rect 124 419 125 420 
<< m2c >>
rect 124 419 125 420 
<< m1 >>
rect 124 419 125 420 
<< m2 >>
rect 124 419 125 420 
<< m1 >>
rect 139 419 140 420 
<< m1 >>
rect 140 419 141 420 
<< m1 >>
rect 141 419 142 420 
<< m1 >>
rect 142 419 143 420 
<< m1 >>
rect 143 419 144 420 
<< m1 >>
rect 144 419 145 420 
<< m1 >>
rect 145 419 146 420 
<< m2 >>
rect 145 419 146 420 
<< m2c >>
rect 145 419 146 420 
<< m1 >>
rect 145 419 146 420 
<< m2 >>
rect 145 419 146 420 
<< m1 >>
rect 150 419 151 420 
<< m2 >>
rect 150 419 151 420 
<< m2c >>
rect 150 419 151 420 
<< m1 >>
rect 150 419 151 420 
<< m2 >>
rect 150 419 151 420 
<< m1 >>
rect 157 419 158 420 
<< m1 >>
rect 169 419 170 420 
<< m1 >>
rect 181 419 182 420 
<< m1 >>
rect 199 419 200 420 
<< m1 >>
rect 208 419 209 420 
<< m1 >>
rect 217 419 218 420 
<< m1 >>
rect 229 419 230 420 
<< m2 >>
rect 253 419 254 420 
<< m2 >>
rect 264 419 265 420 
<< m1 >>
rect 316 419 317 420 
<< m1 >>
rect 322 419 323 420 
<< m1 >>
rect 325 419 326 420 
<< m1 >>
rect 357 419 358 420 
<< m2 >>
rect 357 419 358 420 
<< m2c >>
rect 357 419 358 420 
<< m1 >>
rect 357 419 358 420 
<< m2 >>
rect 357 419 358 420 
<< m2 >>
rect 360 419 361 420 
<< m1 >>
rect 361 419 362 420 
<< m1 >>
rect 379 419 380 420 
<< m2 >>
rect 379 419 380 420 
<< m1 >>
rect 383 419 384 420 
<< m1 >>
rect 385 419 386 420 
<< m1 >>
rect 397 419 398 420 
<< m1 >>
rect 400 419 401 420 
<< m2 >>
rect 400 419 401 420 
<< m2c >>
rect 400 419 401 420 
<< m1 >>
rect 400 419 401 420 
<< m2 >>
rect 400 419 401 420 
<< m2 >>
rect 401 419 402 420 
<< m1 >>
rect 402 419 403 420 
<< m2 >>
rect 402 419 403 420 
<< m2 >>
rect 403 419 404 420 
<< m1 >>
rect 404 419 405 420 
<< m2 >>
rect 404 419 405 420 
<< m2c >>
rect 404 419 405 420 
<< m1 >>
rect 404 419 405 420 
<< m2 >>
rect 404 419 405 420 
<< m2 >>
rect 405 419 406 420 
<< m1 >>
rect 406 419 407 420 
<< m2 >>
rect 406 419 407 420 
<< m2 >>
rect 407 419 408 420 
<< m1 >>
rect 408 419 409 420 
<< m2 >>
rect 408 419 409 420 
<< m2c >>
rect 408 419 409 420 
<< m1 >>
rect 408 419 409 420 
<< m2 >>
rect 408 419 409 420 
<< m1 >>
rect 409 419 410 420 
<< m1 >>
rect 410 419 411 420 
<< m1 >>
rect 411 419 412 420 
<< m1 >>
rect 412 419 413 420 
<< m1 >>
rect 413 419 414 420 
<< m1 >>
rect 414 419 415 420 
<< m2 >>
rect 414 419 415 420 
<< m2c >>
rect 414 419 415 420 
<< m1 >>
rect 414 419 415 420 
<< m2 >>
rect 414 419 415 420 
<< m2 >>
rect 415 419 416 420 
<< m2 >>
rect 417 419 418 420 
<< m2 >>
rect 418 419 419 420 
<< m2 >>
rect 419 419 420 420 
<< m2 >>
rect 420 419 421 420 
<< m2 >>
rect 421 419 422 420 
<< m2 >>
rect 422 419 423 420 
<< m2 >>
rect 423 419 424 420 
<< m2 >>
rect 424 419 425 420 
<< m2 >>
rect 426 419 427 420 
<< m2 >>
rect 427 419 428 420 
<< m2 >>
rect 428 419 429 420 
<< m2 >>
rect 429 419 430 420 
<< m2 >>
rect 430 419 431 420 
<< m2 >>
rect 431 419 432 420 
<< m2 >>
rect 433 419 434 420 
<< m1 >>
rect 466 419 467 420 
<< m2 >>
rect 470 419 471 420 
<< m2 >>
rect 472 419 473 420 
<< m2 >>
rect 474 419 475 420 
<< m2 >>
rect 476 419 477 420 
<< m2 >>
rect 480 419 481 420 
<< m1 >>
rect 486 419 487 420 
<< m1 >>
rect 489 419 490 420 
<< m1 >>
rect 16 420 17 421 
<< m1 >>
rect 19 420 20 421 
<< m1 >>
rect 21 420 22 421 
<< m2 >>
rect 26 420 27 421 
<< m2 >>
rect 28 420 29 421 
<< m2 >>
rect 64 420 65 421 
<< m2 >>
rect 68 420 69 421 
<< m2 >>
rect 73 420 74 421 
<< m1 >>
rect 82 420 83 421 
<< m2 >>
rect 93 420 94 421 
<< m2 >>
rect 96 420 97 421 
<< m1 >>
rect 100 420 101 421 
<< m2 >>
rect 110 420 111 421 
<< m2 >>
rect 114 420 115 421 
<< m2 >>
rect 120 420 121 421 
<< m2 >>
rect 121 420 122 421 
<< m2 >>
rect 122 420 123 421 
<< m2 >>
rect 124 420 125 421 
<< m2 >>
rect 125 420 126 421 
<< m2 >>
rect 126 420 127 421 
<< m2 >>
rect 127 420 128 421 
<< m2 >>
rect 128 420 129 421 
<< m2 >>
rect 129 420 130 421 
<< m2 >>
rect 130 420 131 421 
<< m2 >>
rect 131 420 132 421 
<< m2 >>
rect 132 420 133 421 
<< m2 >>
rect 133 420 134 421 
<< m2 >>
rect 134 420 135 421 
<< m2 >>
rect 135 420 136 421 
<< m2 >>
rect 136 420 137 421 
<< m2 >>
rect 137 420 138 421 
<< m2 >>
rect 138 420 139 421 
<< m2 >>
rect 139 420 140 421 
<< m2 >>
rect 140 420 141 421 
<< m2 >>
rect 145 420 146 421 
<< m2 >>
rect 150 420 151 421 
<< m1 >>
rect 157 420 158 421 
<< m1 >>
rect 169 420 170 421 
<< m1 >>
rect 181 420 182 421 
<< m1 >>
rect 199 420 200 421 
<< m1 >>
rect 208 420 209 421 
<< m1 >>
rect 217 420 218 421 
<< m1 >>
rect 229 420 230 421 
<< m2 >>
rect 253 420 254 421 
<< m2 >>
rect 264 420 265 421 
<< m2 >>
rect 298 420 299 421 
<< m2 >>
rect 299 420 300 421 
<< m1 >>
rect 300 420 301 421 
<< m2 >>
rect 300 420 301 421 
<< m2c >>
rect 300 420 301 421 
<< m1 >>
rect 300 420 301 421 
<< m2 >>
rect 300 420 301 421 
<< m1 >>
rect 301 420 302 421 
<< m1 >>
rect 302 420 303 421 
<< m1 >>
rect 303 420 304 421 
<< m1 >>
rect 304 420 305 421 
<< m1 >>
rect 305 420 306 421 
<< m1 >>
rect 306 420 307 421 
<< m1 >>
rect 307 420 308 421 
<< m1 >>
rect 308 420 309 421 
<< m1 >>
rect 309 420 310 421 
<< m1 >>
rect 310 420 311 421 
<< m1 >>
rect 311 420 312 421 
<< m1 >>
rect 312 420 313 421 
<< m1 >>
rect 313 420 314 421 
<< m1 >>
rect 314 420 315 421 
<< m1 >>
rect 315 420 316 421 
<< m1 >>
rect 316 420 317 421 
<< m1 >>
rect 322 420 323 421 
<< m1 >>
rect 325 420 326 421 
<< m2 >>
rect 357 420 358 421 
<< m2 >>
rect 360 420 361 421 
<< m1 >>
rect 361 420 362 421 
<< m1 >>
rect 379 420 380 421 
<< m2 >>
rect 379 420 380 421 
<< m1 >>
rect 383 420 384 421 
<< m1 >>
rect 385 420 386 421 
<< m1 >>
rect 397 420 398 421 
<< m1 >>
rect 402 420 403 421 
<< m1 >>
rect 406 420 407 421 
<< m2 >>
rect 415 420 416 421 
<< m1 >>
rect 424 420 425 421 
<< m2 >>
rect 424 420 425 421 
<< m2c >>
rect 424 420 425 421 
<< m1 >>
rect 424 420 425 421 
<< m2 >>
rect 424 420 425 421 
<< m1 >>
rect 431 420 432 421 
<< m2 >>
rect 431 420 432 421 
<< m2c >>
rect 431 420 432 421 
<< m1 >>
rect 431 420 432 421 
<< m2 >>
rect 431 420 432 421 
<< m1 >>
rect 433 420 434 421 
<< m2 >>
rect 433 420 434 421 
<< m2c >>
rect 433 420 434 421 
<< m1 >>
rect 433 420 434 421 
<< m2 >>
rect 433 420 434 421 
<< m1 >>
rect 466 420 467 421 
<< m1 >>
rect 470 420 471 421 
<< m2 >>
rect 470 420 471 421 
<< m2c >>
rect 470 420 471 421 
<< m1 >>
rect 470 420 471 421 
<< m2 >>
rect 470 420 471 421 
<< m1 >>
rect 471 420 472 421 
<< m1 >>
rect 472 420 473 421 
<< m2 >>
rect 472 420 473 421 
<< m1 >>
rect 473 420 474 421 
<< m1 >>
rect 474 420 475 421 
<< m2 >>
rect 474 420 475 421 
<< m1 >>
rect 475 420 476 421 
<< m1 >>
rect 476 420 477 421 
<< m2 >>
rect 476 420 477 421 
<< m1 >>
rect 477 420 478 421 
<< m1 >>
rect 478 420 479 421 
<< m1 >>
rect 479 420 480 421 
<< m1 >>
rect 480 420 481 421 
<< m2 >>
rect 480 420 481 421 
<< m1 >>
rect 481 420 482 421 
<< m1 >>
rect 482 420 483 421 
<< m1 >>
rect 483 420 484 421 
<< m1 >>
rect 484 420 485 421 
<< m1 >>
rect 486 420 487 421 
<< m1 >>
rect 489 420 490 421 
<< m1 >>
rect 16 421 17 422 
<< m1 >>
rect 19 421 20 422 
<< m1 >>
rect 21 421 22 422 
<< m1 >>
rect 26 421 27 422 
<< m2 >>
rect 26 421 27 422 
<< m2c >>
rect 26 421 27 422 
<< m1 >>
rect 26 421 27 422 
<< m2 >>
rect 26 421 27 422 
<< m1 >>
rect 28 421 29 422 
<< m2 >>
rect 28 421 29 422 
<< m1 >>
rect 29 421 30 422 
<< m1 >>
rect 30 421 31 422 
<< m1 >>
rect 31 421 32 422 
<< m1 >>
rect 32 421 33 422 
<< m2 >>
rect 32 421 33 422 
<< m2c >>
rect 32 421 33 422 
<< m1 >>
rect 32 421 33 422 
<< m2 >>
rect 32 421 33 422 
<< m2 >>
rect 33 421 34 422 
<< m1 >>
rect 34 421 35 422 
<< m2 >>
rect 34 421 35 422 
<< m1 >>
rect 35 421 36 422 
<< m2 >>
rect 35 421 36 422 
<< m1 >>
rect 36 421 37 422 
<< m2 >>
rect 36 421 37 422 
<< m1 >>
rect 37 421 38 422 
<< m2 >>
rect 37 421 38 422 
<< m1 >>
rect 38 421 39 422 
<< m2 >>
rect 38 421 39 422 
<< m1 >>
rect 39 421 40 422 
<< m2 >>
rect 39 421 40 422 
<< m1 >>
rect 40 421 41 422 
<< m2 >>
rect 40 421 41 422 
<< m1 >>
rect 41 421 42 422 
<< m2 >>
rect 41 421 42 422 
<< m1 >>
rect 42 421 43 422 
<< m2 >>
rect 42 421 43 422 
<< m1 >>
rect 43 421 44 422 
<< m2 >>
rect 43 421 44 422 
<< m1 >>
rect 44 421 45 422 
<< m2 >>
rect 44 421 45 422 
<< m1 >>
rect 45 421 46 422 
<< m2 >>
rect 45 421 46 422 
<< m1 >>
rect 46 421 47 422 
<< m2 >>
rect 46 421 47 422 
<< m1 >>
rect 47 421 48 422 
<< m2 >>
rect 47 421 48 422 
<< m1 >>
rect 48 421 49 422 
<< m2 >>
rect 48 421 49 422 
<< m1 >>
rect 49 421 50 422 
<< m2 >>
rect 49 421 50 422 
<< m1 >>
rect 50 421 51 422 
<< m2 >>
rect 50 421 51 422 
<< m1 >>
rect 51 421 52 422 
<< m2 >>
rect 51 421 52 422 
<< m1 >>
rect 52 421 53 422 
<< m2 >>
rect 52 421 53 422 
<< m1 >>
rect 53 421 54 422 
<< m2 >>
rect 53 421 54 422 
<< m1 >>
rect 54 421 55 422 
<< m2 >>
rect 54 421 55 422 
<< m1 >>
rect 55 421 56 422 
<< m2 >>
rect 55 421 56 422 
<< m1 >>
rect 56 421 57 422 
<< m2 >>
rect 56 421 57 422 
<< m1 >>
rect 57 421 58 422 
<< m2 >>
rect 57 421 58 422 
<< m1 >>
rect 58 421 59 422 
<< m2 >>
rect 58 421 59 422 
<< m1 >>
rect 59 421 60 422 
<< m2 >>
rect 59 421 60 422 
<< m1 >>
rect 60 421 61 422 
<< m2 >>
rect 60 421 61 422 
<< m1 >>
rect 61 421 62 422 
<< m2 >>
rect 61 421 62 422 
<< m1 >>
rect 62 421 63 422 
<< m2 >>
rect 62 421 63 422 
<< m1 >>
rect 63 421 64 422 
<< m2 >>
rect 63 421 64 422 
<< m1 >>
rect 64 421 65 422 
<< m2 >>
rect 64 421 65 422 
<< m1 >>
rect 65 421 66 422 
<< m1 >>
rect 66 421 67 422 
<< m2 >>
rect 66 421 67 422 
<< m1 >>
rect 67 421 68 422 
<< m2 >>
rect 67 421 68 422 
<< m1 >>
rect 68 421 69 422 
<< m2 >>
rect 68 421 69 422 
<< m1 >>
rect 69 421 70 422 
<< m1 >>
rect 70 421 71 422 
<< m1 >>
rect 71 421 72 422 
<< m1 >>
rect 72 421 73 422 
<< m1 >>
rect 73 421 74 422 
<< m2 >>
rect 73 421 74 422 
<< m1 >>
rect 74 421 75 422 
<< m1 >>
rect 75 421 76 422 
<< m1 >>
rect 76 421 77 422 
<< m1 >>
rect 77 421 78 422 
<< m1 >>
rect 78 421 79 422 
<< m1 >>
rect 79 421 80 422 
<< m1 >>
rect 80 421 81 422 
<< m2 >>
rect 80 421 81 422 
<< m2c >>
rect 80 421 81 422 
<< m1 >>
rect 80 421 81 422 
<< m2 >>
rect 80 421 81 422 
<< m2 >>
rect 81 421 82 422 
<< m1 >>
rect 82 421 83 422 
<< m2 >>
rect 82 421 83 422 
<< m2 >>
rect 83 421 84 422 
<< m1 >>
rect 84 421 85 422 
<< m2 >>
rect 84 421 85 422 
<< m2c >>
rect 84 421 85 422 
<< m1 >>
rect 84 421 85 422 
<< m2 >>
rect 84 421 85 422 
<< m1 >>
rect 85 421 86 422 
<< m1 >>
rect 86 421 87 422 
<< m1 >>
rect 87 421 88 422 
<< m1 >>
rect 88 421 89 422 
<< m1 >>
rect 89 421 90 422 
<< m1 >>
rect 90 421 91 422 
<< m1 >>
rect 91 421 92 422 
<< m1 >>
rect 92 421 93 422 
<< m1 >>
rect 93 421 94 422 
<< m2 >>
rect 93 421 94 422 
<< m1 >>
rect 94 421 95 422 
<< m1 >>
rect 95 421 96 422 
<< m1 >>
rect 96 421 97 422 
<< m2 >>
rect 96 421 97 422 
<< m1 >>
rect 97 421 98 422 
<< m1 >>
rect 98 421 99 422 
<< m2 >>
rect 98 421 99 422 
<< m2c >>
rect 98 421 99 422 
<< m1 >>
rect 98 421 99 422 
<< m2 >>
rect 98 421 99 422 
<< m2 >>
rect 99 421 100 422 
<< m1 >>
rect 100 421 101 422 
<< m2 >>
rect 100 421 101 422 
<< m2 >>
rect 101 421 102 422 
<< m1 >>
rect 102 421 103 422 
<< m2 >>
rect 102 421 103 422 
<< m2c >>
rect 102 421 103 422 
<< m1 >>
rect 102 421 103 422 
<< m2 >>
rect 102 421 103 422 
<< m1 >>
rect 103 421 104 422 
<< m1 >>
rect 104 421 105 422 
<< m1 >>
rect 105 421 106 422 
<< m1 >>
rect 106 421 107 422 
<< m1 >>
rect 107 421 108 422 
<< m1 >>
rect 108 421 109 422 
<< m1 >>
rect 109 421 110 422 
<< m1 >>
rect 110 421 111 422 
<< m2 >>
rect 110 421 111 422 
<< m1 >>
rect 111 421 112 422 
<< m1 >>
rect 112 421 113 422 
<< m1 >>
rect 113 421 114 422 
<< m1 >>
rect 114 421 115 422 
<< m2 >>
rect 114 421 115 422 
<< m1 >>
rect 115 421 116 422 
<< m1 >>
rect 116 421 117 422 
<< m1 >>
rect 117 421 118 422 
<< m1 >>
rect 118 421 119 422 
<< m1 >>
rect 119 421 120 422 
<< m1 >>
rect 120 421 121 422 
<< m2 >>
rect 120 421 121 422 
<< m1 >>
rect 121 421 122 422 
<< m1 >>
rect 122 421 123 422 
<< m1 >>
rect 123 421 124 422 
<< m1 >>
rect 124 421 125 422 
<< m1 >>
rect 125 421 126 422 
<< m1 >>
rect 126 421 127 422 
<< m1 >>
rect 127 421 128 422 
<< m1 >>
rect 128 421 129 422 
<< m1 >>
rect 129 421 130 422 
<< m1 >>
rect 130 421 131 422 
<< m1 >>
rect 131 421 132 422 
<< m1 >>
rect 132 421 133 422 
<< m1 >>
rect 133 421 134 422 
<< m1 >>
rect 134 421 135 422 
<< m1 >>
rect 135 421 136 422 
<< m1 >>
rect 136 421 137 422 
<< m1 >>
rect 137 421 138 422 
<< m1 >>
rect 138 421 139 422 
<< m1 >>
rect 139 421 140 422 
<< m1 >>
rect 140 421 141 422 
<< m2 >>
rect 140 421 141 422 
<< m1 >>
rect 141 421 142 422 
<< m1 >>
rect 142 421 143 422 
<< m1 >>
rect 143 421 144 422 
<< m1 >>
rect 144 421 145 422 
<< m1 >>
rect 145 421 146 422 
<< m2 >>
rect 145 421 146 422 
<< m1 >>
rect 146 421 147 422 
<< m1 >>
rect 147 421 148 422 
<< m1 >>
rect 148 421 149 422 
<< m1 >>
rect 149 421 150 422 
<< m1 >>
rect 150 421 151 422 
<< m2 >>
rect 150 421 151 422 
<< m1 >>
rect 151 421 152 422 
<< m1 >>
rect 152 421 153 422 
<< m1 >>
rect 153 421 154 422 
<< m1 >>
rect 154 421 155 422 
<< m1 >>
rect 155 421 156 422 
<< m1 >>
rect 156 421 157 422 
<< m1 >>
rect 157 421 158 422 
<< m2 >>
rect 168 421 169 422 
<< m1 >>
rect 169 421 170 422 
<< m2 >>
rect 169 421 170 422 
<< m2 >>
rect 170 421 171 422 
<< m1 >>
rect 171 421 172 422 
<< m2 >>
rect 171 421 172 422 
<< m1 >>
rect 172 421 173 422 
<< m2 >>
rect 172 421 173 422 
<< m1 >>
rect 173 421 174 422 
<< m2 >>
rect 173 421 174 422 
<< m1 >>
rect 174 421 175 422 
<< m2 >>
rect 174 421 175 422 
<< m1 >>
rect 175 421 176 422 
<< m2 >>
rect 175 421 176 422 
<< m1 >>
rect 176 421 177 422 
<< m2 >>
rect 176 421 177 422 
<< m1 >>
rect 177 421 178 422 
<< m2 >>
rect 177 421 178 422 
<< m1 >>
rect 178 421 179 422 
<< m2 >>
rect 178 421 179 422 
<< m1 >>
rect 179 421 180 422 
<< m2 >>
rect 179 421 180 422 
<< m1 >>
rect 180 421 181 422 
<< m2 >>
rect 180 421 181 422 
<< m1 >>
rect 181 421 182 422 
<< m2 >>
rect 181 421 182 422 
<< m2 >>
rect 182 421 183 422 
<< m1 >>
rect 183 421 184 422 
<< m2 >>
rect 183 421 184 422 
<< m2c >>
rect 183 421 184 422 
<< m1 >>
rect 183 421 184 422 
<< m2 >>
rect 183 421 184 422 
<< m1 >>
rect 184 421 185 422 
<< m1 >>
rect 185 421 186 422 
<< m1 >>
rect 186 421 187 422 
<< m1 >>
rect 187 421 188 422 
<< m1 >>
rect 188 421 189 422 
<< m1 >>
rect 189 421 190 422 
<< m1 >>
rect 190 421 191 422 
<< m1 >>
rect 191 421 192 422 
<< m1 >>
rect 192 421 193 422 
<< m1 >>
rect 193 421 194 422 
<< m1 >>
rect 194 421 195 422 
<< m1 >>
rect 195 421 196 422 
<< m1 >>
rect 196 421 197 422 
<< m1 >>
rect 197 421 198 422 
<< m1 >>
rect 198 421 199 422 
<< m1 >>
rect 199 421 200 422 
<< m1 >>
rect 208 421 209 422 
<< m1 >>
rect 217 421 218 422 
<< m1 >>
rect 229 421 230 422 
<< m1 >>
rect 230 421 231 422 
<< m1 >>
rect 231 421 232 422 
<< m1 >>
rect 232 421 233 422 
<< m1 >>
rect 233 421 234 422 
<< m1 >>
rect 234 421 235 422 
<< m1 >>
rect 235 421 236 422 
<< m1 >>
rect 236 421 237 422 
<< m1 >>
rect 237 421 238 422 
<< m1 >>
rect 238 421 239 422 
<< m1 >>
rect 239 421 240 422 
<< m1 >>
rect 240 421 241 422 
<< m1 >>
rect 241 421 242 422 
<< m1 >>
rect 242 421 243 422 
<< m1 >>
rect 243 421 244 422 
<< m1 >>
rect 244 421 245 422 
<< m1 >>
rect 245 421 246 422 
<< m1 >>
rect 246 421 247 422 
<< m1 >>
rect 247 421 248 422 
<< m1 >>
rect 248 421 249 422 
<< m1 >>
rect 249 421 250 422 
<< m1 >>
rect 250 421 251 422 
<< m1 >>
rect 251 421 252 422 
<< m1 >>
rect 252 421 253 422 
<< m1 >>
rect 253 421 254 422 
<< m2 >>
rect 253 421 254 422 
<< m1 >>
rect 254 421 255 422 
<< m1 >>
rect 255 421 256 422 
<< m1 >>
rect 256 421 257 422 
<< m1 >>
rect 257 421 258 422 
<< m1 >>
rect 258 421 259 422 
<< m1 >>
rect 259 421 260 422 
<< m1 >>
rect 260 421 261 422 
<< m1 >>
rect 261 421 262 422 
<< m1 >>
rect 262 421 263 422 
<< m1 >>
rect 263 421 264 422 
<< m1 >>
rect 264 421 265 422 
<< m2 >>
rect 264 421 265 422 
<< m1 >>
rect 265 421 266 422 
<< m1 >>
rect 266 421 267 422 
<< m1 >>
rect 267 421 268 422 
<< m1 >>
rect 268 421 269 422 
<< m1 >>
rect 269 421 270 422 
<< m1 >>
rect 270 421 271 422 
<< m1 >>
rect 271 421 272 422 
<< m1 >>
rect 272 421 273 422 
<< m1 >>
rect 273 421 274 422 
<< m1 >>
rect 274 421 275 422 
<< m1 >>
rect 275 421 276 422 
<< m1 >>
rect 276 421 277 422 
<< m1 >>
rect 277 421 278 422 
<< m1 >>
rect 278 421 279 422 
<< m1 >>
rect 279 421 280 422 
<< m1 >>
rect 280 421 281 422 
<< m1 >>
rect 281 421 282 422 
<< m1 >>
rect 282 421 283 422 
<< m1 >>
rect 283 421 284 422 
<< m1 >>
rect 284 421 285 422 
<< m1 >>
rect 285 421 286 422 
<< m1 >>
rect 286 421 287 422 
<< m1 >>
rect 287 421 288 422 
<< m1 >>
rect 288 421 289 422 
<< m1 >>
rect 289 421 290 422 
<< m1 >>
rect 290 421 291 422 
<< m1 >>
rect 291 421 292 422 
<< m1 >>
rect 292 421 293 422 
<< m1 >>
rect 293 421 294 422 
<< m1 >>
rect 294 421 295 422 
<< m1 >>
rect 295 421 296 422 
<< m1 >>
rect 296 421 297 422 
<< m1 >>
rect 297 421 298 422 
<< m1 >>
rect 298 421 299 422 
<< m2 >>
rect 298 421 299 422 
<< m1 >>
rect 318 421 319 422 
<< m1 >>
rect 319 421 320 422 
<< m1 >>
rect 320 421 321 422 
<< m2 >>
rect 320 421 321 422 
<< m2c >>
rect 320 421 321 422 
<< m1 >>
rect 320 421 321 422 
<< m2 >>
rect 320 421 321 422 
<< m2 >>
rect 321 421 322 422 
<< m1 >>
rect 322 421 323 422 
<< m2 >>
rect 322 421 323 422 
<< m2 >>
rect 323 421 324 422 
<< m2 >>
rect 324 421 325 422 
<< m1 >>
rect 325 421 326 422 
<< m2 >>
rect 325 421 326 422 
<< m2 >>
rect 326 421 327 422 
<< m1 >>
rect 327 421 328 422 
<< m2 >>
rect 327 421 328 422 
<< m2c >>
rect 327 421 328 422 
<< m1 >>
rect 327 421 328 422 
<< m2 >>
rect 327 421 328 422 
<< m1 >>
rect 328 421 329 422 
<< m1 >>
rect 329 421 330 422 
<< m1 >>
rect 330 421 331 422 
<< m1 >>
rect 331 421 332 422 
<< m1 >>
rect 332 421 333 422 
<< m1 >>
rect 333 421 334 422 
<< m1 >>
rect 334 421 335 422 
<< m1 >>
rect 335 421 336 422 
<< m1 >>
rect 336 421 337 422 
<< m1 >>
rect 337 421 338 422 
<< m1 >>
rect 338 421 339 422 
<< m1 >>
rect 339 421 340 422 
<< m1 >>
rect 340 421 341 422 
<< m1 >>
rect 341 421 342 422 
<< m1 >>
rect 342 421 343 422 
<< m1 >>
rect 343 421 344 422 
<< m1 >>
rect 344 421 345 422 
<< m1 >>
rect 345 421 346 422 
<< m1 >>
rect 346 421 347 422 
<< m1 >>
rect 347 421 348 422 
<< m1 >>
rect 348 421 349 422 
<< m1 >>
rect 349 421 350 422 
<< m1 >>
rect 350 421 351 422 
<< m1 >>
rect 351 421 352 422 
<< m1 >>
rect 352 421 353 422 
<< m1 >>
rect 353 421 354 422 
<< m1 >>
rect 354 421 355 422 
<< m1 >>
rect 355 421 356 422 
<< m1 >>
rect 356 421 357 422 
<< m1 >>
rect 357 421 358 422 
<< m2 >>
rect 357 421 358 422 
<< m1 >>
rect 358 421 359 422 
<< m1 >>
rect 359 421 360 422 
<< m2 >>
rect 359 421 360 422 
<< m2c >>
rect 359 421 360 422 
<< m1 >>
rect 359 421 360 422 
<< m2 >>
rect 359 421 360 422 
<< m2 >>
rect 360 421 361 422 
<< m1 >>
rect 361 421 362 422 
<< m1 >>
rect 379 421 380 422 
<< m2 >>
rect 379 421 380 422 
<< m1 >>
rect 383 421 384 422 
<< m2 >>
rect 383 421 384 422 
<< m2c >>
rect 383 421 384 422 
<< m1 >>
rect 383 421 384 422 
<< m2 >>
rect 383 421 384 422 
<< m2 >>
rect 384 421 385 422 
<< m1 >>
rect 385 421 386 422 
<< m2 >>
rect 385 421 386 422 
<< m2 >>
rect 386 421 387 422 
<< m1 >>
rect 387 421 388 422 
<< m2 >>
rect 387 421 388 422 
<< m2c >>
rect 387 421 388 422 
<< m1 >>
rect 387 421 388 422 
<< m2 >>
rect 387 421 388 422 
<< m1 >>
rect 388 421 389 422 
<< m1 >>
rect 389 421 390 422 
<< m2 >>
rect 389 421 390 422 
<< m2c >>
rect 389 421 390 422 
<< m1 >>
rect 389 421 390 422 
<< m2 >>
rect 389 421 390 422 
<< m2 >>
rect 390 421 391 422 
<< m1 >>
rect 391 421 392 422 
<< m2 >>
rect 391 421 392 422 
<< m1 >>
rect 392 421 393 422 
<< m2 >>
rect 392 421 393 422 
<< m1 >>
rect 393 421 394 422 
<< m2 >>
rect 393 421 394 422 
<< m1 >>
rect 394 421 395 422 
<< m1 >>
rect 395 421 396 422 
<< m2 >>
rect 395 421 396 422 
<< m2c >>
rect 395 421 396 422 
<< m1 >>
rect 395 421 396 422 
<< m2 >>
rect 395 421 396 422 
<< m2 >>
rect 396 421 397 422 
<< m1 >>
rect 397 421 398 422 
<< m2 >>
rect 397 421 398 422 
<< m2 >>
rect 398 421 399 422 
<< m1 >>
rect 399 421 400 422 
<< m2 >>
rect 399 421 400 422 
<< m1 >>
rect 400 421 401 422 
<< m2 >>
rect 400 421 401 422 
<< m2c >>
rect 400 421 401 422 
<< m1 >>
rect 400 421 401 422 
<< m2 >>
rect 400 421 401 422 
<< m2 >>
rect 401 421 402 422 
<< m1 >>
rect 402 421 403 422 
<< m2 >>
rect 402 421 403 422 
<< m2 >>
rect 403 421 404 422 
<< m1 >>
rect 404 421 405 422 
<< m2 >>
rect 404 421 405 422 
<< m2c >>
rect 404 421 405 422 
<< m1 >>
rect 404 421 405 422 
<< m2 >>
rect 404 421 405 422 
<< m2 >>
rect 405 421 406 422 
<< m1 >>
rect 406 421 407 422 
<< m2 >>
rect 406 421 407 422 
<< m2 >>
rect 407 421 408 422 
<< m1 >>
rect 408 421 409 422 
<< m2 >>
rect 408 421 409 422 
<< m2c >>
rect 408 421 409 422 
<< m1 >>
rect 408 421 409 422 
<< m2 >>
rect 408 421 409 422 
<< m1 >>
rect 409 421 410 422 
<< m1 >>
rect 410 421 411 422 
<< m1 >>
rect 411 421 412 422 
<< m1 >>
rect 412 421 413 422 
<< m1 >>
rect 413 421 414 422 
<< m1 >>
rect 414 421 415 422 
<< m1 >>
rect 415 421 416 422 
<< m2 >>
rect 415 421 416 422 
<< m1 >>
rect 416 421 417 422 
<< m1 >>
rect 417 421 418 422 
<< m1 >>
rect 418 421 419 422 
<< m1 >>
rect 419 421 420 422 
<< m1 >>
rect 420 421 421 422 
<< m1 >>
rect 421 421 422 422 
<< m1 >>
rect 422 421 423 422 
<< m1 >>
rect 424 421 425 422 
<< m1 >>
rect 426 421 427 422 
<< m1 >>
rect 427 421 428 422 
<< m1 >>
rect 428 421 429 422 
<< m1 >>
rect 429 421 430 422 
<< m1 >>
rect 431 421 432 422 
<< m1 >>
rect 433 421 434 422 
<< m1 >>
rect 466 421 467 422 
<< m2 >>
rect 472 421 473 422 
<< m2 >>
rect 474 421 475 422 
<< m2 >>
rect 476 421 477 422 
<< m2 >>
rect 480 421 481 422 
<< m1 >>
rect 484 421 485 422 
<< m1 >>
rect 486 421 487 422 
<< m1 >>
rect 489 421 490 422 
<< m1 >>
rect 16 422 17 423 
<< m1 >>
rect 19 422 20 423 
<< m1 >>
rect 21 422 22 423 
<< m1 >>
rect 26 422 27 423 
<< m1 >>
rect 28 422 29 423 
<< m2 >>
rect 28 422 29 423 
<< m1 >>
rect 34 422 35 423 
<< m2 >>
rect 66 422 67 423 
<< m2 >>
rect 73 422 74 423 
<< m1 >>
rect 82 422 83 423 
<< m2 >>
rect 93 422 94 423 
<< m2 >>
rect 96 422 97 423 
<< m1 >>
rect 100 422 101 423 
<< m2 >>
rect 110 422 111 423 
<< m2 >>
rect 114 422 115 423 
<< m2 >>
rect 120 422 121 423 
<< m2 >>
rect 140 422 141 423 
<< m2 >>
rect 145 422 146 423 
<< m2 >>
rect 150 422 151 423 
<< m2 >>
rect 168 422 169 423 
<< m1 >>
rect 169 422 170 423 
<< m1 >>
rect 171 422 172 423 
<< m1 >>
rect 208 422 209 423 
<< m1 >>
rect 217 422 218 423 
<< m2 >>
rect 253 422 254 423 
<< m2 >>
rect 264 422 265 423 
<< m1 >>
rect 298 422 299 423 
<< m2 >>
rect 298 422 299 423 
<< m1 >>
rect 318 422 319 423 
<< m1 >>
rect 322 422 323 423 
<< m1 >>
rect 325 422 326 423 
<< m2 >>
rect 357 422 358 423 
<< m1 >>
rect 361 422 362 423 
<< m1 >>
rect 379 422 380 423 
<< m2 >>
rect 379 422 380 423 
<< m1 >>
rect 385 422 386 423 
<< m1 >>
rect 391 422 392 423 
<< m2 >>
rect 393 422 394 423 
<< m1 >>
rect 397 422 398 423 
<< m1 >>
rect 402 422 403 423 
<< m1 >>
rect 406 422 407 423 
<< m2 >>
rect 415 422 416 423 
<< m2 >>
rect 416 422 417 423 
<< m2 >>
rect 417 422 418 423 
<< m2 >>
rect 418 422 419 423 
<< m2 >>
rect 419 422 420 423 
<< m2 >>
rect 420 422 421 423 
<< m1 >>
rect 422 422 423 423 
<< m2 >>
rect 422 422 423 423 
<< m2c >>
rect 422 422 423 423 
<< m1 >>
rect 422 422 423 423 
<< m2 >>
rect 422 422 423 423 
<< m2 >>
rect 423 422 424 423 
<< m1 >>
rect 424 422 425 423 
<< m2 >>
rect 424 422 425 423 
<< m2 >>
rect 425 422 426 423 
<< m1 >>
rect 426 422 427 423 
<< m2 >>
rect 426 422 427 423 
<< m2c >>
rect 426 422 427 423 
<< m1 >>
rect 426 422 427 423 
<< m2 >>
rect 426 422 427 423 
<< m1 >>
rect 429 422 430 423 
<< m2 >>
rect 429 422 430 423 
<< m2c >>
rect 429 422 430 423 
<< m1 >>
rect 429 422 430 423 
<< m2 >>
rect 429 422 430 423 
<< m2 >>
rect 430 422 431 423 
<< m1 >>
rect 431 422 432 423 
<< m2 >>
rect 431 422 432 423 
<< m2 >>
rect 432 422 433 423 
<< m1 >>
rect 433 422 434 423 
<< m2 >>
rect 433 422 434 423 
<< m2 >>
rect 434 422 435 423 
<< m1 >>
rect 435 422 436 423 
<< m2 >>
rect 435 422 436 423 
<< m2c >>
rect 435 422 436 423 
<< m1 >>
rect 435 422 436 423 
<< m2 >>
rect 435 422 436 423 
<< m1 >>
rect 436 422 437 423 
<< m1 >>
rect 437 422 438 423 
<< m1 >>
rect 438 422 439 423 
<< m1 >>
rect 439 422 440 423 
<< m1 >>
rect 440 422 441 423 
<< m1 >>
rect 441 422 442 423 
<< m1 >>
rect 442 422 443 423 
<< m1 >>
rect 466 422 467 423 
<< m1 >>
rect 472 422 473 423 
<< m2 >>
rect 472 422 473 423 
<< m2c >>
rect 472 422 473 423 
<< m1 >>
rect 472 422 473 423 
<< m2 >>
rect 472 422 473 423 
<< m1 >>
rect 474 422 475 423 
<< m2 >>
rect 474 422 475 423 
<< m2c >>
rect 474 422 475 423 
<< m1 >>
rect 474 422 475 423 
<< m2 >>
rect 474 422 475 423 
<< m1 >>
rect 476 422 477 423 
<< m2 >>
rect 476 422 477 423 
<< m2c >>
rect 476 422 477 423 
<< m1 >>
rect 476 422 477 423 
<< m2 >>
rect 476 422 477 423 
<< m1 >>
rect 477 422 478 423 
<< m1 >>
rect 478 422 479 423 
<< m2 >>
rect 478 422 479 423 
<< m2c >>
rect 478 422 479 423 
<< m1 >>
rect 478 422 479 423 
<< m2 >>
rect 478 422 479 423 
<< m1 >>
rect 480 422 481 423 
<< m2 >>
rect 480 422 481 423 
<< m2c >>
rect 480 422 481 423 
<< m1 >>
rect 480 422 481 423 
<< m2 >>
rect 480 422 481 423 
<< m1 >>
rect 484 422 485 423 
<< m1 >>
rect 486 422 487 423 
<< m2 >>
rect 486 422 487 423 
<< m2c >>
rect 486 422 487 423 
<< m1 >>
rect 486 422 487 423 
<< m2 >>
rect 486 422 487 423 
<< m1 >>
rect 489 422 490 423 
<< m2 >>
rect 489 422 490 423 
<< m2c >>
rect 489 422 490 423 
<< m1 >>
rect 489 422 490 423 
<< m2 >>
rect 489 422 490 423 
<< m1 >>
rect 16 423 17 424 
<< m1 >>
rect 19 423 20 424 
<< m1 >>
rect 21 423 22 424 
<< m1 >>
rect 26 423 27 424 
<< m1 >>
rect 28 423 29 424 
<< m2 >>
rect 28 423 29 424 
<< m1 >>
rect 34 423 35 424 
<< m1 >>
rect 66 423 67 424 
<< m2 >>
rect 66 423 67 424 
<< m2c >>
rect 66 423 67 424 
<< m1 >>
rect 66 423 67 424 
<< m2 >>
rect 66 423 67 424 
<< m1 >>
rect 73 423 74 424 
<< m2 >>
rect 73 423 74 424 
<< m2c >>
rect 73 423 74 424 
<< m1 >>
rect 73 423 74 424 
<< m2 >>
rect 73 423 74 424 
<< m1 >>
rect 82 423 83 424 
<< m1 >>
rect 93 423 94 424 
<< m2 >>
rect 93 423 94 424 
<< m2c >>
rect 93 423 94 424 
<< m1 >>
rect 93 423 94 424 
<< m2 >>
rect 93 423 94 424 
<< m1 >>
rect 96 423 97 424 
<< m2 >>
rect 96 423 97 424 
<< m2c >>
rect 96 423 97 424 
<< m1 >>
rect 96 423 97 424 
<< m2 >>
rect 96 423 97 424 
<< m1 >>
rect 100 423 101 424 
<< m1 >>
rect 110 423 111 424 
<< m2 >>
rect 110 423 111 424 
<< m2c >>
rect 110 423 111 424 
<< m1 >>
rect 110 423 111 424 
<< m2 >>
rect 110 423 111 424 
<< m1 >>
rect 114 423 115 424 
<< m2 >>
rect 114 423 115 424 
<< m2c >>
rect 114 423 115 424 
<< m1 >>
rect 114 423 115 424 
<< m2 >>
rect 114 423 115 424 
<< m1 >>
rect 118 423 119 424 
<< m1 >>
rect 119 423 120 424 
<< m1 >>
rect 120 423 121 424 
<< m2 >>
rect 120 423 121 424 
<< m2c >>
rect 120 423 121 424 
<< m1 >>
rect 120 423 121 424 
<< m2 >>
rect 120 423 121 424 
<< m1 >>
rect 140 423 141 424 
<< m2 >>
rect 140 423 141 424 
<< m2c >>
rect 140 423 141 424 
<< m1 >>
rect 140 423 141 424 
<< m2 >>
rect 140 423 141 424 
<< m1 >>
rect 141 423 142 424 
<< m1 >>
rect 142 423 143 424 
<< m1 >>
rect 143 423 144 424 
<< m1 >>
rect 144 423 145 424 
<< m1 >>
rect 145 423 146 424 
<< m2 >>
rect 145 423 146 424 
<< m1 >>
rect 150 423 151 424 
<< m2 >>
rect 150 423 151 424 
<< m2c >>
rect 150 423 151 424 
<< m1 >>
rect 150 423 151 424 
<< m2 >>
rect 150 423 151 424 
<< m2 >>
rect 168 423 169 424 
<< m1 >>
rect 169 423 170 424 
<< m1 >>
rect 171 423 172 424 
<< m1 >>
rect 208 423 209 424 
<< m1 >>
rect 217 423 218 424 
<< m1 >>
rect 253 423 254 424 
<< m2 >>
rect 253 423 254 424 
<< m2c >>
rect 253 423 254 424 
<< m1 >>
rect 253 423 254 424 
<< m2 >>
rect 253 423 254 424 
<< m1 >>
rect 262 423 263 424 
<< m1 >>
rect 263 423 264 424 
<< m1 >>
rect 264 423 265 424 
<< m2 >>
rect 264 423 265 424 
<< m2c >>
rect 264 423 265 424 
<< m1 >>
rect 264 423 265 424 
<< m2 >>
rect 264 423 265 424 
<< m1 >>
rect 298 423 299 424 
<< m2 >>
rect 298 423 299 424 
<< m1 >>
rect 318 423 319 424 
<< m1 >>
rect 322 423 323 424 
<< m1 >>
rect 323 423 324 424 
<< m1 >>
rect 325 423 326 424 
<< m1 >>
rect 357 423 358 424 
<< m2 >>
rect 357 423 358 424 
<< m2c >>
rect 357 423 358 424 
<< m1 >>
rect 357 423 358 424 
<< m2 >>
rect 357 423 358 424 
<< m1 >>
rect 358 423 359 424 
<< m1 >>
rect 359 423 360 424 
<< m1 >>
rect 361 423 362 424 
<< m1 >>
rect 379 423 380 424 
<< m2 >>
rect 379 423 380 424 
<< m1 >>
rect 385 423 386 424 
<< m1 >>
rect 391 423 392 424 
<< m1 >>
rect 393 423 394 424 
<< m2 >>
rect 393 423 394 424 
<< m2c >>
rect 393 423 394 424 
<< m1 >>
rect 393 423 394 424 
<< m2 >>
rect 393 423 394 424 
<< m1 >>
rect 394 423 395 424 
<< m1 >>
rect 395 423 396 424 
<< m1 >>
rect 397 423 398 424 
<< m1 >>
rect 402 423 403 424 
<< m1 >>
rect 406 423 407 424 
<< m1 >>
rect 420 423 421 424 
<< m2 >>
rect 420 423 421 424 
<< m2c >>
rect 420 423 421 424 
<< m1 >>
rect 420 423 421 424 
<< m2 >>
rect 420 423 421 424 
<< m1 >>
rect 424 423 425 424 
<< m1 >>
rect 431 423 432 424 
<< m1 >>
rect 433 423 434 424 
<< m1 >>
rect 442 423 443 424 
<< m1 >>
rect 466 423 467 424 
<< m1 >>
rect 472 423 473 424 
<< m1 >>
rect 474 423 475 424 
<< m2 >>
rect 478 423 479 424 
<< m1 >>
rect 480 423 481 424 
<< m1 >>
rect 484 423 485 424 
<< m2 >>
rect 486 423 487 424 
<< m2 >>
rect 487 423 488 424 
<< m2 >>
rect 489 423 490 424 
<< m2 >>
rect 490 423 491 424 
<< m2 >>
rect 491 423 492 424 
<< m1 >>
rect 16 424 17 425 
<< m1 >>
rect 19 424 20 425 
<< m1 >>
rect 21 424 22 425 
<< m1 >>
rect 26 424 27 425 
<< m1 >>
rect 28 424 29 425 
<< m2 >>
rect 28 424 29 425 
<< m1 >>
rect 34 424 35 425 
<< m1 >>
rect 55 424 56 425 
<< m1 >>
rect 56 424 57 425 
<< m1 >>
rect 57 424 58 425 
<< m1 >>
rect 58 424 59 425 
<< m1 >>
rect 59 424 60 425 
<< m1 >>
rect 60 424 61 425 
<< m1 >>
rect 61 424 62 425 
<< m1 >>
rect 62 424 63 425 
<< m1 >>
rect 63 424 64 425 
<< m1 >>
rect 64 424 65 425 
<< m1 >>
rect 65 424 66 425 
<< m1 >>
rect 66 424 67 425 
<< m1 >>
rect 73 424 74 425 
<< m1 >>
rect 82 424 83 425 
<< m1 >>
rect 93 424 94 425 
<< m1 >>
rect 96 424 97 425 
<< m1 >>
rect 100 424 101 425 
<< m1 >>
rect 110 424 111 425 
<< m1 >>
rect 114 424 115 425 
<< m1 >>
rect 118 424 119 425 
<< m1 >>
rect 145 424 146 425 
<< m2 >>
rect 145 424 146 425 
<< m1 >>
rect 150 424 151 425 
<< m2 >>
rect 168 424 169 425 
<< m1 >>
rect 169 424 170 425 
<< m1 >>
rect 171 424 172 425 
<< m1 >>
rect 208 424 209 425 
<< m1 >>
rect 217 424 218 425 
<< m1 >>
rect 253 424 254 425 
<< m1 >>
rect 262 424 263 425 
<< m1 >>
rect 286 424 287 425 
<< m1 >>
rect 287 424 288 425 
<< m1 >>
rect 288 424 289 425 
<< m1 >>
rect 289 424 290 425 
<< m1 >>
rect 290 424 291 425 
<< m1 >>
rect 298 424 299 425 
<< m2 >>
rect 298 424 299 425 
<< m1 >>
rect 304 424 305 425 
<< m1 >>
rect 305 424 306 425 
<< m1 >>
rect 306 424 307 425 
<< m1 >>
rect 307 424 308 425 
<< m1 >>
rect 309 424 310 425 
<< m1 >>
rect 310 424 311 425 
<< m1 >>
rect 311 424 312 425 
<< m1 >>
rect 312 424 313 425 
<< m1 >>
rect 313 424 314 425 
<< m1 >>
rect 314 424 315 425 
<< m1 >>
rect 315 424 316 425 
<< m1 >>
rect 316 424 317 425 
<< m1 >>
rect 317 424 318 425 
<< m1 >>
rect 318 424 319 425 
<< m1 >>
rect 323 424 324 425 
<< m2 >>
rect 323 424 324 425 
<< m2c >>
rect 323 424 324 425 
<< m1 >>
rect 323 424 324 425 
<< m2 >>
rect 323 424 324 425 
<< m2 >>
rect 324 424 325 425 
<< m1 >>
rect 325 424 326 425 
<< m2 >>
rect 325 424 326 425 
<< m2 >>
rect 326 424 327 425 
<< m1 >>
rect 359 424 360 425 
<< m2 >>
rect 359 424 360 425 
<< m2c >>
rect 359 424 360 425 
<< m1 >>
rect 359 424 360 425 
<< m2 >>
rect 359 424 360 425 
<< m2 >>
rect 360 424 361 425 
<< m1 >>
rect 361 424 362 425 
<< m2 >>
rect 361 424 362 425 
<< m1 >>
rect 379 424 380 425 
<< m2 >>
rect 379 424 380 425 
<< m1 >>
rect 385 424 386 425 
<< m1 >>
rect 391 424 392 425 
<< m1 >>
rect 395 424 396 425 
<< m2 >>
rect 395 424 396 425 
<< m2c >>
rect 395 424 396 425 
<< m1 >>
rect 395 424 396 425 
<< m2 >>
rect 395 424 396 425 
<< m2 >>
rect 396 424 397 425 
<< m1 >>
rect 397 424 398 425 
<< m2 >>
rect 397 424 398 425 
<< m2 >>
rect 398 424 399 425 
<< m1 >>
rect 402 424 403 425 
<< m1 >>
rect 406 424 407 425 
<< m1 >>
rect 420 424 421 425 
<< m1 >>
rect 424 424 425 425 
<< m1 >>
rect 431 424 432 425 
<< m2 >>
rect 431 424 432 425 
<< m2c >>
rect 431 424 432 425 
<< m1 >>
rect 431 424 432 425 
<< m2 >>
rect 431 424 432 425 
<< m2 >>
rect 432 424 433 425 
<< m1 >>
rect 433 424 434 425 
<< m2 >>
rect 433 424 434 425 
<< m2 >>
rect 434 424 435 425 
<< m1 >>
rect 442 424 443 425 
<< m1 >>
rect 448 424 449 425 
<< m1 >>
rect 449 424 450 425 
<< m1 >>
rect 450 424 451 425 
<< m1 >>
rect 451 424 452 425 
<< m1 >>
rect 452 424 453 425 
<< m1 >>
rect 466 424 467 425 
<< m1 >>
rect 472 424 473 425 
<< m2 >>
rect 473 424 474 425 
<< m1 >>
rect 474 424 475 425 
<< m2 >>
rect 474 424 475 425 
<< m2 >>
rect 475 424 476 425 
<< m1 >>
rect 476 424 477 425 
<< m2 >>
rect 476 424 477 425 
<< m2c >>
rect 476 424 477 425 
<< m1 >>
rect 476 424 477 425 
<< m2 >>
rect 476 424 477 425 
<< m1 >>
rect 477 424 478 425 
<< m1 >>
rect 478 424 479 425 
<< m2 >>
rect 478 424 479 425 
<< m1 >>
rect 479 424 480 425 
<< m1 >>
rect 480 424 481 425 
<< m1 >>
rect 484 424 485 425 
<< m1 >>
rect 487 424 488 425 
<< m2 >>
rect 487 424 488 425 
<< m1 >>
rect 488 424 489 425 
<< m1 >>
rect 489 424 490 425 
<< m1 >>
rect 490 424 491 425 
<< m1 >>
rect 491 424 492 425 
<< m2 >>
rect 491 424 492 425 
<< m1 >>
rect 492 424 493 425 
<< m1 >>
rect 493 424 494 425 
<< m1 >>
rect 494 424 495 425 
<< m1 >>
rect 495 424 496 425 
<< m1 >>
rect 496 424 497 425 
<< m1 >>
rect 497 424 498 425 
<< m1 >>
rect 498 424 499 425 
<< m1 >>
rect 499 424 500 425 
<< m1 >>
rect 16 425 17 426 
<< m1 >>
rect 19 425 20 426 
<< m1 >>
rect 21 425 22 426 
<< m1 >>
rect 26 425 27 426 
<< m1 >>
rect 28 425 29 426 
<< m2 >>
rect 28 425 29 426 
<< m1 >>
rect 34 425 35 426 
<< m1 >>
rect 55 425 56 426 
<< m1 >>
rect 73 425 74 426 
<< m1 >>
rect 82 425 83 426 
<< m1 >>
rect 93 425 94 426 
<< m1 >>
rect 96 425 97 426 
<< m1 >>
rect 100 425 101 426 
<< m1 >>
rect 110 425 111 426 
<< m1 >>
rect 114 425 115 426 
<< m1 >>
rect 118 425 119 426 
<< m1 >>
rect 145 425 146 426 
<< m2 >>
rect 145 425 146 426 
<< m1 >>
rect 150 425 151 426 
<< m2 >>
rect 168 425 169 426 
<< m1 >>
rect 169 425 170 426 
<< m1 >>
rect 171 425 172 426 
<< m1 >>
rect 208 425 209 426 
<< m1 >>
rect 217 425 218 426 
<< m1 >>
rect 253 425 254 426 
<< m2 >>
rect 254 425 255 426 
<< m1 >>
rect 255 425 256 426 
<< m2 >>
rect 255 425 256 426 
<< m2c >>
rect 255 425 256 426 
<< m1 >>
rect 255 425 256 426 
<< m2 >>
rect 255 425 256 426 
<< m1 >>
rect 256 425 257 426 
<< m1 >>
rect 257 425 258 426 
<< m1 >>
rect 258 425 259 426 
<< m1 >>
rect 259 425 260 426 
<< m1 >>
rect 260 425 261 426 
<< m1 >>
rect 261 425 262 426 
<< m1 >>
rect 262 425 263 426 
<< m1 >>
rect 286 425 287 426 
<< m1 >>
rect 290 425 291 426 
<< m1 >>
rect 298 425 299 426 
<< m2 >>
rect 298 425 299 426 
<< m1 >>
rect 304 425 305 426 
<< m1 >>
rect 307 425 308 426 
<< m1 >>
rect 309 425 310 426 
<< m1 >>
rect 325 425 326 426 
<< m2 >>
rect 326 425 327 426 
<< m1 >>
rect 361 425 362 426 
<< m2 >>
rect 361 425 362 426 
<< m1 >>
rect 379 425 380 426 
<< m2 >>
rect 379 425 380 426 
<< m1 >>
rect 385 425 386 426 
<< m1 >>
rect 391 425 392 426 
<< m1 >>
rect 397 425 398 426 
<< m2 >>
rect 398 425 399 426 
<< m1 >>
rect 402 425 403 426 
<< m1 >>
rect 406 425 407 426 
<< m1 >>
rect 420 425 421 426 
<< m1 >>
rect 424 425 425 426 
<< m1 >>
rect 433 425 434 426 
<< m2 >>
rect 434 425 435 426 
<< m1 >>
rect 442 425 443 426 
<< m1 >>
rect 448 425 449 426 
<< m1 >>
rect 452 425 453 426 
<< m1 >>
rect 466 425 467 426 
<< m1 >>
rect 472 425 473 426 
<< m2 >>
rect 473 425 474 426 
<< m1 >>
rect 474 425 475 426 
<< m2 >>
rect 478 425 479 426 
<< m1 >>
rect 484 425 485 426 
<< m1 >>
rect 487 425 488 426 
<< m2 >>
rect 487 425 488 426 
<< m2 >>
rect 491 425 492 426 
<< m1 >>
rect 499 425 500 426 
<< pdiffusion >>
rect 12 426 13 427 
<< pdiffusion >>
rect 13 426 14 427 
<< pdiffusion >>
rect 14 426 15 427 
<< pdiffusion >>
rect 15 426 16 427 
<< m1 >>
rect 16 426 17 427 
<< pdiffusion >>
rect 16 426 17 427 
<< pdiffusion >>
rect 17 426 18 427 
<< m1 >>
rect 19 426 20 427 
<< m1 >>
rect 21 426 22 427 
<< m1 >>
rect 26 426 27 427 
<< m1 >>
rect 28 426 29 427 
<< m2 >>
rect 28 426 29 427 
<< pdiffusion >>
rect 30 426 31 427 
<< pdiffusion >>
rect 31 426 32 427 
<< pdiffusion >>
rect 32 426 33 427 
<< pdiffusion >>
rect 33 426 34 427 
<< m1 >>
rect 34 426 35 427 
<< pdiffusion >>
rect 34 426 35 427 
<< pdiffusion >>
rect 35 426 36 427 
<< pdiffusion >>
rect 48 426 49 427 
<< pdiffusion >>
rect 49 426 50 427 
<< pdiffusion >>
rect 50 426 51 427 
<< pdiffusion >>
rect 51 426 52 427 
<< pdiffusion >>
rect 52 426 53 427 
<< pdiffusion >>
rect 53 426 54 427 
<< m1 >>
rect 55 426 56 427 
<< pdiffusion >>
rect 66 426 67 427 
<< pdiffusion >>
rect 67 426 68 427 
<< pdiffusion >>
rect 68 426 69 427 
<< pdiffusion >>
rect 69 426 70 427 
<< pdiffusion >>
rect 70 426 71 427 
<< pdiffusion >>
rect 71 426 72 427 
<< m1 >>
rect 73 426 74 427 
<< m1 >>
rect 82 426 83 427 
<< pdiffusion >>
rect 84 426 85 427 
<< pdiffusion >>
rect 85 426 86 427 
<< pdiffusion >>
rect 86 426 87 427 
<< pdiffusion >>
rect 87 426 88 427 
<< pdiffusion >>
rect 88 426 89 427 
<< pdiffusion >>
rect 89 426 90 427 
<< m1 >>
rect 93 426 94 427 
<< m1 >>
rect 96 426 97 427 
<< m1 >>
rect 100 426 101 427 
<< pdiffusion >>
rect 102 426 103 427 
<< pdiffusion >>
rect 103 426 104 427 
<< pdiffusion >>
rect 104 426 105 427 
<< pdiffusion >>
rect 105 426 106 427 
<< pdiffusion >>
rect 106 426 107 427 
<< pdiffusion >>
rect 107 426 108 427 
<< m1 >>
rect 110 426 111 427 
<< m1 >>
rect 114 426 115 427 
<< m1 >>
rect 118 426 119 427 
<< pdiffusion >>
rect 120 426 121 427 
<< pdiffusion >>
rect 121 426 122 427 
<< pdiffusion >>
rect 122 426 123 427 
<< pdiffusion >>
rect 123 426 124 427 
<< pdiffusion >>
rect 124 426 125 427 
<< pdiffusion >>
rect 125 426 126 427 
<< pdiffusion >>
rect 138 426 139 427 
<< pdiffusion >>
rect 139 426 140 427 
<< pdiffusion >>
rect 140 426 141 427 
<< pdiffusion >>
rect 141 426 142 427 
<< pdiffusion >>
rect 142 426 143 427 
<< pdiffusion >>
rect 143 426 144 427 
<< m1 >>
rect 145 426 146 427 
<< m2 >>
rect 145 426 146 427 
<< m1 >>
rect 150 426 151 427 
<< pdiffusion >>
rect 156 426 157 427 
<< pdiffusion >>
rect 157 426 158 427 
<< pdiffusion >>
rect 158 426 159 427 
<< pdiffusion >>
rect 159 426 160 427 
<< pdiffusion >>
rect 160 426 161 427 
<< pdiffusion >>
rect 161 426 162 427 
<< m2 >>
rect 168 426 169 427 
<< m1 >>
rect 169 426 170 427 
<< m1 >>
rect 171 426 172 427 
<< pdiffusion >>
rect 174 426 175 427 
<< pdiffusion >>
rect 175 426 176 427 
<< pdiffusion >>
rect 176 426 177 427 
<< pdiffusion >>
rect 177 426 178 427 
<< pdiffusion >>
rect 178 426 179 427 
<< pdiffusion >>
rect 179 426 180 427 
<< pdiffusion >>
rect 192 426 193 427 
<< pdiffusion >>
rect 193 426 194 427 
<< pdiffusion >>
rect 194 426 195 427 
<< pdiffusion >>
rect 195 426 196 427 
<< pdiffusion >>
rect 196 426 197 427 
<< pdiffusion >>
rect 197 426 198 427 
<< m1 >>
rect 208 426 209 427 
<< pdiffusion >>
rect 210 426 211 427 
<< pdiffusion >>
rect 211 426 212 427 
<< pdiffusion >>
rect 212 426 213 427 
<< pdiffusion >>
rect 213 426 214 427 
<< pdiffusion >>
rect 214 426 215 427 
<< pdiffusion >>
rect 215 426 216 427 
<< m1 >>
rect 217 426 218 427 
<< pdiffusion >>
rect 228 426 229 427 
<< pdiffusion >>
rect 229 426 230 427 
<< pdiffusion >>
rect 230 426 231 427 
<< pdiffusion >>
rect 231 426 232 427 
<< pdiffusion >>
rect 232 426 233 427 
<< pdiffusion >>
rect 233 426 234 427 
<< pdiffusion >>
rect 246 426 247 427 
<< pdiffusion >>
rect 247 426 248 427 
<< pdiffusion >>
rect 248 426 249 427 
<< pdiffusion >>
rect 249 426 250 427 
<< pdiffusion >>
rect 250 426 251 427 
<< pdiffusion >>
rect 251 426 252 427 
<< m1 >>
rect 253 426 254 427 
<< m2 >>
rect 254 426 255 427 
<< pdiffusion >>
rect 264 426 265 427 
<< pdiffusion >>
rect 265 426 266 427 
<< pdiffusion >>
rect 266 426 267 427 
<< pdiffusion >>
rect 267 426 268 427 
<< pdiffusion >>
rect 268 426 269 427 
<< pdiffusion >>
rect 269 426 270 427 
<< pdiffusion >>
rect 282 426 283 427 
<< pdiffusion >>
rect 283 426 284 427 
<< pdiffusion >>
rect 284 426 285 427 
<< pdiffusion >>
rect 285 426 286 427 
<< m1 >>
rect 286 426 287 427 
<< pdiffusion >>
rect 286 426 287 427 
<< pdiffusion >>
rect 287 426 288 427 
<< m1 >>
rect 290 426 291 427 
<< m1 >>
rect 298 426 299 427 
<< m2 >>
rect 298 426 299 427 
<< pdiffusion >>
rect 300 426 301 427 
<< pdiffusion >>
rect 301 426 302 427 
<< pdiffusion >>
rect 302 426 303 427 
<< pdiffusion >>
rect 303 426 304 427 
<< m1 >>
rect 304 426 305 427 
<< pdiffusion >>
rect 304 426 305 427 
<< pdiffusion >>
rect 305 426 306 427 
<< m1 >>
rect 307 426 308 427 
<< m1 >>
rect 309 426 310 427 
<< pdiffusion >>
rect 318 426 319 427 
<< pdiffusion >>
rect 319 426 320 427 
<< pdiffusion >>
rect 320 426 321 427 
<< pdiffusion >>
rect 321 426 322 427 
<< pdiffusion >>
rect 322 426 323 427 
<< pdiffusion >>
rect 323 426 324 427 
<< m1 >>
rect 325 426 326 427 
<< m2 >>
rect 326 426 327 427 
<< pdiffusion >>
rect 336 426 337 427 
<< pdiffusion >>
rect 337 426 338 427 
<< pdiffusion >>
rect 338 426 339 427 
<< pdiffusion >>
rect 339 426 340 427 
<< pdiffusion >>
rect 340 426 341 427 
<< pdiffusion >>
rect 341 426 342 427 
<< pdiffusion >>
rect 354 426 355 427 
<< pdiffusion >>
rect 355 426 356 427 
<< pdiffusion >>
rect 356 426 357 427 
<< pdiffusion >>
rect 357 426 358 427 
<< pdiffusion >>
rect 358 426 359 427 
<< pdiffusion >>
rect 359 426 360 427 
<< m1 >>
rect 361 426 362 427 
<< m2 >>
rect 361 426 362 427 
<< pdiffusion >>
rect 372 426 373 427 
<< pdiffusion >>
rect 373 426 374 427 
<< pdiffusion >>
rect 374 426 375 427 
<< pdiffusion >>
rect 375 426 376 427 
<< pdiffusion >>
rect 376 426 377 427 
<< pdiffusion >>
rect 377 426 378 427 
<< m1 >>
rect 379 426 380 427 
<< m2 >>
rect 379 426 380 427 
<< m1 >>
rect 385 426 386 427 
<< pdiffusion >>
rect 390 426 391 427 
<< m1 >>
rect 391 426 392 427 
<< pdiffusion >>
rect 391 426 392 427 
<< pdiffusion >>
rect 392 426 393 427 
<< pdiffusion >>
rect 393 426 394 427 
<< pdiffusion >>
rect 394 426 395 427 
<< pdiffusion >>
rect 395 426 396 427 
<< m1 >>
rect 397 426 398 427 
<< m2 >>
rect 398 426 399 427 
<< m1 >>
rect 402 426 403 427 
<< m1 >>
rect 406 426 407 427 
<< pdiffusion >>
rect 408 426 409 427 
<< pdiffusion >>
rect 409 426 410 427 
<< pdiffusion >>
rect 410 426 411 427 
<< pdiffusion >>
rect 411 426 412 427 
<< pdiffusion >>
rect 412 426 413 427 
<< pdiffusion >>
rect 413 426 414 427 
<< m1 >>
rect 420 426 421 427 
<< m1 >>
rect 424 426 425 427 
<< pdiffusion >>
rect 426 426 427 427 
<< pdiffusion >>
rect 427 426 428 427 
<< pdiffusion >>
rect 428 426 429 427 
<< pdiffusion >>
rect 429 426 430 427 
<< pdiffusion >>
rect 430 426 431 427 
<< pdiffusion >>
rect 431 426 432 427 
<< m1 >>
rect 433 426 434 427 
<< m2 >>
rect 434 426 435 427 
<< m1 >>
rect 442 426 443 427 
<< pdiffusion >>
rect 444 426 445 427 
<< pdiffusion >>
rect 445 426 446 427 
<< pdiffusion >>
rect 446 426 447 427 
<< pdiffusion >>
rect 447 426 448 427 
<< m1 >>
rect 448 426 449 427 
<< pdiffusion >>
rect 448 426 449 427 
<< pdiffusion >>
rect 449 426 450 427 
<< m1 >>
rect 452 426 453 427 
<< pdiffusion >>
rect 462 426 463 427 
<< pdiffusion >>
rect 463 426 464 427 
<< pdiffusion >>
rect 464 426 465 427 
<< pdiffusion >>
rect 465 426 466 427 
<< m1 >>
rect 466 426 467 427 
<< pdiffusion >>
rect 466 426 467 427 
<< pdiffusion >>
rect 467 426 468 427 
<< m1 >>
rect 472 426 473 427 
<< m2 >>
rect 473 426 474 427 
<< m1 >>
rect 474 426 475 427 
<< m1 >>
rect 478 426 479 427 
<< m2 >>
rect 478 426 479 427 
<< m2c >>
rect 478 426 479 427 
<< m1 >>
rect 478 426 479 427 
<< m2 >>
rect 478 426 479 427 
<< pdiffusion >>
rect 480 426 481 427 
<< pdiffusion >>
rect 481 426 482 427 
<< pdiffusion >>
rect 482 426 483 427 
<< pdiffusion >>
rect 483 426 484 427 
<< m1 >>
rect 484 426 485 427 
<< pdiffusion >>
rect 484 426 485 427 
<< pdiffusion >>
rect 485 426 486 427 
<< m1 >>
rect 487 426 488 427 
<< m2 >>
rect 487 426 488 427 
<< m2 >>
rect 488 426 489 427 
<< m1 >>
rect 489 426 490 427 
<< m2 >>
rect 489 426 490 427 
<< m2c >>
rect 489 426 490 427 
<< m1 >>
rect 489 426 490 427 
<< m2 >>
rect 489 426 490 427 
<< m1 >>
rect 491 426 492 427 
<< m2 >>
rect 491 426 492 427 
<< m2c >>
rect 491 426 492 427 
<< m1 >>
rect 491 426 492 427 
<< m2 >>
rect 491 426 492 427 
<< pdiffusion >>
rect 498 426 499 427 
<< m1 >>
rect 499 426 500 427 
<< pdiffusion >>
rect 499 426 500 427 
<< pdiffusion >>
rect 500 426 501 427 
<< pdiffusion >>
rect 501 426 502 427 
<< pdiffusion >>
rect 502 426 503 427 
<< pdiffusion >>
rect 503 426 504 427 
<< pdiffusion >>
rect 516 426 517 427 
<< pdiffusion >>
rect 517 426 518 427 
<< pdiffusion >>
rect 518 426 519 427 
<< pdiffusion >>
rect 519 426 520 427 
<< pdiffusion >>
rect 520 426 521 427 
<< pdiffusion >>
rect 521 426 522 427 
<< pdiffusion >>
rect 12 427 13 428 
<< pdiffusion >>
rect 13 427 14 428 
<< pdiffusion >>
rect 14 427 15 428 
<< pdiffusion >>
rect 15 427 16 428 
<< pdiffusion >>
rect 16 427 17 428 
<< pdiffusion >>
rect 17 427 18 428 
<< m1 >>
rect 19 427 20 428 
<< m1 >>
rect 21 427 22 428 
<< m1 >>
rect 26 427 27 428 
<< m1 >>
rect 28 427 29 428 
<< m2 >>
rect 28 427 29 428 
<< pdiffusion >>
rect 30 427 31 428 
<< pdiffusion >>
rect 31 427 32 428 
<< pdiffusion >>
rect 32 427 33 428 
<< pdiffusion >>
rect 33 427 34 428 
<< pdiffusion >>
rect 34 427 35 428 
<< pdiffusion >>
rect 35 427 36 428 
<< pdiffusion >>
rect 48 427 49 428 
<< pdiffusion >>
rect 49 427 50 428 
<< pdiffusion >>
rect 50 427 51 428 
<< pdiffusion >>
rect 51 427 52 428 
<< pdiffusion >>
rect 52 427 53 428 
<< pdiffusion >>
rect 53 427 54 428 
<< m1 >>
rect 55 427 56 428 
<< pdiffusion >>
rect 66 427 67 428 
<< pdiffusion >>
rect 67 427 68 428 
<< pdiffusion >>
rect 68 427 69 428 
<< pdiffusion >>
rect 69 427 70 428 
<< pdiffusion >>
rect 70 427 71 428 
<< pdiffusion >>
rect 71 427 72 428 
<< m1 >>
rect 73 427 74 428 
<< m1 >>
rect 82 427 83 428 
<< pdiffusion >>
rect 84 427 85 428 
<< pdiffusion >>
rect 85 427 86 428 
<< pdiffusion >>
rect 86 427 87 428 
<< pdiffusion >>
rect 87 427 88 428 
<< pdiffusion >>
rect 88 427 89 428 
<< pdiffusion >>
rect 89 427 90 428 
<< m1 >>
rect 93 427 94 428 
<< m1 >>
rect 96 427 97 428 
<< m1 >>
rect 100 427 101 428 
<< pdiffusion >>
rect 102 427 103 428 
<< pdiffusion >>
rect 103 427 104 428 
<< pdiffusion >>
rect 104 427 105 428 
<< pdiffusion >>
rect 105 427 106 428 
<< pdiffusion >>
rect 106 427 107 428 
<< pdiffusion >>
rect 107 427 108 428 
<< m1 >>
rect 110 427 111 428 
<< m1 >>
rect 114 427 115 428 
<< m1 >>
rect 118 427 119 428 
<< pdiffusion >>
rect 120 427 121 428 
<< pdiffusion >>
rect 121 427 122 428 
<< pdiffusion >>
rect 122 427 123 428 
<< pdiffusion >>
rect 123 427 124 428 
<< pdiffusion >>
rect 124 427 125 428 
<< pdiffusion >>
rect 125 427 126 428 
<< pdiffusion >>
rect 138 427 139 428 
<< pdiffusion >>
rect 139 427 140 428 
<< pdiffusion >>
rect 140 427 141 428 
<< pdiffusion >>
rect 141 427 142 428 
<< pdiffusion >>
rect 142 427 143 428 
<< pdiffusion >>
rect 143 427 144 428 
<< m1 >>
rect 145 427 146 428 
<< m2 >>
rect 145 427 146 428 
<< m1 >>
rect 150 427 151 428 
<< pdiffusion >>
rect 156 427 157 428 
<< pdiffusion >>
rect 157 427 158 428 
<< pdiffusion >>
rect 158 427 159 428 
<< pdiffusion >>
rect 159 427 160 428 
<< pdiffusion >>
rect 160 427 161 428 
<< pdiffusion >>
rect 161 427 162 428 
<< m2 >>
rect 168 427 169 428 
<< m1 >>
rect 169 427 170 428 
<< m1 >>
rect 171 427 172 428 
<< pdiffusion >>
rect 174 427 175 428 
<< pdiffusion >>
rect 175 427 176 428 
<< pdiffusion >>
rect 176 427 177 428 
<< pdiffusion >>
rect 177 427 178 428 
<< pdiffusion >>
rect 178 427 179 428 
<< pdiffusion >>
rect 179 427 180 428 
<< pdiffusion >>
rect 192 427 193 428 
<< pdiffusion >>
rect 193 427 194 428 
<< pdiffusion >>
rect 194 427 195 428 
<< pdiffusion >>
rect 195 427 196 428 
<< pdiffusion >>
rect 196 427 197 428 
<< pdiffusion >>
rect 197 427 198 428 
<< m1 >>
rect 208 427 209 428 
<< pdiffusion >>
rect 210 427 211 428 
<< pdiffusion >>
rect 211 427 212 428 
<< pdiffusion >>
rect 212 427 213 428 
<< pdiffusion >>
rect 213 427 214 428 
<< pdiffusion >>
rect 214 427 215 428 
<< pdiffusion >>
rect 215 427 216 428 
<< m1 >>
rect 217 427 218 428 
<< pdiffusion >>
rect 228 427 229 428 
<< pdiffusion >>
rect 229 427 230 428 
<< pdiffusion >>
rect 230 427 231 428 
<< pdiffusion >>
rect 231 427 232 428 
<< pdiffusion >>
rect 232 427 233 428 
<< pdiffusion >>
rect 233 427 234 428 
<< pdiffusion >>
rect 246 427 247 428 
<< pdiffusion >>
rect 247 427 248 428 
<< pdiffusion >>
rect 248 427 249 428 
<< pdiffusion >>
rect 249 427 250 428 
<< pdiffusion >>
rect 250 427 251 428 
<< pdiffusion >>
rect 251 427 252 428 
<< m1 >>
rect 253 427 254 428 
<< m2 >>
rect 254 427 255 428 
<< pdiffusion >>
rect 264 427 265 428 
<< pdiffusion >>
rect 265 427 266 428 
<< pdiffusion >>
rect 266 427 267 428 
<< pdiffusion >>
rect 267 427 268 428 
<< pdiffusion >>
rect 268 427 269 428 
<< pdiffusion >>
rect 269 427 270 428 
<< pdiffusion >>
rect 282 427 283 428 
<< pdiffusion >>
rect 283 427 284 428 
<< pdiffusion >>
rect 284 427 285 428 
<< pdiffusion >>
rect 285 427 286 428 
<< pdiffusion >>
rect 286 427 287 428 
<< pdiffusion >>
rect 287 427 288 428 
<< m1 >>
rect 290 427 291 428 
<< m1 >>
rect 298 427 299 428 
<< m2 >>
rect 298 427 299 428 
<< pdiffusion >>
rect 300 427 301 428 
<< pdiffusion >>
rect 301 427 302 428 
<< pdiffusion >>
rect 302 427 303 428 
<< pdiffusion >>
rect 303 427 304 428 
<< pdiffusion >>
rect 304 427 305 428 
<< pdiffusion >>
rect 305 427 306 428 
<< m1 >>
rect 307 427 308 428 
<< m1 >>
rect 309 427 310 428 
<< pdiffusion >>
rect 318 427 319 428 
<< pdiffusion >>
rect 319 427 320 428 
<< pdiffusion >>
rect 320 427 321 428 
<< pdiffusion >>
rect 321 427 322 428 
<< pdiffusion >>
rect 322 427 323 428 
<< pdiffusion >>
rect 323 427 324 428 
<< m1 >>
rect 325 427 326 428 
<< m2 >>
rect 326 427 327 428 
<< pdiffusion >>
rect 336 427 337 428 
<< pdiffusion >>
rect 337 427 338 428 
<< pdiffusion >>
rect 338 427 339 428 
<< pdiffusion >>
rect 339 427 340 428 
<< pdiffusion >>
rect 340 427 341 428 
<< pdiffusion >>
rect 341 427 342 428 
<< pdiffusion >>
rect 354 427 355 428 
<< pdiffusion >>
rect 355 427 356 428 
<< pdiffusion >>
rect 356 427 357 428 
<< pdiffusion >>
rect 357 427 358 428 
<< pdiffusion >>
rect 358 427 359 428 
<< pdiffusion >>
rect 359 427 360 428 
<< m1 >>
rect 361 427 362 428 
<< m2 >>
rect 361 427 362 428 
<< pdiffusion >>
rect 372 427 373 428 
<< pdiffusion >>
rect 373 427 374 428 
<< pdiffusion >>
rect 374 427 375 428 
<< pdiffusion >>
rect 375 427 376 428 
<< pdiffusion >>
rect 376 427 377 428 
<< pdiffusion >>
rect 377 427 378 428 
<< m1 >>
rect 379 427 380 428 
<< m2 >>
rect 379 427 380 428 
<< m1 >>
rect 385 427 386 428 
<< pdiffusion >>
rect 390 427 391 428 
<< pdiffusion >>
rect 391 427 392 428 
<< pdiffusion >>
rect 392 427 393 428 
<< pdiffusion >>
rect 393 427 394 428 
<< pdiffusion >>
rect 394 427 395 428 
<< pdiffusion >>
rect 395 427 396 428 
<< m1 >>
rect 397 427 398 428 
<< m2 >>
rect 398 427 399 428 
<< m1 >>
rect 402 427 403 428 
<< m1 >>
rect 406 427 407 428 
<< pdiffusion >>
rect 408 427 409 428 
<< pdiffusion >>
rect 409 427 410 428 
<< pdiffusion >>
rect 410 427 411 428 
<< pdiffusion >>
rect 411 427 412 428 
<< pdiffusion >>
rect 412 427 413 428 
<< pdiffusion >>
rect 413 427 414 428 
<< m1 >>
rect 420 427 421 428 
<< m1 >>
rect 424 427 425 428 
<< pdiffusion >>
rect 426 427 427 428 
<< pdiffusion >>
rect 427 427 428 428 
<< pdiffusion >>
rect 428 427 429 428 
<< pdiffusion >>
rect 429 427 430 428 
<< pdiffusion >>
rect 430 427 431 428 
<< pdiffusion >>
rect 431 427 432 428 
<< m1 >>
rect 433 427 434 428 
<< m2 >>
rect 434 427 435 428 
<< m1 >>
rect 442 427 443 428 
<< pdiffusion >>
rect 444 427 445 428 
<< pdiffusion >>
rect 445 427 446 428 
<< pdiffusion >>
rect 446 427 447 428 
<< pdiffusion >>
rect 447 427 448 428 
<< pdiffusion >>
rect 448 427 449 428 
<< pdiffusion >>
rect 449 427 450 428 
<< m1 >>
rect 452 427 453 428 
<< pdiffusion >>
rect 462 427 463 428 
<< pdiffusion >>
rect 463 427 464 428 
<< pdiffusion >>
rect 464 427 465 428 
<< pdiffusion >>
rect 465 427 466 428 
<< pdiffusion >>
rect 466 427 467 428 
<< pdiffusion >>
rect 467 427 468 428 
<< m1 >>
rect 472 427 473 428 
<< m2 >>
rect 473 427 474 428 
<< m1 >>
rect 474 427 475 428 
<< m1 >>
rect 478 427 479 428 
<< pdiffusion >>
rect 480 427 481 428 
<< pdiffusion >>
rect 481 427 482 428 
<< pdiffusion >>
rect 482 427 483 428 
<< pdiffusion >>
rect 483 427 484 428 
<< pdiffusion >>
rect 484 427 485 428 
<< pdiffusion >>
rect 485 427 486 428 
<< m1 >>
rect 487 427 488 428 
<< m1 >>
rect 489 427 490 428 
<< m1 >>
rect 491 427 492 428 
<< pdiffusion >>
rect 498 427 499 428 
<< pdiffusion >>
rect 499 427 500 428 
<< pdiffusion >>
rect 500 427 501 428 
<< pdiffusion >>
rect 501 427 502 428 
<< pdiffusion >>
rect 502 427 503 428 
<< pdiffusion >>
rect 503 427 504 428 
<< pdiffusion >>
rect 516 427 517 428 
<< pdiffusion >>
rect 517 427 518 428 
<< pdiffusion >>
rect 518 427 519 428 
<< pdiffusion >>
rect 519 427 520 428 
<< pdiffusion >>
rect 520 427 521 428 
<< pdiffusion >>
rect 521 427 522 428 
<< pdiffusion >>
rect 12 428 13 429 
<< pdiffusion >>
rect 13 428 14 429 
<< pdiffusion >>
rect 14 428 15 429 
<< pdiffusion >>
rect 15 428 16 429 
<< pdiffusion >>
rect 16 428 17 429 
<< pdiffusion >>
rect 17 428 18 429 
<< m1 >>
rect 19 428 20 429 
<< m1 >>
rect 21 428 22 429 
<< m1 >>
rect 26 428 27 429 
<< m1 >>
rect 28 428 29 429 
<< m2 >>
rect 28 428 29 429 
<< pdiffusion >>
rect 30 428 31 429 
<< pdiffusion >>
rect 31 428 32 429 
<< pdiffusion >>
rect 32 428 33 429 
<< pdiffusion >>
rect 33 428 34 429 
<< pdiffusion >>
rect 34 428 35 429 
<< pdiffusion >>
rect 35 428 36 429 
<< pdiffusion >>
rect 48 428 49 429 
<< pdiffusion >>
rect 49 428 50 429 
<< pdiffusion >>
rect 50 428 51 429 
<< pdiffusion >>
rect 51 428 52 429 
<< pdiffusion >>
rect 52 428 53 429 
<< pdiffusion >>
rect 53 428 54 429 
<< m1 >>
rect 55 428 56 429 
<< pdiffusion >>
rect 66 428 67 429 
<< pdiffusion >>
rect 67 428 68 429 
<< pdiffusion >>
rect 68 428 69 429 
<< pdiffusion >>
rect 69 428 70 429 
<< pdiffusion >>
rect 70 428 71 429 
<< pdiffusion >>
rect 71 428 72 429 
<< m1 >>
rect 73 428 74 429 
<< m1 >>
rect 82 428 83 429 
<< pdiffusion >>
rect 84 428 85 429 
<< pdiffusion >>
rect 85 428 86 429 
<< pdiffusion >>
rect 86 428 87 429 
<< pdiffusion >>
rect 87 428 88 429 
<< pdiffusion >>
rect 88 428 89 429 
<< pdiffusion >>
rect 89 428 90 429 
<< m1 >>
rect 93 428 94 429 
<< m1 >>
rect 96 428 97 429 
<< m1 >>
rect 100 428 101 429 
<< pdiffusion >>
rect 102 428 103 429 
<< pdiffusion >>
rect 103 428 104 429 
<< pdiffusion >>
rect 104 428 105 429 
<< pdiffusion >>
rect 105 428 106 429 
<< pdiffusion >>
rect 106 428 107 429 
<< pdiffusion >>
rect 107 428 108 429 
<< m1 >>
rect 110 428 111 429 
<< m1 >>
rect 114 428 115 429 
<< m1 >>
rect 118 428 119 429 
<< pdiffusion >>
rect 120 428 121 429 
<< pdiffusion >>
rect 121 428 122 429 
<< pdiffusion >>
rect 122 428 123 429 
<< pdiffusion >>
rect 123 428 124 429 
<< pdiffusion >>
rect 124 428 125 429 
<< pdiffusion >>
rect 125 428 126 429 
<< pdiffusion >>
rect 138 428 139 429 
<< pdiffusion >>
rect 139 428 140 429 
<< pdiffusion >>
rect 140 428 141 429 
<< pdiffusion >>
rect 141 428 142 429 
<< pdiffusion >>
rect 142 428 143 429 
<< pdiffusion >>
rect 143 428 144 429 
<< m1 >>
rect 145 428 146 429 
<< m2 >>
rect 145 428 146 429 
<< m1 >>
rect 150 428 151 429 
<< pdiffusion >>
rect 156 428 157 429 
<< pdiffusion >>
rect 157 428 158 429 
<< pdiffusion >>
rect 158 428 159 429 
<< pdiffusion >>
rect 159 428 160 429 
<< pdiffusion >>
rect 160 428 161 429 
<< pdiffusion >>
rect 161 428 162 429 
<< m2 >>
rect 168 428 169 429 
<< m1 >>
rect 169 428 170 429 
<< m1 >>
rect 171 428 172 429 
<< pdiffusion >>
rect 174 428 175 429 
<< pdiffusion >>
rect 175 428 176 429 
<< pdiffusion >>
rect 176 428 177 429 
<< pdiffusion >>
rect 177 428 178 429 
<< pdiffusion >>
rect 178 428 179 429 
<< pdiffusion >>
rect 179 428 180 429 
<< pdiffusion >>
rect 192 428 193 429 
<< pdiffusion >>
rect 193 428 194 429 
<< pdiffusion >>
rect 194 428 195 429 
<< pdiffusion >>
rect 195 428 196 429 
<< pdiffusion >>
rect 196 428 197 429 
<< pdiffusion >>
rect 197 428 198 429 
<< m1 >>
rect 208 428 209 429 
<< pdiffusion >>
rect 210 428 211 429 
<< pdiffusion >>
rect 211 428 212 429 
<< pdiffusion >>
rect 212 428 213 429 
<< pdiffusion >>
rect 213 428 214 429 
<< pdiffusion >>
rect 214 428 215 429 
<< pdiffusion >>
rect 215 428 216 429 
<< m1 >>
rect 217 428 218 429 
<< pdiffusion >>
rect 228 428 229 429 
<< pdiffusion >>
rect 229 428 230 429 
<< pdiffusion >>
rect 230 428 231 429 
<< pdiffusion >>
rect 231 428 232 429 
<< pdiffusion >>
rect 232 428 233 429 
<< pdiffusion >>
rect 233 428 234 429 
<< pdiffusion >>
rect 246 428 247 429 
<< pdiffusion >>
rect 247 428 248 429 
<< pdiffusion >>
rect 248 428 249 429 
<< pdiffusion >>
rect 249 428 250 429 
<< pdiffusion >>
rect 250 428 251 429 
<< pdiffusion >>
rect 251 428 252 429 
<< m1 >>
rect 253 428 254 429 
<< m2 >>
rect 254 428 255 429 
<< pdiffusion >>
rect 264 428 265 429 
<< pdiffusion >>
rect 265 428 266 429 
<< pdiffusion >>
rect 266 428 267 429 
<< pdiffusion >>
rect 267 428 268 429 
<< pdiffusion >>
rect 268 428 269 429 
<< pdiffusion >>
rect 269 428 270 429 
<< pdiffusion >>
rect 282 428 283 429 
<< pdiffusion >>
rect 283 428 284 429 
<< pdiffusion >>
rect 284 428 285 429 
<< pdiffusion >>
rect 285 428 286 429 
<< pdiffusion >>
rect 286 428 287 429 
<< pdiffusion >>
rect 287 428 288 429 
<< m1 >>
rect 290 428 291 429 
<< m1 >>
rect 298 428 299 429 
<< m2 >>
rect 298 428 299 429 
<< pdiffusion >>
rect 300 428 301 429 
<< pdiffusion >>
rect 301 428 302 429 
<< pdiffusion >>
rect 302 428 303 429 
<< pdiffusion >>
rect 303 428 304 429 
<< pdiffusion >>
rect 304 428 305 429 
<< pdiffusion >>
rect 305 428 306 429 
<< m1 >>
rect 307 428 308 429 
<< m1 >>
rect 309 428 310 429 
<< pdiffusion >>
rect 318 428 319 429 
<< pdiffusion >>
rect 319 428 320 429 
<< pdiffusion >>
rect 320 428 321 429 
<< pdiffusion >>
rect 321 428 322 429 
<< pdiffusion >>
rect 322 428 323 429 
<< pdiffusion >>
rect 323 428 324 429 
<< m1 >>
rect 325 428 326 429 
<< m2 >>
rect 326 428 327 429 
<< pdiffusion >>
rect 336 428 337 429 
<< pdiffusion >>
rect 337 428 338 429 
<< pdiffusion >>
rect 338 428 339 429 
<< pdiffusion >>
rect 339 428 340 429 
<< pdiffusion >>
rect 340 428 341 429 
<< pdiffusion >>
rect 341 428 342 429 
<< pdiffusion >>
rect 354 428 355 429 
<< pdiffusion >>
rect 355 428 356 429 
<< pdiffusion >>
rect 356 428 357 429 
<< pdiffusion >>
rect 357 428 358 429 
<< pdiffusion >>
rect 358 428 359 429 
<< pdiffusion >>
rect 359 428 360 429 
<< m1 >>
rect 361 428 362 429 
<< m2 >>
rect 361 428 362 429 
<< pdiffusion >>
rect 372 428 373 429 
<< pdiffusion >>
rect 373 428 374 429 
<< pdiffusion >>
rect 374 428 375 429 
<< pdiffusion >>
rect 375 428 376 429 
<< pdiffusion >>
rect 376 428 377 429 
<< pdiffusion >>
rect 377 428 378 429 
<< m1 >>
rect 379 428 380 429 
<< m2 >>
rect 379 428 380 429 
<< m1 >>
rect 385 428 386 429 
<< pdiffusion >>
rect 390 428 391 429 
<< pdiffusion >>
rect 391 428 392 429 
<< pdiffusion >>
rect 392 428 393 429 
<< pdiffusion >>
rect 393 428 394 429 
<< pdiffusion >>
rect 394 428 395 429 
<< pdiffusion >>
rect 395 428 396 429 
<< m1 >>
rect 397 428 398 429 
<< m2 >>
rect 398 428 399 429 
<< m1 >>
rect 402 428 403 429 
<< m1 >>
rect 406 428 407 429 
<< pdiffusion >>
rect 408 428 409 429 
<< pdiffusion >>
rect 409 428 410 429 
<< pdiffusion >>
rect 410 428 411 429 
<< pdiffusion >>
rect 411 428 412 429 
<< pdiffusion >>
rect 412 428 413 429 
<< pdiffusion >>
rect 413 428 414 429 
<< m1 >>
rect 420 428 421 429 
<< m1 >>
rect 424 428 425 429 
<< pdiffusion >>
rect 426 428 427 429 
<< pdiffusion >>
rect 427 428 428 429 
<< pdiffusion >>
rect 428 428 429 429 
<< pdiffusion >>
rect 429 428 430 429 
<< pdiffusion >>
rect 430 428 431 429 
<< pdiffusion >>
rect 431 428 432 429 
<< m1 >>
rect 433 428 434 429 
<< m2 >>
rect 434 428 435 429 
<< m1 >>
rect 442 428 443 429 
<< pdiffusion >>
rect 444 428 445 429 
<< pdiffusion >>
rect 445 428 446 429 
<< pdiffusion >>
rect 446 428 447 429 
<< pdiffusion >>
rect 447 428 448 429 
<< pdiffusion >>
rect 448 428 449 429 
<< pdiffusion >>
rect 449 428 450 429 
<< m1 >>
rect 452 428 453 429 
<< pdiffusion >>
rect 462 428 463 429 
<< pdiffusion >>
rect 463 428 464 429 
<< pdiffusion >>
rect 464 428 465 429 
<< pdiffusion >>
rect 465 428 466 429 
<< pdiffusion >>
rect 466 428 467 429 
<< pdiffusion >>
rect 467 428 468 429 
<< m1 >>
rect 472 428 473 429 
<< m2 >>
rect 473 428 474 429 
<< m1 >>
rect 474 428 475 429 
<< m1 >>
rect 478 428 479 429 
<< pdiffusion >>
rect 480 428 481 429 
<< pdiffusion >>
rect 481 428 482 429 
<< pdiffusion >>
rect 482 428 483 429 
<< pdiffusion >>
rect 483 428 484 429 
<< pdiffusion >>
rect 484 428 485 429 
<< pdiffusion >>
rect 485 428 486 429 
<< m1 >>
rect 487 428 488 429 
<< m1 >>
rect 489 428 490 429 
<< m1 >>
rect 491 428 492 429 
<< pdiffusion >>
rect 498 428 499 429 
<< pdiffusion >>
rect 499 428 500 429 
<< pdiffusion >>
rect 500 428 501 429 
<< pdiffusion >>
rect 501 428 502 429 
<< pdiffusion >>
rect 502 428 503 429 
<< pdiffusion >>
rect 503 428 504 429 
<< pdiffusion >>
rect 516 428 517 429 
<< pdiffusion >>
rect 517 428 518 429 
<< pdiffusion >>
rect 518 428 519 429 
<< pdiffusion >>
rect 519 428 520 429 
<< pdiffusion >>
rect 520 428 521 429 
<< pdiffusion >>
rect 521 428 522 429 
<< pdiffusion >>
rect 12 429 13 430 
<< pdiffusion >>
rect 13 429 14 430 
<< pdiffusion >>
rect 14 429 15 430 
<< pdiffusion >>
rect 15 429 16 430 
<< pdiffusion >>
rect 16 429 17 430 
<< pdiffusion >>
rect 17 429 18 430 
<< m1 >>
rect 19 429 20 430 
<< m1 >>
rect 21 429 22 430 
<< m1 >>
rect 26 429 27 430 
<< m1 >>
rect 28 429 29 430 
<< m2 >>
rect 28 429 29 430 
<< pdiffusion >>
rect 30 429 31 430 
<< pdiffusion >>
rect 31 429 32 430 
<< pdiffusion >>
rect 32 429 33 430 
<< pdiffusion >>
rect 33 429 34 430 
<< pdiffusion >>
rect 34 429 35 430 
<< pdiffusion >>
rect 35 429 36 430 
<< pdiffusion >>
rect 48 429 49 430 
<< pdiffusion >>
rect 49 429 50 430 
<< pdiffusion >>
rect 50 429 51 430 
<< pdiffusion >>
rect 51 429 52 430 
<< pdiffusion >>
rect 52 429 53 430 
<< pdiffusion >>
rect 53 429 54 430 
<< m1 >>
rect 55 429 56 430 
<< pdiffusion >>
rect 66 429 67 430 
<< pdiffusion >>
rect 67 429 68 430 
<< pdiffusion >>
rect 68 429 69 430 
<< pdiffusion >>
rect 69 429 70 430 
<< pdiffusion >>
rect 70 429 71 430 
<< pdiffusion >>
rect 71 429 72 430 
<< m1 >>
rect 73 429 74 430 
<< m1 >>
rect 82 429 83 430 
<< pdiffusion >>
rect 84 429 85 430 
<< pdiffusion >>
rect 85 429 86 430 
<< pdiffusion >>
rect 86 429 87 430 
<< pdiffusion >>
rect 87 429 88 430 
<< pdiffusion >>
rect 88 429 89 430 
<< pdiffusion >>
rect 89 429 90 430 
<< m1 >>
rect 93 429 94 430 
<< m1 >>
rect 96 429 97 430 
<< m1 >>
rect 100 429 101 430 
<< pdiffusion >>
rect 102 429 103 430 
<< pdiffusion >>
rect 103 429 104 430 
<< pdiffusion >>
rect 104 429 105 430 
<< pdiffusion >>
rect 105 429 106 430 
<< pdiffusion >>
rect 106 429 107 430 
<< pdiffusion >>
rect 107 429 108 430 
<< m1 >>
rect 110 429 111 430 
<< m1 >>
rect 114 429 115 430 
<< m1 >>
rect 118 429 119 430 
<< pdiffusion >>
rect 120 429 121 430 
<< pdiffusion >>
rect 121 429 122 430 
<< pdiffusion >>
rect 122 429 123 430 
<< pdiffusion >>
rect 123 429 124 430 
<< pdiffusion >>
rect 124 429 125 430 
<< pdiffusion >>
rect 125 429 126 430 
<< pdiffusion >>
rect 138 429 139 430 
<< pdiffusion >>
rect 139 429 140 430 
<< pdiffusion >>
rect 140 429 141 430 
<< pdiffusion >>
rect 141 429 142 430 
<< pdiffusion >>
rect 142 429 143 430 
<< pdiffusion >>
rect 143 429 144 430 
<< m1 >>
rect 145 429 146 430 
<< m2 >>
rect 145 429 146 430 
<< m1 >>
rect 150 429 151 430 
<< pdiffusion >>
rect 156 429 157 430 
<< pdiffusion >>
rect 157 429 158 430 
<< pdiffusion >>
rect 158 429 159 430 
<< pdiffusion >>
rect 159 429 160 430 
<< pdiffusion >>
rect 160 429 161 430 
<< pdiffusion >>
rect 161 429 162 430 
<< m2 >>
rect 168 429 169 430 
<< m1 >>
rect 169 429 170 430 
<< m1 >>
rect 171 429 172 430 
<< pdiffusion >>
rect 174 429 175 430 
<< pdiffusion >>
rect 175 429 176 430 
<< pdiffusion >>
rect 176 429 177 430 
<< pdiffusion >>
rect 177 429 178 430 
<< pdiffusion >>
rect 178 429 179 430 
<< pdiffusion >>
rect 179 429 180 430 
<< pdiffusion >>
rect 192 429 193 430 
<< pdiffusion >>
rect 193 429 194 430 
<< pdiffusion >>
rect 194 429 195 430 
<< pdiffusion >>
rect 195 429 196 430 
<< pdiffusion >>
rect 196 429 197 430 
<< pdiffusion >>
rect 197 429 198 430 
<< m1 >>
rect 208 429 209 430 
<< pdiffusion >>
rect 210 429 211 430 
<< pdiffusion >>
rect 211 429 212 430 
<< pdiffusion >>
rect 212 429 213 430 
<< pdiffusion >>
rect 213 429 214 430 
<< pdiffusion >>
rect 214 429 215 430 
<< pdiffusion >>
rect 215 429 216 430 
<< m1 >>
rect 217 429 218 430 
<< pdiffusion >>
rect 228 429 229 430 
<< pdiffusion >>
rect 229 429 230 430 
<< pdiffusion >>
rect 230 429 231 430 
<< pdiffusion >>
rect 231 429 232 430 
<< pdiffusion >>
rect 232 429 233 430 
<< pdiffusion >>
rect 233 429 234 430 
<< pdiffusion >>
rect 246 429 247 430 
<< pdiffusion >>
rect 247 429 248 430 
<< pdiffusion >>
rect 248 429 249 430 
<< pdiffusion >>
rect 249 429 250 430 
<< pdiffusion >>
rect 250 429 251 430 
<< pdiffusion >>
rect 251 429 252 430 
<< m1 >>
rect 253 429 254 430 
<< m2 >>
rect 254 429 255 430 
<< pdiffusion >>
rect 264 429 265 430 
<< pdiffusion >>
rect 265 429 266 430 
<< pdiffusion >>
rect 266 429 267 430 
<< pdiffusion >>
rect 267 429 268 430 
<< pdiffusion >>
rect 268 429 269 430 
<< pdiffusion >>
rect 269 429 270 430 
<< pdiffusion >>
rect 282 429 283 430 
<< pdiffusion >>
rect 283 429 284 430 
<< pdiffusion >>
rect 284 429 285 430 
<< pdiffusion >>
rect 285 429 286 430 
<< pdiffusion >>
rect 286 429 287 430 
<< pdiffusion >>
rect 287 429 288 430 
<< m1 >>
rect 290 429 291 430 
<< m1 >>
rect 298 429 299 430 
<< m2 >>
rect 298 429 299 430 
<< pdiffusion >>
rect 300 429 301 430 
<< pdiffusion >>
rect 301 429 302 430 
<< pdiffusion >>
rect 302 429 303 430 
<< pdiffusion >>
rect 303 429 304 430 
<< pdiffusion >>
rect 304 429 305 430 
<< pdiffusion >>
rect 305 429 306 430 
<< m1 >>
rect 307 429 308 430 
<< m1 >>
rect 309 429 310 430 
<< pdiffusion >>
rect 318 429 319 430 
<< pdiffusion >>
rect 319 429 320 430 
<< pdiffusion >>
rect 320 429 321 430 
<< pdiffusion >>
rect 321 429 322 430 
<< pdiffusion >>
rect 322 429 323 430 
<< pdiffusion >>
rect 323 429 324 430 
<< m1 >>
rect 325 429 326 430 
<< m2 >>
rect 326 429 327 430 
<< pdiffusion >>
rect 336 429 337 430 
<< pdiffusion >>
rect 337 429 338 430 
<< pdiffusion >>
rect 338 429 339 430 
<< pdiffusion >>
rect 339 429 340 430 
<< pdiffusion >>
rect 340 429 341 430 
<< pdiffusion >>
rect 341 429 342 430 
<< pdiffusion >>
rect 354 429 355 430 
<< pdiffusion >>
rect 355 429 356 430 
<< pdiffusion >>
rect 356 429 357 430 
<< pdiffusion >>
rect 357 429 358 430 
<< pdiffusion >>
rect 358 429 359 430 
<< pdiffusion >>
rect 359 429 360 430 
<< m1 >>
rect 361 429 362 430 
<< m2 >>
rect 361 429 362 430 
<< pdiffusion >>
rect 372 429 373 430 
<< pdiffusion >>
rect 373 429 374 430 
<< pdiffusion >>
rect 374 429 375 430 
<< pdiffusion >>
rect 375 429 376 430 
<< pdiffusion >>
rect 376 429 377 430 
<< pdiffusion >>
rect 377 429 378 430 
<< m1 >>
rect 379 429 380 430 
<< m2 >>
rect 379 429 380 430 
<< m1 >>
rect 385 429 386 430 
<< pdiffusion >>
rect 390 429 391 430 
<< pdiffusion >>
rect 391 429 392 430 
<< pdiffusion >>
rect 392 429 393 430 
<< pdiffusion >>
rect 393 429 394 430 
<< pdiffusion >>
rect 394 429 395 430 
<< pdiffusion >>
rect 395 429 396 430 
<< m1 >>
rect 397 429 398 430 
<< m2 >>
rect 398 429 399 430 
<< m1 >>
rect 402 429 403 430 
<< m1 >>
rect 406 429 407 430 
<< pdiffusion >>
rect 408 429 409 430 
<< pdiffusion >>
rect 409 429 410 430 
<< pdiffusion >>
rect 410 429 411 430 
<< pdiffusion >>
rect 411 429 412 430 
<< pdiffusion >>
rect 412 429 413 430 
<< pdiffusion >>
rect 413 429 414 430 
<< m1 >>
rect 420 429 421 430 
<< m1 >>
rect 424 429 425 430 
<< pdiffusion >>
rect 426 429 427 430 
<< pdiffusion >>
rect 427 429 428 430 
<< pdiffusion >>
rect 428 429 429 430 
<< pdiffusion >>
rect 429 429 430 430 
<< pdiffusion >>
rect 430 429 431 430 
<< pdiffusion >>
rect 431 429 432 430 
<< m1 >>
rect 433 429 434 430 
<< m2 >>
rect 434 429 435 430 
<< m1 >>
rect 442 429 443 430 
<< pdiffusion >>
rect 444 429 445 430 
<< pdiffusion >>
rect 445 429 446 430 
<< pdiffusion >>
rect 446 429 447 430 
<< pdiffusion >>
rect 447 429 448 430 
<< pdiffusion >>
rect 448 429 449 430 
<< pdiffusion >>
rect 449 429 450 430 
<< m1 >>
rect 452 429 453 430 
<< pdiffusion >>
rect 462 429 463 430 
<< pdiffusion >>
rect 463 429 464 430 
<< pdiffusion >>
rect 464 429 465 430 
<< pdiffusion >>
rect 465 429 466 430 
<< pdiffusion >>
rect 466 429 467 430 
<< pdiffusion >>
rect 467 429 468 430 
<< m1 >>
rect 472 429 473 430 
<< m2 >>
rect 473 429 474 430 
<< m1 >>
rect 474 429 475 430 
<< m1 >>
rect 478 429 479 430 
<< pdiffusion >>
rect 480 429 481 430 
<< pdiffusion >>
rect 481 429 482 430 
<< pdiffusion >>
rect 482 429 483 430 
<< pdiffusion >>
rect 483 429 484 430 
<< pdiffusion >>
rect 484 429 485 430 
<< pdiffusion >>
rect 485 429 486 430 
<< m1 >>
rect 487 429 488 430 
<< m1 >>
rect 489 429 490 430 
<< m1 >>
rect 491 429 492 430 
<< pdiffusion >>
rect 498 429 499 430 
<< pdiffusion >>
rect 499 429 500 430 
<< pdiffusion >>
rect 500 429 501 430 
<< pdiffusion >>
rect 501 429 502 430 
<< pdiffusion >>
rect 502 429 503 430 
<< pdiffusion >>
rect 503 429 504 430 
<< pdiffusion >>
rect 516 429 517 430 
<< pdiffusion >>
rect 517 429 518 430 
<< pdiffusion >>
rect 518 429 519 430 
<< pdiffusion >>
rect 519 429 520 430 
<< pdiffusion >>
rect 520 429 521 430 
<< pdiffusion >>
rect 521 429 522 430 
<< pdiffusion >>
rect 12 430 13 431 
<< pdiffusion >>
rect 13 430 14 431 
<< pdiffusion >>
rect 14 430 15 431 
<< pdiffusion >>
rect 15 430 16 431 
<< pdiffusion >>
rect 16 430 17 431 
<< pdiffusion >>
rect 17 430 18 431 
<< m1 >>
rect 19 430 20 431 
<< m1 >>
rect 21 430 22 431 
<< m1 >>
rect 26 430 27 431 
<< m1 >>
rect 28 430 29 431 
<< m2 >>
rect 28 430 29 431 
<< pdiffusion >>
rect 30 430 31 431 
<< pdiffusion >>
rect 31 430 32 431 
<< pdiffusion >>
rect 32 430 33 431 
<< pdiffusion >>
rect 33 430 34 431 
<< pdiffusion >>
rect 34 430 35 431 
<< pdiffusion >>
rect 35 430 36 431 
<< pdiffusion >>
rect 48 430 49 431 
<< pdiffusion >>
rect 49 430 50 431 
<< pdiffusion >>
rect 50 430 51 431 
<< pdiffusion >>
rect 51 430 52 431 
<< pdiffusion >>
rect 52 430 53 431 
<< pdiffusion >>
rect 53 430 54 431 
<< m1 >>
rect 55 430 56 431 
<< pdiffusion >>
rect 66 430 67 431 
<< pdiffusion >>
rect 67 430 68 431 
<< pdiffusion >>
rect 68 430 69 431 
<< pdiffusion >>
rect 69 430 70 431 
<< pdiffusion >>
rect 70 430 71 431 
<< pdiffusion >>
rect 71 430 72 431 
<< m1 >>
rect 73 430 74 431 
<< m1 >>
rect 82 430 83 431 
<< pdiffusion >>
rect 84 430 85 431 
<< pdiffusion >>
rect 85 430 86 431 
<< pdiffusion >>
rect 86 430 87 431 
<< pdiffusion >>
rect 87 430 88 431 
<< pdiffusion >>
rect 88 430 89 431 
<< pdiffusion >>
rect 89 430 90 431 
<< m1 >>
rect 93 430 94 431 
<< m1 >>
rect 96 430 97 431 
<< m1 >>
rect 100 430 101 431 
<< pdiffusion >>
rect 102 430 103 431 
<< pdiffusion >>
rect 103 430 104 431 
<< pdiffusion >>
rect 104 430 105 431 
<< pdiffusion >>
rect 105 430 106 431 
<< pdiffusion >>
rect 106 430 107 431 
<< pdiffusion >>
rect 107 430 108 431 
<< m1 >>
rect 110 430 111 431 
<< m1 >>
rect 114 430 115 431 
<< m1 >>
rect 118 430 119 431 
<< pdiffusion >>
rect 120 430 121 431 
<< pdiffusion >>
rect 121 430 122 431 
<< pdiffusion >>
rect 122 430 123 431 
<< pdiffusion >>
rect 123 430 124 431 
<< pdiffusion >>
rect 124 430 125 431 
<< pdiffusion >>
rect 125 430 126 431 
<< pdiffusion >>
rect 138 430 139 431 
<< pdiffusion >>
rect 139 430 140 431 
<< pdiffusion >>
rect 140 430 141 431 
<< pdiffusion >>
rect 141 430 142 431 
<< pdiffusion >>
rect 142 430 143 431 
<< pdiffusion >>
rect 143 430 144 431 
<< m1 >>
rect 145 430 146 431 
<< m2 >>
rect 145 430 146 431 
<< m1 >>
rect 150 430 151 431 
<< pdiffusion >>
rect 156 430 157 431 
<< pdiffusion >>
rect 157 430 158 431 
<< pdiffusion >>
rect 158 430 159 431 
<< pdiffusion >>
rect 159 430 160 431 
<< pdiffusion >>
rect 160 430 161 431 
<< pdiffusion >>
rect 161 430 162 431 
<< m2 >>
rect 168 430 169 431 
<< m1 >>
rect 169 430 170 431 
<< m1 >>
rect 171 430 172 431 
<< pdiffusion >>
rect 174 430 175 431 
<< pdiffusion >>
rect 175 430 176 431 
<< pdiffusion >>
rect 176 430 177 431 
<< pdiffusion >>
rect 177 430 178 431 
<< pdiffusion >>
rect 178 430 179 431 
<< pdiffusion >>
rect 179 430 180 431 
<< pdiffusion >>
rect 192 430 193 431 
<< pdiffusion >>
rect 193 430 194 431 
<< pdiffusion >>
rect 194 430 195 431 
<< pdiffusion >>
rect 195 430 196 431 
<< pdiffusion >>
rect 196 430 197 431 
<< pdiffusion >>
rect 197 430 198 431 
<< m1 >>
rect 208 430 209 431 
<< pdiffusion >>
rect 210 430 211 431 
<< pdiffusion >>
rect 211 430 212 431 
<< pdiffusion >>
rect 212 430 213 431 
<< pdiffusion >>
rect 213 430 214 431 
<< pdiffusion >>
rect 214 430 215 431 
<< pdiffusion >>
rect 215 430 216 431 
<< m1 >>
rect 217 430 218 431 
<< pdiffusion >>
rect 228 430 229 431 
<< pdiffusion >>
rect 229 430 230 431 
<< pdiffusion >>
rect 230 430 231 431 
<< pdiffusion >>
rect 231 430 232 431 
<< pdiffusion >>
rect 232 430 233 431 
<< pdiffusion >>
rect 233 430 234 431 
<< pdiffusion >>
rect 246 430 247 431 
<< pdiffusion >>
rect 247 430 248 431 
<< pdiffusion >>
rect 248 430 249 431 
<< pdiffusion >>
rect 249 430 250 431 
<< pdiffusion >>
rect 250 430 251 431 
<< pdiffusion >>
rect 251 430 252 431 
<< m1 >>
rect 253 430 254 431 
<< m2 >>
rect 254 430 255 431 
<< pdiffusion >>
rect 264 430 265 431 
<< pdiffusion >>
rect 265 430 266 431 
<< pdiffusion >>
rect 266 430 267 431 
<< pdiffusion >>
rect 267 430 268 431 
<< pdiffusion >>
rect 268 430 269 431 
<< pdiffusion >>
rect 269 430 270 431 
<< pdiffusion >>
rect 282 430 283 431 
<< pdiffusion >>
rect 283 430 284 431 
<< pdiffusion >>
rect 284 430 285 431 
<< pdiffusion >>
rect 285 430 286 431 
<< pdiffusion >>
rect 286 430 287 431 
<< pdiffusion >>
rect 287 430 288 431 
<< m1 >>
rect 290 430 291 431 
<< m1 >>
rect 298 430 299 431 
<< m2 >>
rect 298 430 299 431 
<< pdiffusion >>
rect 300 430 301 431 
<< pdiffusion >>
rect 301 430 302 431 
<< pdiffusion >>
rect 302 430 303 431 
<< pdiffusion >>
rect 303 430 304 431 
<< pdiffusion >>
rect 304 430 305 431 
<< pdiffusion >>
rect 305 430 306 431 
<< m1 >>
rect 307 430 308 431 
<< m1 >>
rect 309 430 310 431 
<< pdiffusion >>
rect 318 430 319 431 
<< pdiffusion >>
rect 319 430 320 431 
<< pdiffusion >>
rect 320 430 321 431 
<< pdiffusion >>
rect 321 430 322 431 
<< pdiffusion >>
rect 322 430 323 431 
<< pdiffusion >>
rect 323 430 324 431 
<< m1 >>
rect 325 430 326 431 
<< m2 >>
rect 326 430 327 431 
<< pdiffusion >>
rect 336 430 337 431 
<< pdiffusion >>
rect 337 430 338 431 
<< pdiffusion >>
rect 338 430 339 431 
<< pdiffusion >>
rect 339 430 340 431 
<< pdiffusion >>
rect 340 430 341 431 
<< pdiffusion >>
rect 341 430 342 431 
<< pdiffusion >>
rect 354 430 355 431 
<< pdiffusion >>
rect 355 430 356 431 
<< pdiffusion >>
rect 356 430 357 431 
<< pdiffusion >>
rect 357 430 358 431 
<< pdiffusion >>
rect 358 430 359 431 
<< pdiffusion >>
rect 359 430 360 431 
<< m1 >>
rect 361 430 362 431 
<< m2 >>
rect 361 430 362 431 
<< pdiffusion >>
rect 372 430 373 431 
<< pdiffusion >>
rect 373 430 374 431 
<< pdiffusion >>
rect 374 430 375 431 
<< pdiffusion >>
rect 375 430 376 431 
<< pdiffusion >>
rect 376 430 377 431 
<< pdiffusion >>
rect 377 430 378 431 
<< m1 >>
rect 379 430 380 431 
<< m2 >>
rect 379 430 380 431 
<< m1 >>
rect 385 430 386 431 
<< pdiffusion >>
rect 390 430 391 431 
<< pdiffusion >>
rect 391 430 392 431 
<< pdiffusion >>
rect 392 430 393 431 
<< pdiffusion >>
rect 393 430 394 431 
<< pdiffusion >>
rect 394 430 395 431 
<< pdiffusion >>
rect 395 430 396 431 
<< m1 >>
rect 397 430 398 431 
<< m2 >>
rect 398 430 399 431 
<< m1 >>
rect 402 430 403 431 
<< m1 >>
rect 406 430 407 431 
<< pdiffusion >>
rect 408 430 409 431 
<< pdiffusion >>
rect 409 430 410 431 
<< pdiffusion >>
rect 410 430 411 431 
<< pdiffusion >>
rect 411 430 412 431 
<< pdiffusion >>
rect 412 430 413 431 
<< pdiffusion >>
rect 413 430 414 431 
<< m1 >>
rect 420 430 421 431 
<< m1 >>
rect 424 430 425 431 
<< pdiffusion >>
rect 426 430 427 431 
<< pdiffusion >>
rect 427 430 428 431 
<< pdiffusion >>
rect 428 430 429 431 
<< pdiffusion >>
rect 429 430 430 431 
<< pdiffusion >>
rect 430 430 431 431 
<< pdiffusion >>
rect 431 430 432 431 
<< m1 >>
rect 433 430 434 431 
<< m2 >>
rect 434 430 435 431 
<< m1 >>
rect 442 430 443 431 
<< pdiffusion >>
rect 444 430 445 431 
<< pdiffusion >>
rect 445 430 446 431 
<< pdiffusion >>
rect 446 430 447 431 
<< pdiffusion >>
rect 447 430 448 431 
<< pdiffusion >>
rect 448 430 449 431 
<< pdiffusion >>
rect 449 430 450 431 
<< m1 >>
rect 452 430 453 431 
<< pdiffusion >>
rect 462 430 463 431 
<< pdiffusion >>
rect 463 430 464 431 
<< pdiffusion >>
rect 464 430 465 431 
<< pdiffusion >>
rect 465 430 466 431 
<< pdiffusion >>
rect 466 430 467 431 
<< pdiffusion >>
rect 467 430 468 431 
<< m1 >>
rect 472 430 473 431 
<< m2 >>
rect 473 430 474 431 
<< m1 >>
rect 474 430 475 431 
<< m1 >>
rect 478 430 479 431 
<< pdiffusion >>
rect 480 430 481 431 
<< pdiffusion >>
rect 481 430 482 431 
<< pdiffusion >>
rect 482 430 483 431 
<< pdiffusion >>
rect 483 430 484 431 
<< pdiffusion >>
rect 484 430 485 431 
<< pdiffusion >>
rect 485 430 486 431 
<< m1 >>
rect 487 430 488 431 
<< m1 >>
rect 489 430 490 431 
<< m1 >>
rect 491 430 492 431 
<< pdiffusion >>
rect 498 430 499 431 
<< pdiffusion >>
rect 499 430 500 431 
<< pdiffusion >>
rect 500 430 501 431 
<< pdiffusion >>
rect 501 430 502 431 
<< pdiffusion >>
rect 502 430 503 431 
<< pdiffusion >>
rect 503 430 504 431 
<< pdiffusion >>
rect 516 430 517 431 
<< pdiffusion >>
rect 517 430 518 431 
<< pdiffusion >>
rect 518 430 519 431 
<< pdiffusion >>
rect 519 430 520 431 
<< pdiffusion >>
rect 520 430 521 431 
<< pdiffusion >>
rect 521 430 522 431 
<< pdiffusion >>
rect 12 431 13 432 
<< pdiffusion >>
rect 13 431 14 432 
<< pdiffusion >>
rect 14 431 15 432 
<< pdiffusion >>
rect 15 431 16 432 
<< pdiffusion >>
rect 16 431 17 432 
<< pdiffusion >>
rect 17 431 18 432 
<< m1 >>
rect 19 431 20 432 
<< m1 >>
rect 21 431 22 432 
<< m1 >>
rect 26 431 27 432 
<< m1 >>
rect 28 431 29 432 
<< m2 >>
rect 28 431 29 432 
<< pdiffusion >>
rect 30 431 31 432 
<< pdiffusion >>
rect 31 431 32 432 
<< pdiffusion >>
rect 32 431 33 432 
<< pdiffusion >>
rect 33 431 34 432 
<< pdiffusion >>
rect 34 431 35 432 
<< pdiffusion >>
rect 35 431 36 432 
<< pdiffusion >>
rect 48 431 49 432 
<< pdiffusion >>
rect 49 431 50 432 
<< pdiffusion >>
rect 50 431 51 432 
<< pdiffusion >>
rect 51 431 52 432 
<< m1 >>
rect 52 431 53 432 
<< pdiffusion >>
rect 52 431 53 432 
<< pdiffusion >>
rect 53 431 54 432 
<< m1 >>
rect 55 431 56 432 
<< pdiffusion >>
rect 66 431 67 432 
<< pdiffusion >>
rect 67 431 68 432 
<< pdiffusion >>
rect 68 431 69 432 
<< pdiffusion >>
rect 69 431 70 432 
<< pdiffusion >>
rect 70 431 71 432 
<< pdiffusion >>
rect 71 431 72 432 
<< m1 >>
rect 73 431 74 432 
<< m1 >>
rect 82 431 83 432 
<< pdiffusion >>
rect 84 431 85 432 
<< pdiffusion >>
rect 85 431 86 432 
<< pdiffusion >>
rect 86 431 87 432 
<< pdiffusion >>
rect 87 431 88 432 
<< m1 >>
rect 88 431 89 432 
<< pdiffusion >>
rect 88 431 89 432 
<< pdiffusion >>
rect 89 431 90 432 
<< m1 >>
rect 93 431 94 432 
<< m2 >>
rect 93 431 94 432 
<< m2c >>
rect 93 431 94 432 
<< m1 >>
rect 93 431 94 432 
<< m2 >>
rect 93 431 94 432 
<< m1 >>
rect 96 431 97 432 
<< m2 >>
rect 96 431 97 432 
<< m2c >>
rect 96 431 97 432 
<< m1 >>
rect 96 431 97 432 
<< m2 >>
rect 96 431 97 432 
<< m1 >>
rect 100 431 101 432 
<< pdiffusion >>
rect 102 431 103 432 
<< pdiffusion >>
rect 103 431 104 432 
<< pdiffusion >>
rect 104 431 105 432 
<< pdiffusion >>
rect 105 431 106 432 
<< pdiffusion >>
rect 106 431 107 432 
<< pdiffusion >>
rect 107 431 108 432 
<< m1 >>
rect 110 431 111 432 
<< m1 >>
rect 114 431 115 432 
<< m1 >>
rect 118 431 119 432 
<< pdiffusion >>
rect 120 431 121 432 
<< pdiffusion >>
rect 121 431 122 432 
<< pdiffusion >>
rect 122 431 123 432 
<< pdiffusion >>
rect 123 431 124 432 
<< pdiffusion >>
rect 124 431 125 432 
<< pdiffusion >>
rect 125 431 126 432 
<< pdiffusion >>
rect 138 431 139 432 
<< pdiffusion >>
rect 139 431 140 432 
<< pdiffusion >>
rect 140 431 141 432 
<< pdiffusion >>
rect 141 431 142 432 
<< pdiffusion >>
rect 142 431 143 432 
<< pdiffusion >>
rect 143 431 144 432 
<< m1 >>
rect 145 431 146 432 
<< m2 >>
rect 145 431 146 432 
<< m1 >>
rect 150 431 151 432 
<< m2 >>
rect 150 431 151 432 
<< m2c >>
rect 150 431 151 432 
<< m1 >>
rect 150 431 151 432 
<< m2 >>
rect 150 431 151 432 
<< pdiffusion >>
rect 156 431 157 432 
<< m1 >>
rect 157 431 158 432 
<< pdiffusion >>
rect 157 431 158 432 
<< pdiffusion >>
rect 158 431 159 432 
<< pdiffusion >>
rect 159 431 160 432 
<< m1 >>
rect 160 431 161 432 
<< pdiffusion >>
rect 160 431 161 432 
<< pdiffusion >>
rect 161 431 162 432 
<< m1 >>
rect 164 431 165 432 
<< m2 >>
rect 164 431 165 432 
<< m2c >>
rect 164 431 165 432 
<< m1 >>
rect 164 431 165 432 
<< m2 >>
rect 164 431 165 432 
<< m1 >>
rect 165 431 166 432 
<< m1 >>
rect 166 431 167 432 
<< m1 >>
rect 167 431 168 432 
<< m2 >>
rect 167 431 168 432 
<< m2c >>
rect 167 431 168 432 
<< m1 >>
rect 167 431 168 432 
<< m2 >>
rect 167 431 168 432 
<< m2 >>
rect 168 431 169 432 
<< m1 >>
rect 169 431 170 432 
<< m1 >>
rect 171 431 172 432 
<< pdiffusion >>
rect 174 431 175 432 
<< pdiffusion >>
rect 175 431 176 432 
<< pdiffusion >>
rect 176 431 177 432 
<< pdiffusion >>
rect 177 431 178 432 
<< pdiffusion >>
rect 178 431 179 432 
<< pdiffusion >>
rect 179 431 180 432 
<< pdiffusion >>
rect 192 431 193 432 
<< m1 >>
rect 193 431 194 432 
<< pdiffusion >>
rect 193 431 194 432 
<< pdiffusion >>
rect 194 431 195 432 
<< pdiffusion >>
rect 195 431 196 432 
<< pdiffusion >>
rect 196 431 197 432 
<< pdiffusion >>
rect 197 431 198 432 
<< m1 >>
rect 208 431 209 432 
<< pdiffusion >>
rect 210 431 211 432 
<< pdiffusion >>
rect 211 431 212 432 
<< pdiffusion >>
rect 212 431 213 432 
<< pdiffusion >>
rect 213 431 214 432 
<< pdiffusion >>
rect 214 431 215 432 
<< pdiffusion >>
rect 215 431 216 432 
<< m1 >>
rect 217 431 218 432 
<< pdiffusion >>
rect 228 431 229 432 
<< pdiffusion >>
rect 229 431 230 432 
<< pdiffusion >>
rect 230 431 231 432 
<< pdiffusion >>
rect 231 431 232 432 
<< pdiffusion >>
rect 232 431 233 432 
<< pdiffusion >>
rect 233 431 234 432 
<< pdiffusion >>
rect 246 431 247 432 
<< m1 >>
rect 247 431 248 432 
<< pdiffusion >>
rect 247 431 248 432 
<< pdiffusion >>
rect 248 431 249 432 
<< pdiffusion >>
rect 249 431 250 432 
<< pdiffusion >>
rect 250 431 251 432 
<< pdiffusion >>
rect 251 431 252 432 
<< m1 >>
rect 253 431 254 432 
<< m2 >>
rect 254 431 255 432 
<< pdiffusion >>
rect 264 431 265 432 
<< pdiffusion >>
rect 265 431 266 432 
<< pdiffusion >>
rect 266 431 267 432 
<< pdiffusion >>
rect 267 431 268 432 
<< pdiffusion >>
rect 268 431 269 432 
<< pdiffusion >>
rect 269 431 270 432 
<< pdiffusion >>
rect 282 431 283 432 
<< pdiffusion >>
rect 283 431 284 432 
<< pdiffusion >>
rect 284 431 285 432 
<< pdiffusion >>
rect 285 431 286 432 
<< m1 >>
rect 286 431 287 432 
<< pdiffusion >>
rect 286 431 287 432 
<< pdiffusion >>
rect 287 431 288 432 
<< m1 >>
rect 290 431 291 432 
<< m1 >>
rect 298 431 299 432 
<< m2 >>
rect 298 431 299 432 
<< pdiffusion >>
rect 300 431 301 432 
<< m1 >>
rect 301 431 302 432 
<< pdiffusion >>
rect 301 431 302 432 
<< pdiffusion >>
rect 302 431 303 432 
<< pdiffusion >>
rect 303 431 304 432 
<< pdiffusion >>
rect 304 431 305 432 
<< pdiffusion >>
rect 305 431 306 432 
<< m1 >>
rect 307 431 308 432 
<< m1 >>
rect 309 431 310 432 
<< pdiffusion >>
rect 318 431 319 432 
<< pdiffusion >>
rect 319 431 320 432 
<< pdiffusion >>
rect 320 431 321 432 
<< pdiffusion >>
rect 321 431 322 432 
<< m1 >>
rect 322 431 323 432 
<< pdiffusion >>
rect 322 431 323 432 
<< pdiffusion >>
rect 323 431 324 432 
<< m1 >>
rect 325 431 326 432 
<< m2 >>
rect 326 431 327 432 
<< pdiffusion >>
rect 336 431 337 432 
<< pdiffusion >>
rect 337 431 338 432 
<< pdiffusion >>
rect 338 431 339 432 
<< pdiffusion >>
rect 339 431 340 432 
<< m1 >>
rect 340 431 341 432 
<< pdiffusion >>
rect 340 431 341 432 
<< pdiffusion >>
rect 341 431 342 432 
<< pdiffusion >>
rect 354 431 355 432 
<< pdiffusion >>
rect 355 431 356 432 
<< pdiffusion >>
rect 356 431 357 432 
<< pdiffusion >>
rect 357 431 358 432 
<< m1 >>
rect 358 431 359 432 
<< pdiffusion >>
rect 358 431 359 432 
<< pdiffusion >>
rect 359 431 360 432 
<< m1 >>
rect 361 431 362 432 
<< m2 >>
rect 361 431 362 432 
<< pdiffusion >>
rect 372 431 373 432 
<< m1 >>
rect 373 431 374 432 
<< pdiffusion >>
rect 373 431 374 432 
<< pdiffusion >>
rect 374 431 375 432 
<< pdiffusion >>
rect 375 431 376 432 
<< pdiffusion >>
rect 376 431 377 432 
<< pdiffusion >>
rect 377 431 378 432 
<< m1 >>
rect 379 431 380 432 
<< m2 >>
rect 379 431 380 432 
<< m1 >>
rect 385 431 386 432 
<< m2 >>
rect 385 431 386 432 
<< m2c >>
rect 385 431 386 432 
<< m1 >>
rect 385 431 386 432 
<< m2 >>
rect 385 431 386 432 
<< pdiffusion >>
rect 390 431 391 432 
<< m1 >>
rect 391 431 392 432 
<< pdiffusion >>
rect 391 431 392 432 
<< pdiffusion >>
rect 392 431 393 432 
<< pdiffusion >>
rect 393 431 394 432 
<< pdiffusion >>
rect 394 431 395 432 
<< pdiffusion >>
rect 395 431 396 432 
<< m1 >>
rect 397 431 398 432 
<< m2 >>
rect 398 431 399 432 
<< m1 >>
rect 402 431 403 432 
<< m1 >>
rect 406 431 407 432 
<< pdiffusion >>
rect 408 431 409 432 
<< pdiffusion >>
rect 409 431 410 432 
<< pdiffusion >>
rect 410 431 411 432 
<< pdiffusion >>
rect 411 431 412 432 
<< pdiffusion >>
rect 412 431 413 432 
<< pdiffusion >>
rect 413 431 414 432 
<< m1 >>
rect 420 431 421 432 
<< m1 >>
rect 424 431 425 432 
<< pdiffusion >>
rect 426 431 427 432 
<< pdiffusion >>
rect 427 431 428 432 
<< pdiffusion >>
rect 428 431 429 432 
<< pdiffusion >>
rect 429 431 430 432 
<< m1 >>
rect 430 431 431 432 
<< pdiffusion >>
rect 430 431 431 432 
<< pdiffusion >>
rect 431 431 432 432 
<< m1 >>
rect 433 431 434 432 
<< m2 >>
rect 434 431 435 432 
<< m1 >>
rect 442 431 443 432 
<< pdiffusion >>
rect 444 431 445 432 
<< pdiffusion >>
rect 445 431 446 432 
<< pdiffusion >>
rect 446 431 447 432 
<< pdiffusion >>
rect 447 431 448 432 
<< m1 >>
rect 448 431 449 432 
<< pdiffusion >>
rect 448 431 449 432 
<< pdiffusion >>
rect 449 431 450 432 
<< m1 >>
rect 452 431 453 432 
<< pdiffusion >>
rect 462 431 463 432 
<< pdiffusion >>
rect 463 431 464 432 
<< pdiffusion >>
rect 464 431 465 432 
<< pdiffusion >>
rect 465 431 466 432 
<< pdiffusion >>
rect 466 431 467 432 
<< pdiffusion >>
rect 467 431 468 432 
<< m1 >>
rect 472 431 473 432 
<< m2 >>
rect 473 431 474 432 
<< m1 >>
rect 474 431 475 432 
<< m1 >>
rect 478 431 479 432 
<< pdiffusion >>
rect 480 431 481 432 
<< pdiffusion >>
rect 481 431 482 432 
<< pdiffusion >>
rect 482 431 483 432 
<< pdiffusion >>
rect 483 431 484 432 
<< pdiffusion >>
rect 484 431 485 432 
<< pdiffusion >>
rect 485 431 486 432 
<< m1 >>
rect 487 431 488 432 
<< m1 >>
rect 489 431 490 432 
<< m1 >>
rect 491 431 492 432 
<< pdiffusion >>
rect 498 431 499 432 
<< pdiffusion >>
rect 499 431 500 432 
<< pdiffusion >>
rect 500 431 501 432 
<< pdiffusion >>
rect 501 431 502 432 
<< pdiffusion >>
rect 502 431 503 432 
<< pdiffusion >>
rect 503 431 504 432 
<< pdiffusion >>
rect 516 431 517 432 
<< pdiffusion >>
rect 517 431 518 432 
<< pdiffusion >>
rect 518 431 519 432 
<< pdiffusion >>
rect 519 431 520 432 
<< m1 >>
rect 520 431 521 432 
<< pdiffusion >>
rect 520 431 521 432 
<< pdiffusion >>
rect 521 431 522 432 
<< m1 >>
rect 19 432 20 433 
<< m1 >>
rect 21 432 22 433 
<< m1 >>
rect 26 432 27 433 
<< m1 >>
rect 28 432 29 433 
<< m2 >>
rect 28 432 29 433 
<< m1 >>
rect 52 432 53 433 
<< m1 >>
rect 55 432 56 433 
<< m1 >>
rect 73 432 74 433 
<< m1 >>
rect 82 432 83 433 
<< m1 >>
rect 88 432 89 433 
<< m2 >>
rect 93 432 94 433 
<< m2 >>
rect 96 432 97 433 
<< m1 >>
rect 100 432 101 433 
<< m1 >>
rect 110 432 111 433 
<< m2 >>
rect 110 432 111 433 
<< m2c >>
rect 110 432 111 433 
<< m1 >>
rect 110 432 111 433 
<< m2 >>
rect 110 432 111 433 
<< m1 >>
rect 114 432 115 433 
<< m2 >>
rect 114 432 115 433 
<< m2c >>
rect 114 432 115 433 
<< m1 >>
rect 114 432 115 433 
<< m2 >>
rect 114 432 115 433 
<< m1 >>
rect 118 432 119 433 
<< m1 >>
rect 145 432 146 433 
<< m2 >>
rect 145 432 146 433 
<< m2 >>
rect 150 432 151 433 
<< m1 >>
rect 157 432 158 433 
<< m1 >>
rect 160 432 161 433 
<< m2 >>
rect 164 432 165 433 
<< m1 >>
rect 169 432 170 433 
<< m1 >>
rect 171 432 172 433 
<< m1 >>
rect 193 432 194 433 
<< m1 >>
rect 208 432 209 433 
<< m1 >>
rect 217 432 218 433 
<< m1 >>
rect 247 432 248 433 
<< m1 >>
rect 253 432 254 433 
<< m2 >>
rect 254 432 255 433 
<< m1 >>
rect 286 432 287 433 
<< m1 >>
rect 290 432 291 433 
<< m1 >>
rect 298 432 299 433 
<< m2 >>
rect 298 432 299 433 
<< m1 >>
rect 301 432 302 433 
<< m1 >>
rect 307 432 308 433 
<< m1 >>
rect 309 432 310 433 
<< m1 >>
rect 322 432 323 433 
<< m1 >>
rect 325 432 326 433 
<< m2 >>
rect 326 432 327 433 
<< m1 >>
rect 340 432 341 433 
<< m1 >>
rect 358 432 359 433 
<< m1 >>
rect 361 432 362 433 
<< m2 >>
rect 361 432 362 433 
<< m1 >>
rect 373 432 374 433 
<< m1 >>
rect 379 432 380 433 
<< m2 >>
rect 379 432 380 433 
<< m2 >>
rect 385 432 386 433 
<< m1 >>
rect 391 432 392 433 
<< m1 >>
rect 397 432 398 433 
<< m2 >>
rect 398 432 399 433 
<< m1 >>
rect 402 432 403 433 
<< m1 >>
rect 406 432 407 433 
<< m1 >>
rect 420 432 421 433 
<< m1 >>
rect 424 432 425 433 
<< m1 >>
rect 430 432 431 433 
<< m1 >>
rect 433 432 434 433 
<< m2 >>
rect 434 432 435 433 
<< m1 >>
rect 442 432 443 433 
<< m1 >>
rect 448 432 449 433 
<< m1 >>
rect 452 432 453 433 
<< m1 >>
rect 472 432 473 433 
<< m2 >>
rect 473 432 474 433 
<< m1 >>
rect 474 432 475 433 
<< m1 >>
rect 478 432 479 433 
<< m1 >>
rect 487 432 488 433 
<< m1 >>
rect 489 432 490 433 
<< m1 >>
rect 491 432 492 433 
<< m1 >>
rect 520 432 521 433 
<< m1 >>
rect 19 433 20 434 
<< m1 >>
rect 21 433 22 434 
<< m1 >>
rect 26 433 27 434 
<< m1 >>
rect 28 433 29 434 
<< m2 >>
rect 28 433 29 434 
<< m1 >>
rect 52 433 53 434 
<< m1 >>
rect 53 433 54 434 
<< m1 >>
rect 54 433 55 434 
<< m1 >>
rect 55 433 56 434 
<< m1 >>
rect 73 433 74 434 
<< m1 >>
rect 82 433 83 434 
<< m1 >>
rect 88 433 89 434 
<< m1 >>
rect 89 433 90 434 
<< m1 >>
rect 90 433 91 434 
<< m1 >>
rect 91 433 92 434 
<< m1 >>
rect 92 433 93 434 
<< m1 >>
rect 93 433 94 434 
<< m2 >>
rect 93 433 94 434 
<< m1 >>
rect 94 433 95 434 
<< m1 >>
rect 95 433 96 434 
<< m1 >>
rect 96 433 97 434 
<< m2 >>
rect 96 433 97 434 
<< m1 >>
rect 97 433 98 434 
<< m1 >>
rect 98 433 99 434 
<< m2 >>
rect 98 433 99 434 
<< m2c >>
rect 98 433 99 434 
<< m1 >>
rect 98 433 99 434 
<< m2 >>
rect 98 433 99 434 
<< m2 >>
rect 99 433 100 434 
<< m1 >>
rect 100 433 101 434 
<< m2 >>
rect 100 433 101 434 
<< m2 >>
rect 101 433 102 434 
<< m1 >>
rect 102 433 103 434 
<< m2 >>
rect 102 433 103 434 
<< m2c >>
rect 102 433 103 434 
<< m1 >>
rect 102 433 103 434 
<< m2 >>
rect 102 433 103 434 
<< m2 >>
rect 110 433 111 434 
<< m2 >>
rect 114 433 115 434 
<< m1 >>
rect 118 433 119 434 
<< m1 >>
rect 145 433 146 434 
<< m2 >>
rect 145 433 146 434 
<< m1 >>
rect 146 433 147 434 
<< m1 >>
rect 147 433 148 434 
<< m1 >>
rect 148 433 149 434 
<< m1 >>
rect 149 433 150 434 
<< m1 >>
rect 150 433 151 434 
<< m2 >>
rect 150 433 151 434 
<< m1 >>
rect 151 433 152 434 
<< m1 >>
rect 152 433 153 434 
<< m1 >>
rect 153 433 154 434 
<< m1 >>
rect 154 433 155 434 
<< m1 >>
rect 155 433 156 434 
<< m1 >>
rect 156 433 157 434 
<< m1 >>
rect 157 433 158 434 
<< m1 >>
rect 160 433 161 434 
<< m2 >>
rect 161 433 162 434 
<< m1 >>
rect 162 433 163 434 
<< m2 >>
rect 162 433 163 434 
<< m2c >>
rect 162 433 163 434 
<< m1 >>
rect 162 433 163 434 
<< m2 >>
rect 162 433 163 434 
<< m1 >>
rect 163 433 164 434 
<< m1 >>
rect 164 433 165 434 
<< m2 >>
rect 164 433 165 434 
<< m1 >>
rect 165 433 166 434 
<< m1 >>
rect 166 433 167 434 
<< m1 >>
rect 167 433 168 434 
<< m2 >>
rect 167 433 168 434 
<< m2c >>
rect 167 433 168 434 
<< m1 >>
rect 167 433 168 434 
<< m2 >>
rect 167 433 168 434 
<< m2 >>
rect 168 433 169 434 
<< m1 >>
rect 169 433 170 434 
<< m2 >>
rect 169 433 170 434 
<< m2 >>
rect 170 433 171 434 
<< m1 >>
rect 171 433 172 434 
<< m2 >>
rect 171 433 172 434 
<< m2c >>
rect 171 433 172 434 
<< m1 >>
rect 171 433 172 434 
<< m2 >>
rect 171 433 172 434 
<< m1 >>
rect 193 433 194 434 
<< m1 >>
rect 208 433 209 434 
<< m1 >>
rect 217 433 218 434 
<< m1 >>
rect 247 433 248 434 
<< m1 >>
rect 251 433 252 434 
<< m2 >>
rect 251 433 252 434 
<< m2c >>
rect 251 433 252 434 
<< m1 >>
rect 251 433 252 434 
<< m2 >>
rect 251 433 252 434 
<< m2 >>
rect 252 433 253 434 
<< m1 >>
rect 253 433 254 434 
<< m2 >>
rect 253 433 254 434 
<< m2 >>
rect 254 433 255 434 
<< m1 >>
rect 286 433 287 434 
<< m1 >>
rect 290 433 291 434 
<< m1 >>
rect 298 433 299 434 
<< m2 >>
rect 298 433 299 434 
<< m1 >>
rect 299 433 300 434 
<< m1 >>
rect 300 433 301 434 
<< m1 >>
rect 301 433 302 434 
<< m1 >>
rect 307 433 308 434 
<< m1 >>
rect 309 433 310 434 
<< m1 >>
rect 322 433 323 434 
<< m1 >>
rect 325 433 326 434 
<< m2 >>
rect 326 433 327 434 
<< m1 >>
rect 327 433 328 434 
<< m2 >>
rect 327 433 328 434 
<< m2c >>
rect 327 433 328 434 
<< m1 >>
rect 327 433 328 434 
<< m2 >>
rect 327 433 328 434 
<< m1 >>
rect 328 433 329 434 
<< m1 >>
rect 329 433 330 434 
<< m1 >>
rect 330 433 331 434 
<< m1 >>
rect 331 433 332 434 
<< m1 >>
rect 332 433 333 434 
<< m1 >>
rect 333 433 334 434 
<< m1 >>
rect 334 433 335 434 
<< m1 >>
rect 335 433 336 434 
<< m1 >>
rect 336 433 337 434 
<< m1 >>
rect 340 433 341 434 
<< m1 >>
rect 358 433 359 434 
<< m1 >>
rect 359 433 360 434 
<< m2 >>
rect 359 433 360 434 
<< m2c >>
rect 359 433 360 434 
<< m1 >>
rect 359 433 360 434 
<< m2 >>
rect 359 433 360 434 
<< m2 >>
rect 360 433 361 434 
<< m1 >>
rect 361 433 362 434 
<< m2 >>
rect 361 433 362 434 
<< m1 >>
rect 362 433 363 434 
<< m1 >>
rect 363 433 364 434 
<< m1 >>
rect 364 433 365 434 
<< m1 >>
rect 365 433 366 434 
<< m1 >>
rect 366 433 367 434 
<< m1 >>
rect 367 433 368 434 
<< m1 >>
rect 368 433 369 434 
<< m1 >>
rect 369 433 370 434 
<< m1 >>
rect 370 433 371 434 
<< m1 >>
rect 371 433 372 434 
<< m1 >>
rect 372 433 373 434 
<< m1 >>
rect 373 433 374 434 
<< m1 >>
rect 379 433 380 434 
<< m2 >>
rect 379 433 380 434 
<< m1 >>
rect 380 433 381 434 
<< m1 >>
rect 381 433 382 434 
<< m1 >>
rect 382 433 383 434 
<< m1 >>
rect 383 433 384 434 
<< m1 >>
rect 384 433 385 434 
<< m1 >>
rect 385 433 386 434 
<< m2 >>
rect 385 433 386 434 
<< m1 >>
rect 386 433 387 434 
<< m1 >>
rect 387 433 388 434 
<< m1 >>
rect 388 433 389 434 
<< m1 >>
rect 389 433 390 434 
<< m1 >>
rect 390 433 391 434 
<< m1 >>
rect 391 433 392 434 
<< m1 >>
rect 397 433 398 434 
<< m2 >>
rect 398 433 399 434 
<< m1 >>
rect 402 433 403 434 
<< m1 >>
rect 406 433 407 434 
<< m1 >>
rect 420 433 421 434 
<< m1 >>
rect 424 433 425 434 
<< m1 >>
rect 430 433 431 434 
<< m1 >>
rect 433 433 434 434 
<< m2 >>
rect 434 433 435 434 
<< m1 >>
rect 442 433 443 434 
<< m1 >>
rect 448 433 449 434 
<< m1 >>
rect 452 433 453 434 
<< m1 >>
rect 472 433 473 434 
<< m2 >>
rect 473 433 474 434 
<< m1 >>
rect 474 433 475 434 
<< m1 >>
rect 478 433 479 434 
<< m1 >>
rect 487 433 488 434 
<< m1 >>
rect 489 433 490 434 
<< m1 >>
rect 491 433 492 434 
<< m1 >>
rect 520 433 521 434 
<< m1 >>
rect 19 434 20 435 
<< m1 >>
rect 21 434 22 435 
<< m1 >>
rect 26 434 27 435 
<< m1 >>
rect 28 434 29 435 
<< m2 >>
rect 28 434 29 435 
<< m1 >>
rect 73 434 74 435 
<< m2 >>
rect 73 434 74 435 
<< m2c >>
rect 73 434 74 435 
<< m1 >>
rect 73 434 74 435 
<< m2 >>
rect 73 434 74 435 
<< m1 >>
rect 82 434 83 435 
<< m2 >>
rect 93 434 94 435 
<< m2 >>
rect 96 434 97 435 
<< m1 >>
rect 100 434 101 435 
<< m1 >>
rect 102 434 103 435 
<< m1 >>
rect 106 434 107 435 
<< m1 >>
rect 107 434 108 435 
<< m1 >>
rect 108 434 109 435 
<< m1 >>
rect 109 434 110 435 
<< m1 >>
rect 110 434 111 435 
<< m2 >>
rect 110 434 111 435 
<< m1 >>
rect 111 434 112 435 
<< m1 >>
rect 112 434 113 435 
<< m1 >>
rect 113 434 114 435 
<< m1 >>
rect 114 434 115 435 
<< m2 >>
rect 114 434 115 435 
<< m1 >>
rect 115 434 116 435 
<< m1 >>
rect 116 434 117 435 
<< m1 >>
rect 117 434 118 435 
<< m1 >>
rect 118 434 119 435 
<< m2 >>
rect 144 434 145 435 
<< m2 >>
rect 145 434 146 435 
<< m2 >>
rect 150 434 151 435 
<< m1 >>
rect 160 434 161 435 
<< m2 >>
rect 161 434 162 435 
<< m2 >>
rect 164 434 165 435 
<< m1 >>
rect 169 434 170 435 
<< m1 >>
rect 193 434 194 435 
<< m1 >>
rect 208 434 209 435 
<< m1 >>
rect 217 434 218 435 
<< m2 >>
rect 217 434 218 435 
<< m2c >>
rect 217 434 218 435 
<< m1 >>
rect 217 434 218 435 
<< m2 >>
rect 217 434 218 435 
<< m1 >>
rect 247 434 248 435 
<< m1 >>
rect 248 434 249 435 
<< m1 >>
rect 249 434 250 435 
<< m2 >>
rect 249 434 250 435 
<< m2c >>
rect 249 434 250 435 
<< m1 >>
rect 249 434 250 435 
<< m2 >>
rect 249 434 250 435 
<< m1 >>
rect 251 434 252 435 
<< m1 >>
rect 253 434 254 435 
<< m1 >>
rect 286 434 287 435 
<< m1 >>
rect 290 434 291 435 
<< m2 >>
rect 298 434 299 435 
<< m1 >>
rect 307 434 308 435 
<< m1 >>
rect 309 434 310 435 
<< m1 >>
rect 322 434 323 435 
<< m1 >>
rect 325 434 326 435 
<< m1 >>
rect 336 434 337 435 
<< m1 >>
rect 340 434 341 435 
<< m2 >>
rect 379 434 380 435 
<< m2 >>
rect 385 434 386 435 
<< m1 >>
rect 397 434 398 435 
<< m2 >>
rect 398 434 399 435 
<< m1 >>
rect 402 434 403 435 
<< m1 >>
rect 406 434 407 435 
<< m1 >>
rect 420 434 421 435 
<< m1 >>
rect 424 434 425 435 
<< m1 >>
rect 430 434 431 435 
<< m1 >>
rect 433 434 434 435 
<< m2 >>
rect 434 434 435 435 
<< m1 >>
rect 442 434 443 435 
<< m1 >>
rect 443 434 444 435 
<< m1 >>
rect 444 434 445 435 
<< m2 >>
rect 444 434 445 435 
<< m2c >>
rect 444 434 445 435 
<< m1 >>
rect 444 434 445 435 
<< m2 >>
rect 444 434 445 435 
<< m1 >>
rect 448 434 449 435 
<< m1 >>
rect 452 434 453 435 
<< m1 >>
rect 472 434 473 435 
<< m2 >>
rect 473 434 474 435 
<< m1 >>
rect 474 434 475 435 
<< m1 >>
rect 478 434 479 435 
<< m2 >>
rect 478 434 479 435 
<< m2c >>
rect 478 434 479 435 
<< m1 >>
rect 478 434 479 435 
<< m2 >>
rect 478 434 479 435 
<< m1 >>
rect 487 434 488 435 
<< m1 >>
rect 489 434 490 435 
<< m1 >>
rect 491 434 492 435 
<< m1 >>
rect 520 434 521 435 
<< m1 >>
rect 19 435 20 436 
<< m1 >>
rect 21 435 22 436 
<< m1 >>
rect 26 435 27 436 
<< m1 >>
rect 28 435 29 436 
<< m2 >>
rect 28 435 29 436 
<< m2 >>
rect 73 435 74 436 
<< m1 >>
rect 82 435 83 436 
<< m1 >>
rect 93 435 94 436 
<< m2 >>
rect 93 435 94 436 
<< m2c >>
rect 93 435 94 436 
<< m1 >>
rect 93 435 94 436 
<< m2 >>
rect 93 435 94 436 
<< m1 >>
rect 94 435 95 436 
<< m1 >>
rect 95 435 96 436 
<< m1 >>
rect 96 435 97 436 
<< m2 >>
rect 96 435 97 436 
<< m1 >>
rect 97 435 98 436 
<< m1 >>
rect 98 435 99 436 
<< m2 >>
rect 98 435 99 436 
<< m2c >>
rect 98 435 99 436 
<< m1 >>
rect 98 435 99 436 
<< m2 >>
rect 98 435 99 436 
<< m2 >>
rect 99 435 100 436 
<< m1 >>
rect 100 435 101 436 
<< m1 >>
rect 102 435 103 436 
<< m1 >>
rect 106 435 107 436 
<< m2 >>
rect 110 435 111 436 
<< m2 >>
rect 114 435 115 436 
<< m1 >>
rect 144 435 145 436 
<< m2 >>
rect 144 435 145 436 
<< m2c >>
rect 144 435 145 436 
<< m1 >>
rect 144 435 145 436 
<< m2 >>
rect 144 435 145 436 
<< m1 >>
rect 150 435 151 436 
<< m2 >>
rect 150 435 151 436 
<< m2c >>
rect 150 435 151 436 
<< m1 >>
rect 150 435 151 436 
<< m2 >>
rect 150 435 151 436 
<< m1 >>
rect 160 435 161 436 
<< m1 >>
rect 161 435 162 436 
<< m2 >>
rect 161 435 162 436 
<< m1 >>
rect 162 435 163 436 
<< m1 >>
rect 163 435 164 436 
<< m1 >>
rect 164 435 165 436 
<< m2 >>
rect 164 435 165 436 
<< m1 >>
rect 165 435 166 436 
<< m1 >>
rect 166 435 167 436 
<< m1 >>
rect 167 435 168 436 
<< m2 >>
rect 167 435 168 436 
<< m2c >>
rect 167 435 168 436 
<< m1 >>
rect 167 435 168 436 
<< m2 >>
rect 167 435 168 436 
<< m2 >>
rect 168 435 169 436 
<< m1 >>
rect 169 435 170 436 
<< m2 >>
rect 169 435 170 436 
<< m2 >>
rect 170 435 171 436 
<< m1 >>
rect 193 435 194 436 
<< m1 >>
rect 208 435 209 436 
<< m2 >>
rect 217 435 218 436 
<< m2 >>
rect 249 435 250 436 
<< m1 >>
rect 251 435 252 436 
<< m1 >>
rect 253 435 254 436 
<< m1 >>
rect 286 435 287 436 
<< m1 >>
rect 290 435 291 436 
<< m2 >>
rect 290 435 291 436 
<< m2c >>
rect 290 435 291 436 
<< m1 >>
rect 290 435 291 436 
<< m2 >>
rect 290 435 291 436 
<< m1 >>
rect 298 435 299 436 
<< m2 >>
rect 298 435 299 436 
<< m2c >>
rect 298 435 299 436 
<< m1 >>
rect 298 435 299 436 
<< m2 >>
rect 298 435 299 436 
<< m1 >>
rect 302 435 303 436 
<< m1 >>
rect 303 435 304 436 
<< m1 >>
rect 304 435 305 436 
<< m1 >>
rect 305 435 306 436 
<< m2 >>
rect 305 435 306 436 
<< m2c >>
rect 305 435 306 436 
<< m1 >>
rect 305 435 306 436 
<< m2 >>
rect 305 435 306 436 
<< m2 >>
rect 306 435 307 436 
<< m1 >>
rect 307 435 308 436 
<< m2 >>
rect 307 435 308 436 
<< m2 >>
rect 308 435 309 436 
<< m1 >>
rect 309 435 310 436 
<< m2 >>
rect 309 435 310 436 
<< m2c >>
rect 309 435 310 436 
<< m1 >>
rect 309 435 310 436 
<< m2 >>
rect 309 435 310 436 
<< m1 >>
rect 322 435 323 436 
<< m1 >>
rect 325 435 326 436 
<< m2 >>
rect 325 435 326 436 
<< m2c >>
rect 325 435 326 436 
<< m1 >>
rect 325 435 326 436 
<< m2 >>
rect 325 435 326 436 
<< m1 >>
rect 336 435 337 436 
<< m2 >>
rect 336 435 337 436 
<< m2c >>
rect 336 435 337 436 
<< m1 >>
rect 336 435 337 436 
<< m2 >>
rect 336 435 337 436 
<< m1 >>
rect 340 435 341 436 
<< m2 >>
rect 340 435 341 436 
<< m2c >>
rect 340 435 341 436 
<< m1 >>
rect 340 435 341 436 
<< m2 >>
rect 340 435 341 436 
<< m1 >>
rect 379 435 380 436 
<< m2 >>
rect 379 435 380 436 
<< m2c >>
rect 379 435 380 436 
<< m1 >>
rect 379 435 380 436 
<< m2 >>
rect 379 435 380 436 
<< m1 >>
rect 385 435 386 436 
<< m2 >>
rect 385 435 386 436 
<< m2c >>
rect 385 435 386 436 
<< m1 >>
rect 385 435 386 436 
<< m2 >>
rect 385 435 386 436 
<< m1 >>
rect 397 435 398 436 
<< m2 >>
rect 398 435 399 436 
<< m1 >>
rect 399 435 400 436 
<< m2 >>
rect 399 435 400 436 
<< m2c >>
rect 399 435 400 436 
<< m1 >>
rect 399 435 400 436 
<< m2 >>
rect 399 435 400 436 
<< m1 >>
rect 400 435 401 436 
<< m1 >>
rect 402 435 403 436 
<< m1 >>
rect 406 435 407 436 
<< m1 >>
rect 420 435 421 436 
<< m1 >>
rect 424 435 425 436 
<< m1 >>
rect 430 435 431 436 
<< m1 >>
rect 433 435 434 436 
<< m2 >>
rect 434 435 435 436 
<< m2 >>
rect 444 435 445 436 
<< m1 >>
rect 448 435 449 436 
<< m1 >>
rect 452 435 453 436 
<< m1 >>
rect 472 435 473 436 
<< m2 >>
rect 473 435 474 436 
<< m1 >>
rect 474 435 475 436 
<< m2 >>
rect 478 435 479 436 
<< m1 >>
rect 487 435 488 436 
<< m1 >>
rect 489 435 490 436 
<< m1 >>
rect 491 435 492 436 
<< m1 >>
rect 520 435 521 436 
<< m1 >>
rect 19 436 20 437 
<< m1 >>
rect 21 436 22 437 
<< m1 >>
rect 26 436 27 437 
<< m1 >>
rect 28 436 29 437 
<< m2 >>
rect 28 436 29 437 
<< m1 >>
rect 49 436 50 437 
<< m1 >>
rect 50 436 51 437 
<< m1 >>
rect 51 436 52 437 
<< m1 >>
rect 52 436 53 437 
<< m1 >>
rect 53 436 54 437 
<< m1 >>
rect 54 436 55 437 
<< m1 >>
rect 55 436 56 437 
<< m1 >>
rect 56 436 57 437 
<< m1 >>
rect 57 436 58 437 
<< m1 >>
rect 58 436 59 437 
<< m1 >>
rect 59 436 60 437 
<< m1 >>
rect 60 436 61 437 
<< m1 >>
rect 61 436 62 437 
<< m1 >>
rect 62 436 63 437 
<< m1 >>
rect 63 436 64 437 
<< m1 >>
rect 64 436 65 437 
<< m1 >>
rect 65 436 66 437 
<< m1 >>
rect 66 436 67 437 
<< m1 >>
rect 67 436 68 437 
<< m1 >>
rect 68 436 69 437 
<< m1 >>
rect 69 436 70 437 
<< m1 >>
rect 70 436 71 437 
<< m1 >>
rect 71 436 72 437 
<< m1 >>
rect 72 436 73 437 
<< m1 >>
rect 73 436 74 437 
<< m2 >>
rect 73 436 74 437 
<< m1 >>
rect 74 436 75 437 
<< m1 >>
rect 75 436 76 437 
<< m1 >>
rect 76 436 77 437 
<< m1 >>
rect 77 436 78 437 
<< m1 >>
rect 78 436 79 437 
<< m1 >>
rect 79 436 80 437 
<< m1 >>
rect 80 436 81 437 
<< m1 >>
rect 81 436 82 437 
<< m1 >>
rect 82 436 83 437 
<< m2 >>
rect 96 436 97 437 
<< m2 >>
rect 99 436 100 437 
<< m1 >>
rect 100 436 101 437 
<< m1 >>
rect 102 436 103 437 
<< m1 >>
rect 103 436 104 437 
<< m1 >>
rect 104 436 105 437 
<< m2 >>
rect 104 436 105 437 
<< m2c >>
rect 104 436 105 437 
<< m1 >>
rect 104 436 105 437 
<< m2 >>
rect 104 436 105 437 
<< m2 >>
rect 105 436 106 437 
<< m1 >>
rect 106 436 107 437 
<< m2 >>
rect 106 436 107 437 
<< m2 >>
rect 107 436 108 437 
<< m1 >>
rect 108 436 109 437 
<< m2 >>
rect 108 436 109 437 
<< m2c >>
rect 108 436 109 437 
<< m1 >>
rect 108 436 109 437 
<< m2 >>
rect 108 436 109 437 
<< m1 >>
rect 109 436 110 437 
<< m1 >>
rect 110 436 111 437 
<< m2 >>
rect 110 436 111 437 
<< m1 >>
rect 111 436 112 437 
<< m1 >>
rect 112 436 113 437 
<< m1 >>
rect 113 436 114 437 
<< m1 >>
rect 114 436 115 437 
<< m2 >>
rect 114 436 115 437 
<< m1 >>
rect 115 436 116 437 
<< m1 >>
rect 116 436 117 437 
<< m1 >>
rect 117 436 118 437 
<< m1 >>
rect 118 436 119 437 
<< m1 >>
rect 119 436 120 437 
<< m1 >>
rect 120 436 121 437 
<< m1 >>
rect 121 436 122 437 
<< m1 >>
rect 122 436 123 437 
<< m1 >>
rect 123 436 124 437 
<< m1 >>
rect 124 436 125 437 
<< m1 >>
rect 125 436 126 437 
<< m1 >>
rect 126 436 127 437 
<< m1 >>
rect 127 436 128 437 
<< m1 >>
rect 128 436 129 437 
<< m1 >>
rect 129 436 130 437 
<< m1 >>
rect 130 436 131 437 
<< m1 >>
rect 131 436 132 437 
<< m1 >>
rect 132 436 133 437 
<< m1 >>
rect 133 436 134 437 
<< m1 >>
rect 134 436 135 437 
<< m1 >>
rect 135 436 136 437 
<< m1 >>
rect 136 436 137 437 
<< m1 >>
rect 137 436 138 437 
<< m1 >>
rect 138 436 139 437 
<< m1 >>
rect 139 436 140 437 
<< m1 >>
rect 140 436 141 437 
<< m1 >>
rect 141 436 142 437 
<< m1 >>
rect 142 436 143 437 
<< m1 >>
rect 143 436 144 437 
<< m1 >>
rect 144 436 145 437 
<< m1 >>
rect 150 436 151 437 
<< m2 >>
rect 161 436 162 437 
<< m2 >>
rect 164 436 165 437 
<< m1 >>
rect 169 436 170 437 
<< m2 >>
rect 170 436 171 437 
<< m1 >>
rect 193 436 194 437 
<< m1 >>
rect 208 436 209 437 
<< m1 >>
rect 211 436 212 437 
<< m1 >>
rect 212 436 213 437 
<< m1 >>
rect 213 436 214 437 
<< m1 >>
rect 214 436 215 437 
<< m1 >>
rect 215 436 216 437 
<< m1 >>
rect 216 436 217 437 
<< m1 >>
rect 217 436 218 437 
<< m2 >>
rect 217 436 218 437 
<< m1 >>
rect 218 436 219 437 
<< m1 >>
rect 219 436 220 437 
<< m1 >>
rect 220 436 221 437 
<< m1 >>
rect 221 436 222 437 
<< m1 >>
rect 222 436 223 437 
<< m1 >>
rect 223 436 224 437 
<< m1 >>
rect 224 436 225 437 
<< m1 >>
rect 225 436 226 437 
<< m1 >>
rect 226 436 227 437 
<< m1 >>
rect 227 436 228 437 
<< m1 >>
rect 228 436 229 437 
<< m1 >>
rect 229 436 230 437 
<< m1 >>
rect 230 436 231 437 
<< m1 >>
rect 231 436 232 437 
<< m1 >>
rect 232 436 233 437 
<< m1 >>
rect 233 436 234 437 
<< m1 >>
rect 234 436 235 437 
<< m1 >>
rect 235 436 236 437 
<< m1 >>
rect 236 436 237 437 
<< m1 >>
rect 237 436 238 437 
<< m1 >>
rect 238 436 239 437 
<< m1 >>
rect 239 436 240 437 
<< m1 >>
rect 240 436 241 437 
<< m1 >>
rect 241 436 242 437 
<< m1 >>
rect 242 436 243 437 
<< m1 >>
rect 243 436 244 437 
<< m1 >>
rect 244 436 245 437 
<< m1 >>
rect 245 436 246 437 
<< m1 >>
rect 246 436 247 437 
<< m1 >>
rect 247 436 248 437 
<< m1 >>
rect 248 436 249 437 
<< m1 >>
rect 249 436 250 437 
<< m2 >>
rect 249 436 250 437 
<< m1 >>
rect 250 436 251 437 
<< m1 >>
rect 251 436 252 437 
<< m1 >>
rect 253 436 254 437 
<< m1 >>
rect 286 436 287 437 
<< m2 >>
rect 290 436 291 437 
<< m1 >>
rect 298 436 299 437 
<< m1 >>
rect 302 436 303 437 
<< m1 >>
rect 307 436 308 437 
<< m1 >>
rect 322 436 323 437 
<< m2 >>
rect 325 436 326 437 
<< m2 >>
rect 336 436 337 437 
<< m2 >>
rect 337 436 338 437 
<< m2 >>
rect 338 436 339 437 
<< m2 >>
rect 339 436 340 437 
<< m2 >>
rect 340 436 341 437 
<< m1 >>
rect 379 436 380 437 
<< m1 >>
rect 385 436 386 437 
<< m1 >>
rect 397 436 398 437 
<< m1 >>
rect 400 436 401 437 
<< m1 >>
rect 402 436 403 437 
<< m1 >>
rect 406 436 407 437 
<< m1 >>
rect 420 436 421 437 
<< m1 >>
rect 424 436 425 437 
<< m1 >>
rect 425 436 426 437 
<< m1 >>
rect 426 436 427 437 
<< m1 >>
rect 427 436 428 437 
<< m1 >>
rect 428 436 429 437 
<< m1 >>
rect 429 436 430 437 
<< m1 >>
rect 430 436 431 437 
<< m1 >>
rect 433 436 434 437 
<< m2 >>
rect 434 436 435 437 
<< m1 >>
rect 435 436 436 437 
<< m2 >>
rect 435 436 436 437 
<< m2c >>
rect 435 436 436 437 
<< m1 >>
rect 435 436 436 437 
<< m2 >>
rect 435 436 436 437 
<< m1 >>
rect 436 436 437 437 
<< m1 >>
rect 437 436 438 437 
<< m1 >>
rect 438 436 439 437 
<< m1 >>
rect 439 436 440 437 
<< m1 >>
rect 440 436 441 437 
<< m1 >>
rect 441 436 442 437 
<< m1 >>
rect 442 436 443 437 
<< m1 >>
rect 443 436 444 437 
<< m1 >>
rect 444 436 445 437 
<< m2 >>
rect 444 436 445 437 
<< m1 >>
rect 445 436 446 437 
<< m1 >>
rect 446 436 447 437 
<< m1 >>
rect 447 436 448 437 
<< m1 >>
rect 448 436 449 437 
<< m1 >>
rect 452 436 453 437 
<< m1 >>
rect 472 436 473 437 
<< m2 >>
rect 473 436 474 437 
<< m1 >>
rect 474 436 475 437 
<< m1 >>
rect 475 436 476 437 
<< m1 >>
rect 476 436 477 437 
<< m1 >>
rect 477 436 478 437 
<< m1 >>
rect 478 436 479 437 
<< m2 >>
rect 478 436 479 437 
<< m1 >>
rect 479 436 480 437 
<< m1 >>
rect 480 436 481 437 
<< m1 >>
rect 481 436 482 437 
<< m1 >>
rect 482 436 483 437 
<< m1 >>
rect 483 436 484 437 
<< m1 >>
rect 484 436 485 437 
<< m1 >>
rect 485 436 486 437 
<< m2 >>
rect 485 436 486 437 
<< m2c >>
rect 485 436 486 437 
<< m1 >>
rect 485 436 486 437 
<< m2 >>
rect 485 436 486 437 
<< m2 >>
rect 486 436 487 437 
<< m1 >>
rect 487 436 488 437 
<< m2 >>
rect 487 436 488 437 
<< m2 >>
rect 488 436 489 437 
<< m1 >>
rect 489 436 490 437 
<< m2 >>
rect 489 436 490 437 
<< m2 >>
rect 490 436 491 437 
<< m1 >>
rect 491 436 492 437 
<< m2 >>
rect 491 436 492 437 
<< m1 >>
rect 492 436 493 437 
<< m2 >>
rect 492 436 493 437 
<< m1 >>
rect 493 436 494 437 
<< m2 >>
rect 493 436 494 437 
<< m1 >>
rect 494 436 495 437 
<< m2 >>
rect 494 436 495 437 
<< m1 >>
rect 495 436 496 437 
<< m2 >>
rect 495 436 496 437 
<< m1 >>
rect 496 436 497 437 
<< m2 >>
rect 496 436 497 437 
<< m1 >>
rect 497 436 498 437 
<< m2 >>
rect 497 436 498 437 
<< m1 >>
rect 498 436 499 437 
<< m2 >>
rect 498 436 499 437 
<< m1 >>
rect 499 436 500 437 
<< m2 >>
rect 499 436 500 437 
<< m1 >>
rect 500 436 501 437 
<< m2 >>
rect 500 436 501 437 
<< m1 >>
rect 501 436 502 437 
<< m2 >>
rect 501 436 502 437 
<< m1 >>
rect 502 436 503 437 
<< m2 >>
rect 502 436 503 437 
<< m2 >>
rect 503 436 504 437 
<< m1 >>
rect 504 436 505 437 
<< m2 >>
rect 504 436 505 437 
<< m2c >>
rect 504 436 505 437 
<< m1 >>
rect 504 436 505 437 
<< m2 >>
rect 504 436 505 437 
<< m1 >>
rect 505 436 506 437 
<< m1 >>
rect 506 436 507 437 
<< m1 >>
rect 507 436 508 437 
<< m1 >>
rect 508 436 509 437 
<< m1 >>
rect 509 436 510 437 
<< m1 >>
rect 510 436 511 437 
<< m1 >>
rect 511 436 512 437 
<< m1 >>
rect 512 436 513 437 
<< m1 >>
rect 513 436 514 437 
<< m1 >>
rect 514 436 515 437 
<< m1 >>
rect 515 436 516 437 
<< m1 >>
rect 516 436 517 437 
<< m1 >>
rect 517 436 518 437 
<< m1 >>
rect 518 436 519 437 
<< m1 >>
rect 519 436 520 437 
<< m1 >>
rect 520 436 521 437 
<< m1 >>
rect 19 437 20 438 
<< m1 >>
rect 21 437 22 438 
<< m1 >>
rect 26 437 27 438 
<< m1 >>
rect 28 437 29 438 
<< m2 >>
rect 28 437 29 438 
<< m1 >>
rect 49 437 50 438 
<< m2 >>
rect 73 437 74 438 
<< m1 >>
rect 96 437 97 438 
<< m2 >>
rect 96 437 97 438 
<< m2c >>
rect 96 437 97 438 
<< m1 >>
rect 96 437 97 438 
<< m2 >>
rect 96 437 97 438 
<< m2 >>
rect 99 437 100 438 
<< m1 >>
rect 100 437 101 438 
<< m1 >>
rect 106 437 107 438 
<< m2 >>
rect 110 437 111 438 
<< m2 >>
rect 114 437 115 438 
<< m2 >>
rect 115 437 116 438 
<< m2 >>
rect 116 437 117 438 
<< m2 >>
rect 117 437 118 438 
<< m2 >>
rect 118 437 119 438 
<< m2 >>
rect 119 437 120 438 
<< m2 >>
rect 120 437 121 438 
<< m2 >>
rect 121 437 122 438 
<< m2 >>
rect 122 437 123 438 
<< m2 >>
rect 123 437 124 438 
<< m2 >>
rect 124 437 125 438 
<< m2 >>
rect 125 437 126 438 
<< m2 >>
rect 126 437 127 438 
<< m2 >>
rect 127 437 128 438 
<< m2 >>
rect 128 437 129 438 
<< m2 >>
rect 129 437 130 438 
<< m2 >>
rect 130 437 131 438 
<< m2 >>
rect 131 437 132 438 
<< m2 >>
rect 132 437 133 438 
<< m2 >>
rect 133 437 134 438 
<< m2 >>
rect 134 437 135 438 
<< m2 >>
rect 135 437 136 438 
<< m2 >>
rect 136 437 137 438 
<< m2 >>
rect 137 437 138 438 
<< m2 >>
rect 138 437 139 438 
<< m2 >>
rect 139 437 140 438 
<< m2 >>
rect 140 437 141 438 
<< m2 >>
rect 141 437 142 438 
<< m2 >>
rect 142 437 143 438 
<< m2 >>
rect 143 437 144 438 
<< m2 >>
rect 144 437 145 438 
<< m2 >>
rect 145 437 146 438 
<< m1 >>
rect 146 437 147 438 
<< m2 >>
rect 146 437 147 438 
<< m2c >>
rect 146 437 147 438 
<< m1 >>
rect 146 437 147 438 
<< m2 >>
rect 146 437 147 438 
<< m1 >>
rect 147 437 148 438 
<< m1 >>
rect 148 437 149 438 
<< m2 >>
rect 148 437 149 438 
<< m2c >>
rect 148 437 149 438 
<< m1 >>
rect 148 437 149 438 
<< m2 >>
rect 148 437 149 438 
<< m2 >>
rect 149 437 150 438 
<< m1 >>
rect 150 437 151 438 
<< m2 >>
rect 150 437 151 438 
<< m2 >>
rect 151 437 152 438 
<< m1 >>
rect 152 437 153 438 
<< m2 >>
rect 152 437 153 438 
<< m2c >>
rect 152 437 153 438 
<< m1 >>
rect 152 437 153 438 
<< m2 >>
rect 152 437 153 438 
<< m1 >>
rect 153 437 154 438 
<< m1 >>
rect 154 437 155 438 
<< m1 >>
rect 155 437 156 438 
<< m1 >>
rect 156 437 157 438 
<< m1 >>
rect 157 437 158 438 
<< m1 >>
rect 158 437 159 438 
<< m1 >>
rect 159 437 160 438 
<< m1 >>
rect 160 437 161 438 
<< m1 >>
rect 161 437 162 438 
<< m2 >>
rect 161 437 162 438 
<< m1 >>
rect 162 437 163 438 
<< m1 >>
rect 163 437 164 438 
<< m1 >>
rect 164 437 165 438 
<< m2 >>
rect 164 437 165 438 
<< m1 >>
rect 165 437 166 438 
<< m1 >>
rect 166 437 167 438 
<< m1 >>
rect 167 437 168 438 
<< m1 >>
rect 168 437 169 438 
<< m1 >>
rect 169 437 170 438 
<< m2 >>
rect 170 437 171 438 
<< m1 >>
rect 193 437 194 438 
<< m1 >>
rect 208 437 209 438 
<< m1 >>
rect 211 437 212 438 
<< m2 >>
rect 217 437 218 438 
<< m2 >>
rect 249 437 250 438 
<< m1 >>
rect 253 437 254 438 
<< m2 >>
rect 285 437 286 438 
<< m1 >>
rect 286 437 287 438 
<< m2 >>
rect 286 437 287 438 
<< m2 >>
rect 287 437 288 438 
<< m1 >>
rect 288 437 289 438 
<< m2 >>
rect 288 437 289 438 
<< m2c >>
rect 288 437 289 438 
<< m1 >>
rect 288 437 289 438 
<< m2 >>
rect 288 437 289 438 
<< m1 >>
rect 289 437 290 438 
<< m1 >>
rect 290 437 291 438 
<< m2 >>
rect 290 437 291 438 
<< m1 >>
rect 291 437 292 438 
<< m1 >>
rect 292 437 293 438 
<< m1 >>
rect 293 437 294 438 
<< m1 >>
rect 294 437 295 438 
<< m1 >>
rect 295 437 296 438 
<< m1 >>
rect 296 437 297 438 
<< m2 >>
rect 296 437 297 438 
<< m2c >>
rect 296 437 297 438 
<< m1 >>
rect 296 437 297 438 
<< m2 >>
rect 296 437 297 438 
<< m2 >>
rect 297 437 298 438 
<< m1 >>
rect 298 437 299 438 
<< m2 >>
rect 298 437 299 438 
<< m2 >>
rect 299 437 300 438 
<< m1 >>
rect 300 437 301 438 
<< m2 >>
rect 300 437 301 438 
<< m2c >>
rect 300 437 301 438 
<< m1 >>
rect 300 437 301 438 
<< m2 >>
rect 300 437 301 438 
<< m1 >>
rect 301 437 302 438 
<< m1 >>
rect 302 437 303 438 
<< m1 >>
rect 307 437 308 438 
<< m2 >>
rect 307 437 308 438 
<< m2c >>
rect 307 437 308 438 
<< m1 >>
rect 307 437 308 438 
<< m2 >>
rect 307 437 308 438 
<< m1 >>
rect 322 437 323 438 
<< m1 >>
rect 323 437 324 438 
<< m1 >>
rect 324 437 325 438 
<< m1 >>
rect 325 437 326 438 
<< m2 >>
rect 325 437 326 438 
<< m1 >>
rect 326 437 327 438 
<< m1 >>
rect 327 437 328 438 
<< m1 >>
rect 328 437 329 438 
<< m1 >>
rect 329 437 330 438 
<< m1 >>
rect 330 437 331 438 
<< m1 >>
rect 331 437 332 438 
<< m1 >>
rect 332 437 333 438 
<< m1 >>
rect 333 437 334 438 
<< m1 >>
rect 334 437 335 438 
<< m1 >>
rect 335 437 336 438 
<< m1 >>
rect 336 437 337 438 
<< m1 >>
rect 337 437 338 438 
<< m1 >>
rect 338 437 339 438 
<< m1 >>
rect 339 437 340 438 
<< m1 >>
rect 340 437 341 438 
<< m1 >>
rect 341 437 342 438 
<< m1 >>
rect 342 437 343 438 
<< m1 >>
rect 343 437 344 438 
<< m1 >>
rect 344 437 345 438 
<< m1 >>
rect 345 437 346 438 
<< m1 >>
rect 346 437 347 438 
<< m1 >>
rect 347 437 348 438 
<< m1 >>
rect 348 437 349 438 
<< m1 >>
rect 349 437 350 438 
<< m1 >>
rect 350 437 351 438 
<< m1 >>
rect 351 437 352 438 
<< m1 >>
rect 352 437 353 438 
<< m1 >>
rect 353 437 354 438 
<< m1 >>
rect 354 437 355 438 
<< m1 >>
rect 355 437 356 438 
<< m1 >>
rect 356 437 357 438 
<< m1 >>
rect 357 437 358 438 
<< m1 >>
rect 358 437 359 438 
<< m1 >>
rect 359 437 360 438 
<< m1 >>
rect 360 437 361 438 
<< m1 >>
rect 361 437 362 438 
<< m2 >>
rect 361 437 362 438 
<< m2c >>
rect 361 437 362 438 
<< m1 >>
rect 361 437 362 438 
<< m2 >>
rect 361 437 362 438 
<< m1 >>
rect 379 437 380 438 
<< m2 >>
rect 379 437 380 438 
<< m2c >>
rect 379 437 380 438 
<< m1 >>
rect 379 437 380 438 
<< m2 >>
rect 379 437 380 438 
<< m1 >>
rect 385 437 386 438 
<< m2 >>
rect 385 437 386 438 
<< m2c >>
rect 385 437 386 438 
<< m1 >>
rect 385 437 386 438 
<< m2 >>
rect 385 437 386 438 
<< m1 >>
rect 397 437 398 438 
<< m2 >>
rect 397 437 398 438 
<< m2c >>
rect 397 437 398 438 
<< m1 >>
rect 397 437 398 438 
<< m2 >>
rect 397 437 398 438 
<< m1 >>
rect 400 437 401 438 
<< m2 >>
rect 400 437 401 438 
<< m2c >>
rect 400 437 401 438 
<< m1 >>
rect 400 437 401 438 
<< m2 >>
rect 400 437 401 438 
<< m1 >>
rect 402 437 403 438 
<< m2 >>
rect 402 437 403 438 
<< m2c >>
rect 402 437 403 438 
<< m1 >>
rect 402 437 403 438 
<< m2 >>
rect 402 437 403 438 
<< m1 >>
rect 406 437 407 438 
<< m2 >>
rect 406 437 407 438 
<< m2c >>
rect 406 437 407 438 
<< m1 >>
rect 406 437 407 438 
<< m2 >>
rect 406 437 407 438 
<< m1 >>
rect 420 437 421 438 
<< m1 >>
rect 421 437 422 438 
<< m1 >>
rect 422 437 423 438 
<< m2 >>
rect 422 437 423 438 
<< m2c >>
rect 422 437 423 438 
<< m1 >>
rect 422 437 423 438 
<< m2 >>
rect 422 437 423 438 
<< m2 >>
rect 423 437 424 438 
<< m2 >>
rect 424 437 425 438 
<< m1 >>
rect 433 437 434 438 
<< m2 >>
rect 444 437 445 438 
<< m1 >>
rect 452 437 453 438 
<< m2 >>
rect 452 437 453 438 
<< m2c >>
rect 452 437 453 438 
<< m1 >>
rect 452 437 453 438 
<< m2 >>
rect 452 437 453 438 
<< m1 >>
rect 472 437 473 438 
<< m2 >>
rect 473 437 474 438 
<< m2 >>
rect 478 437 479 438 
<< m1 >>
rect 487 437 488 438 
<< m1 >>
rect 489 437 490 438 
<< m1 >>
rect 502 437 503 438 
<< m1 >>
rect 19 438 20 439 
<< m1 >>
rect 21 438 22 439 
<< m1 >>
rect 26 438 27 439 
<< m1 >>
rect 28 438 29 439 
<< m2 >>
rect 28 438 29 439 
<< m1 >>
rect 49 438 50 439 
<< m1 >>
rect 73 438 74 439 
<< m2 >>
rect 73 438 74 439 
<< m2c >>
rect 73 438 74 439 
<< m1 >>
rect 73 438 74 439 
<< m2 >>
rect 73 438 74 439 
<< m1 >>
rect 96 438 97 439 
<< m2 >>
rect 99 438 100 439 
<< m1 >>
rect 100 438 101 439 
<< m2 >>
rect 100 438 101 439 
<< m2 >>
rect 101 438 102 439 
<< m1 >>
rect 102 438 103 439 
<< m2 >>
rect 102 438 103 439 
<< m2c >>
rect 102 438 103 439 
<< m1 >>
rect 102 438 103 439 
<< m2 >>
rect 102 438 103 439 
<< m1 >>
rect 103 438 104 439 
<< m1 >>
rect 104 438 105 439 
<< m2 >>
rect 104 438 105 439 
<< m2c >>
rect 104 438 105 439 
<< m1 >>
rect 104 438 105 439 
<< m2 >>
rect 104 438 105 439 
<< m2 >>
rect 105 438 106 439 
<< m1 >>
rect 106 438 107 439 
<< m2 >>
rect 106 438 107 439 
<< m2 >>
rect 107 438 108 439 
<< m1 >>
rect 108 438 109 439 
<< m2 >>
rect 108 438 109 439 
<< m2c >>
rect 108 438 109 439 
<< m1 >>
rect 108 438 109 439 
<< m2 >>
rect 108 438 109 439 
<< m2 >>
rect 110 438 111 439 
<< m1 >>
rect 150 438 151 439 
<< m2 >>
rect 161 438 162 439 
<< m2 >>
rect 164 438 165 439 
<< m2 >>
rect 170 438 171 439 
<< m1 >>
rect 193 438 194 439 
<< m1 >>
rect 208 438 209 439 
<< m1 >>
rect 211 438 212 439 
<< m2 >>
rect 217 438 218 439 
<< m2 >>
rect 249 438 250 439 
<< m1 >>
rect 253 438 254 439 
<< m2 >>
rect 285 438 286 439 
<< m1 >>
rect 286 438 287 439 
<< m2 >>
rect 290 438 291 439 
<< m1 >>
rect 298 438 299 439 
<< m2 >>
rect 307 438 308 439 
<< m2 >>
rect 325 438 326 439 
<< m2 >>
rect 361 438 362 439 
<< m2 >>
rect 379 438 380 439 
<< m2 >>
rect 385 438 386 439 
<< m2 >>
rect 397 438 398 439 
<< m2 >>
rect 400 438 401 439 
<< m2 >>
rect 402 438 403 439 
<< m2 >>
rect 406 438 407 439 
<< m2 >>
rect 424 438 425 439 
<< m1 >>
rect 433 438 434 439 
<< m2 >>
rect 444 438 445 439 
<< m2 >>
rect 452 438 453 439 
<< m2 >>
rect 462 438 463 439 
<< m2 >>
rect 463 438 464 439 
<< m2 >>
rect 464 438 465 439 
<< m2 >>
rect 465 438 466 439 
<< m2 >>
rect 466 438 467 439 
<< m2 >>
rect 467 438 468 439 
<< m2 >>
rect 468 438 469 439 
<< m2 >>
rect 469 438 470 439 
<< m2 >>
rect 470 438 471 439 
<< m2 >>
rect 471 438 472 439 
<< m1 >>
rect 472 438 473 439 
<< m2 >>
rect 472 438 473 439 
<< m2 >>
rect 473 438 474 439 
<< m1 >>
rect 478 438 479 439 
<< m2 >>
rect 478 438 479 439 
<< m2c >>
rect 478 438 479 439 
<< m1 >>
rect 478 438 479 439 
<< m2 >>
rect 478 438 479 439 
<< m1 >>
rect 487 438 488 439 
<< m1 >>
rect 489 438 490 439 
<< m1 >>
rect 502 438 503 439 
<< m1 >>
rect 19 439 20 440 
<< m1 >>
rect 21 439 22 440 
<< m1 >>
rect 26 439 27 440 
<< m1 >>
rect 28 439 29 440 
<< m2 >>
rect 28 439 29 440 
<< m1 >>
rect 49 439 50 440 
<< m1 >>
rect 73 439 74 440 
<< m1 >>
rect 96 439 97 440 
<< m1 >>
rect 100 439 101 440 
<< m1 >>
rect 106 439 107 440 
<< m1 >>
rect 108 439 109 440 
<< m1 >>
rect 109 439 110 440 
<< m1 >>
rect 110 439 111 440 
<< m2 >>
rect 110 439 111 440 
<< m1 >>
rect 111 439 112 440 
<< m2 >>
rect 111 439 112 440 
<< m1 >>
rect 112 439 113 440 
<< m2 >>
rect 112 439 113 440 
<< m1 >>
rect 113 439 114 440 
<< m2 >>
rect 113 439 114 440 
<< m1 >>
rect 114 439 115 440 
<< m2 >>
rect 114 439 115 440 
<< m1 >>
rect 115 439 116 440 
<< m2 >>
rect 115 439 116 440 
<< m1 >>
rect 116 439 117 440 
<< m2 >>
rect 116 439 117 440 
<< m1 >>
rect 117 439 118 440 
<< m2 >>
rect 117 439 118 440 
<< m1 >>
rect 118 439 119 440 
<< m2 >>
rect 118 439 119 440 
<< m1 >>
rect 119 439 120 440 
<< m2 >>
rect 119 439 120 440 
<< m1 >>
rect 120 439 121 440 
<< m2 >>
rect 120 439 121 440 
<< m1 >>
rect 121 439 122 440 
<< m2 >>
rect 121 439 122 440 
<< m1 >>
rect 122 439 123 440 
<< m2 >>
rect 122 439 123 440 
<< m1 >>
rect 123 439 124 440 
<< m1 >>
rect 124 439 125 440 
<< m1 >>
rect 125 439 126 440 
<< m1 >>
rect 126 439 127 440 
<< m1 >>
rect 127 439 128 440 
<< m1 >>
rect 128 439 129 440 
<< m1 >>
rect 129 439 130 440 
<< m1 >>
rect 130 439 131 440 
<< m1 >>
rect 131 439 132 440 
<< m1 >>
rect 132 439 133 440 
<< m1 >>
rect 133 439 134 440 
<< m1 >>
rect 134 439 135 440 
<< m1 >>
rect 135 439 136 440 
<< m1 >>
rect 136 439 137 440 
<< m1 >>
rect 137 439 138 440 
<< m1 >>
rect 138 439 139 440 
<< m1 >>
rect 139 439 140 440 
<< m1 >>
rect 140 439 141 440 
<< m1 >>
rect 141 439 142 440 
<< m1 >>
rect 142 439 143 440 
<< m1 >>
rect 143 439 144 440 
<< m1 >>
rect 144 439 145 440 
<< m1 >>
rect 145 439 146 440 
<< m1 >>
rect 146 439 147 440 
<< m1 >>
rect 147 439 148 440 
<< m1 >>
rect 148 439 149 440 
<< m2 >>
rect 148 439 149 440 
<< m2c >>
rect 148 439 149 440 
<< m1 >>
rect 148 439 149 440 
<< m2 >>
rect 148 439 149 440 
<< m2 >>
rect 149 439 150 440 
<< m1 >>
rect 150 439 151 440 
<< m2 >>
rect 150 439 151 440 
<< m2 >>
rect 151 439 152 440 
<< m1 >>
rect 152 439 153 440 
<< m2 >>
rect 152 439 153 440 
<< m1 >>
rect 153 439 154 440 
<< m2 >>
rect 153 439 154 440 
<< m1 >>
rect 154 439 155 440 
<< m2 >>
rect 154 439 155 440 
<< m1 >>
rect 155 439 156 440 
<< m2 >>
rect 155 439 156 440 
<< m1 >>
rect 156 439 157 440 
<< m2 >>
rect 156 439 157 440 
<< m1 >>
rect 157 439 158 440 
<< m2 >>
rect 157 439 158 440 
<< m1 >>
rect 158 439 159 440 
<< m2 >>
rect 158 439 159 440 
<< m1 >>
rect 159 439 160 440 
<< m2 >>
rect 159 439 160 440 
<< m1 >>
rect 160 439 161 440 
<< m2 >>
rect 160 439 161 440 
<< m1 >>
rect 161 439 162 440 
<< m2 >>
rect 161 439 162 440 
<< m1 >>
rect 162 439 163 440 
<< m1 >>
rect 163 439 164 440 
<< m1 >>
rect 164 439 165 440 
<< m2 >>
rect 164 439 165 440 
<< m1 >>
rect 165 439 166 440 
<< m1 >>
rect 166 439 167 440 
<< m1 >>
rect 167 439 168 440 
<< m1 >>
rect 168 439 169 440 
<< m1 >>
rect 169 439 170 440 
<< m1 >>
rect 170 439 171 440 
<< m2 >>
rect 170 439 171 440 
<< m1 >>
rect 171 439 172 440 
<< m2 >>
rect 171 439 172 440 
<< m1 >>
rect 172 439 173 440 
<< m2 >>
rect 172 439 173 440 
<< m1 >>
rect 173 439 174 440 
<< m2 >>
rect 173 439 174 440 
<< m1 >>
rect 174 439 175 440 
<< m2 >>
rect 174 439 175 440 
<< m1 >>
rect 175 439 176 440 
<< m2 >>
rect 175 439 176 440 
<< m1 >>
rect 176 439 177 440 
<< m2 >>
rect 176 439 177 440 
<< m1 >>
rect 177 439 178 440 
<< m2 >>
rect 177 439 178 440 
<< m1 >>
rect 178 439 179 440 
<< m2 >>
rect 178 439 179 440 
<< m1 >>
rect 179 439 180 440 
<< m2 >>
rect 179 439 180 440 
<< m1 >>
rect 180 439 181 440 
<< m2 >>
rect 180 439 181 440 
<< m1 >>
rect 181 439 182 440 
<< m2 >>
rect 181 439 182 440 
<< m1 >>
rect 182 439 183 440 
<< m2 >>
rect 182 439 183 440 
<< m1 >>
rect 183 439 184 440 
<< m2 >>
rect 183 439 184 440 
<< m1 >>
rect 184 439 185 440 
<< m2 >>
rect 184 439 185 440 
<< m1 >>
rect 185 439 186 440 
<< m2 >>
rect 185 439 186 440 
<< m1 >>
rect 186 439 187 440 
<< m2 >>
rect 186 439 187 440 
<< m1 >>
rect 187 439 188 440 
<< m2 >>
rect 187 439 188 440 
<< m1 >>
rect 188 439 189 440 
<< m2 >>
rect 188 439 189 440 
<< m1 >>
rect 189 439 190 440 
<< m2 >>
rect 189 439 190 440 
<< m1 >>
rect 190 439 191 440 
<< m2 >>
rect 190 439 191 440 
<< m1 >>
rect 191 439 192 440 
<< m2 >>
rect 191 439 192 440 
<< m1 >>
rect 192 439 193 440 
<< m2 >>
rect 192 439 193 440 
<< m1 >>
rect 193 439 194 440 
<< m2 >>
rect 193 439 194 440 
<< m2 >>
rect 194 439 195 440 
<< m2 >>
rect 207 439 208 440 
<< m1 >>
rect 208 439 209 440 
<< m2 >>
rect 208 439 209 440 
<< m2 >>
rect 209 439 210 440 
<< m2 >>
rect 210 439 211 440 
<< m1 >>
rect 211 439 212 440 
<< m2 >>
rect 211 439 212 440 
<< m2 >>
rect 212 439 213 440 
<< m1 >>
rect 213 439 214 440 
<< m2 >>
rect 213 439 214 440 
<< m2c >>
rect 213 439 214 440 
<< m1 >>
rect 213 439 214 440 
<< m2 >>
rect 213 439 214 440 
<< m1 >>
rect 214 439 215 440 
<< m1 >>
rect 215 439 216 440 
<< m1 >>
rect 216 439 217 440 
<< m1 >>
rect 217 439 218 440 
<< m2 >>
rect 217 439 218 440 
<< m1 >>
rect 218 439 219 440 
<< m1 >>
rect 219 439 220 440 
<< m1 >>
rect 220 439 221 440 
<< m1 >>
rect 221 439 222 440 
<< m1 >>
rect 222 439 223 440 
<< m1 >>
rect 223 439 224 440 
<< m1 >>
rect 224 439 225 440 
<< m1 >>
rect 225 439 226 440 
<< m1 >>
rect 226 439 227 440 
<< m1 >>
rect 227 439 228 440 
<< m1 >>
rect 228 439 229 440 
<< m1 >>
rect 229 439 230 440 
<< m1 >>
rect 230 439 231 440 
<< m1 >>
rect 231 439 232 440 
<< m1 >>
rect 232 439 233 440 
<< m1 >>
rect 233 439 234 440 
<< m1 >>
rect 234 439 235 440 
<< m1 >>
rect 235 439 236 440 
<< m1 >>
rect 236 439 237 440 
<< m1 >>
rect 237 439 238 440 
<< m1 >>
rect 238 439 239 440 
<< m1 >>
rect 239 439 240 440 
<< m1 >>
rect 240 439 241 440 
<< m1 >>
rect 241 439 242 440 
<< m1 >>
rect 242 439 243 440 
<< m1 >>
rect 243 439 244 440 
<< m1 >>
rect 244 439 245 440 
<< m1 >>
rect 245 439 246 440 
<< m1 >>
rect 246 439 247 440 
<< m1 >>
rect 247 439 248 440 
<< m1 >>
rect 248 439 249 440 
<< m1 >>
rect 249 439 250 440 
<< m2 >>
rect 249 439 250 440 
<< m1 >>
rect 250 439 251 440 
<< m1 >>
rect 251 439 252 440 
<< m2 >>
rect 251 439 252 440 
<< m2c >>
rect 251 439 252 440 
<< m1 >>
rect 251 439 252 440 
<< m2 >>
rect 251 439 252 440 
<< m2 >>
rect 252 439 253 440 
<< m1 >>
rect 253 439 254 440 
<< m2 >>
rect 253 439 254 440 
<< m2 >>
rect 254 439 255 440 
<< m1 >>
rect 255 439 256 440 
<< m2 >>
rect 255 439 256 440 
<< m2c >>
rect 255 439 256 440 
<< m1 >>
rect 255 439 256 440 
<< m2 >>
rect 255 439 256 440 
<< m1 >>
rect 256 439 257 440 
<< m1 >>
rect 257 439 258 440 
<< m1 >>
rect 258 439 259 440 
<< m1 >>
rect 259 439 260 440 
<< m1 >>
rect 260 439 261 440 
<< m1 >>
rect 261 439 262 440 
<< m1 >>
rect 262 439 263 440 
<< m1 >>
rect 263 439 264 440 
<< m1 >>
rect 264 439 265 440 
<< m1 >>
rect 265 439 266 440 
<< m1 >>
rect 266 439 267 440 
<< m1 >>
rect 267 439 268 440 
<< m1 >>
rect 268 439 269 440 
<< m1 >>
rect 269 439 270 440 
<< m1 >>
rect 270 439 271 440 
<< m1 >>
rect 271 439 272 440 
<< m1 >>
rect 272 439 273 440 
<< m1 >>
rect 273 439 274 440 
<< m1 >>
rect 274 439 275 440 
<< m1 >>
rect 275 439 276 440 
<< m1 >>
rect 276 439 277 440 
<< m1 >>
rect 277 439 278 440 
<< m1 >>
rect 278 439 279 440 
<< m1 >>
rect 279 439 280 440 
<< m1 >>
rect 280 439 281 440 
<< m1 >>
rect 281 439 282 440 
<< m1 >>
rect 282 439 283 440 
<< m1 >>
rect 283 439 284 440 
<< m1 >>
rect 284 439 285 440 
<< m2 >>
rect 284 439 285 440 
<< m2c >>
rect 284 439 285 440 
<< m1 >>
rect 284 439 285 440 
<< m2 >>
rect 284 439 285 440 
<< m2 >>
rect 285 439 286 440 
<< m1 >>
rect 286 439 287 440 
<< m1 >>
rect 287 439 288 440 
<< m1 >>
rect 288 439 289 440 
<< m1 >>
rect 289 439 290 440 
<< m1 >>
rect 290 439 291 440 
<< m2 >>
rect 290 439 291 440 
<< m1 >>
rect 291 439 292 440 
<< m1 >>
rect 292 439 293 440 
<< m1 >>
rect 293 439 294 440 
<< m1 >>
rect 294 439 295 440 
<< m1 >>
rect 295 439 296 440 
<< m1 >>
rect 296 439 297 440 
<< m2 >>
rect 296 439 297 440 
<< m2c >>
rect 296 439 297 440 
<< m1 >>
rect 296 439 297 440 
<< m2 >>
rect 296 439 297 440 
<< m2 >>
rect 297 439 298 440 
<< m1 >>
rect 298 439 299 440 
<< m2 >>
rect 298 439 299 440 
<< m2 >>
rect 299 439 300 440 
<< m1 >>
rect 300 439 301 440 
<< m2 >>
rect 300 439 301 440 
<< m2c >>
rect 300 439 301 440 
<< m1 >>
rect 300 439 301 440 
<< m2 >>
rect 300 439 301 440 
<< m1 >>
rect 301 439 302 440 
<< m1 >>
rect 302 439 303 440 
<< m1 >>
rect 303 439 304 440 
<< m1 >>
rect 304 439 305 440 
<< m1 >>
rect 305 439 306 440 
<< m1 >>
rect 306 439 307 440 
<< m1 >>
rect 307 439 308 440 
<< m2 >>
rect 307 439 308 440 
<< m1 >>
rect 308 439 309 440 
<< m1 >>
rect 309 439 310 440 
<< m1 >>
rect 310 439 311 440 
<< m1 >>
rect 311 439 312 440 
<< m1 >>
rect 312 439 313 440 
<< m1 >>
rect 313 439 314 440 
<< m1 >>
rect 314 439 315 440 
<< m1 >>
rect 315 439 316 440 
<< m1 >>
rect 316 439 317 440 
<< m1 >>
rect 317 439 318 440 
<< m1 >>
rect 318 439 319 440 
<< m1 >>
rect 319 439 320 440 
<< m1 >>
rect 320 439 321 440 
<< m1 >>
rect 321 439 322 440 
<< m1 >>
rect 322 439 323 440 
<< m1 >>
rect 323 439 324 440 
<< m1 >>
rect 324 439 325 440 
<< m1 >>
rect 325 439 326 440 
<< m2 >>
rect 325 439 326 440 
<< m1 >>
rect 326 439 327 440 
<< m1 >>
rect 327 439 328 440 
<< m1 >>
rect 328 439 329 440 
<< m1 >>
rect 329 439 330 440 
<< m1 >>
rect 330 439 331 440 
<< m1 >>
rect 331 439 332 440 
<< m1 >>
rect 332 439 333 440 
<< m1 >>
rect 333 439 334 440 
<< m1 >>
rect 334 439 335 440 
<< m1 >>
rect 335 439 336 440 
<< m1 >>
rect 336 439 337 440 
<< m1 >>
rect 337 439 338 440 
<< m1 >>
rect 338 439 339 440 
<< m1 >>
rect 339 439 340 440 
<< m1 >>
rect 340 439 341 440 
<< m1 >>
rect 341 439 342 440 
<< m1 >>
rect 342 439 343 440 
<< m1 >>
rect 343 439 344 440 
<< m1 >>
rect 344 439 345 440 
<< m1 >>
rect 345 439 346 440 
<< m1 >>
rect 346 439 347 440 
<< m1 >>
rect 347 439 348 440 
<< m1 >>
rect 348 439 349 440 
<< m1 >>
rect 349 439 350 440 
<< m1 >>
rect 350 439 351 440 
<< m1 >>
rect 351 439 352 440 
<< m1 >>
rect 352 439 353 440 
<< m1 >>
rect 353 439 354 440 
<< m1 >>
rect 354 439 355 440 
<< m1 >>
rect 355 439 356 440 
<< m1 >>
rect 356 439 357 440 
<< m1 >>
rect 357 439 358 440 
<< m1 >>
rect 358 439 359 440 
<< m1 >>
rect 359 439 360 440 
<< m1 >>
rect 360 439 361 440 
<< m1 >>
rect 361 439 362 440 
<< m2 >>
rect 361 439 362 440 
<< m1 >>
rect 362 439 363 440 
<< m1 >>
rect 363 439 364 440 
<< m1 >>
rect 364 439 365 440 
<< m1 >>
rect 365 439 366 440 
<< m1 >>
rect 366 439 367 440 
<< m1 >>
rect 367 439 368 440 
<< m1 >>
rect 368 439 369 440 
<< m1 >>
rect 369 439 370 440 
<< m1 >>
rect 370 439 371 440 
<< m1 >>
rect 371 439 372 440 
<< m1 >>
rect 372 439 373 440 
<< m1 >>
rect 373 439 374 440 
<< m1 >>
rect 374 439 375 440 
<< m1 >>
rect 375 439 376 440 
<< m1 >>
rect 376 439 377 440 
<< m1 >>
rect 377 439 378 440 
<< m1 >>
rect 378 439 379 440 
<< m1 >>
rect 379 439 380 440 
<< m2 >>
rect 379 439 380 440 
<< m1 >>
rect 380 439 381 440 
<< m1 >>
rect 381 439 382 440 
<< m1 >>
rect 382 439 383 440 
<< m1 >>
rect 383 439 384 440 
<< m1 >>
rect 384 439 385 440 
<< m1 >>
rect 385 439 386 440 
<< m2 >>
rect 385 439 386 440 
<< m1 >>
rect 386 439 387 440 
<< m1 >>
rect 387 439 388 440 
<< m1 >>
rect 388 439 389 440 
<< m1 >>
rect 389 439 390 440 
<< m1 >>
rect 390 439 391 440 
<< m1 >>
rect 391 439 392 440 
<< m1 >>
rect 392 439 393 440 
<< m1 >>
rect 393 439 394 440 
<< m1 >>
rect 394 439 395 440 
<< m1 >>
rect 395 439 396 440 
<< m1 >>
rect 396 439 397 440 
<< m1 >>
rect 397 439 398 440 
<< m2 >>
rect 397 439 398 440 
<< m1 >>
rect 398 439 399 440 
<< m1 >>
rect 399 439 400 440 
<< m1 >>
rect 400 439 401 440 
<< m2 >>
rect 400 439 401 440 
<< m1 >>
rect 401 439 402 440 
<< m1 >>
rect 402 439 403 440 
<< m2 >>
rect 402 439 403 440 
<< m1 >>
rect 403 439 404 440 
<< m1 >>
rect 404 439 405 440 
<< m1 >>
rect 405 439 406 440 
<< m1 >>
rect 406 439 407 440 
<< m2 >>
rect 406 439 407 440 
<< m1 >>
rect 407 439 408 440 
<< m1 >>
rect 408 439 409 440 
<< m1 >>
rect 409 439 410 440 
<< m1 >>
rect 410 439 411 440 
<< m1 >>
rect 411 439 412 440 
<< m1 >>
rect 412 439 413 440 
<< m1 >>
rect 413 439 414 440 
<< m1 >>
rect 414 439 415 440 
<< m1 >>
rect 415 439 416 440 
<< m1 >>
rect 416 439 417 440 
<< m1 >>
rect 417 439 418 440 
<< m1 >>
rect 418 439 419 440 
<< m1 >>
rect 419 439 420 440 
<< m1 >>
rect 420 439 421 440 
<< m1 >>
rect 421 439 422 440 
<< m1 >>
rect 422 439 423 440 
<< m1 >>
rect 423 439 424 440 
<< m1 >>
rect 424 439 425 440 
<< m2 >>
rect 424 439 425 440 
<< m1 >>
rect 425 439 426 440 
<< m1 >>
rect 426 439 427 440 
<< m1 >>
rect 427 439 428 440 
<< m1 >>
rect 428 439 429 440 
<< m1 >>
rect 429 439 430 440 
<< m1 >>
rect 430 439 431 440 
<< m1 >>
rect 431 439 432 440 
<< m2 >>
rect 431 439 432 440 
<< m2c >>
rect 431 439 432 440 
<< m1 >>
rect 431 439 432 440 
<< m2 >>
rect 431 439 432 440 
<< m2 >>
rect 432 439 433 440 
<< m1 >>
rect 433 439 434 440 
<< m2 >>
rect 433 439 434 440 
<< m2 >>
rect 434 439 435 440 
<< m1 >>
rect 435 439 436 440 
<< m2 >>
rect 435 439 436 440 
<< m2c >>
rect 435 439 436 440 
<< m1 >>
rect 435 439 436 440 
<< m2 >>
rect 435 439 436 440 
<< m1 >>
rect 436 439 437 440 
<< m1 >>
rect 437 439 438 440 
<< m1 >>
rect 438 439 439 440 
<< m1 >>
rect 439 439 440 440 
<< m1 >>
rect 440 439 441 440 
<< m1 >>
rect 441 439 442 440 
<< m1 >>
rect 442 439 443 440 
<< m1 >>
rect 443 439 444 440 
<< m1 >>
rect 444 439 445 440 
<< m2 >>
rect 444 439 445 440 
<< m1 >>
rect 445 439 446 440 
<< m2 >>
rect 445 439 446 440 
<< m1 >>
rect 446 439 447 440 
<< m2 >>
rect 446 439 447 440 
<< m1 >>
rect 447 439 448 440 
<< m2 >>
rect 447 439 448 440 
<< m1 >>
rect 448 439 449 440 
<< m2 >>
rect 448 439 449 440 
<< m2 >>
rect 449 439 450 440 
<< m1 >>
rect 450 439 451 440 
<< m2 >>
rect 450 439 451 440 
<< m2c >>
rect 450 439 451 440 
<< m1 >>
rect 450 439 451 440 
<< m2 >>
rect 450 439 451 440 
<< m1 >>
rect 451 439 452 440 
<< m1 >>
rect 452 439 453 440 
<< m2 >>
rect 452 439 453 440 
<< m1 >>
rect 453 439 454 440 
<< m1 >>
rect 454 439 455 440 
<< m1 >>
rect 455 439 456 440 
<< m1 >>
rect 456 439 457 440 
<< m1 >>
rect 457 439 458 440 
<< m1 >>
rect 458 439 459 440 
<< m1 >>
rect 459 439 460 440 
<< m1 >>
rect 460 439 461 440 
<< m1 >>
rect 461 439 462 440 
<< m1 >>
rect 462 439 463 440 
<< m2 >>
rect 462 439 463 440 
<< m1 >>
rect 463 439 464 440 
<< m1 >>
rect 464 439 465 440 
<< m1 >>
rect 465 439 466 440 
<< m1 >>
rect 466 439 467 440 
<< m1 >>
rect 467 439 468 440 
<< m1 >>
rect 468 439 469 440 
<< m1 >>
rect 469 439 470 440 
<< m1 >>
rect 470 439 471 440 
<< m1 >>
rect 472 439 473 440 
<< m1 >>
rect 478 439 479 440 
<< m1 >>
rect 487 439 488 440 
<< m1 >>
rect 489 439 490 440 
<< m1 >>
rect 502 439 503 440 
<< m1 >>
rect 19 440 20 441 
<< m1 >>
rect 21 440 22 441 
<< m1 >>
rect 26 440 27 441 
<< m1 >>
rect 28 440 29 441 
<< m2 >>
rect 28 440 29 441 
<< m1 >>
rect 49 440 50 441 
<< m1 >>
rect 73 440 74 441 
<< m1 >>
rect 96 440 97 441 
<< m1 >>
rect 97 440 98 441 
<< m1 >>
rect 98 440 99 441 
<< m2 >>
rect 98 440 99 441 
<< m2c >>
rect 98 440 99 441 
<< m1 >>
rect 98 440 99 441 
<< m2 >>
rect 98 440 99 441 
<< m2 >>
rect 99 440 100 441 
<< m1 >>
rect 100 440 101 441 
<< m1 >>
rect 106 440 107 441 
<< m2 >>
rect 122 440 123 441 
<< m1 >>
rect 150 440 151 441 
<< m1 >>
rect 152 440 153 441 
<< m2 >>
rect 164 440 165 441 
<< m2 >>
rect 194 440 195 441 
<< m2 >>
rect 207 440 208 441 
<< m1 >>
rect 208 440 209 441 
<< m1 >>
rect 211 440 212 441 
<< m2 >>
rect 217 440 218 441 
<< m2 >>
rect 249 440 250 441 
<< m1 >>
rect 253 440 254 441 
<< m2 >>
rect 289 440 290 441 
<< m2 >>
rect 290 440 291 441 
<< m1 >>
rect 298 440 299 441 
<< m2 >>
rect 307 440 308 441 
<< m2 >>
rect 325 440 326 441 
<< m2 >>
rect 361 440 362 441 
<< m2 >>
rect 379 440 380 441 
<< m2 >>
rect 385 440 386 441 
<< m2 >>
rect 397 440 398 441 
<< m2 >>
rect 400 440 401 441 
<< m2 >>
rect 402 440 403 441 
<< m2 >>
rect 406 440 407 441 
<< m2 >>
rect 424 440 425 441 
<< m1 >>
rect 433 440 434 441 
<< m1 >>
rect 448 440 449 441 
<< m2 >>
rect 452 440 453 441 
<< m2 >>
rect 462 440 463 441 
<< m1 >>
rect 470 440 471 441 
<< m1 >>
rect 472 440 473 441 
<< m1 >>
rect 478 440 479 441 
<< m1 >>
rect 487 440 488 441 
<< m1 >>
rect 489 440 490 441 
<< m1 >>
rect 502 440 503 441 
<< m1 >>
rect 19 441 20 442 
<< m1 >>
rect 21 441 22 442 
<< m1 >>
rect 26 441 27 442 
<< m1 >>
rect 28 441 29 442 
<< m2 >>
rect 28 441 29 442 
<< m1 >>
rect 49 441 50 442 
<< m1 >>
rect 73 441 74 442 
<< m2 >>
rect 99 441 100 442 
<< m1 >>
rect 100 441 101 442 
<< m1 >>
rect 106 441 107 442 
<< m1 >>
rect 122 441 123 442 
<< m2 >>
rect 122 441 123 442 
<< m2c >>
rect 122 441 123 442 
<< m1 >>
rect 122 441 123 442 
<< m2 >>
rect 122 441 123 442 
<< m1 >>
rect 123 441 124 442 
<< m1 >>
rect 124 441 125 442 
<< m1 >>
rect 125 441 126 442 
<< m1 >>
rect 126 441 127 442 
<< m1 >>
rect 127 441 128 442 
<< m1 >>
rect 128 441 129 442 
<< m1 >>
rect 129 441 130 442 
<< m1 >>
rect 130 441 131 442 
<< m1 >>
rect 131 441 132 442 
<< m1 >>
rect 132 441 133 442 
<< m1 >>
rect 133 441 134 442 
<< m1 >>
rect 134 441 135 442 
<< m1 >>
rect 135 441 136 442 
<< m1 >>
rect 136 441 137 442 
<< m1 >>
rect 137 441 138 442 
<< m1 >>
rect 138 441 139 442 
<< m1 >>
rect 139 441 140 442 
<< m1 >>
rect 140 441 141 442 
<< m1 >>
rect 141 441 142 442 
<< m1 >>
rect 142 441 143 442 
<< m1 >>
rect 143 441 144 442 
<< m1 >>
rect 144 441 145 442 
<< m1 >>
rect 145 441 146 442 
<< m1 >>
rect 146 441 147 442 
<< m1 >>
rect 147 441 148 442 
<< m1 >>
rect 148 441 149 442 
<< m2 >>
rect 148 441 149 442 
<< m2c >>
rect 148 441 149 442 
<< m1 >>
rect 148 441 149 442 
<< m2 >>
rect 148 441 149 442 
<< m2 >>
rect 149 441 150 442 
<< m1 >>
rect 150 441 151 442 
<< m2 >>
rect 150 441 151 442 
<< m2 >>
rect 151 441 152 442 
<< m1 >>
rect 152 441 153 442 
<< m2 >>
rect 152 441 153 442 
<< m2 >>
rect 153 441 154 442 
<< m1 >>
rect 154 441 155 442 
<< m2 >>
rect 154 441 155 442 
<< m2c >>
rect 154 441 155 442 
<< m1 >>
rect 154 441 155 442 
<< m2 >>
rect 154 441 155 442 
<< m2 >>
rect 164 441 165 442 
<< m1 >>
rect 193 441 194 442 
<< m1 >>
rect 194 441 195 442 
<< m2 >>
rect 194 441 195 442 
<< m1 >>
rect 195 441 196 442 
<< m2 >>
rect 195 441 196 442 
<< m1 >>
rect 196 441 197 442 
<< m2 >>
rect 196 441 197 442 
<< m1 >>
rect 197 441 198 442 
<< m2 >>
rect 197 441 198 442 
<< m1 >>
rect 198 441 199 442 
<< m2 >>
rect 198 441 199 442 
<< m1 >>
rect 199 441 200 442 
<< m2 >>
rect 199 441 200 442 
<< m1 >>
rect 200 441 201 442 
<< m2 >>
rect 200 441 201 442 
<< m1 >>
rect 201 441 202 442 
<< m2 >>
rect 201 441 202 442 
<< m1 >>
rect 202 441 203 442 
<< m2 >>
rect 202 441 203 442 
<< m1 >>
rect 203 441 204 442 
<< m2 >>
rect 203 441 204 442 
<< m1 >>
rect 204 441 205 442 
<< m2 >>
rect 204 441 205 442 
<< m1 >>
rect 205 441 206 442 
<< m1 >>
rect 206 441 207 442 
<< m2 >>
rect 206 441 207 442 
<< m2c >>
rect 206 441 207 442 
<< m1 >>
rect 206 441 207 442 
<< m2 >>
rect 206 441 207 442 
<< m2 >>
rect 207 441 208 442 
<< m1 >>
rect 208 441 209 442 
<< m1 >>
rect 211 441 212 442 
<< m1 >>
rect 217 441 218 442 
<< m2 >>
rect 217 441 218 442 
<< m2c >>
rect 217 441 218 442 
<< m1 >>
rect 217 441 218 442 
<< m2 >>
rect 217 441 218 442 
<< m1 >>
rect 249 441 250 442 
<< m2 >>
rect 249 441 250 442 
<< m2c >>
rect 249 441 250 442 
<< m1 >>
rect 249 441 250 442 
<< m2 >>
rect 249 441 250 442 
<< m1 >>
rect 250 441 251 442 
<< m1 >>
rect 251 441 252 442 
<< m1 >>
rect 253 441 254 442 
<< m1 >>
rect 289 441 290 442 
<< m2 >>
rect 289 441 290 442 
<< m2c >>
rect 289 441 290 442 
<< m1 >>
rect 289 441 290 442 
<< m2 >>
rect 289 441 290 442 
<< m1 >>
rect 298 441 299 442 
<< m1 >>
rect 307 441 308 442 
<< m2 >>
rect 307 441 308 442 
<< m2c >>
rect 307 441 308 442 
<< m1 >>
rect 307 441 308 442 
<< m2 >>
rect 307 441 308 442 
<< m1 >>
rect 325 441 326 442 
<< m2 >>
rect 325 441 326 442 
<< m2c >>
rect 325 441 326 442 
<< m1 >>
rect 325 441 326 442 
<< m2 >>
rect 325 441 326 442 
<< m1 >>
rect 361 441 362 442 
<< m2 >>
rect 361 441 362 442 
<< m2c >>
rect 361 441 362 442 
<< m1 >>
rect 361 441 362 442 
<< m2 >>
rect 361 441 362 442 
<< m1 >>
rect 379 441 380 442 
<< m2 >>
rect 379 441 380 442 
<< m2c >>
rect 379 441 380 442 
<< m1 >>
rect 379 441 380 442 
<< m2 >>
rect 379 441 380 442 
<< m1 >>
rect 380 441 381 442 
<< m1 >>
rect 381 441 382 442 
<< m2 >>
rect 385 441 386 442 
<< m1 >>
rect 397 441 398 442 
<< m2 >>
rect 397 441 398 442 
<< m2c >>
rect 397 441 398 442 
<< m1 >>
rect 397 441 398 442 
<< m2 >>
rect 397 441 398 442 
<< m1 >>
rect 400 441 401 442 
<< m2 >>
rect 400 441 401 442 
<< m2c >>
rect 400 441 401 442 
<< m1 >>
rect 400 441 401 442 
<< m2 >>
rect 400 441 401 442 
<< m1 >>
rect 402 441 403 442 
<< m2 >>
rect 402 441 403 442 
<< m2c >>
rect 402 441 403 442 
<< m1 >>
rect 402 441 403 442 
<< m2 >>
rect 402 441 403 442 
<< m1 >>
rect 406 441 407 442 
<< m2 >>
rect 406 441 407 442 
<< m2c >>
rect 406 441 407 442 
<< m1 >>
rect 406 441 407 442 
<< m2 >>
rect 406 441 407 442 
<< m1 >>
rect 424 441 425 442 
<< m2 >>
rect 424 441 425 442 
<< m2c >>
rect 424 441 425 442 
<< m1 >>
rect 424 441 425 442 
<< m2 >>
rect 424 441 425 442 
<< m1 >>
rect 433 441 434 442 
<< m1 >>
rect 448 441 449 442 
<< m1 >>
rect 452 441 453 442 
<< m2 >>
rect 452 441 453 442 
<< m2c >>
rect 452 441 453 442 
<< m1 >>
rect 452 441 453 442 
<< m2 >>
rect 452 441 453 442 
<< m1 >>
rect 460 441 461 442 
<< m1 >>
rect 461 441 462 442 
<< m1 >>
rect 462 441 463 442 
<< m2 >>
rect 462 441 463 442 
<< m2c >>
rect 462 441 463 442 
<< m1 >>
rect 462 441 463 442 
<< m2 >>
rect 462 441 463 442 
<< m1 >>
rect 470 441 471 442 
<< m1 >>
rect 472 441 473 442 
<< m1 >>
rect 478 441 479 442 
<< m1 >>
rect 487 441 488 442 
<< m1 >>
rect 489 441 490 442 
<< m1 >>
rect 502 441 503 442 
<< m1 >>
rect 19 442 20 443 
<< m1 >>
rect 21 442 22 443 
<< m1 >>
rect 26 442 27 443 
<< m1 >>
rect 28 442 29 443 
<< m2 >>
rect 28 442 29 443 
<< m1 >>
rect 49 442 50 443 
<< m1 >>
rect 55 442 56 443 
<< m1 >>
rect 56 442 57 443 
<< m1 >>
rect 57 442 58 443 
<< m1 >>
rect 58 442 59 443 
<< m1 >>
rect 59 442 60 443 
<< m1 >>
rect 60 442 61 443 
<< m1 >>
rect 61 442 62 443 
<< m1 >>
rect 62 442 63 443 
<< m1 >>
rect 63 442 64 443 
<< m1 >>
rect 64 442 65 443 
<< m1 >>
rect 65 442 66 443 
<< m1 >>
rect 66 442 67 443 
<< m1 >>
rect 67 442 68 443 
<< m1 >>
rect 73 442 74 443 
<< m2 >>
rect 99 442 100 443 
<< m1 >>
rect 100 442 101 443 
<< m1 >>
rect 106 442 107 443 
<< m1 >>
rect 150 442 151 443 
<< m1 >>
rect 152 442 153 443 
<< m1 >>
rect 154 442 155 443 
<< m1 >>
rect 160 442 161 443 
<< m1 >>
rect 161 442 162 443 
<< m1 >>
rect 162 442 163 443 
<< m1 >>
rect 163 442 164 443 
<< m1 >>
rect 164 442 165 443 
<< m2 >>
rect 164 442 165 443 
<< m1 >>
rect 165 442 166 443 
<< m1 >>
rect 166 442 167 443 
<< m1 >>
rect 167 442 168 443 
<< m1 >>
rect 168 442 169 443 
<< m1 >>
rect 169 442 170 443 
<< m1 >>
rect 170 442 171 443 
<< m1 >>
rect 172 442 173 443 
<< m1 >>
rect 173 442 174 443 
<< m1 >>
rect 174 442 175 443 
<< m1 >>
rect 175 442 176 443 
<< m1 >>
rect 193 442 194 443 
<< m2 >>
rect 204 442 205 443 
<< m1 >>
rect 208 442 209 443 
<< m1 >>
rect 211 442 212 443 
<< m1 >>
rect 217 442 218 443 
<< m1 >>
rect 251 442 252 443 
<< m2 >>
rect 251 442 252 443 
<< m2c >>
rect 251 442 252 443 
<< m1 >>
rect 251 442 252 443 
<< m2 >>
rect 251 442 252 443 
<< m2 >>
rect 252 442 253 443 
<< m1 >>
rect 253 442 254 443 
<< m2 >>
rect 253 442 254 443 
<< m2 >>
rect 254 442 255 443 
<< m1 >>
rect 289 442 290 443 
<< m1 >>
rect 298 442 299 443 
<< m1 >>
rect 307 442 308 443 
<< m1 >>
rect 325 442 326 443 
<< m1 >>
rect 361 442 362 443 
<< m1 >>
rect 381 442 382 443 
<< m2 >>
rect 382 442 383 443 
<< m1 >>
rect 383 442 384 443 
<< m2 >>
rect 383 442 384 443 
<< m2c >>
rect 383 442 384 443 
<< m1 >>
rect 383 442 384 443 
<< m2 >>
rect 383 442 384 443 
<< m1 >>
rect 384 442 385 443 
<< m1 >>
rect 385 442 386 443 
<< m2 >>
rect 385 442 386 443 
<< m1 >>
rect 386 442 387 443 
<< m1 >>
rect 387 442 388 443 
<< m1 >>
rect 388 442 389 443 
<< m1 >>
rect 389 442 390 443 
<< m1 >>
rect 390 442 391 443 
<< m1 >>
rect 391 442 392 443 
<< m1 >>
rect 397 442 398 443 
<< m1 >>
rect 400 442 401 443 
<< m1 >>
rect 402 442 403 443 
<< m1 >>
rect 406 442 407 443 
<< m1 >>
rect 424 442 425 443 
<< m1 >>
rect 433 442 434 443 
<< m2 >>
rect 434 442 435 443 
<< m1 >>
rect 435 442 436 443 
<< m2 >>
rect 435 442 436 443 
<< m2c >>
rect 435 442 436 443 
<< m1 >>
rect 435 442 436 443 
<< m2 >>
rect 435 442 436 443 
<< m1 >>
rect 436 442 437 443 
<< m1 >>
rect 437 442 438 443 
<< m1 >>
rect 438 442 439 443 
<< m1 >>
rect 439 442 440 443 
<< m1 >>
rect 440 442 441 443 
<< m1 >>
rect 441 442 442 443 
<< m1 >>
rect 442 442 443 443 
<< m1 >>
rect 443 442 444 443 
<< m1 >>
rect 444 442 445 443 
<< m1 >>
rect 445 442 446 443 
<< m1 >>
rect 448 442 449 443 
<< m1 >>
rect 452 442 453 443 
<< m1 >>
rect 460 442 461 443 
<< m1 >>
rect 470 442 471 443 
<< m1 >>
rect 472 442 473 443 
<< m1 >>
rect 478 442 479 443 
<< m1 >>
rect 487 442 488 443 
<< m1 >>
rect 489 442 490 443 
<< m1 >>
rect 502 442 503 443 
<< m1 >>
rect 19 443 20 444 
<< m1 >>
rect 21 443 22 444 
<< m1 >>
rect 26 443 27 444 
<< m1 >>
rect 28 443 29 444 
<< m2 >>
rect 28 443 29 444 
<< m1 >>
rect 49 443 50 444 
<< m1 >>
rect 55 443 56 444 
<< m1 >>
rect 67 443 68 444 
<< m1 >>
rect 73 443 74 444 
<< m2 >>
rect 99 443 100 444 
<< m1 >>
rect 100 443 101 444 
<< m1 >>
rect 106 443 107 444 
<< m1 >>
rect 150 443 151 444 
<< m1 >>
rect 152 443 153 444 
<< m1 >>
rect 154 443 155 444 
<< m1 >>
rect 160 443 161 444 
<< m2 >>
rect 163 443 164 444 
<< m2 >>
rect 164 443 165 444 
<< m1 >>
rect 170 443 171 444 
<< m1 >>
rect 172 443 173 444 
<< m1 >>
rect 175 443 176 444 
<< m1 >>
rect 193 443 194 444 
<< m1 >>
rect 204 443 205 444 
<< m2 >>
rect 204 443 205 444 
<< m2c >>
rect 204 443 205 444 
<< m1 >>
rect 204 443 205 444 
<< m2 >>
rect 204 443 205 444 
<< m1 >>
rect 208 443 209 444 
<< m1 >>
rect 211 443 212 444 
<< m1 >>
rect 217 443 218 444 
<< m1 >>
rect 253 443 254 444 
<< m2 >>
rect 254 443 255 444 
<< m1 >>
rect 289 443 290 444 
<< m1 >>
rect 298 443 299 444 
<< m1 >>
rect 307 443 308 444 
<< m1 >>
rect 325 443 326 444 
<< m1 >>
rect 361 443 362 444 
<< m1 >>
rect 379 443 380 444 
<< m2 >>
rect 379 443 380 444 
<< m2c >>
rect 379 443 380 444 
<< m1 >>
rect 379 443 380 444 
<< m2 >>
rect 379 443 380 444 
<< m2 >>
rect 380 443 381 444 
<< m1 >>
rect 381 443 382 444 
<< m2 >>
rect 381 443 382 444 
<< m2 >>
rect 382 443 383 444 
<< m2 >>
rect 385 443 386 444 
<< m1 >>
rect 391 443 392 444 
<< m1 >>
rect 397 443 398 444 
<< m1 >>
rect 400 443 401 444 
<< m1 >>
rect 402 443 403 444 
<< m1 >>
rect 406 443 407 444 
<< m1 >>
rect 424 443 425 444 
<< m1 >>
rect 433 443 434 444 
<< m2 >>
rect 434 443 435 444 
<< m1 >>
rect 445 443 446 444 
<< m1 >>
rect 448 443 449 444 
<< m1 >>
rect 452 443 453 444 
<< m2 >>
rect 453 443 454 444 
<< m1 >>
rect 454 443 455 444 
<< m2 >>
rect 454 443 455 444 
<< m2c >>
rect 454 443 455 444 
<< m1 >>
rect 454 443 455 444 
<< m2 >>
rect 454 443 455 444 
<< m1 >>
rect 455 443 456 444 
<< m1 >>
rect 456 443 457 444 
<< m1 >>
rect 457 443 458 444 
<< m1 >>
rect 458 443 459 444 
<< m1 >>
rect 459 443 460 444 
<< m1 >>
rect 460 443 461 444 
<< m1 >>
rect 470 443 471 444 
<< m1 >>
rect 472 443 473 444 
<< m1 >>
rect 478 443 479 444 
<< m1 >>
rect 487 443 488 444 
<< m1 >>
rect 489 443 490 444 
<< m1 >>
rect 502 443 503 444 
<< pdiffusion >>
rect 12 444 13 445 
<< pdiffusion >>
rect 13 444 14 445 
<< pdiffusion >>
rect 14 444 15 445 
<< pdiffusion >>
rect 15 444 16 445 
<< pdiffusion >>
rect 16 444 17 445 
<< pdiffusion >>
rect 17 444 18 445 
<< m1 >>
rect 19 444 20 445 
<< m1 >>
rect 21 444 22 445 
<< m1 >>
rect 26 444 27 445 
<< m1 >>
rect 28 444 29 445 
<< m2 >>
rect 28 444 29 445 
<< pdiffusion >>
rect 30 444 31 445 
<< pdiffusion >>
rect 31 444 32 445 
<< pdiffusion >>
rect 32 444 33 445 
<< pdiffusion >>
rect 33 444 34 445 
<< pdiffusion >>
rect 34 444 35 445 
<< pdiffusion >>
rect 35 444 36 445 
<< pdiffusion >>
rect 48 444 49 445 
<< m1 >>
rect 49 444 50 445 
<< pdiffusion >>
rect 49 444 50 445 
<< pdiffusion >>
rect 50 444 51 445 
<< pdiffusion >>
rect 51 444 52 445 
<< pdiffusion >>
rect 52 444 53 445 
<< pdiffusion >>
rect 53 444 54 445 
<< m1 >>
rect 55 444 56 445 
<< pdiffusion >>
rect 66 444 67 445 
<< m1 >>
rect 67 444 68 445 
<< pdiffusion >>
rect 67 444 68 445 
<< pdiffusion >>
rect 68 444 69 445 
<< pdiffusion >>
rect 69 444 70 445 
<< pdiffusion >>
rect 70 444 71 445 
<< pdiffusion >>
rect 71 444 72 445 
<< m1 >>
rect 73 444 74 445 
<< pdiffusion >>
rect 84 444 85 445 
<< pdiffusion >>
rect 85 444 86 445 
<< pdiffusion >>
rect 86 444 87 445 
<< pdiffusion >>
rect 87 444 88 445 
<< pdiffusion >>
rect 88 444 89 445 
<< pdiffusion >>
rect 89 444 90 445 
<< m2 >>
rect 99 444 100 445 
<< m1 >>
rect 100 444 101 445 
<< pdiffusion >>
rect 102 444 103 445 
<< pdiffusion >>
rect 103 444 104 445 
<< pdiffusion >>
rect 104 444 105 445 
<< pdiffusion >>
rect 105 444 106 445 
<< m1 >>
rect 106 444 107 445 
<< pdiffusion >>
rect 106 444 107 445 
<< pdiffusion >>
rect 107 444 108 445 
<< pdiffusion >>
rect 120 444 121 445 
<< pdiffusion >>
rect 121 444 122 445 
<< pdiffusion >>
rect 122 444 123 445 
<< pdiffusion >>
rect 123 444 124 445 
<< pdiffusion >>
rect 124 444 125 445 
<< pdiffusion >>
rect 125 444 126 445 
<< m1 >>
rect 150 444 151 445 
<< m1 >>
rect 152 444 153 445 
<< m1 >>
rect 154 444 155 445 
<< pdiffusion >>
rect 156 444 157 445 
<< pdiffusion >>
rect 157 444 158 445 
<< pdiffusion >>
rect 158 444 159 445 
<< pdiffusion >>
rect 159 444 160 445 
<< m1 >>
rect 160 444 161 445 
<< pdiffusion >>
rect 160 444 161 445 
<< pdiffusion >>
rect 161 444 162 445 
<< m1 >>
rect 163 444 164 445 
<< m2 >>
rect 163 444 164 445 
<< m2c >>
rect 163 444 164 445 
<< m1 >>
rect 163 444 164 445 
<< m2 >>
rect 163 444 164 445 
<< m1 >>
rect 170 444 171 445 
<< m1 >>
rect 172 444 173 445 
<< pdiffusion >>
rect 174 444 175 445 
<< m1 >>
rect 175 444 176 445 
<< pdiffusion >>
rect 175 444 176 445 
<< pdiffusion >>
rect 176 444 177 445 
<< pdiffusion >>
rect 177 444 178 445 
<< pdiffusion >>
rect 178 444 179 445 
<< pdiffusion >>
rect 179 444 180 445 
<< pdiffusion >>
rect 192 444 193 445 
<< m1 >>
rect 193 444 194 445 
<< pdiffusion >>
rect 193 444 194 445 
<< pdiffusion >>
rect 194 444 195 445 
<< pdiffusion >>
rect 195 444 196 445 
<< pdiffusion >>
rect 196 444 197 445 
<< pdiffusion >>
rect 197 444 198 445 
<< m1 >>
rect 204 444 205 445 
<< m1 >>
rect 208 444 209 445 
<< pdiffusion >>
rect 210 444 211 445 
<< m1 >>
rect 211 444 212 445 
<< pdiffusion >>
rect 211 444 212 445 
<< pdiffusion >>
rect 212 444 213 445 
<< pdiffusion >>
rect 213 444 214 445 
<< pdiffusion >>
rect 214 444 215 445 
<< pdiffusion >>
rect 215 444 216 445 
<< m1 >>
rect 217 444 218 445 
<< pdiffusion >>
rect 228 444 229 445 
<< pdiffusion >>
rect 229 444 230 445 
<< pdiffusion >>
rect 230 444 231 445 
<< pdiffusion >>
rect 231 444 232 445 
<< pdiffusion >>
rect 232 444 233 445 
<< pdiffusion >>
rect 233 444 234 445 
<< pdiffusion >>
rect 246 444 247 445 
<< pdiffusion >>
rect 247 444 248 445 
<< pdiffusion >>
rect 248 444 249 445 
<< pdiffusion >>
rect 249 444 250 445 
<< pdiffusion >>
rect 250 444 251 445 
<< pdiffusion >>
rect 251 444 252 445 
<< m1 >>
rect 253 444 254 445 
<< m2 >>
rect 254 444 255 445 
<< pdiffusion >>
rect 264 444 265 445 
<< pdiffusion >>
rect 265 444 266 445 
<< pdiffusion >>
rect 266 444 267 445 
<< pdiffusion >>
rect 267 444 268 445 
<< pdiffusion >>
rect 268 444 269 445 
<< pdiffusion >>
rect 269 444 270 445 
<< pdiffusion >>
rect 282 444 283 445 
<< pdiffusion >>
rect 283 444 284 445 
<< pdiffusion >>
rect 284 444 285 445 
<< pdiffusion >>
rect 285 444 286 445 
<< pdiffusion >>
rect 286 444 287 445 
<< pdiffusion >>
rect 287 444 288 445 
<< m1 >>
rect 289 444 290 445 
<< m1 >>
rect 298 444 299 445 
<< pdiffusion >>
rect 300 444 301 445 
<< pdiffusion >>
rect 301 444 302 445 
<< pdiffusion >>
rect 302 444 303 445 
<< pdiffusion >>
rect 303 444 304 445 
<< pdiffusion >>
rect 304 444 305 445 
<< pdiffusion >>
rect 305 444 306 445 
<< m1 >>
rect 307 444 308 445 
<< pdiffusion >>
rect 318 444 319 445 
<< pdiffusion >>
rect 319 444 320 445 
<< pdiffusion >>
rect 320 444 321 445 
<< pdiffusion >>
rect 321 444 322 445 
<< pdiffusion >>
rect 322 444 323 445 
<< pdiffusion >>
rect 323 444 324 445 
<< m1 >>
rect 325 444 326 445 
<< pdiffusion >>
rect 336 444 337 445 
<< pdiffusion >>
rect 337 444 338 445 
<< pdiffusion >>
rect 338 444 339 445 
<< pdiffusion >>
rect 339 444 340 445 
<< pdiffusion >>
rect 340 444 341 445 
<< pdiffusion >>
rect 341 444 342 445 
<< pdiffusion >>
rect 354 444 355 445 
<< pdiffusion >>
rect 355 444 356 445 
<< pdiffusion >>
rect 356 444 357 445 
<< pdiffusion >>
rect 357 444 358 445 
<< pdiffusion >>
rect 358 444 359 445 
<< pdiffusion >>
rect 359 444 360 445 
<< m1 >>
rect 361 444 362 445 
<< pdiffusion >>
rect 372 444 373 445 
<< pdiffusion >>
rect 373 444 374 445 
<< pdiffusion >>
rect 374 444 375 445 
<< pdiffusion >>
rect 375 444 376 445 
<< pdiffusion >>
rect 376 444 377 445 
<< pdiffusion >>
rect 377 444 378 445 
<< m1 >>
rect 379 444 380 445 
<< m1 >>
rect 381 444 382 445 
<< m1 >>
rect 385 444 386 445 
<< m2 >>
rect 385 444 386 445 
<< m2c >>
rect 385 444 386 445 
<< m1 >>
rect 385 444 386 445 
<< m2 >>
rect 385 444 386 445 
<< pdiffusion >>
rect 390 444 391 445 
<< m1 >>
rect 391 444 392 445 
<< pdiffusion >>
rect 391 444 392 445 
<< pdiffusion >>
rect 392 444 393 445 
<< pdiffusion >>
rect 393 444 394 445 
<< pdiffusion >>
rect 394 444 395 445 
<< pdiffusion >>
rect 395 444 396 445 
<< m1 >>
rect 397 444 398 445 
<< m1 >>
rect 400 444 401 445 
<< m1 >>
rect 402 444 403 445 
<< m1 >>
rect 406 444 407 445 
<< pdiffusion >>
rect 408 444 409 445 
<< pdiffusion >>
rect 409 444 410 445 
<< pdiffusion >>
rect 410 444 411 445 
<< pdiffusion >>
rect 411 444 412 445 
<< pdiffusion >>
rect 412 444 413 445 
<< pdiffusion >>
rect 413 444 414 445 
<< m1 >>
rect 424 444 425 445 
<< pdiffusion >>
rect 426 444 427 445 
<< pdiffusion >>
rect 427 444 428 445 
<< pdiffusion >>
rect 428 444 429 445 
<< pdiffusion >>
rect 429 444 430 445 
<< pdiffusion >>
rect 430 444 431 445 
<< pdiffusion >>
rect 431 444 432 445 
<< m1 >>
rect 433 444 434 445 
<< m2 >>
rect 434 444 435 445 
<< pdiffusion >>
rect 444 444 445 445 
<< m1 >>
rect 445 444 446 445 
<< pdiffusion >>
rect 445 444 446 445 
<< pdiffusion >>
rect 446 444 447 445 
<< pdiffusion >>
rect 447 444 448 445 
<< m1 >>
rect 448 444 449 445 
<< pdiffusion >>
rect 448 444 449 445 
<< pdiffusion >>
rect 449 444 450 445 
<< m1 >>
rect 452 444 453 445 
<< m2 >>
rect 453 444 454 445 
<< pdiffusion >>
rect 462 444 463 445 
<< pdiffusion >>
rect 463 444 464 445 
<< pdiffusion >>
rect 464 444 465 445 
<< pdiffusion >>
rect 465 444 466 445 
<< pdiffusion >>
rect 466 444 467 445 
<< pdiffusion >>
rect 467 444 468 445 
<< m1 >>
rect 470 444 471 445 
<< m1 >>
rect 472 444 473 445 
<< m1 >>
rect 478 444 479 445 
<< pdiffusion >>
rect 480 444 481 445 
<< pdiffusion >>
rect 481 444 482 445 
<< pdiffusion >>
rect 482 444 483 445 
<< pdiffusion >>
rect 483 444 484 445 
<< pdiffusion >>
rect 484 444 485 445 
<< pdiffusion >>
rect 485 444 486 445 
<< m1 >>
rect 487 444 488 445 
<< m1 >>
rect 489 444 490 445 
<< pdiffusion >>
rect 498 444 499 445 
<< pdiffusion >>
rect 499 444 500 445 
<< pdiffusion >>
rect 500 444 501 445 
<< pdiffusion >>
rect 501 444 502 445 
<< m1 >>
rect 502 444 503 445 
<< pdiffusion >>
rect 502 444 503 445 
<< pdiffusion >>
rect 503 444 504 445 
<< pdiffusion >>
rect 516 444 517 445 
<< pdiffusion >>
rect 517 444 518 445 
<< pdiffusion >>
rect 518 444 519 445 
<< pdiffusion >>
rect 519 444 520 445 
<< pdiffusion >>
rect 520 444 521 445 
<< pdiffusion >>
rect 521 444 522 445 
<< pdiffusion >>
rect 12 445 13 446 
<< pdiffusion >>
rect 13 445 14 446 
<< pdiffusion >>
rect 14 445 15 446 
<< pdiffusion >>
rect 15 445 16 446 
<< pdiffusion >>
rect 16 445 17 446 
<< pdiffusion >>
rect 17 445 18 446 
<< m1 >>
rect 19 445 20 446 
<< m1 >>
rect 21 445 22 446 
<< m1 >>
rect 26 445 27 446 
<< m1 >>
rect 28 445 29 446 
<< m2 >>
rect 28 445 29 446 
<< pdiffusion >>
rect 30 445 31 446 
<< pdiffusion >>
rect 31 445 32 446 
<< pdiffusion >>
rect 32 445 33 446 
<< pdiffusion >>
rect 33 445 34 446 
<< pdiffusion >>
rect 34 445 35 446 
<< pdiffusion >>
rect 35 445 36 446 
<< pdiffusion >>
rect 48 445 49 446 
<< pdiffusion >>
rect 49 445 50 446 
<< pdiffusion >>
rect 50 445 51 446 
<< pdiffusion >>
rect 51 445 52 446 
<< pdiffusion >>
rect 52 445 53 446 
<< pdiffusion >>
rect 53 445 54 446 
<< m1 >>
rect 55 445 56 446 
<< pdiffusion >>
rect 66 445 67 446 
<< pdiffusion >>
rect 67 445 68 446 
<< pdiffusion >>
rect 68 445 69 446 
<< pdiffusion >>
rect 69 445 70 446 
<< pdiffusion >>
rect 70 445 71 446 
<< pdiffusion >>
rect 71 445 72 446 
<< m1 >>
rect 73 445 74 446 
<< pdiffusion >>
rect 84 445 85 446 
<< pdiffusion >>
rect 85 445 86 446 
<< pdiffusion >>
rect 86 445 87 446 
<< pdiffusion >>
rect 87 445 88 446 
<< pdiffusion >>
rect 88 445 89 446 
<< pdiffusion >>
rect 89 445 90 446 
<< m2 >>
rect 99 445 100 446 
<< m1 >>
rect 100 445 101 446 
<< pdiffusion >>
rect 102 445 103 446 
<< pdiffusion >>
rect 103 445 104 446 
<< pdiffusion >>
rect 104 445 105 446 
<< pdiffusion >>
rect 105 445 106 446 
<< pdiffusion >>
rect 106 445 107 446 
<< pdiffusion >>
rect 107 445 108 446 
<< pdiffusion >>
rect 120 445 121 446 
<< pdiffusion >>
rect 121 445 122 446 
<< pdiffusion >>
rect 122 445 123 446 
<< pdiffusion >>
rect 123 445 124 446 
<< pdiffusion >>
rect 124 445 125 446 
<< pdiffusion >>
rect 125 445 126 446 
<< m1 >>
rect 150 445 151 446 
<< m1 >>
rect 152 445 153 446 
<< m1 >>
rect 154 445 155 446 
<< pdiffusion >>
rect 156 445 157 446 
<< pdiffusion >>
rect 157 445 158 446 
<< pdiffusion >>
rect 158 445 159 446 
<< pdiffusion >>
rect 159 445 160 446 
<< pdiffusion >>
rect 160 445 161 446 
<< pdiffusion >>
rect 161 445 162 446 
<< m1 >>
rect 163 445 164 446 
<< m1 >>
rect 170 445 171 446 
<< m1 >>
rect 172 445 173 446 
<< pdiffusion >>
rect 174 445 175 446 
<< pdiffusion >>
rect 175 445 176 446 
<< pdiffusion >>
rect 176 445 177 446 
<< pdiffusion >>
rect 177 445 178 446 
<< pdiffusion >>
rect 178 445 179 446 
<< pdiffusion >>
rect 179 445 180 446 
<< pdiffusion >>
rect 192 445 193 446 
<< pdiffusion >>
rect 193 445 194 446 
<< pdiffusion >>
rect 194 445 195 446 
<< pdiffusion >>
rect 195 445 196 446 
<< pdiffusion >>
rect 196 445 197 446 
<< pdiffusion >>
rect 197 445 198 446 
<< m1 >>
rect 204 445 205 446 
<< m1 >>
rect 208 445 209 446 
<< pdiffusion >>
rect 210 445 211 446 
<< pdiffusion >>
rect 211 445 212 446 
<< pdiffusion >>
rect 212 445 213 446 
<< pdiffusion >>
rect 213 445 214 446 
<< pdiffusion >>
rect 214 445 215 446 
<< pdiffusion >>
rect 215 445 216 446 
<< m1 >>
rect 217 445 218 446 
<< pdiffusion >>
rect 228 445 229 446 
<< pdiffusion >>
rect 229 445 230 446 
<< pdiffusion >>
rect 230 445 231 446 
<< pdiffusion >>
rect 231 445 232 446 
<< pdiffusion >>
rect 232 445 233 446 
<< pdiffusion >>
rect 233 445 234 446 
<< pdiffusion >>
rect 246 445 247 446 
<< pdiffusion >>
rect 247 445 248 446 
<< pdiffusion >>
rect 248 445 249 446 
<< pdiffusion >>
rect 249 445 250 446 
<< pdiffusion >>
rect 250 445 251 446 
<< pdiffusion >>
rect 251 445 252 446 
<< m1 >>
rect 253 445 254 446 
<< m2 >>
rect 254 445 255 446 
<< pdiffusion >>
rect 264 445 265 446 
<< pdiffusion >>
rect 265 445 266 446 
<< pdiffusion >>
rect 266 445 267 446 
<< pdiffusion >>
rect 267 445 268 446 
<< pdiffusion >>
rect 268 445 269 446 
<< pdiffusion >>
rect 269 445 270 446 
<< pdiffusion >>
rect 282 445 283 446 
<< pdiffusion >>
rect 283 445 284 446 
<< pdiffusion >>
rect 284 445 285 446 
<< pdiffusion >>
rect 285 445 286 446 
<< pdiffusion >>
rect 286 445 287 446 
<< pdiffusion >>
rect 287 445 288 446 
<< m1 >>
rect 289 445 290 446 
<< m1 >>
rect 298 445 299 446 
<< pdiffusion >>
rect 300 445 301 446 
<< pdiffusion >>
rect 301 445 302 446 
<< pdiffusion >>
rect 302 445 303 446 
<< pdiffusion >>
rect 303 445 304 446 
<< pdiffusion >>
rect 304 445 305 446 
<< pdiffusion >>
rect 305 445 306 446 
<< m1 >>
rect 307 445 308 446 
<< pdiffusion >>
rect 318 445 319 446 
<< pdiffusion >>
rect 319 445 320 446 
<< pdiffusion >>
rect 320 445 321 446 
<< pdiffusion >>
rect 321 445 322 446 
<< pdiffusion >>
rect 322 445 323 446 
<< pdiffusion >>
rect 323 445 324 446 
<< m1 >>
rect 325 445 326 446 
<< pdiffusion >>
rect 336 445 337 446 
<< pdiffusion >>
rect 337 445 338 446 
<< pdiffusion >>
rect 338 445 339 446 
<< pdiffusion >>
rect 339 445 340 446 
<< pdiffusion >>
rect 340 445 341 446 
<< pdiffusion >>
rect 341 445 342 446 
<< pdiffusion >>
rect 354 445 355 446 
<< pdiffusion >>
rect 355 445 356 446 
<< pdiffusion >>
rect 356 445 357 446 
<< pdiffusion >>
rect 357 445 358 446 
<< pdiffusion >>
rect 358 445 359 446 
<< pdiffusion >>
rect 359 445 360 446 
<< m1 >>
rect 361 445 362 446 
<< pdiffusion >>
rect 372 445 373 446 
<< pdiffusion >>
rect 373 445 374 446 
<< pdiffusion >>
rect 374 445 375 446 
<< pdiffusion >>
rect 375 445 376 446 
<< pdiffusion >>
rect 376 445 377 446 
<< pdiffusion >>
rect 377 445 378 446 
<< m1 >>
rect 379 445 380 446 
<< m1 >>
rect 381 445 382 446 
<< m1 >>
rect 385 445 386 446 
<< pdiffusion >>
rect 390 445 391 446 
<< pdiffusion >>
rect 391 445 392 446 
<< pdiffusion >>
rect 392 445 393 446 
<< pdiffusion >>
rect 393 445 394 446 
<< pdiffusion >>
rect 394 445 395 446 
<< pdiffusion >>
rect 395 445 396 446 
<< m1 >>
rect 397 445 398 446 
<< m1 >>
rect 400 445 401 446 
<< m1 >>
rect 402 445 403 446 
<< m1 >>
rect 406 445 407 446 
<< pdiffusion >>
rect 408 445 409 446 
<< pdiffusion >>
rect 409 445 410 446 
<< pdiffusion >>
rect 410 445 411 446 
<< pdiffusion >>
rect 411 445 412 446 
<< pdiffusion >>
rect 412 445 413 446 
<< pdiffusion >>
rect 413 445 414 446 
<< m1 >>
rect 424 445 425 446 
<< pdiffusion >>
rect 426 445 427 446 
<< pdiffusion >>
rect 427 445 428 446 
<< pdiffusion >>
rect 428 445 429 446 
<< pdiffusion >>
rect 429 445 430 446 
<< pdiffusion >>
rect 430 445 431 446 
<< pdiffusion >>
rect 431 445 432 446 
<< m1 >>
rect 433 445 434 446 
<< m2 >>
rect 434 445 435 446 
<< pdiffusion >>
rect 444 445 445 446 
<< pdiffusion >>
rect 445 445 446 446 
<< pdiffusion >>
rect 446 445 447 446 
<< pdiffusion >>
rect 447 445 448 446 
<< pdiffusion >>
rect 448 445 449 446 
<< pdiffusion >>
rect 449 445 450 446 
<< m1 >>
rect 452 445 453 446 
<< m2 >>
rect 453 445 454 446 
<< pdiffusion >>
rect 462 445 463 446 
<< pdiffusion >>
rect 463 445 464 446 
<< pdiffusion >>
rect 464 445 465 446 
<< pdiffusion >>
rect 465 445 466 446 
<< pdiffusion >>
rect 466 445 467 446 
<< pdiffusion >>
rect 467 445 468 446 
<< m1 >>
rect 470 445 471 446 
<< m1 >>
rect 472 445 473 446 
<< m1 >>
rect 478 445 479 446 
<< pdiffusion >>
rect 480 445 481 446 
<< pdiffusion >>
rect 481 445 482 446 
<< pdiffusion >>
rect 482 445 483 446 
<< pdiffusion >>
rect 483 445 484 446 
<< pdiffusion >>
rect 484 445 485 446 
<< pdiffusion >>
rect 485 445 486 446 
<< m1 >>
rect 487 445 488 446 
<< m1 >>
rect 489 445 490 446 
<< pdiffusion >>
rect 498 445 499 446 
<< pdiffusion >>
rect 499 445 500 446 
<< pdiffusion >>
rect 500 445 501 446 
<< pdiffusion >>
rect 501 445 502 446 
<< pdiffusion >>
rect 502 445 503 446 
<< pdiffusion >>
rect 503 445 504 446 
<< pdiffusion >>
rect 516 445 517 446 
<< pdiffusion >>
rect 517 445 518 446 
<< pdiffusion >>
rect 518 445 519 446 
<< pdiffusion >>
rect 519 445 520 446 
<< pdiffusion >>
rect 520 445 521 446 
<< pdiffusion >>
rect 521 445 522 446 
<< pdiffusion >>
rect 12 446 13 447 
<< pdiffusion >>
rect 13 446 14 447 
<< pdiffusion >>
rect 14 446 15 447 
<< pdiffusion >>
rect 15 446 16 447 
<< pdiffusion >>
rect 16 446 17 447 
<< pdiffusion >>
rect 17 446 18 447 
<< m1 >>
rect 19 446 20 447 
<< m1 >>
rect 21 446 22 447 
<< m1 >>
rect 26 446 27 447 
<< m1 >>
rect 28 446 29 447 
<< m2 >>
rect 28 446 29 447 
<< pdiffusion >>
rect 30 446 31 447 
<< pdiffusion >>
rect 31 446 32 447 
<< pdiffusion >>
rect 32 446 33 447 
<< pdiffusion >>
rect 33 446 34 447 
<< pdiffusion >>
rect 34 446 35 447 
<< pdiffusion >>
rect 35 446 36 447 
<< pdiffusion >>
rect 48 446 49 447 
<< pdiffusion >>
rect 49 446 50 447 
<< pdiffusion >>
rect 50 446 51 447 
<< pdiffusion >>
rect 51 446 52 447 
<< pdiffusion >>
rect 52 446 53 447 
<< pdiffusion >>
rect 53 446 54 447 
<< m1 >>
rect 55 446 56 447 
<< pdiffusion >>
rect 66 446 67 447 
<< pdiffusion >>
rect 67 446 68 447 
<< pdiffusion >>
rect 68 446 69 447 
<< pdiffusion >>
rect 69 446 70 447 
<< pdiffusion >>
rect 70 446 71 447 
<< pdiffusion >>
rect 71 446 72 447 
<< m1 >>
rect 73 446 74 447 
<< pdiffusion >>
rect 84 446 85 447 
<< pdiffusion >>
rect 85 446 86 447 
<< pdiffusion >>
rect 86 446 87 447 
<< pdiffusion >>
rect 87 446 88 447 
<< pdiffusion >>
rect 88 446 89 447 
<< pdiffusion >>
rect 89 446 90 447 
<< m2 >>
rect 99 446 100 447 
<< m1 >>
rect 100 446 101 447 
<< pdiffusion >>
rect 102 446 103 447 
<< pdiffusion >>
rect 103 446 104 447 
<< pdiffusion >>
rect 104 446 105 447 
<< pdiffusion >>
rect 105 446 106 447 
<< pdiffusion >>
rect 106 446 107 447 
<< pdiffusion >>
rect 107 446 108 447 
<< pdiffusion >>
rect 120 446 121 447 
<< pdiffusion >>
rect 121 446 122 447 
<< pdiffusion >>
rect 122 446 123 447 
<< pdiffusion >>
rect 123 446 124 447 
<< pdiffusion >>
rect 124 446 125 447 
<< pdiffusion >>
rect 125 446 126 447 
<< m1 >>
rect 150 446 151 447 
<< m1 >>
rect 152 446 153 447 
<< m1 >>
rect 154 446 155 447 
<< pdiffusion >>
rect 156 446 157 447 
<< pdiffusion >>
rect 157 446 158 447 
<< pdiffusion >>
rect 158 446 159 447 
<< pdiffusion >>
rect 159 446 160 447 
<< pdiffusion >>
rect 160 446 161 447 
<< pdiffusion >>
rect 161 446 162 447 
<< m1 >>
rect 163 446 164 447 
<< m1 >>
rect 170 446 171 447 
<< m1 >>
rect 172 446 173 447 
<< pdiffusion >>
rect 174 446 175 447 
<< pdiffusion >>
rect 175 446 176 447 
<< pdiffusion >>
rect 176 446 177 447 
<< pdiffusion >>
rect 177 446 178 447 
<< pdiffusion >>
rect 178 446 179 447 
<< pdiffusion >>
rect 179 446 180 447 
<< pdiffusion >>
rect 192 446 193 447 
<< pdiffusion >>
rect 193 446 194 447 
<< pdiffusion >>
rect 194 446 195 447 
<< pdiffusion >>
rect 195 446 196 447 
<< pdiffusion >>
rect 196 446 197 447 
<< pdiffusion >>
rect 197 446 198 447 
<< m1 >>
rect 204 446 205 447 
<< m1 >>
rect 208 446 209 447 
<< pdiffusion >>
rect 210 446 211 447 
<< pdiffusion >>
rect 211 446 212 447 
<< pdiffusion >>
rect 212 446 213 447 
<< pdiffusion >>
rect 213 446 214 447 
<< pdiffusion >>
rect 214 446 215 447 
<< pdiffusion >>
rect 215 446 216 447 
<< m1 >>
rect 217 446 218 447 
<< pdiffusion >>
rect 228 446 229 447 
<< pdiffusion >>
rect 229 446 230 447 
<< pdiffusion >>
rect 230 446 231 447 
<< pdiffusion >>
rect 231 446 232 447 
<< pdiffusion >>
rect 232 446 233 447 
<< pdiffusion >>
rect 233 446 234 447 
<< pdiffusion >>
rect 246 446 247 447 
<< pdiffusion >>
rect 247 446 248 447 
<< pdiffusion >>
rect 248 446 249 447 
<< pdiffusion >>
rect 249 446 250 447 
<< pdiffusion >>
rect 250 446 251 447 
<< pdiffusion >>
rect 251 446 252 447 
<< m1 >>
rect 253 446 254 447 
<< m2 >>
rect 254 446 255 447 
<< pdiffusion >>
rect 264 446 265 447 
<< pdiffusion >>
rect 265 446 266 447 
<< pdiffusion >>
rect 266 446 267 447 
<< pdiffusion >>
rect 267 446 268 447 
<< pdiffusion >>
rect 268 446 269 447 
<< pdiffusion >>
rect 269 446 270 447 
<< pdiffusion >>
rect 282 446 283 447 
<< pdiffusion >>
rect 283 446 284 447 
<< pdiffusion >>
rect 284 446 285 447 
<< pdiffusion >>
rect 285 446 286 447 
<< pdiffusion >>
rect 286 446 287 447 
<< pdiffusion >>
rect 287 446 288 447 
<< m1 >>
rect 289 446 290 447 
<< m1 >>
rect 298 446 299 447 
<< pdiffusion >>
rect 300 446 301 447 
<< pdiffusion >>
rect 301 446 302 447 
<< pdiffusion >>
rect 302 446 303 447 
<< pdiffusion >>
rect 303 446 304 447 
<< pdiffusion >>
rect 304 446 305 447 
<< pdiffusion >>
rect 305 446 306 447 
<< m1 >>
rect 307 446 308 447 
<< pdiffusion >>
rect 318 446 319 447 
<< pdiffusion >>
rect 319 446 320 447 
<< pdiffusion >>
rect 320 446 321 447 
<< pdiffusion >>
rect 321 446 322 447 
<< pdiffusion >>
rect 322 446 323 447 
<< pdiffusion >>
rect 323 446 324 447 
<< m1 >>
rect 325 446 326 447 
<< pdiffusion >>
rect 336 446 337 447 
<< pdiffusion >>
rect 337 446 338 447 
<< pdiffusion >>
rect 338 446 339 447 
<< pdiffusion >>
rect 339 446 340 447 
<< pdiffusion >>
rect 340 446 341 447 
<< pdiffusion >>
rect 341 446 342 447 
<< pdiffusion >>
rect 354 446 355 447 
<< pdiffusion >>
rect 355 446 356 447 
<< pdiffusion >>
rect 356 446 357 447 
<< pdiffusion >>
rect 357 446 358 447 
<< pdiffusion >>
rect 358 446 359 447 
<< pdiffusion >>
rect 359 446 360 447 
<< m1 >>
rect 361 446 362 447 
<< pdiffusion >>
rect 372 446 373 447 
<< pdiffusion >>
rect 373 446 374 447 
<< pdiffusion >>
rect 374 446 375 447 
<< pdiffusion >>
rect 375 446 376 447 
<< pdiffusion >>
rect 376 446 377 447 
<< pdiffusion >>
rect 377 446 378 447 
<< m1 >>
rect 379 446 380 447 
<< m1 >>
rect 381 446 382 447 
<< m1 >>
rect 385 446 386 447 
<< pdiffusion >>
rect 390 446 391 447 
<< pdiffusion >>
rect 391 446 392 447 
<< pdiffusion >>
rect 392 446 393 447 
<< pdiffusion >>
rect 393 446 394 447 
<< pdiffusion >>
rect 394 446 395 447 
<< pdiffusion >>
rect 395 446 396 447 
<< m1 >>
rect 397 446 398 447 
<< m1 >>
rect 400 446 401 447 
<< m1 >>
rect 402 446 403 447 
<< m1 >>
rect 406 446 407 447 
<< pdiffusion >>
rect 408 446 409 447 
<< pdiffusion >>
rect 409 446 410 447 
<< pdiffusion >>
rect 410 446 411 447 
<< pdiffusion >>
rect 411 446 412 447 
<< pdiffusion >>
rect 412 446 413 447 
<< pdiffusion >>
rect 413 446 414 447 
<< m1 >>
rect 424 446 425 447 
<< pdiffusion >>
rect 426 446 427 447 
<< pdiffusion >>
rect 427 446 428 447 
<< pdiffusion >>
rect 428 446 429 447 
<< pdiffusion >>
rect 429 446 430 447 
<< pdiffusion >>
rect 430 446 431 447 
<< pdiffusion >>
rect 431 446 432 447 
<< m1 >>
rect 433 446 434 447 
<< m2 >>
rect 434 446 435 447 
<< pdiffusion >>
rect 444 446 445 447 
<< pdiffusion >>
rect 445 446 446 447 
<< pdiffusion >>
rect 446 446 447 447 
<< pdiffusion >>
rect 447 446 448 447 
<< pdiffusion >>
rect 448 446 449 447 
<< pdiffusion >>
rect 449 446 450 447 
<< m1 >>
rect 452 446 453 447 
<< m2 >>
rect 453 446 454 447 
<< pdiffusion >>
rect 462 446 463 447 
<< pdiffusion >>
rect 463 446 464 447 
<< pdiffusion >>
rect 464 446 465 447 
<< pdiffusion >>
rect 465 446 466 447 
<< pdiffusion >>
rect 466 446 467 447 
<< pdiffusion >>
rect 467 446 468 447 
<< m1 >>
rect 470 446 471 447 
<< m1 >>
rect 472 446 473 447 
<< m1 >>
rect 478 446 479 447 
<< pdiffusion >>
rect 480 446 481 447 
<< pdiffusion >>
rect 481 446 482 447 
<< pdiffusion >>
rect 482 446 483 447 
<< pdiffusion >>
rect 483 446 484 447 
<< pdiffusion >>
rect 484 446 485 447 
<< pdiffusion >>
rect 485 446 486 447 
<< m1 >>
rect 487 446 488 447 
<< m1 >>
rect 489 446 490 447 
<< pdiffusion >>
rect 498 446 499 447 
<< pdiffusion >>
rect 499 446 500 447 
<< pdiffusion >>
rect 500 446 501 447 
<< pdiffusion >>
rect 501 446 502 447 
<< pdiffusion >>
rect 502 446 503 447 
<< pdiffusion >>
rect 503 446 504 447 
<< pdiffusion >>
rect 516 446 517 447 
<< pdiffusion >>
rect 517 446 518 447 
<< pdiffusion >>
rect 518 446 519 447 
<< pdiffusion >>
rect 519 446 520 447 
<< pdiffusion >>
rect 520 446 521 447 
<< pdiffusion >>
rect 521 446 522 447 
<< pdiffusion >>
rect 12 447 13 448 
<< pdiffusion >>
rect 13 447 14 448 
<< pdiffusion >>
rect 14 447 15 448 
<< pdiffusion >>
rect 15 447 16 448 
<< pdiffusion >>
rect 16 447 17 448 
<< pdiffusion >>
rect 17 447 18 448 
<< m1 >>
rect 19 447 20 448 
<< m1 >>
rect 21 447 22 448 
<< m1 >>
rect 26 447 27 448 
<< m1 >>
rect 28 447 29 448 
<< m2 >>
rect 28 447 29 448 
<< pdiffusion >>
rect 30 447 31 448 
<< pdiffusion >>
rect 31 447 32 448 
<< pdiffusion >>
rect 32 447 33 448 
<< pdiffusion >>
rect 33 447 34 448 
<< pdiffusion >>
rect 34 447 35 448 
<< pdiffusion >>
rect 35 447 36 448 
<< pdiffusion >>
rect 48 447 49 448 
<< pdiffusion >>
rect 49 447 50 448 
<< pdiffusion >>
rect 50 447 51 448 
<< pdiffusion >>
rect 51 447 52 448 
<< pdiffusion >>
rect 52 447 53 448 
<< pdiffusion >>
rect 53 447 54 448 
<< m1 >>
rect 55 447 56 448 
<< pdiffusion >>
rect 66 447 67 448 
<< pdiffusion >>
rect 67 447 68 448 
<< pdiffusion >>
rect 68 447 69 448 
<< pdiffusion >>
rect 69 447 70 448 
<< pdiffusion >>
rect 70 447 71 448 
<< pdiffusion >>
rect 71 447 72 448 
<< m1 >>
rect 73 447 74 448 
<< pdiffusion >>
rect 84 447 85 448 
<< pdiffusion >>
rect 85 447 86 448 
<< pdiffusion >>
rect 86 447 87 448 
<< pdiffusion >>
rect 87 447 88 448 
<< pdiffusion >>
rect 88 447 89 448 
<< pdiffusion >>
rect 89 447 90 448 
<< m2 >>
rect 99 447 100 448 
<< m1 >>
rect 100 447 101 448 
<< pdiffusion >>
rect 102 447 103 448 
<< pdiffusion >>
rect 103 447 104 448 
<< pdiffusion >>
rect 104 447 105 448 
<< pdiffusion >>
rect 105 447 106 448 
<< pdiffusion >>
rect 106 447 107 448 
<< pdiffusion >>
rect 107 447 108 448 
<< pdiffusion >>
rect 120 447 121 448 
<< pdiffusion >>
rect 121 447 122 448 
<< pdiffusion >>
rect 122 447 123 448 
<< pdiffusion >>
rect 123 447 124 448 
<< pdiffusion >>
rect 124 447 125 448 
<< pdiffusion >>
rect 125 447 126 448 
<< m1 >>
rect 150 447 151 448 
<< m1 >>
rect 152 447 153 448 
<< m1 >>
rect 154 447 155 448 
<< pdiffusion >>
rect 156 447 157 448 
<< pdiffusion >>
rect 157 447 158 448 
<< pdiffusion >>
rect 158 447 159 448 
<< pdiffusion >>
rect 159 447 160 448 
<< pdiffusion >>
rect 160 447 161 448 
<< pdiffusion >>
rect 161 447 162 448 
<< m1 >>
rect 163 447 164 448 
<< m1 >>
rect 170 447 171 448 
<< m1 >>
rect 172 447 173 448 
<< pdiffusion >>
rect 174 447 175 448 
<< pdiffusion >>
rect 175 447 176 448 
<< pdiffusion >>
rect 176 447 177 448 
<< pdiffusion >>
rect 177 447 178 448 
<< pdiffusion >>
rect 178 447 179 448 
<< pdiffusion >>
rect 179 447 180 448 
<< pdiffusion >>
rect 192 447 193 448 
<< pdiffusion >>
rect 193 447 194 448 
<< pdiffusion >>
rect 194 447 195 448 
<< pdiffusion >>
rect 195 447 196 448 
<< pdiffusion >>
rect 196 447 197 448 
<< pdiffusion >>
rect 197 447 198 448 
<< m1 >>
rect 204 447 205 448 
<< m1 >>
rect 208 447 209 448 
<< pdiffusion >>
rect 210 447 211 448 
<< pdiffusion >>
rect 211 447 212 448 
<< pdiffusion >>
rect 212 447 213 448 
<< pdiffusion >>
rect 213 447 214 448 
<< pdiffusion >>
rect 214 447 215 448 
<< pdiffusion >>
rect 215 447 216 448 
<< m1 >>
rect 217 447 218 448 
<< pdiffusion >>
rect 228 447 229 448 
<< pdiffusion >>
rect 229 447 230 448 
<< pdiffusion >>
rect 230 447 231 448 
<< pdiffusion >>
rect 231 447 232 448 
<< pdiffusion >>
rect 232 447 233 448 
<< pdiffusion >>
rect 233 447 234 448 
<< pdiffusion >>
rect 246 447 247 448 
<< pdiffusion >>
rect 247 447 248 448 
<< pdiffusion >>
rect 248 447 249 448 
<< pdiffusion >>
rect 249 447 250 448 
<< pdiffusion >>
rect 250 447 251 448 
<< pdiffusion >>
rect 251 447 252 448 
<< m1 >>
rect 253 447 254 448 
<< m2 >>
rect 254 447 255 448 
<< pdiffusion >>
rect 264 447 265 448 
<< pdiffusion >>
rect 265 447 266 448 
<< pdiffusion >>
rect 266 447 267 448 
<< pdiffusion >>
rect 267 447 268 448 
<< pdiffusion >>
rect 268 447 269 448 
<< pdiffusion >>
rect 269 447 270 448 
<< pdiffusion >>
rect 282 447 283 448 
<< pdiffusion >>
rect 283 447 284 448 
<< pdiffusion >>
rect 284 447 285 448 
<< pdiffusion >>
rect 285 447 286 448 
<< pdiffusion >>
rect 286 447 287 448 
<< pdiffusion >>
rect 287 447 288 448 
<< m1 >>
rect 289 447 290 448 
<< m1 >>
rect 298 447 299 448 
<< pdiffusion >>
rect 300 447 301 448 
<< pdiffusion >>
rect 301 447 302 448 
<< pdiffusion >>
rect 302 447 303 448 
<< pdiffusion >>
rect 303 447 304 448 
<< pdiffusion >>
rect 304 447 305 448 
<< pdiffusion >>
rect 305 447 306 448 
<< m1 >>
rect 307 447 308 448 
<< pdiffusion >>
rect 318 447 319 448 
<< pdiffusion >>
rect 319 447 320 448 
<< pdiffusion >>
rect 320 447 321 448 
<< pdiffusion >>
rect 321 447 322 448 
<< pdiffusion >>
rect 322 447 323 448 
<< pdiffusion >>
rect 323 447 324 448 
<< m1 >>
rect 325 447 326 448 
<< pdiffusion >>
rect 336 447 337 448 
<< pdiffusion >>
rect 337 447 338 448 
<< pdiffusion >>
rect 338 447 339 448 
<< pdiffusion >>
rect 339 447 340 448 
<< pdiffusion >>
rect 340 447 341 448 
<< pdiffusion >>
rect 341 447 342 448 
<< pdiffusion >>
rect 354 447 355 448 
<< pdiffusion >>
rect 355 447 356 448 
<< pdiffusion >>
rect 356 447 357 448 
<< pdiffusion >>
rect 357 447 358 448 
<< pdiffusion >>
rect 358 447 359 448 
<< pdiffusion >>
rect 359 447 360 448 
<< m1 >>
rect 361 447 362 448 
<< pdiffusion >>
rect 372 447 373 448 
<< pdiffusion >>
rect 373 447 374 448 
<< pdiffusion >>
rect 374 447 375 448 
<< pdiffusion >>
rect 375 447 376 448 
<< pdiffusion >>
rect 376 447 377 448 
<< pdiffusion >>
rect 377 447 378 448 
<< m1 >>
rect 379 447 380 448 
<< m1 >>
rect 381 447 382 448 
<< m1 >>
rect 385 447 386 448 
<< pdiffusion >>
rect 390 447 391 448 
<< pdiffusion >>
rect 391 447 392 448 
<< pdiffusion >>
rect 392 447 393 448 
<< pdiffusion >>
rect 393 447 394 448 
<< pdiffusion >>
rect 394 447 395 448 
<< pdiffusion >>
rect 395 447 396 448 
<< m1 >>
rect 397 447 398 448 
<< m1 >>
rect 400 447 401 448 
<< m2 >>
rect 400 447 401 448 
<< m2c >>
rect 400 447 401 448 
<< m1 >>
rect 400 447 401 448 
<< m2 >>
rect 400 447 401 448 
<< m2 >>
rect 401 447 402 448 
<< m1 >>
rect 402 447 403 448 
<< m2 >>
rect 402 447 403 448 
<< m2 >>
rect 403 447 404 448 
<< m1 >>
rect 404 447 405 448 
<< m2 >>
rect 404 447 405 448 
<< m2c >>
rect 404 447 405 448 
<< m1 >>
rect 404 447 405 448 
<< m2 >>
rect 404 447 405 448 
<< m1 >>
rect 406 447 407 448 
<< pdiffusion >>
rect 408 447 409 448 
<< pdiffusion >>
rect 409 447 410 448 
<< pdiffusion >>
rect 410 447 411 448 
<< pdiffusion >>
rect 411 447 412 448 
<< pdiffusion >>
rect 412 447 413 448 
<< pdiffusion >>
rect 413 447 414 448 
<< m1 >>
rect 424 447 425 448 
<< pdiffusion >>
rect 426 447 427 448 
<< pdiffusion >>
rect 427 447 428 448 
<< pdiffusion >>
rect 428 447 429 448 
<< pdiffusion >>
rect 429 447 430 448 
<< pdiffusion >>
rect 430 447 431 448 
<< pdiffusion >>
rect 431 447 432 448 
<< m1 >>
rect 433 447 434 448 
<< m2 >>
rect 434 447 435 448 
<< pdiffusion >>
rect 444 447 445 448 
<< pdiffusion >>
rect 445 447 446 448 
<< pdiffusion >>
rect 446 447 447 448 
<< pdiffusion >>
rect 447 447 448 448 
<< pdiffusion >>
rect 448 447 449 448 
<< pdiffusion >>
rect 449 447 450 448 
<< m1 >>
rect 452 447 453 448 
<< m2 >>
rect 453 447 454 448 
<< pdiffusion >>
rect 462 447 463 448 
<< pdiffusion >>
rect 463 447 464 448 
<< pdiffusion >>
rect 464 447 465 448 
<< pdiffusion >>
rect 465 447 466 448 
<< pdiffusion >>
rect 466 447 467 448 
<< pdiffusion >>
rect 467 447 468 448 
<< m1 >>
rect 470 447 471 448 
<< m1 >>
rect 472 447 473 448 
<< m1 >>
rect 478 447 479 448 
<< pdiffusion >>
rect 480 447 481 448 
<< pdiffusion >>
rect 481 447 482 448 
<< pdiffusion >>
rect 482 447 483 448 
<< pdiffusion >>
rect 483 447 484 448 
<< pdiffusion >>
rect 484 447 485 448 
<< pdiffusion >>
rect 485 447 486 448 
<< m1 >>
rect 487 447 488 448 
<< m1 >>
rect 489 447 490 448 
<< pdiffusion >>
rect 498 447 499 448 
<< pdiffusion >>
rect 499 447 500 448 
<< pdiffusion >>
rect 500 447 501 448 
<< pdiffusion >>
rect 501 447 502 448 
<< pdiffusion >>
rect 502 447 503 448 
<< pdiffusion >>
rect 503 447 504 448 
<< pdiffusion >>
rect 516 447 517 448 
<< pdiffusion >>
rect 517 447 518 448 
<< pdiffusion >>
rect 518 447 519 448 
<< pdiffusion >>
rect 519 447 520 448 
<< pdiffusion >>
rect 520 447 521 448 
<< pdiffusion >>
rect 521 447 522 448 
<< pdiffusion >>
rect 12 448 13 449 
<< pdiffusion >>
rect 13 448 14 449 
<< pdiffusion >>
rect 14 448 15 449 
<< pdiffusion >>
rect 15 448 16 449 
<< pdiffusion >>
rect 16 448 17 449 
<< pdiffusion >>
rect 17 448 18 449 
<< m1 >>
rect 19 448 20 449 
<< m1 >>
rect 21 448 22 449 
<< m1 >>
rect 26 448 27 449 
<< m1 >>
rect 28 448 29 449 
<< m2 >>
rect 28 448 29 449 
<< pdiffusion >>
rect 30 448 31 449 
<< pdiffusion >>
rect 31 448 32 449 
<< pdiffusion >>
rect 32 448 33 449 
<< pdiffusion >>
rect 33 448 34 449 
<< pdiffusion >>
rect 34 448 35 449 
<< pdiffusion >>
rect 35 448 36 449 
<< pdiffusion >>
rect 48 448 49 449 
<< pdiffusion >>
rect 49 448 50 449 
<< pdiffusion >>
rect 50 448 51 449 
<< pdiffusion >>
rect 51 448 52 449 
<< pdiffusion >>
rect 52 448 53 449 
<< pdiffusion >>
rect 53 448 54 449 
<< m1 >>
rect 55 448 56 449 
<< pdiffusion >>
rect 66 448 67 449 
<< pdiffusion >>
rect 67 448 68 449 
<< pdiffusion >>
rect 68 448 69 449 
<< pdiffusion >>
rect 69 448 70 449 
<< pdiffusion >>
rect 70 448 71 449 
<< pdiffusion >>
rect 71 448 72 449 
<< m1 >>
rect 73 448 74 449 
<< pdiffusion >>
rect 84 448 85 449 
<< pdiffusion >>
rect 85 448 86 449 
<< pdiffusion >>
rect 86 448 87 449 
<< pdiffusion >>
rect 87 448 88 449 
<< pdiffusion >>
rect 88 448 89 449 
<< pdiffusion >>
rect 89 448 90 449 
<< m2 >>
rect 99 448 100 449 
<< m1 >>
rect 100 448 101 449 
<< pdiffusion >>
rect 102 448 103 449 
<< pdiffusion >>
rect 103 448 104 449 
<< pdiffusion >>
rect 104 448 105 449 
<< pdiffusion >>
rect 105 448 106 449 
<< pdiffusion >>
rect 106 448 107 449 
<< pdiffusion >>
rect 107 448 108 449 
<< pdiffusion >>
rect 120 448 121 449 
<< pdiffusion >>
rect 121 448 122 449 
<< pdiffusion >>
rect 122 448 123 449 
<< pdiffusion >>
rect 123 448 124 449 
<< pdiffusion >>
rect 124 448 125 449 
<< pdiffusion >>
rect 125 448 126 449 
<< m1 >>
rect 150 448 151 449 
<< m1 >>
rect 152 448 153 449 
<< m1 >>
rect 154 448 155 449 
<< pdiffusion >>
rect 156 448 157 449 
<< pdiffusion >>
rect 157 448 158 449 
<< pdiffusion >>
rect 158 448 159 449 
<< pdiffusion >>
rect 159 448 160 449 
<< pdiffusion >>
rect 160 448 161 449 
<< pdiffusion >>
rect 161 448 162 449 
<< m1 >>
rect 163 448 164 449 
<< m1 >>
rect 170 448 171 449 
<< m1 >>
rect 172 448 173 449 
<< pdiffusion >>
rect 174 448 175 449 
<< pdiffusion >>
rect 175 448 176 449 
<< pdiffusion >>
rect 176 448 177 449 
<< pdiffusion >>
rect 177 448 178 449 
<< pdiffusion >>
rect 178 448 179 449 
<< pdiffusion >>
rect 179 448 180 449 
<< pdiffusion >>
rect 192 448 193 449 
<< pdiffusion >>
rect 193 448 194 449 
<< pdiffusion >>
rect 194 448 195 449 
<< pdiffusion >>
rect 195 448 196 449 
<< pdiffusion >>
rect 196 448 197 449 
<< pdiffusion >>
rect 197 448 198 449 
<< m1 >>
rect 204 448 205 449 
<< m1 >>
rect 208 448 209 449 
<< pdiffusion >>
rect 210 448 211 449 
<< pdiffusion >>
rect 211 448 212 449 
<< pdiffusion >>
rect 212 448 213 449 
<< pdiffusion >>
rect 213 448 214 449 
<< pdiffusion >>
rect 214 448 215 449 
<< pdiffusion >>
rect 215 448 216 449 
<< m1 >>
rect 217 448 218 449 
<< pdiffusion >>
rect 228 448 229 449 
<< pdiffusion >>
rect 229 448 230 449 
<< pdiffusion >>
rect 230 448 231 449 
<< pdiffusion >>
rect 231 448 232 449 
<< pdiffusion >>
rect 232 448 233 449 
<< pdiffusion >>
rect 233 448 234 449 
<< pdiffusion >>
rect 246 448 247 449 
<< pdiffusion >>
rect 247 448 248 449 
<< pdiffusion >>
rect 248 448 249 449 
<< pdiffusion >>
rect 249 448 250 449 
<< pdiffusion >>
rect 250 448 251 449 
<< pdiffusion >>
rect 251 448 252 449 
<< m1 >>
rect 253 448 254 449 
<< m2 >>
rect 254 448 255 449 
<< pdiffusion >>
rect 264 448 265 449 
<< pdiffusion >>
rect 265 448 266 449 
<< pdiffusion >>
rect 266 448 267 449 
<< pdiffusion >>
rect 267 448 268 449 
<< pdiffusion >>
rect 268 448 269 449 
<< pdiffusion >>
rect 269 448 270 449 
<< pdiffusion >>
rect 282 448 283 449 
<< pdiffusion >>
rect 283 448 284 449 
<< pdiffusion >>
rect 284 448 285 449 
<< pdiffusion >>
rect 285 448 286 449 
<< pdiffusion >>
rect 286 448 287 449 
<< pdiffusion >>
rect 287 448 288 449 
<< m1 >>
rect 289 448 290 449 
<< m1 >>
rect 298 448 299 449 
<< pdiffusion >>
rect 300 448 301 449 
<< pdiffusion >>
rect 301 448 302 449 
<< pdiffusion >>
rect 302 448 303 449 
<< pdiffusion >>
rect 303 448 304 449 
<< pdiffusion >>
rect 304 448 305 449 
<< pdiffusion >>
rect 305 448 306 449 
<< m1 >>
rect 307 448 308 449 
<< pdiffusion >>
rect 318 448 319 449 
<< pdiffusion >>
rect 319 448 320 449 
<< pdiffusion >>
rect 320 448 321 449 
<< pdiffusion >>
rect 321 448 322 449 
<< pdiffusion >>
rect 322 448 323 449 
<< pdiffusion >>
rect 323 448 324 449 
<< m1 >>
rect 325 448 326 449 
<< pdiffusion >>
rect 336 448 337 449 
<< pdiffusion >>
rect 337 448 338 449 
<< pdiffusion >>
rect 338 448 339 449 
<< pdiffusion >>
rect 339 448 340 449 
<< pdiffusion >>
rect 340 448 341 449 
<< pdiffusion >>
rect 341 448 342 449 
<< pdiffusion >>
rect 354 448 355 449 
<< pdiffusion >>
rect 355 448 356 449 
<< pdiffusion >>
rect 356 448 357 449 
<< pdiffusion >>
rect 357 448 358 449 
<< pdiffusion >>
rect 358 448 359 449 
<< pdiffusion >>
rect 359 448 360 449 
<< m1 >>
rect 361 448 362 449 
<< pdiffusion >>
rect 372 448 373 449 
<< pdiffusion >>
rect 373 448 374 449 
<< pdiffusion >>
rect 374 448 375 449 
<< pdiffusion >>
rect 375 448 376 449 
<< pdiffusion >>
rect 376 448 377 449 
<< pdiffusion >>
rect 377 448 378 449 
<< m1 >>
rect 379 448 380 449 
<< m1 >>
rect 381 448 382 449 
<< m1 >>
rect 385 448 386 449 
<< pdiffusion >>
rect 390 448 391 449 
<< pdiffusion >>
rect 391 448 392 449 
<< pdiffusion >>
rect 392 448 393 449 
<< pdiffusion >>
rect 393 448 394 449 
<< pdiffusion >>
rect 394 448 395 449 
<< pdiffusion >>
rect 395 448 396 449 
<< m1 >>
rect 397 448 398 449 
<< m1 >>
rect 402 448 403 449 
<< m1 >>
rect 404 448 405 449 
<< m1 >>
rect 406 448 407 449 
<< pdiffusion >>
rect 408 448 409 449 
<< pdiffusion >>
rect 409 448 410 449 
<< pdiffusion >>
rect 410 448 411 449 
<< pdiffusion >>
rect 411 448 412 449 
<< pdiffusion >>
rect 412 448 413 449 
<< pdiffusion >>
rect 413 448 414 449 
<< m1 >>
rect 424 448 425 449 
<< pdiffusion >>
rect 426 448 427 449 
<< pdiffusion >>
rect 427 448 428 449 
<< pdiffusion >>
rect 428 448 429 449 
<< pdiffusion >>
rect 429 448 430 449 
<< pdiffusion >>
rect 430 448 431 449 
<< pdiffusion >>
rect 431 448 432 449 
<< m1 >>
rect 433 448 434 449 
<< m2 >>
rect 434 448 435 449 
<< pdiffusion >>
rect 444 448 445 449 
<< pdiffusion >>
rect 445 448 446 449 
<< pdiffusion >>
rect 446 448 447 449 
<< pdiffusion >>
rect 447 448 448 449 
<< pdiffusion >>
rect 448 448 449 449 
<< pdiffusion >>
rect 449 448 450 449 
<< m1 >>
rect 452 448 453 449 
<< m2 >>
rect 453 448 454 449 
<< pdiffusion >>
rect 462 448 463 449 
<< pdiffusion >>
rect 463 448 464 449 
<< pdiffusion >>
rect 464 448 465 449 
<< pdiffusion >>
rect 465 448 466 449 
<< pdiffusion >>
rect 466 448 467 449 
<< pdiffusion >>
rect 467 448 468 449 
<< m1 >>
rect 470 448 471 449 
<< m1 >>
rect 472 448 473 449 
<< m1 >>
rect 478 448 479 449 
<< pdiffusion >>
rect 480 448 481 449 
<< pdiffusion >>
rect 481 448 482 449 
<< pdiffusion >>
rect 482 448 483 449 
<< pdiffusion >>
rect 483 448 484 449 
<< pdiffusion >>
rect 484 448 485 449 
<< pdiffusion >>
rect 485 448 486 449 
<< m1 >>
rect 487 448 488 449 
<< m1 >>
rect 489 448 490 449 
<< pdiffusion >>
rect 498 448 499 449 
<< pdiffusion >>
rect 499 448 500 449 
<< pdiffusion >>
rect 500 448 501 449 
<< pdiffusion >>
rect 501 448 502 449 
<< pdiffusion >>
rect 502 448 503 449 
<< pdiffusion >>
rect 503 448 504 449 
<< pdiffusion >>
rect 516 448 517 449 
<< pdiffusion >>
rect 517 448 518 449 
<< pdiffusion >>
rect 518 448 519 449 
<< pdiffusion >>
rect 519 448 520 449 
<< pdiffusion >>
rect 520 448 521 449 
<< pdiffusion >>
rect 521 448 522 449 
<< pdiffusion >>
rect 12 449 13 450 
<< pdiffusion >>
rect 13 449 14 450 
<< pdiffusion >>
rect 14 449 15 450 
<< pdiffusion >>
rect 15 449 16 450 
<< pdiffusion >>
rect 16 449 17 450 
<< pdiffusion >>
rect 17 449 18 450 
<< m1 >>
rect 19 449 20 450 
<< m1 >>
rect 21 449 22 450 
<< m1 >>
rect 26 449 27 450 
<< m1 >>
rect 28 449 29 450 
<< m2 >>
rect 28 449 29 450 
<< pdiffusion >>
rect 30 449 31 450 
<< pdiffusion >>
rect 31 449 32 450 
<< pdiffusion >>
rect 32 449 33 450 
<< pdiffusion >>
rect 33 449 34 450 
<< pdiffusion >>
rect 34 449 35 450 
<< pdiffusion >>
rect 35 449 36 450 
<< pdiffusion >>
rect 48 449 49 450 
<< pdiffusion >>
rect 49 449 50 450 
<< pdiffusion >>
rect 50 449 51 450 
<< pdiffusion >>
rect 51 449 52 450 
<< pdiffusion >>
rect 52 449 53 450 
<< pdiffusion >>
rect 53 449 54 450 
<< m1 >>
rect 55 449 56 450 
<< pdiffusion >>
rect 66 449 67 450 
<< pdiffusion >>
rect 67 449 68 450 
<< pdiffusion >>
rect 68 449 69 450 
<< pdiffusion >>
rect 69 449 70 450 
<< pdiffusion >>
rect 70 449 71 450 
<< pdiffusion >>
rect 71 449 72 450 
<< m1 >>
rect 73 449 74 450 
<< pdiffusion >>
rect 84 449 85 450 
<< pdiffusion >>
rect 85 449 86 450 
<< pdiffusion >>
rect 86 449 87 450 
<< pdiffusion >>
rect 87 449 88 450 
<< pdiffusion >>
rect 88 449 89 450 
<< pdiffusion >>
rect 89 449 90 450 
<< m2 >>
rect 99 449 100 450 
<< m1 >>
rect 100 449 101 450 
<< pdiffusion >>
rect 102 449 103 450 
<< pdiffusion >>
rect 103 449 104 450 
<< pdiffusion >>
rect 104 449 105 450 
<< pdiffusion >>
rect 105 449 106 450 
<< pdiffusion >>
rect 106 449 107 450 
<< pdiffusion >>
rect 107 449 108 450 
<< pdiffusion >>
rect 120 449 121 450 
<< pdiffusion >>
rect 121 449 122 450 
<< pdiffusion >>
rect 122 449 123 450 
<< pdiffusion >>
rect 123 449 124 450 
<< pdiffusion >>
rect 124 449 125 450 
<< pdiffusion >>
rect 125 449 126 450 
<< m1 >>
rect 150 449 151 450 
<< m1 >>
rect 152 449 153 450 
<< m1 >>
rect 154 449 155 450 
<< pdiffusion >>
rect 156 449 157 450 
<< pdiffusion >>
rect 157 449 158 450 
<< pdiffusion >>
rect 158 449 159 450 
<< pdiffusion >>
rect 159 449 160 450 
<< pdiffusion >>
rect 160 449 161 450 
<< pdiffusion >>
rect 161 449 162 450 
<< m1 >>
rect 163 449 164 450 
<< m1 >>
rect 170 449 171 450 
<< m1 >>
rect 172 449 173 450 
<< pdiffusion >>
rect 174 449 175 450 
<< pdiffusion >>
rect 175 449 176 450 
<< pdiffusion >>
rect 176 449 177 450 
<< pdiffusion >>
rect 177 449 178 450 
<< pdiffusion >>
rect 178 449 179 450 
<< pdiffusion >>
rect 179 449 180 450 
<< pdiffusion >>
rect 192 449 193 450 
<< pdiffusion >>
rect 193 449 194 450 
<< pdiffusion >>
rect 194 449 195 450 
<< pdiffusion >>
rect 195 449 196 450 
<< m1 >>
rect 196 449 197 450 
<< pdiffusion >>
rect 196 449 197 450 
<< pdiffusion >>
rect 197 449 198 450 
<< m1 >>
rect 204 449 205 450 
<< m1 >>
rect 205 449 206 450 
<< m1 >>
rect 206 449 207 450 
<< m2 >>
rect 206 449 207 450 
<< m2c >>
rect 206 449 207 450 
<< m1 >>
rect 206 449 207 450 
<< m2 >>
rect 206 449 207 450 
<< m2 >>
rect 207 449 208 450 
<< m1 >>
rect 208 449 209 450 
<< m2 >>
rect 208 449 209 450 
<< pdiffusion >>
rect 210 449 211 450 
<< pdiffusion >>
rect 211 449 212 450 
<< pdiffusion >>
rect 212 449 213 450 
<< pdiffusion >>
rect 213 449 214 450 
<< pdiffusion >>
rect 214 449 215 450 
<< pdiffusion >>
rect 215 449 216 450 
<< m1 >>
rect 217 449 218 450 
<< pdiffusion >>
rect 228 449 229 450 
<< m1 >>
rect 229 449 230 450 
<< pdiffusion >>
rect 229 449 230 450 
<< pdiffusion >>
rect 230 449 231 450 
<< pdiffusion >>
rect 231 449 232 450 
<< pdiffusion >>
rect 232 449 233 450 
<< pdiffusion >>
rect 233 449 234 450 
<< pdiffusion >>
rect 246 449 247 450 
<< pdiffusion >>
rect 247 449 248 450 
<< pdiffusion >>
rect 248 449 249 450 
<< pdiffusion >>
rect 249 449 250 450 
<< pdiffusion >>
rect 250 449 251 450 
<< pdiffusion >>
rect 251 449 252 450 
<< m1 >>
rect 253 449 254 450 
<< m2 >>
rect 254 449 255 450 
<< pdiffusion >>
rect 264 449 265 450 
<< pdiffusion >>
rect 265 449 266 450 
<< pdiffusion >>
rect 266 449 267 450 
<< pdiffusion >>
rect 267 449 268 450 
<< pdiffusion >>
rect 268 449 269 450 
<< pdiffusion >>
rect 269 449 270 450 
<< pdiffusion >>
rect 282 449 283 450 
<< m1 >>
rect 283 449 284 450 
<< pdiffusion >>
rect 283 449 284 450 
<< pdiffusion >>
rect 284 449 285 450 
<< pdiffusion >>
rect 285 449 286 450 
<< pdiffusion >>
rect 286 449 287 450 
<< pdiffusion >>
rect 287 449 288 450 
<< m1 >>
rect 289 449 290 450 
<< m1 >>
rect 298 449 299 450 
<< pdiffusion >>
rect 300 449 301 450 
<< pdiffusion >>
rect 301 449 302 450 
<< pdiffusion >>
rect 302 449 303 450 
<< pdiffusion >>
rect 303 449 304 450 
<< pdiffusion >>
rect 304 449 305 450 
<< pdiffusion >>
rect 305 449 306 450 
<< m1 >>
rect 307 449 308 450 
<< pdiffusion >>
rect 318 449 319 450 
<< m1 >>
rect 319 449 320 450 
<< pdiffusion >>
rect 319 449 320 450 
<< pdiffusion >>
rect 320 449 321 450 
<< pdiffusion >>
rect 321 449 322 450 
<< pdiffusion >>
rect 322 449 323 450 
<< pdiffusion >>
rect 323 449 324 450 
<< m1 >>
rect 325 449 326 450 
<< pdiffusion >>
rect 336 449 337 450 
<< pdiffusion >>
rect 337 449 338 450 
<< pdiffusion >>
rect 338 449 339 450 
<< pdiffusion >>
rect 339 449 340 450 
<< pdiffusion >>
rect 340 449 341 450 
<< pdiffusion >>
rect 341 449 342 450 
<< pdiffusion >>
rect 354 449 355 450 
<< pdiffusion >>
rect 355 449 356 450 
<< pdiffusion >>
rect 356 449 357 450 
<< pdiffusion >>
rect 357 449 358 450 
<< pdiffusion >>
rect 358 449 359 450 
<< pdiffusion >>
rect 359 449 360 450 
<< m1 >>
rect 361 449 362 450 
<< pdiffusion >>
rect 372 449 373 450 
<< m1 >>
rect 373 449 374 450 
<< pdiffusion >>
rect 373 449 374 450 
<< pdiffusion >>
rect 374 449 375 450 
<< pdiffusion >>
rect 375 449 376 450 
<< pdiffusion >>
rect 376 449 377 450 
<< pdiffusion >>
rect 377 449 378 450 
<< m1 >>
rect 379 449 380 450 
<< m1 >>
rect 381 449 382 450 
<< m1 >>
rect 385 449 386 450 
<< pdiffusion >>
rect 390 449 391 450 
<< pdiffusion >>
rect 391 449 392 450 
<< pdiffusion >>
rect 392 449 393 450 
<< pdiffusion >>
rect 393 449 394 450 
<< m1 >>
rect 394 449 395 450 
<< pdiffusion >>
rect 394 449 395 450 
<< pdiffusion >>
rect 395 449 396 450 
<< m1 >>
rect 397 449 398 450 
<< m2 >>
rect 397 449 398 450 
<< m2c >>
rect 397 449 398 450 
<< m1 >>
rect 397 449 398 450 
<< m2 >>
rect 397 449 398 450 
<< m1 >>
rect 402 449 403 450 
<< m2 >>
rect 402 449 403 450 
<< m2c >>
rect 402 449 403 450 
<< m1 >>
rect 402 449 403 450 
<< m2 >>
rect 402 449 403 450 
<< m1 >>
rect 404 449 405 450 
<< m2 >>
rect 404 449 405 450 
<< m2c >>
rect 404 449 405 450 
<< m1 >>
rect 404 449 405 450 
<< m2 >>
rect 404 449 405 450 
<< m2 >>
rect 405 449 406 450 
<< m1 >>
rect 406 449 407 450 
<< m2 >>
rect 406 449 407 450 
<< pdiffusion >>
rect 408 449 409 450 
<< pdiffusion >>
rect 409 449 410 450 
<< pdiffusion >>
rect 410 449 411 450 
<< pdiffusion >>
rect 411 449 412 450 
<< pdiffusion >>
rect 412 449 413 450 
<< pdiffusion >>
rect 413 449 414 450 
<< m1 >>
rect 424 449 425 450 
<< pdiffusion >>
rect 426 449 427 450 
<< pdiffusion >>
rect 427 449 428 450 
<< pdiffusion >>
rect 428 449 429 450 
<< pdiffusion >>
rect 429 449 430 450 
<< pdiffusion >>
rect 430 449 431 450 
<< pdiffusion >>
rect 431 449 432 450 
<< m1 >>
rect 433 449 434 450 
<< m2 >>
rect 434 449 435 450 
<< pdiffusion >>
rect 444 449 445 450 
<< pdiffusion >>
rect 445 449 446 450 
<< pdiffusion >>
rect 446 449 447 450 
<< pdiffusion >>
rect 447 449 448 450 
<< pdiffusion >>
rect 448 449 449 450 
<< pdiffusion >>
rect 449 449 450 450 
<< m1 >>
rect 452 449 453 450 
<< m2 >>
rect 453 449 454 450 
<< pdiffusion >>
rect 462 449 463 450 
<< pdiffusion >>
rect 463 449 464 450 
<< pdiffusion >>
rect 464 449 465 450 
<< pdiffusion >>
rect 465 449 466 450 
<< pdiffusion >>
rect 466 449 467 450 
<< pdiffusion >>
rect 467 449 468 450 
<< m1 >>
rect 470 449 471 450 
<< m1 >>
rect 472 449 473 450 
<< m1 >>
rect 478 449 479 450 
<< m2 >>
rect 478 449 479 450 
<< m2c >>
rect 478 449 479 450 
<< m1 >>
rect 478 449 479 450 
<< m2 >>
rect 478 449 479 450 
<< pdiffusion >>
rect 480 449 481 450 
<< m1 >>
rect 481 449 482 450 
<< pdiffusion >>
rect 481 449 482 450 
<< pdiffusion >>
rect 482 449 483 450 
<< pdiffusion >>
rect 483 449 484 450 
<< pdiffusion >>
rect 484 449 485 450 
<< pdiffusion >>
rect 485 449 486 450 
<< m1 >>
rect 487 449 488 450 
<< m1 >>
rect 489 449 490 450 
<< pdiffusion >>
rect 498 449 499 450 
<< pdiffusion >>
rect 499 449 500 450 
<< pdiffusion >>
rect 500 449 501 450 
<< pdiffusion >>
rect 501 449 502 450 
<< pdiffusion >>
rect 502 449 503 450 
<< pdiffusion >>
rect 503 449 504 450 
<< pdiffusion >>
rect 516 449 517 450 
<< pdiffusion >>
rect 517 449 518 450 
<< pdiffusion >>
rect 518 449 519 450 
<< pdiffusion >>
rect 519 449 520 450 
<< pdiffusion >>
rect 520 449 521 450 
<< pdiffusion >>
rect 521 449 522 450 
<< m1 >>
rect 19 450 20 451 
<< m1 >>
rect 21 450 22 451 
<< m1 >>
rect 26 450 27 451 
<< m1 >>
rect 28 450 29 451 
<< m2 >>
rect 28 450 29 451 
<< m1 >>
rect 55 450 56 451 
<< m1 >>
rect 73 450 74 451 
<< m2 >>
rect 99 450 100 451 
<< m1 >>
rect 100 450 101 451 
<< m1 >>
rect 150 450 151 451 
<< m1 >>
rect 152 450 153 451 
<< m1 >>
rect 154 450 155 451 
<< m1 >>
rect 163 450 164 451 
<< m2 >>
rect 163 450 164 451 
<< m2c >>
rect 163 450 164 451 
<< m1 >>
rect 163 450 164 451 
<< m2 >>
rect 163 450 164 451 
<< m1 >>
rect 170 450 171 451 
<< m2 >>
rect 170 450 171 451 
<< m2c >>
rect 170 450 171 451 
<< m1 >>
rect 170 450 171 451 
<< m2 >>
rect 170 450 171 451 
<< m2 >>
rect 171 450 172 451 
<< m1 >>
rect 172 450 173 451 
<< m2 >>
rect 172 450 173 451 
<< m1 >>
rect 196 450 197 451 
<< m1 >>
rect 208 450 209 451 
<< m2 >>
rect 208 450 209 451 
<< m1 >>
rect 217 450 218 451 
<< m1 >>
rect 229 450 230 451 
<< m1 >>
rect 253 450 254 451 
<< m2 >>
rect 254 450 255 451 
<< m1 >>
rect 283 450 284 451 
<< m1 >>
rect 289 450 290 451 
<< m1 >>
rect 298 450 299 451 
<< m1 >>
rect 307 450 308 451 
<< m1 >>
rect 319 450 320 451 
<< m1 >>
rect 325 450 326 451 
<< m1 >>
rect 361 450 362 451 
<< m1 >>
rect 373 450 374 451 
<< m1 >>
rect 379 450 380 451 
<< m1 >>
rect 381 450 382 451 
<< m1 >>
rect 385 450 386 451 
<< m1 >>
rect 394 450 395 451 
<< m2 >>
rect 397 450 398 451 
<< m2 >>
rect 402 450 403 451 
<< m1 >>
rect 406 450 407 451 
<< m2 >>
rect 406 450 407 451 
<< m1 >>
rect 424 450 425 451 
<< m1 >>
rect 433 450 434 451 
<< m2 >>
rect 434 450 435 451 
<< m1 >>
rect 452 450 453 451 
<< m2 >>
rect 453 450 454 451 
<< m1 >>
rect 470 450 471 451 
<< m1 >>
rect 472 450 473 451 
<< m2 >>
rect 478 450 479 451 
<< m1 >>
rect 481 450 482 451 
<< m1 >>
rect 487 450 488 451 
<< m1 >>
rect 489 450 490 451 
<< m1 >>
rect 19 451 20 452 
<< m1 >>
rect 21 451 22 452 
<< m1 >>
rect 26 451 27 452 
<< m1 >>
rect 28 451 29 452 
<< m2 >>
rect 28 451 29 452 
<< m2 >>
rect 29 451 30 452 
<< m1 >>
rect 30 451 31 452 
<< m2 >>
rect 30 451 31 452 
<< m2c >>
rect 30 451 31 452 
<< m1 >>
rect 30 451 31 452 
<< m2 >>
rect 30 451 31 452 
<< m1 >>
rect 55 451 56 452 
<< m1 >>
rect 73 451 74 452 
<< m2 >>
rect 99 451 100 452 
<< m1 >>
rect 100 451 101 452 
<< m1 >>
rect 150 451 151 452 
<< m1 >>
rect 152 451 153 452 
<< m1 >>
rect 154 451 155 452 
<< m2 >>
rect 163 451 164 452 
<< m1 >>
rect 172 451 173 452 
<< m2 >>
rect 172 451 173 452 
<< m1 >>
rect 196 451 197 452 
<< m2 >>
rect 197 451 198 452 
<< m1 >>
rect 198 451 199 452 
<< m2 >>
rect 198 451 199 452 
<< m2c >>
rect 198 451 199 452 
<< m1 >>
rect 198 451 199 452 
<< m2 >>
rect 198 451 199 452 
<< m1 >>
rect 199 451 200 452 
<< m1 >>
rect 200 451 201 452 
<< m1 >>
rect 201 451 202 452 
<< m1 >>
rect 202 451 203 452 
<< m1 >>
rect 203 451 204 452 
<< m1 >>
rect 204 451 205 452 
<< m1 >>
rect 205 451 206 452 
<< m1 >>
rect 206 451 207 452 
<< m1 >>
rect 207 451 208 452 
<< m1 >>
rect 208 451 209 452 
<< m2 >>
rect 208 451 209 452 
<< m1 >>
rect 217 451 218 452 
<< m1 >>
rect 229 451 230 452 
<< m1 >>
rect 253 451 254 452 
<< m2 >>
rect 254 451 255 452 
<< m1 >>
rect 283 451 284 452 
<< m1 >>
rect 289 451 290 452 
<< m1 >>
rect 298 451 299 452 
<< m1 >>
rect 307 451 308 452 
<< m1 >>
rect 319 451 320 452 
<< m1 >>
rect 325 451 326 452 
<< m1 >>
rect 361 451 362 452 
<< m1 >>
rect 373 451 374 452 
<< m1 >>
rect 379 451 380 452 
<< m1 >>
rect 381 451 382 452 
<< m1 >>
rect 385 451 386 452 
<< m1 >>
rect 394 451 395 452 
<< m1 >>
rect 395 451 396 452 
<< m1 >>
rect 396 451 397 452 
<< m1 >>
rect 397 451 398 452 
<< m2 >>
rect 397 451 398 452 
<< m1 >>
rect 398 451 399 452 
<< m1 >>
rect 399 451 400 452 
<< m1 >>
rect 400 451 401 452 
<< m1 >>
rect 401 451 402 452 
<< m1 >>
rect 402 451 403 452 
<< m2 >>
rect 402 451 403 452 
<< m1 >>
rect 403 451 404 452 
<< m1 >>
rect 404 451 405 452 
<< m1 >>
rect 405 451 406 452 
<< m1 >>
rect 406 451 407 452 
<< m2 >>
rect 406 451 407 452 
<< m1 >>
rect 424 451 425 452 
<< m1 >>
rect 431 451 432 452 
<< m2 >>
rect 431 451 432 452 
<< m2c >>
rect 431 451 432 452 
<< m1 >>
rect 431 451 432 452 
<< m2 >>
rect 431 451 432 452 
<< m2 >>
rect 432 451 433 452 
<< m1 >>
rect 433 451 434 452 
<< m2 >>
rect 433 451 434 452 
<< m2 >>
rect 434 451 435 452 
<< m1 >>
rect 450 451 451 452 
<< m2 >>
rect 450 451 451 452 
<< m2c >>
rect 450 451 451 452 
<< m1 >>
rect 450 451 451 452 
<< m2 >>
rect 450 451 451 452 
<< m2 >>
rect 451 451 452 452 
<< m1 >>
rect 452 451 453 452 
<< m2 >>
rect 452 451 453 452 
<< m2 >>
rect 453 451 454 452 
<< m1 >>
rect 470 451 471 452 
<< m2 >>
rect 470 451 471 452 
<< m2c >>
rect 470 451 471 452 
<< m1 >>
rect 470 451 471 452 
<< m2 >>
rect 470 451 471 452 
<< m2 >>
rect 471 451 472 452 
<< m1 >>
rect 472 451 473 452 
<< m2 >>
rect 472 451 473 452 
<< m2 >>
rect 473 451 474 452 
<< m1 >>
rect 474 451 475 452 
<< m2 >>
rect 474 451 475 452 
<< m2c >>
rect 474 451 475 452 
<< m1 >>
rect 474 451 475 452 
<< m2 >>
rect 474 451 475 452 
<< m1 >>
rect 475 451 476 452 
<< m1 >>
rect 476 451 477 452 
<< m1 >>
rect 477 451 478 452 
<< m1 >>
rect 478 451 479 452 
<< m2 >>
rect 478 451 479 452 
<< m1 >>
rect 479 451 480 452 
<< m1 >>
rect 480 451 481 452 
<< m1 >>
rect 481 451 482 452 
<< m1 >>
rect 487 451 488 452 
<< m1 >>
rect 489 451 490 452 
<< m1 >>
rect 19 452 20 453 
<< m1 >>
rect 21 452 22 453 
<< m1 >>
rect 26 452 27 453 
<< m1 >>
rect 28 452 29 453 
<< m1 >>
rect 30 452 31 453 
<< m1 >>
rect 55 452 56 453 
<< m1 >>
rect 73 452 74 453 
<< m2 >>
rect 99 452 100 453 
<< m1 >>
rect 100 452 101 453 
<< m1 >>
rect 150 452 151 453 
<< m1 >>
rect 152 452 153 453 
<< m1 >>
rect 154 452 155 453 
<< m1 >>
rect 160 452 161 453 
<< m1 >>
rect 161 452 162 453 
<< m1 >>
rect 162 452 163 453 
<< m1 >>
rect 163 452 164 453 
<< m2 >>
rect 163 452 164 453 
<< m1 >>
rect 164 452 165 453 
<< m1 >>
rect 165 452 166 453 
<< m1 >>
rect 166 452 167 453 
<< m1 >>
rect 167 452 168 453 
<< m1 >>
rect 168 452 169 453 
<< m1 >>
rect 169 452 170 453 
<< m1 >>
rect 170 452 171 453 
<< m1 >>
rect 171 452 172 453 
<< m1 >>
rect 172 452 173 453 
<< m2 >>
rect 172 452 173 453 
<< m1 >>
rect 194 452 195 453 
<< m2 >>
rect 194 452 195 453 
<< m2c >>
rect 194 452 195 453 
<< m1 >>
rect 194 452 195 453 
<< m2 >>
rect 194 452 195 453 
<< m2 >>
rect 195 452 196 453 
<< m1 >>
rect 196 452 197 453 
<< m2 >>
rect 196 452 197 453 
<< m2 >>
rect 197 452 198 453 
<< m2 >>
rect 208 452 209 453 
<< m2 >>
rect 209 452 210 453 
<< m1 >>
rect 210 452 211 453 
<< m2 >>
rect 210 452 211 453 
<< m2c >>
rect 210 452 211 453 
<< m1 >>
rect 210 452 211 453 
<< m2 >>
rect 210 452 211 453 
<< m1 >>
rect 217 452 218 453 
<< m1 >>
rect 229 452 230 453 
<< m1 >>
rect 253 452 254 453 
<< m2 >>
rect 254 452 255 453 
<< m1 >>
rect 283 452 284 453 
<< m2 >>
rect 283 452 284 453 
<< m2c >>
rect 283 452 284 453 
<< m1 >>
rect 283 452 284 453 
<< m2 >>
rect 283 452 284 453 
<< m1 >>
rect 289 452 290 453 
<< m1 >>
rect 298 452 299 453 
<< m1 >>
rect 307 452 308 453 
<< m1 >>
rect 319 452 320 453 
<< m1 >>
rect 320 452 321 453 
<< m1 >>
rect 321 452 322 453 
<< m1 >>
rect 322 452 323 453 
<< m1 >>
rect 323 452 324 453 
<< m1 >>
rect 324 452 325 453 
<< m1 >>
rect 325 452 326 453 
<< m1 >>
rect 361 452 362 453 
<< m1 >>
rect 373 452 374 453 
<< m1 >>
rect 374 452 375 453 
<< m1 >>
rect 375 452 376 453 
<< m1 >>
rect 376 452 377 453 
<< m1 >>
rect 377 452 378 453 
<< m2 >>
rect 377 452 378 453 
<< m2c >>
rect 377 452 378 453 
<< m1 >>
rect 377 452 378 453 
<< m2 >>
rect 377 452 378 453 
<< m2 >>
rect 378 452 379 453 
<< m1 >>
rect 379 452 380 453 
<< m2 >>
rect 379 452 380 453 
<< m2 >>
rect 380 452 381 453 
<< m1 >>
rect 381 452 382 453 
<< m2 >>
rect 381 452 382 453 
<< m2 >>
rect 382 452 383 453 
<< m1 >>
rect 383 452 384 453 
<< m2 >>
rect 383 452 384 453 
<< m2c >>
rect 383 452 384 453 
<< m1 >>
rect 383 452 384 453 
<< m2 >>
rect 383 452 384 453 
<< m1 >>
rect 384 452 385 453 
<< m1 >>
rect 385 452 386 453 
<< m2 >>
rect 397 452 398 453 
<< m2 >>
rect 402 452 403 453 
<< m2 >>
rect 406 452 407 453 
<< m1 >>
rect 424 452 425 453 
<< m1 >>
rect 425 452 426 453 
<< m1 >>
rect 426 452 427 453 
<< m2 >>
rect 426 452 427 453 
<< m2c >>
rect 426 452 427 453 
<< m1 >>
rect 426 452 427 453 
<< m2 >>
rect 426 452 427 453 
<< m1 >>
rect 431 452 432 453 
<< m1 >>
rect 433 452 434 453 
<< m1 >>
rect 450 452 451 453 
<< m1 >>
rect 452 452 453 453 
<< m1 >>
rect 472 452 473 453 
<< m2 >>
rect 478 452 479 453 
<< m1 >>
rect 487 452 488 453 
<< m1 >>
rect 489 452 490 453 
<< m1 >>
rect 19 453 20 454 
<< m1 >>
rect 21 453 22 454 
<< m1 >>
rect 26 453 27 454 
<< m2 >>
rect 26 453 27 454 
<< m2c >>
rect 26 453 27 454 
<< m1 >>
rect 26 453 27 454 
<< m2 >>
rect 26 453 27 454 
<< m2 >>
rect 27 453 28 454 
<< m1 >>
rect 28 453 29 454 
<< m1 >>
rect 30 453 31 454 
<< m1 >>
rect 55 453 56 454 
<< m1 >>
rect 73 453 74 454 
<< m2 >>
rect 99 453 100 454 
<< m1 >>
rect 100 453 101 454 
<< m1 >>
rect 150 453 151 454 
<< m1 >>
rect 152 453 153 454 
<< m1 >>
rect 154 453 155 454 
<< m2 >>
rect 159 453 160 454 
<< m1 >>
rect 160 453 161 454 
<< m2 >>
rect 160 453 161 454 
<< m2 >>
rect 161 453 162 454 
<< m2 >>
rect 162 453 163 454 
<< m2 >>
rect 163 453 164 454 
<< m2 >>
rect 172 453 173 454 
<< m1 >>
rect 194 453 195 454 
<< m1 >>
rect 196 453 197 454 
<< m1 >>
rect 210 453 211 454 
<< m1 >>
rect 217 453 218 454 
<< m1 >>
rect 229 453 230 454 
<< m1 >>
rect 253 453 254 454 
<< m2 >>
rect 254 453 255 454 
<< m2 >>
rect 283 453 284 454 
<< m1 >>
rect 289 453 290 454 
<< m1 >>
rect 298 453 299 454 
<< m1 >>
rect 307 453 308 454 
<< m1 >>
rect 361 453 362 454 
<< m1 >>
rect 379 453 380 454 
<< m1 >>
rect 381 453 382 454 
<< m2 >>
rect 397 453 398 454 
<< m2 >>
rect 402 453 403 454 
<< m2 >>
rect 406 453 407 454 
<< m2 >>
rect 426 453 427 454 
<< m1 >>
rect 431 453 432 454 
<< m1 >>
rect 433 453 434 454 
<< m1 >>
rect 450 453 451 454 
<< m1 >>
rect 452 453 453 454 
<< m1 >>
rect 470 453 471 454 
<< m2 >>
rect 470 453 471 454 
<< m2c >>
rect 470 453 471 454 
<< m1 >>
rect 470 453 471 454 
<< m2 >>
rect 470 453 471 454 
<< m2 >>
rect 471 453 472 454 
<< m1 >>
rect 472 453 473 454 
<< m2 >>
rect 472 453 473 454 
<< m2 >>
rect 473 453 474 454 
<< m1 >>
rect 474 453 475 454 
<< m2 >>
rect 474 453 475 454 
<< m2c >>
rect 474 453 475 454 
<< m1 >>
rect 474 453 475 454 
<< m2 >>
rect 474 453 475 454 
<< m1 >>
rect 475 453 476 454 
<< m1 >>
rect 476 453 477 454 
<< m1 >>
rect 477 453 478 454 
<< m1 >>
rect 478 453 479 454 
<< m2 >>
rect 478 453 479 454 
<< m2c >>
rect 478 453 479 454 
<< m1 >>
rect 478 453 479 454 
<< m2 >>
rect 478 453 479 454 
<< m1 >>
rect 487 453 488 454 
<< m1 >>
rect 489 453 490 454 
<< m1 >>
rect 19 454 20 455 
<< m1 >>
rect 21 454 22 455 
<< m2 >>
rect 27 454 28 455 
<< m1 >>
rect 28 454 29 455 
<< m2 >>
rect 28 454 29 455 
<< m2 >>
rect 29 454 30 455 
<< m1 >>
rect 30 454 31 455 
<< m2 >>
rect 30 454 31 455 
<< m2 >>
rect 31 454 32 455 
<< m1 >>
rect 32 454 33 455 
<< m2 >>
rect 32 454 33 455 
<< m2c >>
rect 32 454 33 455 
<< m1 >>
rect 32 454 33 455 
<< m2 >>
rect 32 454 33 455 
<< m1 >>
rect 33 454 34 455 
<< m1 >>
rect 34 454 35 455 
<< m1 >>
rect 35 454 36 455 
<< m1 >>
rect 36 454 37 455 
<< m1 >>
rect 37 454 38 455 
<< m1 >>
rect 38 454 39 455 
<< m1 >>
rect 39 454 40 455 
<< m1 >>
rect 40 454 41 455 
<< m1 >>
rect 41 454 42 455 
<< m1 >>
rect 42 454 43 455 
<< m1 >>
rect 43 454 44 455 
<< m1 >>
rect 44 454 45 455 
<< m1 >>
rect 45 454 46 455 
<< m1 >>
rect 46 454 47 455 
<< m1 >>
rect 47 454 48 455 
<< m1 >>
rect 48 454 49 455 
<< m1 >>
rect 49 454 50 455 
<< m1 >>
rect 50 454 51 455 
<< m1 >>
rect 51 454 52 455 
<< m1 >>
rect 52 454 53 455 
<< m1 >>
rect 53 454 54 455 
<< m1 >>
rect 54 454 55 455 
<< m1 >>
rect 55 454 56 455 
<< m1 >>
rect 73 454 74 455 
<< m2 >>
rect 99 454 100 455 
<< m1 >>
rect 100 454 101 455 
<< m2 >>
rect 100 454 101 455 
<< m2 >>
rect 101 454 102 455 
<< m2 >>
rect 102 454 103 455 
<< m1 >>
rect 103 454 104 455 
<< m2 >>
rect 103 454 104 455 
<< m1 >>
rect 104 454 105 455 
<< m2 >>
rect 104 454 105 455 
<< m1 >>
rect 105 454 106 455 
<< m2 >>
rect 105 454 106 455 
<< m1 >>
rect 106 454 107 455 
<< m2 >>
rect 106 454 107 455 
<< m1 >>
rect 107 454 108 455 
<< m2 >>
rect 107 454 108 455 
<< m1 >>
rect 108 454 109 455 
<< m2 >>
rect 108 454 109 455 
<< m1 >>
rect 109 454 110 455 
<< m2 >>
rect 109 454 110 455 
<< m1 >>
rect 110 454 111 455 
<< m2 >>
rect 110 454 111 455 
<< m1 >>
rect 111 454 112 455 
<< m2 >>
rect 111 454 112 455 
<< m1 >>
rect 112 454 113 455 
<< m2 >>
rect 112 454 113 455 
<< m1 >>
rect 113 454 114 455 
<< m2 >>
rect 113 454 114 455 
<< m1 >>
rect 114 454 115 455 
<< m2 >>
rect 114 454 115 455 
<< m1 >>
rect 115 454 116 455 
<< m2 >>
rect 115 454 116 455 
<< m1 >>
rect 116 454 117 455 
<< m2 >>
rect 116 454 117 455 
<< m1 >>
rect 117 454 118 455 
<< m2 >>
rect 117 454 118 455 
<< m1 >>
rect 118 454 119 455 
<< m2 >>
rect 118 454 119 455 
<< m1 >>
rect 119 454 120 455 
<< m2 >>
rect 119 454 120 455 
<< m1 >>
rect 120 454 121 455 
<< m2 >>
rect 120 454 121 455 
<< m1 >>
rect 121 454 122 455 
<< m2 >>
rect 121 454 122 455 
<< m1 >>
rect 122 454 123 455 
<< m2 >>
rect 122 454 123 455 
<< m1 >>
rect 123 454 124 455 
<< m2 >>
rect 123 454 124 455 
<< m1 >>
rect 124 454 125 455 
<< m2 >>
rect 124 454 125 455 
<< m1 >>
rect 125 454 126 455 
<< m2 >>
rect 125 454 126 455 
<< m1 >>
rect 126 454 127 455 
<< m2 >>
rect 126 454 127 455 
<< m1 >>
rect 127 454 128 455 
<< m2 >>
rect 127 454 128 455 
<< m1 >>
rect 128 454 129 455 
<< m2 >>
rect 128 454 129 455 
<< m1 >>
rect 129 454 130 455 
<< m2 >>
rect 129 454 130 455 
<< m1 >>
rect 130 454 131 455 
<< m2 >>
rect 130 454 131 455 
<< m1 >>
rect 131 454 132 455 
<< m2 >>
rect 131 454 132 455 
<< m1 >>
rect 132 454 133 455 
<< m2 >>
rect 132 454 133 455 
<< m1 >>
rect 133 454 134 455 
<< m2 >>
rect 133 454 134 455 
<< m1 >>
rect 134 454 135 455 
<< m2 >>
rect 134 454 135 455 
<< m1 >>
rect 135 454 136 455 
<< m2 >>
rect 135 454 136 455 
<< m1 >>
rect 136 454 137 455 
<< m2 >>
rect 136 454 137 455 
<< m1 >>
rect 137 454 138 455 
<< m2 >>
rect 137 454 138 455 
<< m1 >>
rect 138 454 139 455 
<< m2 >>
rect 138 454 139 455 
<< m1 >>
rect 139 454 140 455 
<< m2 >>
rect 139 454 140 455 
<< m1 >>
rect 140 454 141 455 
<< m2 >>
rect 140 454 141 455 
<< m1 >>
rect 141 454 142 455 
<< m2 >>
rect 141 454 142 455 
<< m1 >>
rect 142 454 143 455 
<< m2 >>
rect 142 454 143 455 
<< m1 >>
rect 143 454 144 455 
<< m2 >>
rect 143 454 144 455 
<< m1 >>
rect 144 454 145 455 
<< m2 >>
rect 144 454 145 455 
<< m1 >>
rect 145 454 146 455 
<< m2 >>
rect 145 454 146 455 
<< m1 >>
rect 146 454 147 455 
<< m2 >>
rect 146 454 147 455 
<< m1 >>
rect 147 454 148 455 
<< m2 >>
rect 147 454 148 455 
<< m1 >>
rect 148 454 149 455 
<< m2 >>
rect 148 454 149 455 
<< m1 >>
rect 149 454 150 455 
<< m2 >>
rect 149 454 150 455 
<< m1 >>
rect 150 454 151 455 
<< m2 >>
rect 150 454 151 455 
<< m2 >>
rect 151 454 152 455 
<< m1 >>
rect 152 454 153 455 
<< m1 >>
rect 154 454 155 455 
<< m1 >>
rect 155 454 156 455 
<< m1 >>
rect 156 454 157 455 
<< m1 >>
rect 157 454 158 455 
<< m1 >>
rect 158 454 159 455 
<< m2 >>
rect 158 454 159 455 
<< m2c >>
rect 158 454 159 455 
<< m1 >>
rect 158 454 159 455 
<< m2 >>
rect 158 454 159 455 
<< m2 >>
rect 159 454 160 455 
<< m1 >>
rect 160 454 161 455 
<< m1 >>
rect 172 454 173 455 
<< m2 >>
rect 172 454 173 455 
<< m1 >>
rect 173 454 174 455 
<< m1 >>
rect 174 454 175 455 
<< m1 >>
rect 175 454 176 455 
<< m1 >>
rect 176 454 177 455 
<< m1 >>
rect 177 454 178 455 
<< m1 >>
rect 178 454 179 455 
<< m1 >>
rect 179 454 180 455 
<< m1 >>
rect 180 454 181 455 
<< m1 >>
rect 181 454 182 455 
<< m1 >>
rect 182 454 183 455 
<< m1 >>
rect 183 454 184 455 
<< m1 >>
rect 184 454 185 455 
<< m1 >>
rect 185 454 186 455 
<< m1 >>
rect 186 454 187 455 
<< m1 >>
rect 187 454 188 455 
<< m1 >>
rect 188 454 189 455 
<< m1 >>
rect 189 454 190 455 
<< m1 >>
rect 190 454 191 455 
<< m1 >>
rect 191 454 192 455 
<< m1 >>
rect 192 454 193 455 
<< m1 >>
rect 193 454 194 455 
<< m1 >>
rect 194 454 195 455 
<< m1 >>
rect 196 454 197 455 
<< m2 >>
rect 209 454 210 455 
<< m1 >>
rect 210 454 211 455 
<< m2 >>
rect 210 454 211 455 
<< m2 >>
rect 211 454 212 455 
<< m1 >>
rect 212 454 213 455 
<< m2 >>
rect 212 454 213 455 
<< m2c >>
rect 212 454 213 455 
<< m1 >>
rect 212 454 213 455 
<< m2 >>
rect 212 454 213 455 
<< m1 >>
rect 213 454 214 455 
<< m1 >>
rect 214 454 215 455 
<< m1 >>
rect 215 454 216 455 
<< m1 >>
rect 216 454 217 455 
<< m1 >>
rect 217 454 218 455 
<< m1 >>
rect 229 454 230 455 
<< m1 >>
rect 253 454 254 455 
<< m2 >>
rect 254 454 255 455 
<< m1 >>
rect 255 454 256 455 
<< m2 >>
rect 255 454 256 455 
<< m2c >>
rect 255 454 256 455 
<< m1 >>
rect 255 454 256 455 
<< m2 >>
rect 255 454 256 455 
<< m1 >>
rect 256 454 257 455 
<< m1 >>
rect 257 454 258 455 
<< m1 >>
rect 258 454 259 455 
<< m1 >>
rect 259 454 260 455 
<< m1 >>
rect 260 454 261 455 
<< m1 >>
rect 261 454 262 455 
<< m1 >>
rect 262 454 263 455 
<< m1 >>
rect 263 454 264 455 
<< m1 >>
rect 264 454 265 455 
<< m1 >>
rect 265 454 266 455 
<< m1 >>
rect 266 454 267 455 
<< m1 >>
rect 267 454 268 455 
<< m1 >>
rect 268 454 269 455 
<< m1 >>
rect 269 454 270 455 
<< m1 >>
rect 270 454 271 455 
<< m1 >>
rect 271 454 272 455 
<< m1 >>
rect 272 454 273 455 
<< m1 >>
rect 273 454 274 455 
<< m1 >>
rect 274 454 275 455 
<< m1 >>
rect 275 454 276 455 
<< m1 >>
rect 276 454 277 455 
<< m1 >>
rect 277 454 278 455 
<< m1 >>
rect 278 454 279 455 
<< m1 >>
rect 279 454 280 455 
<< m1 >>
rect 280 454 281 455 
<< m1 >>
rect 281 454 282 455 
<< m1 >>
rect 282 454 283 455 
<< m1 >>
rect 283 454 284 455 
<< m2 >>
rect 283 454 284 455 
<< m1 >>
rect 284 454 285 455 
<< m1 >>
rect 285 454 286 455 
<< m1 >>
rect 286 454 287 455 
<< m1 >>
rect 287 454 288 455 
<< m2 >>
rect 287 454 288 455 
<< m2c >>
rect 287 454 288 455 
<< m1 >>
rect 287 454 288 455 
<< m2 >>
rect 287 454 288 455 
<< m2 >>
rect 288 454 289 455 
<< m1 >>
rect 289 454 290 455 
<< m2 >>
rect 289 454 290 455 
<< m2 >>
rect 290 454 291 455 
<< m1 >>
rect 291 454 292 455 
<< m2 >>
rect 291 454 292 455 
<< m2c >>
rect 291 454 292 455 
<< m1 >>
rect 291 454 292 455 
<< m2 >>
rect 291 454 292 455 
<< m1 >>
rect 292 454 293 455 
<< m1 >>
rect 293 454 294 455 
<< m1 >>
rect 294 454 295 455 
<< m1 >>
rect 295 454 296 455 
<< m1 >>
rect 296 454 297 455 
<< m2 >>
rect 296 454 297 455 
<< m2c >>
rect 296 454 297 455 
<< m1 >>
rect 296 454 297 455 
<< m2 >>
rect 296 454 297 455 
<< m2 >>
rect 297 454 298 455 
<< m1 >>
rect 298 454 299 455 
<< m2 >>
rect 298 454 299 455 
<< m2 >>
rect 299 454 300 455 
<< m1 >>
rect 300 454 301 455 
<< m2 >>
rect 300 454 301 455 
<< m2c >>
rect 300 454 301 455 
<< m1 >>
rect 300 454 301 455 
<< m2 >>
rect 300 454 301 455 
<< m1 >>
rect 301 454 302 455 
<< m1 >>
rect 302 454 303 455 
<< m1 >>
rect 303 454 304 455 
<< m1 >>
rect 304 454 305 455 
<< m1 >>
rect 305 454 306 455 
<< m2 >>
rect 305 454 306 455 
<< m2c >>
rect 305 454 306 455 
<< m1 >>
rect 305 454 306 455 
<< m2 >>
rect 305 454 306 455 
<< m2 >>
rect 306 454 307 455 
<< m1 >>
rect 307 454 308 455 
<< m2 >>
rect 307 454 308 455 
<< m2 >>
rect 308 454 309 455 
<< m1 >>
rect 309 454 310 455 
<< m2 >>
rect 309 454 310 455 
<< m2c >>
rect 309 454 310 455 
<< m1 >>
rect 309 454 310 455 
<< m2 >>
rect 309 454 310 455 
<< m1 >>
rect 310 454 311 455 
<< m1 >>
rect 311 454 312 455 
<< m1 >>
rect 312 454 313 455 
<< m1 >>
rect 313 454 314 455 
<< m1 >>
rect 314 454 315 455 
<< m1 >>
rect 315 454 316 455 
<< m1 >>
rect 316 454 317 455 
<< m1 >>
rect 317 454 318 455 
<< m1 >>
rect 318 454 319 455 
<< m1 >>
rect 319 454 320 455 
<< m1 >>
rect 320 454 321 455 
<< m1 >>
rect 321 454 322 455 
<< m1 >>
rect 322 454 323 455 
<< m1 >>
rect 323 454 324 455 
<< m1 >>
rect 324 454 325 455 
<< m1 >>
rect 325 454 326 455 
<< m1 >>
rect 326 454 327 455 
<< m1 >>
rect 327 454 328 455 
<< m1 >>
rect 328 454 329 455 
<< m1 >>
rect 329 454 330 455 
<< m1 >>
rect 330 454 331 455 
<< m1 >>
rect 331 454 332 455 
<< m1 >>
rect 332 454 333 455 
<< m1 >>
rect 333 454 334 455 
<< m1 >>
rect 334 454 335 455 
<< m1 >>
rect 335 454 336 455 
<< m1 >>
rect 336 454 337 455 
<< m1 >>
rect 337 454 338 455 
<< m1 >>
rect 338 454 339 455 
<< m1 >>
rect 339 454 340 455 
<< m1 >>
rect 340 454 341 455 
<< m1 >>
rect 341 454 342 455 
<< m1 >>
rect 342 454 343 455 
<< m1 >>
rect 343 454 344 455 
<< m1 >>
rect 344 454 345 455 
<< m1 >>
rect 345 454 346 455 
<< m1 >>
rect 346 454 347 455 
<< m1 >>
rect 347 454 348 455 
<< m1 >>
rect 348 454 349 455 
<< m1 >>
rect 349 454 350 455 
<< m1 >>
rect 350 454 351 455 
<< m1 >>
rect 351 454 352 455 
<< m1 >>
rect 352 454 353 455 
<< m1 >>
rect 353 454 354 455 
<< m1 >>
rect 354 454 355 455 
<< m1 >>
rect 355 454 356 455 
<< m1 >>
rect 356 454 357 455 
<< m1 >>
rect 357 454 358 455 
<< m1 >>
rect 358 454 359 455 
<< m1 >>
rect 359 454 360 455 
<< m2 >>
rect 359 454 360 455 
<< m2c >>
rect 359 454 360 455 
<< m1 >>
rect 359 454 360 455 
<< m2 >>
rect 359 454 360 455 
<< m2 >>
rect 360 454 361 455 
<< m1 >>
rect 361 454 362 455 
<< m2 >>
rect 361 454 362 455 
<< m2 >>
rect 362 454 363 455 
<< m1 >>
rect 363 454 364 455 
<< m2 >>
rect 363 454 364 455 
<< m2c >>
rect 363 454 364 455 
<< m1 >>
rect 363 454 364 455 
<< m2 >>
rect 363 454 364 455 
<< m1 >>
rect 364 454 365 455 
<< m1 >>
rect 365 454 366 455 
<< m1 >>
rect 366 454 367 455 
<< m1 >>
rect 367 454 368 455 
<< m1 >>
rect 368 454 369 455 
<< m1 >>
rect 369 454 370 455 
<< m1 >>
rect 370 454 371 455 
<< m1 >>
rect 371 454 372 455 
<< m1 >>
rect 372 454 373 455 
<< m1 >>
rect 373 454 374 455 
<< m1 >>
rect 374 454 375 455 
<< m1 >>
rect 375 454 376 455 
<< m1 >>
rect 376 454 377 455 
<< m1 >>
rect 377 454 378 455 
<< m1 >>
rect 378 454 379 455 
<< m1 >>
rect 379 454 380 455 
<< m1 >>
rect 381 454 382 455 
<< m1 >>
rect 394 454 395 455 
<< m1 >>
rect 395 454 396 455 
<< m1 >>
rect 396 454 397 455 
<< m1 >>
rect 397 454 398 455 
<< m2 >>
rect 397 454 398 455 
<< m1 >>
rect 398 454 399 455 
<< m1 >>
rect 399 454 400 455 
<< m1 >>
rect 400 454 401 455 
<< m1 >>
rect 401 454 402 455 
<< m1 >>
rect 402 454 403 455 
<< m2 >>
rect 402 454 403 455 
<< m1 >>
rect 403 454 404 455 
<< m1 >>
rect 404 454 405 455 
<< m1 >>
rect 405 454 406 455 
<< m1 >>
rect 406 454 407 455 
<< m2 >>
rect 406 454 407 455 
<< m1 >>
rect 407 454 408 455 
<< m1 >>
rect 408 454 409 455 
<< m1 >>
rect 409 454 410 455 
<< m1 >>
rect 410 454 411 455 
<< m1 >>
rect 411 454 412 455 
<< m1 >>
rect 412 454 413 455 
<< m1 >>
rect 413 454 414 455 
<< m1 >>
rect 414 454 415 455 
<< m1 >>
rect 415 454 416 455 
<< m1 >>
rect 416 454 417 455 
<< m1 >>
rect 417 454 418 455 
<< m1 >>
rect 418 454 419 455 
<< m1 >>
rect 419 454 420 455 
<< m1 >>
rect 420 454 421 455 
<< m1 >>
rect 421 454 422 455 
<< m1 >>
rect 422 454 423 455 
<< m1 >>
rect 423 454 424 455 
<< m1 >>
rect 424 454 425 455 
<< m1 >>
rect 425 454 426 455 
<< m1 >>
rect 426 454 427 455 
<< m2 >>
rect 426 454 427 455 
<< m1 >>
rect 427 454 428 455 
<< m2 >>
rect 427 454 428 455 
<< m1 >>
rect 428 454 429 455 
<< m2 >>
rect 428 454 429 455 
<< m1 >>
rect 429 454 430 455 
<< m2 >>
rect 429 454 430 455 
<< m1 >>
rect 430 454 431 455 
<< m2 >>
rect 430 454 431 455 
<< m1 >>
rect 431 454 432 455 
<< m2 >>
rect 431 454 432 455 
<< m2 >>
rect 432 454 433 455 
<< m1 >>
rect 433 454 434 455 
<< m2 >>
rect 433 454 434 455 
<< m2 >>
rect 434 454 435 455 
<< m1 >>
rect 435 454 436 455 
<< m2 >>
rect 435 454 436 455 
<< m2c >>
rect 435 454 436 455 
<< m1 >>
rect 435 454 436 455 
<< m2 >>
rect 435 454 436 455 
<< m1 >>
rect 436 454 437 455 
<< m1 >>
rect 437 454 438 455 
<< m1 >>
rect 438 454 439 455 
<< m1 >>
rect 439 454 440 455 
<< m1 >>
rect 440 454 441 455 
<< m1 >>
rect 441 454 442 455 
<< m1 >>
rect 442 454 443 455 
<< m1 >>
rect 443 454 444 455 
<< m1 >>
rect 444 454 445 455 
<< m1 >>
rect 445 454 446 455 
<< m1 >>
rect 446 454 447 455 
<< m1 >>
rect 447 454 448 455 
<< m1 >>
rect 448 454 449 455 
<< m1 >>
rect 449 454 450 455 
<< m1 >>
rect 450 454 451 455 
<< m1 >>
rect 452 454 453 455 
<< m2 >>
rect 453 454 454 455 
<< m1 >>
rect 454 454 455 455 
<< m2 >>
rect 454 454 455 455 
<< m2c >>
rect 454 454 455 455 
<< m1 >>
rect 454 454 455 455 
<< m2 >>
rect 454 454 455 455 
<< m1 >>
rect 455 454 456 455 
<< m1 >>
rect 456 454 457 455 
<< m1 >>
rect 457 454 458 455 
<< m1 >>
rect 458 454 459 455 
<< m1 >>
rect 459 454 460 455 
<< m1 >>
rect 460 454 461 455 
<< m1 >>
rect 461 454 462 455 
<< m1 >>
rect 462 454 463 455 
<< m1 >>
rect 463 454 464 455 
<< m1 >>
rect 464 454 465 455 
<< m1 >>
rect 465 454 466 455 
<< m1 >>
rect 466 454 467 455 
<< m1 >>
rect 467 454 468 455 
<< m1 >>
rect 468 454 469 455 
<< m1 >>
rect 469 454 470 455 
<< m1 >>
rect 470 454 471 455 
<< m1 >>
rect 472 454 473 455 
<< m1 >>
rect 487 454 488 455 
<< m1 >>
rect 489 454 490 455 
<< m1 >>
rect 19 455 20 456 
<< m1 >>
rect 21 455 22 456 
<< m1 >>
rect 28 455 29 456 
<< m1 >>
rect 30 455 31 456 
<< m1 >>
rect 73 455 74 456 
<< m1 >>
rect 100 455 101 456 
<< m1 >>
rect 103 455 104 456 
<< m2 >>
rect 151 455 152 456 
<< m1 >>
rect 152 455 153 456 
<< m1 >>
rect 160 455 161 456 
<< m1 >>
rect 172 455 173 456 
<< m2 >>
rect 172 455 173 456 
<< m1 >>
rect 196 455 197 456 
<< m2 >>
rect 209 455 210 456 
<< m1 >>
rect 210 455 211 456 
<< m1 >>
rect 229 455 230 456 
<< m1 >>
rect 253 455 254 456 
<< m2 >>
rect 283 455 284 456 
<< m1 >>
rect 289 455 290 456 
<< m1 >>
rect 298 455 299 456 
<< m1 >>
rect 307 455 308 456 
<< m1 >>
rect 361 455 362 456 
<< m1 >>
rect 381 455 382 456 
<< m1 >>
rect 394 455 395 456 
<< m2 >>
rect 397 455 398 456 
<< m2 >>
rect 402 455 403 456 
<< m2 >>
rect 406 455 407 456 
<< m1 >>
rect 433 455 434 456 
<< m1 >>
rect 452 455 453 456 
<< m2 >>
rect 453 455 454 456 
<< m1 >>
rect 472 455 473 456 
<< m1 >>
rect 487 455 488 456 
<< m1 >>
rect 489 455 490 456 
<< m1 >>
rect 19 456 20 457 
<< m1 >>
rect 21 456 22 457 
<< m1 >>
rect 28 456 29 457 
<< m1 >>
rect 30 456 31 457 
<< m1 >>
rect 73 456 74 457 
<< m1 >>
rect 100 456 101 457 
<< m1 >>
rect 103 456 104 457 
<< m2 >>
rect 151 456 152 457 
<< m1 >>
rect 152 456 153 457 
<< m2 >>
rect 152 456 153 457 
<< m2 >>
rect 153 456 154 457 
<< m1 >>
rect 154 456 155 457 
<< m2 >>
rect 154 456 155 457 
<< m2c >>
rect 154 456 155 457 
<< m1 >>
rect 154 456 155 457 
<< m2 >>
rect 154 456 155 457 
<< m1 >>
rect 155 456 156 457 
<< m1 >>
rect 156 456 157 457 
<< m1 >>
rect 157 456 158 457 
<< m1 >>
rect 158 456 159 457 
<< m2 >>
rect 158 456 159 457 
<< m2c >>
rect 158 456 159 457 
<< m1 >>
rect 158 456 159 457 
<< m2 >>
rect 158 456 159 457 
<< m2 >>
rect 159 456 160 457 
<< m1 >>
rect 160 456 161 457 
<< m2 >>
rect 160 456 161 457 
<< m2 >>
rect 161 456 162 457 
<< m1 >>
rect 162 456 163 457 
<< m2 >>
rect 162 456 163 457 
<< m2c >>
rect 162 456 163 457 
<< m1 >>
rect 162 456 163 457 
<< m2 >>
rect 162 456 163 457 
<< m1 >>
rect 163 456 164 457 
<< m1 >>
rect 172 456 173 457 
<< m2 >>
rect 172 456 173 457 
<< m1 >>
rect 196 456 197 457 
<< m2 >>
rect 209 456 210 457 
<< m1 >>
rect 210 456 211 457 
<< m1 >>
rect 211 456 212 457 
<< m1 >>
rect 212 456 213 457 
<< m1 >>
rect 213 456 214 457 
<< m1 >>
rect 214 456 215 457 
<< m1 >>
rect 215 456 216 457 
<< m1 >>
rect 216 456 217 457 
<< m1 >>
rect 217 456 218 457 
<< m1 >>
rect 218 456 219 457 
<< m1 >>
rect 219 456 220 457 
<< m1 >>
rect 220 456 221 457 
<< m1 >>
rect 221 456 222 457 
<< m1 >>
rect 222 456 223 457 
<< m1 >>
rect 223 456 224 457 
<< m1 >>
rect 224 456 225 457 
<< m1 >>
rect 225 456 226 457 
<< m1 >>
rect 226 456 227 457 
<< m1 >>
rect 227 456 228 457 
<< m2 >>
rect 227 456 228 457 
<< m2c >>
rect 227 456 228 457 
<< m1 >>
rect 227 456 228 457 
<< m2 >>
rect 227 456 228 457 
<< m2 >>
rect 228 456 229 457 
<< m1 >>
rect 229 456 230 457 
<< m2 >>
rect 229 456 230 457 
<< m2 >>
rect 230 456 231 457 
<< m1 >>
rect 231 456 232 457 
<< m2 >>
rect 231 456 232 457 
<< m2c >>
rect 231 456 232 457 
<< m1 >>
rect 231 456 232 457 
<< m2 >>
rect 231 456 232 457 
<< m1 >>
rect 232 456 233 457 
<< m1 >>
rect 233 456 234 457 
<< m1 >>
rect 234 456 235 457 
<< m1 >>
rect 235 456 236 457 
<< m1 >>
rect 236 456 237 457 
<< m1 >>
rect 237 456 238 457 
<< m1 >>
rect 238 456 239 457 
<< m1 >>
rect 239 456 240 457 
<< m1 >>
rect 240 456 241 457 
<< m1 >>
rect 241 456 242 457 
<< m1 >>
rect 242 456 243 457 
<< m1 >>
rect 243 456 244 457 
<< m1 >>
rect 244 456 245 457 
<< m1 >>
rect 245 456 246 457 
<< m1 >>
rect 246 456 247 457 
<< m1 >>
rect 247 456 248 457 
<< m1 >>
rect 248 456 249 457 
<< m1 >>
rect 249 456 250 457 
<< m1 >>
rect 250 456 251 457 
<< m1 >>
rect 251 456 252 457 
<< m2 >>
rect 251 456 252 457 
<< m2c >>
rect 251 456 252 457 
<< m1 >>
rect 251 456 252 457 
<< m2 >>
rect 251 456 252 457 
<< m2 >>
rect 252 456 253 457 
<< m1 >>
rect 253 456 254 457 
<< m2 >>
rect 253 456 254 457 
<< m2 >>
rect 254 456 255 457 
<< m1 >>
rect 255 456 256 457 
<< m2 >>
rect 255 456 256 457 
<< m2c >>
rect 255 456 256 457 
<< m1 >>
rect 255 456 256 457 
<< m2 >>
rect 255 456 256 457 
<< m1 >>
rect 256 456 257 457 
<< m1 >>
rect 257 456 258 457 
<< m1 >>
rect 258 456 259 457 
<< m1 >>
rect 259 456 260 457 
<< m1 >>
rect 260 456 261 457 
<< m1 >>
rect 261 456 262 457 
<< m1 >>
rect 262 456 263 457 
<< m1 >>
rect 263 456 264 457 
<< m1 >>
rect 264 456 265 457 
<< m1 >>
rect 265 456 266 457 
<< m1 >>
rect 266 456 267 457 
<< m1 >>
rect 267 456 268 457 
<< m1 >>
rect 268 456 269 457 
<< m1 >>
rect 269 456 270 457 
<< m1 >>
rect 270 456 271 457 
<< m1 >>
rect 271 456 272 457 
<< m1 >>
rect 272 456 273 457 
<< m1 >>
rect 273 456 274 457 
<< m1 >>
rect 274 456 275 457 
<< m1 >>
rect 275 456 276 457 
<< m1 >>
rect 276 456 277 457 
<< m1 >>
rect 277 456 278 457 
<< m1 >>
rect 278 456 279 457 
<< m1 >>
rect 279 456 280 457 
<< m1 >>
rect 280 456 281 457 
<< m1 >>
rect 281 456 282 457 
<< m1 >>
rect 282 456 283 457 
<< m1 >>
rect 283 456 284 457 
<< m2 >>
rect 283 456 284 457 
<< m2c >>
rect 283 456 284 457 
<< m1 >>
rect 283 456 284 457 
<< m2 >>
rect 283 456 284 457 
<< m1 >>
rect 289 456 290 457 
<< m1 >>
rect 298 456 299 457 
<< m1 >>
rect 307 456 308 457 
<< m1 >>
rect 361 456 362 457 
<< m1 >>
rect 381 456 382 457 
<< m1 >>
rect 394 456 395 457 
<< m1 >>
rect 397 456 398 457 
<< m2 >>
rect 397 456 398 457 
<< m2c >>
rect 397 456 398 457 
<< m1 >>
rect 397 456 398 457 
<< m2 >>
rect 397 456 398 457 
<< m1 >>
rect 398 456 399 457 
<< m1 >>
rect 399 456 400 457 
<< m1 >>
rect 400 456 401 457 
<< m1 >>
rect 401 456 402 457 
<< m1 >>
rect 402 456 403 457 
<< m2 >>
rect 402 456 403 457 
<< m1 >>
rect 403 456 404 457 
<< m1 >>
rect 404 456 405 457 
<< m1 >>
rect 405 456 406 457 
<< m1 >>
rect 406 456 407 457 
<< m2 >>
rect 406 456 407 457 
<< m1 >>
rect 407 456 408 457 
<< m2 >>
rect 407 456 408 457 
<< m1 >>
rect 408 456 409 457 
<< m2 >>
rect 408 456 409 457 
<< m1 >>
rect 409 456 410 457 
<< m2 >>
rect 409 456 410 457 
<< m2 >>
rect 410 456 411 457 
<< m1 >>
rect 411 456 412 457 
<< m2 >>
rect 411 456 412 457 
<< m2c >>
rect 411 456 412 457 
<< m1 >>
rect 411 456 412 457 
<< m2 >>
rect 411 456 412 457 
<< m1 >>
rect 412 456 413 457 
<< m1 >>
rect 413 456 414 457 
<< m1 >>
rect 414 456 415 457 
<< m1 >>
rect 415 456 416 457 
<< m1 >>
rect 416 456 417 457 
<< m1 >>
rect 417 456 418 457 
<< m1 >>
rect 418 456 419 457 
<< m1 >>
rect 419 456 420 457 
<< m1 >>
rect 420 456 421 457 
<< m1 >>
rect 421 456 422 457 
<< m1 >>
rect 422 456 423 457 
<< m1 >>
rect 423 456 424 457 
<< m1 >>
rect 424 456 425 457 
<< m1 >>
rect 425 456 426 457 
<< m1 >>
rect 426 456 427 457 
<< m1 >>
rect 427 456 428 457 
<< m1 >>
rect 428 456 429 457 
<< m1 >>
rect 429 456 430 457 
<< m1 >>
rect 430 456 431 457 
<< m1 >>
rect 431 456 432 457 
<< m2 >>
rect 431 456 432 457 
<< m2c >>
rect 431 456 432 457 
<< m1 >>
rect 431 456 432 457 
<< m2 >>
rect 431 456 432 457 
<< m2 >>
rect 432 456 433 457 
<< m1 >>
rect 433 456 434 457 
<< m2 >>
rect 433 456 434 457 
<< m2 >>
rect 434 456 435 457 
<< m1 >>
rect 435 456 436 457 
<< m2 >>
rect 435 456 436 457 
<< m2c >>
rect 435 456 436 457 
<< m1 >>
rect 435 456 436 457 
<< m2 >>
rect 435 456 436 457 
<< m1 >>
rect 436 456 437 457 
<< m1 >>
rect 437 456 438 457 
<< m1 >>
rect 438 456 439 457 
<< m1 >>
rect 439 456 440 457 
<< m1 >>
rect 440 456 441 457 
<< m1 >>
rect 441 456 442 457 
<< m1 >>
rect 442 456 443 457 
<< m1 >>
rect 443 456 444 457 
<< m1 >>
rect 444 456 445 457 
<< m1 >>
rect 445 456 446 457 
<< m1 >>
rect 446 456 447 457 
<< m1 >>
rect 447 456 448 457 
<< m1 >>
rect 448 456 449 457 
<< m1 >>
rect 449 456 450 457 
<< m1 >>
rect 450 456 451 457 
<< m2 >>
rect 450 456 451 457 
<< m2c >>
rect 450 456 451 457 
<< m1 >>
rect 450 456 451 457 
<< m2 >>
rect 450 456 451 457 
<< m2 >>
rect 451 456 452 457 
<< m1 >>
rect 452 456 453 457 
<< m2 >>
rect 452 456 453 457 
<< m2 >>
rect 453 456 454 457 
<< m1 >>
rect 472 456 473 457 
<< m1 >>
rect 487 456 488 457 
<< m1 >>
rect 489 456 490 457 
<< m1 >>
rect 19 457 20 458 
<< m1 >>
rect 21 457 22 458 
<< m1 >>
rect 28 457 29 458 
<< m1 >>
rect 30 457 31 458 
<< m1 >>
rect 73 457 74 458 
<< m1 >>
rect 100 457 101 458 
<< m1 >>
rect 103 457 104 458 
<< m1 >>
rect 152 457 153 458 
<< m1 >>
rect 160 457 161 458 
<< m1 >>
rect 163 457 164 458 
<< m1 >>
rect 172 457 173 458 
<< m2 >>
rect 172 457 173 458 
<< m1 >>
rect 196 457 197 458 
<< m2 >>
rect 209 457 210 458 
<< m1 >>
rect 229 457 230 458 
<< m1 >>
rect 253 457 254 458 
<< m1 >>
rect 289 457 290 458 
<< m1 >>
rect 298 457 299 458 
<< m1 >>
rect 307 457 308 458 
<< m1 >>
rect 352 457 353 458 
<< m1 >>
rect 353 457 354 458 
<< m1 >>
rect 354 457 355 458 
<< m1 >>
rect 355 457 356 458 
<< m1 >>
rect 356 457 357 458 
<< m1 >>
rect 357 457 358 458 
<< m1 >>
rect 358 457 359 458 
<< m1 >>
rect 359 457 360 458 
<< m1 >>
rect 361 457 362 458 
<< m1 >>
rect 381 457 382 458 
<< m1 >>
rect 394 457 395 458 
<< m2 >>
rect 402 457 403 458 
<< m1 >>
rect 409 457 410 458 
<< m1 >>
rect 433 457 434 458 
<< m1 >>
rect 452 457 453 458 
<< m1 >>
rect 472 457 473 458 
<< m1 >>
rect 487 457 488 458 
<< m1 >>
rect 489 457 490 458 
<< m1 >>
rect 19 458 20 459 
<< m1 >>
rect 21 458 22 459 
<< m1 >>
rect 28 458 29 459 
<< m1 >>
rect 30 458 31 459 
<< m1 >>
rect 73 458 74 459 
<< m1 >>
rect 100 458 101 459 
<< m1 >>
rect 103 458 104 459 
<< m1 >>
rect 152 458 153 459 
<< m1 >>
rect 160 458 161 459 
<< m1 >>
rect 163 458 164 459 
<< m1 >>
rect 172 458 173 459 
<< m2 >>
rect 172 458 173 459 
<< m1 >>
rect 196 458 197 459 
<< m2 >>
rect 209 458 210 459 
<< m1 >>
rect 229 458 230 459 
<< m1 >>
rect 253 458 254 459 
<< m1 >>
rect 289 458 290 459 
<< m1 >>
rect 298 458 299 459 
<< m1 >>
rect 307 458 308 459 
<< m1 >>
rect 352 458 353 459 
<< m1 >>
rect 359 458 360 459 
<< m1 >>
rect 361 458 362 459 
<< m1 >>
rect 381 458 382 459 
<< m1 >>
rect 394 458 395 459 
<< m1 >>
rect 402 458 403 459 
<< m2 >>
rect 402 458 403 459 
<< m2c >>
rect 402 458 403 459 
<< m1 >>
rect 402 458 403 459 
<< m2 >>
rect 402 458 403 459 
<< m1 >>
rect 409 458 410 459 
<< m1 >>
rect 433 458 434 459 
<< m1 >>
rect 451 458 452 459 
<< m2 >>
rect 451 458 452 459 
<< m2c >>
rect 451 458 452 459 
<< m1 >>
rect 451 458 452 459 
<< m2 >>
rect 451 458 452 459 
<< m1 >>
rect 452 458 453 459 
<< m1 >>
rect 472 458 473 459 
<< m1 >>
rect 487 458 488 459 
<< m1 >>
rect 489 458 490 459 
<< m1 >>
rect 19 459 20 460 
<< m1 >>
rect 21 459 22 460 
<< m1 >>
rect 28 459 29 460 
<< m1 >>
rect 30 459 31 460 
<< m1 >>
rect 73 459 74 460 
<< m1 >>
rect 100 459 101 460 
<< m1 >>
rect 103 459 104 460 
<< m1 >>
rect 152 459 153 460 
<< m1 >>
rect 160 459 161 460 
<< m1 >>
rect 163 459 164 460 
<< m1 >>
rect 172 459 173 460 
<< m2 >>
rect 172 459 173 460 
<< m1 >>
rect 196 459 197 460 
<< m1 >>
rect 197 459 198 460 
<< m1 >>
rect 198 459 199 460 
<< m1 >>
rect 199 459 200 460 
<< m1 >>
rect 200 459 201 460 
<< m1 >>
rect 201 459 202 460 
<< m1 >>
rect 202 459 203 460 
<< m1 >>
rect 203 459 204 460 
<< m1 >>
rect 204 459 205 460 
<< m1 >>
rect 205 459 206 460 
<< m1 >>
rect 206 459 207 460 
<< m1 >>
rect 207 459 208 460 
<< m1 >>
rect 208 459 209 460 
<< m2 >>
rect 209 459 210 460 
<< m1 >>
rect 229 459 230 460 
<< m1 >>
rect 253 459 254 460 
<< m1 >>
rect 289 459 290 460 
<< m1 >>
rect 298 459 299 460 
<< m1 >>
rect 307 459 308 460 
<< m1 >>
rect 352 459 353 460 
<< m1 >>
rect 359 459 360 460 
<< m1 >>
rect 361 459 362 460 
<< m1 >>
rect 381 459 382 460 
<< m1 >>
rect 394 459 395 460 
<< m1 >>
rect 402 459 403 460 
<< m1 >>
rect 409 459 410 460 
<< m1 >>
rect 433 459 434 460 
<< m2 >>
rect 451 459 452 460 
<< m1 >>
rect 472 459 473 460 
<< m1 >>
rect 487 459 488 460 
<< m1 >>
rect 489 459 490 460 
<< m1 >>
rect 19 460 20 461 
<< m1 >>
rect 21 460 22 461 
<< m1 >>
rect 28 460 29 461 
<< m1 >>
rect 30 460 31 461 
<< m1 >>
rect 73 460 74 461 
<< m1 >>
rect 100 460 101 461 
<< m1 >>
rect 103 460 104 461 
<< m1 >>
rect 136 460 137 461 
<< m1 >>
rect 137 460 138 461 
<< m1 >>
rect 138 460 139 461 
<< m1 >>
rect 139 460 140 461 
<< m1 >>
rect 152 460 153 461 
<< m1 >>
rect 160 460 161 461 
<< m1 >>
rect 163 460 164 461 
<< m1 >>
rect 172 460 173 461 
<< m2 >>
rect 172 460 173 461 
<< m2 >>
rect 199 460 200 461 
<< m2 >>
rect 200 460 201 461 
<< m2 >>
rect 201 460 202 461 
<< m2 >>
rect 202 460 203 461 
<< m2 >>
rect 203 460 204 461 
<< m2 >>
rect 204 460 205 461 
<< m2 >>
rect 205 460 206 461 
<< m2 >>
rect 206 460 207 461 
<< m2 >>
rect 207 460 208 461 
<< m1 >>
rect 208 460 209 461 
<< m2 >>
rect 208 460 209 461 
<< m2 >>
rect 209 460 210 461 
<< m1 >>
rect 229 460 230 461 
<< m1 >>
rect 253 460 254 461 
<< m1 >>
rect 289 460 290 461 
<< m1 >>
rect 298 460 299 461 
<< m1 >>
rect 307 460 308 461 
<< m1 >>
rect 352 460 353 461 
<< m1 >>
rect 359 460 360 461 
<< m2 >>
rect 359 460 360 461 
<< m2c >>
rect 359 460 360 461 
<< m1 >>
rect 359 460 360 461 
<< m2 >>
rect 359 460 360 461 
<< m2 >>
rect 360 460 361 461 
<< m1 >>
rect 361 460 362 461 
<< m2 >>
rect 361 460 362 461 
<< m2 >>
rect 362 460 363 461 
<< m1 >>
rect 381 460 382 461 
<< m1 >>
rect 394 460 395 461 
<< m1 >>
rect 402 460 403 461 
<< m1 >>
rect 409 460 410 461 
<< m1 >>
rect 433 460 434 461 
<< m1 >>
rect 448 460 449 461 
<< m1 >>
rect 449 460 450 461 
<< m1 >>
rect 450 460 451 461 
<< m1 >>
rect 451 460 452 461 
<< m2 >>
rect 451 460 452 461 
<< m1 >>
rect 472 460 473 461 
<< m1 >>
rect 487 460 488 461 
<< m1 >>
rect 489 460 490 461 
<< m1 >>
rect 19 461 20 462 
<< m1 >>
rect 21 461 22 462 
<< m1 >>
rect 28 461 29 462 
<< m1 >>
rect 30 461 31 462 
<< m1 >>
rect 73 461 74 462 
<< m1 >>
rect 100 461 101 462 
<< m1 >>
rect 103 461 104 462 
<< m1 >>
rect 136 461 137 462 
<< m1 >>
rect 139 461 140 462 
<< m1 >>
rect 152 461 153 462 
<< m1 >>
rect 160 461 161 462 
<< m1 >>
rect 163 461 164 462 
<< m1 >>
rect 172 461 173 462 
<< m2 >>
rect 172 461 173 462 
<< m1 >>
rect 199 461 200 462 
<< m2 >>
rect 199 461 200 462 
<< m2c >>
rect 199 461 200 462 
<< m1 >>
rect 199 461 200 462 
<< m2 >>
rect 199 461 200 462 
<< m1 >>
rect 208 461 209 462 
<< m1 >>
rect 229 461 230 462 
<< m1 >>
rect 253 461 254 462 
<< m1 >>
rect 289 461 290 462 
<< m1 >>
rect 298 461 299 462 
<< m1 >>
rect 307 461 308 462 
<< m1 >>
rect 352 461 353 462 
<< m1 >>
rect 361 461 362 462 
<< m2 >>
rect 362 461 363 462 
<< m1 >>
rect 381 461 382 462 
<< m1 >>
rect 394 461 395 462 
<< m1 >>
rect 402 461 403 462 
<< m1 >>
rect 409 461 410 462 
<< m1 >>
rect 433 461 434 462 
<< m1 >>
rect 448 461 449 462 
<< m1 >>
rect 451 461 452 462 
<< m2 >>
rect 451 461 452 462 
<< m1 >>
rect 472 461 473 462 
<< m1 >>
rect 487 461 488 462 
<< m1 >>
rect 489 461 490 462 
<< pdiffusion >>
rect 12 462 13 463 
<< pdiffusion >>
rect 13 462 14 463 
<< pdiffusion >>
rect 14 462 15 463 
<< pdiffusion >>
rect 15 462 16 463 
<< pdiffusion >>
rect 16 462 17 463 
<< pdiffusion >>
rect 17 462 18 463 
<< m1 >>
rect 19 462 20 463 
<< m1 >>
rect 21 462 22 463 
<< m1 >>
rect 28 462 29 463 
<< m1 >>
rect 30 462 31 463 
<< pdiffusion >>
rect 48 462 49 463 
<< pdiffusion >>
rect 49 462 50 463 
<< pdiffusion >>
rect 50 462 51 463 
<< pdiffusion >>
rect 51 462 52 463 
<< pdiffusion >>
rect 52 462 53 463 
<< pdiffusion >>
rect 53 462 54 463 
<< pdiffusion >>
rect 66 462 67 463 
<< pdiffusion >>
rect 67 462 68 463 
<< pdiffusion >>
rect 68 462 69 463 
<< pdiffusion >>
rect 69 462 70 463 
<< pdiffusion >>
rect 70 462 71 463 
<< pdiffusion >>
rect 71 462 72 463 
<< m1 >>
rect 73 462 74 463 
<< pdiffusion >>
rect 84 462 85 463 
<< pdiffusion >>
rect 85 462 86 463 
<< pdiffusion >>
rect 86 462 87 463 
<< pdiffusion >>
rect 87 462 88 463 
<< pdiffusion >>
rect 88 462 89 463 
<< pdiffusion >>
rect 89 462 90 463 
<< m1 >>
rect 100 462 101 463 
<< pdiffusion >>
rect 102 462 103 463 
<< m1 >>
rect 103 462 104 463 
<< pdiffusion >>
rect 103 462 104 463 
<< pdiffusion >>
rect 104 462 105 463 
<< pdiffusion >>
rect 105 462 106 463 
<< pdiffusion >>
rect 106 462 107 463 
<< pdiffusion >>
rect 107 462 108 463 
<< pdiffusion >>
rect 120 462 121 463 
<< pdiffusion >>
rect 121 462 122 463 
<< pdiffusion >>
rect 122 462 123 463 
<< pdiffusion >>
rect 123 462 124 463 
<< pdiffusion >>
rect 124 462 125 463 
<< pdiffusion >>
rect 125 462 126 463 
<< m1 >>
rect 136 462 137 463 
<< pdiffusion >>
rect 138 462 139 463 
<< m1 >>
rect 139 462 140 463 
<< pdiffusion >>
rect 139 462 140 463 
<< pdiffusion >>
rect 140 462 141 463 
<< pdiffusion >>
rect 141 462 142 463 
<< pdiffusion >>
rect 142 462 143 463 
<< pdiffusion >>
rect 143 462 144 463 
<< m1 >>
rect 152 462 153 463 
<< pdiffusion >>
rect 156 462 157 463 
<< pdiffusion >>
rect 157 462 158 463 
<< pdiffusion >>
rect 158 462 159 463 
<< pdiffusion >>
rect 159 462 160 463 
<< m1 >>
rect 160 462 161 463 
<< pdiffusion >>
rect 160 462 161 463 
<< pdiffusion >>
rect 161 462 162 463 
<< m1 >>
rect 163 462 164 463 
<< m1 >>
rect 172 462 173 463 
<< m2 >>
rect 172 462 173 463 
<< pdiffusion >>
rect 174 462 175 463 
<< pdiffusion >>
rect 175 462 176 463 
<< pdiffusion >>
rect 176 462 177 463 
<< pdiffusion >>
rect 177 462 178 463 
<< pdiffusion >>
rect 178 462 179 463 
<< pdiffusion >>
rect 179 462 180 463 
<< pdiffusion >>
rect 192 462 193 463 
<< pdiffusion >>
rect 193 462 194 463 
<< pdiffusion >>
rect 194 462 195 463 
<< pdiffusion >>
rect 195 462 196 463 
<< pdiffusion >>
rect 196 462 197 463 
<< pdiffusion >>
rect 197 462 198 463 
<< m1 >>
rect 199 462 200 463 
<< m1 >>
rect 208 462 209 463 
<< pdiffusion >>
rect 210 462 211 463 
<< pdiffusion >>
rect 211 462 212 463 
<< pdiffusion >>
rect 212 462 213 463 
<< pdiffusion >>
rect 213 462 214 463 
<< pdiffusion >>
rect 214 462 215 463 
<< pdiffusion >>
rect 215 462 216 463 
<< pdiffusion >>
rect 228 462 229 463 
<< m1 >>
rect 229 462 230 463 
<< pdiffusion >>
rect 229 462 230 463 
<< pdiffusion >>
rect 230 462 231 463 
<< pdiffusion >>
rect 231 462 232 463 
<< pdiffusion >>
rect 232 462 233 463 
<< pdiffusion >>
rect 233 462 234 463 
<< pdiffusion >>
rect 246 462 247 463 
<< pdiffusion >>
rect 247 462 248 463 
<< pdiffusion >>
rect 248 462 249 463 
<< pdiffusion >>
rect 249 462 250 463 
<< pdiffusion >>
rect 250 462 251 463 
<< pdiffusion >>
rect 251 462 252 463 
<< m1 >>
rect 253 462 254 463 
<< pdiffusion >>
rect 264 462 265 463 
<< pdiffusion >>
rect 265 462 266 463 
<< pdiffusion >>
rect 266 462 267 463 
<< pdiffusion >>
rect 267 462 268 463 
<< pdiffusion >>
rect 268 462 269 463 
<< pdiffusion >>
rect 269 462 270 463 
<< pdiffusion >>
rect 282 462 283 463 
<< pdiffusion >>
rect 283 462 284 463 
<< pdiffusion >>
rect 284 462 285 463 
<< pdiffusion >>
rect 285 462 286 463 
<< pdiffusion >>
rect 286 462 287 463 
<< pdiffusion >>
rect 287 462 288 463 
<< m1 >>
rect 289 462 290 463 
<< m1 >>
rect 298 462 299 463 
<< pdiffusion >>
rect 300 462 301 463 
<< pdiffusion >>
rect 301 462 302 463 
<< pdiffusion >>
rect 302 462 303 463 
<< pdiffusion >>
rect 303 462 304 463 
<< pdiffusion >>
rect 304 462 305 463 
<< pdiffusion >>
rect 305 462 306 463 
<< m1 >>
rect 307 462 308 463 
<< pdiffusion >>
rect 318 462 319 463 
<< pdiffusion >>
rect 319 462 320 463 
<< pdiffusion >>
rect 320 462 321 463 
<< pdiffusion >>
rect 321 462 322 463 
<< pdiffusion >>
rect 322 462 323 463 
<< pdiffusion >>
rect 323 462 324 463 
<< pdiffusion >>
rect 336 462 337 463 
<< pdiffusion >>
rect 337 462 338 463 
<< pdiffusion >>
rect 338 462 339 463 
<< pdiffusion >>
rect 339 462 340 463 
<< pdiffusion >>
rect 340 462 341 463 
<< pdiffusion >>
rect 341 462 342 463 
<< m1 >>
rect 352 462 353 463 
<< pdiffusion >>
rect 354 462 355 463 
<< pdiffusion >>
rect 355 462 356 463 
<< pdiffusion >>
rect 356 462 357 463 
<< pdiffusion >>
rect 357 462 358 463 
<< pdiffusion >>
rect 358 462 359 463 
<< pdiffusion >>
rect 359 462 360 463 
<< m1 >>
rect 361 462 362 463 
<< m2 >>
rect 362 462 363 463 
<< pdiffusion >>
rect 372 462 373 463 
<< pdiffusion >>
rect 373 462 374 463 
<< pdiffusion >>
rect 374 462 375 463 
<< pdiffusion >>
rect 375 462 376 463 
<< pdiffusion >>
rect 376 462 377 463 
<< pdiffusion >>
rect 377 462 378 463 
<< m1 >>
rect 381 462 382 463 
<< pdiffusion >>
rect 390 462 391 463 
<< pdiffusion >>
rect 391 462 392 463 
<< pdiffusion >>
rect 392 462 393 463 
<< pdiffusion >>
rect 393 462 394 463 
<< m1 >>
rect 394 462 395 463 
<< pdiffusion >>
rect 394 462 395 463 
<< pdiffusion >>
rect 395 462 396 463 
<< m1 >>
rect 402 462 403 463 
<< pdiffusion >>
rect 408 462 409 463 
<< m1 >>
rect 409 462 410 463 
<< pdiffusion >>
rect 409 462 410 463 
<< pdiffusion >>
rect 410 462 411 463 
<< pdiffusion >>
rect 411 462 412 463 
<< pdiffusion >>
rect 412 462 413 463 
<< pdiffusion >>
rect 413 462 414 463 
<< pdiffusion >>
rect 426 462 427 463 
<< pdiffusion >>
rect 427 462 428 463 
<< pdiffusion >>
rect 428 462 429 463 
<< pdiffusion >>
rect 429 462 430 463 
<< pdiffusion >>
rect 430 462 431 463 
<< pdiffusion >>
rect 431 462 432 463 
<< m1 >>
rect 433 462 434 463 
<< pdiffusion >>
rect 444 462 445 463 
<< pdiffusion >>
rect 445 462 446 463 
<< pdiffusion >>
rect 446 462 447 463 
<< pdiffusion >>
rect 447 462 448 463 
<< m1 >>
rect 448 462 449 463 
<< pdiffusion >>
rect 448 462 449 463 
<< pdiffusion >>
rect 449 462 450 463 
<< m1 >>
rect 451 462 452 463 
<< m2 >>
rect 451 462 452 463 
<< pdiffusion >>
rect 462 462 463 463 
<< pdiffusion >>
rect 463 462 464 463 
<< pdiffusion >>
rect 464 462 465 463 
<< pdiffusion >>
rect 465 462 466 463 
<< pdiffusion >>
rect 466 462 467 463 
<< pdiffusion >>
rect 467 462 468 463 
<< m1 >>
rect 472 462 473 463 
<< pdiffusion >>
rect 480 462 481 463 
<< pdiffusion >>
rect 481 462 482 463 
<< pdiffusion >>
rect 482 462 483 463 
<< pdiffusion >>
rect 483 462 484 463 
<< pdiffusion >>
rect 484 462 485 463 
<< pdiffusion >>
rect 485 462 486 463 
<< m1 >>
rect 487 462 488 463 
<< m1 >>
rect 489 462 490 463 
<< pdiffusion >>
rect 498 462 499 463 
<< pdiffusion >>
rect 499 462 500 463 
<< pdiffusion >>
rect 500 462 501 463 
<< pdiffusion >>
rect 501 462 502 463 
<< pdiffusion >>
rect 502 462 503 463 
<< pdiffusion >>
rect 503 462 504 463 
<< pdiffusion >>
rect 516 462 517 463 
<< pdiffusion >>
rect 517 462 518 463 
<< pdiffusion >>
rect 518 462 519 463 
<< pdiffusion >>
rect 519 462 520 463 
<< pdiffusion >>
rect 520 462 521 463 
<< pdiffusion >>
rect 521 462 522 463 
<< pdiffusion >>
rect 12 463 13 464 
<< pdiffusion >>
rect 13 463 14 464 
<< pdiffusion >>
rect 14 463 15 464 
<< pdiffusion >>
rect 15 463 16 464 
<< pdiffusion >>
rect 16 463 17 464 
<< pdiffusion >>
rect 17 463 18 464 
<< m1 >>
rect 19 463 20 464 
<< m1 >>
rect 21 463 22 464 
<< m1 >>
rect 28 463 29 464 
<< m1 >>
rect 30 463 31 464 
<< pdiffusion >>
rect 48 463 49 464 
<< pdiffusion >>
rect 49 463 50 464 
<< pdiffusion >>
rect 50 463 51 464 
<< pdiffusion >>
rect 51 463 52 464 
<< pdiffusion >>
rect 52 463 53 464 
<< pdiffusion >>
rect 53 463 54 464 
<< pdiffusion >>
rect 66 463 67 464 
<< pdiffusion >>
rect 67 463 68 464 
<< pdiffusion >>
rect 68 463 69 464 
<< pdiffusion >>
rect 69 463 70 464 
<< pdiffusion >>
rect 70 463 71 464 
<< pdiffusion >>
rect 71 463 72 464 
<< m1 >>
rect 73 463 74 464 
<< pdiffusion >>
rect 84 463 85 464 
<< pdiffusion >>
rect 85 463 86 464 
<< pdiffusion >>
rect 86 463 87 464 
<< pdiffusion >>
rect 87 463 88 464 
<< pdiffusion >>
rect 88 463 89 464 
<< pdiffusion >>
rect 89 463 90 464 
<< m1 >>
rect 100 463 101 464 
<< pdiffusion >>
rect 102 463 103 464 
<< pdiffusion >>
rect 103 463 104 464 
<< pdiffusion >>
rect 104 463 105 464 
<< pdiffusion >>
rect 105 463 106 464 
<< pdiffusion >>
rect 106 463 107 464 
<< pdiffusion >>
rect 107 463 108 464 
<< pdiffusion >>
rect 120 463 121 464 
<< pdiffusion >>
rect 121 463 122 464 
<< pdiffusion >>
rect 122 463 123 464 
<< pdiffusion >>
rect 123 463 124 464 
<< pdiffusion >>
rect 124 463 125 464 
<< pdiffusion >>
rect 125 463 126 464 
<< m1 >>
rect 136 463 137 464 
<< pdiffusion >>
rect 138 463 139 464 
<< pdiffusion >>
rect 139 463 140 464 
<< pdiffusion >>
rect 140 463 141 464 
<< pdiffusion >>
rect 141 463 142 464 
<< pdiffusion >>
rect 142 463 143 464 
<< pdiffusion >>
rect 143 463 144 464 
<< m1 >>
rect 152 463 153 464 
<< pdiffusion >>
rect 156 463 157 464 
<< pdiffusion >>
rect 157 463 158 464 
<< pdiffusion >>
rect 158 463 159 464 
<< pdiffusion >>
rect 159 463 160 464 
<< pdiffusion >>
rect 160 463 161 464 
<< pdiffusion >>
rect 161 463 162 464 
<< m1 >>
rect 163 463 164 464 
<< m1 >>
rect 172 463 173 464 
<< m2 >>
rect 172 463 173 464 
<< pdiffusion >>
rect 174 463 175 464 
<< pdiffusion >>
rect 175 463 176 464 
<< pdiffusion >>
rect 176 463 177 464 
<< pdiffusion >>
rect 177 463 178 464 
<< pdiffusion >>
rect 178 463 179 464 
<< pdiffusion >>
rect 179 463 180 464 
<< pdiffusion >>
rect 192 463 193 464 
<< pdiffusion >>
rect 193 463 194 464 
<< pdiffusion >>
rect 194 463 195 464 
<< pdiffusion >>
rect 195 463 196 464 
<< pdiffusion >>
rect 196 463 197 464 
<< pdiffusion >>
rect 197 463 198 464 
<< m1 >>
rect 199 463 200 464 
<< m1 >>
rect 208 463 209 464 
<< pdiffusion >>
rect 210 463 211 464 
<< pdiffusion >>
rect 211 463 212 464 
<< pdiffusion >>
rect 212 463 213 464 
<< pdiffusion >>
rect 213 463 214 464 
<< pdiffusion >>
rect 214 463 215 464 
<< pdiffusion >>
rect 215 463 216 464 
<< pdiffusion >>
rect 228 463 229 464 
<< pdiffusion >>
rect 229 463 230 464 
<< pdiffusion >>
rect 230 463 231 464 
<< pdiffusion >>
rect 231 463 232 464 
<< pdiffusion >>
rect 232 463 233 464 
<< pdiffusion >>
rect 233 463 234 464 
<< pdiffusion >>
rect 246 463 247 464 
<< pdiffusion >>
rect 247 463 248 464 
<< pdiffusion >>
rect 248 463 249 464 
<< pdiffusion >>
rect 249 463 250 464 
<< pdiffusion >>
rect 250 463 251 464 
<< pdiffusion >>
rect 251 463 252 464 
<< m1 >>
rect 253 463 254 464 
<< pdiffusion >>
rect 264 463 265 464 
<< pdiffusion >>
rect 265 463 266 464 
<< pdiffusion >>
rect 266 463 267 464 
<< pdiffusion >>
rect 267 463 268 464 
<< pdiffusion >>
rect 268 463 269 464 
<< pdiffusion >>
rect 269 463 270 464 
<< pdiffusion >>
rect 282 463 283 464 
<< pdiffusion >>
rect 283 463 284 464 
<< pdiffusion >>
rect 284 463 285 464 
<< pdiffusion >>
rect 285 463 286 464 
<< pdiffusion >>
rect 286 463 287 464 
<< pdiffusion >>
rect 287 463 288 464 
<< m1 >>
rect 289 463 290 464 
<< m1 >>
rect 298 463 299 464 
<< pdiffusion >>
rect 300 463 301 464 
<< pdiffusion >>
rect 301 463 302 464 
<< pdiffusion >>
rect 302 463 303 464 
<< pdiffusion >>
rect 303 463 304 464 
<< pdiffusion >>
rect 304 463 305 464 
<< pdiffusion >>
rect 305 463 306 464 
<< m1 >>
rect 307 463 308 464 
<< pdiffusion >>
rect 318 463 319 464 
<< pdiffusion >>
rect 319 463 320 464 
<< pdiffusion >>
rect 320 463 321 464 
<< pdiffusion >>
rect 321 463 322 464 
<< pdiffusion >>
rect 322 463 323 464 
<< pdiffusion >>
rect 323 463 324 464 
<< pdiffusion >>
rect 336 463 337 464 
<< pdiffusion >>
rect 337 463 338 464 
<< pdiffusion >>
rect 338 463 339 464 
<< pdiffusion >>
rect 339 463 340 464 
<< pdiffusion >>
rect 340 463 341 464 
<< pdiffusion >>
rect 341 463 342 464 
<< m1 >>
rect 352 463 353 464 
<< pdiffusion >>
rect 354 463 355 464 
<< pdiffusion >>
rect 355 463 356 464 
<< pdiffusion >>
rect 356 463 357 464 
<< pdiffusion >>
rect 357 463 358 464 
<< pdiffusion >>
rect 358 463 359 464 
<< pdiffusion >>
rect 359 463 360 464 
<< m1 >>
rect 361 463 362 464 
<< m2 >>
rect 362 463 363 464 
<< pdiffusion >>
rect 372 463 373 464 
<< pdiffusion >>
rect 373 463 374 464 
<< pdiffusion >>
rect 374 463 375 464 
<< pdiffusion >>
rect 375 463 376 464 
<< pdiffusion >>
rect 376 463 377 464 
<< pdiffusion >>
rect 377 463 378 464 
<< m1 >>
rect 381 463 382 464 
<< pdiffusion >>
rect 390 463 391 464 
<< pdiffusion >>
rect 391 463 392 464 
<< pdiffusion >>
rect 392 463 393 464 
<< pdiffusion >>
rect 393 463 394 464 
<< pdiffusion >>
rect 394 463 395 464 
<< pdiffusion >>
rect 395 463 396 464 
<< m1 >>
rect 402 463 403 464 
<< pdiffusion >>
rect 408 463 409 464 
<< pdiffusion >>
rect 409 463 410 464 
<< pdiffusion >>
rect 410 463 411 464 
<< pdiffusion >>
rect 411 463 412 464 
<< pdiffusion >>
rect 412 463 413 464 
<< pdiffusion >>
rect 413 463 414 464 
<< pdiffusion >>
rect 426 463 427 464 
<< pdiffusion >>
rect 427 463 428 464 
<< pdiffusion >>
rect 428 463 429 464 
<< pdiffusion >>
rect 429 463 430 464 
<< pdiffusion >>
rect 430 463 431 464 
<< pdiffusion >>
rect 431 463 432 464 
<< m1 >>
rect 433 463 434 464 
<< pdiffusion >>
rect 444 463 445 464 
<< pdiffusion >>
rect 445 463 446 464 
<< pdiffusion >>
rect 446 463 447 464 
<< pdiffusion >>
rect 447 463 448 464 
<< pdiffusion >>
rect 448 463 449 464 
<< pdiffusion >>
rect 449 463 450 464 
<< m1 >>
rect 451 463 452 464 
<< m2 >>
rect 451 463 452 464 
<< pdiffusion >>
rect 462 463 463 464 
<< pdiffusion >>
rect 463 463 464 464 
<< pdiffusion >>
rect 464 463 465 464 
<< pdiffusion >>
rect 465 463 466 464 
<< pdiffusion >>
rect 466 463 467 464 
<< pdiffusion >>
rect 467 463 468 464 
<< m1 >>
rect 472 463 473 464 
<< pdiffusion >>
rect 480 463 481 464 
<< pdiffusion >>
rect 481 463 482 464 
<< pdiffusion >>
rect 482 463 483 464 
<< pdiffusion >>
rect 483 463 484 464 
<< pdiffusion >>
rect 484 463 485 464 
<< pdiffusion >>
rect 485 463 486 464 
<< m1 >>
rect 487 463 488 464 
<< m1 >>
rect 489 463 490 464 
<< pdiffusion >>
rect 498 463 499 464 
<< pdiffusion >>
rect 499 463 500 464 
<< pdiffusion >>
rect 500 463 501 464 
<< pdiffusion >>
rect 501 463 502 464 
<< pdiffusion >>
rect 502 463 503 464 
<< pdiffusion >>
rect 503 463 504 464 
<< pdiffusion >>
rect 516 463 517 464 
<< pdiffusion >>
rect 517 463 518 464 
<< pdiffusion >>
rect 518 463 519 464 
<< pdiffusion >>
rect 519 463 520 464 
<< pdiffusion >>
rect 520 463 521 464 
<< pdiffusion >>
rect 521 463 522 464 
<< pdiffusion >>
rect 12 464 13 465 
<< pdiffusion >>
rect 13 464 14 465 
<< pdiffusion >>
rect 14 464 15 465 
<< pdiffusion >>
rect 15 464 16 465 
<< pdiffusion >>
rect 16 464 17 465 
<< pdiffusion >>
rect 17 464 18 465 
<< m1 >>
rect 19 464 20 465 
<< m1 >>
rect 21 464 22 465 
<< m1 >>
rect 28 464 29 465 
<< m1 >>
rect 30 464 31 465 
<< pdiffusion >>
rect 48 464 49 465 
<< pdiffusion >>
rect 49 464 50 465 
<< pdiffusion >>
rect 50 464 51 465 
<< pdiffusion >>
rect 51 464 52 465 
<< pdiffusion >>
rect 52 464 53 465 
<< pdiffusion >>
rect 53 464 54 465 
<< pdiffusion >>
rect 66 464 67 465 
<< pdiffusion >>
rect 67 464 68 465 
<< pdiffusion >>
rect 68 464 69 465 
<< pdiffusion >>
rect 69 464 70 465 
<< pdiffusion >>
rect 70 464 71 465 
<< pdiffusion >>
rect 71 464 72 465 
<< m1 >>
rect 73 464 74 465 
<< pdiffusion >>
rect 84 464 85 465 
<< pdiffusion >>
rect 85 464 86 465 
<< pdiffusion >>
rect 86 464 87 465 
<< pdiffusion >>
rect 87 464 88 465 
<< pdiffusion >>
rect 88 464 89 465 
<< pdiffusion >>
rect 89 464 90 465 
<< m1 >>
rect 100 464 101 465 
<< pdiffusion >>
rect 102 464 103 465 
<< pdiffusion >>
rect 103 464 104 465 
<< pdiffusion >>
rect 104 464 105 465 
<< pdiffusion >>
rect 105 464 106 465 
<< pdiffusion >>
rect 106 464 107 465 
<< pdiffusion >>
rect 107 464 108 465 
<< pdiffusion >>
rect 120 464 121 465 
<< pdiffusion >>
rect 121 464 122 465 
<< pdiffusion >>
rect 122 464 123 465 
<< pdiffusion >>
rect 123 464 124 465 
<< pdiffusion >>
rect 124 464 125 465 
<< pdiffusion >>
rect 125 464 126 465 
<< m1 >>
rect 136 464 137 465 
<< pdiffusion >>
rect 138 464 139 465 
<< pdiffusion >>
rect 139 464 140 465 
<< pdiffusion >>
rect 140 464 141 465 
<< pdiffusion >>
rect 141 464 142 465 
<< pdiffusion >>
rect 142 464 143 465 
<< pdiffusion >>
rect 143 464 144 465 
<< m1 >>
rect 152 464 153 465 
<< pdiffusion >>
rect 156 464 157 465 
<< pdiffusion >>
rect 157 464 158 465 
<< pdiffusion >>
rect 158 464 159 465 
<< pdiffusion >>
rect 159 464 160 465 
<< pdiffusion >>
rect 160 464 161 465 
<< pdiffusion >>
rect 161 464 162 465 
<< m1 >>
rect 163 464 164 465 
<< m1 >>
rect 172 464 173 465 
<< m2 >>
rect 172 464 173 465 
<< pdiffusion >>
rect 174 464 175 465 
<< pdiffusion >>
rect 175 464 176 465 
<< pdiffusion >>
rect 176 464 177 465 
<< pdiffusion >>
rect 177 464 178 465 
<< pdiffusion >>
rect 178 464 179 465 
<< pdiffusion >>
rect 179 464 180 465 
<< pdiffusion >>
rect 192 464 193 465 
<< pdiffusion >>
rect 193 464 194 465 
<< pdiffusion >>
rect 194 464 195 465 
<< pdiffusion >>
rect 195 464 196 465 
<< pdiffusion >>
rect 196 464 197 465 
<< pdiffusion >>
rect 197 464 198 465 
<< m1 >>
rect 199 464 200 465 
<< m1 >>
rect 208 464 209 465 
<< pdiffusion >>
rect 210 464 211 465 
<< pdiffusion >>
rect 211 464 212 465 
<< pdiffusion >>
rect 212 464 213 465 
<< pdiffusion >>
rect 213 464 214 465 
<< pdiffusion >>
rect 214 464 215 465 
<< pdiffusion >>
rect 215 464 216 465 
<< pdiffusion >>
rect 228 464 229 465 
<< pdiffusion >>
rect 229 464 230 465 
<< pdiffusion >>
rect 230 464 231 465 
<< pdiffusion >>
rect 231 464 232 465 
<< pdiffusion >>
rect 232 464 233 465 
<< pdiffusion >>
rect 233 464 234 465 
<< pdiffusion >>
rect 246 464 247 465 
<< pdiffusion >>
rect 247 464 248 465 
<< pdiffusion >>
rect 248 464 249 465 
<< pdiffusion >>
rect 249 464 250 465 
<< pdiffusion >>
rect 250 464 251 465 
<< pdiffusion >>
rect 251 464 252 465 
<< m1 >>
rect 253 464 254 465 
<< pdiffusion >>
rect 264 464 265 465 
<< pdiffusion >>
rect 265 464 266 465 
<< pdiffusion >>
rect 266 464 267 465 
<< pdiffusion >>
rect 267 464 268 465 
<< pdiffusion >>
rect 268 464 269 465 
<< pdiffusion >>
rect 269 464 270 465 
<< pdiffusion >>
rect 282 464 283 465 
<< pdiffusion >>
rect 283 464 284 465 
<< pdiffusion >>
rect 284 464 285 465 
<< pdiffusion >>
rect 285 464 286 465 
<< pdiffusion >>
rect 286 464 287 465 
<< pdiffusion >>
rect 287 464 288 465 
<< m1 >>
rect 289 464 290 465 
<< m1 >>
rect 298 464 299 465 
<< pdiffusion >>
rect 300 464 301 465 
<< pdiffusion >>
rect 301 464 302 465 
<< pdiffusion >>
rect 302 464 303 465 
<< pdiffusion >>
rect 303 464 304 465 
<< pdiffusion >>
rect 304 464 305 465 
<< pdiffusion >>
rect 305 464 306 465 
<< m1 >>
rect 307 464 308 465 
<< pdiffusion >>
rect 318 464 319 465 
<< pdiffusion >>
rect 319 464 320 465 
<< pdiffusion >>
rect 320 464 321 465 
<< pdiffusion >>
rect 321 464 322 465 
<< pdiffusion >>
rect 322 464 323 465 
<< pdiffusion >>
rect 323 464 324 465 
<< pdiffusion >>
rect 336 464 337 465 
<< pdiffusion >>
rect 337 464 338 465 
<< pdiffusion >>
rect 338 464 339 465 
<< pdiffusion >>
rect 339 464 340 465 
<< pdiffusion >>
rect 340 464 341 465 
<< pdiffusion >>
rect 341 464 342 465 
<< m1 >>
rect 352 464 353 465 
<< pdiffusion >>
rect 354 464 355 465 
<< pdiffusion >>
rect 355 464 356 465 
<< pdiffusion >>
rect 356 464 357 465 
<< pdiffusion >>
rect 357 464 358 465 
<< pdiffusion >>
rect 358 464 359 465 
<< pdiffusion >>
rect 359 464 360 465 
<< m1 >>
rect 361 464 362 465 
<< m2 >>
rect 362 464 363 465 
<< pdiffusion >>
rect 372 464 373 465 
<< pdiffusion >>
rect 373 464 374 465 
<< pdiffusion >>
rect 374 464 375 465 
<< pdiffusion >>
rect 375 464 376 465 
<< pdiffusion >>
rect 376 464 377 465 
<< pdiffusion >>
rect 377 464 378 465 
<< m1 >>
rect 381 464 382 465 
<< pdiffusion >>
rect 390 464 391 465 
<< pdiffusion >>
rect 391 464 392 465 
<< pdiffusion >>
rect 392 464 393 465 
<< pdiffusion >>
rect 393 464 394 465 
<< pdiffusion >>
rect 394 464 395 465 
<< pdiffusion >>
rect 395 464 396 465 
<< m1 >>
rect 402 464 403 465 
<< pdiffusion >>
rect 408 464 409 465 
<< pdiffusion >>
rect 409 464 410 465 
<< pdiffusion >>
rect 410 464 411 465 
<< pdiffusion >>
rect 411 464 412 465 
<< pdiffusion >>
rect 412 464 413 465 
<< pdiffusion >>
rect 413 464 414 465 
<< pdiffusion >>
rect 426 464 427 465 
<< pdiffusion >>
rect 427 464 428 465 
<< pdiffusion >>
rect 428 464 429 465 
<< pdiffusion >>
rect 429 464 430 465 
<< pdiffusion >>
rect 430 464 431 465 
<< pdiffusion >>
rect 431 464 432 465 
<< m1 >>
rect 433 464 434 465 
<< pdiffusion >>
rect 444 464 445 465 
<< pdiffusion >>
rect 445 464 446 465 
<< pdiffusion >>
rect 446 464 447 465 
<< pdiffusion >>
rect 447 464 448 465 
<< pdiffusion >>
rect 448 464 449 465 
<< pdiffusion >>
rect 449 464 450 465 
<< m1 >>
rect 451 464 452 465 
<< m2 >>
rect 451 464 452 465 
<< pdiffusion >>
rect 462 464 463 465 
<< pdiffusion >>
rect 463 464 464 465 
<< pdiffusion >>
rect 464 464 465 465 
<< pdiffusion >>
rect 465 464 466 465 
<< pdiffusion >>
rect 466 464 467 465 
<< pdiffusion >>
rect 467 464 468 465 
<< m1 >>
rect 472 464 473 465 
<< pdiffusion >>
rect 480 464 481 465 
<< pdiffusion >>
rect 481 464 482 465 
<< pdiffusion >>
rect 482 464 483 465 
<< pdiffusion >>
rect 483 464 484 465 
<< pdiffusion >>
rect 484 464 485 465 
<< pdiffusion >>
rect 485 464 486 465 
<< m1 >>
rect 487 464 488 465 
<< m1 >>
rect 489 464 490 465 
<< pdiffusion >>
rect 498 464 499 465 
<< pdiffusion >>
rect 499 464 500 465 
<< pdiffusion >>
rect 500 464 501 465 
<< pdiffusion >>
rect 501 464 502 465 
<< pdiffusion >>
rect 502 464 503 465 
<< pdiffusion >>
rect 503 464 504 465 
<< pdiffusion >>
rect 516 464 517 465 
<< pdiffusion >>
rect 517 464 518 465 
<< pdiffusion >>
rect 518 464 519 465 
<< pdiffusion >>
rect 519 464 520 465 
<< pdiffusion >>
rect 520 464 521 465 
<< pdiffusion >>
rect 521 464 522 465 
<< pdiffusion >>
rect 12 465 13 466 
<< pdiffusion >>
rect 13 465 14 466 
<< pdiffusion >>
rect 14 465 15 466 
<< pdiffusion >>
rect 15 465 16 466 
<< pdiffusion >>
rect 16 465 17 466 
<< pdiffusion >>
rect 17 465 18 466 
<< m1 >>
rect 19 465 20 466 
<< m1 >>
rect 21 465 22 466 
<< m1 >>
rect 28 465 29 466 
<< m1 >>
rect 30 465 31 466 
<< pdiffusion >>
rect 48 465 49 466 
<< pdiffusion >>
rect 49 465 50 466 
<< pdiffusion >>
rect 50 465 51 466 
<< pdiffusion >>
rect 51 465 52 466 
<< pdiffusion >>
rect 52 465 53 466 
<< pdiffusion >>
rect 53 465 54 466 
<< pdiffusion >>
rect 66 465 67 466 
<< pdiffusion >>
rect 67 465 68 466 
<< pdiffusion >>
rect 68 465 69 466 
<< pdiffusion >>
rect 69 465 70 466 
<< pdiffusion >>
rect 70 465 71 466 
<< pdiffusion >>
rect 71 465 72 466 
<< m1 >>
rect 73 465 74 466 
<< pdiffusion >>
rect 84 465 85 466 
<< pdiffusion >>
rect 85 465 86 466 
<< pdiffusion >>
rect 86 465 87 466 
<< pdiffusion >>
rect 87 465 88 466 
<< pdiffusion >>
rect 88 465 89 466 
<< pdiffusion >>
rect 89 465 90 466 
<< m1 >>
rect 100 465 101 466 
<< pdiffusion >>
rect 102 465 103 466 
<< pdiffusion >>
rect 103 465 104 466 
<< pdiffusion >>
rect 104 465 105 466 
<< pdiffusion >>
rect 105 465 106 466 
<< pdiffusion >>
rect 106 465 107 466 
<< pdiffusion >>
rect 107 465 108 466 
<< pdiffusion >>
rect 120 465 121 466 
<< pdiffusion >>
rect 121 465 122 466 
<< pdiffusion >>
rect 122 465 123 466 
<< pdiffusion >>
rect 123 465 124 466 
<< pdiffusion >>
rect 124 465 125 466 
<< pdiffusion >>
rect 125 465 126 466 
<< m1 >>
rect 136 465 137 466 
<< pdiffusion >>
rect 138 465 139 466 
<< pdiffusion >>
rect 139 465 140 466 
<< pdiffusion >>
rect 140 465 141 466 
<< pdiffusion >>
rect 141 465 142 466 
<< pdiffusion >>
rect 142 465 143 466 
<< pdiffusion >>
rect 143 465 144 466 
<< m1 >>
rect 152 465 153 466 
<< pdiffusion >>
rect 156 465 157 466 
<< pdiffusion >>
rect 157 465 158 466 
<< pdiffusion >>
rect 158 465 159 466 
<< pdiffusion >>
rect 159 465 160 466 
<< pdiffusion >>
rect 160 465 161 466 
<< pdiffusion >>
rect 161 465 162 466 
<< m1 >>
rect 163 465 164 466 
<< m1 >>
rect 172 465 173 466 
<< m2 >>
rect 172 465 173 466 
<< pdiffusion >>
rect 174 465 175 466 
<< pdiffusion >>
rect 175 465 176 466 
<< pdiffusion >>
rect 176 465 177 466 
<< pdiffusion >>
rect 177 465 178 466 
<< pdiffusion >>
rect 178 465 179 466 
<< pdiffusion >>
rect 179 465 180 466 
<< pdiffusion >>
rect 192 465 193 466 
<< pdiffusion >>
rect 193 465 194 466 
<< pdiffusion >>
rect 194 465 195 466 
<< pdiffusion >>
rect 195 465 196 466 
<< pdiffusion >>
rect 196 465 197 466 
<< pdiffusion >>
rect 197 465 198 466 
<< m1 >>
rect 199 465 200 466 
<< m1 >>
rect 208 465 209 466 
<< pdiffusion >>
rect 210 465 211 466 
<< pdiffusion >>
rect 211 465 212 466 
<< pdiffusion >>
rect 212 465 213 466 
<< pdiffusion >>
rect 213 465 214 466 
<< pdiffusion >>
rect 214 465 215 466 
<< pdiffusion >>
rect 215 465 216 466 
<< pdiffusion >>
rect 228 465 229 466 
<< pdiffusion >>
rect 229 465 230 466 
<< pdiffusion >>
rect 230 465 231 466 
<< pdiffusion >>
rect 231 465 232 466 
<< pdiffusion >>
rect 232 465 233 466 
<< pdiffusion >>
rect 233 465 234 466 
<< pdiffusion >>
rect 246 465 247 466 
<< pdiffusion >>
rect 247 465 248 466 
<< pdiffusion >>
rect 248 465 249 466 
<< pdiffusion >>
rect 249 465 250 466 
<< pdiffusion >>
rect 250 465 251 466 
<< pdiffusion >>
rect 251 465 252 466 
<< m1 >>
rect 253 465 254 466 
<< pdiffusion >>
rect 264 465 265 466 
<< pdiffusion >>
rect 265 465 266 466 
<< pdiffusion >>
rect 266 465 267 466 
<< pdiffusion >>
rect 267 465 268 466 
<< pdiffusion >>
rect 268 465 269 466 
<< pdiffusion >>
rect 269 465 270 466 
<< pdiffusion >>
rect 282 465 283 466 
<< pdiffusion >>
rect 283 465 284 466 
<< pdiffusion >>
rect 284 465 285 466 
<< pdiffusion >>
rect 285 465 286 466 
<< pdiffusion >>
rect 286 465 287 466 
<< pdiffusion >>
rect 287 465 288 466 
<< m1 >>
rect 289 465 290 466 
<< m1 >>
rect 298 465 299 466 
<< pdiffusion >>
rect 300 465 301 466 
<< pdiffusion >>
rect 301 465 302 466 
<< pdiffusion >>
rect 302 465 303 466 
<< pdiffusion >>
rect 303 465 304 466 
<< pdiffusion >>
rect 304 465 305 466 
<< pdiffusion >>
rect 305 465 306 466 
<< m1 >>
rect 307 465 308 466 
<< pdiffusion >>
rect 318 465 319 466 
<< pdiffusion >>
rect 319 465 320 466 
<< pdiffusion >>
rect 320 465 321 466 
<< pdiffusion >>
rect 321 465 322 466 
<< pdiffusion >>
rect 322 465 323 466 
<< pdiffusion >>
rect 323 465 324 466 
<< pdiffusion >>
rect 336 465 337 466 
<< pdiffusion >>
rect 337 465 338 466 
<< pdiffusion >>
rect 338 465 339 466 
<< pdiffusion >>
rect 339 465 340 466 
<< pdiffusion >>
rect 340 465 341 466 
<< pdiffusion >>
rect 341 465 342 466 
<< m1 >>
rect 352 465 353 466 
<< pdiffusion >>
rect 354 465 355 466 
<< pdiffusion >>
rect 355 465 356 466 
<< pdiffusion >>
rect 356 465 357 466 
<< pdiffusion >>
rect 357 465 358 466 
<< pdiffusion >>
rect 358 465 359 466 
<< pdiffusion >>
rect 359 465 360 466 
<< m1 >>
rect 361 465 362 466 
<< m2 >>
rect 362 465 363 466 
<< pdiffusion >>
rect 372 465 373 466 
<< pdiffusion >>
rect 373 465 374 466 
<< pdiffusion >>
rect 374 465 375 466 
<< pdiffusion >>
rect 375 465 376 466 
<< pdiffusion >>
rect 376 465 377 466 
<< pdiffusion >>
rect 377 465 378 466 
<< m1 >>
rect 381 465 382 466 
<< pdiffusion >>
rect 390 465 391 466 
<< pdiffusion >>
rect 391 465 392 466 
<< pdiffusion >>
rect 392 465 393 466 
<< pdiffusion >>
rect 393 465 394 466 
<< pdiffusion >>
rect 394 465 395 466 
<< pdiffusion >>
rect 395 465 396 466 
<< m1 >>
rect 402 465 403 466 
<< pdiffusion >>
rect 408 465 409 466 
<< pdiffusion >>
rect 409 465 410 466 
<< pdiffusion >>
rect 410 465 411 466 
<< pdiffusion >>
rect 411 465 412 466 
<< pdiffusion >>
rect 412 465 413 466 
<< pdiffusion >>
rect 413 465 414 466 
<< pdiffusion >>
rect 426 465 427 466 
<< pdiffusion >>
rect 427 465 428 466 
<< pdiffusion >>
rect 428 465 429 466 
<< pdiffusion >>
rect 429 465 430 466 
<< pdiffusion >>
rect 430 465 431 466 
<< pdiffusion >>
rect 431 465 432 466 
<< m1 >>
rect 433 465 434 466 
<< pdiffusion >>
rect 444 465 445 466 
<< pdiffusion >>
rect 445 465 446 466 
<< pdiffusion >>
rect 446 465 447 466 
<< pdiffusion >>
rect 447 465 448 466 
<< pdiffusion >>
rect 448 465 449 466 
<< pdiffusion >>
rect 449 465 450 466 
<< m1 >>
rect 451 465 452 466 
<< m2 >>
rect 451 465 452 466 
<< pdiffusion >>
rect 462 465 463 466 
<< pdiffusion >>
rect 463 465 464 466 
<< pdiffusion >>
rect 464 465 465 466 
<< pdiffusion >>
rect 465 465 466 466 
<< pdiffusion >>
rect 466 465 467 466 
<< pdiffusion >>
rect 467 465 468 466 
<< m1 >>
rect 472 465 473 466 
<< pdiffusion >>
rect 480 465 481 466 
<< pdiffusion >>
rect 481 465 482 466 
<< pdiffusion >>
rect 482 465 483 466 
<< pdiffusion >>
rect 483 465 484 466 
<< pdiffusion >>
rect 484 465 485 466 
<< pdiffusion >>
rect 485 465 486 466 
<< m1 >>
rect 487 465 488 466 
<< m1 >>
rect 489 465 490 466 
<< pdiffusion >>
rect 498 465 499 466 
<< pdiffusion >>
rect 499 465 500 466 
<< pdiffusion >>
rect 500 465 501 466 
<< pdiffusion >>
rect 501 465 502 466 
<< pdiffusion >>
rect 502 465 503 466 
<< pdiffusion >>
rect 503 465 504 466 
<< pdiffusion >>
rect 516 465 517 466 
<< pdiffusion >>
rect 517 465 518 466 
<< pdiffusion >>
rect 518 465 519 466 
<< pdiffusion >>
rect 519 465 520 466 
<< pdiffusion >>
rect 520 465 521 466 
<< pdiffusion >>
rect 521 465 522 466 
<< pdiffusion >>
rect 12 466 13 467 
<< pdiffusion >>
rect 13 466 14 467 
<< pdiffusion >>
rect 14 466 15 467 
<< pdiffusion >>
rect 15 466 16 467 
<< pdiffusion >>
rect 16 466 17 467 
<< pdiffusion >>
rect 17 466 18 467 
<< m1 >>
rect 19 466 20 467 
<< m1 >>
rect 21 466 22 467 
<< m1 >>
rect 28 466 29 467 
<< m1 >>
rect 30 466 31 467 
<< pdiffusion >>
rect 48 466 49 467 
<< pdiffusion >>
rect 49 466 50 467 
<< pdiffusion >>
rect 50 466 51 467 
<< pdiffusion >>
rect 51 466 52 467 
<< pdiffusion >>
rect 52 466 53 467 
<< pdiffusion >>
rect 53 466 54 467 
<< pdiffusion >>
rect 66 466 67 467 
<< pdiffusion >>
rect 67 466 68 467 
<< pdiffusion >>
rect 68 466 69 467 
<< pdiffusion >>
rect 69 466 70 467 
<< pdiffusion >>
rect 70 466 71 467 
<< pdiffusion >>
rect 71 466 72 467 
<< m1 >>
rect 73 466 74 467 
<< pdiffusion >>
rect 84 466 85 467 
<< pdiffusion >>
rect 85 466 86 467 
<< pdiffusion >>
rect 86 466 87 467 
<< pdiffusion >>
rect 87 466 88 467 
<< pdiffusion >>
rect 88 466 89 467 
<< pdiffusion >>
rect 89 466 90 467 
<< m1 >>
rect 100 466 101 467 
<< pdiffusion >>
rect 102 466 103 467 
<< pdiffusion >>
rect 103 466 104 467 
<< pdiffusion >>
rect 104 466 105 467 
<< pdiffusion >>
rect 105 466 106 467 
<< pdiffusion >>
rect 106 466 107 467 
<< pdiffusion >>
rect 107 466 108 467 
<< pdiffusion >>
rect 120 466 121 467 
<< pdiffusion >>
rect 121 466 122 467 
<< pdiffusion >>
rect 122 466 123 467 
<< pdiffusion >>
rect 123 466 124 467 
<< pdiffusion >>
rect 124 466 125 467 
<< pdiffusion >>
rect 125 466 126 467 
<< m1 >>
rect 136 466 137 467 
<< pdiffusion >>
rect 138 466 139 467 
<< pdiffusion >>
rect 139 466 140 467 
<< pdiffusion >>
rect 140 466 141 467 
<< pdiffusion >>
rect 141 466 142 467 
<< pdiffusion >>
rect 142 466 143 467 
<< pdiffusion >>
rect 143 466 144 467 
<< m1 >>
rect 152 466 153 467 
<< pdiffusion >>
rect 156 466 157 467 
<< pdiffusion >>
rect 157 466 158 467 
<< pdiffusion >>
rect 158 466 159 467 
<< pdiffusion >>
rect 159 466 160 467 
<< pdiffusion >>
rect 160 466 161 467 
<< pdiffusion >>
rect 161 466 162 467 
<< m1 >>
rect 163 466 164 467 
<< m1 >>
rect 172 466 173 467 
<< m2 >>
rect 172 466 173 467 
<< pdiffusion >>
rect 174 466 175 467 
<< pdiffusion >>
rect 175 466 176 467 
<< pdiffusion >>
rect 176 466 177 467 
<< pdiffusion >>
rect 177 466 178 467 
<< pdiffusion >>
rect 178 466 179 467 
<< pdiffusion >>
rect 179 466 180 467 
<< pdiffusion >>
rect 192 466 193 467 
<< pdiffusion >>
rect 193 466 194 467 
<< pdiffusion >>
rect 194 466 195 467 
<< pdiffusion >>
rect 195 466 196 467 
<< pdiffusion >>
rect 196 466 197 467 
<< pdiffusion >>
rect 197 466 198 467 
<< m1 >>
rect 199 466 200 467 
<< m1 >>
rect 208 466 209 467 
<< pdiffusion >>
rect 210 466 211 467 
<< pdiffusion >>
rect 211 466 212 467 
<< pdiffusion >>
rect 212 466 213 467 
<< pdiffusion >>
rect 213 466 214 467 
<< pdiffusion >>
rect 214 466 215 467 
<< pdiffusion >>
rect 215 466 216 467 
<< pdiffusion >>
rect 228 466 229 467 
<< pdiffusion >>
rect 229 466 230 467 
<< pdiffusion >>
rect 230 466 231 467 
<< pdiffusion >>
rect 231 466 232 467 
<< pdiffusion >>
rect 232 466 233 467 
<< pdiffusion >>
rect 233 466 234 467 
<< pdiffusion >>
rect 246 466 247 467 
<< pdiffusion >>
rect 247 466 248 467 
<< pdiffusion >>
rect 248 466 249 467 
<< pdiffusion >>
rect 249 466 250 467 
<< pdiffusion >>
rect 250 466 251 467 
<< pdiffusion >>
rect 251 466 252 467 
<< m1 >>
rect 253 466 254 467 
<< pdiffusion >>
rect 264 466 265 467 
<< pdiffusion >>
rect 265 466 266 467 
<< pdiffusion >>
rect 266 466 267 467 
<< pdiffusion >>
rect 267 466 268 467 
<< pdiffusion >>
rect 268 466 269 467 
<< pdiffusion >>
rect 269 466 270 467 
<< pdiffusion >>
rect 282 466 283 467 
<< pdiffusion >>
rect 283 466 284 467 
<< pdiffusion >>
rect 284 466 285 467 
<< pdiffusion >>
rect 285 466 286 467 
<< pdiffusion >>
rect 286 466 287 467 
<< pdiffusion >>
rect 287 466 288 467 
<< m1 >>
rect 289 466 290 467 
<< m1 >>
rect 298 466 299 467 
<< pdiffusion >>
rect 300 466 301 467 
<< pdiffusion >>
rect 301 466 302 467 
<< pdiffusion >>
rect 302 466 303 467 
<< pdiffusion >>
rect 303 466 304 467 
<< pdiffusion >>
rect 304 466 305 467 
<< pdiffusion >>
rect 305 466 306 467 
<< m1 >>
rect 307 466 308 467 
<< pdiffusion >>
rect 318 466 319 467 
<< pdiffusion >>
rect 319 466 320 467 
<< pdiffusion >>
rect 320 466 321 467 
<< pdiffusion >>
rect 321 466 322 467 
<< pdiffusion >>
rect 322 466 323 467 
<< pdiffusion >>
rect 323 466 324 467 
<< pdiffusion >>
rect 336 466 337 467 
<< pdiffusion >>
rect 337 466 338 467 
<< pdiffusion >>
rect 338 466 339 467 
<< pdiffusion >>
rect 339 466 340 467 
<< pdiffusion >>
rect 340 466 341 467 
<< pdiffusion >>
rect 341 466 342 467 
<< m1 >>
rect 352 466 353 467 
<< pdiffusion >>
rect 354 466 355 467 
<< pdiffusion >>
rect 355 466 356 467 
<< pdiffusion >>
rect 356 466 357 467 
<< pdiffusion >>
rect 357 466 358 467 
<< pdiffusion >>
rect 358 466 359 467 
<< pdiffusion >>
rect 359 466 360 467 
<< m1 >>
rect 361 466 362 467 
<< m2 >>
rect 362 466 363 467 
<< pdiffusion >>
rect 372 466 373 467 
<< pdiffusion >>
rect 373 466 374 467 
<< pdiffusion >>
rect 374 466 375 467 
<< pdiffusion >>
rect 375 466 376 467 
<< pdiffusion >>
rect 376 466 377 467 
<< pdiffusion >>
rect 377 466 378 467 
<< m1 >>
rect 381 466 382 467 
<< pdiffusion >>
rect 390 466 391 467 
<< pdiffusion >>
rect 391 466 392 467 
<< pdiffusion >>
rect 392 466 393 467 
<< pdiffusion >>
rect 393 466 394 467 
<< pdiffusion >>
rect 394 466 395 467 
<< pdiffusion >>
rect 395 466 396 467 
<< m1 >>
rect 402 466 403 467 
<< pdiffusion >>
rect 408 466 409 467 
<< pdiffusion >>
rect 409 466 410 467 
<< pdiffusion >>
rect 410 466 411 467 
<< pdiffusion >>
rect 411 466 412 467 
<< pdiffusion >>
rect 412 466 413 467 
<< pdiffusion >>
rect 413 466 414 467 
<< pdiffusion >>
rect 426 466 427 467 
<< pdiffusion >>
rect 427 466 428 467 
<< pdiffusion >>
rect 428 466 429 467 
<< pdiffusion >>
rect 429 466 430 467 
<< pdiffusion >>
rect 430 466 431 467 
<< pdiffusion >>
rect 431 466 432 467 
<< m1 >>
rect 433 466 434 467 
<< pdiffusion >>
rect 444 466 445 467 
<< pdiffusion >>
rect 445 466 446 467 
<< pdiffusion >>
rect 446 466 447 467 
<< pdiffusion >>
rect 447 466 448 467 
<< pdiffusion >>
rect 448 466 449 467 
<< pdiffusion >>
rect 449 466 450 467 
<< m1 >>
rect 451 466 452 467 
<< m2 >>
rect 451 466 452 467 
<< pdiffusion >>
rect 462 466 463 467 
<< pdiffusion >>
rect 463 466 464 467 
<< pdiffusion >>
rect 464 466 465 467 
<< pdiffusion >>
rect 465 466 466 467 
<< pdiffusion >>
rect 466 466 467 467 
<< pdiffusion >>
rect 467 466 468 467 
<< m1 >>
rect 472 466 473 467 
<< pdiffusion >>
rect 480 466 481 467 
<< pdiffusion >>
rect 481 466 482 467 
<< pdiffusion >>
rect 482 466 483 467 
<< pdiffusion >>
rect 483 466 484 467 
<< pdiffusion >>
rect 484 466 485 467 
<< pdiffusion >>
rect 485 466 486 467 
<< m1 >>
rect 487 466 488 467 
<< m1 >>
rect 489 466 490 467 
<< pdiffusion >>
rect 498 466 499 467 
<< pdiffusion >>
rect 499 466 500 467 
<< pdiffusion >>
rect 500 466 501 467 
<< pdiffusion >>
rect 501 466 502 467 
<< pdiffusion >>
rect 502 466 503 467 
<< pdiffusion >>
rect 503 466 504 467 
<< pdiffusion >>
rect 516 466 517 467 
<< pdiffusion >>
rect 517 466 518 467 
<< pdiffusion >>
rect 518 466 519 467 
<< pdiffusion >>
rect 519 466 520 467 
<< pdiffusion >>
rect 520 466 521 467 
<< pdiffusion >>
rect 521 466 522 467 
<< pdiffusion >>
rect 12 467 13 468 
<< pdiffusion >>
rect 13 467 14 468 
<< pdiffusion >>
rect 14 467 15 468 
<< pdiffusion >>
rect 15 467 16 468 
<< m1 >>
rect 16 467 17 468 
<< pdiffusion >>
rect 16 467 17 468 
<< pdiffusion >>
rect 17 467 18 468 
<< m1 >>
rect 19 467 20 468 
<< m1 >>
rect 21 467 22 468 
<< m1 >>
rect 28 467 29 468 
<< m1 >>
rect 30 467 31 468 
<< pdiffusion >>
rect 48 467 49 468 
<< pdiffusion >>
rect 49 467 50 468 
<< pdiffusion >>
rect 50 467 51 468 
<< pdiffusion >>
rect 51 467 52 468 
<< pdiffusion >>
rect 52 467 53 468 
<< pdiffusion >>
rect 53 467 54 468 
<< pdiffusion >>
rect 66 467 67 468 
<< pdiffusion >>
rect 67 467 68 468 
<< pdiffusion >>
rect 68 467 69 468 
<< pdiffusion >>
rect 69 467 70 468 
<< m1 >>
rect 70 467 71 468 
<< pdiffusion >>
rect 70 467 71 468 
<< pdiffusion >>
rect 71 467 72 468 
<< m1 >>
rect 73 467 74 468 
<< pdiffusion >>
rect 84 467 85 468 
<< pdiffusion >>
rect 85 467 86 468 
<< pdiffusion >>
rect 86 467 87 468 
<< pdiffusion >>
rect 87 467 88 468 
<< m1 >>
rect 88 467 89 468 
<< pdiffusion >>
rect 88 467 89 468 
<< pdiffusion >>
rect 89 467 90 468 
<< m1 >>
rect 100 467 101 468 
<< pdiffusion >>
rect 102 467 103 468 
<< pdiffusion >>
rect 103 467 104 468 
<< pdiffusion >>
rect 104 467 105 468 
<< pdiffusion >>
rect 105 467 106 468 
<< pdiffusion >>
rect 106 467 107 468 
<< pdiffusion >>
rect 107 467 108 468 
<< pdiffusion >>
rect 120 467 121 468 
<< pdiffusion >>
rect 121 467 122 468 
<< pdiffusion >>
rect 122 467 123 468 
<< pdiffusion >>
rect 123 467 124 468 
<< pdiffusion >>
rect 124 467 125 468 
<< pdiffusion >>
rect 125 467 126 468 
<< m1 >>
rect 136 467 137 468 
<< pdiffusion >>
rect 138 467 139 468 
<< pdiffusion >>
rect 139 467 140 468 
<< pdiffusion >>
rect 140 467 141 468 
<< pdiffusion >>
rect 141 467 142 468 
<< m1 >>
rect 142 467 143 468 
<< pdiffusion >>
rect 142 467 143 468 
<< pdiffusion >>
rect 143 467 144 468 
<< m1 >>
rect 152 467 153 468 
<< pdiffusion >>
rect 156 467 157 468 
<< pdiffusion >>
rect 157 467 158 468 
<< pdiffusion >>
rect 158 467 159 468 
<< pdiffusion >>
rect 159 467 160 468 
<< pdiffusion >>
rect 160 467 161 468 
<< pdiffusion >>
rect 161 467 162 468 
<< m1 >>
rect 163 467 164 468 
<< m1 >>
rect 172 467 173 468 
<< m2 >>
rect 172 467 173 468 
<< pdiffusion >>
rect 174 467 175 468 
<< m1 >>
rect 175 467 176 468 
<< pdiffusion >>
rect 175 467 176 468 
<< pdiffusion >>
rect 176 467 177 468 
<< pdiffusion >>
rect 177 467 178 468 
<< pdiffusion >>
rect 178 467 179 468 
<< pdiffusion >>
rect 179 467 180 468 
<< pdiffusion >>
rect 192 467 193 468 
<< pdiffusion >>
rect 193 467 194 468 
<< pdiffusion >>
rect 194 467 195 468 
<< pdiffusion >>
rect 195 467 196 468 
<< pdiffusion >>
rect 196 467 197 468 
<< pdiffusion >>
rect 197 467 198 468 
<< m1 >>
rect 199 467 200 468 
<< m1 >>
rect 208 467 209 468 
<< pdiffusion >>
rect 210 467 211 468 
<< pdiffusion >>
rect 211 467 212 468 
<< pdiffusion >>
rect 212 467 213 468 
<< pdiffusion >>
rect 213 467 214 468 
<< pdiffusion >>
rect 214 467 215 468 
<< pdiffusion >>
rect 215 467 216 468 
<< pdiffusion >>
rect 228 467 229 468 
<< pdiffusion >>
rect 229 467 230 468 
<< pdiffusion >>
rect 230 467 231 468 
<< pdiffusion >>
rect 231 467 232 468 
<< pdiffusion >>
rect 232 467 233 468 
<< pdiffusion >>
rect 233 467 234 468 
<< pdiffusion >>
rect 246 467 247 468 
<< pdiffusion >>
rect 247 467 248 468 
<< pdiffusion >>
rect 248 467 249 468 
<< pdiffusion >>
rect 249 467 250 468 
<< pdiffusion >>
rect 250 467 251 468 
<< pdiffusion >>
rect 251 467 252 468 
<< m1 >>
rect 253 467 254 468 
<< pdiffusion >>
rect 264 467 265 468 
<< pdiffusion >>
rect 265 467 266 468 
<< pdiffusion >>
rect 266 467 267 468 
<< pdiffusion >>
rect 267 467 268 468 
<< pdiffusion >>
rect 268 467 269 468 
<< pdiffusion >>
rect 269 467 270 468 
<< pdiffusion >>
rect 282 467 283 468 
<< pdiffusion >>
rect 283 467 284 468 
<< pdiffusion >>
rect 284 467 285 468 
<< pdiffusion >>
rect 285 467 286 468 
<< m1 >>
rect 286 467 287 468 
<< pdiffusion >>
rect 286 467 287 468 
<< pdiffusion >>
rect 287 467 288 468 
<< m1 >>
rect 289 467 290 468 
<< m2 >>
rect 289 467 290 468 
<< m2c >>
rect 289 467 290 468 
<< m1 >>
rect 289 467 290 468 
<< m2 >>
rect 289 467 290 468 
<< m1 >>
rect 298 467 299 468 
<< pdiffusion >>
rect 300 467 301 468 
<< pdiffusion >>
rect 301 467 302 468 
<< pdiffusion >>
rect 302 467 303 468 
<< pdiffusion >>
rect 303 467 304 468 
<< pdiffusion >>
rect 304 467 305 468 
<< pdiffusion >>
rect 305 467 306 468 
<< m1 >>
rect 307 467 308 468 
<< pdiffusion >>
rect 318 467 319 468 
<< pdiffusion >>
rect 319 467 320 468 
<< pdiffusion >>
rect 320 467 321 468 
<< pdiffusion >>
rect 321 467 322 468 
<< pdiffusion >>
rect 322 467 323 468 
<< pdiffusion >>
rect 323 467 324 468 
<< pdiffusion >>
rect 336 467 337 468 
<< pdiffusion >>
rect 337 467 338 468 
<< pdiffusion >>
rect 338 467 339 468 
<< pdiffusion >>
rect 339 467 340 468 
<< pdiffusion >>
rect 340 467 341 468 
<< pdiffusion >>
rect 341 467 342 468 
<< m1 >>
rect 352 467 353 468 
<< pdiffusion >>
rect 354 467 355 468 
<< m1 >>
rect 355 467 356 468 
<< pdiffusion >>
rect 355 467 356 468 
<< pdiffusion >>
rect 356 467 357 468 
<< pdiffusion >>
rect 357 467 358 468 
<< m1 >>
rect 358 467 359 468 
<< pdiffusion >>
rect 358 467 359 468 
<< pdiffusion >>
rect 359 467 360 468 
<< m1 >>
rect 361 467 362 468 
<< m2 >>
rect 362 467 363 468 
<< pdiffusion >>
rect 372 467 373 468 
<< m1 >>
rect 373 467 374 468 
<< pdiffusion >>
rect 373 467 374 468 
<< pdiffusion >>
rect 374 467 375 468 
<< m1 >>
rect 375 467 376 468 
<< m2 >>
rect 375 467 376 468 
<< m2c >>
rect 375 467 376 468 
<< m1 >>
rect 375 467 376 468 
<< m2 >>
rect 375 467 376 468 
<< pdiffusion >>
rect 375 467 376 468 
<< m1 >>
rect 376 467 377 468 
<< pdiffusion >>
rect 376 467 377 468 
<< pdiffusion >>
rect 377 467 378 468 
<< m1 >>
rect 381 467 382 468 
<< pdiffusion >>
rect 390 467 391 468 
<< pdiffusion >>
rect 391 467 392 468 
<< pdiffusion >>
rect 392 467 393 468 
<< pdiffusion >>
rect 393 467 394 468 
<< m1 >>
rect 394 467 395 468 
<< pdiffusion >>
rect 394 467 395 468 
<< pdiffusion >>
rect 395 467 396 468 
<< m1 >>
rect 402 467 403 468 
<< pdiffusion >>
rect 408 467 409 468 
<< pdiffusion >>
rect 409 467 410 468 
<< pdiffusion >>
rect 410 467 411 468 
<< pdiffusion >>
rect 411 467 412 468 
<< pdiffusion >>
rect 412 467 413 468 
<< pdiffusion >>
rect 413 467 414 468 
<< pdiffusion >>
rect 426 467 427 468 
<< pdiffusion >>
rect 427 467 428 468 
<< pdiffusion >>
rect 428 467 429 468 
<< pdiffusion >>
rect 429 467 430 468 
<< pdiffusion >>
rect 430 467 431 468 
<< pdiffusion >>
rect 431 467 432 468 
<< m1 >>
rect 433 467 434 468 
<< pdiffusion >>
rect 444 467 445 468 
<< m1 >>
rect 445 467 446 468 
<< pdiffusion >>
rect 445 467 446 468 
<< pdiffusion >>
rect 446 467 447 468 
<< pdiffusion >>
rect 447 467 448 468 
<< pdiffusion >>
rect 448 467 449 468 
<< pdiffusion >>
rect 449 467 450 468 
<< m1 >>
rect 451 467 452 468 
<< m2 >>
rect 451 467 452 468 
<< pdiffusion >>
rect 462 467 463 468 
<< pdiffusion >>
rect 463 467 464 468 
<< pdiffusion >>
rect 464 467 465 468 
<< pdiffusion >>
rect 465 467 466 468 
<< pdiffusion >>
rect 466 467 467 468 
<< pdiffusion >>
rect 467 467 468 468 
<< m1 >>
rect 472 467 473 468 
<< pdiffusion >>
rect 480 467 481 468 
<< pdiffusion >>
rect 481 467 482 468 
<< pdiffusion >>
rect 482 467 483 468 
<< pdiffusion >>
rect 483 467 484 468 
<< pdiffusion >>
rect 484 467 485 468 
<< pdiffusion >>
rect 485 467 486 468 
<< m1 >>
rect 487 467 488 468 
<< m1 >>
rect 489 467 490 468 
<< pdiffusion >>
rect 498 467 499 468 
<< pdiffusion >>
rect 499 467 500 468 
<< pdiffusion >>
rect 500 467 501 468 
<< pdiffusion >>
rect 501 467 502 468 
<< pdiffusion >>
rect 502 467 503 468 
<< pdiffusion >>
rect 503 467 504 468 
<< pdiffusion >>
rect 516 467 517 468 
<< pdiffusion >>
rect 517 467 518 468 
<< pdiffusion >>
rect 518 467 519 468 
<< pdiffusion >>
rect 519 467 520 468 
<< pdiffusion >>
rect 520 467 521 468 
<< pdiffusion >>
rect 521 467 522 468 
<< m1 >>
rect 16 468 17 469 
<< m1 >>
rect 19 468 20 469 
<< m1 >>
rect 21 468 22 469 
<< m1 >>
rect 28 468 29 469 
<< m1 >>
rect 30 468 31 469 
<< m1 >>
rect 70 468 71 469 
<< m1 >>
rect 73 468 74 469 
<< m1 >>
rect 88 468 89 469 
<< m1 >>
rect 100 468 101 469 
<< m1 >>
rect 136 468 137 469 
<< m1 >>
rect 142 468 143 469 
<< m1 >>
rect 145 468 146 469 
<< m2 >>
rect 145 468 146 469 
<< m2c >>
rect 145 468 146 469 
<< m1 >>
rect 145 468 146 469 
<< m2 >>
rect 145 468 146 469 
<< m1 >>
rect 146 468 147 469 
<< m1 >>
rect 147 468 148 469 
<< m1 >>
rect 148 468 149 469 
<< m1 >>
rect 149 468 150 469 
<< m1 >>
rect 150 468 151 469 
<< m1 >>
rect 151 468 152 469 
<< m1 >>
rect 152 468 153 469 
<< m1 >>
rect 163 468 164 469 
<< m1 >>
rect 172 468 173 469 
<< m2 >>
rect 172 468 173 469 
<< m1 >>
rect 175 468 176 469 
<< m1 >>
rect 199 468 200 469 
<< m1 >>
rect 208 468 209 469 
<< m1 >>
rect 253 468 254 469 
<< m1 >>
rect 286 468 287 469 
<< m2 >>
rect 289 468 290 469 
<< m1 >>
rect 298 468 299 469 
<< m1 >>
rect 307 468 308 469 
<< m1 >>
rect 352 468 353 469 
<< m1 >>
rect 355 468 356 469 
<< m1 >>
rect 358 468 359 469 
<< m1 >>
rect 361 468 362 469 
<< m2 >>
rect 362 468 363 469 
<< m1 >>
rect 373 468 374 469 
<< m1 >>
rect 376 468 377 469 
<< m2 >>
rect 376 468 377 469 
<< m1 >>
rect 381 468 382 469 
<< m1 >>
rect 394 468 395 469 
<< m1 >>
rect 402 468 403 469 
<< m1 >>
rect 433 468 434 469 
<< m1 >>
rect 445 468 446 469 
<< m1 >>
rect 451 468 452 469 
<< m2 >>
rect 451 468 452 469 
<< m1 >>
rect 472 468 473 469 
<< m1 >>
rect 487 468 488 469 
<< m1 >>
rect 489 468 490 469 
<< m1 >>
rect 16 469 17 470 
<< m1 >>
rect 17 469 18 470 
<< m1 >>
rect 18 469 19 470 
<< m1 >>
rect 19 469 20 470 
<< m1 >>
rect 21 469 22 470 
<< m1 >>
rect 28 469 29 470 
<< m1 >>
rect 30 469 31 470 
<< m1 >>
rect 70 469 71 470 
<< m1 >>
rect 73 469 74 470 
<< m1 >>
rect 88 469 89 470 
<< m1 >>
rect 100 469 101 470 
<< m1 >>
rect 136 469 137 470 
<< m1 >>
rect 142 469 143 470 
<< m2 >>
rect 145 469 146 470 
<< m1 >>
rect 163 469 164 470 
<< m1 >>
rect 172 469 173 470 
<< m2 >>
rect 172 469 173 470 
<< m2 >>
rect 173 469 174 470 
<< m1 >>
rect 174 469 175 470 
<< m2 >>
rect 174 469 175 470 
<< m2c >>
rect 174 469 175 470 
<< m1 >>
rect 174 469 175 470 
<< m2 >>
rect 174 469 175 470 
<< m1 >>
rect 175 469 176 470 
<< m1 >>
rect 199 469 200 470 
<< m1 >>
rect 208 469 209 470 
<< m1 >>
rect 253 469 254 470 
<< m1 >>
rect 286 469 287 470 
<< m1 >>
rect 287 469 288 470 
<< m1 >>
rect 288 469 289 470 
<< m1 >>
rect 289 469 290 470 
<< m2 >>
rect 289 469 290 470 
<< m1 >>
rect 290 469 291 470 
<< m1 >>
rect 291 469 292 470 
<< m1 >>
rect 292 469 293 470 
<< m1 >>
rect 293 469 294 470 
<< m1 >>
rect 294 469 295 470 
<< m1 >>
rect 295 469 296 470 
<< m1 >>
rect 296 469 297 470 
<< m1 >>
rect 297 469 298 470 
<< m1 >>
rect 298 469 299 470 
<< m1 >>
rect 307 469 308 470 
<< m1 >>
rect 352 469 353 470 
<< m1 >>
rect 355 469 356 470 
<< m1 >>
rect 358 469 359 470 
<< m1 >>
rect 359 469 360 470 
<< m1 >>
rect 360 469 361 470 
<< m1 >>
rect 361 469 362 470 
<< m2 >>
rect 362 469 363 470 
<< m1 >>
rect 373 469 374 470 
<< m2 >>
rect 376 469 377 470 
<< m1 >>
rect 381 469 382 470 
<< m1 >>
rect 394 469 395 470 
<< m2 >>
rect 395 469 396 470 
<< m1 >>
rect 396 469 397 470 
<< m2 >>
rect 396 469 397 470 
<< m2c >>
rect 396 469 397 470 
<< m1 >>
rect 396 469 397 470 
<< m2 >>
rect 396 469 397 470 
<< m1 >>
rect 397 469 398 470 
<< m1 >>
rect 398 469 399 470 
<< m1 >>
rect 399 469 400 470 
<< m1 >>
rect 400 469 401 470 
<< m1 >>
rect 401 469 402 470 
<< m1 >>
rect 402 469 403 470 
<< m1 >>
rect 433 469 434 470 
<< m1 >>
rect 445 469 446 470 
<< m1 >>
rect 451 469 452 470 
<< m2 >>
rect 451 469 452 470 
<< m1 >>
rect 472 469 473 470 
<< m1 >>
rect 487 469 488 470 
<< m1 >>
rect 489 469 490 470 
<< m1 >>
rect 21 470 22 471 
<< m1 >>
rect 28 470 29 471 
<< m1 >>
rect 30 470 31 471 
<< m1 >>
rect 70 470 71 471 
<< m1 >>
rect 73 470 74 471 
<< m1 >>
rect 88 470 89 471 
<< m1 >>
rect 89 470 90 471 
<< m1 >>
rect 90 470 91 471 
<< m1 >>
rect 91 470 92 471 
<< m1 >>
rect 92 470 93 471 
<< m1 >>
rect 93 470 94 471 
<< m1 >>
rect 94 470 95 471 
<< m1 >>
rect 95 470 96 471 
<< m1 >>
rect 96 470 97 471 
<< m1 >>
rect 97 470 98 471 
<< m1 >>
rect 98 470 99 471 
<< m2 >>
rect 98 470 99 471 
<< m2c >>
rect 98 470 99 471 
<< m1 >>
rect 98 470 99 471 
<< m2 >>
rect 98 470 99 471 
<< m2 >>
rect 99 470 100 471 
<< m1 >>
rect 100 470 101 471 
<< m2 >>
rect 100 470 101 471 
<< m2 >>
rect 101 470 102 471 
<< m1 >>
rect 136 470 137 471 
<< m1 >>
rect 142 470 143 471 
<< m1 >>
rect 143 470 144 471 
<< m1 >>
rect 144 470 145 471 
<< m1 >>
rect 145 470 146 471 
<< m2 >>
rect 145 470 146 471 
<< m1 >>
rect 146 470 147 471 
<< m1 >>
rect 147 470 148 471 
<< m1 >>
rect 148 470 149 471 
<< m1 >>
rect 149 470 150 471 
<< m1 >>
rect 150 470 151 471 
<< m1 >>
rect 151 470 152 471 
<< m1 >>
rect 152 470 153 471 
<< m1 >>
rect 153 470 154 471 
<< m1 >>
rect 154 470 155 471 
<< m1 >>
rect 155 470 156 471 
<< m1 >>
rect 156 470 157 471 
<< m1 >>
rect 163 470 164 471 
<< m1 >>
rect 172 470 173 471 
<< m1 >>
rect 199 470 200 471 
<< m1 >>
rect 208 470 209 471 
<< m1 >>
rect 253 470 254 471 
<< m2 >>
rect 286 470 287 471 
<< m2 >>
rect 287 470 288 471 
<< m2 >>
rect 288 470 289 471 
<< m2 >>
rect 289 470 290 471 
<< m1 >>
rect 307 470 308 471 
<< m1 >>
rect 352 470 353 471 
<< m1 >>
rect 355 470 356 471 
<< m2 >>
rect 362 470 363 471 
<< m1 >>
rect 363 470 364 471 
<< m2 >>
rect 363 470 364 471 
<< m2c >>
rect 363 470 364 471 
<< m1 >>
rect 363 470 364 471 
<< m2 >>
rect 363 470 364 471 
<< m1 >>
rect 364 470 365 471 
<< m1 >>
rect 365 470 366 471 
<< m1 >>
rect 366 470 367 471 
<< m1 >>
rect 367 470 368 471 
<< m1 >>
rect 368 470 369 471 
<< m1 >>
rect 369 470 370 471 
<< m1 >>
rect 370 470 371 471 
<< m1 >>
rect 371 470 372 471 
<< m1 >>
rect 373 470 374 471 
<< m1 >>
rect 374 470 375 471 
<< m1 >>
rect 375 470 376 471 
<< m1 >>
rect 376 470 377 471 
<< m2 >>
rect 376 470 377 471 
<< m1 >>
rect 377 470 378 471 
<< m1 >>
rect 378 470 379 471 
<< m1 >>
rect 379 470 380 471 
<< m1 >>
rect 381 470 382 471 
<< m1 >>
rect 394 470 395 471 
<< m2 >>
rect 395 470 396 471 
<< m1 >>
rect 433 470 434 471 
<< m1 >>
rect 445 470 446 471 
<< m1 >>
rect 446 470 447 471 
<< m1 >>
rect 447 470 448 471 
<< m1 >>
rect 448 470 449 471 
<< m1 >>
rect 449 470 450 471 
<< m2 >>
rect 449 470 450 471 
<< m2c >>
rect 449 470 450 471 
<< m1 >>
rect 449 470 450 471 
<< m2 >>
rect 449 470 450 471 
<< m2 >>
rect 450 470 451 471 
<< m1 >>
rect 451 470 452 471 
<< m2 >>
rect 451 470 452 471 
<< m1 >>
rect 472 470 473 471 
<< m1 >>
rect 487 470 488 471 
<< m1 >>
rect 489 470 490 471 
<< m1 >>
rect 21 471 22 472 
<< m1 >>
rect 28 471 29 472 
<< m1 >>
rect 30 471 31 472 
<< m1 >>
rect 70 471 71 472 
<< m1 >>
rect 73 471 74 472 
<< m1 >>
rect 100 471 101 472 
<< m2 >>
rect 101 471 102 472 
<< m1 >>
rect 136 471 137 472 
<< m2 >>
rect 140 471 141 472 
<< m2 >>
rect 141 471 142 472 
<< m2 >>
rect 142 471 143 472 
<< m2 >>
rect 143 471 144 472 
<< m2 >>
rect 144 471 145 472 
<< m2 >>
rect 145 471 146 472 
<< m1 >>
rect 156 471 157 472 
<< m1 >>
rect 163 471 164 472 
<< m1 >>
rect 164 471 165 472 
<< m1 >>
rect 165 471 166 472 
<< m1 >>
rect 166 471 167 472 
<< m1 >>
rect 167 471 168 472 
<< m1 >>
rect 168 471 169 472 
<< m1 >>
rect 169 471 170 472 
<< m1 >>
rect 170 471 171 472 
<< m2 >>
rect 170 471 171 472 
<< m2c >>
rect 170 471 171 472 
<< m1 >>
rect 170 471 171 472 
<< m2 >>
rect 170 471 171 472 
<< m2 >>
rect 171 471 172 472 
<< m1 >>
rect 172 471 173 472 
<< m2 >>
rect 172 471 173 472 
<< m2 >>
rect 173 471 174 472 
<< m1 >>
rect 174 471 175 472 
<< m2 >>
rect 174 471 175 472 
<< m2c >>
rect 174 471 175 472 
<< m1 >>
rect 174 471 175 472 
<< m2 >>
rect 174 471 175 472 
<< m1 >>
rect 199 471 200 472 
<< m1 >>
rect 208 471 209 472 
<< m1 >>
rect 253 471 254 472 
<< m1 >>
rect 286 471 287 472 
<< m2 >>
rect 286 471 287 472 
<< m2c >>
rect 286 471 287 472 
<< m1 >>
rect 286 471 287 472 
<< m2 >>
rect 286 471 287 472 
<< m1 >>
rect 307 471 308 472 
<< m1 >>
rect 352 471 353 472 
<< m1 >>
rect 355 471 356 472 
<< m1 >>
rect 371 471 372 472 
<< m2 >>
rect 376 471 377 472 
<< m1 >>
rect 379 471 380 472 
<< m1 >>
rect 381 471 382 472 
<< m1 >>
rect 394 471 395 472 
<< m2 >>
rect 395 471 396 472 
<< m1 >>
rect 433 471 434 472 
<< m1 >>
rect 451 471 452 472 
<< m1 >>
rect 472 471 473 472 
<< m1 >>
rect 487 471 488 472 
<< m1 >>
rect 489 471 490 472 
<< m1 >>
rect 21 472 22 473 
<< m1 >>
rect 28 472 29 473 
<< m1 >>
rect 30 472 31 473 
<< m1 >>
rect 31 472 32 473 
<< m1 >>
rect 32 472 33 473 
<< m1 >>
rect 33 472 34 473 
<< m1 >>
rect 34 472 35 473 
<< m1 >>
rect 35 472 36 473 
<< m1 >>
rect 36 472 37 473 
<< m1 >>
rect 37 472 38 473 
<< m1 >>
rect 38 472 39 473 
<< m1 >>
rect 39 472 40 473 
<< m1 >>
rect 40 472 41 473 
<< m1 >>
rect 41 472 42 473 
<< m1 >>
rect 42 472 43 473 
<< m1 >>
rect 43 472 44 473 
<< m1 >>
rect 44 472 45 473 
<< m1 >>
rect 45 472 46 473 
<< m1 >>
rect 46 472 47 473 
<< m1 >>
rect 47 472 48 473 
<< m1 >>
rect 48 472 49 473 
<< m1 >>
rect 49 472 50 473 
<< m1 >>
rect 70 472 71 473 
<< m1 >>
rect 73 472 74 473 
<< m1 >>
rect 85 472 86 473 
<< m1 >>
rect 86 472 87 473 
<< m1 >>
rect 87 472 88 473 
<< m1 >>
rect 88 472 89 473 
<< m1 >>
rect 89 472 90 473 
<< m1 >>
rect 90 472 91 473 
<< m1 >>
rect 91 472 92 473 
<< m1 >>
rect 92 472 93 473 
<< m1 >>
rect 93 472 94 473 
<< m1 >>
rect 94 472 95 473 
<< m1 >>
rect 95 472 96 473 
<< m1 >>
rect 96 472 97 473 
<< m1 >>
rect 97 472 98 473 
<< m1 >>
rect 98 472 99 473 
<< m1 >>
rect 99 472 100 473 
<< m1 >>
rect 100 472 101 473 
<< m2 >>
rect 101 472 102 473 
<< m1 >>
rect 136 472 137 473 
<< m1 >>
rect 137 472 138 473 
<< m1 >>
rect 138 472 139 473 
<< m1 >>
rect 139 472 140 473 
<< m1 >>
rect 140 472 141 473 
<< m2 >>
rect 140 472 141 473 
<< m1 >>
rect 141 472 142 473 
<< m1 >>
rect 142 472 143 473 
<< m1 >>
rect 156 472 157 473 
<< m1 >>
rect 172 472 173 473 
<< m1 >>
rect 174 472 175 473 
<< m1 >>
rect 175 472 176 473 
<< m1 >>
rect 176 472 177 473 
<< m1 >>
rect 177 472 178 473 
<< m1 >>
rect 178 472 179 473 
<< m1 >>
rect 179 472 180 473 
<< m1 >>
rect 180 472 181 473 
<< m1 >>
rect 181 472 182 473 
<< m1 >>
rect 182 472 183 473 
<< m1 >>
rect 183 472 184 473 
<< m1 >>
rect 184 472 185 473 
<< m1 >>
rect 185 472 186 473 
<< m1 >>
rect 186 472 187 473 
<< m1 >>
rect 187 472 188 473 
<< m1 >>
rect 188 472 189 473 
<< m1 >>
rect 189 472 190 473 
<< m1 >>
rect 190 472 191 473 
<< m1 >>
rect 191 472 192 473 
<< m1 >>
rect 192 472 193 473 
<< m1 >>
rect 193 472 194 473 
<< m1 >>
rect 194 472 195 473 
<< m1 >>
rect 195 472 196 473 
<< m1 >>
rect 196 472 197 473 
<< m1 >>
rect 197 472 198 473 
<< m1 >>
rect 198 472 199 473 
<< m1 >>
rect 199 472 200 473 
<< m1 >>
rect 208 472 209 473 
<< m1 >>
rect 253 472 254 473 
<< m1 >>
rect 286 472 287 473 
<< m1 >>
rect 307 472 308 473 
<< m1 >>
rect 352 472 353 473 
<< m1 >>
rect 355 472 356 473 
<< m1 >>
rect 371 472 372 473 
<< m1 >>
rect 372 472 373 473 
<< m1 >>
rect 373 472 374 473 
<< m1 >>
rect 374 472 375 473 
<< m1 >>
rect 375 472 376 473 
<< m1 >>
rect 376 472 377 473 
<< m2 >>
rect 376 472 377 473 
<< m2c >>
rect 376 472 377 473 
<< m1 >>
rect 376 472 377 473 
<< m2 >>
rect 376 472 377 473 
<< m1 >>
rect 379 472 380 473 
<< m1 >>
rect 381 472 382 473 
<< m1 >>
rect 394 472 395 473 
<< m2 >>
rect 395 472 396 473 
<< m1 >>
rect 433 472 434 473 
<< m1 >>
rect 451 472 452 473 
<< m1 >>
rect 472 472 473 473 
<< m1 >>
rect 487 472 488 473 
<< m1 >>
rect 489 472 490 473 
<< m1 >>
rect 21 473 22 474 
<< m1 >>
rect 28 473 29 474 
<< m1 >>
rect 49 473 50 474 
<< m1 >>
rect 70 473 71 474 
<< m1 >>
rect 73 473 74 474 
<< m1 >>
rect 85 473 86 474 
<< m2 >>
rect 101 473 102 474 
<< m1 >>
rect 102 473 103 474 
<< m2 >>
rect 102 473 103 474 
<< m2c >>
rect 102 473 103 474 
<< m1 >>
rect 102 473 103 474 
<< m2 >>
rect 102 473 103 474 
<< m1 >>
rect 103 473 104 474 
<< m1 >>
rect 104 473 105 474 
<< m1 >>
rect 105 473 106 474 
<< m1 >>
rect 106 473 107 474 
<< m1 >>
rect 107 473 108 474 
<< m1 >>
rect 108 473 109 474 
<< m1 >>
rect 109 473 110 474 
<< m1 >>
rect 110 473 111 474 
<< m1 >>
rect 111 473 112 474 
<< m1 >>
rect 112 473 113 474 
<< m1 >>
rect 113 473 114 474 
<< m1 >>
rect 114 473 115 474 
<< m1 >>
rect 115 473 116 474 
<< m1 >>
rect 116 473 117 474 
<< m1 >>
rect 117 473 118 474 
<< m1 >>
rect 118 473 119 474 
<< m1 >>
rect 119 473 120 474 
<< m1 >>
rect 120 473 121 474 
<< m1 >>
rect 121 473 122 474 
<< m2 >>
rect 135 473 136 474 
<< m2 >>
rect 136 473 137 474 
<< m2 >>
rect 137 473 138 474 
<< m2 >>
rect 138 473 139 474 
<< m2 >>
rect 139 473 140 474 
<< m2 >>
rect 140 473 141 474 
<< m1 >>
rect 142 473 143 474 
<< m1 >>
rect 156 473 157 474 
<< m1 >>
rect 172 473 173 474 
<< m1 >>
rect 208 473 209 474 
<< m1 >>
rect 253 473 254 474 
<< m1 >>
rect 255 473 256 474 
<< m1 >>
rect 256 473 257 474 
<< m1 >>
rect 257 473 258 474 
<< m1 >>
rect 258 473 259 474 
<< m1 >>
rect 259 473 260 474 
<< m1 >>
rect 260 473 261 474 
<< m1 >>
rect 261 473 262 474 
<< m1 >>
rect 262 473 263 474 
<< m1 >>
rect 263 473 264 474 
<< m1 >>
rect 264 473 265 474 
<< m1 >>
rect 265 473 266 474 
<< m1 >>
rect 266 473 267 474 
<< m1 >>
rect 267 473 268 474 
<< m1 >>
rect 268 473 269 474 
<< m1 >>
rect 269 473 270 474 
<< m1 >>
rect 270 473 271 474 
<< m1 >>
rect 271 473 272 474 
<< m1 >>
rect 272 473 273 474 
<< m1 >>
rect 273 473 274 474 
<< m1 >>
rect 274 473 275 474 
<< m1 >>
rect 275 473 276 474 
<< m1 >>
rect 276 473 277 474 
<< m1 >>
rect 277 473 278 474 
<< m1 >>
rect 278 473 279 474 
<< m1 >>
rect 279 473 280 474 
<< m1 >>
rect 280 473 281 474 
<< m1 >>
rect 281 473 282 474 
<< m1 >>
rect 282 473 283 474 
<< m1 >>
rect 283 473 284 474 
<< m1 >>
rect 284 473 285 474 
<< m2 >>
rect 284 473 285 474 
<< m2c >>
rect 284 473 285 474 
<< m1 >>
rect 284 473 285 474 
<< m2 >>
rect 284 473 285 474 
<< m2 >>
rect 285 473 286 474 
<< m1 >>
rect 286 473 287 474 
<< m2 >>
rect 286 473 287 474 
<< m2 >>
rect 287 473 288 474 
<< m1 >>
rect 288 473 289 474 
<< m2 >>
rect 288 473 289 474 
<< m2c >>
rect 288 473 289 474 
<< m1 >>
rect 288 473 289 474 
<< m2 >>
rect 288 473 289 474 
<< m1 >>
rect 289 473 290 474 
<< m1 >>
rect 290 473 291 474 
<< m2 >>
rect 290 473 291 474 
<< m2c >>
rect 290 473 291 474 
<< m1 >>
rect 290 473 291 474 
<< m2 >>
rect 290 473 291 474 
<< m1 >>
rect 307 473 308 474 
<< m1 >>
rect 352 473 353 474 
<< m2 >>
rect 352 473 353 474 
<< m2c >>
rect 352 473 353 474 
<< m1 >>
rect 352 473 353 474 
<< m2 >>
rect 352 473 353 474 
<< m1 >>
rect 355 473 356 474 
<< m2 >>
rect 355 473 356 474 
<< m2c >>
rect 355 473 356 474 
<< m1 >>
rect 355 473 356 474 
<< m2 >>
rect 355 473 356 474 
<< m1 >>
rect 379 473 380 474 
<< m1 >>
rect 381 473 382 474 
<< m1 >>
rect 394 473 395 474 
<< m2 >>
rect 395 473 396 474 
<< m1 >>
rect 433 473 434 474 
<< m1 >>
rect 451 473 452 474 
<< m1 >>
rect 472 473 473 474 
<< m1 >>
rect 487 473 488 474 
<< m1 >>
rect 489 473 490 474 
<< m1 >>
rect 21 474 22 475 
<< m1 >>
rect 28 474 29 475 
<< m1 >>
rect 49 474 50 475 
<< m1 >>
rect 70 474 71 475 
<< m1 >>
rect 73 474 74 475 
<< m1 >>
rect 85 474 86 475 
<< m1 >>
rect 121 474 122 475 
<< m1 >>
rect 135 474 136 475 
<< m2 >>
rect 135 474 136 475 
<< m2c >>
rect 135 474 136 475 
<< m1 >>
rect 135 474 136 475 
<< m2 >>
rect 135 474 136 475 
<< m1 >>
rect 142 474 143 475 
<< m1 >>
rect 156 474 157 475 
<< m1 >>
rect 172 474 173 475 
<< m1 >>
rect 208 474 209 475 
<< m1 >>
rect 253 474 254 475 
<< m1 >>
rect 255 474 256 475 
<< m1 >>
rect 286 474 287 475 
<< m2 >>
rect 290 474 291 475 
<< m2 >>
rect 291 474 292 475 
<< m2 >>
rect 292 474 293 475 
<< m2 >>
rect 293 474 294 475 
<< m2 >>
rect 294 474 295 475 
<< m2 >>
rect 295 474 296 475 
<< m2 >>
rect 296 474 297 475 
<< m2 >>
rect 297 474 298 475 
<< m2 >>
rect 298 474 299 475 
<< m2 >>
rect 299 474 300 475 
<< m2 >>
rect 300 474 301 475 
<< m2 >>
rect 301 474 302 475 
<< m2 >>
rect 302 474 303 475 
<< m1 >>
rect 307 474 308 475 
<< m2 >>
rect 352 474 353 475 
<< m2 >>
rect 355 474 356 475 
<< m2 >>
rect 356 474 357 475 
<< m1 >>
rect 379 474 380 475 
<< m1 >>
rect 381 474 382 475 
<< m2 >>
rect 390 474 391 475 
<< m2 >>
rect 391 474 392 475 
<< m2 >>
rect 392 474 393 475 
<< m2 >>
rect 393 474 394 475 
<< m1 >>
rect 394 474 395 475 
<< m2 >>
rect 394 474 395 475 
<< m2 >>
rect 395 474 396 475 
<< m1 >>
rect 433 474 434 475 
<< m1 >>
rect 451 474 452 475 
<< m1 >>
rect 472 474 473 475 
<< m1 >>
rect 487 474 488 475 
<< m1 >>
rect 489 474 490 475 
<< m1 >>
rect 21 475 22 476 
<< m1 >>
rect 28 475 29 476 
<< m1 >>
rect 49 475 50 476 
<< m1 >>
rect 70 475 71 476 
<< m1 >>
rect 73 475 74 476 
<< m1 >>
rect 85 475 86 476 
<< m1 >>
rect 121 475 122 476 
<< m1 >>
rect 135 475 136 476 
<< m1 >>
rect 142 475 143 476 
<< m1 >>
rect 156 475 157 476 
<< m1 >>
rect 157 475 158 476 
<< m1 >>
rect 158 475 159 476 
<< m1 >>
rect 159 475 160 476 
<< m1 >>
rect 160 475 161 476 
<< m1 >>
rect 161 475 162 476 
<< m1 >>
rect 162 475 163 476 
<< m1 >>
rect 163 475 164 476 
<< m1 >>
rect 164 475 165 476 
<< m1 >>
rect 165 475 166 476 
<< m1 >>
rect 166 475 167 476 
<< m1 >>
rect 167 475 168 476 
<< m1 >>
rect 168 475 169 476 
<< m1 >>
rect 169 475 170 476 
<< m1 >>
rect 170 475 171 476 
<< m2 >>
rect 170 475 171 476 
<< m2c >>
rect 170 475 171 476 
<< m1 >>
rect 170 475 171 476 
<< m2 >>
rect 170 475 171 476 
<< m2 >>
rect 171 475 172 476 
<< m1 >>
rect 172 475 173 476 
<< m2 >>
rect 172 475 173 476 
<< m2 >>
rect 173 475 174 476 
<< m1 >>
rect 174 475 175 476 
<< m2 >>
rect 174 475 175 476 
<< m2c >>
rect 174 475 175 476 
<< m1 >>
rect 174 475 175 476 
<< m2 >>
rect 174 475 175 476 
<< m1 >>
rect 175 475 176 476 
<< m1 >>
rect 176 475 177 476 
<< m1 >>
rect 177 475 178 476 
<< m1 >>
rect 178 475 179 476 
<< m2 >>
rect 178 475 179 476 
<< m2c >>
rect 178 475 179 476 
<< m1 >>
rect 178 475 179 476 
<< m2 >>
rect 178 475 179 476 
<< m1 >>
rect 208 475 209 476 
<< m1 >>
rect 253 475 254 476 
<< m1 >>
rect 255 475 256 476 
<< m1 >>
rect 271 475 272 476 
<< m1 >>
rect 272 475 273 476 
<< m1 >>
rect 273 475 274 476 
<< m1 >>
rect 274 475 275 476 
<< m1 >>
rect 275 475 276 476 
<< m1 >>
rect 276 475 277 476 
<< m1 >>
rect 277 475 278 476 
<< m1 >>
rect 278 475 279 476 
<< m1 >>
rect 279 475 280 476 
<< m1 >>
rect 280 475 281 476 
<< m1 >>
rect 281 475 282 476 
<< m1 >>
rect 282 475 283 476 
<< m1 >>
rect 283 475 284 476 
<< m1 >>
rect 284 475 285 476 
<< m2 >>
rect 284 475 285 476 
<< m2c >>
rect 284 475 285 476 
<< m1 >>
rect 284 475 285 476 
<< m2 >>
rect 284 475 285 476 
<< m2 >>
rect 285 475 286 476 
<< m1 >>
rect 286 475 287 476 
<< m2 >>
rect 286 475 287 476 
<< m2 >>
rect 287 475 288 476 
<< m1 >>
rect 288 475 289 476 
<< m2 >>
rect 288 475 289 476 
<< m2c >>
rect 288 475 289 476 
<< m1 >>
rect 288 475 289 476 
<< m2 >>
rect 288 475 289 476 
<< m1 >>
rect 289 475 290 476 
<< m1 >>
rect 290 475 291 476 
<< m1 >>
rect 291 475 292 476 
<< m1 >>
rect 292 475 293 476 
<< m1 >>
rect 293 475 294 476 
<< m1 >>
rect 294 475 295 476 
<< m1 >>
rect 295 475 296 476 
<< m1 >>
rect 296 475 297 476 
<< m1 >>
rect 297 475 298 476 
<< m1 >>
rect 298 475 299 476 
<< m1 >>
rect 299 475 300 476 
<< m1 >>
rect 300 475 301 476 
<< m1 >>
rect 301 475 302 476 
<< m1 >>
rect 302 475 303 476 
<< m2 >>
rect 302 475 303 476 
<< m1 >>
rect 303 475 304 476 
<< m1 >>
rect 304 475 305 476 
<< m1 >>
rect 305 475 306 476 
<< m2 >>
rect 305 475 306 476 
<< m2c >>
rect 305 475 306 476 
<< m1 >>
rect 305 475 306 476 
<< m2 >>
rect 305 475 306 476 
<< m2 >>
rect 306 475 307 476 
<< m1 >>
rect 307 475 308 476 
<< m2 >>
rect 307 475 308 476 
<< m2 >>
rect 308 475 309 476 
<< m1 >>
rect 309 475 310 476 
<< m2 >>
rect 309 475 310 476 
<< m2c >>
rect 309 475 310 476 
<< m1 >>
rect 309 475 310 476 
<< m2 >>
rect 309 475 310 476 
<< m1 >>
rect 310 475 311 476 
<< m1 >>
rect 311 475 312 476 
<< m1 >>
rect 312 475 313 476 
<< m1 >>
rect 313 475 314 476 
<< m1 >>
rect 314 475 315 476 
<< m1 >>
rect 315 475 316 476 
<< m1 >>
rect 316 475 317 476 
<< m1 >>
rect 317 475 318 476 
<< m1 >>
rect 318 475 319 476 
<< m1 >>
rect 319 475 320 476 
<< m1 >>
rect 320 475 321 476 
<< m1 >>
rect 321 475 322 476 
<< m1 >>
rect 322 475 323 476 
<< m1 >>
rect 323 475 324 476 
<< m1 >>
rect 324 475 325 476 
<< m1 >>
rect 325 475 326 476 
<< m1 >>
rect 326 475 327 476 
<< m1 >>
rect 327 475 328 476 
<< m1 >>
rect 328 475 329 476 
<< m1 >>
rect 329 475 330 476 
<< m1 >>
rect 330 475 331 476 
<< m1 >>
rect 331 475 332 476 
<< m1 >>
rect 332 475 333 476 
<< m1 >>
rect 333 475 334 476 
<< m1 >>
rect 334 475 335 476 
<< m1 >>
rect 335 475 336 476 
<< m1 >>
rect 336 475 337 476 
<< m1 >>
rect 337 475 338 476 
<< m1 >>
rect 338 475 339 476 
<< m1 >>
rect 339 475 340 476 
<< m1 >>
rect 340 475 341 476 
<< m1 >>
rect 341 475 342 476 
<< m1 >>
rect 342 475 343 476 
<< m1 >>
rect 343 475 344 476 
<< m1 >>
rect 344 475 345 476 
<< m1 >>
rect 345 475 346 476 
<< m1 >>
rect 346 475 347 476 
<< m1 >>
rect 347 475 348 476 
<< m1 >>
rect 348 475 349 476 
<< m1 >>
rect 349 475 350 476 
<< m1 >>
rect 350 475 351 476 
<< m1 >>
rect 351 475 352 476 
<< m1 >>
rect 352 475 353 476 
<< m2 >>
rect 352 475 353 476 
<< m1 >>
rect 353 475 354 476 
<< m1 >>
rect 354 475 355 476 
<< m1 >>
rect 355 475 356 476 
<< m1 >>
rect 356 475 357 476 
<< m2 >>
rect 356 475 357 476 
<< m1 >>
rect 357 475 358 476 
<< m1 >>
rect 358 475 359 476 
<< m1 >>
rect 359 475 360 476 
<< m1 >>
rect 360 475 361 476 
<< m1 >>
rect 361 475 362 476 
<< m1 >>
rect 362 475 363 476 
<< m1 >>
rect 363 475 364 476 
<< m1 >>
rect 364 475 365 476 
<< m1 >>
rect 365 475 366 476 
<< m1 >>
rect 366 475 367 476 
<< m1 >>
rect 367 475 368 476 
<< m1 >>
rect 368 475 369 476 
<< m1 >>
rect 369 475 370 476 
<< m1 >>
rect 370 475 371 476 
<< m1 >>
rect 371 475 372 476 
<< m1 >>
rect 372 475 373 476 
<< m1 >>
rect 373 475 374 476 
<< m1 >>
rect 374 475 375 476 
<< m1 >>
rect 375 475 376 476 
<< m1 >>
rect 376 475 377 476 
<< m1 >>
rect 377 475 378 476 
<< m2 >>
rect 377 475 378 476 
<< m2c >>
rect 377 475 378 476 
<< m1 >>
rect 377 475 378 476 
<< m2 >>
rect 377 475 378 476 
<< m2 >>
rect 378 475 379 476 
<< m1 >>
rect 379 475 380 476 
<< m2 >>
rect 379 475 380 476 
<< m2 >>
rect 380 475 381 476 
<< m1 >>
rect 381 475 382 476 
<< m2 >>
rect 381 475 382 476 
<< m2 >>
rect 382 475 383 476 
<< m1 >>
rect 383 475 384 476 
<< m2 >>
rect 383 475 384 476 
<< m2c >>
rect 383 475 384 476 
<< m1 >>
rect 383 475 384 476 
<< m2 >>
rect 383 475 384 476 
<< m1 >>
rect 384 475 385 476 
<< m1 >>
rect 385 475 386 476 
<< m1 >>
rect 386 475 387 476 
<< m1 >>
rect 387 475 388 476 
<< m1 >>
rect 388 475 389 476 
<< m1 >>
rect 389 475 390 476 
<< m1 >>
rect 390 475 391 476 
<< m2 >>
rect 390 475 391 476 
<< m1 >>
rect 391 475 392 476 
<< m1 >>
rect 392 475 393 476 
<< m1 >>
rect 393 475 394 476 
<< m1 >>
rect 394 475 395 476 
<< m1 >>
rect 433 475 434 476 
<< m1 >>
rect 451 475 452 476 
<< m1 >>
rect 472 475 473 476 
<< m1 >>
rect 487 475 488 476 
<< m1 >>
rect 489 475 490 476 
<< m1 >>
rect 21 476 22 477 
<< m1 >>
rect 28 476 29 477 
<< m1 >>
rect 49 476 50 477 
<< m1 >>
rect 70 476 71 477 
<< m1 >>
rect 73 476 74 477 
<< m1 >>
rect 85 476 86 477 
<< m1 >>
rect 121 476 122 477 
<< m1 >>
rect 135 476 136 477 
<< m1 >>
rect 142 476 143 477 
<< m1 >>
rect 172 476 173 477 
<< m2 >>
rect 178 476 179 477 
<< m1 >>
rect 208 476 209 477 
<< m1 >>
rect 253 476 254 477 
<< m1 >>
rect 255 476 256 477 
<< m1 >>
rect 271 476 272 477 
<< m1 >>
rect 286 476 287 477 
<< m2 >>
rect 302 476 303 477 
<< m1 >>
rect 307 476 308 477 
<< m2 >>
rect 352 476 353 477 
<< m2 >>
rect 356 476 357 477 
<< m1 >>
rect 379 476 380 477 
<< m1 >>
rect 381 476 382 477 
<< m2 >>
rect 390 476 391 477 
<< m1 >>
rect 433 476 434 477 
<< m1 >>
rect 451 476 452 477 
<< m1 >>
rect 472 476 473 477 
<< m1 >>
rect 487 476 488 477 
<< m1 >>
rect 489 476 490 477 
<< m1 >>
rect 21 477 22 478 
<< m1 >>
rect 28 477 29 478 
<< m1 >>
rect 49 477 50 478 
<< m1 >>
rect 70 477 71 478 
<< m1 >>
rect 73 477 74 478 
<< m1 >>
rect 85 477 86 478 
<< m1 >>
rect 121 477 122 478 
<< m1 >>
rect 135 477 136 478 
<< m1 >>
rect 142 477 143 478 
<< m1 >>
rect 172 477 173 478 
<< m1 >>
rect 175 477 176 478 
<< m1 >>
rect 176 477 177 478 
<< m1 >>
rect 177 477 178 478 
<< m1 >>
rect 178 477 179 478 
<< m2 >>
rect 178 477 179 478 
<< m1 >>
rect 179 477 180 478 
<< m1 >>
rect 180 477 181 478 
<< m1 >>
rect 181 477 182 478 
<< m1 >>
rect 208 477 209 478 
<< m1 >>
rect 247 477 248 478 
<< m1 >>
rect 248 477 249 478 
<< m1 >>
rect 249 477 250 478 
<< m1 >>
rect 250 477 251 478 
<< m1 >>
rect 251 477 252 478 
<< m2 >>
rect 251 477 252 478 
<< m2c >>
rect 251 477 252 478 
<< m1 >>
rect 251 477 252 478 
<< m2 >>
rect 251 477 252 478 
<< m2 >>
rect 252 477 253 478 
<< m1 >>
rect 253 477 254 478 
<< m2 >>
rect 253 477 254 478 
<< m2 >>
rect 254 477 255 478 
<< m1 >>
rect 255 477 256 478 
<< m2 >>
rect 255 477 256 478 
<< m2c >>
rect 255 477 256 478 
<< m1 >>
rect 255 477 256 478 
<< m2 >>
rect 255 477 256 478 
<< m1 >>
rect 271 477 272 478 
<< m1 >>
rect 286 477 287 478 
<< m1 >>
rect 302 477 303 478 
<< m2 >>
rect 302 477 303 478 
<< m2c >>
rect 302 477 303 478 
<< m1 >>
rect 302 477 303 478 
<< m2 >>
rect 302 477 303 478 
<< m1 >>
rect 303 477 304 478 
<< m1 >>
rect 304 477 305 478 
<< m1 >>
rect 307 477 308 478 
<< m1 >>
rect 337 477 338 478 
<< m1 >>
rect 338 477 339 478 
<< m1 >>
rect 339 477 340 478 
<< m1 >>
rect 340 477 341 478 
<< m1 >>
rect 341 477 342 478 
<< m1 >>
rect 342 477 343 478 
<< m1 >>
rect 343 477 344 478 
<< m1 >>
rect 344 477 345 478 
<< m1 >>
rect 345 477 346 478 
<< m1 >>
rect 346 477 347 478 
<< m1 >>
rect 347 477 348 478 
<< m1 >>
rect 348 477 349 478 
<< m1 >>
rect 349 477 350 478 
<< m1 >>
rect 350 477 351 478 
<< m1 >>
rect 351 477 352 478 
<< m1 >>
rect 352 477 353 478 
<< m2 >>
rect 352 477 353 478 
<< m2c >>
rect 352 477 353 478 
<< m1 >>
rect 352 477 353 478 
<< m2 >>
rect 352 477 353 478 
<< m1 >>
rect 356 477 357 478 
<< m2 >>
rect 356 477 357 478 
<< m2c >>
rect 356 477 357 478 
<< m1 >>
rect 356 477 357 478 
<< m2 >>
rect 356 477 357 478 
<< m1 >>
rect 357 477 358 478 
<< m1 >>
rect 358 477 359 478 
<< m1 >>
rect 359 477 360 478 
<< m1 >>
rect 360 477 361 478 
<< m1 >>
rect 361 477 362 478 
<< m1 >>
rect 379 477 380 478 
<< m1 >>
rect 381 477 382 478 
<< m2 >>
rect 382 477 383 478 
<< m1 >>
rect 383 477 384 478 
<< m2 >>
rect 383 477 384 478 
<< m2c >>
rect 383 477 384 478 
<< m1 >>
rect 383 477 384 478 
<< m2 >>
rect 383 477 384 478 
<< m1 >>
rect 384 477 385 478 
<< m1 >>
rect 385 477 386 478 
<< m1 >>
rect 386 477 387 478 
<< m1 >>
rect 387 477 388 478 
<< m1 >>
rect 388 477 389 478 
<< m1 >>
rect 389 477 390 478 
<< m1 >>
rect 390 477 391 478 
<< m2 >>
rect 390 477 391 478 
<< m2c >>
rect 390 477 391 478 
<< m1 >>
rect 390 477 391 478 
<< m2 >>
rect 390 477 391 478 
<< m1 >>
rect 433 477 434 478 
<< m1 >>
rect 451 477 452 478 
<< m1 >>
rect 472 477 473 478 
<< m1 >>
rect 487 477 488 478 
<< m1 >>
rect 489 477 490 478 
<< m1 >>
rect 21 478 22 479 
<< m1 >>
rect 28 478 29 479 
<< m1 >>
rect 49 478 50 479 
<< m1 >>
rect 70 478 71 479 
<< m1 >>
rect 73 478 74 479 
<< m1 >>
rect 85 478 86 479 
<< m1 >>
rect 121 478 122 479 
<< m1 >>
rect 135 478 136 479 
<< m1 >>
rect 142 478 143 479 
<< m1 >>
rect 172 478 173 479 
<< m1 >>
rect 175 478 176 479 
<< m2 >>
rect 178 478 179 479 
<< m1 >>
rect 181 478 182 479 
<< m1 >>
rect 208 478 209 479 
<< m1 >>
rect 247 478 248 479 
<< m1 >>
rect 253 478 254 479 
<< m1 >>
rect 271 478 272 479 
<< m1 >>
rect 286 478 287 479 
<< m1 >>
rect 304 478 305 479 
<< m1 >>
rect 307 478 308 479 
<< m1 >>
rect 337 478 338 479 
<< m1 >>
rect 361 478 362 479 
<< m1 >>
rect 379 478 380 479 
<< m1 >>
rect 381 478 382 479 
<< m2 >>
rect 382 478 383 479 
<< m1 >>
rect 394 478 395 479 
<< m1 >>
rect 395 478 396 479 
<< m1 >>
rect 396 478 397 479 
<< m1 >>
rect 397 478 398 479 
<< m1 >>
rect 398 478 399 479 
<< m1 >>
rect 399 478 400 479 
<< m1 >>
rect 400 478 401 479 
<< m1 >>
rect 401 478 402 479 
<< m1 >>
rect 402 478 403 479 
<< m1 >>
rect 403 478 404 479 
<< m1 >>
rect 404 478 405 479 
<< m1 >>
rect 405 478 406 479 
<< m1 >>
rect 406 478 407 479 
<< m1 >>
rect 433 478 434 479 
<< m1 >>
rect 451 478 452 479 
<< m1 >>
rect 472 478 473 479 
<< m1 >>
rect 484 478 485 479 
<< m1 >>
rect 485 478 486 479 
<< m2 >>
rect 485 478 486 479 
<< m2c >>
rect 485 478 486 479 
<< m1 >>
rect 485 478 486 479 
<< m2 >>
rect 485 478 486 479 
<< m2 >>
rect 486 478 487 479 
<< m1 >>
rect 487 478 488 479 
<< m2 >>
rect 487 478 488 479 
<< m2 >>
rect 488 478 489 479 
<< m1 >>
rect 489 478 490 479 
<< m2 >>
rect 489 478 490 479 
<< m2 >>
rect 490 478 491 479 
<< m1 >>
rect 491 478 492 479 
<< m2 >>
rect 491 478 492 479 
<< m2c >>
rect 491 478 492 479 
<< m1 >>
rect 491 478 492 479 
<< m2 >>
rect 491 478 492 479 
<< m1 >>
rect 492 478 493 479 
<< m1 >>
rect 493 478 494 479 
<< m1 >>
rect 494 478 495 479 
<< m1 >>
rect 495 478 496 479 
<< m1 >>
rect 496 478 497 479 
<< m1 >>
rect 497 478 498 479 
<< m1 >>
rect 498 478 499 479 
<< m1 >>
rect 499 478 500 479 
<< m1 >>
rect 21 479 22 480 
<< m1 >>
rect 28 479 29 480 
<< m1 >>
rect 49 479 50 480 
<< m1 >>
rect 70 479 71 480 
<< m1 >>
rect 73 479 74 480 
<< m1 >>
rect 85 479 86 480 
<< m1 >>
rect 121 479 122 480 
<< m1 >>
rect 135 479 136 480 
<< m1 >>
rect 142 479 143 480 
<< m1 >>
rect 172 479 173 480 
<< m1 >>
rect 175 479 176 480 
<< m1 >>
rect 178 479 179 480 
<< m2 >>
rect 178 479 179 480 
<< m1 >>
rect 181 479 182 480 
<< m1 >>
rect 208 479 209 480 
<< m1 >>
rect 247 479 248 480 
<< m1 >>
rect 253 479 254 480 
<< m1 >>
rect 271 479 272 480 
<< m1 >>
rect 286 479 287 480 
<< m1 >>
rect 304 479 305 480 
<< m1 >>
rect 307 479 308 480 
<< m1 >>
rect 337 479 338 480 
<< m1 >>
rect 361 479 362 480 
<< m1 >>
rect 379 479 380 480 
<< m1 >>
rect 381 479 382 480 
<< m2 >>
rect 382 479 383 480 
<< m1 >>
rect 394 479 395 480 
<< m1 >>
rect 406 479 407 480 
<< m1 >>
rect 433 479 434 480 
<< m1 >>
rect 451 479 452 480 
<< m1 >>
rect 472 479 473 480 
<< m1 >>
rect 484 479 485 480 
<< m1 >>
rect 487 479 488 480 
<< m1 >>
rect 489 479 490 480 
<< m1 >>
rect 499 479 500 480 
<< pdiffusion >>
rect 12 480 13 481 
<< pdiffusion >>
rect 13 480 14 481 
<< pdiffusion >>
rect 14 480 15 481 
<< pdiffusion >>
rect 15 480 16 481 
<< pdiffusion >>
rect 16 480 17 481 
<< pdiffusion >>
rect 17 480 18 481 
<< m1 >>
rect 21 480 22 481 
<< m1 >>
rect 28 480 29 481 
<< pdiffusion >>
rect 30 480 31 481 
<< pdiffusion >>
rect 31 480 32 481 
<< pdiffusion >>
rect 32 480 33 481 
<< pdiffusion >>
rect 33 480 34 481 
<< pdiffusion >>
rect 34 480 35 481 
<< pdiffusion >>
rect 35 480 36 481 
<< pdiffusion >>
rect 48 480 49 481 
<< m1 >>
rect 49 480 50 481 
<< pdiffusion >>
rect 49 480 50 481 
<< pdiffusion >>
rect 50 480 51 481 
<< pdiffusion >>
rect 51 480 52 481 
<< pdiffusion >>
rect 52 480 53 481 
<< pdiffusion >>
rect 53 480 54 481 
<< pdiffusion >>
rect 66 480 67 481 
<< pdiffusion >>
rect 67 480 68 481 
<< pdiffusion >>
rect 68 480 69 481 
<< pdiffusion >>
rect 69 480 70 481 
<< m1 >>
rect 70 480 71 481 
<< pdiffusion >>
rect 70 480 71 481 
<< pdiffusion >>
rect 71 480 72 481 
<< m1 >>
rect 73 480 74 481 
<< pdiffusion >>
rect 84 480 85 481 
<< m1 >>
rect 85 480 86 481 
<< pdiffusion >>
rect 85 480 86 481 
<< pdiffusion >>
rect 86 480 87 481 
<< pdiffusion >>
rect 87 480 88 481 
<< pdiffusion >>
rect 88 480 89 481 
<< pdiffusion >>
rect 89 480 90 481 
<< pdiffusion >>
rect 102 480 103 481 
<< pdiffusion >>
rect 103 480 104 481 
<< pdiffusion >>
rect 104 480 105 481 
<< pdiffusion >>
rect 105 480 106 481 
<< pdiffusion >>
rect 106 480 107 481 
<< pdiffusion >>
rect 107 480 108 481 
<< pdiffusion >>
rect 120 480 121 481 
<< m1 >>
rect 121 480 122 481 
<< pdiffusion >>
rect 121 480 122 481 
<< pdiffusion >>
rect 122 480 123 481 
<< pdiffusion >>
rect 123 480 124 481 
<< pdiffusion >>
rect 124 480 125 481 
<< pdiffusion >>
rect 125 480 126 481 
<< m1 >>
rect 135 480 136 481 
<< pdiffusion >>
rect 138 480 139 481 
<< pdiffusion >>
rect 139 480 140 481 
<< pdiffusion >>
rect 140 480 141 481 
<< pdiffusion >>
rect 141 480 142 481 
<< m1 >>
rect 142 480 143 481 
<< pdiffusion >>
rect 142 480 143 481 
<< pdiffusion >>
rect 143 480 144 481 
<< pdiffusion >>
rect 156 480 157 481 
<< pdiffusion >>
rect 157 480 158 481 
<< pdiffusion >>
rect 158 480 159 481 
<< pdiffusion >>
rect 159 480 160 481 
<< pdiffusion >>
rect 160 480 161 481 
<< pdiffusion >>
rect 161 480 162 481 
<< m1 >>
rect 172 480 173 481 
<< pdiffusion >>
rect 174 480 175 481 
<< m1 >>
rect 175 480 176 481 
<< pdiffusion >>
rect 175 480 176 481 
<< pdiffusion >>
rect 176 480 177 481 
<< m1 >>
rect 177 480 178 481 
<< m2 >>
rect 177 480 178 481 
<< m2c >>
rect 177 480 178 481 
<< m1 >>
rect 177 480 178 481 
<< m2 >>
rect 177 480 178 481 
<< pdiffusion >>
rect 177 480 178 481 
<< m1 >>
rect 178 480 179 481 
<< pdiffusion >>
rect 178 480 179 481 
<< pdiffusion >>
rect 179 480 180 481 
<< m1 >>
rect 181 480 182 481 
<< pdiffusion >>
rect 192 480 193 481 
<< pdiffusion >>
rect 193 480 194 481 
<< pdiffusion >>
rect 194 480 195 481 
<< pdiffusion >>
rect 195 480 196 481 
<< pdiffusion >>
rect 196 480 197 481 
<< pdiffusion >>
rect 197 480 198 481 
<< m1 >>
rect 208 480 209 481 
<< pdiffusion >>
rect 210 480 211 481 
<< pdiffusion >>
rect 211 480 212 481 
<< pdiffusion >>
rect 212 480 213 481 
<< pdiffusion >>
rect 213 480 214 481 
<< pdiffusion >>
rect 214 480 215 481 
<< pdiffusion >>
rect 215 480 216 481 
<< pdiffusion >>
rect 228 480 229 481 
<< pdiffusion >>
rect 229 480 230 481 
<< pdiffusion >>
rect 230 480 231 481 
<< pdiffusion >>
rect 231 480 232 481 
<< pdiffusion >>
rect 232 480 233 481 
<< pdiffusion >>
rect 233 480 234 481 
<< pdiffusion >>
rect 246 480 247 481 
<< m1 >>
rect 247 480 248 481 
<< pdiffusion >>
rect 247 480 248 481 
<< pdiffusion >>
rect 248 480 249 481 
<< pdiffusion >>
rect 249 480 250 481 
<< pdiffusion >>
rect 250 480 251 481 
<< pdiffusion >>
rect 251 480 252 481 
<< m1 >>
rect 253 480 254 481 
<< pdiffusion >>
rect 264 480 265 481 
<< pdiffusion >>
rect 265 480 266 481 
<< pdiffusion >>
rect 266 480 267 481 
<< pdiffusion >>
rect 267 480 268 481 
<< pdiffusion >>
rect 268 480 269 481 
<< pdiffusion >>
rect 269 480 270 481 
<< m1 >>
rect 271 480 272 481 
<< pdiffusion >>
rect 282 480 283 481 
<< pdiffusion >>
rect 283 480 284 481 
<< pdiffusion >>
rect 284 480 285 481 
<< pdiffusion >>
rect 285 480 286 481 
<< m1 >>
rect 286 480 287 481 
<< pdiffusion >>
rect 286 480 287 481 
<< pdiffusion >>
rect 287 480 288 481 
<< pdiffusion >>
rect 300 480 301 481 
<< pdiffusion >>
rect 301 480 302 481 
<< pdiffusion >>
rect 302 480 303 481 
<< pdiffusion >>
rect 303 480 304 481 
<< m1 >>
rect 304 480 305 481 
<< pdiffusion >>
rect 304 480 305 481 
<< pdiffusion >>
rect 305 480 306 481 
<< m1 >>
rect 307 480 308 481 
<< pdiffusion >>
rect 318 480 319 481 
<< pdiffusion >>
rect 319 480 320 481 
<< pdiffusion >>
rect 320 480 321 481 
<< pdiffusion >>
rect 321 480 322 481 
<< pdiffusion >>
rect 322 480 323 481 
<< pdiffusion >>
rect 323 480 324 481 
<< pdiffusion >>
rect 336 480 337 481 
<< m1 >>
rect 337 480 338 481 
<< pdiffusion >>
rect 337 480 338 481 
<< pdiffusion >>
rect 338 480 339 481 
<< pdiffusion >>
rect 339 480 340 481 
<< pdiffusion >>
rect 340 480 341 481 
<< pdiffusion >>
rect 341 480 342 481 
<< pdiffusion >>
rect 354 480 355 481 
<< pdiffusion >>
rect 355 480 356 481 
<< pdiffusion >>
rect 356 480 357 481 
<< pdiffusion >>
rect 357 480 358 481 
<< pdiffusion >>
rect 358 480 359 481 
<< pdiffusion >>
rect 359 480 360 481 
<< m1 >>
rect 361 480 362 481 
<< pdiffusion >>
rect 372 480 373 481 
<< pdiffusion >>
rect 373 480 374 481 
<< pdiffusion >>
rect 374 480 375 481 
<< pdiffusion >>
rect 375 480 376 481 
<< pdiffusion >>
rect 376 480 377 481 
<< pdiffusion >>
rect 377 480 378 481 
<< m1 >>
rect 379 480 380 481 
<< m1 >>
rect 381 480 382 481 
<< m2 >>
rect 382 480 383 481 
<< pdiffusion >>
rect 390 480 391 481 
<< pdiffusion >>
rect 391 480 392 481 
<< pdiffusion >>
rect 392 480 393 481 
<< pdiffusion >>
rect 393 480 394 481 
<< m1 >>
rect 394 480 395 481 
<< pdiffusion >>
rect 394 480 395 481 
<< pdiffusion >>
rect 395 480 396 481 
<< m1 >>
rect 406 480 407 481 
<< pdiffusion >>
rect 408 480 409 481 
<< pdiffusion >>
rect 409 480 410 481 
<< pdiffusion >>
rect 410 480 411 481 
<< pdiffusion >>
rect 411 480 412 481 
<< pdiffusion >>
rect 412 480 413 481 
<< pdiffusion >>
rect 413 480 414 481 
<< pdiffusion >>
rect 426 480 427 481 
<< pdiffusion >>
rect 427 480 428 481 
<< pdiffusion >>
rect 428 480 429 481 
<< pdiffusion >>
rect 429 480 430 481 
<< pdiffusion >>
rect 430 480 431 481 
<< pdiffusion >>
rect 431 480 432 481 
<< m1 >>
rect 433 480 434 481 
<< pdiffusion >>
rect 444 480 445 481 
<< pdiffusion >>
rect 445 480 446 481 
<< pdiffusion >>
rect 446 480 447 481 
<< pdiffusion >>
rect 447 480 448 481 
<< pdiffusion >>
rect 448 480 449 481 
<< pdiffusion >>
rect 449 480 450 481 
<< m1 >>
rect 451 480 452 481 
<< pdiffusion >>
rect 462 480 463 481 
<< pdiffusion >>
rect 463 480 464 481 
<< pdiffusion >>
rect 464 480 465 481 
<< pdiffusion >>
rect 465 480 466 481 
<< pdiffusion >>
rect 466 480 467 481 
<< pdiffusion >>
rect 467 480 468 481 
<< m1 >>
rect 472 480 473 481 
<< pdiffusion >>
rect 480 480 481 481 
<< pdiffusion >>
rect 481 480 482 481 
<< pdiffusion >>
rect 482 480 483 481 
<< pdiffusion >>
rect 483 480 484 481 
<< m1 >>
rect 484 480 485 481 
<< pdiffusion >>
rect 484 480 485 481 
<< pdiffusion >>
rect 485 480 486 481 
<< m1 >>
rect 487 480 488 481 
<< m1 >>
rect 489 480 490 481 
<< pdiffusion >>
rect 498 480 499 481 
<< m1 >>
rect 499 480 500 481 
<< pdiffusion >>
rect 499 480 500 481 
<< pdiffusion >>
rect 500 480 501 481 
<< pdiffusion >>
rect 501 480 502 481 
<< pdiffusion >>
rect 502 480 503 481 
<< pdiffusion >>
rect 503 480 504 481 
<< pdiffusion >>
rect 516 480 517 481 
<< pdiffusion >>
rect 517 480 518 481 
<< pdiffusion >>
rect 518 480 519 481 
<< pdiffusion >>
rect 519 480 520 481 
<< pdiffusion >>
rect 520 480 521 481 
<< pdiffusion >>
rect 521 480 522 481 
<< pdiffusion >>
rect 12 481 13 482 
<< pdiffusion >>
rect 13 481 14 482 
<< pdiffusion >>
rect 14 481 15 482 
<< pdiffusion >>
rect 15 481 16 482 
<< pdiffusion >>
rect 16 481 17 482 
<< pdiffusion >>
rect 17 481 18 482 
<< m1 >>
rect 21 481 22 482 
<< m1 >>
rect 28 481 29 482 
<< pdiffusion >>
rect 30 481 31 482 
<< pdiffusion >>
rect 31 481 32 482 
<< pdiffusion >>
rect 32 481 33 482 
<< pdiffusion >>
rect 33 481 34 482 
<< pdiffusion >>
rect 34 481 35 482 
<< pdiffusion >>
rect 35 481 36 482 
<< pdiffusion >>
rect 48 481 49 482 
<< pdiffusion >>
rect 49 481 50 482 
<< pdiffusion >>
rect 50 481 51 482 
<< pdiffusion >>
rect 51 481 52 482 
<< pdiffusion >>
rect 52 481 53 482 
<< pdiffusion >>
rect 53 481 54 482 
<< pdiffusion >>
rect 66 481 67 482 
<< pdiffusion >>
rect 67 481 68 482 
<< pdiffusion >>
rect 68 481 69 482 
<< pdiffusion >>
rect 69 481 70 482 
<< pdiffusion >>
rect 70 481 71 482 
<< pdiffusion >>
rect 71 481 72 482 
<< m1 >>
rect 73 481 74 482 
<< pdiffusion >>
rect 84 481 85 482 
<< pdiffusion >>
rect 85 481 86 482 
<< pdiffusion >>
rect 86 481 87 482 
<< pdiffusion >>
rect 87 481 88 482 
<< pdiffusion >>
rect 88 481 89 482 
<< pdiffusion >>
rect 89 481 90 482 
<< pdiffusion >>
rect 102 481 103 482 
<< pdiffusion >>
rect 103 481 104 482 
<< pdiffusion >>
rect 104 481 105 482 
<< pdiffusion >>
rect 105 481 106 482 
<< pdiffusion >>
rect 106 481 107 482 
<< pdiffusion >>
rect 107 481 108 482 
<< pdiffusion >>
rect 120 481 121 482 
<< pdiffusion >>
rect 121 481 122 482 
<< pdiffusion >>
rect 122 481 123 482 
<< pdiffusion >>
rect 123 481 124 482 
<< pdiffusion >>
rect 124 481 125 482 
<< pdiffusion >>
rect 125 481 126 482 
<< m1 >>
rect 135 481 136 482 
<< pdiffusion >>
rect 138 481 139 482 
<< pdiffusion >>
rect 139 481 140 482 
<< pdiffusion >>
rect 140 481 141 482 
<< pdiffusion >>
rect 141 481 142 482 
<< pdiffusion >>
rect 142 481 143 482 
<< pdiffusion >>
rect 143 481 144 482 
<< pdiffusion >>
rect 156 481 157 482 
<< pdiffusion >>
rect 157 481 158 482 
<< pdiffusion >>
rect 158 481 159 482 
<< pdiffusion >>
rect 159 481 160 482 
<< pdiffusion >>
rect 160 481 161 482 
<< pdiffusion >>
rect 161 481 162 482 
<< m1 >>
rect 172 481 173 482 
<< pdiffusion >>
rect 174 481 175 482 
<< pdiffusion >>
rect 175 481 176 482 
<< pdiffusion >>
rect 176 481 177 482 
<< pdiffusion >>
rect 177 481 178 482 
<< pdiffusion >>
rect 178 481 179 482 
<< pdiffusion >>
rect 179 481 180 482 
<< m1 >>
rect 181 481 182 482 
<< pdiffusion >>
rect 192 481 193 482 
<< pdiffusion >>
rect 193 481 194 482 
<< pdiffusion >>
rect 194 481 195 482 
<< pdiffusion >>
rect 195 481 196 482 
<< pdiffusion >>
rect 196 481 197 482 
<< pdiffusion >>
rect 197 481 198 482 
<< m1 >>
rect 208 481 209 482 
<< pdiffusion >>
rect 210 481 211 482 
<< pdiffusion >>
rect 211 481 212 482 
<< pdiffusion >>
rect 212 481 213 482 
<< pdiffusion >>
rect 213 481 214 482 
<< pdiffusion >>
rect 214 481 215 482 
<< pdiffusion >>
rect 215 481 216 482 
<< pdiffusion >>
rect 228 481 229 482 
<< pdiffusion >>
rect 229 481 230 482 
<< pdiffusion >>
rect 230 481 231 482 
<< pdiffusion >>
rect 231 481 232 482 
<< pdiffusion >>
rect 232 481 233 482 
<< pdiffusion >>
rect 233 481 234 482 
<< pdiffusion >>
rect 246 481 247 482 
<< pdiffusion >>
rect 247 481 248 482 
<< pdiffusion >>
rect 248 481 249 482 
<< pdiffusion >>
rect 249 481 250 482 
<< pdiffusion >>
rect 250 481 251 482 
<< pdiffusion >>
rect 251 481 252 482 
<< m1 >>
rect 253 481 254 482 
<< pdiffusion >>
rect 264 481 265 482 
<< pdiffusion >>
rect 265 481 266 482 
<< pdiffusion >>
rect 266 481 267 482 
<< pdiffusion >>
rect 267 481 268 482 
<< pdiffusion >>
rect 268 481 269 482 
<< pdiffusion >>
rect 269 481 270 482 
<< m1 >>
rect 271 481 272 482 
<< pdiffusion >>
rect 282 481 283 482 
<< pdiffusion >>
rect 283 481 284 482 
<< pdiffusion >>
rect 284 481 285 482 
<< pdiffusion >>
rect 285 481 286 482 
<< pdiffusion >>
rect 286 481 287 482 
<< pdiffusion >>
rect 287 481 288 482 
<< pdiffusion >>
rect 300 481 301 482 
<< pdiffusion >>
rect 301 481 302 482 
<< pdiffusion >>
rect 302 481 303 482 
<< pdiffusion >>
rect 303 481 304 482 
<< pdiffusion >>
rect 304 481 305 482 
<< pdiffusion >>
rect 305 481 306 482 
<< m1 >>
rect 307 481 308 482 
<< pdiffusion >>
rect 318 481 319 482 
<< pdiffusion >>
rect 319 481 320 482 
<< pdiffusion >>
rect 320 481 321 482 
<< pdiffusion >>
rect 321 481 322 482 
<< pdiffusion >>
rect 322 481 323 482 
<< pdiffusion >>
rect 323 481 324 482 
<< pdiffusion >>
rect 336 481 337 482 
<< pdiffusion >>
rect 337 481 338 482 
<< pdiffusion >>
rect 338 481 339 482 
<< pdiffusion >>
rect 339 481 340 482 
<< pdiffusion >>
rect 340 481 341 482 
<< pdiffusion >>
rect 341 481 342 482 
<< pdiffusion >>
rect 354 481 355 482 
<< pdiffusion >>
rect 355 481 356 482 
<< pdiffusion >>
rect 356 481 357 482 
<< pdiffusion >>
rect 357 481 358 482 
<< pdiffusion >>
rect 358 481 359 482 
<< pdiffusion >>
rect 359 481 360 482 
<< m1 >>
rect 361 481 362 482 
<< pdiffusion >>
rect 372 481 373 482 
<< pdiffusion >>
rect 373 481 374 482 
<< pdiffusion >>
rect 374 481 375 482 
<< pdiffusion >>
rect 375 481 376 482 
<< pdiffusion >>
rect 376 481 377 482 
<< pdiffusion >>
rect 377 481 378 482 
<< m1 >>
rect 379 481 380 482 
<< m1 >>
rect 381 481 382 482 
<< m2 >>
rect 382 481 383 482 
<< pdiffusion >>
rect 390 481 391 482 
<< pdiffusion >>
rect 391 481 392 482 
<< pdiffusion >>
rect 392 481 393 482 
<< pdiffusion >>
rect 393 481 394 482 
<< pdiffusion >>
rect 394 481 395 482 
<< pdiffusion >>
rect 395 481 396 482 
<< m1 >>
rect 406 481 407 482 
<< pdiffusion >>
rect 408 481 409 482 
<< pdiffusion >>
rect 409 481 410 482 
<< pdiffusion >>
rect 410 481 411 482 
<< pdiffusion >>
rect 411 481 412 482 
<< pdiffusion >>
rect 412 481 413 482 
<< pdiffusion >>
rect 413 481 414 482 
<< pdiffusion >>
rect 426 481 427 482 
<< pdiffusion >>
rect 427 481 428 482 
<< pdiffusion >>
rect 428 481 429 482 
<< pdiffusion >>
rect 429 481 430 482 
<< pdiffusion >>
rect 430 481 431 482 
<< pdiffusion >>
rect 431 481 432 482 
<< m1 >>
rect 433 481 434 482 
<< pdiffusion >>
rect 444 481 445 482 
<< pdiffusion >>
rect 445 481 446 482 
<< pdiffusion >>
rect 446 481 447 482 
<< pdiffusion >>
rect 447 481 448 482 
<< pdiffusion >>
rect 448 481 449 482 
<< pdiffusion >>
rect 449 481 450 482 
<< m1 >>
rect 451 481 452 482 
<< pdiffusion >>
rect 462 481 463 482 
<< pdiffusion >>
rect 463 481 464 482 
<< pdiffusion >>
rect 464 481 465 482 
<< pdiffusion >>
rect 465 481 466 482 
<< pdiffusion >>
rect 466 481 467 482 
<< pdiffusion >>
rect 467 481 468 482 
<< m1 >>
rect 472 481 473 482 
<< pdiffusion >>
rect 480 481 481 482 
<< pdiffusion >>
rect 481 481 482 482 
<< pdiffusion >>
rect 482 481 483 482 
<< pdiffusion >>
rect 483 481 484 482 
<< pdiffusion >>
rect 484 481 485 482 
<< pdiffusion >>
rect 485 481 486 482 
<< m1 >>
rect 487 481 488 482 
<< m1 >>
rect 489 481 490 482 
<< pdiffusion >>
rect 498 481 499 482 
<< pdiffusion >>
rect 499 481 500 482 
<< pdiffusion >>
rect 500 481 501 482 
<< pdiffusion >>
rect 501 481 502 482 
<< pdiffusion >>
rect 502 481 503 482 
<< pdiffusion >>
rect 503 481 504 482 
<< pdiffusion >>
rect 516 481 517 482 
<< pdiffusion >>
rect 517 481 518 482 
<< pdiffusion >>
rect 518 481 519 482 
<< pdiffusion >>
rect 519 481 520 482 
<< pdiffusion >>
rect 520 481 521 482 
<< pdiffusion >>
rect 521 481 522 482 
<< pdiffusion >>
rect 12 482 13 483 
<< pdiffusion >>
rect 13 482 14 483 
<< pdiffusion >>
rect 14 482 15 483 
<< pdiffusion >>
rect 15 482 16 483 
<< pdiffusion >>
rect 16 482 17 483 
<< pdiffusion >>
rect 17 482 18 483 
<< m1 >>
rect 21 482 22 483 
<< m1 >>
rect 28 482 29 483 
<< pdiffusion >>
rect 30 482 31 483 
<< pdiffusion >>
rect 31 482 32 483 
<< pdiffusion >>
rect 32 482 33 483 
<< pdiffusion >>
rect 33 482 34 483 
<< pdiffusion >>
rect 34 482 35 483 
<< pdiffusion >>
rect 35 482 36 483 
<< pdiffusion >>
rect 48 482 49 483 
<< pdiffusion >>
rect 49 482 50 483 
<< pdiffusion >>
rect 50 482 51 483 
<< pdiffusion >>
rect 51 482 52 483 
<< pdiffusion >>
rect 52 482 53 483 
<< pdiffusion >>
rect 53 482 54 483 
<< pdiffusion >>
rect 66 482 67 483 
<< pdiffusion >>
rect 67 482 68 483 
<< pdiffusion >>
rect 68 482 69 483 
<< pdiffusion >>
rect 69 482 70 483 
<< pdiffusion >>
rect 70 482 71 483 
<< pdiffusion >>
rect 71 482 72 483 
<< m1 >>
rect 73 482 74 483 
<< pdiffusion >>
rect 84 482 85 483 
<< pdiffusion >>
rect 85 482 86 483 
<< pdiffusion >>
rect 86 482 87 483 
<< pdiffusion >>
rect 87 482 88 483 
<< pdiffusion >>
rect 88 482 89 483 
<< pdiffusion >>
rect 89 482 90 483 
<< pdiffusion >>
rect 102 482 103 483 
<< pdiffusion >>
rect 103 482 104 483 
<< pdiffusion >>
rect 104 482 105 483 
<< pdiffusion >>
rect 105 482 106 483 
<< pdiffusion >>
rect 106 482 107 483 
<< pdiffusion >>
rect 107 482 108 483 
<< pdiffusion >>
rect 120 482 121 483 
<< pdiffusion >>
rect 121 482 122 483 
<< pdiffusion >>
rect 122 482 123 483 
<< pdiffusion >>
rect 123 482 124 483 
<< pdiffusion >>
rect 124 482 125 483 
<< pdiffusion >>
rect 125 482 126 483 
<< m1 >>
rect 135 482 136 483 
<< pdiffusion >>
rect 138 482 139 483 
<< pdiffusion >>
rect 139 482 140 483 
<< pdiffusion >>
rect 140 482 141 483 
<< pdiffusion >>
rect 141 482 142 483 
<< pdiffusion >>
rect 142 482 143 483 
<< pdiffusion >>
rect 143 482 144 483 
<< pdiffusion >>
rect 156 482 157 483 
<< pdiffusion >>
rect 157 482 158 483 
<< pdiffusion >>
rect 158 482 159 483 
<< pdiffusion >>
rect 159 482 160 483 
<< pdiffusion >>
rect 160 482 161 483 
<< pdiffusion >>
rect 161 482 162 483 
<< m1 >>
rect 172 482 173 483 
<< pdiffusion >>
rect 174 482 175 483 
<< pdiffusion >>
rect 175 482 176 483 
<< pdiffusion >>
rect 176 482 177 483 
<< pdiffusion >>
rect 177 482 178 483 
<< pdiffusion >>
rect 178 482 179 483 
<< pdiffusion >>
rect 179 482 180 483 
<< m1 >>
rect 181 482 182 483 
<< pdiffusion >>
rect 192 482 193 483 
<< pdiffusion >>
rect 193 482 194 483 
<< pdiffusion >>
rect 194 482 195 483 
<< pdiffusion >>
rect 195 482 196 483 
<< pdiffusion >>
rect 196 482 197 483 
<< pdiffusion >>
rect 197 482 198 483 
<< m1 >>
rect 208 482 209 483 
<< pdiffusion >>
rect 210 482 211 483 
<< pdiffusion >>
rect 211 482 212 483 
<< pdiffusion >>
rect 212 482 213 483 
<< pdiffusion >>
rect 213 482 214 483 
<< pdiffusion >>
rect 214 482 215 483 
<< pdiffusion >>
rect 215 482 216 483 
<< pdiffusion >>
rect 228 482 229 483 
<< pdiffusion >>
rect 229 482 230 483 
<< pdiffusion >>
rect 230 482 231 483 
<< pdiffusion >>
rect 231 482 232 483 
<< pdiffusion >>
rect 232 482 233 483 
<< pdiffusion >>
rect 233 482 234 483 
<< pdiffusion >>
rect 246 482 247 483 
<< pdiffusion >>
rect 247 482 248 483 
<< pdiffusion >>
rect 248 482 249 483 
<< pdiffusion >>
rect 249 482 250 483 
<< pdiffusion >>
rect 250 482 251 483 
<< pdiffusion >>
rect 251 482 252 483 
<< m1 >>
rect 253 482 254 483 
<< pdiffusion >>
rect 264 482 265 483 
<< pdiffusion >>
rect 265 482 266 483 
<< pdiffusion >>
rect 266 482 267 483 
<< pdiffusion >>
rect 267 482 268 483 
<< pdiffusion >>
rect 268 482 269 483 
<< pdiffusion >>
rect 269 482 270 483 
<< m1 >>
rect 271 482 272 483 
<< pdiffusion >>
rect 282 482 283 483 
<< pdiffusion >>
rect 283 482 284 483 
<< pdiffusion >>
rect 284 482 285 483 
<< pdiffusion >>
rect 285 482 286 483 
<< pdiffusion >>
rect 286 482 287 483 
<< pdiffusion >>
rect 287 482 288 483 
<< pdiffusion >>
rect 300 482 301 483 
<< pdiffusion >>
rect 301 482 302 483 
<< pdiffusion >>
rect 302 482 303 483 
<< pdiffusion >>
rect 303 482 304 483 
<< pdiffusion >>
rect 304 482 305 483 
<< pdiffusion >>
rect 305 482 306 483 
<< m1 >>
rect 307 482 308 483 
<< pdiffusion >>
rect 318 482 319 483 
<< pdiffusion >>
rect 319 482 320 483 
<< pdiffusion >>
rect 320 482 321 483 
<< pdiffusion >>
rect 321 482 322 483 
<< pdiffusion >>
rect 322 482 323 483 
<< pdiffusion >>
rect 323 482 324 483 
<< pdiffusion >>
rect 336 482 337 483 
<< pdiffusion >>
rect 337 482 338 483 
<< pdiffusion >>
rect 338 482 339 483 
<< pdiffusion >>
rect 339 482 340 483 
<< pdiffusion >>
rect 340 482 341 483 
<< pdiffusion >>
rect 341 482 342 483 
<< pdiffusion >>
rect 354 482 355 483 
<< pdiffusion >>
rect 355 482 356 483 
<< pdiffusion >>
rect 356 482 357 483 
<< pdiffusion >>
rect 357 482 358 483 
<< pdiffusion >>
rect 358 482 359 483 
<< pdiffusion >>
rect 359 482 360 483 
<< m1 >>
rect 361 482 362 483 
<< pdiffusion >>
rect 372 482 373 483 
<< pdiffusion >>
rect 373 482 374 483 
<< pdiffusion >>
rect 374 482 375 483 
<< pdiffusion >>
rect 375 482 376 483 
<< pdiffusion >>
rect 376 482 377 483 
<< pdiffusion >>
rect 377 482 378 483 
<< m1 >>
rect 379 482 380 483 
<< m1 >>
rect 381 482 382 483 
<< m2 >>
rect 382 482 383 483 
<< pdiffusion >>
rect 390 482 391 483 
<< pdiffusion >>
rect 391 482 392 483 
<< pdiffusion >>
rect 392 482 393 483 
<< pdiffusion >>
rect 393 482 394 483 
<< pdiffusion >>
rect 394 482 395 483 
<< pdiffusion >>
rect 395 482 396 483 
<< m1 >>
rect 406 482 407 483 
<< pdiffusion >>
rect 408 482 409 483 
<< pdiffusion >>
rect 409 482 410 483 
<< pdiffusion >>
rect 410 482 411 483 
<< pdiffusion >>
rect 411 482 412 483 
<< pdiffusion >>
rect 412 482 413 483 
<< pdiffusion >>
rect 413 482 414 483 
<< pdiffusion >>
rect 426 482 427 483 
<< pdiffusion >>
rect 427 482 428 483 
<< pdiffusion >>
rect 428 482 429 483 
<< pdiffusion >>
rect 429 482 430 483 
<< pdiffusion >>
rect 430 482 431 483 
<< pdiffusion >>
rect 431 482 432 483 
<< m1 >>
rect 433 482 434 483 
<< pdiffusion >>
rect 444 482 445 483 
<< pdiffusion >>
rect 445 482 446 483 
<< pdiffusion >>
rect 446 482 447 483 
<< pdiffusion >>
rect 447 482 448 483 
<< pdiffusion >>
rect 448 482 449 483 
<< pdiffusion >>
rect 449 482 450 483 
<< m1 >>
rect 451 482 452 483 
<< pdiffusion >>
rect 462 482 463 483 
<< pdiffusion >>
rect 463 482 464 483 
<< pdiffusion >>
rect 464 482 465 483 
<< pdiffusion >>
rect 465 482 466 483 
<< pdiffusion >>
rect 466 482 467 483 
<< pdiffusion >>
rect 467 482 468 483 
<< m1 >>
rect 472 482 473 483 
<< pdiffusion >>
rect 480 482 481 483 
<< pdiffusion >>
rect 481 482 482 483 
<< pdiffusion >>
rect 482 482 483 483 
<< pdiffusion >>
rect 483 482 484 483 
<< pdiffusion >>
rect 484 482 485 483 
<< pdiffusion >>
rect 485 482 486 483 
<< m1 >>
rect 487 482 488 483 
<< m1 >>
rect 489 482 490 483 
<< pdiffusion >>
rect 498 482 499 483 
<< pdiffusion >>
rect 499 482 500 483 
<< pdiffusion >>
rect 500 482 501 483 
<< pdiffusion >>
rect 501 482 502 483 
<< pdiffusion >>
rect 502 482 503 483 
<< pdiffusion >>
rect 503 482 504 483 
<< pdiffusion >>
rect 516 482 517 483 
<< pdiffusion >>
rect 517 482 518 483 
<< pdiffusion >>
rect 518 482 519 483 
<< pdiffusion >>
rect 519 482 520 483 
<< pdiffusion >>
rect 520 482 521 483 
<< pdiffusion >>
rect 521 482 522 483 
<< pdiffusion >>
rect 12 483 13 484 
<< pdiffusion >>
rect 13 483 14 484 
<< pdiffusion >>
rect 14 483 15 484 
<< pdiffusion >>
rect 15 483 16 484 
<< pdiffusion >>
rect 16 483 17 484 
<< pdiffusion >>
rect 17 483 18 484 
<< m1 >>
rect 21 483 22 484 
<< m1 >>
rect 28 483 29 484 
<< pdiffusion >>
rect 30 483 31 484 
<< pdiffusion >>
rect 31 483 32 484 
<< pdiffusion >>
rect 32 483 33 484 
<< pdiffusion >>
rect 33 483 34 484 
<< pdiffusion >>
rect 34 483 35 484 
<< pdiffusion >>
rect 35 483 36 484 
<< pdiffusion >>
rect 48 483 49 484 
<< pdiffusion >>
rect 49 483 50 484 
<< pdiffusion >>
rect 50 483 51 484 
<< pdiffusion >>
rect 51 483 52 484 
<< pdiffusion >>
rect 52 483 53 484 
<< pdiffusion >>
rect 53 483 54 484 
<< pdiffusion >>
rect 66 483 67 484 
<< pdiffusion >>
rect 67 483 68 484 
<< pdiffusion >>
rect 68 483 69 484 
<< pdiffusion >>
rect 69 483 70 484 
<< pdiffusion >>
rect 70 483 71 484 
<< pdiffusion >>
rect 71 483 72 484 
<< m1 >>
rect 73 483 74 484 
<< pdiffusion >>
rect 84 483 85 484 
<< pdiffusion >>
rect 85 483 86 484 
<< pdiffusion >>
rect 86 483 87 484 
<< pdiffusion >>
rect 87 483 88 484 
<< pdiffusion >>
rect 88 483 89 484 
<< pdiffusion >>
rect 89 483 90 484 
<< pdiffusion >>
rect 102 483 103 484 
<< pdiffusion >>
rect 103 483 104 484 
<< pdiffusion >>
rect 104 483 105 484 
<< pdiffusion >>
rect 105 483 106 484 
<< pdiffusion >>
rect 106 483 107 484 
<< pdiffusion >>
rect 107 483 108 484 
<< pdiffusion >>
rect 120 483 121 484 
<< pdiffusion >>
rect 121 483 122 484 
<< pdiffusion >>
rect 122 483 123 484 
<< pdiffusion >>
rect 123 483 124 484 
<< pdiffusion >>
rect 124 483 125 484 
<< pdiffusion >>
rect 125 483 126 484 
<< m1 >>
rect 135 483 136 484 
<< pdiffusion >>
rect 138 483 139 484 
<< pdiffusion >>
rect 139 483 140 484 
<< pdiffusion >>
rect 140 483 141 484 
<< pdiffusion >>
rect 141 483 142 484 
<< pdiffusion >>
rect 142 483 143 484 
<< pdiffusion >>
rect 143 483 144 484 
<< pdiffusion >>
rect 156 483 157 484 
<< pdiffusion >>
rect 157 483 158 484 
<< pdiffusion >>
rect 158 483 159 484 
<< pdiffusion >>
rect 159 483 160 484 
<< pdiffusion >>
rect 160 483 161 484 
<< pdiffusion >>
rect 161 483 162 484 
<< m1 >>
rect 172 483 173 484 
<< pdiffusion >>
rect 174 483 175 484 
<< pdiffusion >>
rect 175 483 176 484 
<< pdiffusion >>
rect 176 483 177 484 
<< pdiffusion >>
rect 177 483 178 484 
<< pdiffusion >>
rect 178 483 179 484 
<< pdiffusion >>
rect 179 483 180 484 
<< m1 >>
rect 181 483 182 484 
<< pdiffusion >>
rect 192 483 193 484 
<< pdiffusion >>
rect 193 483 194 484 
<< pdiffusion >>
rect 194 483 195 484 
<< pdiffusion >>
rect 195 483 196 484 
<< pdiffusion >>
rect 196 483 197 484 
<< pdiffusion >>
rect 197 483 198 484 
<< m1 >>
rect 208 483 209 484 
<< pdiffusion >>
rect 210 483 211 484 
<< pdiffusion >>
rect 211 483 212 484 
<< pdiffusion >>
rect 212 483 213 484 
<< pdiffusion >>
rect 213 483 214 484 
<< pdiffusion >>
rect 214 483 215 484 
<< pdiffusion >>
rect 215 483 216 484 
<< pdiffusion >>
rect 228 483 229 484 
<< pdiffusion >>
rect 229 483 230 484 
<< pdiffusion >>
rect 230 483 231 484 
<< pdiffusion >>
rect 231 483 232 484 
<< pdiffusion >>
rect 232 483 233 484 
<< pdiffusion >>
rect 233 483 234 484 
<< pdiffusion >>
rect 246 483 247 484 
<< pdiffusion >>
rect 247 483 248 484 
<< pdiffusion >>
rect 248 483 249 484 
<< pdiffusion >>
rect 249 483 250 484 
<< pdiffusion >>
rect 250 483 251 484 
<< pdiffusion >>
rect 251 483 252 484 
<< m1 >>
rect 253 483 254 484 
<< pdiffusion >>
rect 264 483 265 484 
<< pdiffusion >>
rect 265 483 266 484 
<< pdiffusion >>
rect 266 483 267 484 
<< pdiffusion >>
rect 267 483 268 484 
<< pdiffusion >>
rect 268 483 269 484 
<< pdiffusion >>
rect 269 483 270 484 
<< m1 >>
rect 271 483 272 484 
<< pdiffusion >>
rect 282 483 283 484 
<< pdiffusion >>
rect 283 483 284 484 
<< pdiffusion >>
rect 284 483 285 484 
<< pdiffusion >>
rect 285 483 286 484 
<< pdiffusion >>
rect 286 483 287 484 
<< pdiffusion >>
rect 287 483 288 484 
<< pdiffusion >>
rect 300 483 301 484 
<< pdiffusion >>
rect 301 483 302 484 
<< pdiffusion >>
rect 302 483 303 484 
<< pdiffusion >>
rect 303 483 304 484 
<< pdiffusion >>
rect 304 483 305 484 
<< pdiffusion >>
rect 305 483 306 484 
<< m1 >>
rect 307 483 308 484 
<< pdiffusion >>
rect 318 483 319 484 
<< pdiffusion >>
rect 319 483 320 484 
<< pdiffusion >>
rect 320 483 321 484 
<< pdiffusion >>
rect 321 483 322 484 
<< pdiffusion >>
rect 322 483 323 484 
<< pdiffusion >>
rect 323 483 324 484 
<< pdiffusion >>
rect 336 483 337 484 
<< pdiffusion >>
rect 337 483 338 484 
<< pdiffusion >>
rect 338 483 339 484 
<< pdiffusion >>
rect 339 483 340 484 
<< pdiffusion >>
rect 340 483 341 484 
<< pdiffusion >>
rect 341 483 342 484 
<< pdiffusion >>
rect 354 483 355 484 
<< pdiffusion >>
rect 355 483 356 484 
<< pdiffusion >>
rect 356 483 357 484 
<< pdiffusion >>
rect 357 483 358 484 
<< pdiffusion >>
rect 358 483 359 484 
<< pdiffusion >>
rect 359 483 360 484 
<< m1 >>
rect 361 483 362 484 
<< pdiffusion >>
rect 372 483 373 484 
<< pdiffusion >>
rect 373 483 374 484 
<< pdiffusion >>
rect 374 483 375 484 
<< pdiffusion >>
rect 375 483 376 484 
<< pdiffusion >>
rect 376 483 377 484 
<< pdiffusion >>
rect 377 483 378 484 
<< m1 >>
rect 379 483 380 484 
<< m1 >>
rect 381 483 382 484 
<< m2 >>
rect 382 483 383 484 
<< pdiffusion >>
rect 390 483 391 484 
<< pdiffusion >>
rect 391 483 392 484 
<< pdiffusion >>
rect 392 483 393 484 
<< pdiffusion >>
rect 393 483 394 484 
<< pdiffusion >>
rect 394 483 395 484 
<< pdiffusion >>
rect 395 483 396 484 
<< m1 >>
rect 406 483 407 484 
<< pdiffusion >>
rect 408 483 409 484 
<< pdiffusion >>
rect 409 483 410 484 
<< pdiffusion >>
rect 410 483 411 484 
<< pdiffusion >>
rect 411 483 412 484 
<< pdiffusion >>
rect 412 483 413 484 
<< pdiffusion >>
rect 413 483 414 484 
<< pdiffusion >>
rect 426 483 427 484 
<< pdiffusion >>
rect 427 483 428 484 
<< pdiffusion >>
rect 428 483 429 484 
<< pdiffusion >>
rect 429 483 430 484 
<< pdiffusion >>
rect 430 483 431 484 
<< pdiffusion >>
rect 431 483 432 484 
<< m1 >>
rect 433 483 434 484 
<< pdiffusion >>
rect 444 483 445 484 
<< pdiffusion >>
rect 445 483 446 484 
<< pdiffusion >>
rect 446 483 447 484 
<< pdiffusion >>
rect 447 483 448 484 
<< pdiffusion >>
rect 448 483 449 484 
<< pdiffusion >>
rect 449 483 450 484 
<< m1 >>
rect 451 483 452 484 
<< pdiffusion >>
rect 462 483 463 484 
<< pdiffusion >>
rect 463 483 464 484 
<< pdiffusion >>
rect 464 483 465 484 
<< pdiffusion >>
rect 465 483 466 484 
<< pdiffusion >>
rect 466 483 467 484 
<< pdiffusion >>
rect 467 483 468 484 
<< m1 >>
rect 472 483 473 484 
<< pdiffusion >>
rect 480 483 481 484 
<< pdiffusion >>
rect 481 483 482 484 
<< pdiffusion >>
rect 482 483 483 484 
<< pdiffusion >>
rect 483 483 484 484 
<< pdiffusion >>
rect 484 483 485 484 
<< pdiffusion >>
rect 485 483 486 484 
<< m1 >>
rect 487 483 488 484 
<< m1 >>
rect 489 483 490 484 
<< pdiffusion >>
rect 498 483 499 484 
<< pdiffusion >>
rect 499 483 500 484 
<< pdiffusion >>
rect 500 483 501 484 
<< pdiffusion >>
rect 501 483 502 484 
<< pdiffusion >>
rect 502 483 503 484 
<< pdiffusion >>
rect 503 483 504 484 
<< pdiffusion >>
rect 516 483 517 484 
<< pdiffusion >>
rect 517 483 518 484 
<< pdiffusion >>
rect 518 483 519 484 
<< pdiffusion >>
rect 519 483 520 484 
<< pdiffusion >>
rect 520 483 521 484 
<< pdiffusion >>
rect 521 483 522 484 
<< pdiffusion >>
rect 12 484 13 485 
<< pdiffusion >>
rect 13 484 14 485 
<< pdiffusion >>
rect 14 484 15 485 
<< pdiffusion >>
rect 15 484 16 485 
<< pdiffusion >>
rect 16 484 17 485 
<< pdiffusion >>
rect 17 484 18 485 
<< m1 >>
rect 21 484 22 485 
<< m1 >>
rect 28 484 29 485 
<< pdiffusion >>
rect 30 484 31 485 
<< pdiffusion >>
rect 31 484 32 485 
<< pdiffusion >>
rect 32 484 33 485 
<< pdiffusion >>
rect 33 484 34 485 
<< pdiffusion >>
rect 34 484 35 485 
<< pdiffusion >>
rect 35 484 36 485 
<< pdiffusion >>
rect 48 484 49 485 
<< pdiffusion >>
rect 49 484 50 485 
<< pdiffusion >>
rect 50 484 51 485 
<< pdiffusion >>
rect 51 484 52 485 
<< pdiffusion >>
rect 52 484 53 485 
<< pdiffusion >>
rect 53 484 54 485 
<< pdiffusion >>
rect 66 484 67 485 
<< pdiffusion >>
rect 67 484 68 485 
<< pdiffusion >>
rect 68 484 69 485 
<< pdiffusion >>
rect 69 484 70 485 
<< pdiffusion >>
rect 70 484 71 485 
<< pdiffusion >>
rect 71 484 72 485 
<< m1 >>
rect 73 484 74 485 
<< pdiffusion >>
rect 84 484 85 485 
<< pdiffusion >>
rect 85 484 86 485 
<< pdiffusion >>
rect 86 484 87 485 
<< pdiffusion >>
rect 87 484 88 485 
<< pdiffusion >>
rect 88 484 89 485 
<< pdiffusion >>
rect 89 484 90 485 
<< pdiffusion >>
rect 102 484 103 485 
<< pdiffusion >>
rect 103 484 104 485 
<< pdiffusion >>
rect 104 484 105 485 
<< pdiffusion >>
rect 105 484 106 485 
<< pdiffusion >>
rect 106 484 107 485 
<< pdiffusion >>
rect 107 484 108 485 
<< pdiffusion >>
rect 120 484 121 485 
<< pdiffusion >>
rect 121 484 122 485 
<< pdiffusion >>
rect 122 484 123 485 
<< pdiffusion >>
rect 123 484 124 485 
<< pdiffusion >>
rect 124 484 125 485 
<< pdiffusion >>
rect 125 484 126 485 
<< m1 >>
rect 135 484 136 485 
<< pdiffusion >>
rect 138 484 139 485 
<< pdiffusion >>
rect 139 484 140 485 
<< pdiffusion >>
rect 140 484 141 485 
<< pdiffusion >>
rect 141 484 142 485 
<< pdiffusion >>
rect 142 484 143 485 
<< pdiffusion >>
rect 143 484 144 485 
<< pdiffusion >>
rect 156 484 157 485 
<< pdiffusion >>
rect 157 484 158 485 
<< pdiffusion >>
rect 158 484 159 485 
<< pdiffusion >>
rect 159 484 160 485 
<< pdiffusion >>
rect 160 484 161 485 
<< pdiffusion >>
rect 161 484 162 485 
<< m1 >>
rect 172 484 173 485 
<< pdiffusion >>
rect 174 484 175 485 
<< pdiffusion >>
rect 175 484 176 485 
<< pdiffusion >>
rect 176 484 177 485 
<< pdiffusion >>
rect 177 484 178 485 
<< pdiffusion >>
rect 178 484 179 485 
<< pdiffusion >>
rect 179 484 180 485 
<< m1 >>
rect 181 484 182 485 
<< pdiffusion >>
rect 192 484 193 485 
<< pdiffusion >>
rect 193 484 194 485 
<< pdiffusion >>
rect 194 484 195 485 
<< pdiffusion >>
rect 195 484 196 485 
<< pdiffusion >>
rect 196 484 197 485 
<< pdiffusion >>
rect 197 484 198 485 
<< m1 >>
rect 208 484 209 485 
<< pdiffusion >>
rect 210 484 211 485 
<< pdiffusion >>
rect 211 484 212 485 
<< pdiffusion >>
rect 212 484 213 485 
<< pdiffusion >>
rect 213 484 214 485 
<< pdiffusion >>
rect 214 484 215 485 
<< pdiffusion >>
rect 215 484 216 485 
<< pdiffusion >>
rect 228 484 229 485 
<< pdiffusion >>
rect 229 484 230 485 
<< pdiffusion >>
rect 230 484 231 485 
<< pdiffusion >>
rect 231 484 232 485 
<< pdiffusion >>
rect 232 484 233 485 
<< pdiffusion >>
rect 233 484 234 485 
<< pdiffusion >>
rect 246 484 247 485 
<< pdiffusion >>
rect 247 484 248 485 
<< pdiffusion >>
rect 248 484 249 485 
<< pdiffusion >>
rect 249 484 250 485 
<< pdiffusion >>
rect 250 484 251 485 
<< pdiffusion >>
rect 251 484 252 485 
<< m1 >>
rect 253 484 254 485 
<< pdiffusion >>
rect 264 484 265 485 
<< pdiffusion >>
rect 265 484 266 485 
<< pdiffusion >>
rect 266 484 267 485 
<< pdiffusion >>
rect 267 484 268 485 
<< pdiffusion >>
rect 268 484 269 485 
<< pdiffusion >>
rect 269 484 270 485 
<< m1 >>
rect 271 484 272 485 
<< pdiffusion >>
rect 282 484 283 485 
<< pdiffusion >>
rect 283 484 284 485 
<< pdiffusion >>
rect 284 484 285 485 
<< pdiffusion >>
rect 285 484 286 485 
<< pdiffusion >>
rect 286 484 287 485 
<< pdiffusion >>
rect 287 484 288 485 
<< pdiffusion >>
rect 300 484 301 485 
<< pdiffusion >>
rect 301 484 302 485 
<< pdiffusion >>
rect 302 484 303 485 
<< pdiffusion >>
rect 303 484 304 485 
<< pdiffusion >>
rect 304 484 305 485 
<< pdiffusion >>
rect 305 484 306 485 
<< m1 >>
rect 307 484 308 485 
<< pdiffusion >>
rect 318 484 319 485 
<< pdiffusion >>
rect 319 484 320 485 
<< pdiffusion >>
rect 320 484 321 485 
<< pdiffusion >>
rect 321 484 322 485 
<< pdiffusion >>
rect 322 484 323 485 
<< pdiffusion >>
rect 323 484 324 485 
<< pdiffusion >>
rect 336 484 337 485 
<< pdiffusion >>
rect 337 484 338 485 
<< pdiffusion >>
rect 338 484 339 485 
<< pdiffusion >>
rect 339 484 340 485 
<< pdiffusion >>
rect 340 484 341 485 
<< pdiffusion >>
rect 341 484 342 485 
<< pdiffusion >>
rect 354 484 355 485 
<< pdiffusion >>
rect 355 484 356 485 
<< pdiffusion >>
rect 356 484 357 485 
<< pdiffusion >>
rect 357 484 358 485 
<< pdiffusion >>
rect 358 484 359 485 
<< pdiffusion >>
rect 359 484 360 485 
<< m1 >>
rect 361 484 362 485 
<< pdiffusion >>
rect 372 484 373 485 
<< pdiffusion >>
rect 373 484 374 485 
<< pdiffusion >>
rect 374 484 375 485 
<< pdiffusion >>
rect 375 484 376 485 
<< pdiffusion >>
rect 376 484 377 485 
<< pdiffusion >>
rect 377 484 378 485 
<< m1 >>
rect 379 484 380 485 
<< m1 >>
rect 381 484 382 485 
<< m2 >>
rect 382 484 383 485 
<< pdiffusion >>
rect 390 484 391 485 
<< pdiffusion >>
rect 391 484 392 485 
<< pdiffusion >>
rect 392 484 393 485 
<< pdiffusion >>
rect 393 484 394 485 
<< pdiffusion >>
rect 394 484 395 485 
<< pdiffusion >>
rect 395 484 396 485 
<< m1 >>
rect 406 484 407 485 
<< pdiffusion >>
rect 408 484 409 485 
<< pdiffusion >>
rect 409 484 410 485 
<< pdiffusion >>
rect 410 484 411 485 
<< pdiffusion >>
rect 411 484 412 485 
<< pdiffusion >>
rect 412 484 413 485 
<< pdiffusion >>
rect 413 484 414 485 
<< pdiffusion >>
rect 426 484 427 485 
<< pdiffusion >>
rect 427 484 428 485 
<< pdiffusion >>
rect 428 484 429 485 
<< pdiffusion >>
rect 429 484 430 485 
<< pdiffusion >>
rect 430 484 431 485 
<< pdiffusion >>
rect 431 484 432 485 
<< m1 >>
rect 433 484 434 485 
<< pdiffusion >>
rect 444 484 445 485 
<< pdiffusion >>
rect 445 484 446 485 
<< pdiffusion >>
rect 446 484 447 485 
<< pdiffusion >>
rect 447 484 448 485 
<< pdiffusion >>
rect 448 484 449 485 
<< pdiffusion >>
rect 449 484 450 485 
<< m1 >>
rect 451 484 452 485 
<< pdiffusion >>
rect 462 484 463 485 
<< pdiffusion >>
rect 463 484 464 485 
<< pdiffusion >>
rect 464 484 465 485 
<< pdiffusion >>
rect 465 484 466 485 
<< pdiffusion >>
rect 466 484 467 485 
<< pdiffusion >>
rect 467 484 468 485 
<< m1 >>
rect 472 484 473 485 
<< pdiffusion >>
rect 480 484 481 485 
<< pdiffusion >>
rect 481 484 482 485 
<< pdiffusion >>
rect 482 484 483 485 
<< pdiffusion >>
rect 483 484 484 485 
<< pdiffusion >>
rect 484 484 485 485 
<< pdiffusion >>
rect 485 484 486 485 
<< m1 >>
rect 487 484 488 485 
<< m1 >>
rect 489 484 490 485 
<< pdiffusion >>
rect 498 484 499 485 
<< pdiffusion >>
rect 499 484 500 485 
<< pdiffusion >>
rect 500 484 501 485 
<< pdiffusion >>
rect 501 484 502 485 
<< pdiffusion >>
rect 502 484 503 485 
<< pdiffusion >>
rect 503 484 504 485 
<< pdiffusion >>
rect 516 484 517 485 
<< pdiffusion >>
rect 517 484 518 485 
<< pdiffusion >>
rect 518 484 519 485 
<< pdiffusion >>
rect 519 484 520 485 
<< pdiffusion >>
rect 520 484 521 485 
<< pdiffusion >>
rect 521 484 522 485 
<< pdiffusion >>
rect 12 485 13 486 
<< pdiffusion >>
rect 13 485 14 486 
<< pdiffusion >>
rect 14 485 15 486 
<< pdiffusion >>
rect 15 485 16 486 
<< m1 >>
rect 16 485 17 486 
<< pdiffusion >>
rect 16 485 17 486 
<< pdiffusion >>
rect 17 485 18 486 
<< m1 >>
rect 21 485 22 486 
<< m1 >>
rect 28 485 29 486 
<< pdiffusion >>
rect 30 485 31 486 
<< pdiffusion >>
rect 31 485 32 486 
<< pdiffusion >>
rect 32 485 33 486 
<< pdiffusion >>
rect 33 485 34 486 
<< pdiffusion >>
rect 34 485 35 486 
<< pdiffusion >>
rect 35 485 36 486 
<< pdiffusion >>
rect 48 485 49 486 
<< pdiffusion >>
rect 49 485 50 486 
<< pdiffusion >>
rect 50 485 51 486 
<< pdiffusion >>
rect 51 485 52 486 
<< pdiffusion >>
rect 52 485 53 486 
<< pdiffusion >>
rect 53 485 54 486 
<< pdiffusion >>
rect 66 485 67 486 
<< pdiffusion >>
rect 67 485 68 486 
<< pdiffusion >>
rect 68 485 69 486 
<< pdiffusion >>
rect 69 485 70 486 
<< pdiffusion >>
rect 70 485 71 486 
<< pdiffusion >>
rect 71 485 72 486 
<< m1 >>
rect 73 485 74 486 
<< pdiffusion >>
rect 84 485 85 486 
<< pdiffusion >>
rect 85 485 86 486 
<< pdiffusion >>
rect 86 485 87 486 
<< pdiffusion >>
rect 87 485 88 486 
<< pdiffusion >>
rect 88 485 89 486 
<< pdiffusion >>
rect 89 485 90 486 
<< pdiffusion >>
rect 102 485 103 486 
<< pdiffusion >>
rect 103 485 104 486 
<< pdiffusion >>
rect 104 485 105 486 
<< pdiffusion >>
rect 105 485 106 486 
<< pdiffusion >>
rect 106 485 107 486 
<< pdiffusion >>
rect 107 485 108 486 
<< pdiffusion >>
rect 120 485 121 486 
<< pdiffusion >>
rect 121 485 122 486 
<< pdiffusion >>
rect 122 485 123 486 
<< pdiffusion >>
rect 123 485 124 486 
<< m1 >>
rect 124 485 125 486 
<< pdiffusion >>
rect 124 485 125 486 
<< pdiffusion >>
rect 125 485 126 486 
<< m1 >>
rect 135 485 136 486 
<< pdiffusion >>
rect 138 485 139 486 
<< pdiffusion >>
rect 139 485 140 486 
<< pdiffusion >>
rect 140 485 141 486 
<< pdiffusion >>
rect 141 485 142 486 
<< pdiffusion >>
rect 142 485 143 486 
<< pdiffusion >>
rect 143 485 144 486 
<< pdiffusion >>
rect 156 485 157 486 
<< m1 >>
rect 157 485 158 486 
<< pdiffusion >>
rect 157 485 158 486 
<< pdiffusion >>
rect 158 485 159 486 
<< pdiffusion >>
rect 159 485 160 486 
<< pdiffusion >>
rect 160 485 161 486 
<< pdiffusion >>
rect 161 485 162 486 
<< m1 >>
rect 172 485 173 486 
<< pdiffusion >>
rect 174 485 175 486 
<< pdiffusion >>
rect 175 485 176 486 
<< pdiffusion >>
rect 176 485 177 486 
<< pdiffusion >>
rect 177 485 178 486 
<< pdiffusion >>
rect 178 485 179 486 
<< pdiffusion >>
rect 179 485 180 486 
<< m1 >>
rect 181 485 182 486 
<< pdiffusion >>
rect 192 485 193 486 
<< pdiffusion >>
rect 193 485 194 486 
<< pdiffusion >>
rect 194 485 195 486 
<< pdiffusion >>
rect 195 485 196 486 
<< pdiffusion >>
rect 196 485 197 486 
<< pdiffusion >>
rect 197 485 198 486 
<< m1 >>
rect 208 485 209 486 
<< pdiffusion >>
rect 210 485 211 486 
<< pdiffusion >>
rect 211 485 212 486 
<< pdiffusion >>
rect 212 485 213 486 
<< pdiffusion >>
rect 213 485 214 486 
<< pdiffusion >>
rect 214 485 215 486 
<< pdiffusion >>
rect 215 485 216 486 
<< pdiffusion >>
rect 228 485 229 486 
<< pdiffusion >>
rect 229 485 230 486 
<< pdiffusion >>
rect 230 485 231 486 
<< pdiffusion >>
rect 231 485 232 486 
<< pdiffusion >>
rect 232 485 233 486 
<< pdiffusion >>
rect 233 485 234 486 
<< pdiffusion >>
rect 246 485 247 486 
<< pdiffusion >>
rect 247 485 248 486 
<< pdiffusion >>
rect 248 485 249 486 
<< pdiffusion >>
rect 249 485 250 486 
<< pdiffusion >>
rect 250 485 251 486 
<< pdiffusion >>
rect 251 485 252 486 
<< m1 >>
rect 253 485 254 486 
<< pdiffusion >>
rect 264 485 265 486 
<< pdiffusion >>
rect 265 485 266 486 
<< pdiffusion >>
rect 266 485 267 486 
<< pdiffusion >>
rect 267 485 268 486 
<< m1 >>
rect 268 485 269 486 
<< pdiffusion >>
rect 268 485 269 486 
<< pdiffusion >>
rect 269 485 270 486 
<< m1 >>
rect 271 485 272 486 
<< pdiffusion >>
rect 282 485 283 486 
<< pdiffusion >>
rect 283 485 284 486 
<< pdiffusion >>
rect 284 485 285 486 
<< pdiffusion >>
rect 285 485 286 486 
<< m1 >>
rect 286 485 287 486 
<< pdiffusion >>
rect 286 485 287 486 
<< pdiffusion >>
rect 287 485 288 486 
<< pdiffusion >>
rect 300 485 301 486 
<< pdiffusion >>
rect 301 485 302 486 
<< pdiffusion >>
rect 302 485 303 486 
<< pdiffusion >>
rect 303 485 304 486 
<< pdiffusion >>
rect 304 485 305 486 
<< pdiffusion >>
rect 305 485 306 486 
<< m1 >>
rect 307 485 308 486 
<< pdiffusion >>
rect 318 485 319 486 
<< pdiffusion >>
rect 319 485 320 486 
<< pdiffusion >>
rect 320 485 321 486 
<< pdiffusion >>
rect 321 485 322 486 
<< pdiffusion >>
rect 322 485 323 486 
<< pdiffusion >>
rect 323 485 324 486 
<< pdiffusion >>
rect 336 485 337 486 
<< pdiffusion >>
rect 337 485 338 486 
<< pdiffusion >>
rect 338 485 339 486 
<< pdiffusion >>
rect 339 485 340 486 
<< pdiffusion >>
rect 340 485 341 486 
<< pdiffusion >>
rect 341 485 342 486 
<< pdiffusion >>
rect 354 485 355 486 
<< pdiffusion >>
rect 355 485 356 486 
<< pdiffusion >>
rect 356 485 357 486 
<< pdiffusion >>
rect 357 485 358 486 
<< pdiffusion >>
rect 358 485 359 486 
<< pdiffusion >>
rect 359 485 360 486 
<< m1 >>
rect 361 485 362 486 
<< pdiffusion >>
rect 372 485 373 486 
<< pdiffusion >>
rect 373 485 374 486 
<< pdiffusion >>
rect 374 485 375 486 
<< pdiffusion >>
rect 375 485 376 486 
<< pdiffusion >>
rect 376 485 377 486 
<< pdiffusion >>
rect 377 485 378 486 
<< m1 >>
rect 379 485 380 486 
<< m1 >>
rect 381 485 382 486 
<< m2 >>
rect 382 485 383 486 
<< pdiffusion >>
rect 390 485 391 486 
<< pdiffusion >>
rect 391 485 392 486 
<< pdiffusion >>
rect 392 485 393 486 
<< pdiffusion >>
rect 393 485 394 486 
<< pdiffusion >>
rect 394 485 395 486 
<< pdiffusion >>
rect 395 485 396 486 
<< m1 >>
rect 406 485 407 486 
<< pdiffusion >>
rect 408 485 409 486 
<< pdiffusion >>
rect 409 485 410 486 
<< pdiffusion >>
rect 410 485 411 486 
<< pdiffusion >>
rect 411 485 412 486 
<< pdiffusion >>
rect 412 485 413 486 
<< pdiffusion >>
rect 413 485 414 486 
<< pdiffusion >>
rect 426 485 427 486 
<< pdiffusion >>
rect 427 485 428 486 
<< pdiffusion >>
rect 428 485 429 486 
<< pdiffusion >>
rect 429 485 430 486 
<< pdiffusion >>
rect 430 485 431 486 
<< pdiffusion >>
rect 431 485 432 486 
<< m1 >>
rect 433 485 434 486 
<< pdiffusion >>
rect 444 485 445 486 
<< pdiffusion >>
rect 445 485 446 486 
<< pdiffusion >>
rect 446 485 447 486 
<< pdiffusion >>
rect 447 485 448 486 
<< pdiffusion >>
rect 448 485 449 486 
<< pdiffusion >>
rect 449 485 450 486 
<< m1 >>
rect 451 485 452 486 
<< pdiffusion >>
rect 462 485 463 486 
<< pdiffusion >>
rect 463 485 464 486 
<< pdiffusion >>
rect 464 485 465 486 
<< pdiffusion >>
rect 465 485 466 486 
<< m1 >>
rect 466 485 467 486 
<< pdiffusion >>
rect 466 485 467 486 
<< pdiffusion >>
rect 467 485 468 486 
<< m1 >>
rect 472 485 473 486 
<< pdiffusion >>
rect 480 485 481 486 
<< pdiffusion >>
rect 481 485 482 486 
<< pdiffusion >>
rect 482 485 483 486 
<< pdiffusion >>
rect 483 485 484 486 
<< pdiffusion >>
rect 484 485 485 486 
<< pdiffusion >>
rect 485 485 486 486 
<< m1 >>
rect 487 485 488 486 
<< m1 >>
rect 489 485 490 486 
<< pdiffusion >>
rect 498 485 499 486 
<< pdiffusion >>
rect 499 485 500 486 
<< pdiffusion >>
rect 500 485 501 486 
<< pdiffusion >>
rect 501 485 502 486 
<< pdiffusion >>
rect 502 485 503 486 
<< pdiffusion >>
rect 503 485 504 486 
<< pdiffusion >>
rect 516 485 517 486 
<< pdiffusion >>
rect 517 485 518 486 
<< pdiffusion >>
rect 518 485 519 486 
<< pdiffusion >>
rect 519 485 520 486 
<< m1 >>
rect 520 485 521 486 
<< pdiffusion >>
rect 520 485 521 486 
<< pdiffusion >>
rect 521 485 522 486 
<< m1 >>
rect 16 486 17 487 
<< m1 >>
rect 21 486 22 487 
<< m1 >>
rect 28 486 29 487 
<< m1 >>
rect 73 486 74 487 
<< m1 >>
rect 124 486 125 487 
<< m1 >>
rect 135 486 136 487 
<< m1 >>
rect 157 486 158 487 
<< m1 >>
rect 172 486 173 487 
<< m1 >>
rect 181 486 182 487 
<< m1 >>
rect 208 486 209 487 
<< m1 >>
rect 253 486 254 487 
<< m1 >>
rect 268 486 269 487 
<< m1 >>
rect 271 486 272 487 
<< m1 >>
rect 286 486 287 487 
<< m1 >>
rect 307 486 308 487 
<< m1 >>
rect 361 486 362 487 
<< m1 >>
rect 379 486 380 487 
<< m1 >>
rect 381 486 382 487 
<< m2 >>
rect 382 486 383 487 
<< m1 >>
rect 406 486 407 487 
<< m1 >>
rect 433 486 434 487 
<< m1 >>
rect 451 486 452 487 
<< m1 >>
rect 466 486 467 487 
<< m1 >>
rect 472 486 473 487 
<< m1 >>
rect 487 486 488 487 
<< m1 >>
rect 489 486 490 487 
<< m1 >>
rect 520 486 521 487 
<< m1 >>
rect 16 487 17 488 
<< m1 >>
rect 17 487 18 488 
<< m1 >>
rect 18 487 19 488 
<< m1 >>
rect 19 487 20 488 
<< m1 >>
rect 20 487 21 488 
<< m1 >>
rect 21 487 22 488 
<< m1 >>
rect 28 487 29 488 
<< m1 >>
rect 73 487 74 488 
<< m1 >>
rect 124 487 125 488 
<< m1 >>
rect 125 487 126 488 
<< m1 >>
rect 126 487 127 488 
<< m1 >>
rect 127 487 128 488 
<< m1 >>
rect 128 487 129 488 
<< m1 >>
rect 129 487 130 488 
<< m1 >>
rect 130 487 131 488 
<< m1 >>
rect 131 487 132 488 
<< m1 >>
rect 132 487 133 488 
<< m1 >>
rect 133 487 134 488 
<< m1 >>
rect 134 487 135 488 
<< m1 >>
rect 135 487 136 488 
<< m1 >>
rect 157 487 158 488 
<< m1 >>
rect 172 487 173 488 
<< m1 >>
rect 181 487 182 488 
<< m1 >>
rect 208 487 209 488 
<< m1 >>
rect 253 487 254 488 
<< m1 >>
rect 268 487 269 488 
<< m1 >>
rect 269 487 270 488 
<< m1 >>
rect 270 487 271 488 
<< m1 >>
rect 271 487 272 488 
<< m1 >>
rect 286 487 287 488 
<< m1 >>
rect 307 487 308 488 
<< m1 >>
rect 361 487 362 488 
<< m1 >>
rect 379 487 380 488 
<< m1 >>
rect 381 487 382 488 
<< m2 >>
rect 382 487 383 488 
<< m1 >>
rect 406 487 407 488 
<< m1 >>
rect 433 487 434 488 
<< m1 >>
rect 451 487 452 488 
<< m1 >>
rect 466 487 467 488 
<< m1 >>
rect 472 487 473 488 
<< m1 >>
rect 487 487 488 488 
<< m1 >>
rect 489 487 490 488 
<< m1 >>
rect 520 487 521 488 
<< m1 >>
rect 521 487 522 488 
<< m1 >>
rect 522 487 523 488 
<< m1 >>
rect 523 487 524 488 
<< m1 >>
rect 28 488 29 489 
<< m1 >>
rect 73 488 74 489 
<< m1 >>
rect 157 488 158 489 
<< m1 >>
rect 158 488 159 489 
<< m1 >>
rect 159 488 160 489 
<< m1 >>
rect 160 488 161 489 
<< m1 >>
rect 161 488 162 489 
<< m1 >>
rect 162 488 163 489 
<< m1 >>
rect 163 488 164 489 
<< m1 >>
rect 164 488 165 489 
<< m1 >>
rect 165 488 166 489 
<< m1 >>
rect 166 488 167 489 
<< m1 >>
rect 167 488 168 489 
<< m1 >>
rect 168 488 169 489 
<< m1 >>
rect 169 488 170 489 
<< m1 >>
rect 170 488 171 489 
<< m1 >>
rect 171 488 172 489 
<< m1 >>
rect 172 488 173 489 
<< m1 >>
rect 181 488 182 489 
<< m1 >>
rect 208 488 209 489 
<< m1 >>
rect 209 488 210 489 
<< m1 >>
rect 210 488 211 489 
<< m2 >>
rect 210 488 211 489 
<< m2c >>
rect 210 488 211 489 
<< m1 >>
rect 210 488 211 489 
<< m2 >>
rect 210 488 211 489 
<< m1 >>
rect 253 488 254 489 
<< m2 >>
rect 253 488 254 489 
<< m2c >>
rect 253 488 254 489 
<< m1 >>
rect 253 488 254 489 
<< m2 >>
rect 253 488 254 489 
<< m1 >>
rect 286 488 287 489 
<< m1 >>
rect 307 488 308 489 
<< m1 >>
rect 361 488 362 489 
<< m2 >>
rect 361 488 362 489 
<< m2c >>
rect 361 488 362 489 
<< m1 >>
rect 361 488 362 489 
<< m2 >>
rect 361 488 362 489 
<< m1 >>
rect 379 488 380 489 
<< m1 >>
rect 381 488 382 489 
<< m2 >>
rect 382 488 383 489 
<< m1 >>
rect 406 488 407 489 
<< m1 >>
rect 433 488 434 489 
<< m1 >>
rect 451 488 452 489 
<< m2 >>
rect 451 488 452 489 
<< m2c >>
rect 451 488 452 489 
<< m1 >>
rect 451 488 452 489 
<< m2 >>
rect 451 488 452 489 
<< m1 >>
rect 466 488 467 489 
<< m1 >>
rect 472 488 473 489 
<< m1 >>
rect 487 488 488 489 
<< m1 >>
rect 489 488 490 489 
<< m1 >>
rect 523 488 524 489 
<< m1 >>
rect 28 489 29 490 
<< m1 >>
rect 73 489 74 490 
<< m1 >>
rect 181 489 182 490 
<< m2 >>
rect 210 489 211 490 
<< m2 >>
rect 253 489 254 490 
<< m1 >>
rect 286 489 287 490 
<< m1 >>
rect 307 489 308 490 
<< m2 >>
rect 361 489 362 490 
<< m1 >>
rect 379 489 380 490 
<< m1 >>
rect 381 489 382 490 
<< m2 >>
rect 382 489 383 490 
<< m1 >>
rect 406 489 407 490 
<< m1 >>
rect 433 489 434 490 
<< m2 >>
rect 451 489 452 490 
<< m1 >>
rect 466 489 467 490 
<< m1 >>
rect 472 489 473 490 
<< m1 >>
rect 487 489 488 490 
<< m1 >>
rect 489 489 490 490 
<< m1 >>
rect 523 489 524 490 
<< m1 >>
rect 28 490 29 491 
<< m1 >>
rect 73 490 74 491 
<< m1 >>
rect 181 490 182 491 
<< m1 >>
rect 182 490 183 491 
<< m1 >>
rect 183 490 184 491 
<< m1 >>
rect 184 490 185 491 
<< m1 >>
rect 185 490 186 491 
<< m1 >>
rect 186 490 187 491 
<< m1 >>
rect 187 490 188 491 
<< m1 >>
rect 188 490 189 491 
<< m1 >>
rect 189 490 190 491 
<< m1 >>
rect 190 490 191 491 
<< m1 >>
rect 191 490 192 491 
<< m1 >>
rect 192 490 193 491 
<< m1 >>
rect 193 490 194 491 
<< m1 >>
rect 194 490 195 491 
<< m1 >>
rect 195 490 196 491 
<< m1 >>
rect 196 490 197 491 
<< m1 >>
rect 197 490 198 491 
<< m1 >>
rect 198 490 199 491 
<< m1 >>
rect 199 490 200 491 
<< m1 >>
rect 200 490 201 491 
<< m1 >>
rect 201 490 202 491 
<< m1 >>
rect 202 490 203 491 
<< m1 >>
rect 203 490 204 491 
<< m1 >>
rect 204 490 205 491 
<< m1 >>
rect 205 490 206 491 
<< m1 >>
rect 206 490 207 491 
<< m1 >>
rect 207 490 208 491 
<< m1 >>
rect 208 490 209 491 
<< m1 >>
rect 209 490 210 491 
<< m1 >>
rect 210 490 211 491 
<< m2 >>
rect 210 490 211 491 
<< m1 >>
rect 211 490 212 491 
<< m2 >>
rect 211 490 212 491 
<< m2 >>
rect 212 490 213 491 
<< m1 >>
rect 213 490 214 491 
<< m2 >>
rect 213 490 214 491 
<< m2c >>
rect 213 490 214 491 
<< m1 >>
rect 213 490 214 491 
<< m2 >>
rect 213 490 214 491 
<< m1 >>
rect 214 490 215 491 
<< m1 >>
rect 215 490 216 491 
<< m1 >>
rect 216 490 217 491 
<< m1 >>
rect 217 490 218 491 
<< m1 >>
rect 218 490 219 491 
<< m1 >>
rect 219 490 220 491 
<< m1 >>
rect 220 490 221 491 
<< m1 >>
rect 221 490 222 491 
<< m1 >>
rect 222 490 223 491 
<< m1 >>
rect 223 490 224 491 
<< m1 >>
rect 224 490 225 491 
<< m1 >>
rect 225 490 226 491 
<< m1 >>
rect 226 490 227 491 
<< m1 >>
rect 227 490 228 491 
<< m1 >>
rect 228 490 229 491 
<< m1 >>
rect 229 490 230 491 
<< m1 >>
rect 230 490 231 491 
<< m1 >>
rect 231 490 232 491 
<< m1 >>
rect 232 490 233 491 
<< m1 >>
rect 233 490 234 491 
<< m1 >>
rect 234 490 235 491 
<< m1 >>
rect 235 490 236 491 
<< m1 >>
rect 236 490 237 491 
<< m1 >>
rect 237 490 238 491 
<< m1 >>
rect 238 490 239 491 
<< m1 >>
rect 239 490 240 491 
<< m1 >>
rect 240 490 241 491 
<< m1 >>
rect 241 490 242 491 
<< m1 >>
rect 242 490 243 491 
<< m1 >>
rect 243 490 244 491 
<< m1 >>
rect 244 490 245 491 
<< m1 >>
rect 245 490 246 491 
<< m1 >>
rect 246 490 247 491 
<< m1 >>
rect 247 490 248 491 
<< m1 >>
rect 248 490 249 491 
<< m1 >>
rect 249 490 250 491 
<< m1 >>
rect 250 490 251 491 
<< m1 >>
rect 251 490 252 491 
<< m1 >>
rect 252 490 253 491 
<< m1 >>
rect 253 490 254 491 
<< m2 >>
rect 253 490 254 491 
<< m1 >>
rect 254 490 255 491 
<< m1 >>
rect 255 490 256 491 
<< m1 >>
rect 256 490 257 491 
<< m1 >>
rect 257 490 258 491 
<< m1 >>
rect 258 490 259 491 
<< m1 >>
rect 259 490 260 491 
<< m1 >>
rect 260 490 261 491 
<< m1 >>
rect 261 490 262 491 
<< m1 >>
rect 262 490 263 491 
<< m1 >>
rect 263 490 264 491 
<< m1 >>
rect 264 490 265 491 
<< m1 >>
rect 265 490 266 491 
<< m1 >>
rect 266 490 267 491 
<< m1 >>
rect 267 490 268 491 
<< m1 >>
rect 268 490 269 491 
<< m1 >>
rect 269 490 270 491 
<< m1 >>
rect 270 490 271 491 
<< m1 >>
rect 271 490 272 491 
<< m1 >>
rect 272 490 273 491 
<< m1 >>
rect 273 490 274 491 
<< m1 >>
rect 274 490 275 491 
<< m1 >>
rect 275 490 276 491 
<< m1 >>
rect 276 490 277 491 
<< m1 >>
rect 277 490 278 491 
<< m1 >>
rect 278 490 279 491 
<< m1 >>
rect 279 490 280 491 
<< m1 >>
rect 280 490 281 491 
<< m1 >>
rect 281 490 282 491 
<< m1 >>
rect 282 490 283 491 
<< m1 >>
rect 283 490 284 491 
<< m1 >>
rect 284 490 285 491 
<< m1 >>
rect 285 490 286 491 
<< m1 >>
rect 286 490 287 491 
<< m1 >>
rect 307 490 308 491 
<< m1 >>
rect 308 490 309 491 
<< m1 >>
rect 309 490 310 491 
<< m1 >>
rect 310 490 311 491 
<< m1 >>
rect 311 490 312 491 
<< m1 >>
rect 312 490 313 491 
<< m1 >>
rect 313 490 314 491 
<< m1 >>
rect 314 490 315 491 
<< m1 >>
rect 315 490 316 491 
<< m1 >>
rect 316 490 317 491 
<< m1 >>
rect 317 490 318 491 
<< m1 >>
rect 318 490 319 491 
<< m1 >>
rect 319 490 320 491 
<< m1 >>
rect 320 490 321 491 
<< m1 >>
rect 321 490 322 491 
<< m1 >>
rect 322 490 323 491 
<< m1 >>
rect 323 490 324 491 
<< m1 >>
rect 324 490 325 491 
<< m1 >>
rect 325 490 326 491 
<< m1 >>
rect 326 490 327 491 
<< m1 >>
rect 327 490 328 491 
<< m1 >>
rect 328 490 329 491 
<< m1 >>
rect 329 490 330 491 
<< m1 >>
rect 330 490 331 491 
<< m1 >>
rect 331 490 332 491 
<< m1 >>
rect 332 490 333 491 
<< m1 >>
rect 333 490 334 491 
<< m1 >>
rect 334 490 335 491 
<< m1 >>
rect 335 490 336 491 
<< m1 >>
rect 336 490 337 491 
<< m1 >>
rect 337 490 338 491 
<< m1 >>
rect 338 490 339 491 
<< m1 >>
rect 339 490 340 491 
<< m1 >>
rect 340 490 341 491 
<< m1 >>
rect 341 490 342 491 
<< m1 >>
rect 342 490 343 491 
<< m1 >>
rect 343 490 344 491 
<< m1 >>
rect 344 490 345 491 
<< m1 >>
rect 345 490 346 491 
<< m1 >>
rect 346 490 347 491 
<< m1 >>
rect 347 490 348 491 
<< m1 >>
rect 348 490 349 491 
<< m1 >>
rect 349 490 350 491 
<< m1 >>
rect 350 490 351 491 
<< m1 >>
rect 351 490 352 491 
<< m1 >>
rect 352 490 353 491 
<< m1 >>
rect 353 490 354 491 
<< m1 >>
rect 354 490 355 491 
<< m1 >>
rect 355 490 356 491 
<< m1 >>
rect 356 490 357 491 
<< m1 >>
rect 357 490 358 491 
<< m1 >>
rect 358 490 359 491 
<< m1 >>
rect 359 490 360 491 
<< m1 >>
rect 360 490 361 491 
<< m1 >>
rect 361 490 362 491 
<< m2 >>
rect 361 490 362 491 
<< m1 >>
rect 362 490 363 491 
<< m1 >>
rect 363 490 364 491 
<< m1 >>
rect 364 490 365 491 
<< m1 >>
rect 365 490 366 491 
<< m1 >>
rect 366 490 367 491 
<< m1 >>
rect 367 490 368 491 
<< m1 >>
rect 368 490 369 491 
<< m1 >>
rect 369 490 370 491 
<< m1 >>
rect 370 490 371 491 
<< m1 >>
rect 371 490 372 491 
<< m1 >>
rect 372 490 373 491 
<< m1 >>
rect 373 490 374 491 
<< m1 >>
rect 379 490 380 491 
<< m1 >>
rect 381 490 382 491 
<< m2 >>
rect 382 490 383 491 
<< m1 >>
rect 406 490 407 491 
<< m1 >>
rect 433 490 434 491 
<< m1 >>
rect 434 490 435 491 
<< m1 >>
rect 435 490 436 491 
<< m1 >>
rect 436 490 437 491 
<< m1 >>
rect 437 490 438 491 
<< m1 >>
rect 438 490 439 491 
<< m1 >>
rect 439 490 440 491 
<< m1 >>
rect 440 490 441 491 
<< m1 >>
rect 441 490 442 491 
<< m1 >>
rect 442 490 443 491 
<< m1 >>
rect 443 490 444 491 
<< m1 >>
rect 444 490 445 491 
<< m1 >>
rect 445 490 446 491 
<< m1 >>
rect 446 490 447 491 
<< m1 >>
rect 447 490 448 491 
<< m1 >>
rect 448 490 449 491 
<< m1 >>
rect 449 490 450 491 
<< m1 >>
rect 450 490 451 491 
<< m1 >>
rect 451 490 452 491 
<< m2 >>
rect 451 490 452 491 
<< m1 >>
rect 452 490 453 491 
<< m1 >>
rect 453 490 454 491 
<< m1 >>
rect 454 490 455 491 
<< m1 >>
rect 455 490 456 491 
<< m1 >>
rect 456 490 457 491 
<< m1 >>
rect 457 490 458 491 
<< m1 >>
rect 458 490 459 491 
<< m1 >>
rect 459 490 460 491 
<< m1 >>
rect 460 490 461 491 
<< m1 >>
rect 461 490 462 491 
<< m1 >>
rect 462 490 463 491 
<< m1 >>
rect 463 490 464 491 
<< m1 >>
rect 464 490 465 491 
<< m1 >>
rect 465 490 466 491 
<< m1 >>
rect 466 490 467 491 
<< m1 >>
rect 472 490 473 491 
<< m1 >>
rect 487 490 488 491 
<< m1 >>
rect 489 490 490 491 
<< m1 >>
rect 523 490 524 491 
<< m1 >>
rect 28 491 29 492 
<< m1 >>
rect 73 491 74 492 
<< m1 >>
rect 211 491 212 492 
<< m2 >>
rect 253 491 254 492 
<< m2 >>
rect 361 491 362 492 
<< m1 >>
rect 373 491 374 492 
<< m1 >>
rect 379 491 380 492 
<< m1 >>
rect 381 491 382 492 
<< m2 >>
rect 382 491 383 492 
<< m1 >>
rect 406 491 407 492 
<< m2 >>
rect 451 491 452 492 
<< m1 >>
rect 472 491 473 492 
<< m1 >>
rect 487 491 488 492 
<< m1 >>
rect 489 491 490 492 
<< m1 >>
rect 523 491 524 492 
<< m1 >>
rect 28 492 29 493 
<< m1 >>
rect 73 492 74 493 
<< m1 >>
rect 211 492 212 493 
<< m1 >>
rect 253 492 254 493 
<< m2 >>
rect 253 492 254 493 
<< m2c >>
rect 253 492 254 493 
<< m1 >>
rect 253 492 254 493 
<< m2 >>
rect 253 492 254 493 
<< m1 >>
rect 361 492 362 493 
<< m2 >>
rect 361 492 362 493 
<< m2c >>
rect 361 492 362 493 
<< m1 >>
rect 361 492 362 493 
<< m2 >>
rect 361 492 362 493 
<< m1 >>
rect 373 492 374 493 
<< m1 >>
rect 379 492 380 493 
<< m1 >>
rect 381 492 382 493 
<< m2 >>
rect 382 492 383 493 
<< m1 >>
rect 406 492 407 493 
<< m1 >>
rect 451 492 452 493 
<< m2 >>
rect 451 492 452 493 
<< m2c >>
rect 451 492 452 493 
<< m1 >>
rect 451 492 452 493 
<< m2 >>
rect 451 492 452 493 
<< m1 >>
rect 472 492 473 493 
<< m1 >>
rect 487 492 488 493 
<< m1 >>
rect 489 492 490 493 
<< m1 >>
rect 523 492 524 493 
<< m1 >>
rect 28 493 29 494 
<< m1 >>
rect 73 493 74 494 
<< m1 >>
rect 211 493 212 494 
<< m1 >>
rect 253 493 254 494 
<< m1 >>
rect 361 493 362 494 
<< m1 >>
rect 373 493 374 494 
<< m1 >>
rect 379 493 380 494 
<< m1 >>
rect 381 493 382 494 
<< m2 >>
rect 382 493 383 494 
<< m1 >>
rect 406 493 407 494 
<< m1 >>
rect 451 493 452 494 
<< m1 >>
rect 472 493 473 494 
<< m1 >>
rect 487 493 488 494 
<< m1 >>
rect 489 493 490 494 
<< m1 >>
rect 523 493 524 494 
<< m1 >>
rect 28 494 29 495 
<< m1 >>
rect 73 494 74 495 
<< m1 >>
rect 211 494 212 495 
<< m1 >>
rect 253 494 254 495 
<< m1 >>
rect 361 494 362 495 
<< m1 >>
rect 373 494 374 495 
<< m1 >>
rect 379 494 380 495 
<< m1 >>
rect 381 494 382 495 
<< m2 >>
rect 382 494 383 495 
<< m1 >>
rect 406 494 407 495 
<< m1 >>
rect 451 494 452 495 
<< m1 >>
rect 472 494 473 495 
<< m1 >>
rect 487 494 488 495 
<< m1 >>
rect 489 494 490 495 
<< m1 >>
rect 523 494 524 495 
<< m1 >>
rect 28 495 29 496 
<< m1 >>
rect 73 495 74 496 
<< m1 >>
rect 103 495 104 496 
<< m1 >>
rect 104 495 105 496 
<< m1 >>
rect 105 495 106 496 
<< m1 >>
rect 106 495 107 496 
<< m1 >>
rect 107 495 108 496 
<< m1 >>
rect 108 495 109 496 
<< m1 >>
rect 109 495 110 496 
<< m1 >>
rect 110 495 111 496 
<< m1 >>
rect 111 495 112 496 
<< m1 >>
rect 112 495 113 496 
<< m1 >>
rect 113 495 114 496 
<< m1 >>
rect 114 495 115 496 
<< m1 >>
rect 115 495 116 496 
<< m1 >>
rect 116 495 117 496 
<< m1 >>
rect 117 495 118 496 
<< m1 >>
rect 118 495 119 496 
<< m1 >>
rect 175 495 176 496 
<< m1 >>
rect 176 495 177 496 
<< m1 >>
rect 177 495 178 496 
<< m1 >>
rect 178 495 179 496 
<< m1 >>
rect 179 495 180 496 
<< m1 >>
rect 180 495 181 496 
<< m1 >>
rect 181 495 182 496 
<< m1 >>
rect 182 495 183 496 
<< m1 >>
rect 183 495 184 496 
<< m1 >>
rect 184 495 185 496 
<< m1 >>
rect 185 495 186 496 
<< m1 >>
rect 186 495 187 496 
<< m1 >>
rect 187 495 188 496 
<< m1 >>
rect 188 495 189 496 
<< m1 >>
rect 189 495 190 496 
<< m1 >>
rect 190 495 191 496 
<< m1 >>
rect 211 495 212 496 
<< m1 >>
rect 253 495 254 496 
<< m1 >>
rect 361 495 362 496 
<< m1 >>
rect 373 495 374 496 
<< m1 >>
rect 379 495 380 496 
<< m1 >>
rect 381 495 382 496 
<< m2 >>
rect 382 495 383 496 
<< m1 >>
rect 406 495 407 496 
<< m1 >>
rect 451 495 452 496 
<< m1 >>
rect 472 495 473 496 
<< m1 >>
rect 487 495 488 496 
<< m1 >>
rect 489 495 490 496 
<< m1 >>
rect 523 495 524 496 
<< m1 >>
rect 28 496 29 497 
<< m1 >>
rect 34 496 35 497 
<< m1 >>
rect 35 496 36 497 
<< m1 >>
rect 36 496 37 497 
<< m1 >>
rect 37 496 38 497 
<< m1 >>
rect 73 496 74 497 
<< m1 >>
rect 88 496 89 497 
<< m1 >>
rect 89 496 90 497 
<< m1 >>
rect 90 496 91 497 
<< m1 >>
rect 91 496 92 497 
<< m1 >>
rect 92 496 93 497 
<< m1 >>
rect 93 496 94 497 
<< m1 >>
rect 94 496 95 497 
<< m1 >>
rect 95 496 96 497 
<< m1 >>
rect 96 496 97 497 
<< m1 >>
rect 97 496 98 497 
<< m1 >>
rect 98 496 99 497 
<< m1 >>
rect 99 496 100 497 
<< m1 >>
rect 100 496 101 497 
<< m1 >>
rect 103 496 104 497 
<< m1 >>
rect 118 496 119 497 
<< m1 >>
rect 175 496 176 497 
<< m1 >>
rect 190 496 191 497 
<< m2 >>
rect 190 496 191 497 
<< m2 >>
rect 191 496 192 497 
<< m1 >>
rect 192 496 193 497 
<< m2 >>
rect 192 496 193 497 
<< m2c >>
rect 192 496 193 497 
<< m1 >>
rect 192 496 193 497 
<< m2 >>
rect 192 496 193 497 
<< m1 >>
rect 193 496 194 497 
<< m1 >>
rect 211 496 212 497 
<< m1 >>
rect 253 496 254 497 
<< m1 >>
rect 361 496 362 497 
<< m1 >>
rect 373 496 374 497 
<< m1 >>
rect 379 496 380 497 
<< m1 >>
rect 381 496 382 497 
<< m2 >>
rect 382 496 383 497 
<< m1 >>
rect 406 496 407 497 
<< m1 >>
rect 451 496 452 497 
<< m1 >>
rect 472 496 473 497 
<< m1 >>
rect 487 496 488 497 
<< m1 >>
rect 489 496 490 497 
<< m1 >>
rect 523 496 524 497 
<< m1 >>
rect 28 497 29 498 
<< m1 >>
rect 34 497 35 498 
<< m1 >>
rect 37 497 38 498 
<< m1 >>
rect 73 497 74 498 
<< m1 >>
rect 88 497 89 498 
<< m1 >>
rect 100 497 101 498 
<< m1 >>
rect 103 497 104 498 
<< m1 >>
rect 118 497 119 498 
<< m1 >>
rect 175 497 176 498 
<< m1 >>
rect 186 497 187 498 
<< m1 >>
rect 187 497 188 498 
<< m1 >>
rect 188 497 189 498 
<< m2 >>
rect 188 497 189 498 
<< m2c >>
rect 188 497 189 498 
<< m1 >>
rect 188 497 189 498 
<< m2 >>
rect 188 497 189 498 
<< m2 >>
rect 189 497 190 498 
<< m1 >>
rect 190 497 191 498 
<< m2 >>
rect 190 497 191 498 
<< m1 >>
rect 193 497 194 498 
<< m1 >>
rect 211 497 212 498 
<< m1 >>
rect 253 497 254 498 
<< m1 >>
rect 361 497 362 498 
<< m1 >>
rect 373 497 374 498 
<< m1 >>
rect 379 497 380 498 
<< m1 >>
rect 381 497 382 498 
<< m2 >>
rect 382 497 383 498 
<< m1 >>
rect 406 497 407 498 
<< m1 >>
rect 451 497 452 498 
<< m1 >>
rect 472 497 473 498 
<< m1 >>
rect 487 497 488 498 
<< m1 >>
rect 489 497 490 498 
<< m1 >>
rect 523 497 524 498 
<< pdiffusion >>
rect 12 498 13 499 
<< pdiffusion >>
rect 13 498 14 499 
<< pdiffusion >>
rect 14 498 15 499 
<< pdiffusion >>
rect 15 498 16 499 
<< pdiffusion >>
rect 16 498 17 499 
<< pdiffusion >>
rect 17 498 18 499 
<< m1 >>
rect 28 498 29 499 
<< pdiffusion >>
rect 30 498 31 499 
<< pdiffusion >>
rect 31 498 32 499 
<< pdiffusion >>
rect 32 498 33 499 
<< pdiffusion >>
rect 33 498 34 499 
<< m1 >>
rect 34 498 35 499 
<< pdiffusion >>
rect 34 498 35 499 
<< pdiffusion >>
rect 35 498 36 499 
<< m1 >>
rect 37 498 38 499 
<< pdiffusion >>
rect 48 498 49 499 
<< pdiffusion >>
rect 49 498 50 499 
<< pdiffusion >>
rect 50 498 51 499 
<< pdiffusion >>
rect 51 498 52 499 
<< pdiffusion >>
rect 52 498 53 499 
<< pdiffusion >>
rect 53 498 54 499 
<< pdiffusion >>
rect 66 498 67 499 
<< pdiffusion >>
rect 67 498 68 499 
<< pdiffusion >>
rect 68 498 69 499 
<< pdiffusion >>
rect 69 498 70 499 
<< pdiffusion >>
rect 70 498 71 499 
<< pdiffusion >>
rect 71 498 72 499 
<< m1 >>
rect 73 498 74 499 
<< pdiffusion >>
rect 84 498 85 499 
<< pdiffusion >>
rect 85 498 86 499 
<< pdiffusion >>
rect 86 498 87 499 
<< pdiffusion >>
rect 87 498 88 499 
<< m1 >>
rect 88 498 89 499 
<< pdiffusion >>
rect 88 498 89 499 
<< pdiffusion >>
rect 89 498 90 499 
<< m1 >>
rect 100 498 101 499 
<< pdiffusion >>
rect 102 498 103 499 
<< m1 >>
rect 103 498 104 499 
<< pdiffusion >>
rect 103 498 104 499 
<< pdiffusion >>
rect 104 498 105 499 
<< pdiffusion >>
rect 105 498 106 499 
<< pdiffusion >>
rect 106 498 107 499 
<< pdiffusion >>
rect 107 498 108 499 
<< m1 >>
rect 118 498 119 499 
<< pdiffusion >>
rect 120 498 121 499 
<< pdiffusion >>
rect 121 498 122 499 
<< pdiffusion >>
rect 122 498 123 499 
<< pdiffusion >>
rect 123 498 124 499 
<< pdiffusion >>
rect 124 498 125 499 
<< pdiffusion >>
rect 125 498 126 499 
<< pdiffusion >>
rect 138 498 139 499 
<< pdiffusion >>
rect 139 498 140 499 
<< pdiffusion >>
rect 140 498 141 499 
<< pdiffusion >>
rect 141 498 142 499 
<< pdiffusion >>
rect 142 498 143 499 
<< pdiffusion >>
rect 143 498 144 499 
<< pdiffusion >>
rect 174 498 175 499 
<< m1 >>
rect 175 498 176 499 
<< pdiffusion >>
rect 175 498 176 499 
<< pdiffusion >>
rect 176 498 177 499 
<< pdiffusion >>
rect 177 498 178 499 
<< pdiffusion >>
rect 178 498 179 499 
<< pdiffusion >>
rect 179 498 180 499 
<< m1 >>
rect 186 498 187 499 
<< m1 >>
rect 190 498 191 499 
<< pdiffusion >>
rect 192 498 193 499 
<< m1 >>
rect 193 498 194 499 
<< pdiffusion >>
rect 193 498 194 499 
<< pdiffusion >>
rect 194 498 195 499 
<< pdiffusion >>
rect 195 498 196 499 
<< pdiffusion >>
rect 196 498 197 499 
<< pdiffusion >>
rect 197 498 198 499 
<< pdiffusion >>
rect 210 498 211 499 
<< m1 >>
rect 211 498 212 499 
<< pdiffusion >>
rect 211 498 212 499 
<< pdiffusion >>
rect 212 498 213 499 
<< pdiffusion >>
rect 213 498 214 499 
<< pdiffusion >>
rect 214 498 215 499 
<< pdiffusion >>
rect 215 498 216 499 
<< pdiffusion >>
rect 228 498 229 499 
<< pdiffusion >>
rect 229 498 230 499 
<< pdiffusion >>
rect 230 498 231 499 
<< pdiffusion >>
rect 231 498 232 499 
<< pdiffusion >>
rect 232 498 233 499 
<< pdiffusion >>
rect 233 498 234 499 
<< pdiffusion >>
rect 246 498 247 499 
<< pdiffusion >>
rect 247 498 248 499 
<< pdiffusion >>
rect 248 498 249 499 
<< pdiffusion >>
rect 249 498 250 499 
<< pdiffusion >>
rect 250 498 251 499 
<< pdiffusion >>
rect 251 498 252 499 
<< m1 >>
rect 253 498 254 499 
<< pdiffusion >>
rect 264 498 265 499 
<< pdiffusion >>
rect 265 498 266 499 
<< pdiffusion >>
rect 266 498 267 499 
<< pdiffusion >>
rect 267 498 268 499 
<< pdiffusion >>
rect 268 498 269 499 
<< pdiffusion >>
rect 269 498 270 499 
<< pdiffusion >>
rect 282 498 283 499 
<< pdiffusion >>
rect 283 498 284 499 
<< pdiffusion >>
rect 284 498 285 499 
<< pdiffusion >>
rect 285 498 286 499 
<< pdiffusion >>
rect 286 498 287 499 
<< pdiffusion >>
rect 287 498 288 499 
<< pdiffusion >>
rect 318 498 319 499 
<< pdiffusion >>
rect 319 498 320 499 
<< pdiffusion >>
rect 320 498 321 499 
<< pdiffusion >>
rect 321 498 322 499 
<< pdiffusion >>
rect 322 498 323 499 
<< pdiffusion >>
rect 323 498 324 499 
<< pdiffusion >>
rect 336 498 337 499 
<< pdiffusion >>
rect 337 498 338 499 
<< pdiffusion >>
rect 338 498 339 499 
<< pdiffusion >>
rect 339 498 340 499 
<< pdiffusion >>
rect 340 498 341 499 
<< pdiffusion >>
rect 341 498 342 499 
<< pdiffusion >>
rect 354 498 355 499 
<< pdiffusion >>
rect 355 498 356 499 
<< pdiffusion >>
rect 356 498 357 499 
<< pdiffusion >>
rect 357 498 358 499 
<< pdiffusion >>
rect 358 498 359 499 
<< pdiffusion >>
rect 359 498 360 499 
<< m1 >>
rect 361 498 362 499 
<< pdiffusion >>
rect 372 498 373 499 
<< m1 >>
rect 373 498 374 499 
<< pdiffusion >>
rect 373 498 374 499 
<< pdiffusion >>
rect 374 498 375 499 
<< pdiffusion >>
rect 375 498 376 499 
<< pdiffusion >>
rect 376 498 377 499 
<< pdiffusion >>
rect 377 498 378 499 
<< m1 >>
rect 379 498 380 499 
<< m1 >>
rect 381 498 382 499 
<< m2 >>
rect 382 498 383 499 
<< pdiffusion >>
rect 390 498 391 499 
<< pdiffusion >>
rect 391 498 392 499 
<< pdiffusion >>
rect 392 498 393 499 
<< pdiffusion >>
rect 393 498 394 499 
<< pdiffusion >>
rect 394 498 395 499 
<< pdiffusion >>
rect 395 498 396 499 
<< m1 >>
rect 406 498 407 499 
<< pdiffusion >>
rect 408 498 409 499 
<< pdiffusion >>
rect 409 498 410 499 
<< pdiffusion >>
rect 410 498 411 499 
<< pdiffusion >>
rect 411 498 412 499 
<< pdiffusion >>
rect 412 498 413 499 
<< pdiffusion >>
rect 413 498 414 499 
<< pdiffusion >>
rect 444 498 445 499 
<< pdiffusion >>
rect 445 498 446 499 
<< pdiffusion >>
rect 446 498 447 499 
<< pdiffusion >>
rect 447 498 448 499 
<< pdiffusion >>
rect 448 498 449 499 
<< pdiffusion >>
rect 449 498 450 499 
<< m1 >>
rect 451 498 452 499 
<< pdiffusion >>
rect 462 498 463 499 
<< pdiffusion >>
rect 463 498 464 499 
<< pdiffusion >>
rect 464 498 465 499 
<< pdiffusion >>
rect 465 498 466 499 
<< pdiffusion >>
rect 466 498 467 499 
<< pdiffusion >>
rect 467 498 468 499 
<< m1 >>
rect 472 498 473 499 
<< pdiffusion >>
rect 480 498 481 499 
<< pdiffusion >>
rect 481 498 482 499 
<< pdiffusion >>
rect 482 498 483 499 
<< pdiffusion >>
rect 483 498 484 499 
<< pdiffusion >>
rect 484 498 485 499 
<< pdiffusion >>
rect 485 498 486 499 
<< m1 >>
rect 487 498 488 499 
<< m1 >>
rect 489 498 490 499 
<< pdiffusion >>
rect 498 498 499 499 
<< pdiffusion >>
rect 499 498 500 499 
<< pdiffusion >>
rect 500 498 501 499 
<< pdiffusion >>
rect 501 498 502 499 
<< pdiffusion >>
rect 502 498 503 499 
<< pdiffusion >>
rect 503 498 504 499 
<< pdiffusion >>
rect 516 498 517 499 
<< pdiffusion >>
rect 517 498 518 499 
<< pdiffusion >>
rect 518 498 519 499 
<< pdiffusion >>
rect 519 498 520 499 
<< pdiffusion >>
rect 520 498 521 499 
<< pdiffusion >>
rect 521 498 522 499 
<< m1 >>
rect 523 498 524 499 
<< pdiffusion >>
rect 12 499 13 500 
<< pdiffusion >>
rect 13 499 14 500 
<< pdiffusion >>
rect 14 499 15 500 
<< pdiffusion >>
rect 15 499 16 500 
<< pdiffusion >>
rect 16 499 17 500 
<< pdiffusion >>
rect 17 499 18 500 
<< m1 >>
rect 28 499 29 500 
<< pdiffusion >>
rect 30 499 31 500 
<< pdiffusion >>
rect 31 499 32 500 
<< pdiffusion >>
rect 32 499 33 500 
<< pdiffusion >>
rect 33 499 34 500 
<< pdiffusion >>
rect 34 499 35 500 
<< pdiffusion >>
rect 35 499 36 500 
<< m1 >>
rect 37 499 38 500 
<< pdiffusion >>
rect 48 499 49 500 
<< pdiffusion >>
rect 49 499 50 500 
<< pdiffusion >>
rect 50 499 51 500 
<< pdiffusion >>
rect 51 499 52 500 
<< pdiffusion >>
rect 52 499 53 500 
<< pdiffusion >>
rect 53 499 54 500 
<< pdiffusion >>
rect 66 499 67 500 
<< pdiffusion >>
rect 67 499 68 500 
<< pdiffusion >>
rect 68 499 69 500 
<< pdiffusion >>
rect 69 499 70 500 
<< pdiffusion >>
rect 70 499 71 500 
<< pdiffusion >>
rect 71 499 72 500 
<< m1 >>
rect 73 499 74 500 
<< pdiffusion >>
rect 84 499 85 500 
<< pdiffusion >>
rect 85 499 86 500 
<< pdiffusion >>
rect 86 499 87 500 
<< pdiffusion >>
rect 87 499 88 500 
<< pdiffusion >>
rect 88 499 89 500 
<< pdiffusion >>
rect 89 499 90 500 
<< m1 >>
rect 100 499 101 500 
<< pdiffusion >>
rect 102 499 103 500 
<< pdiffusion >>
rect 103 499 104 500 
<< pdiffusion >>
rect 104 499 105 500 
<< pdiffusion >>
rect 105 499 106 500 
<< pdiffusion >>
rect 106 499 107 500 
<< pdiffusion >>
rect 107 499 108 500 
<< m1 >>
rect 118 499 119 500 
<< pdiffusion >>
rect 120 499 121 500 
<< pdiffusion >>
rect 121 499 122 500 
<< pdiffusion >>
rect 122 499 123 500 
<< pdiffusion >>
rect 123 499 124 500 
<< pdiffusion >>
rect 124 499 125 500 
<< pdiffusion >>
rect 125 499 126 500 
<< pdiffusion >>
rect 138 499 139 500 
<< pdiffusion >>
rect 139 499 140 500 
<< pdiffusion >>
rect 140 499 141 500 
<< pdiffusion >>
rect 141 499 142 500 
<< pdiffusion >>
rect 142 499 143 500 
<< pdiffusion >>
rect 143 499 144 500 
<< pdiffusion >>
rect 174 499 175 500 
<< pdiffusion >>
rect 175 499 176 500 
<< pdiffusion >>
rect 176 499 177 500 
<< pdiffusion >>
rect 177 499 178 500 
<< pdiffusion >>
rect 178 499 179 500 
<< pdiffusion >>
rect 179 499 180 500 
<< m1 >>
rect 186 499 187 500 
<< m1 >>
rect 190 499 191 500 
<< pdiffusion >>
rect 192 499 193 500 
<< pdiffusion >>
rect 193 499 194 500 
<< pdiffusion >>
rect 194 499 195 500 
<< pdiffusion >>
rect 195 499 196 500 
<< pdiffusion >>
rect 196 499 197 500 
<< pdiffusion >>
rect 197 499 198 500 
<< pdiffusion >>
rect 210 499 211 500 
<< pdiffusion >>
rect 211 499 212 500 
<< pdiffusion >>
rect 212 499 213 500 
<< pdiffusion >>
rect 213 499 214 500 
<< pdiffusion >>
rect 214 499 215 500 
<< pdiffusion >>
rect 215 499 216 500 
<< pdiffusion >>
rect 228 499 229 500 
<< pdiffusion >>
rect 229 499 230 500 
<< pdiffusion >>
rect 230 499 231 500 
<< pdiffusion >>
rect 231 499 232 500 
<< pdiffusion >>
rect 232 499 233 500 
<< pdiffusion >>
rect 233 499 234 500 
<< pdiffusion >>
rect 246 499 247 500 
<< pdiffusion >>
rect 247 499 248 500 
<< pdiffusion >>
rect 248 499 249 500 
<< pdiffusion >>
rect 249 499 250 500 
<< pdiffusion >>
rect 250 499 251 500 
<< pdiffusion >>
rect 251 499 252 500 
<< m1 >>
rect 253 499 254 500 
<< pdiffusion >>
rect 264 499 265 500 
<< pdiffusion >>
rect 265 499 266 500 
<< pdiffusion >>
rect 266 499 267 500 
<< pdiffusion >>
rect 267 499 268 500 
<< pdiffusion >>
rect 268 499 269 500 
<< pdiffusion >>
rect 269 499 270 500 
<< pdiffusion >>
rect 282 499 283 500 
<< pdiffusion >>
rect 283 499 284 500 
<< pdiffusion >>
rect 284 499 285 500 
<< pdiffusion >>
rect 285 499 286 500 
<< pdiffusion >>
rect 286 499 287 500 
<< pdiffusion >>
rect 287 499 288 500 
<< pdiffusion >>
rect 318 499 319 500 
<< pdiffusion >>
rect 319 499 320 500 
<< pdiffusion >>
rect 320 499 321 500 
<< pdiffusion >>
rect 321 499 322 500 
<< pdiffusion >>
rect 322 499 323 500 
<< pdiffusion >>
rect 323 499 324 500 
<< pdiffusion >>
rect 336 499 337 500 
<< pdiffusion >>
rect 337 499 338 500 
<< pdiffusion >>
rect 338 499 339 500 
<< pdiffusion >>
rect 339 499 340 500 
<< pdiffusion >>
rect 340 499 341 500 
<< pdiffusion >>
rect 341 499 342 500 
<< pdiffusion >>
rect 354 499 355 500 
<< pdiffusion >>
rect 355 499 356 500 
<< pdiffusion >>
rect 356 499 357 500 
<< pdiffusion >>
rect 357 499 358 500 
<< pdiffusion >>
rect 358 499 359 500 
<< pdiffusion >>
rect 359 499 360 500 
<< m1 >>
rect 361 499 362 500 
<< pdiffusion >>
rect 372 499 373 500 
<< pdiffusion >>
rect 373 499 374 500 
<< pdiffusion >>
rect 374 499 375 500 
<< pdiffusion >>
rect 375 499 376 500 
<< pdiffusion >>
rect 376 499 377 500 
<< pdiffusion >>
rect 377 499 378 500 
<< m1 >>
rect 379 499 380 500 
<< m1 >>
rect 381 499 382 500 
<< m2 >>
rect 382 499 383 500 
<< pdiffusion >>
rect 390 499 391 500 
<< pdiffusion >>
rect 391 499 392 500 
<< pdiffusion >>
rect 392 499 393 500 
<< pdiffusion >>
rect 393 499 394 500 
<< pdiffusion >>
rect 394 499 395 500 
<< pdiffusion >>
rect 395 499 396 500 
<< m1 >>
rect 406 499 407 500 
<< pdiffusion >>
rect 408 499 409 500 
<< pdiffusion >>
rect 409 499 410 500 
<< pdiffusion >>
rect 410 499 411 500 
<< pdiffusion >>
rect 411 499 412 500 
<< pdiffusion >>
rect 412 499 413 500 
<< pdiffusion >>
rect 413 499 414 500 
<< pdiffusion >>
rect 444 499 445 500 
<< pdiffusion >>
rect 445 499 446 500 
<< pdiffusion >>
rect 446 499 447 500 
<< pdiffusion >>
rect 447 499 448 500 
<< pdiffusion >>
rect 448 499 449 500 
<< pdiffusion >>
rect 449 499 450 500 
<< m1 >>
rect 451 499 452 500 
<< pdiffusion >>
rect 462 499 463 500 
<< pdiffusion >>
rect 463 499 464 500 
<< pdiffusion >>
rect 464 499 465 500 
<< pdiffusion >>
rect 465 499 466 500 
<< pdiffusion >>
rect 466 499 467 500 
<< pdiffusion >>
rect 467 499 468 500 
<< m1 >>
rect 472 499 473 500 
<< pdiffusion >>
rect 480 499 481 500 
<< pdiffusion >>
rect 481 499 482 500 
<< pdiffusion >>
rect 482 499 483 500 
<< pdiffusion >>
rect 483 499 484 500 
<< pdiffusion >>
rect 484 499 485 500 
<< pdiffusion >>
rect 485 499 486 500 
<< m1 >>
rect 487 499 488 500 
<< m1 >>
rect 489 499 490 500 
<< pdiffusion >>
rect 498 499 499 500 
<< pdiffusion >>
rect 499 499 500 500 
<< pdiffusion >>
rect 500 499 501 500 
<< pdiffusion >>
rect 501 499 502 500 
<< pdiffusion >>
rect 502 499 503 500 
<< pdiffusion >>
rect 503 499 504 500 
<< pdiffusion >>
rect 516 499 517 500 
<< pdiffusion >>
rect 517 499 518 500 
<< pdiffusion >>
rect 518 499 519 500 
<< pdiffusion >>
rect 519 499 520 500 
<< pdiffusion >>
rect 520 499 521 500 
<< pdiffusion >>
rect 521 499 522 500 
<< m1 >>
rect 523 499 524 500 
<< pdiffusion >>
rect 12 500 13 501 
<< pdiffusion >>
rect 13 500 14 501 
<< pdiffusion >>
rect 14 500 15 501 
<< pdiffusion >>
rect 15 500 16 501 
<< pdiffusion >>
rect 16 500 17 501 
<< pdiffusion >>
rect 17 500 18 501 
<< m1 >>
rect 28 500 29 501 
<< pdiffusion >>
rect 30 500 31 501 
<< pdiffusion >>
rect 31 500 32 501 
<< pdiffusion >>
rect 32 500 33 501 
<< pdiffusion >>
rect 33 500 34 501 
<< pdiffusion >>
rect 34 500 35 501 
<< pdiffusion >>
rect 35 500 36 501 
<< m1 >>
rect 37 500 38 501 
<< pdiffusion >>
rect 48 500 49 501 
<< pdiffusion >>
rect 49 500 50 501 
<< pdiffusion >>
rect 50 500 51 501 
<< pdiffusion >>
rect 51 500 52 501 
<< pdiffusion >>
rect 52 500 53 501 
<< pdiffusion >>
rect 53 500 54 501 
<< pdiffusion >>
rect 66 500 67 501 
<< pdiffusion >>
rect 67 500 68 501 
<< pdiffusion >>
rect 68 500 69 501 
<< pdiffusion >>
rect 69 500 70 501 
<< pdiffusion >>
rect 70 500 71 501 
<< pdiffusion >>
rect 71 500 72 501 
<< m1 >>
rect 73 500 74 501 
<< pdiffusion >>
rect 84 500 85 501 
<< pdiffusion >>
rect 85 500 86 501 
<< pdiffusion >>
rect 86 500 87 501 
<< pdiffusion >>
rect 87 500 88 501 
<< pdiffusion >>
rect 88 500 89 501 
<< pdiffusion >>
rect 89 500 90 501 
<< m1 >>
rect 100 500 101 501 
<< pdiffusion >>
rect 102 500 103 501 
<< pdiffusion >>
rect 103 500 104 501 
<< pdiffusion >>
rect 104 500 105 501 
<< pdiffusion >>
rect 105 500 106 501 
<< pdiffusion >>
rect 106 500 107 501 
<< pdiffusion >>
rect 107 500 108 501 
<< m1 >>
rect 118 500 119 501 
<< pdiffusion >>
rect 120 500 121 501 
<< pdiffusion >>
rect 121 500 122 501 
<< pdiffusion >>
rect 122 500 123 501 
<< pdiffusion >>
rect 123 500 124 501 
<< pdiffusion >>
rect 124 500 125 501 
<< pdiffusion >>
rect 125 500 126 501 
<< pdiffusion >>
rect 138 500 139 501 
<< pdiffusion >>
rect 139 500 140 501 
<< pdiffusion >>
rect 140 500 141 501 
<< pdiffusion >>
rect 141 500 142 501 
<< pdiffusion >>
rect 142 500 143 501 
<< pdiffusion >>
rect 143 500 144 501 
<< pdiffusion >>
rect 174 500 175 501 
<< pdiffusion >>
rect 175 500 176 501 
<< pdiffusion >>
rect 176 500 177 501 
<< pdiffusion >>
rect 177 500 178 501 
<< pdiffusion >>
rect 178 500 179 501 
<< pdiffusion >>
rect 179 500 180 501 
<< m1 >>
rect 186 500 187 501 
<< m1 >>
rect 190 500 191 501 
<< pdiffusion >>
rect 192 500 193 501 
<< pdiffusion >>
rect 193 500 194 501 
<< pdiffusion >>
rect 194 500 195 501 
<< pdiffusion >>
rect 195 500 196 501 
<< pdiffusion >>
rect 196 500 197 501 
<< pdiffusion >>
rect 197 500 198 501 
<< pdiffusion >>
rect 210 500 211 501 
<< pdiffusion >>
rect 211 500 212 501 
<< pdiffusion >>
rect 212 500 213 501 
<< pdiffusion >>
rect 213 500 214 501 
<< pdiffusion >>
rect 214 500 215 501 
<< pdiffusion >>
rect 215 500 216 501 
<< pdiffusion >>
rect 228 500 229 501 
<< pdiffusion >>
rect 229 500 230 501 
<< pdiffusion >>
rect 230 500 231 501 
<< pdiffusion >>
rect 231 500 232 501 
<< pdiffusion >>
rect 232 500 233 501 
<< pdiffusion >>
rect 233 500 234 501 
<< pdiffusion >>
rect 246 500 247 501 
<< pdiffusion >>
rect 247 500 248 501 
<< pdiffusion >>
rect 248 500 249 501 
<< pdiffusion >>
rect 249 500 250 501 
<< pdiffusion >>
rect 250 500 251 501 
<< pdiffusion >>
rect 251 500 252 501 
<< m1 >>
rect 253 500 254 501 
<< pdiffusion >>
rect 264 500 265 501 
<< pdiffusion >>
rect 265 500 266 501 
<< pdiffusion >>
rect 266 500 267 501 
<< pdiffusion >>
rect 267 500 268 501 
<< pdiffusion >>
rect 268 500 269 501 
<< pdiffusion >>
rect 269 500 270 501 
<< pdiffusion >>
rect 282 500 283 501 
<< pdiffusion >>
rect 283 500 284 501 
<< pdiffusion >>
rect 284 500 285 501 
<< pdiffusion >>
rect 285 500 286 501 
<< pdiffusion >>
rect 286 500 287 501 
<< pdiffusion >>
rect 287 500 288 501 
<< pdiffusion >>
rect 318 500 319 501 
<< pdiffusion >>
rect 319 500 320 501 
<< pdiffusion >>
rect 320 500 321 501 
<< pdiffusion >>
rect 321 500 322 501 
<< pdiffusion >>
rect 322 500 323 501 
<< pdiffusion >>
rect 323 500 324 501 
<< pdiffusion >>
rect 336 500 337 501 
<< pdiffusion >>
rect 337 500 338 501 
<< pdiffusion >>
rect 338 500 339 501 
<< pdiffusion >>
rect 339 500 340 501 
<< pdiffusion >>
rect 340 500 341 501 
<< pdiffusion >>
rect 341 500 342 501 
<< pdiffusion >>
rect 354 500 355 501 
<< pdiffusion >>
rect 355 500 356 501 
<< pdiffusion >>
rect 356 500 357 501 
<< pdiffusion >>
rect 357 500 358 501 
<< pdiffusion >>
rect 358 500 359 501 
<< pdiffusion >>
rect 359 500 360 501 
<< m1 >>
rect 361 500 362 501 
<< pdiffusion >>
rect 372 500 373 501 
<< pdiffusion >>
rect 373 500 374 501 
<< pdiffusion >>
rect 374 500 375 501 
<< pdiffusion >>
rect 375 500 376 501 
<< pdiffusion >>
rect 376 500 377 501 
<< pdiffusion >>
rect 377 500 378 501 
<< m1 >>
rect 379 500 380 501 
<< m1 >>
rect 381 500 382 501 
<< m2 >>
rect 382 500 383 501 
<< pdiffusion >>
rect 390 500 391 501 
<< pdiffusion >>
rect 391 500 392 501 
<< pdiffusion >>
rect 392 500 393 501 
<< pdiffusion >>
rect 393 500 394 501 
<< pdiffusion >>
rect 394 500 395 501 
<< pdiffusion >>
rect 395 500 396 501 
<< m1 >>
rect 406 500 407 501 
<< pdiffusion >>
rect 408 500 409 501 
<< pdiffusion >>
rect 409 500 410 501 
<< pdiffusion >>
rect 410 500 411 501 
<< pdiffusion >>
rect 411 500 412 501 
<< pdiffusion >>
rect 412 500 413 501 
<< pdiffusion >>
rect 413 500 414 501 
<< pdiffusion >>
rect 444 500 445 501 
<< pdiffusion >>
rect 445 500 446 501 
<< pdiffusion >>
rect 446 500 447 501 
<< pdiffusion >>
rect 447 500 448 501 
<< pdiffusion >>
rect 448 500 449 501 
<< pdiffusion >>
rect 449 500 450 501 
<< m1 >>
rect 451 500 452 501 
<< pdiffusion >>
rect 462 500 463 501 
<< pdiffusion >>
rect 463 500 464 501 
<< pdiffusion >>
rect 464 500 465 501 
<< pdiffusion >>
rect 465 500 466 501 
<< pdiffusion >>
rect 466 500 467 501 
<< pdiffusion >>
rect 467 500 468 501 
<< m1 >>
rect 472 500 473 501 
<< pdiffusion >>
rect 480 500 481 501 
<< pdiffusion >>
rect 481 500 482 501 
<< pdiffusion >>
rect 482 500 483 501 
<< pdiffusion >>
rect 483 500 484 501 
<< pdiffusion >>
rect 484 500 485 501 
<< pdiffusion >>
rect 485 500 486 501 
<< m1 >>
rect 487 500 488 501 
<< m1 >>
rect 489 500 490 501 
<< pdiffusion >>
rect 498 500 499 501 
<< pdiffusion >>
rect 499 500 500 501 
<< pdiffusion >>
rect 500 500 501 501 
<< pdiffusion >>
rect 501 500 502 501 
<< pdiffusion >>
rect 502 500 503 501 
<< pdiffusion >>
rect 503 500 504 501 
<< pdiffusion >>
rect 516 500 517 501 
<< pdiffusion >>
rect 517 500 518 501 
<< pdiffusion >>
rect 518 500 519 501 
<< pdiffusion >>
rect 519 500 520 501 
<< pdiffusion >>
rect 520 500 521 501 
<< pdiffusion >>
rect 521 500 522 501 
<< m1 >>
rect 523 500 524 501 
<< pdiffusion >>
rect 12 501 13 502 
<< pdiffusion >>
rect 13 501 14 502 
<< pdiffusion >>
rect 14 501 15 502 
<< pdiffusion >>
rect 15 501 16 502 
<< pdiffusion >>
rect 16 501 17 502 
<< pdiffusion >>
rect 17 501 18 502 
<< m1 >>
rect 28 501 29 502 
<< pdiffusion >>
rect 30 501 31 502 
<< pdiffusion >>
rect 31 501 32 502 
<< pdiffusion >>
rect 32 501 33 502 
<< pdiffusion >>
rect 33 501 34 502 
<< pdiffusion >>
rect 34 501 35 502 
<< pdiffusion >>
rect 35 501 36 502 
<< m1 >>
rect 37 501 38 502 
<< pdiffusion >>
rect 48 501 49 502 
<< pdiffusion >>
rect 49 501 50 502 
<< pdiffusion >>
rect 50 501 51 502 
<< pdiffusion >>
rect 51 501 52 502 
<< pdiffusion >>
rect 52 501 53 502 
<< pdiffusion >>
rect 53 501 54 502 
<< pdiffusion >>
rect 66 501 67 502 
<< pdiffusion >>
rect 67 501 68 502 
<< pdiffusion >>
rect 68 501 69 502 
<< pdiffusion >>
rect 69 501 70 502 
<< pdiffusion >>
rect 70 501 71 502 
<< pdiffusion >>
rect 71 501 72 502 
<< m1 >>
rect 73 501 74 502 
<< pdiffusion >>
rect 84 501 85 502 
<< pdiffusion >>
rect 85 501 86 502 
<< pdiffusion >>
rect 86 501 87 502 
<< pdiffusion >>
rect 87 501 88 502 
<< pdiffusion >>
rect 88 501 89 502 
<< pdiffusion >>
rect 89 501 90 502 
<< m1 >>
rect 100 501 101 502 
<< pdiffusion >>
rect 102 501 103 502 
<< pdiffusion >>
rect 103 501 104 502 
<< pdiffusion >>
rect 104 501 105 502 
<< pdiffusion >>
rect 105 501 106 502 
<< pdiffusion >>
rect 106 501 107 502 
<< pdiffusion >>
rect 107 501 108 502 
<< m1 >>
rect 118 501 119 502 
<< pdiffusion >>
rect 120 501 121 502 
<< pdiffusion >>
rect 121 501 122 502 
<< pdiffusion >>
rect 122 501 123 502 
<< pdiffusion >>
rect 123 501 124 502 
<< pdiffusion >>
rect 124 501 125 502 
<< pdiffusion >>
rect 125 501 126 502 
<< pdiffusion >>
rect 138 501 139 502 
<< pdiffusion >>
rect 139 501 140 502 
<< pdiffusion >>
rect 140 501 141 502 
<< pdiffusion >>
rect 141 501 142 502 
<< pdiffusion >>
rect 142 501 143 502 
<< pdiffusion >>
rect 143 501 144 502 
<< pdiffusion >>
rect 174 501 175 502 
<< pdiffusion >>
rect 175 501 176 502 
<< pdiffusion >>
rect 176 501 177 502 
<< pdiffusion >>
rect 177 501 178 502 
<< pdiffusion >>
rect 178 501 179 502 
<< pdiffusion >>
rect 179 501 180 502 
<< m1 >>
rect 186 501 187 502 
<< m1 >>
rect 190 501 191 502 
<< pdiffusion >>
rect 192 501 193 502 
<< pdiffusion >>
rect 193 501 194 502 
<< pdiffusion >>
rect 194 501 195 502 
<< pdiffusion >>
rect 195 501 196 502 
<< pdiffusion >>
rect 196 501 197 502 
<< pdiffusion >>
rect 197 501 198 502 
<< pdiffusion >>
rect 210 501 211 502 
<< pdiffusion >>
rect 211 501 212 502 
<< pdiffusion >>
rect 212 501 213 502 
<< pdiffusion >>
rect 213 501 214 502 
<< pdiffusion >>
rect 214 501 215 502 
<< pdiffusion >>
rect 215 501 216 502 
<< pdiffusion >>
rect 228 501 229 502 
<< pdiffusion >>
rect 229 501 230 502 
<< pdiffusion >>
rect 230 501 231 502 
<< pdiffusion >>
rect 231 501 232 502 
<< pdiffusion >>
rect 232 501 233 502 
<< pdiffusion >>
rect 233 501 234 502 
<< pdiffusion >>
rect 246 501 247 502 
<< pdiffusion >>
rect 247 501 248 502 
<< pdiffusion >>
rect 248 501 249 502 
<< pdiffusion >>
rect 249 501 250 502 
<< pdiffusion >>
rect 250 501 251 502 
<< pdiffusion >>
rect 251 501 252 502 
<< m1 >>
rect 253 501 254 502 
<< pdiffusion >>
rect 264 501 265 502 
<< pdiffusion >>
rect 265 501 266 502 
<< pdiffusion >>
rect 266 501 267 502 
<< pdiffusion >>
rect 267 501 268 502 
<< pdiffusion >>
rect 268 501 269 502 
<< pdiffusion >>
rect 269 501 270 502 
<< pdiffusion >>
rect 282 501 283 502 
<< pdiffusion >>
rect 283 501 284 502 
<< pdiffusion >>
rect 284 501 285 502 
<< pdiffusion >>
rect 285 501 286 502 
<< pdiffusion >>
rect 286 501 287 502 
<< pdiffusion >>
rect 287 501 288 502 
<< pdiffusion >>
rect 318 501 319 502 
<< pdiffusion >>
rect 319 501 320 502 
<< pdiffusion >>
rect 320 501 321 502 
<< pdiffusion >>
rect 321 501 322 502 
<< pdiffusion >>
rect 322 501 323 502 
<< pdiffusion >>
rect 323 501 324 502 
<< pdiffusion >>
rect 336 501 337 502 
<< pdiffusion >>
rect 337 501 338 502 
<< pdiffusion >>
rect 338 501 339 502 
<< pdiffusion >>
rect 339 501 340 502 
<< pdiffusion >>
rect 340 501 341 502 
<< pdiffusion >>
rect 341 501 342 502 
<< pdiffusion >>
rect 354 501 355 502 
<< pdiffusion >>
rect 355 501 356 502 
<< pdiffusion >>
rect 356 501 357 502 
<< pdiffusion >>
rect 357 501 358 502 
<< pdiffusion >>
rect 358 501 359 502 
<< pdiffusion >>
rect 359 501 360 502 
<< m1 >>
rect 361 501 362 502 
<< pdiffusion >>
rect 372 501 373 502 
<< pdiffusion >>
rect 373 501 374 502 
<< pdiffusion >>
rect 374 501 375 502 
<< pdiffusion >>
rect 375 501 376 502 
<< pdiffusion >>
rect 376 501 377 502 
<< pdiffusion >>
rect 377 501 378 502 
<< m1 >>
rect 379 501 380 502 
<< m1 >>
rect 381 501 382 502 
<< m2 >>
rect 382 501 383 502 
<< pdiffusion >>
rect 390 501 391 502 
<< pdiffusion >>
rect 391 501 392 502 
<< pdiffusion >>
rect 392 501 393 502 
<< pdiffusion >>
rect 393 501 394 502 
<< pdiffusion >>
rect 394 501 395 502 
<< pdiffusion >>
rect 395 501 396 502 
<< m1 >>
rect 406 501 407 502 
<< pdiffusion >>
rect 408 501 409 502 
<< pdiffusion >>
rect 409 501 410 502 
<< pdiffusion >>
rect 410 501 411 502 
<< pdiffusion >>
rect 411 501 412 502 
<< pdiffusion >>
rect 412 501 413 502 
<< pdiffusion >>
rect 413 501 414 502 
<< pdiffusion >>
rect 444 501 445 502 
<< pdiffusion >>
rect 445 501 446 502 
<< pdiffusion >>
rect 446 501 447 502 
<< pdiffusion >>
rect 447 501 448 502 
<< pdiffusion >>
rect 448 501 449 502 
<< pdiffusion >>
rect 449 501 450 502 
<< m1 >>
rect 451 501 452 502 
<< pdiffusion >>
rect 462 501 463 502 
<< pdiffusion >>
rect 463 501 464 502 
<< pdiffusion >>
rect 464 501 465 502 
<< pdiffusion >>
rect 465 501 466 502 
<< pdiffusion >>
rect 466 501 467 502 
<< pdiffusion >>
rect 467 501 468 502 
<< m1 >>
rect 472 501 473 502 
<< pdiffusion >>
rect 480 501 481 502 
<< pdiffusion >>
rect 481 501 482 502 
<< pdiffusion >>
rect 482 501 483 502 
<< pdiffusion >>
rect 483 501 484 502 
<< pdiffusion >>
rect 484 501 485 502 
<< pdiffusion >>
rect 485 501 486 502 
<< m1 >>
rect 487 501 488 502 
<< m1 >>
rect 489 501 490 502 
<< pdiffusion >>
rect 498 501 499 502 
<< pdiffusion >>
rect 499 501 500 502 
<< pdiffusion >>
rect 500 501 501 502 
<< pdiffusion >>
rect 501 501 502 502 
<< pdiffusion >>
rect 502 501 503 502 
<< pdiffusion >>
rect 503 501 504 502 
<< pdiffusion >>
rect 516 501 517 502 
<< pdiffusion >>
rect 517 501 518 502 
<< pdiffusion >>
rect 518 501 519 502 
<< pdiffusion >>
rect 519 501 520 502 
<< pdiffusion >>
rect 520 501 521 502 
<< pdiffusion >>
rect 521 501 522 502 
<< m1 >>
rect 523 501 524 502 
<< pdiffusion >>
rect 12 502 13 503 
<< pdiffusion >>
rect 13 502 14 503 
<< pdiffusion >>
rect 14 502 15 503 
<< pdiffusion >>
rect 15 502 16 503 
<< pdiffusion >>
rect 16 502 17 503 
<< pdiffusion >>
rect 17 502 18 503 
<< m1 >>
rect 28 502 29 503 
<< pdiffusion >>
rect 30 502 31 503 
<< pdiffusion >>
rect 31 502 32 503 
<< pdiffusion >>
rect 32 502 33 503 
<< pdiffusion >>
rect 33 502 34 503 
<< pdiffusion >>
rect 34 502 35 503 
<< pdiffusion >>
rect 35 502 36 503 
<< m1 >>
rect 37 502 38 503 
<< pdiffusion >>
rect 48 502 49 503 
<< pdiffusion >>
rect 49 502 50 503 
<< pdiffusion >>
rect 50 502 51 503 
<< pdiffusion >>
rect 51 502 52 503 
<< pdiffusion >>
rect 52 502 53 503 
<< pdiffusion >>
rect 53 502 54 503 
<< pdiffusion >>
rect 66 502 67 503 
<< pdiffusion >>
rect 67 502 68 503 
<< pdiffusion >>
rect 68 502 69 503 
<< pdiffusion >>
rect 69 502 70 503 
<< pdiffusion >>
rect 70 502 71 503 
<< pdiffusion >>
rect 71 502 72 503 
<< m1 >>
rect 73 502 74 503 
<< pdiffusion >>
rect 84 502 85 503 
<< pdiffusion >>
rect 85 502 86 503 
<< pdiffusion >>
rect 86 502 87 503 
<< pdiffusion >>
rect 87 502 88 503 
<< pdiffusion >>
rect 88 502 89 503 
<< pdiffusion >>
rect 89 502 90 503 
<< m1 >>
rect 100 502 101 503 
<< pdiffusion >>
rect 102 502 103 503 
<< pdiffusion >>
rect 103 502 104 503 
<< pdiffusion >>
rect 104 502 105 503 
<< pdiffusion >>
rect 105 502 106 503 
<< pdiffusion >>
rect 106 502 107 503 
<< pdiffusion >>
rect 107 502 108 503 
<< m1 >>
rect 118 502 119 503 
<< pdiffusion >>
rect 120 502 121 503 
<< pdiffusion >>
rect 121 502 122 503 
<< pdiffusion >>
rect 122 502 123 503 
<< pdiffusion >>
rect 123 502 124 503 
<< pdiffusion >>
rect 124 502 125 503 
<< pdiffusion >>
rect 125 502 126 503 
<< pdiffusion >>
rect 138 502 139 503 
<< pdiffusion >>
rect 139 502 140 503 
<< pdiffusion >>
rect 140 502 141 503 
<< pdiffusion >>
rect 141 502 142 503 
<< pdiffusion >>
rect 142 502 143 503 
<< pdiffusion >>
rect 143 502 144 503 
<< pdiffusion >>
rect 174 502 175 503 
<< pdiffusion >>
rect 175 502 176 503 
<< pdiffusion >>
rect 176 502 177 503 
<< pdiffusion >>
rect 177 502 178 503 
<< pdiffusion >>
rect 178 502 179 503 
<< pdiffusion >>
rect 179 502 180 503 
<< m1 >>
rect 186 502 187 503 
<< m1 >>
rect 190 502 191 503 
<< pdiffusion >>
rect 192 502 193 503 
<< pdiffusion >>
rect 193 502 194 503 
<< pdiffusion >>
rect 194 502 195 503 
<< pdiffusion >>
rect 195 502 196 503 
<< pdiffusion >>
rect 196 502 197 503 
<< pdiffusion >>
rect 197 502 198 503 
<< pdiffusion >>
rect 210 502 211 503 
<< pdiffusion >>
rect 211 502 212 503 
<< pdiffusion >>
rect 212 502 213 503 
<< pdiffusion >>
rect 213 502 214 503 
<< pdiffusion >>
rect 214 502 215 503 
<< pdiffusion >>
rect 215 502 216 503 
<< pdiffusion >>
rect 228 502 229 503 
<< pdiffusion >>
rect 229 502 230 503 
<< pdiffusion >>
rect 230 502 231 503 
<< pdiffusion >>
rect 231 502 232 503 
<< pdiffusion >>
rect 232 502 233 503 
<< pdiffusion >>
rect 233 502 234 503 
<< pdiffusion >>
rect 246 502 247 503 
<< pdiffusion >>
rect 247 502 248 503 
<< pdiffusion >>
rect 248 502 249 503 
<< pdiffusion >>
rect 249 502 250 503 
<< pdiffusion >>
rect 250 502 251 503 
<< pdiffusion >>
rect 251 502 252 503 
<< m1 >>
rect 253 502 254 503 
<< pdiffusion >>
rect 264 502 265 503 
<< pdiffusion >>
rect 265 502 266 503 
<< pdiffusion >>
rect 266 502 267 503 
<< pdiffusion >>
rect 267 502 268 503 
<< pdiffusion >>
rect 268 502 269 503 
<< pdiffusion >>
rect 269 502 270 503 
<< pdiffusion >>
rect 282 502 283 503 
<< pdiffusion >>
rect 283 502 284 503 
<< pdiffusion >>
rect 284 502 285 503 
<< pdiffusion >>
rect 285 502 286 503 
<< pdiffusion >>
rect 286 502 287 503 
<< pdiffusion >>
rect 287 502 288 503 
<< pdiffusion >>
rect 318 502 319 503 
<< pdiffusion >>
rect 319 502 320 503 
<< pdiffusion >>
rect 320 502 321 503 
<< pdiffusion >>
rect 321 502 322 503 
<< pdiffusion >>
rect 322 502 323 503 
<< pdiffusion >>
rect 323 502 324 503 
<< pdiffusion >>
rect 336 502 337 503 
<< pdiffusion >>
rect 337 502 338 503 
<< pdiffusion >>
rect 338 502 339 503 
<< pdiffusion >>
rect 339 502 340 503 
<< pdiffusion >>
rect 340 502 341 503 
<< pdiffusion >>
rect 341 502 342 503 
<< pdiffusion >>
rect 354 502 355 503 
<< pdiffusion >>
rect 355 502 356 503 
<< pdiffusion >>
rect 356 502 357 503 
<< pdiffusion >>
rect 357 502 358 503 
<< pdiffusion >>
rect 358 502 359 503 
<< pdiffusion >>
rect 359 502 360 503 
<< m1 >>
rect 361 502 362 503 
<< pdiffusion >>
rect 372 502 373 503 
<< pdiffusion >>
rect 373 502 374 503 
<< pdiffusion >>
rect 374 502 375 503 
<< pdiffusion >>
rect 375 502 376 503 
<< pdiffusion >>
rect 376 502 377 503 
<< pdiffusion >>
rect 377 502 378 503 
<< m1 >>
rect 379 502 380 503 
<< m1 >>
rect 381 502 382 503 
<< m2 >>
rect 382 502 383 503 
<< pdiffusion >>
rect 390 502 391 503 
<< pdiffusion >>
rect 391 502 392 503 
<< pdiffusion >>
rect 392 502 393 503 
<< pdiffusion >>
rect 393 502 394 503 
<< pdiffusion >>
rect 394 502 395 503 
<< pdiffusion >>
rect 395 502 396 503 
<< m1 >>
rect 406 502 407 503 
<< pdiffusion >>
rect 408 502 409 503 
<< pdiffusion >>
rect 409 502 410 503 
<< pdiffusion >>
rect 410 502 411 503 
<< pdiffusion >>
rect 411 502 412 503 
<< pdiffusion >>
rect 412 502 413 503 
<< pdiffusion >>
rect 413 502 414 503 
<< pdiffusion >>
rect 444 502 445 503 
<< pdiffusion >>
rect 445 502 446 503 
<< pdiffusion >>
rect 446 502 447 503 
<< pdiffusion >>
rect 447 502 448 503 
<< pdiffusion >>
rect 448 502 449 503 
<< pdiffusion >>
rect 449 502 450 503 
<< m1 >>
rect 451 502 452 503 
<< pdiffusion >>
rect 462 502 463 503 
<< pdiffusion >>
rect 463 502 464 503 
<< pdiffusion >>
rect 464 502 465 503 
<< pdiffusion >>
rect 465 502 466 503 
<< pdiffusion >>
rect 466 502 467 503 
<< pdiffusion >>
rect 467 502 468 503 
<< m1 >>
rect 472 502 473 503 
<< pdiffusion >>
rect 480 502 481 503 
<< pdiffusion >>
rect 481 502 482 503 
<< pdiffusion >>
rect 482 502 483 503 
<< pdiffusion >>
rect 483 502 484 503 
<< pdiffusion >>
rect 484 502 485 503 
<< pdiffusion >>
rect 485 502 486 503 
<< m1 >>
rect 487 502 488 503 
<< m1 >>
rect 489 502 490 503 
<< pdiffusion >>
rect 498 502 499 503 
<< pdiffusion >>
rect 499 502 500 503 
<< pdiffusion >>
rect 500 502 501 503 
<< pdiffusion >>
rect 501 502 502 503 
<< pdiffusion >>
rect 502 502 503 503 
<< pdiffusion >>
rect 503 502 504 503 
<< pdiffusion >>
rect 516 502 517 503 
<< pdiffusion >>
rect 517 502 518 503 
<< pdiffusion >>
rect 518 502 519 503 
<< pdiffusion >>
rect 519 502 520 503 
<< pdiffusion >>
rect 520 502 521 503 
<< pdiffusion >>
rect 521 502 522 503 
<< m1 >>
rect 523 502 524 503 
<< pdiffusion >>
rect 12 503 13 504 
<< m1 >>
rect 13 503 14 504 
<< pdiffusion >>
rect 13 503 14 504 
<< pdiffusion >>
rect 14 503 15 504 
<< pdiffusion >>
rect 15 503 16 504 
<< pdiffusion >>
rect 16 503 17 504 
<< pdiffusion >>
rect 17 503 18 504 
<< m1 >>
rect 28 503 29 504 
<< pdiffusion >>
rect 30 503 31 504 
<< pdiffusion >>
rect 31 503 32 504 
<< pdiffusion >>
rect 32 503 33 504 
<< pdiffusion >>
rect 33 503 34 504 
<< pdiffusion >>
rect 34 503 35 504 
<< pdiffusion >>
rect 35 503 36 504 
<< m1 >>
rect 37 503 38 504 
<< pdiffusion >>
rect 48 503 49 504 
<< m1 >>
rect 49 503 50 504 
<< pdiffusion >>
rect 49 503 50 504 
<< pdiffusion >>
rect 50 503 51 504 
<< pdiffusion >>
rect 51 503 52 504 
<< pdiffusion >>
rect 52 503 53 504 
<< pdiffusion >>
rect 53 503 54 504 
<< pdiffusion >>
rect 66 503 67 504 
<< pdiffusion >>
rect 67 503 68 504 
<< pdiffusion >>
rect 68 503 69 504 
<< pdiffusion >>
rect 69 503 70 504 
<< pdiffusion >>
rect 70 503 71 504 
<< pdiffusion >>
rect 71 503 72 504 
<< m1 >>
rect 73 503 74 504 
<< pdiffusion >>
rect 84 503 85 504 
<< pdiffusion >>
rect 85 503 86 504 
<< pdiffusion >>
rect 86 503 87 504 
<< pdiffusion >>
rect 87 503 88 504 
<< pdiffusion >>
rect 88 503 89 504 
<< pdiffusion >>
rect 89 503 90 504 
<< m1 >>
rect 100 503 101 504 
<< pdiffusion >>
rect 102 503 103 504 
<< pdiffusion >>
rect 103 503 104 504 
<< pdiffusion >>
rect 104 503 105 504 
<< pdiffusion >>
rect 105 503 106 504 
<< pdiffusion >>
rect 106 503 107 504 
<< pdiffusion >>
rect 107 503 108 504 
<< m1 >>
rect 118 503 119 504 
<< pdiffusion >>
rect 120 503 121 504 
<< pdiffusion >>
rect 121 503 122 504 
<< pdiffusion >>
rect 122 503 123 504 
<< pdiffusion >>
rect 123 503 124 504 
<< pdiffusion >>
rect 124 503 125 504 
<< pdiffusion >>
rect 125 503 126 504 
<< pdiffusion >>
rect 138 503 139 504 
<< pdiffusion >>
rect 139 503 140 504 
<< pdiffusion >>
rect 140 503 141 504 
<< pdiffusion >>
rect 141 503 142 504 
<< m1 >>
rect 142 503 143 504 
<< pdiffusion >>
rect 142 503 143 504 
<< pdiffusion >>
rect 143 503 144 504 
<< pdiffusion >>
rect 174 503 175 504 
<< pdiffusion >>
rect 175 503 176 504 
<< pdiffusion >>
rect 176 503 177 504 
<< pdiffusion >>
rect 177 503 178 504 
<< pdiffusion >>
rect 178 503 179 504 
<< pdiffusion >>
rect 179 503 180 504 
<< m1 >>
rect 186 503 187 504 
<< m1 >>
rect 190 503 191 504 
<< pdiffusion >>
rect 192 503 193 504 
<< pdiffusion >>
rect 193 503 194 504 
<< pdiffusion >>
rect 194 503 195 504 
<< pdiffusion >>
rect 195 503 196 504 
<< pdiffusion >>
rect 196 503 197 504 
<< pdiffusion >>
rect 197 503 198 504 
<< pdiffusion >>
rect 210 503 211 504 
<< pdiffusion >>
rect 211 503 212 504 
<< pdiffusion >>
rect 212 503 213 504 
<< pdiffusion >>
rect 213 503 214 504 
<< pdiffusion >>
rect 214 503 215 504 
<< pdiffusion >>
rect 215 503 216 504 
<< pdiffusion >>
rect 228 503 229 504 
<< pdiffusion >>
rect 229 503 230 504 
<< pdiffusion >>
rect 230 503 231 504 
<< pdiffusion >>
rect 231 503 232 504 
<< pdiffusion >>
rect 232 503 233 504 
<< pdiffusion >>
rect 233 503 234 504 
<< pdiffusion >>
rect 246 503 247 504 
<< pdiffusion >>
rect 247 503 248 504 
<< pdiffusion >>
rect 248 503 249 504 
<< pdiffusion >>
rect 249 503 250 504 
<< m1 >>
rect 250 503 251 504 
<< pdiffusion >>
rect 250 503 251 504 
<< pdiffusion >>
rect 251 503 252 504 
<< m1 >>
rect 253 503 254 504 
<< pdiffusion >>
rect 264 503 265 504 
<< pdiffusion >>
rect 265 503 266 504 
<< pdiffusion >>
rect 266 503 267 504 
<< pdiffusion >>
rect 267 503 268 504 
<< pdiffusion >>
rect 268 503 269 504 
<< pdiffusion >>
rect 269 503 270 504 
<< pdiffusion >>
rect 282 503 283 504 
<< pdiffusion >>
rect 283 503 284 504 
<< pdiffusion >>
rect 284 503 285 504 
<< pdiffusion >>
rect 285 503 286 504 
<< pdiffusion >>
rect 286 503 287 504 
<< pdiffusion >>
rect 287 503 288 504 
<< pdiffusion >>
rect 318 503 319 504 
<< m1 >>
rect 319 503 320 504 
<< pdiffusion >>
rect 319 503 320 504 
<< pdiffusion >>
rect 320 503 321 504 
<< pdiffusion >>
rect 321 503 322 504 
<< pdiffusion >>
rect 322 503 323 504 
<< pdiffusion >>
rect 323 503 324 504 
<< pdiffusion >>
rect 336 503 337 504 
<< pdiffusion >>
rect 337 503 338 504 
<< pdiffusion >>
rect 338 503 339 504 
<< pdiffusion >>
rect 339 503 340 504 
<< pdiffusion >>
rect 340 503 341 504 
<< pdiffusion >>
rect 341 503 342 504 
<< pdiffusion >>
rect 354 503 355 504 
<< pdiffusion >>
rect 355 503 356 504 
<< pdiffusion >>
rect 356 503 357 504 
<< pdiffusion >>
rect 357 503 358 504 
<< pdiffusion >>
rect 358 503 359 504 
<< pdiffusion >>
rect 359 503 360 504 
<< m1 >>
rect 361 503 362 504 
<< pdiffusion >>
rect 372 503 373 504 
<< pdiffusion >>
rect 373 503 374 504 
<< pdiffusion >>
rect 374 503 375 504 
<< pdiffusion >>
rect 375 503 376 504 
<< pdiffusion >>
rect 376 503 377 504 
<< pdiffusion >>
rect 377 503 378 504 
<< m1 >>
rect 379 503 380 504 
<< m1 >>
rect 381 503 382 504 
<< m2 >>
rect 382 503 383 504 
<< pdiffusion >>
rect 390 503 391 504 
<< pdiffusion >>
rect 391 503 392 504 
<< pdiffusion >>
rect 392 503 393 504 
<< pdiffusion >>
rect 393 503 394 504 
<< pdiffusion >>
rect 394 503 395 504 
<< pdiffusion >>
rect 395 503 396 504 
<< m1 >>
rect 406 503 407 504 
<< pdiffusion >>
rect 408 503 409 504 
<< m1 >>
rect 409 503 410 504 
<< pdiffusion >>
rect 409 503 410 504 
<< pdiffusion >>
rect 410 503 411 504 
<< pdiffusion >>
rect 411 503 412 504 
<< pdiffusion >>
rect 412 503 413 504 
<< pdiffusion >>
rect 413 503 414 504 
<< pdiffusion >>
rect 444 503 445 504 
<< pdiffusion >>
rect 445 503 446 504 
<< pdiffusion >>
rect 446 503 447 504 
<< pdiffusion >>
rect 447 503 448 504 
<< pdiffusion >>
rect 448 503 449 504 
<< pdiffusion >>
rect 449 503 450 504 
<< m1 >>
rect 451 503 452 504 
<< pdiffusion >>
rect 462 503 463 504 
<< pdiffusion >>
rect 463 503 464 504 
<< pdiffusion >>
rect 464 503 465 504 
<< pdiffusion >>
rect 465 503 466 504 
<< pdiffusion >>
rect 466 503 467 504 
<< pdiffusion >>
rect 467 503 468 504 
<< m1 >>
rect 472 503 473 504 
<< pdiffusion >>
rect 480 503 481 504 
<< pdiffusion >>
rect 481 503 482 504 
<< pdiffusion >>
rect 482 503 483 504 
<< pdiffusion >>
rect 483 503 484 504 
<< pdiffusion >>
rect 484 503 485 504 
<< pdiffusion >>
rect 485 503 486 504 
<< m1 >>
rect 487 503 488 504 
<< m1 >>
rect 489 503 490 504 
<< pdiffusion >>
rect 498 503 499 504 
<< pdiffusion >>
rect 499 503 500 504 
<< pdiffusion >>
rect 500 503 501 504 
<< pdiffusion >>
rect 501 503 502 504 
<< m1 >>
rect 502 503 503 504 
<< pdiffusion >>
rect 502 503 503 504 
<< pdiffusion >>
rect 503 503 504 504 
<< pdiffusion >>
rect 516 503 517 504 
<< pdiffusion >>
rect 517 503 518 504 
<< pdiffusion >>
rect 518 503 519 504 
<< pdiffusion >>
rect 519 503 520 504 
<< m1 >>
rect 520 503 521 504 
<< pdiffusion >>
rect 520 503 521 504 
<< pdiffusion >>
rect 521 503 522 504 
<< m1 >>
rect 523 503 524 504 
<< m1 >>
rect 13 504 14 505 
<< m1 >>
rect 28 504 29 505 
<< m1 >>
rect 37 504 38 505 
<< m1 >>
rect 49 504 50 505 
<< m1 >>
rect 73 504 74 505 
<< m1 >>
rect 100 504 101 505 
<< m1 >>
rect 118 504 119 505 
<< m1 >>
rect 142 504 143 505 
<< m1 >>
rect 186 504 187 505 
<< m1 >>
rect 190 504 191 505 
<< m1 >>
rect 250 504 251 505 
<< m1 >>
rect 253 504 254 505 
<< m1 >>
rect 319 504 320 505 
<< m1 >>
rect 361 504 362 505 
<< m1 >>
rect 379 504 380 505 
<< m1 >>
rect 381 504 382 505 
<< m2 >>
rect 382 504 383 505 
<< m1 >>
rect 406 504 407 505 
<< m1 >>
rect 409 504 410 505 
<< m1 >>
rect 451 504 452 505 
<< m1 >>
rect 472 504 473 505 
<< m1 >>
rect 487 504 488 505 
<< m1 >>
rect 489 504 490 505 
<< m1 >>
rect 502 504 503 505 
<< m1 >>
rect 520 504 521 505 
<< m1 >>
rect 523 504 524 505 
<< m1 >>
rect 13 505 14 506 
<< m1 >>
rect 28 505 29 506 
<< m1 >>
rect 37 505 38 506 
<< m1 >>
rect 38 505 39 506 
<< m1 >>
rect 39 505 40 506 
<< m1 >>
rect 40 505 41 506 
<< m1 >>
rect 41 505 42 506 
<< m1 >>
rect 42 505 43 506 
<< m1 >>
rect 43 505 44 506 
<< m1 >>
rect 44 505 45 506 
<< m1 >>
rect 45 505 46 506 
<< m1 >>
rect 46 505 47 506 
<< m1 >>
rect 47 505 48 506 
<< m1 >>
rect 48 505 49 506 
<< m1 >>
rect 49 505 50 506 
<< m1 >>
rect 73 505 74 506 
<< m1 >>
rect 100 505 101 506 
<< m1 >>
rect 118 505 119 506 
<< m1 >>
rect 142 505 143 506 
<< m1 >>
rect 186 505 187 506 
<< m1 >>
rect 190 505 191 506 
<< m1 >>
rect 250 505 251 506 
<< m1 >>
rect 251 505 252 506 
<< m1 >>
rect 252 505 253 506 
<< m1 >>
rect 253 505 254 506 
<< m1 >>
rect 319 505 320 506 
<< m1 >>
rect 361 505 362 506 
<< m1 >>
rect 377 505 378 506 
<< m2 >>
rect 377 505 378 506 
<< m2c >>
rect 377 505 378 506 
<< m1 >>
rect 377 505 378 506 
<< m2 >>
rect 377 505 378 506 
<< m2 >>
rect 378 505 379 506 
<< m1 >>
rect 379 505 380 506 
<< m2 >>
rect 379 505 380 506 
<< m2 >>
rect 380 505 381 506 
<< m1 >>
rect 381 505 382 506 
<< m2 >>
rect 381 505 382 506 
<< m2 >>
rect 382 505 383 506 
<< m1 >>
rect 406 505 407 506 
<< m1 >>
rect 407 505 408 506 
<< m1 >>
rect 408 505 409 506 
<< m1 >>
rect 409 505 410 506 
<< m1 >>
rect 451 505 452 506 
<< m1 >>
rect 472 505 473 506 
<< m1 >>
rect 487 505 488 506 
<< m1 >>
rect 489 505 490 506 
<< m1 >>
rect 502 505 503 506 
<< m1 >>
rect 520 505 521 506 
<< m1 >>
rect 521 505 522 506 
<< m1 >>
rect 522 505 523 506 
<< m1 >>
rect 523 505 524 506 
<< m1 >>
rect 13 506 14 507 
<< m1 >>
rect 14 506 15 507 
<< m1 >>
rect 15 506 16 507 
<< m1 >>
rect 16 506 17 507 
<< m1 >>
rect 17 506 18 507 
<< m1 >>
rect 18 506 19 507 
<< m1 >>
rect 19 506 20 507 
<< m1 >>
rect 20 506 21 507 
<< m1 >>
rect 21 506 22 507 
<< m1 >>
rect 22 506 23 507 
<< m1 >>
rect 23 506 24 507 
<< m1 >>
rect 24 506 25 507 
<< m1 >>
rect 25 506 26 507 
<< m1 >>
rect 26 506 27 507 
<< m1 >>
rect 27 506 28 507 
<< m1 >>
rect 28 506 29 507 
<< m1 >>
rect 70 506 71 507 
<< m1 >>
rect 71 506 72 507 
<< m1 >>
rect 72 506 73 507 
<< m1 >>
rect 73 506 74 507 
<< m1 >>
rect 100 506 101 507 
<< m1 >>
rect 118 506 119 507 
<< m1 >>
rect 142 506 143 507 
<< m1 >>
rect 186 506 187 507 
<< m1 >>
rect 190 506 191 507 
<< m1 >>
rect 319 506 320 507 
<< m1 >>
rect 361 506 362 507 
<< m1 >>
rect 377 506 378 507 
<< m1 >>
rect 379 506 380 507 
<< m1 >>
rect 381 506 382 507 
<< m1 >>
rect 451 506 452 507 
<< m1 >>
rect 472 506 473 507 
<< m1 >>
rect 487 506 488 507 
<< m1 >>
rect 489 506 490 507 
<< m1 >>
rect 502 506 503 507 
<< m1 >>
rect 70 507 71 508 
<< m1 >>
rect 100 507 101 508 
<< m1 >>
rect 118 507 119 508 
<< m1 >>
rect 142 507 143 508 
<< m1 >>
rect 186 507 187 508 
<< m1 >>
rect 190 507 191 508 
<< m1 >>
rect 319 507 320 508 
<< m1 >>
rect 361 507 362 508 
<< m1 >>
rect 377 507 378 508 
<< m1 >>
rect 379 507 380 508 
<< m1 >>
rect 381 507 382 508 
<< m1 >>
rect 451 507 452 508 
<< m1 >>
rect 472 507 473 508 
<< m1 >>
rect 487 507 488 508 
<< m1 >>
rect 489 507 490 508 
<< m1 >>
rect 502 507 503 508 
<< m1 >>
rect 70 508 71 509 
<< m1 >>
rect 100 508 101 509 
<< m1 >>
rect 118 508 119 509 
<< m1 >>
rect 124 508 125 509 
<< m1 >>
rect 125 508 126 509 
<< m1 >>
rect 126 508 127 509 
<< m1 >>
rect 127 508 128 509 
<< m1 >>
rect 128 508 129 509 
<< m1 >>
rect 129 508 130 509 
<< m1 >>
rect 130 508 131 509 
<< m1 >>
rect 131 508 132 509 
<< m1 >>
rect 132 508 133 509 
<< m1 >>
rect 133 508 134 509 
<< m1 >>
rect 134 508 135 509 
<< m1 >>
rect 135 508 136 509 
<< m1 >>
rect 136 508 137 509 
<< m1 >>
rect 137 508 138 509 
<< m1 >>
rect 138 508 139 509 
<< m1 >>
rect 139 508 140 509 
<< m1 >>
rect 140 508 141 509 
<< m1 >>
rect 141 508 142 509 
<< m1 >>
rect 142 508 143 509 
<< m1 >>
rect 186 508 187 509 
<< m1 >>
rect 190 508 191 509 
<< m1 >>
rect 319 508 320 509 
<< m1 >>
rect 361 508 362 509 
<< m1 >>
rect 377 508 378 509 
<< m1 >>
rect 379 508 380 509 
<< m1 >>
rect 381 508 382 509 
<< m1 >>
rect 451 508 452 509 
<< m1 >>
rect 472 508 473 509 
<< m1 >>
rect 487 508 488 509 
<< m1 >>
rect 489 508 490 509 
<< m1 >>
rect 490 508 491 509 
<< m1 >>
rect 491 508 492 509 
<< m1 >>
rect 492 508 493 509 
<< m1 >>
rect 493 508 494 509 
<< m1 >>
rect 494 508 495 509 
<< m1 >>
rect 495 508 496 509 
<< m1 >>
rect 496 508 497 509 
<< m1 >>
rect 497 508 498 509 
<< m1 >>
rect 498 508 499 509 
<< m1 >>
rect 499 508 500 509 
<< m1 >>
rect 500 508 501 509 
<< m1 >>
rect 501 508 502 509 
<< m1 >>
rect 502 508 503 509 
<< m1 >>
rect 70 509 71 510 
<< m1 >>
rect 100 509 101 510 
<< m1 >>
rect 118 509 119 510 
<< m1 >>
rect 124 509 125 510 
<< m1 >>
rect 186 509 187 510 
<< m2 >>
rect 186 509 187 510 
<< m2c >>
rect 186 509 187 510 
<< m1 >>
rect 186 509 187 510 
<< m2 >>
rect 186 509 187 510 
<< m1 >>
rect 190 509 191 510 
<< m1 >>
rect 319 509 320 510 
<< m2 >>
rect 319 509 320 510 
<< m2c >>
rect 319 509 320 510 
<< m1 >>
rect 319 509 320 510 
<< m2 >>
rect 319 509 320 510 
<< m1 >>
rect 361 509 362 510 
<< m2 >>
rect 361 509 362 510 
<< m2c >>
rect 361 509 362 510 
<< m1 >>
rect 361 509 362 510 
<< m2 >>
rect 361 509 362 510 
<< m1 >>
rect 377 509 378 510 
<< m2 >>
rect 377 509 378 510 
<< m2c >>
rect 377 509 378 510 
<< m1 >>
rect 377 509 378 510 
<< m2 >>
rect 377 509 378 510 
<< m1 >>
rect 379 509 380 510 
<< m2 >>
rect 379 509 380 510 
<< m2c >>
rect 379 509 380 510 
<< m1 >>
rect 379 509 380 510 
<< m2 >>
rect 379 509 380 510 
<< m1 >>
rect 381 509 382 510 
<< m2 >>
rect 381 509 382 510 
<< m2c >>
rect 381 509 382 510 
<< m1 >>
rect 381 509 382 510 
<< m2 >>
rect 381 509 382 510 
<< m1 >>
rect 451 509 452 510 
<< m2 >>
rect 451 509 452 510 
<< m2c >>
rect 451 509 452 510 
<< m1 >>
rect 451 509 452 510 
<< m2 >>
rect 451 509 452 510 
<< m1 >>
rect 472 509 473 510 
<< m2 >>
rect 472 509 473 510 
<< m2c >>
rect 472 509 473 510 
<< m1 >>
rect 472 509 473 510 
<< m2 >>
rect 472 509 473 510 
<< m1 >>
rect 487 509 488 510 
<< m1 >>
rect 70 510 71 511 
<< m1 >>
rect 100 510 101 511 
<< m1 >>
rect 118 510 119 511 
<< m1 >>
rect 124 510 125 511 
<< m2 >>
rect 186 510 187 511 
<< m1 >>
rect 190 510 191 511 
<< m2 >>
rect 319 510 320 511 
<< m2 >>
rect 320 510 321 511 
<< m2 >>
rect 361 510 362 511 
<< m2 >>
rect 372 510 373 511 
<< m2 >>
rect 373 510 374 511 
<< m2 >>
rect 374 510 375 511 
<< m2 >>
rect 375 510 376 511 
<< m2 >>
rect 376 510 377 511 
<< m2 >>
rect 377 510 378 511 
<< m2 >>
rect 379 510 380 511 
<< m2 >>
rect 381 510 382 511 
<< m2 >>
rect 382 510 383 511 
<< m2 >>
rect 383 510 384 511 
<< m2 >>
rect 384 510 385 511 
<< m2 >>
rect 385 510 386 511 
<< m2 >>
rect 386 510 387 511 
<< m2 >>
rect 387 510 388 511 
<< m2 >>
rect 388 510 389 511 
<< m2 >>
rect 389 510 390 511 
<< m2 >>
rect 390 510 391 511 
<< m2 >>
rect 391 510 392 511 
<< m2 >>
rect 392 510 393 511 
<< m2 >>
rect 393 510 394 511 
<< m2 >>
rect 394 510 395 511 
<< m2 >>
rect 395 510 396 511 
<< m2 >>
rect 396 510 397 511 
<< m2 >>
rect 397 510 398 511 
<< m2 >>
rect 398 510 399 511 
<< m2 >>
rect 399 510 400 511 
<< m2 >>
rect 400 510 401 511 
<< m2 >>
rect 401 510 402 511 
<< m2 >>
rect 402 510 403 511 
<< m2 >>
rect 403 510 404 511 
<< m2 >>
rect 404 510 405 511 
<< m2 >>
rect 405 510 406 511 
<< m2 >>
rect 406 510 407 511 
<< m2 >>
rect 407 510 408 511 
<< m2 >>
rect 408 510 409 511 
<< m2 >>
rect 409 510 410 511 
<< m2 >>
rect 410 510 411 511 
<< m2 >>
rect 411 510 412 511 
<< m2 >>
rect 412 510 413 511 
<< m2 >>
rect 413 510 414 511 
<< m2 >>
rect 414 510 415 511 
<< m2 >>
rect 415 510 416 511 
<< m2 >>
rect 416 510 417 511 
<< m2 >>
rect 417 510 418 511 
<< m2 >>
rect 418 510 419 511 
<< m2 >>
rect 419 510 420 511 
<< m2 >>
rect 420 510 421 511 
<< m2 >>
rect 421 510 422 511 
<< m2 >>
rect 422 510 423 511 
<< m2 >>
rect 423 510 424 511 
<< m2 >>
rect 424 510 425 511 
<< m2 >>
rect 425 510 426 511 
<< m2 >>
rect 426 510 427 511 
<< m2 >>
rect 427 510 428 511 
<< m2 >>
rect 428 510 429 511 
<< m2 >>
rect 429 510 430 511 
<< m2 >>
rect 430 510 431 511 
<< m2 >>
rect 431 510 432 511 
<< m2 >>
rect 432 510 433 511 
<< m2 >>
rect 433 510 434 511 
<< m2 >>
rect 434 510 435 511 
<< m2 >>
rect 435 510 436 511 
<< m2 >>
rect 436 510 437 511 
<< m2 >>
rect 437 510 438 511 
<< m2 >>
rect 438 510 439 511 
<< m2 >>
rect 439 510 440 511 
<< m2 >>
rect 440 510 441 511 
<< m2 >>
rect 441 510 442 511 
<< m2 >>
rect 442 510 443 511 
<< m2 >>
rect 443 510 444 511 
<< m2 >>
rect 444 510 445 511 
<< m2 >>
rect 445 510 446 511 
<< m2 >>
rect 446 510 447 511 
<< m2 >>
rect 451 510 452 511 
<< m2 >>
rect 472 510 473 511 
<< m1 >>
rect 487 510 488 511 
<< m1 >>
rect 19 511 20 512 
<< m1 >>
rect 20 511 21 512 
<< m1 >>
rect 21 511 22 512 
<< m1 >>
rect 22 511 23 512 
<< m1 >>
rect 23 511 24 512 
<< m1 >>
rect 24 511 25 512 
<< m1 >>
rect 25 511 26 512 
<< m1 >>
rect 26 511 27 512 
<< m1 >>
rect 27 511 28 512 
<< m1 >>
rect 28 511 29 512 
<< m1 >>
rect 29 511 30 512 
<< m1 >>
rect 30 511 31 512 
<< m1 >>
rect 31 511 32 512 
<< m1 >>
rect 32 511 33 512 
<< m1 >>
rect 33 511 34 512 
<< m1 >>
rect 34 511 35 512 
<< m1 >>
rect 70 511 71 512 
<< m1 >>
rect 100 511 101 512 
<< m1 >>
rect 118 511 119 512 
<< m1 >>
rect 119 511 120 512 
<< m1 >>
rect 120 511 121 512 
<< m1 >>
rect 121 511 122 512 
<< m1 >>
rect 122 511 123 512 
<< m2 >>
rect 122 511 123 512 
<< m2c >>
rect 122 511 123 512 
<< m1 >>
rect 122 511 123 512 
<< m2 >>
rect 122 511 123 512 
<< m2 >>
rect 123 511 124 512 
<< m1 >>
rect 124 511 125 512 
<< m2 >>
rect 124 511 125 512 
<< m2 >>
rect 125 511 126 512 
<< m1 >>
rect 126 511 127 512 
<< m2 >>
rect 126 511 127 512 
<< m2c >>
rect 126 511 127 512 
<< m1 >>
rect 126 511 127 512 
<< m2 >>
rect 126 511 127 512 
<< m1 >>
rect 127 511 128 512 
<< m1 >>
rect 128 511 129 512 
<< m1 >>
rect 129 511 130 512 
<< m1 >>
rect 130 511 131 512 
<< m1 >>
rect 131 511 132 512 
<< m1 >>
rect 132 511 133 512 
<< m1 >>
rect 133 511 134 512 
<< m1 >>
rect 134 511 135 512 
<< m1 >>
rect 135 511 136 512 
<< m1 >>
rect 136 511 137 512 
<< m1 >>
rect 137 511 138 512 
<< m1 >>
rect 138 511 139 512 
<< m1 >>
rect 139 511 140 512 
<< m1 >>
rect 140 511 141 512 
<< m1 >>
rect 141 511 142 512 
<< m1 >>
rect 142 511 143 512 
<< m1 >>
rect 143 511 144 512 
<< m1 >>
rect 144 511 145 512 
<< m1 >>
rect 145 511 146 512 
<< m1 >>
rect 146 511 147 512 
<< m1 >>
rect 147 511 148 512 
<< m1 >>
rect 148 511 149 512 
<< m1 >>
rect 149 511 150 512 
<< m1 >>
rect 150 511 151 512 
<< m1 >>
rect 151 511 152 512 
<< m1 >>
rect 152 511 153 512 
<< m1 >>
rect 153 511 154 512 
<< m1 >>
rect 154 511 155 512 
<< m1 >>
rect 155 511 156 512 
<< m1 >>
rect 156 511 157 512 
<< m1 >>
rect 157 511 158 512 
<< m1 >>
rect 158 511 159 512 
<< m1 >>
rect 159 511 160 512 
<< m1 >>
rect 160 511 161 512 
<< m1 >>
rect 161 511 162 512 
<< m1 >>
rect 162 511 163 512 
<< m1 >>
rect 163 511 164 512 
<< m1 >>
rect 164 511 165 512 
<< m1 >>
rect 165 511 166 512 
<< m1 >>
rect 166 511 167 512 
<< m1 >>
rect 167 511 168 512 
<< m1 >>
rect 168 511 169 512 
<< m1 >>
rect 169 511 170 512 
<< m1 >>
rect 170 511 171 512 
<< m1 >>
rect 171 511 172 512 
<< m1 >>
rect 172 511 173 512 
<< m1 >>
rect 173 511 174 512 
<< m1 >>
rect 174 511 175 512 
<< m1 >>
rect 175 511 176 512 
<< m1 >>
rect 176 511 177 512 
<< m1 >>
rect 177 511 178 512 
<< m1 >>
rect 178 511 179 512 
<< m1 >>
rect 179 511 180 512 
<< m1 >>
rect 180 511 181 512 
<< m1 >>
rect 181 511 182 512 
<< m1 >>
rect 182 511 183 512 
<< m1 >>
rect 183 511 184 512 
<< m1 >>
rect 184 511 185 512 
<< m1 >>
rect 185 511 186 512 
<< m1 >>
rect 186 511 187 512 
<< m2 >>
rect 186 511 187 512 
<< m1 >>
rect 187 511 188 512 
<< m1 >>
rect 188 511 189 512 
<< m2 >>
rect 188 511 189 512 
<< m2c >>
rect 188 511 189 512 
<< m1 >>
rect 188 511 189 512 
<< m2 >>
rect 188 511 189 512 
<< m2 >>
rect 189 511 190 512 
<< m1 >>
rect 190 511 191 512 
<< m2 >>
rect 190 511 191 512 
<< m1 >>
rect 191 511 192 512 
<< m2 >>
rect 191 511 192 512 
<< m1 >>
rect 192 511 193 512 
<< m2 >>
rect 192 511 193 512 
<< m1 >>
rect 193 511 194 512 
<< m2 >>
rect 193 511 194 512 
<< m1 >>
rect 194 511 195 512 
<< m2 >>
rect 194 511 195 512 
<< m1 >>
rect 195 511 196 512 
<< m2 >>
rect 195 511 196 512 
<< m1 >>
rect 196 511 197 512 
<< m2 >>
rect 196 511 197 512 
<< m1 >>
rect 197 511 198 512 
<< m2 >>
rect 197 511 198 512 
<< m1 >>
rect 198 511 199 512 
<< m2 >>
rect 198 511 199 512 
<< m1 >>
rect 199 511 200 512 
<< m2 >>
rect 199 511 200 512 
<< m1 >>
rect 200 511 201 512 
<< m2 >>
rect 200 511 201 512 
<< m1 >>
rect 201 511 202 512 
<< m2 >>
rect 201 511 202 512 
<< m1 >>
rect 202 511 203 512 
<< m2 >>
rect 202 511 203 512 
<< m1 >>
rect 203 511 204 512 
<< m2 >>
rect 203 511 204 512 
<< m1 >>
rect 204 511 205 512 
<< m2 >>
rect 204 511 205 512 
<< m1 >>
rect 205 511 206 512 
<< m2 >>
rect 205 511 206 512 
<< m1 >>
rect 206 511 207 512 
<< m2 >>
rect 206 511 207 512 
<< m1 >>
rect 207 511 208 512 
<< m2 >>
rect 207 511 208 512 
<< m1 >>
rect 208 511 209 512 
<< m2 >>
rect 208 511 209 512 
<< m1 >>
rect 209 511 210 512 
<< m2 >>
rect 209 511 210 512 
<< m1 >>
rect 210 511 211 512 
<< m2 >>
rect 210 511 211 512 
<< m1 >>
rect 211 511 212 512 
<< m2 >>
rect 211 511 212 512 
<< m1 >>
rect 212 511 213 512 
<< m2 >>
rect 212 511 213 512 
<< m1 >>
rect 213 511 214 512 
<< m2 >>
rect 213 511 214 512 
<< m1 >>
rect 214 511 215 512 
<< m2 >>
rect 214 511 215 512 
<< m1 >>
rect 215 511 216 512 
<< m2 >>
rect 215 511 216 512 
<< m1 >>
rect 216 511 217 512 
<< m2 >>
rect 216 511 217 512 
<< m1 >>
rect 217 511 218 512 
<< m2 >>
rect 217 511 218 512 
<< m1 >>
rect 218 511 219 512 
<< m2 >>
rect 218 511 219 512 
<< m1 >>
rect 219 511 220 512 
<< m2 >>
rect 219 511 220 512 
<< m1 >>
rect 220 511 221 512 
<< m2 >>
rect 220 511 221 512 
<< m1 >>
rect 221 511 222 512 
<< m2 >>
rect 221 511 222 512 
<< m1 >>
rect 222 511 223 512 
<< m2 >>
rect 222 511 223 512 
<< m1 >>
rect 223 511 224 512 
<< m2 >>
rect 223 511 224 512 
<< m1 >>
rect 224 511 225 512 
<< m2 >>
rect 224 511 225 512 
<< m1 >>
rect 225 511 226 512 
<< m2 >>
rect 225 511 226 512 
<< m1 >>
rect 226 511 227 512 
<< m2 >>
rect 226 511 227 512 
<< m2 >>
rect 227 511 228 512 
<< m1 >>
rect 228 511 229 512 
<< m2 >>
rect 228 511 229 512 
<< m2c >>
rect 228 511 229 512 
<< m1 >>
rect 228 511 229 512 
<< m2 >>
rect 228 511 229 512 
<< m1 >>
rect 229 511 230 512 
<< m1 >>
rect 230 511 231 512 
<< m1 >>
rect 231 511 232 512 
<< m1 >>
rect 232 511 233 512 
<< m1 >>
rect 233 511 234 512 
<< m1 >>
rect 234 511 235 512 
<< m1 >>
rect 235 511 236 512 
<< m1 >>
rect 236 511 237 512 
<< m1 >>
rect 237 511 238 512 
<< m1 >>
rect 238 511 239 512 
<< m1 >>
rect 239 511 240 512 
<< m1 >>
rect 240 511 241 512 
<< m1 >>
rect 241 511 242 512 
<< m1 >>
rect 242 511 243 512 
<< m1 >>
rect 243 511 244 512 
<< m1 >>
rect 244 511 245 512 
<< m1 >>
rect 245 511 246 512 
<< m1 >>
rect 246 511 247 512 
<< m1 >>
rect 247 511 248 512 
<< m1 >>
rect 248 511 249 512 
<< m1 >>
rect 249 511 250 512 
<< m1 >>
rect 250 511 251 512 
<< m1 >>
rect 251 511 252 512 
<< m1 >>
rect 252 511 253 512 
<< m1 >>
rect 253 511 254 512 
<< m1 >>
rect 254 511 255 512 
<< m1 >>
rect 255 511 256 512 
<< m1 >>
rect 256 511 257 512 
<< m1 >>
rect 257 511 258 512 
<< m1 >>
rect 258 511 259 512 
<< m1 >>
rect 259 511 260 512 
<< m1 >>
rect 260 511 261 512 
<< m1 >>
rect 261 511 262 512 
<< m1 >>
rect 262 511 263 512 
<< m1 >>
rect 268 511 269 512 
<< m1 >>
rect 269 511 270 512 
<< m1 >>
rect 270 511 271 512 
<< m1 >>
rect 271 511 272 512 
<< m1 >>
rect 272 511 273 512 
<< m1 >>
rect 273 511 274 512 
<< m1 >>
rect 274 511 275 512 
<< m1 >>
rect 275 511 276 512 
<< m1 >>
rect 276 511 277 512 
<< m1 >>
rect 277 511 278 512 
<< m1 >>
rect 278 511 279 512 
<< m1 >>
rect 279 511 280 512 
<< m1 >>
rect 280 511 281 512 
<< m1 >>
rect 281 511 282 512 
<< m1 >>
rect 282 511 283 512 
<< m1 >>
rect 283 511 284 512 
<< m1 >>
rect 284 511 285 512 
<< m1 >>
rect 285 511 286 512 
<< m1 >>
rect 286 511 287 512 
<< m1 >>
rect 287 511 288 512 
<< m1 >>
rect 288 511 289 512 
<< m1 >>
rect 289 511 290 512 
<< m1 >>
rect 290 511 291 512 
<< m1 >>
rect 291 511 292 512 
<< m1 >>
rect 292 511 293 512 
<< m1 >>
rect 293 511 294 512 
<< m1 >>
rect 294 511 295 512 
<< m1 >>
rect 295 511 296 512 
<< m1 >>
rect 296 511 297 512 
<< m1 >>
rect 297 511 298 512 
<< m1 >>
rect 298 511 299 512 
<< m1 >>
rect 299 511 300 512 
<< m1 >>
rect 300 511 301 512 
<< m1 >>
rect 301 511 302 512 
<< m1 >>
rect 302 511 303 512 
<< m1 >>
rect 303 511 304 512 
<< m1 >>
rect 304 511 305 512 
<< m1 >>
rect 305 511 306 512 
<< m1 >>
rect 306 511 307 512 
<< m1 >>
rect 307 511 308 512 
<< m1 >>
rect 308 511 309 512 
<< m1 >>
rect 309 511 310 512 
<< m1 >>
rect 310 511 311 512 
<< m1 >>
rect 311 511 312 512 
<< m1 >>
rect 312 511 313 512 
<< m1 >>
rect 313 511 314 512 
<< m1 >>
rect 314 511 315 512 
<< m1 >>
rect 315 511 316 512 
<< m1 >>
rect 316 511 317 512 
<< m1 >>
rect 317 511 318 512 
<< m1 >>
rect 318 511 319 512 
<< m1 >>
rect 319 511 320 512 
<< m1 >>
rect 320 511 321 512 
<< m2 >>
rect 320 511 321 512 
<< m1 >>
rect 321 511 322 512 
<< m1 >>
rect 322 511 323 512 
<< m1 >>
rect 323 511 324 512 
<< m1 >>
rect 324 511 325 512 
<< m1 >>
rect 325 511 326 512 
<< m1 >>
rect 326 511 327 512 
<< m1 >>
rect 327 511 328 512 
<< m1 >>
rect 328 511 329 512 
<< m1 >>
rect 329 511 330 512 
<< m1 >>
rect 330 511 331 512 
<< m1 >>
rect 331 511 332 512 
<< m1 >>
rect 332 511 333 512 
<< m1 >>
rect 333 511 334 512 
<< m1 >>
rect 334 511 335 512 
<< m1 >>
rect 335 511 336 512 
<< m1 >>
rect 336 511 337 512 
<< m1 >>
rect 337 511 338 512 
<< m1 >>
rect 338 511 339 512 
<< m1 >>
rect 339 511 340 512 
<< m1 >>
rect 340 511 341 512 
<< m1 >>
rect 341 511 342 512 
<< m1 >>
rect 342 511 343 512 
<< m1 >>
rect 343 511 344 512 
<< m1 >>
rect 344 511 345 512 
<< m1 >>
rect 345 511 346 512 
<< m1 >>
rect 346 511 347 512 
<< m1 >>
rect 347 511 348 512 
<< m1 >>
rect 348 511 349 512 
<< m1 >>
rect 349 511 350 512 
<< m1 >>
rect 350 511 351 512 
<< m1 >>
rect 351 511 352 512 
<< m1 >>
rect 352 511 353 512 
<< m1 >>
rect 353 511 354 512 
<< m1 >>
rect 354 511 355 512 
<< m1 >>
rect 355 511 356 512 
<< m1 >>
rect 356 511 357 512 
<< m1 >>
rect 357 511 358 512 
<< m1 >>
rect 358 511 359 512 
<< m1 >>
rect 359 511 360 512 
<< m1 >>
rect 360 511 361 512 
<< m1 >>
rect 361 511 362 512 
<< m2 >>
rect 361 511 362 512 
<< m1 >>
rect 362 511 363 512 
<< m1 >>
rect 363 511 364 512 
<< m1 >>
rect 364 511 365 512 
<< m1 >>
rect 365 511 366 512 
<< m1 >>
rect 366 511 367 512 
<< m1 >>
rect 367 511 368 512 
<< m1 >>
rect 368 511 369 512 
<< m1 >>
rect 369 511 370 512 
<< m1 >>
rect 370 511 371 512 
<< m1 >>
rect 371 511 372 512 
<< m1 >>
rect 372 511 373 512 
<< m2 >>
rect 372 511 373 512 
<< m1 >>
rect 373 511 374 512 
<< m1 >>
rect 374 511 375 512 
<< m1 >>
rect 375 511 376 512 
<< m1 >>
rect 376 511 377 512 
<< m1 >>
rect 377 511 378 512 
<< m1 >>
rect 378 511 379 512 
<< m1 >>
rect 379 511 380 512 
<< m2 >>
rect 379 511 380 512 
<< m1 >>
rect 380 511 381 512 
<< m1 >>
rect 381 511 382 512 
<< m1 >>
rect 382 511 383 512 
<< m1 >>
rect 383 511 384 512 
<< m1 >>
rect 384 511 385 512 
<< m1 >>
rect 385 511 386 512 
<< m1 >>
rect 386 511 387 512 
<< m1 >>
rect 387 511 388 512 
<< m1 >>
rect 388 511 389 512 
<< m1 >>
rect 389 511 390 512 
<< m1 >>
rect 390 511 391 512 
<< m1 >>
rect 391 511 392 512 
<< m1 >>
rect 392 511 393 512 
<< m1 >>
rect 393 511 394 512 
<< m1 >>
rect 394 511 395 512 
<< m1 >>
rect 395 511 396 512 
<< m1 >>
rect 396 511 397 512 
<< m1 >>
rect 397 511 398 512 
<< m1 >>
rect 398 511 399 512 
<< m1 >>
rect 399 511 400 512 
<< m1 >>
rect 400 511 401 512 
<< m1 >>
rect 401 511 402 512 
<< m1 >>
rect 402 511 403 512 
<< m1 >>
rect 403 511 404 512 
<< m1 >>
rect 404 511 405 512 
<< m1 >>
rect 405 511 406 512 
<< m1 >>
rect 406 511 407 512 
<< m1 >>
rect 407 511 408 512 
<< m1 >>
rect 408 511 409 512 
<< m1 >>
rect 409 511 410 512 
<< m1 >>
rect 410 511 411 512 
<< m1 >>
rect 411 511 412 512 
<< m1 >>
rect 412 511 413 512 
<< m1 >>
rect 413 511 414 512 
<< m1 >>
rect 414 511 415 512 
<< m1 >>
rect 415 511 416 512 
<< m1 >>
rect 416 511 417 512 
<< m1 >>
rect 417 511 418 512 
<< m1 >>
rect 418 511 419 512 
<< m1 >>
rect 419 511 420 512 
<< m1 >>
rect 420 511 421 512 
<< m1 >>
rect 421 511 422 512 
<< m1 >>
rect 422 511 423 512 
<< m1 >>
rect 423 511 424 512 
<< m1 >>
rect 424 511 425 512 
<< m1 >>
rect 425 511 426 512 
<< m1 >>
rect 426 511 427 512 
<< m1 >>
rect 427 511 428 512 
<< m1 >>
rect 428 511 429 512 
<< m1 >>
rect 429 511 430 512 
<< m1 >>
rect 430 511 431 512 
<< m1 >>
rect 431 511 432 512 
<< m1 >>
rect 432 511 433 512 
<< m1 >>
rect 433 511 434 512 
<< m1 >>
rect 434 511 435 512 
<< m1 >>
rect 435 511 436 512 
<< m1 >>
rect 436 511 437 512 
<< m1 >>
rect 437 511 438 512 
<< m1 >>
rect 438 511 439 512 
<< m1 >>
rect 439 511 440 512 
<< m1 >>
rect 440 511 441 512 
<< m1 >>
rect 441 511 442 512 
<< m1 >>
rect 442 511 443 512 
<< m1 >>
rect 443 511 444 512 
<< m1 >>
rect 444 511 445 512 
<< m1 >>
rect 445 511 446 512 
<< m1 >>
rect 446 511 447 512 
<< m2 >>
rect 446 511 447 512 
<< m1 >>
rect 447 511 448 512 
<< m1 >>
rect 448 511 449 512 
<< m1 >>
rect 449 511 450 512 
<< m1 >>
rect 450 511 451 512 
<< m1 >>
rect 451 511 452 512 
<< m2 >>
rect 451 511 452 512 
<< m1 >>
rect 452 511 453 512 
<< m1 >>
rect 453 511 454 512 
<< m1 >>
rect 454 511 455 512 
<< m1 >>
rect 455 511 456 512 
<< m1 >>
rect 456 511 457 512 
<< m1 >>
rect 457 511 458 512 
<< m1 >>
rect 458 511 459 512 
<< m1 >>
rect 459 511 460 512 
<< m1 >>
rect 460 511 461 512 
<< m1 >>
rect 461 511 462 512 
<< m1 >>
rect 462 511 463 512 
<< m1 >>
rect 463 511 464 512 
<< m1 >>
rect 464 511 465 512 
<< m1 >>
rect 465 511 466 512 
<< m1 >>
rect 466 511 467 512 
<< m1 >>
rect 467 511 468 512 
<< m1 >>
rect 468 511 469 512 
<< m1 >>
rect 469 511 470 512 
<< m1 >>
rect 470 511 471 512 
<< m1 >>
rect 471 511 472 512 
<< m1 >>
rect 472 511 473 512 
<< m2 >>
rect 472 511 473 512 
<< m1 >>
rect 473 511 474 512 
<< m1 >>
rect 474 511 475 512 
<< m1 >>
rect 475 511 476 512 
<< m1 >>
rect 476 511 477 512 
<< m1 >>
rect 477 511 478 512 
<< m1 >>
rect 478 511 479 512 
<< m1 >>
rect 479 511 480 512 
<< m1 >>
rect 480 511 481 512 
<< m1 >>
rect 481 511 482 512 
<< m1 >>
rect 482 511 483 512 
<< m1 >>
rect 483 511 484 512 
<< m1 >>
rect 484 511 485 512 
<< m1 >>
rect 485 511 486 512 
<< m1 >>
rect 486 511 487 512 
<< m1 >>
rect 487 511 488 512 
<< m1 >>
rect 19 512 20 513 
<< m1 >>
rect 34 512 35 513 
<< m1 >>
rect 70 512 71 513 
<< m1 >>
rect 100 512 101 513 
<< m1 >>
rect 124 512 125 513 
<< m2 >>
rect 186 512 187 513 
<< m1 >>
rect 226 512 227 513 
<< m1 >>
rect 262 512 263 513 
<< m1 >>
rect 268 512 269 513 
<< m2 >>
rect 320 512 321 513 
<< m2 >>
rect 361 512 362 513 
<< m2 >>
rect 372 512 373 513 
<< m2 >>
rect 379 512 380 513 
<< m2 >>
rect 446 512 447 513 
<< m2 >>
rect 451 512 452 513 
<< m2 >>
rect 472 512 473 513 
<< m1 >>
rect 19 513 20 514 
<< m1 >>
rect 34 513 35 514 
<< m1 >>
rect 70 513 71 514 
<< m1 >>
rect 100 513 101 514 
<< m1 >>
rect 124 513 125 514 
<< m1 >>
rect 186 513 187 514 
<< m2 >>
rect 186 513 187 514 
<< m2c >>
rect 186 513 187 514 
<< m1 >>
rect 186 513 187 514 
<< m2 >>
rect 186 513 187 514 
<< m1 >>
rect 226 513 227 514 
<< m1 >>
rect 262 513 263 514 
<< m1 >>
rect 268 513 269 514 
<< m1 >>
rect 320 513 321 514 
<< m2 >>
rect 320 513 321 514 
<< m2c >>
rect 320 513 321 514 
<< m1 >>
rect 320 513 321 514 
<< m2 >>
rect 320 513 321 514 
<< m1 >>
rect 321 513 322 514 
<< m1 >>
rect 322 513 323 514 
<< m1 >>
rect 323 513 324 514 
<< m1 >>
rect 324 513 325 514 
<< m1 >>
rect 325 513 326 514 
<< m1 >>
rect 361 513 362 514 
<< m2 >>
rect 361 513 362 514 
<< m2c >>
rect 361 513 362 514 
<< m1 >>
rect 361 513 362 514 
<< m2 >>
rect 361 513 362 514 
<< m1 >>
rect 370 513 371 514 
<< m1 >>
rect 371 513 372 514 
<< m1 >>
rect 372 513 373 514 
<< m2 >>
rect 372 513 373 514 
<< m2c >>
rect 372 513 373 514 
<< m1 >>
rect 372 513 373 514 
<< m2 >>
rect 372 513 373 514 
<< m1 >>
rect 379 513 380 514 
<< m2 >>
rect 379 513 380 514 
<< m2c >>
rect 379 513 380 514 
<< m1 >>
rect 379 513 380 514 
<< m2 >>
rect 379 513 380 514 
<< m1 >>
rect 446 513 447 514 
<< m2 >>
rect 446 513 447 514 
<< m2c >>
rect 446 513 447 514 
<< m1 >>
rect 446 513 447 514 
<< m2 >>
rect 446 513 447 514 
<< m1 >>
rect 447 513 448 514 
<< m1 >>
rect 448 513 449 514 
<< m1 >>
rect 451 513 452 514 
<< m2 >>
rect 451 513 452 514 
<< m2c >>
rect 451 513 452 514 
<< m1 >>
rect 451 513 452 514 
<< m2 >>
rect 451 513 452 514 
<< m1 >>
rect 472 513 473 514 
<< m2 >>
rect 472 513 473 514 
<< m2c >>
rect 472 513 473 514 
<< m1 >>
rect 472 513 473 514 
<< m2 >>
rect 472 513 473 514 
<< m1 >>
rect 19 514 20 515 
<< m1 >>
rect 34 514 35 515 
<< m1 >>
rect 70 514 71 515 
<< m1 >>
rect 100 514 101 515 
<< m1 >>
rect 124 514 125 515 
<< m1 >>
rect 186 514 187 515 
<< m1 >>
rect 226 514 227 515 
<< m1 >>
rect 262 514 263 515 
<< m1 >>
rect 268 514 269 515 
<< m1 >>
rect 325 514 326 515 
<< m1 >>
rect 361 514 362 515 
<< m1 >>
rect 370 514 371 515 
<< m1 >>
rect 379 514 380 515 
<< m1 >>
rect 394 514 395 515 
<< m1 >>
rect 395 514 396 515 
<< m1 >>
rect 396 514 397 515 
<< m1 >>
rect 397 514 398 515 
<< m1 >>
rect 448 514 449 515 
<< m1 >>
rect 451 514 452 515 
<< m1 >>
rect 472 514 473 515 
<< m1 >>
rect 19 515 20 516 
<< m1 >>
rect 34 515 35 516 
<< m1 >>
rect 70 515 71 516 
<< m1 >>
rect 100 515 101 516 
<< m1 >>
rect 124 515 125 516 
<< m1 >>
rect 186 515 187 516 
<< m1 >>
rect 226 515 227 516 
<< m1 >>
rect 262 515 263 516 
<< m1 >>
rect 268 515 269 516 
<< m1 >>
rect 325 515 326 516 
<< m1 >>
rect 361 515 362 516 
<< m1 >>
rect 370 515 371 516 
<< m1 >>
rect 379 515 380 516 
<< m1 >>
rect 394 515 395 516 
<< m1 >>
rect 397 515 398 516 
<< m1 >>
rect 448 515 449 516 
<< m1 >>
rect 451 515 452 516 
<< m1 >>
rect 472 515 473 516 
<< pdiffusion >>
rect 12 516 13 517 
<< pdiffusion >>
rect 13 516 14 517 
<< pdiffusion >>
rect 14 516 15 517 
<< pdiffusion >>
rect 15 516 16 517 
<< pdiffusion >>
rect 16 516 17 517 
<< pdiffusion >>
rect 17 516 18 517 
<< m1 >>
rect 19 516 20 517 
<< pdiffusion >>
rect 30 516 31 517 
<< pdiffusion >>
rect 31 516 32 517 
<< pdiffusion >>
rect 32 516 33 517 
<< pdiffusion >>
rect 33 516 34 517 
<< m1 >>
rect 34 516 35 517 
<< pdiffusion >>
rect 34 516 35 517 
<< pdiffusion >>
rect 35 516 36 517 
<< pdiffusion >>
rect 48 516 49 517 
<< pdiffusion >>
rect 49 516 50 517 
<< pdiffusion >>
rect 50 516 51 517 
<< pdiffusion >>
rect 51 516 52 517 
<< pdiffusion >>
rect 52 516 53 517 
<< pdiffusion >>
rect 53 516 54 517 
<< pdiffusion >>
rect 66 516 67 517 
<< pdiffusion >>
rect 67 516 68 517 
<< pdiffusion >>
rect 68 516 69 517 
<< pdiffusion >>
rect 69 516 70 517 
<< m1 >>
rect 70 516 71 517 
<< pdiffusion >>
rect 70 516 71 517 
<< pdiffusion >>
rect 71 516 72 517 
<< pdiffusion >>
rect 84 516 85 517 
<< pdiffusion >>
rect 85 516 86 517 
<< pdiffusion >>
rect 86 516 87 517 
<< pdiffusion >>
rect 87 516 88 517 
<< pdiffusion >>
rect 88 516 89 517 
<< pdiffusion >>
rect 89 516 90 517 
<< m1 >>
rect 100 516 101 517 
<< pdiffusion >>
rect 102 516 103 517 
<< pdiffusion >>
rect 103 516 104 517 
<< pdiffusion >>
rect 104 516 105 517 
<< pdiffusion >>
rect 105 516 106 517 
<< pdiffusion >>
rect 106 516 107 517 
<< pdiffusion >>
rect 107 516 108 517 
<< pdiffusion >>
rect 120 516 121 517 
<< pdiffusion >>
rect 121 516 122 517 
<< pdiffusion >>
rect 122 516 123 517 
<< pdiffusion >>
rect 123 516 124 517 
<< m1 >>
rect 124 516 125 517 
<< pdiffusion >>
rect 124 516 125 517 
<< pdiffusion >>
rect 125 516 126 517 
<< pdiffusion >>
rect 138 516 139 517 
<< pdiffusion >>
rect 139 516 140 517 
<< pdiffusion >>
rect 140 516 141 517 
<< pdiffusion >>
rect 141 516 142 517 
<< pdiffusion >>
rect 142 516 143 517 
<< pdiffusion >>
rect 143 516 144 517 
<< pdiffusion >>
rect 156 516 157 517 
<< pdiffusion >>
rect 157 516 158 517 
<< pdiffusion >>
rect 158 516 159 517 
<< pdiffusion >>
rect 159 516 160 517 
<< pdiffusion >>
rect 160 516 161 517 
<< pdiffusion >>
rect 161 516 162 517 
<< pdiffusion >>
rect 174 516 175 517 
<< pdiffusion >>
rect 175 516 176 517 
<< pdiffusion >>
rect 176 516 177 517 
<< pdiffusion >>
rect 177 516 178 517 
<< pdiffusion >>
rect 178 516 179 517 
<< pdiffusion >>
rect 179 516 180 517 
<< m1 >>
rect 186 516 187 517 
<< pdiffusion >>
rect 192 516 193 517 
<< pdiffusion >>
rect 193 516 194 517 
<< pdiffusion >>
rect 194 516 195 517 
<< pdiffusion >>
rect 195 516 196 517 
<< pdiffusion >>
rect 196 516 197 517 
<< pdiffusion >>
rect 197 516 198 517 
<< m1 >>
rect 226 516 227 517 
<< pdiffusion >>
rect 228 516 229 517 
<< pdiffusion >>
rect 229 516 230 517 
<< pdiffusion >>
rect 230 516 231 517 
<< pdiffusion >>
rect 231 516 232 517 
<< pdiffusion >>
rect 232 516 233 517 
<< pdiffusion >>
rect 233 516 234 517 
<< pdiffusion >>
rect 246 516 247 517 
<< pdiffusion >>
rect 247 516 248 517 
<< pdiffusion >>
rect 248 516 249 517 
<< pdiffusion >>
rect 249 516 250 517 
<< pdiffusion >>
rect 250 516 251 517 
<< pdiffusion >>
rect 251 516 252 517 
<< m1 >>
rect 262 516 263 517 
<< pdiffusion >>
rect 264 516 265 517 
<< pdiffusion >>
rect 265 516 266 517 
<< pdiffusion >>
rect 266 516 267 517 
<< pdiffusion >>
rect 267 516 268 517 
<< m1 >>
rect 268 516 269 517 
<< pdiffusion >>
rect 268 516 269 517 
<< pdiffusion >>
rect 269 516 270 517 
<< pdiffusion >>
rect 282 516 283 517 
<< pdiffusion >>
rect 283 516 284 517 
<< pdiffusion >>
rect 284 516 285 517 
<< pdiffusion >>
rect 285 516 286 517 
<< pdiffusion >>
rect 286 516 287 517 
<< pdiffusion >>
rect 287 516 288 517 
<< pdiffusion >>
rect 300 516 301 517 
<< pdiffusion >>
rect 301 516 302 517 
<< pdiffusion >>
rect 302 516 303 517 
<< pdiffusion >>
rect 303 516 304 517 
<< pdiffusion >>
rect 304 516 305 517 
<< pdiffusion >>
rect 305 516 306 517 
<< pdiffusion >>
rect 318 516 319 517 
<< pdiffusion >>
rect 319 516 320 517 
<< pdiffusion >>
rect 320 516 321 517 
<< pdiffusion >>
rect 321 516 322 517 
<< pdiffusion >>
rect 322 516 323 517 
<< pdiffusion >>
rect 323 516 324 517 
<< m1 >>
rect 325 516 326 517 
<< pdiffusion >>
rect 336 516 337 517 
<< pdiffusion >>
rect 337 516 338 517 
<< pdiffusion >>
rect 338 516 339 517 
<< pdiffusion >>
rect 339 516 340 517 
<< pdiffusion >>
rect 340 516 341 517 
<< pdiffusion >>
rect 341 516 342 517 
<< pdiffusion >>
rect 354 516 355 517 
<< pdiffusion >>
rect 355 516 356 517 
<< pdiffusion >>
rect 356 516 357 517 
<< pdiffusion >>
rect 357 516 358 517 
<< pdiffusion >>
rect 358 516 359 517 
<< pdiffusion >>
rect 359 516 360 517 
<< m1 >>
rect 361 516 362 517 
<< m1 >>
rect 370 516 371 517 
<< pdiffusion >>
rect 372 516 373 517 
<< pdiffusion >>
rect 373 516 374 517 
<< pdiffusion >>
rect 374 516 375 517 
<< pdiffusion >>
rect 375 516 376 517 
<< pdiffusion >>
rect 376 516 377 517 
<< pdiffusion >>
rect 377 516 378 517 
<< m1 >>
rect 379 516 380 517 
<< pdiffusion >>
rect 390 516 391 517 
<< pdiffusion >>
rect 391 516 392 517 
<< pdiffusion >>
rect 392 516 393 517 
<< pdiffusion >>
rect 393 516 394 517 
<< m1 >>
rect 394 516 395 517 
<< pdiffusion >>
rect 394 516 395 517 
<< pdiffusion >>
rect 395 516 396 517 
<< m1 >>
rect 397 516 398 517 
<< pdiffusion >>
rect 408 516 409 517 
<< pdiffusion >>
rect 409 516 410 517 
<< pdiffusion >>
rect 410 516 411 517 
<< pdiffusion >>
rect 411 516 412 517 
<< pdiffusion >>
rect 412 516 413 517 
<< pdiffusion >>
rect 413 516 414 517 
<< pdiffusion >>
rect 426 516 427 517 
<< pdiffusion >>
rect 427 516 428 517 
<< pdiffusion >>
rect 428 516 429 517 
<< pdiffusion >>
rect 429 516 430 517 
<< pdiffusion >>
rect 430 516 431 517 
<< pdiffusion >>
rect 431 516 432 517 
<< pdiffusion >>
rect 444 516 445 517 
<< pdiffusion >>
rect 445 516 446 517 
<< pdiffusion >>
rect 446 516 447 517 
<< pdiffusion >>
rect 447 516 448 517 
<< m1 >>
rect 448 516 449 517 
<< pdiffusion >>
rect 448 516 449 517 
<< pdiffusion >>
rect 449 516 450 517 
<< m1 >>
rect 451 516 452 517 
<< pdiffusion >>
rect 462 516 463 517 
<< pdiffusion >>
rect 463 516 464 517 
<< pdiffusion >>
rect 464 516 465 517 
<< pdiffusion >>
rect 465 516 466 517 
<< pdiffusion >>
rect 466 516 467 517 
<< pdiffusion >>
rect 467 516 468 517 
<< m1 >>
rect 472 516 473 517 
<< pdiffusion >>
rect 480 516 481 517 
<< pdiffusion >>
rect 481 516 482 517 
<< pdiffusion >>
rect 482 516 483 517 
<< pdiffusion >>
rect 483 516 484 517 
<< pdiffusion >>
rect 484 516 485 517 
<< pdiffusion >>
rect 485 516 486 517 
<< pdiffusion >>
rect 498 516 499 517 
<< pdiffusion >>
rect 499 516 500 517 
<< pdiffusion >>
rect 500 516 501 517 
<< pdiffusion >>
rect 501 516 502 517 
<< pdiffusion >>
rect 502 516 503 517 
<< pdiffusion >>
rect 503 516 504 517 
<< pdiffusion >>
rect 516 516 517 517 
<< pdiffusion >>
rect 517 516 518 517 
<< pdiffusion >>
rect 518 516 519 517 
<< pdiffusion >>
rect 519 516 520 517 
<< pdiffusion >>
rect 520 516 521 517 
<< pdiffusion >>
rect 521 516 522 517 
<< pdiffusion >>
rect 12 517 13 518 
<< pdiffusion >>
rect 13 517 14 518 
<< pdiffusion >>
rect 14 517 15 518 
<< pdiffusion >>
rect 15 517 16 518 
<< pdiffusion >>
rect 16 517 17 518 
<< pdiffusion >>
rect 17 517 18 518 
<< m1 >>
rect 19 517 20 518 
<< pdiffusion >>
rect 30 517 31 518 
<< pdiffusion >>
rect 31 517 32 518 
<< pdiffusion >>
rect 32 517 33 518 
<< pdiffusion >>
rect 33 517 34 518 
<< pdiffusion >>
rect 34 517 35 518 
<< pdiffusion >>
rect 35 517 36 518 
<< pdiffusion >>
rect 48 517 49 518 
<< pdiffusion >>
rect 49 517 50 518 
<< pdiffusion >>
rect 50 517 51 518 
<< pdiffusion >>
rect 51 517 52 518 
<< pdiffusion >>
rect 52 517 53 518 
<< pdiffusion >>
rect 53 517 54 518 
<< pdiffusion >>
rect 66 517 67 518 
<< pdiffusion >>
rect 67 517 68 518 
<< pdiffusion >>
rect 68 517 69 518 
<< pdiffusion >>
rect 69 517 70 518 
<< pdiffusion >>
rect 70 517 71 518 
<< pdiffusion >>
rect 71 517 72 518 
<< pdiffusion >>
rect 84 517 85 518 
<< pdiffusion >>
rect 85 517 86 518 
<< pdiffusion >>
rect 86 517 87 518 
<< pdiffusion >>
rect 87 517 88 518 
<< pdiffusion >>
rect 88 517 89 518 
<< pdiffusion >>
rect 89 517 90 518 
<< m1 >>
rect 100 517 101 518 
<< pdiffusion >>
rect 102 517 103 518 
<< pdiffusion >>
rect 103 517 104 518 
<< pdiffusion >>
rect 104 517 105 518 
<< pdiffusion >>
rect 105 517 106 518 
<< pdiffusion >>
rect 106 517 107 518 
<< pdiffusion >>
rect 107 517 108 518 
<< pdiffusion >>
rect 120 517 121 518 
<< pdiffusion >>
rect 121 517 122 518 
<< pdiffusion >>
rect 122 517 123 518 
<< pdiffusion >>
rect 123 517 124 518 
<< pdiffusion >>
rect 124 517 125 518 
<< pdiffusion >>
rect 125 517 126 518 
<< pdiffusion >>
rect 138 517 139 518 
<< pdiffusion >>
rect 139 517 140 518 
<< pdiffusion >>
rect 140 517 141 518 
<< pdiffusion >>
rect 141 517 142 518 
<< pdiffusion >>
rect 142 517 143 518 
<< pdiffusion >>
rect 143 517 144 518 
<< pdiffusion >>
rect 156 517 157 518 
<< pdiffusion >>
rect 157 517 158 518 
<< pdiffusion >>
rect 158 517 159 518 
<< pdiffusion >>
rect 159 517 160 518 
<< pdiffusion >>
rect 160 517 161 518 
<< pdiffusion >>
rect 161 517 162 518 
<< pdiffusion >>
rect 174 517 175 518 
<< pdiffusion >>
rect 175 517 176 518 
<< pdiffusion >>
rect 176 517 177 518 
<< pdiffusion >>
rect 177 517 178 518 
<< pdiffusion >>
rect 178 517 179 518 
<< pdiffusion >>
rect 179 517 180 518 
<< m1 >>
rect 186 517 187 518 
<< pdiffusion >>
rect 192 517 193 518 
<< pdiffusion >>
rect 193 517 194 518 
<< pdiffusion >>
rect 194 517 195 518 
<< pdiffusion >>
rect 195 517 196 518 
<< pdiffusion >>
rect 196 517 197 518 
<< pdiffusion >>
rect 197 517 198 518 
<< m1 >>
rect 226 517 227 518 
<< pdiffusion >>
rect 228 517 229 518 
<< pdiffusion >>
rect 229 517 230 518 
<< pdiffusion >>
rect 230 517 231 518 
<< pdiffusion >>
rect 231 517 232 518 
<< pdiffusion >>
rect 232 517 233 518 
<< pdiffusion >>
rect 233 517 234 518 
<< pdiffusion >>
rect 246 517 247 518 
<< pdiffusion >>
rect 247 517 248 518 
<< pdiffusion >>
rect 248 517 249 518 
<< pdiffusion >>
rect 249 517 250 518 
<< pdiffusion >>
rect 250 517 251 518 
<< pdiffusion >>
rect 251 517 252 518 
<< m1 >>
rect 262 517 263 518 
<< pdiffusion >>
rect 264 517 265 518 
<< pdiffusion >>
rect 265 517 266 518 
<< pdiffusion >>
rect 266 517 267 518 
<< pdiffusion >>
rect 267 517 268 518 
<< pdiffusion >>
rect 268 517 269 518 
<< pdiffusion >>
rect 269 517 270 518 
<< pdiffusion >>
rect 282 517 283 518 
<< pdiffusion >>
rect 283 517 284 518 
<< pdiffusion >>
rect 284 517 285 518 
<< pdiffusion >>
rect 285 517 286 518 
<< pdiffusion >>
rect 286 517 287 518 
<< pdiffusion >>
rect 287 517 288 518 
<< pdiffusion >>
rect 300 517 301 518 
<< pdiffusion >>
rect 301 517 302 518 
<< pdiffusion >>
rect 302 517 303 518 
<< pdiffusion >>
rect 303 517 304 518 
<< pdiffusion >>
rect 304 517 305 518 
<< pdiffusion >>
rect 305 517 306 518 
<< pdiffusion >>
rect 318 517 319 518 
<< pdiffusion >>
rect 319 517 320 518 
<< pdiffusion >>
rect 320 517 321 518 
<< pdiffusion >>
rect 321 517 322 518 
<< pdiffusion >>
rect 322 517 323 518 
<< pdiffusion >>
rect 323 517 324 518 
<< m1 >>
rect 325 517 326 518 
<< pdiffusion >>
rect 336 517 337 518 
<< pdiffusion >>
rect 337 517 338 518 
<< pdiffusion >>
rect 338 517 339 518 
<< pdiffusion >>
rect 339 517 340 518 
<< pdiffusion >>
rect 340 517 341 518 
<< pdiffusion >>
rect 341 517 342 518 
<< pdiffusion >>
rect 354 517 355 518 
<< pdiffusion >>
rect 355 517 356 518 
<< pdiffusion >>
rect 356 517 357 518 
<< pdiffusion >>
rect 357 517 358 518 
<< pdiffusion >>
rect 358 517 359 518 
<< pdiffusion >>
rect 359 517 360 518 
<< m1 >>
rect 361 517 362 518 
<< m1 >>
rect 370 517 371 518 
<< pdiffusion >>
rect 372 517 373 518 
<< pdiffusion >>
rect 373 517 374 518 
<< pdiffusion >>
rect 374 517 375 518 
<< pdiffusion >>
rect 375 517 376 518 
<< pdiffusion >>
rect 376 517 377 518 
<< pdiffusion >>
rect 377 517 378 518 
<< m1 >>
rect 379 517 380 518 
<< pdiffusion >>
rect 390 517 391 518 
<< pdiffusion >>
rect 391 517 392 518 
<< pdiffusion >>
rect 392 517 393 518 
<< pdiffusion >>
rect 393 517 394 518 
<< pdiffusion >>
rect 394 517 395 518 
<< pdiffusion >>
rect 395 517 396 518 
<< m1 >>
rect 397 517 398 518 
<< pdiffusion >>
rect 408 517 409 518 
<< pdiffusion >>
rect 409 517 410 518 
<< pdiffusion >>
rect 410 517 411 518 
<< pdiffusion >>
rect 411 517 412 518 
<< pdiffusion >>
rect 412 517 413 518 
<< pdiffusion >>
rect 413 517 414 518 
<< pdiffusion >>
rect 426 517 427 518 
<< pdiffusion >>
rect 427 517 428 518 
<< pdiffusion >>
rect 428 517 429 518 
<< pdiffusion >>
rect 429 517 430 518 
<< pdiffusion >>
rect 430 517 431 518 
<< pdiffusion >>
rect 431 517 432 518 
<< pdiffusion >>
rect 444 517 445 518 
<< pdiffusion >>
rect 445 517 446 518 
<< pdiffusion >>
rect 446 517 447 518 
<< pdiffusion >>
rect 447 517 448 518 
<< pdiffusion >>
rect 448 517 449 518 
<< pdiffusion >>
rect 449 517 450 518 
<< m1 >>
rect 451 517 452 518 
<< pdiffusion >>
rect 462 517 463 518 
<< pdiffusion >>
rect 463 517 464 518 
<< pdiffusion >>
rect 464 517 465 518 
<< pdiffusion >>
rect 465 517 466 518 
<< pdiffusion >>
rect 466 517 467 518 
<< pdiffusion >>
rect 467 517 468 518 
<< m1 >>
rect 472 517 473 518 
<< pdiffusion >>
rect 480 517 481 518 
<< pdiffusion >>
rect 481 517 482 518 
<< pdiffusion >>
rect 482 517 483 518 
<< pdiffusion >>
rect 483 517 484 518 
<< pdiffusion >>
rect 484 517 485 518 
<< pdiffusion >>
rect 485 517 486 518 
<< pdiffusion >>
rect 498 517 499 518 
<< pdiffusion >>
rect 499 517 500 518 
<< pdiffusion >>
rect 500 517 501 518 
<< pdiffusion >>
rect 501 517 502 518 
<< pdiffusion >>
rect 502 517 503 518 
<< pdiffusion >>
rect 503 517 504 518 
<< pdiffusion >>
rect 516 517 517 518 
<< pdiffusion >>
rect 517 517 518 518 
<< pdiffusion >>
rect 518 517 519 518 
<< pdiffusion >>
rect 519 517 520 518 
<< pdiffusion >>
rect 520 517 521 518 
<< pdiffusion >>
rect 521 517 522 518 
<< pdiffusion >>
rect 12 518 13 519 
<< pdiffusion >>
rect 13 518 14 519 
<< pdiffusion >>
rect 14 518 15 519 
<< pdiffusion >>
rect 15 518 16 519 
<< pdiffusion >>
rect 16 518 17 519 
<< pdiffusion >>
rect 17 518 18 519 
<< m1 >>
rect 19 518 20 519 
<< pdiffusion >>
rect 30 518 31 519 
<< pdiffusion >>
rect 31 518 32 519 
<< pdiffusion >>
rect 32 518 33 519 
<< pdiffusion >>
rect 33 518 34 519 
<< pdiffusion >>
rect 34 518 35 519 
<< pdiffusion >>
rect 35 518 36 519 
<< pdiffusion >>
rect 48 518 49 519 
<< pdiffusion >>
rect 49 518 50 519 
<< pdiffusion >>
rect 50 518 51 519 
<< pdiffusion >>
rect 51 518 52 519 
<< pdiffusion >>
rect 52 518 53 519 
<< pdiffusion >>
rect 53 518 54 519 
<< pdiffusion >>
rect 66 518 67 519 
<< pdiffusion >>
rect 67 518 68 519 
<< pdiffusion >>
rect 68 518 69 519 
<< pdiffusion >>
rect 69 518 70 519 
<< pdiffusion >>
rect 70 518 71 519 
<< pdiffusion >>
rect 71 518 72 519 
<< pdiffusion >>
rect 84 518 85 519 
<< pdiffusion >>
rect 85 518 86 519 
<< pdiffusion >>
rect 86 518 87 519 
<< pdiffusion >>
rect 87 518 88 519 
<< pdiffusion >>
rect 88 518 89 519 
<< pdiffusion >>
rect 89 518 90 519 
<< m1 >>
rect 100 518 101 519 
<< pdiffusion >>
rect 102 518 103 519 
<< pdiffusion >>
rect 103 518 104 519 
<< pdiffusion >>
rect 104 518 105 519 
<< pdiffusion >>
rect 105 518 106 519 
<< pdiffusion >>
rect 106 518 107 519 
<< pdiffusion >>
rect 107 518 108 519 
<< pdiffusion >>
rect 120 518 121 519 
<< pdiffusion >>
rect 121 518 122 519 
<< pdiffusion >>
rect 122 518 123 519 
<< pdiffusion >>
rect 123 518 124 519 
<< pdiffusion >>
rect 124 518 125 519 
<< pdiffusion >>
rect 125 518 126 519 
<< pdiffusion >>
rect 138 518 139 519 
<< pdiffusion >>
rect 139 518 140 519 
<< pdiffusion >>
rect 140 518 141 519 
<< pdiffusion >>
rect 141 518 142 519 
<< pdiffusion >>
rect 142 518 143 519 
<< pdiffusion >>
rect 143 518 144 519 
<< pdiffusion >>
rect 156 518 157 519 
<< pdiffusion >>
rect 157 518 158 519 
<< pdiffusion >>
rect 158 518 159 519 
<< pdiffusion >>
rect 159 518 160 519 
<< pdiffusion >>
rect 160 518 161 519 
<< pdiffusion >>
rect 161 518 162 519 
<< pdiffusion >>
rect 174 518 175 519 
<< pdiffusion >>
rect 175 518 176 519 
<< pdiffusion >>
rect 176 518 177 519 
<< pdiffusion >>
rect 177 518 178 519 
<< pdiffusion >>
rect 178 518 179 519 
<< pdiffusion >>
rect 179 518 180 519 
<< m1 >>
rect 186 518 187 519 
<< pdiffusion >>
rect 192 518 193 519 
<< pdiffusion >>
rect 193 518 194 519 
<< pdiffusion >>
rect 194 518 195 519 
<< pdiffusion >>
rect 195 518 196 519 
<< pdiffusion >>
rect 196 518 197 519 
<< pdiffusion >>
rect 197 518 198 519 
<< m1 >>
rect 226 518 227 519 
<< pdiffusion >>
rect 228 518 229 519 
<< pdiffusion >>
rect 229 518 230 519 
<< pdiffusion >>
rect 230 518 231 519 
<< pdiffusion >>
rect 231 518 232 519 
<< pdiffusion >>
rect 232 518 233 519 
<< pdiffusion >>
rect 233 518 234 519 
<< pdiffusion >>
rect 246 518 247 519 
<< pdiffusion >>
rect 247 518 248 519 
<< pdiffusion >>
rect 248 518 249 519 
<< pdiffusion >>
rect 249 518 250 519 
<< pdiffusion >>
rect 250 518 251 519 
<< pdiffusion >>
rect 251 518 252 519 
<< m1 >>
rect 262 518 263 519 
<< pdiffusion >>
rect 264 518 265 519 
<< pdiffusion >>
rect 265 518 266 519 
<< pdiffusion >>
rect 266 518 267 519 
<< pdiffusion >>
rect 267 518 268 519 
<< pdiffusion >>
rect 268 518 269 519 
<< pdiffusion >>
rect 269 518 270 519 
<< pdiffusion >>
rect 282 518 283 519 
<< pdiffusion >>
rect 283 518 284 519 
<< pdiffusion >>
rect 284 518 285 519 
<< pdiffusion >>
rect 285 518 286 519 
<< pdiffusion >>
rect 286 518 287 519 
<< pdiffusion >>
rect 287 518 288 519 
<< pdiffusion >>
rect 300 518 301 519 
<< pdiffusion >>
rect 301 518 302 519 
<< pdiffusion >>
rect 302 518 303 519 
<< pdiffusion >>
rect 303 518 304 519 
<< pdiffusion >>
rect 304 518 305 519 
<< pdiffusion >>
rect 305 518 306 519 
<< pdiffusion >>
rect 318 518 319 519 
<< pdiffusion >>
rect 319 518 320 519 
<< pdiffusion >>
rect 320 518 321 519 
<< pdiffusion >>
rect 321 518 322 519 
<< pdiffusion >>
rect 322 518 323 519 
<< pdiffusion >>
rect 323 518 324 519 
<< m1 >>
rect 325 518 326 519 
<< pdiffusion >>
rect 336 518 337 519 
<< pdiffusion >>
rect 337 518 338 519 
<< pdiffusion >>
rect 338 518 339 519 
<< pdiffusion >>
rect 339 518 340 519 
<< pdiffusion >>
rect 340 518 341 519 
<< pdiffusion >>
rect 341 518 342 519 
<< pdiffusion >>
rect 354 518 355 519 
<< pdiffusion >>
rect 355 518 356 519 
<< pdiffusion >>
rect 356 518 357 519 
<< pdiffusion >>
rect 357 518 358 519 
<< pdiffusion >>
rect 358 518 359 519 
<< pdiffusion >>
rect 359 518 360 519 
<< m1 >>
rect 361 518 362 519 
<< m1 >>
rect 370 518 371 519 
<< pdiffusion >>
rect 372 518 373 519 
<< pdiffusion >>
rect 373 518 374 519 
<< pdiffusion >>
rect 374 518 375 519 
<< pdiffusion >>
rect 375 518 376 519 
<< pdiffusion >>
rect 376 518 377 519 
<< pdiffusion >>
rect 377 518 378 519 
<< m1 >>
rect 379 518 380 519 
<< pdiffusion >>
rect 390 518 391 519 
<< pdiffusion >>
rect 391 518 392 519 
<< pdiffusion >>
rect 392 518 393 519 
<< pdiffusion >>
rect 393 518 394 519 
<< pdiffusion >>
rect 394 518 395 519 
<< pdiffusion >>
rect 395 518 396 519 
<< m1 >>
rect 397 518 398 519 
<< pdiffusion >>
rect 408 518 409 519 
<< pdiffusion >>
rect 409 518 410 519 
<< pdiffusion >>
rect 410 518 411 519 
<< pdiffusion >>
rect 411 518 412 519 
<< pdiffusion >>
rect 412 518 413 519 
<< pdiffusion >>
rect 413 518 414 519 
<< pdiffusion >>
rect 426 518 427 519 
<< pdiffusion >>
rect 427 518 428 519 
<< pdiffusion >>
rect 428 518 429 519 
<< pdiffusion >>
rect 429 518 430 519 
<< pdiffusion >>
rect 430 518 431 519 
<< pdiffusion >>
rect 431 518 432 519 
<< pdiffusion >>
rect 444 518 445 519 
<< pdiffusion >>
rect 445 518 446 519 
<< pdiffusion >>
rect 446 518 447 519 
<< pdiffusion >>
rect 447 518 448 519 
<< pdiffusion >>
rect 448 518 449 519 
<< pdiffusion >>
rect 449 518 450 519 
<< m1 >>
rect 451 518 452 519 
<< pdiffusion >>
rect 462 518 463 519 
<< pdiffusion >>
rect 463 518 464 519 
<< pdiffusion >>
rect 464 518 465 519 
<< pdiffusion >>
rect 465 518 466 519 
<< pdiffusion >>
rect 466 518 467 519 
<< pdiffusion >>
rect 467 518 468 519 
<< m1 >>
rect 472 518 473 519 
<< pdiffusion >>
rect 480 518 481 519 
<< pdiffusion >>
rect 481 518 482 519 
<< pdiffusion >>
rect 482 518 483 519 
<< pdiffusion >>
rect 483 518 484 519 
<< pdiffusion >>
rect 484 518 485 519 
<< pdiffusion >>
rect 485 518 486 519 
<< pdiffusion >>
rect 498 518 499 519 
<< pdiffusion >>
rect 499 518 500 519 
<< pdiffusion >>
rect 500 518 501 519 
<< pdiffusion >>
rect 501 518 502 519 
<< pdiffusion >>
rect 502 518 503 519 
<< pdiffusion >>
rect 503 518 504 519 
<< pdiffusion >>
rect 516 518 517 519 
<< pdiffusion >>
rect 517 518 518 519 
<< pdiffusion >>
rect 518 518 519 519 
<< pdiffusion >>
rect 519 518 520 519 
<< pdiffusion >>
rect 520 518 521 519 
<< pdiffusion >>
rect 521 518 522 519 
<< pdiffusion >>
rect 12 519 13 520 
<< pdiffusion >>
rect 13 519 14 520 
<< pdiffusion >>
rect 14 519 15 520 
<< pdiffusion >>
rect 15 519 16 520 
<< pdiffusion >>
rect 16 519 17 520 
<< pdiffusion >>
rect 17 519 18 520 
<< m1 >>
rect 19 519 20 520 
<< pdiffusion >>
rect 30 519 31 520 
<< pdiffusion >>
rect 31 519 32 520 
<< pdiffusion >>
rect 32 519 33 520 
<< pdiffusion >>
rect 33 519 34 520 
<< pdiffusion >>
rect 34 519 35 520 
<< pdiffusion >>
rect 35 519 36 520 
<< pdiffusion >>
rect 48 519 49 520 
<< pdiffusion >>
rect 49 519 50 520 
<< pdiffusion >>
rect 50 519 51 520 
<< pdiffusion >>
rect 51 519 52 520 
<< pdiffusion >>
rect 52 519 53 520 
<< pdiffusion >>
rect 53 519 54 520 
<< pdiffusion >>
rect 66 519 67 520 
<< pdiffusion >>
rect 67 519 68 520 
<< pdiffusion >>
rect 68 519 69 520 
<< pdiffusion >>
rect 69 519 70 520 
<< pdiffusion >>
rect 70 519 71 520 
<< pdiffusion >>
rect 71 519 72 520 
<< pdiffusion >>
rect 84 519 85 520 
<< pdiffusion >>
rect 85 519 86 520 
<< pdiffusion >>
rect 86 519 87 520 
<< pdiffusion >>
rect 87 519 88 520 
<< pdiffusion >>
rect 88 519 89 520 
<< pdiffusion >>
rect 89 519 90 520 
<< m1 >>
rect 100 519 101 520 
<< pdiffusion >>
rect 102 519 103 520 
<< pdiffusion >>
rect 103 519 104 520 
<< pdiffusion >>
rect 104 519 105 520 
<< pdiffusion >>
rect 105 519 106 520 
<< pdiffusion >>
rect 106 519 107 520 
<< pdiffusion >>
rect 107 519 108 520 
<< pdiffusion >>
rect 120 519 121 520 
<< pdiffusion >>
rect 121 519 122 520 
<< pdiffusion >>
rect 122 519 123 520 
<< pdiffusion >>
rect 123 519 124 520 
<< pdiffusion >>
rect 124 519 125 520 
<< pdiffusion >>
rect 125 519 126 520 
<< pdiffusion >>
rect 138 519 139 520 
<< pdiffusion >>
rect 139 519 140 520 
<< pdiffusion >>
rect 140 519 141 520 
<< pdiffusion >>
rect 141 519 142 520 
<< pdiffusion >>
rect 142 519 143 520 
<< pdiffusion >>
rect 143 519 144 520 
<< pdiffusion >>
rect 156 519 157 520 
<< pdiffusion >>
rect 157 519 158 520 
<< pdiffusion >>
rect 158 519 159 520 
<< pdiffusion >>
rect 159 519 160 520 
<< pdiffusion >>
rect 160 519 161 520 
<< pdiffusion >>
rect 161 519 162 520 
<< pdiffusion >>
rect 174 519 175 520 
<< pdiffusion >>
rect 175 519 176 520 
<< pdiffusion >>
rect 176 519 177 520 
<< pdiffusion >>
rect 177 519 178 520 
<< pdiffusion >>
rect 178 519 179 520 
<< pdiffusion >>
rect 179 519 180 520 
<< m1 >>
rect 186 519 187 520 
<< pdiffusion >>
rect 192 519 193 520 
<< pdiffusion >>
rect 193 519 194 520 
<< pdiffusion >>
rect 194 519 195 520 
<< pdiffusion >>
rect 195 519 196 520 
<< pdiffusion >>
rect 196 519 197 520 
<< pdiffusion >>
rect 197 519 198 520 
<< m1 >>
rect 226 519 227 520 
<< pdiffusion >>
rect 228 519 229 520 
<< pdiffusion >>
rect 229 519 230 520 
<< pdiffusion >>
rect 230 519 231 520 
<< pdiffusion >>
rect 231 519 232 520 
<< pdiffusion >>
rect 232 519 233 520 
<< pdiffusion >>
rect 233 519 234 520 
<< pdiffusion >>
rect 246 519 247 520 
<< pdiffusion >>
rect 247 519 248 520 
<< pdiffusion >>
rect 248 519 249 520 
<< pdiffusion >>
rect 249 519 250 520 
<< pdiffusion >>
rect 250 519 251 520 
<< pdiffusion >>
rect 251 519 252 520 
<< m1 >>
rect 262 519 263 520 
<< pdiffusion >>
rect 264 519 265 520 
<< pdiffusion >>
rect 265 519 266 520 
<< pdiffusion >>
rect 266 519 267 520 
<< pdiffusion >>
rect 267 519 268 520 
<< pdiffusion >>
rect 268 519 269 520 
<< pdiffusion >>
rect 269 519 270 520 
<< pdiffusion >>
rect 282 519 283 520 
<< pdiffusion >>
rect 283 519 284 520 
<< pdiffusion >>
rect 284 519 285 520 
<< pdiffusion >>
rect 285 519 286 520 
<< pdiffusion >>
rect 286 519 287 520 
<< pdiffusion >>
rect 287 519 288 520 
<< pdiffusion >>
rect 300 519 301 520 
<< pdiffusion >>
rect 301 519 302 520 
<< pdiffusion >>
rect 302 519 303 520 
<< pdiffusion >>
rect 303 519 304 520 
<< pdiffusion >>
rect 304 519 305 520 
<< pdiffusion >>
rect 305 519 306 520 
<< pdiffusion >>
rect 318 519 319 520 
<< pdiffusion >>
rect 319 519 320 520 
<< pdiffusion >>
rect 320 519 321 520 
<< pdiffusion >>
rect 321 519 322 520 
<< pdiffusion >>
rect 322 519 323 520 
<< pdiffusion >>
rect 323 519 324 520 
<< m1 >>
rect 325 519 326 520 
<< pdiffusion >>
rect 336 519 337 520 
<< pdiffusion >>
rect 337 519 338 520 
<< pdiffusion >>
rect 338 519 339 520 
<< pdiffusion >>
rect 339 519 340 520 
<< pdiffusion >>
rect 340 519 341 520 
<< pdiffusion >>
rect 341 519 342 520 
<< pdiffusion >>
rect 354 519 355 520 
<< pdiffusion >>
rect 355 519 356 520 
<< pdiffusion >>
rect 356 519 357 520 
<< pdiffusion >>
rect 357 519 358 520 
<< pdiffusion >>
rect 358 519 359 520 
<< pdiffusion >>
rect 359 519 360 520 
<< m1 >>
rect 361 519 362 520 
<< m1 >>
rect 370 519 371 520 
<< pdiffusion >>
rect 372 519 373 520 
<< pdiffusion >>
rect 373 519 374 520 
<< pdiffusion >>
rect 374 519 375 520 
<< pdiffusion >>
rect 375 519 376 520 
<< pdiffusion >>
rect 376 519 377 520 
<< pdiffusion >>
rect 377 519 378 520 
<< m1 >>
rect 379 519 380 520 
<< pdiffusion >>
rect 390 519 391 520 
<< pdiffusion >>
rect 391 519 392 520 
<< pdiffusion >>
rect 392 519 393 520 
<< pdiffusion >>
rect 393 519 394 520 
<< pdiffusion >>
rect 394 519 395 520 
<< pdiffusion >>
rect 395 519 396 520 
<< m1 >>
rect 397 519 398 520 
<< pdiffusion >>
rect 408 519 409 520 
<< pdiffusion >>
rect 409 519 410 520 
<< pdiffusion >>
rect 410 519 411 520 
<< pdiffusion >>
rect 411 519 412 520 
<< pdiffusion >>
rect 412 519 413 520 
<< pdiffusion >>
rect 413 519 414 520 
<< pdiffusion >>
rect 426 519 427 520 
<< pdiffusion >>
rect 427 519 428 520 
<< pdiffusion >>
rect 428 519 429 520 
<< pdiffusion >>
rect 429 519 430 520 
<< pdiffusion >>
rect 430 519 431 520 
<< pdiffusion >>
rect 431 519 432 520 
<< pdiffusion >>
rect 444 519 445 520 
<< pdiffusion >>
rect 445 519 446 520 
<< pdiffusion >>
rect 446 519 447 520 
<< pdiffusion >>
rect 447 519 448 520 
<< pdiffusion >>
rect 448 519 449 520 
<< pdiffusion >>
rect 449 519 450 520 
<< m1 >>
rect 451 519 452 520 
<< pdiffusion >>
rect 462 519 463 520 
<< pdiffusion >>
rect 463 519 464 520 
<< pdiffusion >>
rect 464 519 465 520 
<< pdiffusion >>
rect 465 519 466 520 
<< pdiffusion >>
rect 466 519 467 520 
<< pdiffusion >>
rect 467 519 468 520 
<< m1 >>
rect 472 519 473 520 
<< pdiffusion >>
rect 480 519 481 520 
<< pdiffusion >>
rect 481 519 482 520 
<< pdiffusion >>
rect 482 519 483 520 
<< pdiffusion >>
rect 483 519 484 520 
<< pdiffusion >>
rect 484 519 485 520 
<< pdiffusion >>
rect 485 519 486 520 
<< pdiffusion >>
rect 498 519 499 520 
<< pdiffusion >>
rect 499 519 500 520 
<< pdiffusion >>
rect 500 519 501 520 
<< pdiffusion >>
rect 501 519 502 520 
<< pdiffusion >>
rect 502 519 503 520 
<< pdiffusion >>
rect 503 519 504 520 
<< pdiffusion >>
rect 516 519 517 520 
<< pdiffusion >>
rect 517 519 518 520 
<< pdiffusion >>
rect 518 519 519 520 
<< pdiffusion >>
rect 519 519 520 520 
<< pdiffusion >>
rect 520 519 521 520 
<< pdiffusion >>
rect 521 519 522 520 
<< pdiffusion >>
rect 12 520 13 521 
<< pdiffusion >>
rect 13 520 14 521 
<< pdiffusion >>
rect 14 520 15 521 
<< pdiffusion >>
rect 15 520 16 521 
<< pdiffusion >>
rect 16 520 17 521 
<< pdiffusion >>
rect 17 520 18 521 
<< m1 >>
rect 19 520 20 521 
<< pdiffusion >>
rect 30 520 31 521 
<< pdiffusion >>
rect 31 520 32 521 
<< pdiffusion >>
rect 32 520 33 521 
<< pdiffusion >>
rect 33 520 34 521 
<< pdiffusion >>
rect 34 520 35 521 
<< pdiffusion >>
rect 35 520 36 521 
<< pdiffusion >>
rect 48 520 49 521 
<< pdiffusion >>
rect 49 520 50 521 
<< pdiffusion >>
rect 50 520 51 521 
<< pdiffusion >>
rect 51 520 52 521 
<< pdiffusion >>
rect 52 520 53 521 
<< pdiffusion >>
rect 53 520 54 521 
<< pdiffusion >>
rect 66 520 67 521 
<< pdiffusion >>
rect 67 520 68 521 
<< pdiffusion >>
rect 68 520 69 521 
<< pdiffusion >>
rect 69 520 70 521 
<< pdiffusion >>
rect 70 520 71 521 
<< pdiffusion >>
rect 71 520 72 521 
<< pdiffusion >>
rect 84 520 85 521 
<< pdiffusion >>
rect 85 520 86 521 
<< pdiffusion >>
rect 86 520 87 521 
<< pdiffusion >>
rect 87 520 88 521 
<< pdiffusion >>
rect 88 520 89 521 
<< pdiffusion >>
rect 89 520 90 521 
<< m1 >>
rect 100 520 101 521 
<< pdiffusion >>
rect 102 520 103 521 
<< pdiffusion >>
rect 103 520 104 521 
<< pdiffusion >>
rect 104 520 105 521 
<< pdiffusion >>
rect 105 520 106 521 
<< pdiffusion >>
rect 106 520 107 521 
<< pdiffusion >>
rect 107 520 108 521 
<< pdiffusion >>
rect 120 520 121 521 
<< pdiffusion >>
rect 121 520 122 521 
<< pdiffusion >>
rect 122 520 123 521 
<< pdiffusion >>
rect 123 520 124 521 
<< pdiffusion >>
rect 124 520 125 521 
<< pdiffusion >>
rect 125 520 126 521 
<< pdiffusion >>
rect 138 520 139 521 
<< pdiffusion >>
rect 139 520 140 521 
<< pdiffusion >>
rect 140 520 141 521 
<< pdiffusion >>
rect 141 520 142 521 
<< pdiffusion >>
rect 142 520 143 521 
<< pdiffusion >>
rect 143 520 144 521 
<< pdiffusion >>
rect 156 520 157 521 
<< pdiffusion >>
rect 157 520 158 521 
<< pdiffusion >>
rect 158 520 159 521 
<< pdiffusion >>
rect 159 520 160 521 
<< pdiffusion >>
rect 160 520 161 521 
<< pdiffusion >>
rect 161 520 162 521 
<< pdiffusion >>
rect 174 520 175 521 
<< pdiffusion >>
rect 175 520 176 521 
<< pdiffusion >>
rect 176 520 177 521 
<< pdiffusion >>
rect 177 520 178 521 
<< pdiffusion >>
rect 178 520 179 521 
<< pdiffusion >>
rect 179 520 180 521 
<< m1 >>
rect 186 520 187 521 
<< pdiffusion >>
rect 192 520 193 521 
<< pdiffusion >>
rect 193 520 194 521 
<< pdiffusion >>
rect 194 520 195 521 
<< pdiffusion >>
rect 195 520 196 521 
<< pdiffusion >>
rect 196 520 197 521 
<< pdiffusion >>
rect 197 520 198 521 
<< m1 >>
rect 226 520 227 521 
<< pdiffusion >>
rect 228 520 229 521 
<< pdiffusion >>
rect 229 520 230 521 
<< pdiffusion >>
rect 230 520 231 521 
<< pdiffusion >>
rect 231 520 232 521 
<< pdiffusion >>
rect 232 520 233 521 
<< pdiffusion >>
rect 233 520 234 521 
<< pdiffusion >>
rect 246 520 247 521 
<< pdiffusion >>
rect 247 520 248 521 
<< pdiffusion >>
rect 248 520 249 521 
<< pdiffusion >>
rect 249 520 250 521 
<< pdiffusion >>
rect 250 520 251 521 
<< pdiffusion >>
rect 251 520 252 521 
<< m1 >>
rect 262 520 263 521 
<< pdiffusion >>
rect 264 520 265 521 
<< pdiffusion >>
rect 265 520 266 521 
<< pdiffusion >>
rect 266 520 267 521 
<< pdiffusion >>
rect 267 520 268 521 
<< pdiffusion >>
rect 268 520 269 521 
<< pdiffusion >>
rect 269 520 270 521 
<< pdiffusion >>
rect 282 520 283 521 
<< pdiffusion >>
rect 283 520 284 521 
<< pdiffusion >>
rect 284 520 285 521 
<< pdiffusion >>
rect 285 520 286 521 
<< pdiffusion >>
rect 286 520 287 521 
<< pdiffusion >>
rect 287 520 288 521 
<< pdiffusion >>
rect 300 520 301 521 
<< pdiffusion >>
rect 301 520 302 521 
<< pdiffusion >>
rect 302 520 303 521 
<< pdiffusion >>
rect 303 520 304 521 
<< pdiffusion >>
rect 304 520 305 521 
<< pdiffusion >>
rect 305 520 306 521 
<< pdiffusion >>
rect 318 520 319 521 
<< pdiffusion >>
rect 319 520 320 521 
<< pdiffusion >>
rect 320 520 321 521 
<< pdiffusion >>
rect 321 520 322 521 
<< pdiffusion >>
rect 322 520 323 521 
<< pdiffusion >>
rect 323 520 324 521 
<< m1 >>
rect 325 520 326 521 
<< pdiffusion >>
rect 336 520 337 521 
<< pdiffusion >>
rect 337 520 338 521 
<< pdiffusion >>
rect 338 520 339 521 
<< pdiffusion >>
rect 339 520 340 521 
<< pdiffusion >>
rect 340 520 341 521 
<< pdiffusion >>
rect 341 520 342 521 
<< pdiffusion >>
rect 354 520 355 521 
<< pdiffusion >>
rect 355 520 356 521 
<< pdiffusion >>
rect 356 520 357 521 
<< pdiffusion >>
rect 357 520 358 521 
<< pdiffusion >>
rect 358 520 359 521 
<< pdiffusion >>
rect 359 520 360 521 
<< m1 >>
rect 361 520 362 521 
<< m1 >>
rect 370 520 371 521 
<< pdiffusion >>
rect 372 520 373 521 
<< pdiffusion >>
rect 373 520 374 521 
<< pdiffusion >>
rect 374 520 375 521 
<< pdiffusion >>
rect 375 520 376 521 
<< pdiffusion >>
rect 376 520 377 521 
<< pdiffusion >>
rect 377 520 378 521 
<< m1 >>
rect 379 520 380 521 
<< pdiffusion >>
rect 390 520 391 521 
<< pdiffusion >>
rect 391 520 392 521 
<< pdiffusion >>
rect 392 520 393 521 
<< pdiffusion >>
rect 393 520 394 521 
<< pdiffusion >>
rect 394 520 395 521 
<< pdiffusion >>
rect 395 520 396 521 
<< m1 >>
rect 397 520 398 521 
<< pdiffusion >>
rect 408 520 409 521 
<< pdiffusion >>
rect 409 520 410 521 
<< pdiffusion >>
rect 410 520 411 521 
<< pdiffusion >>
rect 411 520 412 521 
<< pdiffusion >>
rect 412 520 413 521 
<< pdiffusion >>
rect 413 520 414 521 
<< pdiffusion >>
rect 426 520 427 521 
<< pdiffusion >>
rect 427 520 428 521 
<< pdiffusion >>
rect 428 520 429 521 
<< pdiffusion >>
rect 429 520 430 521 
<< pdiffusion >>
rect 430 520 431 521 
<< pdiffusion >>
rect 431 520 432 521 
<< pdiffusion >>
rect 444 520 445 521 
<< pdiffusion >>
rect 445 520 446 521 
<< pdiffusion >>
rect 446 520 447 521 
<< pdiffusion >>
rect 447 520 448 521 
<< pdiffusion >>
rect 448 520 449 521 
<< pdiffusion >>
rect 449 520 450 521 
<< m1 >>
rect 451 520 452 521 
<< pdiffusion >>
rect 462 520 463 521 
<< pdiffusion >>
rect 463 520 464 521 
<< pdiffusion >>
rect 464 520 465 521 
<< pdiffusion >>
rect 465 520 466 521 
<< pdiffusion >>
rect 466 520 467 521 
<< pdiffusion >>
rect 467 520 468 521 
<< m1 >>
rect 472 520 473 521 
<< pdiffusion >>
rect 480 520 481 521 
<< pdiffusion >>
rect 481 520 482 521 
<< pdiffusion >>
rect 482 520 483 521 
<< pdiffusion >>
rect 483 520 484 521 
<< pdiffusion >>
rect 484 520 485 521 
<< pdiffusion >>
rect 485 520 486 521 
<< pdiffusion >>
rect 498 520 499 521 
<< pdiffusion >>
rect 499 520 500 521 
<< pdiffusion >>
rect 500 520 501 521 
<< pdiffusion >>
rect 501 520 502 521 
<< pdiffusion >>
rect 502 520 503 521 
<< pdiffusion >>
rect 503 520 504 521 
<< pdiffusion >>
rect 516 520 517 521 
<< pdiffusion >>
rect 517 520 518 521 
<< pdiffusion >>
rect 518 520 519 521 
<< pdiffusion >>
rect 519 520 520 521 
<< pdiffusion >>
rect 520 520 521 521 
<< pdiffusion >>
rect 521 520 522 521 
<< pdiffusion >>
rect 12 521 13 522 
<< pdiffusion >>
rect 13 521 14 522 
<< pdiffusion >>
rect 14 521 15 522 
<< pdiffusion >>
rect 15 521 16 522 
<< m1 >>
rect 16 521 17 522 
<< pdiffusion >>
rect 16 521 17 522 
<< pdiffusion >>
rect 17 521 18 522 
<< m1 >>
rect 19 521 20 522 
<< pdiffusion >>
rect 30 521 31 522 
<< pdiffusion >>
rect 31 521 32 522 
<< pdiffusion >>
rect 32 521 33 522 
<< pdiffusion >>
rect 33 521 34 522 
<< pdiffusion >>
rect 34 521 35 522 
<< pdiffusion >>
rect 35 521 36 522 
<< pdiffusion >>
rect 48 521 49 522 
<< pdiffusion >>
rect 49 521 50 522 
<< pdiffusion >>
rect 50 521 51 522 
<< pdiffusion >>
rect 51 521 52 522 
<< pdiffusion >>
rect 52 521 53 522 
<< pdiffusion >>
rect 53 521 54 522 
<< pdiffusion >>
rect 66 521 67 522 
<< pdiffusion >>
rect 67 521 68 522 
<< pdiffusion >>
rect 68 521 69 522 
<< pdiffusion >>
rect 69 521 70 522 
<< pdiffusion >>
rect 70 521 71 522 
<< pdiffusion >>
rect 71 521 72 522 
<< pdiffusion >>
rect 84 521 85 522 
<< pdiffusion >>
rect 85 521 86 522 
<< pdiffusion >>
rect 86 521 87 522 
<< pdiffusion >>
rect 87 521 88 522 
<< pdiffusion >>
rect 88 521 89 522 
<< pdiffusion >>
rect 89 521 90 522 
<< m1 >>
rect 100 521 101 522 
<< pdiffusion >>
rect 102 521 103 522 
<< m1 >>
rect 103 521 104 522 
<< pdiffusion >>
rect 103 521 104 522 
<< pdiffusion >>
rect 104 521 105 522 
<< pdiffusion >>
rect 105 521 106 522 
<< pdiffusion >>
rect 106 521 107 522 
<< pdiffusion >>
rect 107 521 108 522 
<< pdiffusion >>
rect 120 521 121 522 
<< pdiffusion >>
rect 121 521 122 522 
<< pdiffusion >>
rect 122 521 123 522 
<< pdiffusion >>
rect 123 521 124 522 
<< pdiffusion >>
rect 124 521 125 522 
<< pdiffusion >>
rect 125 521 126 522 
<< pdiffusion >>
rect 138 521 139 522 
<< pdiffusion >>
rect 139 521 140 522 
<< pdiffusion >>
rect 140 521 141 522 
<< pdiffusion >>
rect 141 521 142 522 
<< pdiffusion >>
rect 142 521 143 522 
<< pdiffusion >>
rect 143 521 144 522 
<< pdiffusion >>
rect 156 521 157 522 
<< pdiffusion >>
rect 157 521 158 522 
<< pdiffusion >>
rect 158 521 159 522 
<< pdiffusion >>
rect 159 521 160 522 
<< pdiffusion >>
rect 160 521 161 522 
<< pdiffusion >>
rect 161 521 162 522 
<< pdiffusion >>
rect 174 521 175 522 
<< pdiffusion >>
rect 175 521 176 522 
<< pdiffusion >>
rect 176 521 177 522 
<< pdiffusion >>
rect 177 521 178 522 
<< pdiffusion >>
rect 178 521 179 522 
<< pdiffusion >>
rect 179 521 180 522 
<< m1 >>
rect 186 521 187 522 
<< pdiffusion >>
rect 192 521 193 522 
<< pdiffusion >>
rect 193 521 194 522 
<< pdiffusion >>
rect 194 521 195 522 
<< pdiffusion >>
rect 195 521 196 522 
<< m1 >>
rect 196 521 197 522 
<< pdiffusion >>
rect 196 521 197 522 
<< pdiffusion >>
rect 197 521 198 522 
<< m1 >>
rect 226 521 227 522 
<< pdiffusion >>
rect 228 521 229 522 
<< m1 >>
rect 229 521 230 522 
<< pdiffusion >>
rect 229 521 230 522 
<< pdiffusion >>
rect 230 521 231 522 
<< pdiffusion >>
rect 231 521 232 522 
<< pdiffusion >>
rect 232 521 233 522 
<< pdiffusion >>
rect 233 521 234 522 
<< pdiffusion >>
rect 246 521 247 522 
<< pdiffusion >>
rect 247 521 248 522 
<< pdiffusion >>
rect 248 521 249 522 
<< pdiffusion >>
rect 249 521 250 522 
<< pdiffusion >>
rect 250 521 251 522 
<< pdiffusion >>
rect 251 521 252 522 
<< m1 >>
rect 262 521 263 522 
<< pdiffusion >>
rect 264 521 265 522 
<< m1 >>
rect 265 521 266 522 
<< pdiffusion >>
rect 265 521 266 522 
<< pdiffusion >>
rect 266 521 267 522 
<< pdiffusion >>
rect 267 521 268 522 
<< pdiffusion >>
rect 268 521 269 522 
<< pdiffusion >>
rect 269 521 270 522 
<< pdiffusion >>
rect 282 521 283 522 
<< pdiffusion >>
rect 283 521 284 522 
<< pdiffusion >>
rect 284 521 285 522 
<< pdiffusion >>
rect 285 521 286 522 
<< pdiffusion >>
rect 286 521 287 522 
<< pdiffusion >>
rect 287 521 288 522 
<< pdiffusion >>
rect 300 521 301 522 
<< pdiffusion >>
rect 301 521 302 522 
<< pdiffusion >>
rect 302 521 303 522 
<< pdiffusion >>
rect 303 521 304 522 
<< pdiffusion >>
rect 304 521 305 522 
<< pdiffusion >>
rect 305 521 306 522 
<< pdiffusion >>
rect 318 521 319 522 
<< pdiffusion >>
rect 319 521 320 522 
<< pdiffusion >>
rect 320 521 321 522 
<< pdiffusion >>
rect 321 521 322 522 
<< pdiffusion >>
rect 322 521 323 522 
<< pdiffusion >>
rect 323 521 324 522 
<< m1 >>
rect 325 521 326 522 
<< pdiffusion >>
rect 336 521 337 522 
<< m1 >>
rect 337 521 338 522 
<< pdiffusion >>
rect 337 521 338 522 
<< pdiffusion >>
rect 338 521 339 522 
<< pdiffusion >>
rect 339 521 340 522 
<< pdiffusion >>
rect 340 521 341 522 
<< pdiffusion >>
rect 341 521 342 522 
<< pdiffusion >>
rect 354 521 355 522 
<< pdiffusion >>
rect 355 521 356 522 
<< pdiffusion >>
rect 356 521 357 522 
<< pdiffusion >>
rect 357 521 358 522 
<< pdiffusion >>
rect 358 521 359 522 
<< pdiffusion >>
rect 359 521 360 522 
<< m1 >>
rect 361 521 362 522 
<< m1 >>
rect 370 521 371 522 
<< pdiffusion >>
rect 372 521 373 522 
<< pdiffusion >>
rect 373 521 374 522 
<< pdiffusion >>
rect 374 521 375 522 
<< pdiffusion >>
rect 375 521 376 522 
<< pdiffusion >>
rect 376 521 377 522 
<< pdiffusion >>
rect 377 521 378 522 
<< m1 >>
rect 379 521 380 522 
<< pdiffusion >>
rect 390 521 391 522 
<< pdiffusion >>
rect 391 521 392 522 
<< pdiffusion >>
rect 392 521 393 522 
<< pdiffusion >>
rect 393 521 394 522 
<< pdiffusion >>
rect 394 521 395 522 
<< pdiffusion >>
rect 395 521 396 522 
<< m1 >>
rect 397 521 398 522 
<< pdiffusion >>
rect 408 521 409 522 
<< pdiffusion >>
rect 409 521 410 522 
<< pdiffusion >>
rect 410 521 411 522 
<< pdiffusion >>
rect 411 521 412 522 
<< m1 >>
rect 412 521 413 522 
<< pdiffusion >>
rect 412 521 413 522 
<< pdiffusion >>
rect 413 521 414 522 
<< pdiffusion >>
rect 426 521 427 522 
<< pdiffusion >>
rect 427 521 428 522 
<< pdiffusion >>
rect 428 521 429 522 
<< pdiffusion >>
rect 429 521 430 522 
<< m1 >>
rect 430 521 431 522 
<< pdiffusion >>
rect 430 521 431 522 
<< pdiffusion >>
rect 431 521 432 522 
<< pdiffusion >>
rect 444 521 445 522 
<< pdiffusion >>
rect 445 521 446 522 
<< pdiffusion >>
rect 446 521 447 522 
<< pdiffusion >>
rect 447 521 448 522 
<< pdiffusion >>
rect 448 521 449 522 
<< pdiffusion >>
rect 449 521 450 522 
<< m1 >>
rect 451 521 452 522 
<< pdiffusion >>
rect 462 521 463 522 
<< m1 >>
rect 463 521 464 522 
<< pdiffusion >>
rect 463 521 464 522 
<< pdiffusion >>
rect 464 521 465 522 
<< pdiffusion >>
rect 465 521 466 522 
<< pdiffusion >>
rect 466 521 467 522 
<< pdiffusion >>
rect 467 521 468 522 
<< m1 >>
rect 472 521 473 522 
<< pdiffusion >>
rect 480 521 481 522 
<< m1 >>
rect 481 521 482 522 
<< pdiffusion >>
rect 481 521 482 522 
<< pdiffusion >>
rect 482 521 483 522 
<< pdiffusion >>
rect 483 521 484 522 
<< pdiffusion >>
rect 484 521 485 522 
<< pdiffusion >>
rect 485 521 486 522 
<< pdiffusion >>
rect 498 521 499 522 
<< pdiffusion >>
rect 499 521 500 522 
<< pdiffusion >>
rect 500 521 501 522 
<< pdiffusion >>
rect 501 521 502 522 
<< pdiffusion >>
rect 502 521 503 522 
<< pdiffusion >>
rect 503 521 504 522 
<< pdiffusion >>
rect 516 521 517 522 
<< pdiffusion >>
rect 517 521 518 522 
<< pdiffusion >>
rect 518 521 519 522 
<< pdiffusion >>
rect 519 521 520 522 
<< pdiffusion >>
rect 520 521 521 522 
<< pdiffusion >>
rect 521 521 522 522 
<< m1 >>
rect 16 522 17 523 
<< m1 >>
rect 19 522 20 523 
<< m1 >>
rect 100 522 101 523 
<< m1 >>
rect 103 522 104 523 
<< m1 >>
rect 186 522 187 523 
<< m1 >>
rect 196 522 197 523 
<< m1 >>
rect 226 522 227 523 
<< m1 >>
rect 229 522 230 523 
<< m1 >>
rect 262 522 263 523 
<< m1 >>
rect 265 522 266 523 
<< m1 >>
rect 325 522 326 523 
<< m1 >>
rect 337 522 338 523 
<< m1 >>
rect 361 522 362 523 
<< m1 >>
rect 370 522 371 523 
<< m1 >>
rect 379 522 380 523 
<< m1 >>
rect 397 522 398 523 
<< m1 >>
rect 412 522 413 523 
<< m1 >>
rect 430 522 431 523 
<< m1 >>
rect 451 522 452 523 
<< m1 >>
rect 463 522 464 523 
<< m1 >>
rect 472 522 473 523 
<< m1 >>
rect 481 522 482 523 
<< m1 >>
rect 16 523 17 524 
<< m1 >>
rect 17 523 18 524 
<< m1 >>
rect 18 523 19 524 
<< m1 >>
rect 19 523 20 524 
<< m1 >>
rect 100 523 101 524 
<< m1 >>
rect 101 523 102 524 
<< m1 >>
rect 102 523 103 524 
<< m1 >>
rect 103 523 104 524 
<< m1 >>
rect 186 523 187 524 
<< m1 >>
rect 196 523 197 524 
<< m1 >>
rect 226 523 227 524 
<< m1 >>
rect 227 523 228 524 
<< m1 >>
rect 228 523 229 524 
<< m1 >>
rect 229 523 230 524 
<< m1 >>
rect 262 523 263 524 
<< m1 >>
rect 263 523 264 524 
<< m1 >>
rect 264 523 265 524 
<< m1 >>
rect 265 523 266 524 
<< m1 >>
rect 325 523 326 524 
<< m1 >>
rect 326 523 327 524 
<< m1 >>
rect 327 523 328 524 
<< m1 >>
rect 328 523 329 524 
<< m1 >>
rect 329 523 330 524 
<< m1 >>
rect 330 523 331 524 
<< m1 >>
rect 331 523 332 524 
<< m1 >>
rect 332 523 333 524 
<< m1 >>
rect 333 523 334 524 
<< m1 >>
rect 334 523 335 524 
<< m1 >>
rect 335 523 336 524 
<< m1 >>
rect 336 523 337 524 
<< m1 >>
rect 337 523 338 524 
<< m1 >>
rect 361 523 362 524 
<< m1 >>
rect 370 523 371 524 
<< m1 >>
rect 379 523 380 524 
<< m1 >>
rect 397 523 398 524 
<< m1 >>
rect 412 523 413 524 
<< m1 >>
rect 430 523 431 524 
<< m1 >>
rect 451 523 452 524 
<< m1 >>
rect 452 523 453 524 
<< m1 >>
rect 453 523 454 524 
<< m1 >>
rect 454 523 455 524 
<< m1 >>
rect 455 523 456 524 
<< m1 >>
rect 456 523 457 524 
<< m1 >>
rect 457 523 458 524 
<< m1 >>
rect 458 523 459 524 
<< m1 >>
rect 459 523 460 524 
<< m1 >>
rect 460 523 461 524 
<< m1 >>
rect 461 523 462 524 
<< m1 >>
rect 462 523 463 524 
<< m1 >>
rect 463 523 464 524 
<< m1 >>
rect 472 523 473 524 
<< m1 >>
rect 473 523 474 524 
<< m1 >>
rect 474 523 475 524 
<< m1 >>
rect 475 523 476 524 
<< m1 >>
rect 476 523 477 524 
<< m1 >>
rect 477 523 478 524 
<< m1 >>
rect 478 523 479 524 
<< m1 >>
rect 479 523 480 524 
<< m1 >>
rect 480 523 481 524 
<< m1 >>
rect 481 523 482 524 
<< m1 >>
rect 186 524 187 525 
<< m1 >>
rect 196 524 197 525 
<< m1 >>
rect 361 524 362 525 
<< m1 >>
rect 370 524 371 525 
<< m1 >>
rect 379 524 380 525 
<< m1 >>
rect 392 524 393 525 
<< m2 >>
rect 392 524 393 525 
<< m2c >>
rect 392 524 393 525 
<< m1 >>
rect 392 524 393 525 
<< m2 >>
rect 392 524 393 525 
<< m1 >>
rect 393 524 394 525 
<< m1 >>
rect 394 524 395 525 
<< m1 >>
rect 395 524 396 525 
<< m1 >>
rect 396 524 397 525 
<< m1 >>
rect 397 524 398 525 
<< m1 >>
rect 412 524 413 525 
<< m1 >>
rect 430 524 431 525 
<< m1 >>
rect 186 525 187 526 
<< m1 >>
rect 196 525 197 526 
<< m1 >>
rect 361 525 362 526 
<< m1 >>
rect 370 525 371 526 
<< m1 >>
rect 379 525 380 526 
<< m2 >>
rect 392 525 393 526 
<< m1 >>
rect 412 525 413 526 
<< m1 >>
rect 430 525 431 526 
<< m1 >>
rect 186 526 187 527 
<< m1 >>
rect 187 526 188 527 
<< m1 >>
rect 188 526 189 527 
<< m1 >>
rect 189 526 190 527 
<< m1 >>
rect 190 526 191 527 
<< m1 >>
rect 191 526 192 527 
<< m1 >>
rect 192 526 193 527 
<< m1 >>
rect 193 526 194 527 
<< m1 >>
rect 194 526 195 527 
<< m1 >>
rect 195 526 196 527 
<< m1 >>
rect 196 526 197 527 
<< m1 >>
rect 361 526 362 527 
<< m1 >>
rect 370 526 371 527 
<< m1 >>
rect 371 526 372 527 
<< m1 >>
rect 372 526 373 527 
<< m1 >>
rect 373 526 374 527 
<< m1 >>
rect 374 526 375 527 
<< m1 >>
rect 375 526 376 527 
<< m1 >>
rect 376 526 377 527 
<< m1 >>
rect 377 526 378 527 
<< m2 >>
rect 377 526 378 527 
<< m2c >>
rect 377 526 378 527 
<< m1 >>
rect 377 526 378 527 
<< m2 >>
rect 377 526 378 527 
<< m2 >>
rect 378 526 379 527 
<< m1 >>
rect 379 526 380 527 
<< m2 >>
rect 379 526 380 527 
<< m1 >>
rect 380 526 381 527 
<< m2 >>
rect 380 526 381 527 
<< m1 >>
rect 381 526 382 527 
<< m2 >>
rect 381 526 382 527 
<< m1 >>
rect 382 526 383 527 
<< m2 >>
rect 382 526 383 527 
<< m1 >>
rect 383 526 384 527 
<< m2 >>
rect 383 526 384 527 
<< m1 >>
rect 384 526 385 527 
<< m2 >>
rect 384 526 385 527 
<< m1 >>
rect 385 526 386 527 
<< m2 >>
rect 385 526 386 527 
<< m1 >>
rect 386 526 387 527 
<< m2 >>
rect 386 526 387 527 
<< m1 >>
rect 387 526 388 527 
<< m2 >>
rect 387 526 388 527 
<< m1 >>
rect 388 526 389 527 
<< m2 >>
rect 388 526 389 527 
<< m1 >>
rect 389 526 390 527 
<< m2 >>
rect 389 526 390 527 
<< m1 >>
rect 390 526 391 527 
<< m2 >>
rect 390 526 391 527 
<< m1 >>
rect 391 526 392 527 
<< m2 >>
rect 391 526 392 527 
<< m1 >>
rect 392 526 393 527 
<< m2 >>
rect 392 526 393 527 
<< m1 >>
rect 393 526 394 527 
<< m1 >>
rect 394 526 395 527 
<< m1 >>
rect 395 526 396 527 
<< m1 >>
rect 396 526 397 527 
<< m1 >>
rect 397 526 398 527 
<< m1 >>
rect 398 526 399 527 
<< m1 >>
rect 399 526 400 527 
<< m1 >>
rect 400 526 401 527 
<< m1 >>
rect 401 526 402 527 
<< m1 >>
rect 402 526 403 527 
<< m1 >>
rect 403 526 404 527 
<< m1 >>
rect 404 526 405 527 
<< m1 >>
rect 405 526 406 527 
<< m1 >>
rect 406 526 407 527 
<< m1 >>
rect 407 526 408 527 
<< m1 >>
rect 408 526 409 527 
<< m1 >>
rect 409 526 410 527 
<< m1 >>
rect 410 526 411 527 
<< m1 >>
rect 411 526 412 527 
<< m1 >>
rect 412 526 413 527 
<< m1 >>
rect 430 526 431 527 
<< m1 >>
rect 361 527 362 528 
<< m1 >>
rect 430 527 431 528 
<< m1 >>
rect 361 528 362 529 
<< m1 >>
rect 362 528 363 529 
<< m1 >>
rect 363 528 364 529 
<< m1 >>
rect 364 528 365 529 
<< m1 >>
rect 365 528 366 529 
<< m1 >>
rect 366 528 367 529 
<< m1 >>
rect 367 528 368 529 
<< m1 >>
rect 368 528 369 529 
<< m1 >>
rect 369 528 370 529 
<< m1 >>
rect 370 528 371 529 
<< m1 >>
rect 371 528 372 529 
<< m1 >>
rect 372 528 373 529 
<< m1 >>
rect 373 528 374 529 
<< m1 >>
rect 374 528 375 529 
<< m1 >>
rect 375 528 376 529 
<< m1 >>
rect 376 528 377 529 
<< m1 >>
rect 377 528 378 529 
<< m1 >>
rect 378 528 379 529 
<< m1 >>
rect 379 528 380 529 
<< m1 >>
rect 380 528 381 529 
<< m1 >>
rect 381 528 382 529 
<< m1 >>
rect 382 528 383 529 
<< m1 >>
rect 383 528 384 529 
<< m1 >>
rect 384 528 385 529 
<< m1 >>
rect 385 528 386 529 
<< m1 >>
rect 386 528 387 529 
<< m1 >>
rect 387 528 388 529 
<< m1 >>
rect 388 528 389 529 
<< m1 >>
rect 389 528 390 529 
<< m1 >>
rect 390 528 391 529 
<< m1 >>
rect 391 528 392 529 
<< m1 >>
rect 392 528 393 529 
<< m1 >>
rect 393 528 394 529 
<< m1 >>
rect 394 528 395 529 
<< m1 >>
rect 395 528 396 529 
<< m1 >>
rect 396 528 397 529 
<< m1 >>
rect 397 528 398 529 
<< m1 >>
rect 398 528 399 529 
<< m1 >>
rect 399 528 400 529 
<< m1 >>
rect 400 528 401 529 
<< m1 >>
rect 401 528 402 529 
<< m1 >>
rect 402 528 403 529 
<< m1 >>
rect 403 528 404 529 
<< m1 >>
rect 404 528 405 529 
<< m1 >>
rect 405 528 406 529 
<< m1 >>
rect 406 528 407 529 
<< m1 >>
rect 407 528 408 529 
<< m1 >>
rect 408 528 409 529 
<< m1 >>
rect 409 528 410 529 
<< m1 >>
rect 410 528 411 529 
<< m1 >>
rect 411 528 412 529 
<< m1 >>
rect 412 528 413 529 
<< m1 >>
rect 413 528 414 529 
<< m1 >>
rect 414 528 415 529 
<< m1 >>
rect 415 528 416 529 
<< m1 >>
rect 416 528 417 529 
<< m1 >>
rect 417 528 418 529 
<< m1 >>
rect 418 528 419 529 
<< m1 >>
rect 419 528 420 529 
<< m1 >>
rect 420 528 421 529 
<< m1 >>
rect 421 528 422 529 
<< m1 >>
rect 422 528 423 529 
<< m1 >>
rect 423 528 424 529 
<< m1 >>
rect 424 528 425 529 
<< m1 >>
rect 425 528 426 529 
<< m1 >>
rect 426 528 427 529 
<< m1 >>
rect 427 528 428 529 
<< m1 >>
rect 428 528 429 529 
<< m1 >>
rect 429 528 430 529 
<< m1 >>
rect 430 528 431 529 
<< labels >>
rlabel pdiffusion 391 192 392 193  0 t = 1
rlabel pdiffusion 394 192 395 193  0 t = 2
rlabel pdiffusion 391 197 392 198  0 t = 3
rlabel pdiffusion 394 197 395 198  0 t = 4
rlabel pdiffusion 390 192 396 198 0 cell no = 1
<< m1 >>
rect 391 192 392 193 
rect 394 192 395 193 
rect 391 197 392 198 
rect 394 197 395 198 
<< m2 >>
rect 391 192 392 193 
rect 394 192 395 193 
rect 391 197 392 198 
rect 394 197 395 198 
<< m2c >>
rect 391 192 392 193 
rect 394 192 395 193 
rect 391 197 392 198 
rect 394 197 395 198 
<< labels >>
rlabel pdiffusion 49 138 50 139  0 t = 1
rlabel pdiffusion 52 138 53 139  0 t = 2
rlabel pdiffusion 49 143 50 144  0 t = 3
rlabel pdiffusion 52 143 53 144  0 t = 4
rlabel pdiffusion 48 138 54 144 0 cell no = 2
<< m1 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2 >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< m2c >>
rect 49 138 50 139 
rect 52 138 53 139 
rect 49 143 50 144 
rect 52 143 53 144 
<< labels >>
rlabel pdiffusion 103 156 104 157  0 t = 1
rlabel pdiffusion 106 156 107 157  0 t = 2
rlabel pdiffusion 103 161 104 162  0 t = 3
rlabel pdiffusion 106 161 107 162  0 t = 4
rlabel pdiffusion 102 156 108 162 0 cell no = 3
<< m1 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2 >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< m2c >>
rect 103 156 104 157 
rect 106 156 107 157 
rect 103 161 104 162 
rect 106 161 107 162 
<< labels >>
rlabel pdiffusion 103 516 104 517  0 t = 1
rlabel pdiffusion 106 516 107 517  0 t = 2
rlabel pdiffusion 103 521 104 522  0 t = 3
rlabel pdiffusion 106 521 107 522  0 t = 4
rlabel pdiffusion 102 516 108 522 0 cell no = 4
<< m1 >>
rect 103 516 104 517 
rect 106 516 107 517 
rect 103 521 104 522 
rect 106 521 107 522 
<< m2 >>
rect 103 516 104 517 
rect 106 516 107 517 
rect 103 521 104 522 
rect 106 521 107 522 
<< m2c >>
rect 103 516 104 517 
rect 106 516 107 517 
rect 103 521 104 522 
rect 106 521 107 522 
<< labels >>
rlabel pdiffusion 139 12 140 13  0 t = 1
rlabel pdiffusion 142 12 143 13  0 t = 2
rlabel pdiffusion 139 17 140 18  0 t = 3
rlabel pdiffusion 142 17 143 18  0 t = 4
rlabel pdiffusion 138 12 144 18 0 cell no = 5
<< m1 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2 >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< m2c >>
rect 139 12 140 13 
rect 142 12 143 13 
rect 139 17 140 18 
rect 142 17 143 18 
<< labels >>
rlabel pdiffusion 247 12 248 13  0 t = 1
rlabel pdiffusion 250 12 251 13  0 t = 2
rlabel pdiffusion 247 17 248 18  0 t = 3
rlabel pdiffusion 250 17 251 18  0 t = 4
rlabel pdiffusion 246 12 252 18 0 cell no = 6
<< m1 >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< m2 >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< m2c >>
rect 247 12 248 13 
rect 250 12 251 13 
rect 247 17 248 18 
rect 250 17 251 18 
<< labels >>
rlabel pdiffusion 31 84 32 85  0 t = 1
rlabel pdiffusion 34 84 35 85  0 t = 2
rlabel pdiffusion 31 89 32 90  0 t = 3
rlabel pdiffusion 34 89 35 90  0 t = 4
rlabel pdiffusion 30 84 36 90 0 cell no = 7
<< m1 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2 >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< m2c >>
rect 31 84 32 85 
rect 34 84 35 85 
rect 31 89 32 90 
rect 34 89 35 90 
<< labels >>
rlabel pdiffusion 13 84 14 85  0 t = 1
rlabel pdiffusion 16 84 17 85  0 t = 2
rlabel pdiffusion 13 89 14 90  0 t = 3
rlabel pdiffusion 16 89 17 90  0 t = 4
rlabel pdiffusion 12 84 18 90 0 cell no = 8
<< m1 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2 >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< m2c >>
rect 13 84 14 85 
rect 16 84 17 85 
rect 13 89 14 90 
rect 16 89 17 90 
<< labels >>
rlabel pdiffusion 49 228 50 229  0 t = 1
rlabel pdiffusion 52 228 53 229  0 t = 2
rlabel pdiffusion 49 233 50 234  0 t = 3
rlabel pdiffusion 52 233 53 234  0 t = 4
rlabel pdiffusion 48 228 54 234 0 cell no = 9
<< m1 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2 >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< m2c >>
rect 49 228 50 229 
rect 52 228 53 229 
rect 49 233 50 234 
rect 52 233 53 234 
<< labels >>
rlabel pdiffusion 157 102 158 103  0 t = 1
rlabel pdiffusion 160 102 161 103  0 t = 2
rlabel pdiffusion 157 107 158 108  0 t = 3
rlabel pdiffusion 160 107 161 108  0 t = 4
rlabel pdiffusion 156 102 162 108 0 cell no = 10
<< m1 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2 >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< m2c >>
rect 157 102 158 103 
rect 160 102 161 103 
rect 157 107 158 108 
rect 160 107 161 108 
<< labels >>
rlabel pdiffusion 391 120 392 121  0 t = 1
rlabel pdiffusion 394 120 395 121  0 t = 2
rlabel pdiffusion 391 125 392 126  0 t = 3
rlabel pdiffusion 394 125 395 126  0 t = 4
rlabel pdiffusion 390 120 396 126 0 cell no = 11
<< m1 >>
rect 391 120 392 121 
rect 394 120 395 121 
rect 391 125 392 126 
rect 394 125 395 126 
<< m2 >>
rect 391 120 392 121 
rect 394 120 395 121 
rect 391 125 392 126 
rect 394 125 395 126 
<< m2c >>
rect 391 120 392 121 
rect 394 120 395 121 
rect 391 125 392 126 
rect 394 125 395 126 
<< labels >>
rlabel pdiffusion 355 84 356 85  0 t = 1
rlabel pdiffusion 358 84 359 85  0 t = 2
rlabel pdiffusion 355 89 356 90  0 t = 3
rlabel pdiffusion 358 89 359 90  0 t = 4
rlabel pdiffusion 354 84 360 90 0 cell no = 12
<< m1 >>
rect 355 84 356 85 
rect 358 84 359 85 
rect 355 89 356 90 
rect 358 89 359 90 
<< m2 >>
rect 355 84 356 85 
rect 358 84 359 85 
rect 355 89 356 90 
rect 358 89 359 90 
<< m2c >>
rect 355 84 356 85 
rect 358 84 359 85 
rect 355 89 356 90 
rect 358 89 359 90 
<< labels >>
rlabel pdiffusion 247 48 248 49  0 t = 1
rlabel pdiffusion 250 48 251 49  0 t = 2
rlabel pdiffusion 247 53 248 54  0 t = 3
rlabel pdiffusion 250 53 251 54  0 t = 4
rlabel pdiffusion 246 48 252 54 0 cell no = 13
<< m1 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2 >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< m2c >>
rect 247 48 248 49 
rect 250 48 251 49 
rect 247 53 248 54 
rect 250 53 251 54 
<< labels >>
rlabel pdiffusion 427 12 428 13  0 t = 1
rlabel pdiffusion 430 12 431 13  0 t = 2
rlabel pdiffusion 427 17 428 18  0 t = 3
rlabel pdiffusion 430 17 431 18  0 t = 4
rlabel pdiffusion 426 12 432 18 0 cell no = 14
<< m1 >>
rect 427 12 428 13 
rect 430 12 431 13 
rect 427 17 428 18 
rect 430 17 431 18 
<< m2 >>
rect 427 12 428 13 
rect 430 12 431 13 
rect 427 17 428 18 
rect 430 17 431 18 
<< m2c >>
rect 427 12 428 13 
rect 430 12 431 13 
rect 427 17 428 18 
rect 430 17 431 18 
<< labels >>
rlabel pdiffusion 319 12 320 13  0 t = 1
rlabel pdiffusion 322 12 323 13  0 t = 2
rlabel pdiffusion 319 17 320 18  0 t = 3
rlabel pdiffusion 322 17 323 18  0 t = 4
rlabel pdiffusion 318 12 324 18 0 cell no = 15
<< m1 >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< m2 >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< m2c >>
rect 319 12 320 13 
rect 322 12 323 13 
rect 319 17 320 18 
rect 322 17 323 18 
<< labels >>
rlabel pdiffusion 373 12 374 13  0 t = 1
rlabel pdiffusion 376 12 377 13  0 t = 2
rlabel pdiffusion 373 17 374 18  0 t = 3
rlabel pdiffusion 376 17 377 18  0 t = 4
rlabel pdiffusion 372 12 378 18 0 cell no = 16
<< m1 >>
rect 373 12 374 13 
rect 376 12 377 13 
rect 373 17 374 18 
rect 376 17 377 18 
<< m2 >>
rect 373 12 374 13 
rect 376 12 377 13 
rect 373 17 374 18 
rect 376 17 377 18 
<< m2c >>
rect 373 12 374 13 
rect 376 12 377 13 
rect 373 17 374 18 
rect 376 17 377 18 
<< labels >>
rlabel pdiffusion 319 48 320 49  0 t = 1
rlabel pdiffusion 322 48 323 49  0 t = 2
rlabel pdiffusion 319 53 320 54  0 t = 3
rlabel pdiffusion 322 53 323 54  0 t = 4
rlabel pdiffusion 318 48 324 54 0 cell no = 17
<< m1 >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< m2 >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< m2c >>
rect 319 48 320 49 
rect 322 48 323 49 
rect 319 53 320 54 
rect 322 53 323 54 
<< labels >>
rlabel pdiffusion 265 102 266 103  0 t = 1
rlabel pdiffusion 268 102 269 103  0 t = 2
rlabel pdiffusion 265 107 266 108  0 t = 3
rlabel pdiffusion 268 107 269 108  0 t = 4
rlabel pdiffusion 264 102 270 108 0 cell no = 18
<< m1 >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< m2 >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< m2c >>
rect 265 102 266 103 
rect 268 102 269 103 
rect 265 107 266 108 
rect 268 107 269 108 
<< labels >>
rlabel pdiffusion 391 12 392 13  0 t = 1
rlabel pdiffusion 394 12 395 13  0 t = 2
rlabel pdiffusion 391 17 392 18  0 t = 3
rlabel pdiffusion 394 17 395 18  0 t = 4
rlabel pdiffusion 390 12 396 18 0 cell no = 19
<< m1 >>
rect 391 12 392 13 
rect 394 12 395 13 
rect 391 17 392 18 
rect 394 17 395 18 
<< m2 >>
rect 391 12 392 13 
rect 394 12 395 13 
rect 391 17 392 18 
rect 394 17 395 18 
<< m2c >>
rect 391 12 392 13 
rect 394 12 395 13 
rect 391 17 392 18 
rect 394 17 395 18 
<< labels >>
rlabel pdiffusion 193 138 194 139  0 t = 1
rlabel pdiffusion 196 138 197 139  0 t = 2
rlabel pdiffusion 193 143 194 144  0 t = 3
rlabel pdiffusion 196 143 197 144  0 t = 4
rlabel pdiffusion 192 138 198 144 0 cell no = 20
<< m1 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2 >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< m2c >>
rect 193 138 194 139 
rect 196 138 197 139 
rect 193 143 194 144 
rect 196 143 197 144 
<< labels >>
rlabel pdiffusion 409 30 410 31  0 t = 1
rlabel pdiffusion 412 30 413 31  0 t = 2
rlabel pdiffusion 409 35 410 36  0 t = 3
rlabel pdiffusion 412 35 413 36  0 t = 4
rlabel pdiffusion 408 30 414 36 0 cell no = 21
<< m1 >>
rect 409 30 410 31 
rect 412 30 413 31 
rect 409 35 410 36 
rect 412 35 413 36 
<< m2 >>
rect 409 30 410 31 
rect 412 30 413 31 
rect 409 35 410 36 
rect 412 35 413 36 
<< m2c >>
rect 409 30 410 31 
rect 412 30 413 31 
rect 409 35 410 36 
rect 412 35 413 36 
<< labels >>
rlabel pdiffusion 445 48 446 49  0 t = 1
rlabel pdiffusion 448 48 449 49  0 t = 2
rlabel pdiffusion 445 53 446 54  0 t = 3
rlabel pdiffusion 448 53 449 54  0 t = 4
rlabel pdiffusion 444 48 450 54 0 cell no = 22
<< m1 >>
rect 445 48 446 49 
rect 448 48 449 49 
rect 445 53 446 54 
rect 448 53 449 54 
<< m2 >>
rect 445 48 446 49 
rect 448 48 449 49 
rect 445 53 446 54 
rect 448 53 449 54 
<< m2c >>
rect 445 48 446 49 
rect 448 48 449 49 
rect 445 53 446 54 
rect 448 53 449 54 
<< labels >>
rlabel pdiffusion 481 102 482 103  0 t = 1
rlabel pdiffusion 484 102 485 103  0 t = 2
rlabel pdiffusion 481 107 482 108  0 t = 3
rlabel pdiffusion 484 107 485 108  0 t = 4
rlabel pdiffusion 480 102 486 108 0 cell no = 23
<< m1 >>
rect 481 102 482 103 
rect 484 102 485 103 
rect 481 107 482 108 
rect 484 107 485 108 
<< m2 >>
rect 481 102 482 103 
rect 484 102 485 103 
rect 481 107 482 108 
rect 484 107 485 108 
<< m2c >>
rect 481 102 482 103 
rect 484 102 485 103 
rect 481 107 482 108 
rect 484 107 485 108 
<< labels >>
rlabel pdiffusion 445 30 446 31  0 t = 1
rlabel pdiffusion 448 30 449 31  0 t = 2
rlabel pdiffusion 445 35 446 36  0 t = 3
rlabel pdiffusion 448 35 449 36  0 t = 4
rlabel pdiffusion 444 30 450 36 0 cell no = 24
<< m1 >>
rect 445 30 446 31 
rect 448 30 449 31 
rect 445 35 446 36 
rect 448 35 449 36 
<< m2 >>
rect 445 30 446 31 
rect 448 30 449 31 
rect 445 35 446 36 
rect 448 35 449 36 
<< m2c >>
rect 445 30 446 31 
rect 448 30 449 31 
rect 445 35 446 36 
rect 448 35 449 36 
<< labels >>
rlabel pdiffusion 391 30 392 31  0 t = 1
rlabel pdiffusion 394 30 395 31  0 t = 2
rlabel pdiffusion 391 35 392 36  0 t = 3
rlabel pdiffusion 394 35 395 36  0 t = 4
rlabel pdiffusion 390 30 396 36 0 cell no = 25
<< m1 >>
rect 391 30 392 31 
rect 394 30 395 31 
rect 391 35 392 36 
rect 394 35 395 36 
<< m2 >>
rect 391 30 392 31 
rect 394 30 395 31 
rect 391 35 392 36 
rect 394 35 395 36 
<< m2c >>
rect 391 30 392 31 
rect 394 30 395 31 
rect 391 35 392 36 
rect 394 35 395 36 
<< labels >>
rlabel pdiffusion 283 336 284 337  0 t = 1
rlabel pdiffusion 286 336 287 337  0 t = 2
rlabel pdiffusion 283 341 284 342  0 t = 3
rlabel pdiffusion 286 341 287 342  0 t = 4
rlabel pdiffusion 282 336 288 342 0 cell no = 26
<< m1 >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< m2 >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< m2c >>
rect 283 336 284 337 
rect 286 336 287 337 
rect 283 341 284 342 
rect 286 341 287 342 
<< labels >>
rlabel pdiffusion 355 138 356 139  0 t = 1
rlabel pdiffusion 358 138 359 139  0 t = 2
rlabel pdiffusion 355 143 356 144  0 t = 3
rlabel pdiffusion 358 143 359 144  0 t = 4
rlabel pdiffusion 354 138 360 144 0 cell no = 27
<< m1 >>
rect 355 138 356 139 
rect 358 138 359 139 
rect 355 143 356 144 
rect 358 143 359 144 
<< m2 >>
rect 355 138 356 139 
rect 358 138 359 139 
rect 355 143 356 144 
rect 358 143 359 144 
<< m2c >>
rect 355 138 356 139 
rect 358 138 359 139 
rect 355 143 356 144 
rect 358 143 359 144 
<< labels >>
rlabel pdiffusion 499 156 500 157  0 t = 1
rlabel pdiffusion 502 156 503 157  0 t = 2
rlabel pdiffusion 499 161 500 162  0 t = 3
rlabel pdiffusion 502 161 503 162  0 t = 4
rlabel pdiffusion 498 156 504 162 0 cell no = 28
<< m1 >>
rect 499 156 500 157 
rect 502 156 503 157 
rect 499 161 500 162 
rect 502 161 503 162 
<< m2 >>
rect 499 156 500 157 
rect 502 156 503 157 
rect 499 161 500 162 
rect 502 161 503 162 
<< m2c >>
rect 499 156 500 157 
rect 502 156 503 157 
rect 499 161 500 162 
rect 502 161 503 162 
<< labels >>
rlabel pdiffusion 49 102 50 103  0 t = 1
rlabel pdiffusion 52 102 53 103  0 t = 2
rlabel pdiffusion 49 107 50 108  0 t = 3
rlabel pdiffusion 52 107 53 108  0 t = 4
rlabel pdiffusion 48 102 54 108 0 cell no = 29
<< m1 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2 >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< m2c >>
rect 49 102 50 103 
rect 52 102 53 103 
rect 49 107 50 108 
rect 52 107 53 108 
<< labels >>
rlabel pdiffusion 49 30 50 31  0 t = 1
rlabel pdiffusion 52 30 53 31  0 t = 2
rlabel pdiffusion 49 35 50 36  0 t = 3
rlabel pdiffusion 52 35 53 36  0 t = 4
rlabel pdiffusion 48 30 54 36 0 cell no = 30
<< m1 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2 >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< m2c >>
rect 49 30 50 31 
rect 52 30 53 31 
rect 49 35 50 36 
rect 52 35 53 36 
<< labels >>
rlabel pdiffusion 13 174 14 175  0 t = 1
rlabel pdiffusion 16 174 17 175  0 t = 2
rlabel pdiffusion 13 179 14 180  0 t = 3
rlabel pdiffusion 16 179 17 180  0 t = 4
rlabel pdiffusion 12 174 18 180 0 cell no = 31
<< m1 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2 >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< m2c >>
rect 13 174 14 175 
rect 16 174 17 175 
rect 13 179 14 180 
rect 16 179 17 180 
<< labels >>
rlabel pdiffusion 67 48 68 49  0 t = 1
rlabel pdiffusion 70 48 71 49  0 t = 2
rlabel pdiffusion 67 53 68 54  0 t = 3
rlabel pdiffusion 70 53 71 54  0 t = 4
rlabel pdiffusion 66 48 72 54 0 cell no = 32
<< m1 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2 >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< m2c >>
rect 67 48 68 49 
rect 70 48 71 49 
rect 67 53 68 54 
rect 70 53 71 54 
<< labels >>
rlabel pdiffusion 103 66 104 67  0 t = 1
rlabel pdiffusion 106 66 107 67  0 t = 2
rlabel pdiffusion 103 71 104 72  0 t = 3
rlabel pdiffusion 106 71 107 72  0 t = 4
rlabel pdiffusion 102 66 108 72 0 cell no = 33
<< m1 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2 >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< m2c >>
rect 103 66 104 67 
rect 106 66 107 67 
rect 103 71 104 72 
rect 106 71 107 72 
<< labels >>
rlabel pdiffusion 103 30 104 31  0 t = 1
rlabel pdiffusion 106 30 107 31  0 t = 2
rlabel pdiffusion 103 35 104 36  0 t = 3
rlabel pdiffusion 106 35 107 36  0 t = 4
rlabel pdiffusion 102 30 108 36 0 cell no = 34
<< m1 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2 >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< m2c >>
rect 103 30 104 31 
rect 106 30 107 31 
rect 103 35 104 36 
rect 106 35 107 36 
<< labels >>
rlabel pdiffusion 157 66 158 67  0 t = 1
rlabel pdiffusion 160 66 161 67  0 t = 2
rlabel pdiffusion 157 71 158 72  0 t = 3
rlabel pdiffusion 160 71 161 72  0 t = 4
rlabel pdiffusion 156 66 162 72 0 cell no = 35
<< m1 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2 >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< m2c >>
rect 157 66 158 67 
rect 160 66 161 67 
rect 157 71 158 72 
rect 160 71 161 72 
<< labels >>
rlabel pdiffusion 193 372 194 373  0 t = 1
rlabel pdiffusion 196 372 197 373  0 t = 2
rlabel pdiffusion 193 377 194 378  0 t = 3
rlabel pdiffusion 196 377 197 378  0 t = 4
rlabel pdiffusion 192 372 198 378 0 cell no = 36
<< m1 >>
rect 193 372 194 373 
rect 196 372 197 373 
rect 193 377 194 378 
rect 196 377 197 378 
<< m2 >>
rect 193 372 194 373 
rect 196 372 197 373 
rect 193 377 194 378 
rect 196 377 197 378 
<< m2c >>
rect 193 372 194 373 
rect 196 372 197 373 
rect 193 377 194 378 
rect 196 377 197 378 
<< labels >>
rlabel pdiffusion 229 102 230 103  0 t = 1
rlabel pdiffusion 232 102 233 103  0 t = 2
rlabel pdiffusion 229 107 230 108  0 t = 3
rlabel pdiffusion 232 107 233 108  0 t = 4
rlabel pdiffusion 228 102 234 108 0 cell no = 37
<< m1 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2 >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< m2c >>
rect 229 102 230 103 
rect 232 102 233 103 
rect 229 107 230 108 
rect 232 107 233 108 
<< labels >>
rlabel pdiffusion 337 12 338 13  0 t = 1
rlabel pdiffusion 340 12 341 13  0 t = 2
rlabel pdiffusion 337 17 338 18  0 t = 3
rlabel pdiffusion 340 17 341 18  0 t = 4
rlabel pdiffusion 336 12 342 18 0 cell no = 38
<< m1 >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< m2 >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< m2c >>
rect 337 12 338 13 
rect 340 12 341 13 
rect 337 17 338 18 
rect 340 17 341 18 
<< labels >>
rlabel pdiffusion 247 120 248 121  0 t = 1
rlabel pdiffusion 250 120 251 121  0 t = 2
rlabel pdiffusion 247 125 248 126  0 t = 3
rlabel pdiffusion 250 125 251 126  0 t = 4
rlabel pdiffusion 246 120 252 126 0 cell no = 39
<< m1 >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< m2 >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< m2c >>
rect 247 120 248 121 
rect 250 120 251 121 
rect 247 125 248 126 
rect 250 125 251 126 
<< labels >>
rlabel pdiffusion 283 282 284 283  0 t = 1
rlabel pdiffusion 286 282 287 283  0 t = 2
rlabel pdiffusion 283 287 284 288  0 t = 3
rlabel pdiffusion 286 287 287 288  0 t = 4
rlabel pdiffusion 282 282 288 288 0 cell no = 40
<< m1 >>
rect 283 282 284 283 
rect 286 282 287 283 
rect 283 287 284 288 
rect 286 287 287 288 
<< m2 >>
rect 283 282 284 283 
rect 286 282 287 283 
rect 283 287 284 288 
rect 286 287 287 288 
<< m2c >>
rect 283 282 284 283 
rect 286 282 287 283 
rect 283 287 284 288 
rect 286 287 287 288 
<< labels >>
rlabel pdiffusion 13 516 14 517  0 t = 1
rlabel pdiffusion 16 516 17 517  0 t = 2
rlabel pdiffusion 13 521 14 522  0 t = 3
rlabel pdiffusion 16 521 17 522  0 t = 4
rlabel pdiffusion 12 516 18 522 0 cell no = 41
<< m1 >>
rect 13 516 14 517 
rect 16 516 17 517 
rect 13 521 14 522 
rect 16 521 17 522 
<< m2 >>
rect 13 516 14 517 
rect 16 516 17 517 
rect 13 521 14 522 
rect 16 521 17 522 
<< m2c >>
rect 13 516 14 517 
rect 16 516 17 517 
rect 13 521 14 522 
rect 16 521 17 522 
<< labels >>
rlabel pdiffusion 157 12 158 13  0 t = 1
rlabel pdiffusion 160 12 161 13  0 t = 2
rlabel pdiffusion 157 17 158 18  0 t = 3
rlabel pdiffusion 160 17 161 18  0 t = 4
rlabel pdiffusion 156 12 162 18 0 cell no = 42
<< m1 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2 >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< m2c >>
rect 157 12 158 13 
rect 160 12 161 13 
rect 157 17 158 18 
rect 160 17 161 18 
<< labels >>
rlabel pdiffusion 265 12 266 13  0 t = 1
rlabel pdiffusion 268 12 269 13  0 t = 2
rlabel pdiffusion 265 17 266 18  0 t = 3
rlabel pdiffusion 268 17 269 18  0 t = 4
rlabel pdiffusion 264 12 270 18 0 cell no = 43
<< m1 >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< m2 >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< m2c >>
rect 265 12 266 13 
rect 268 12 269 13 
rect 265 17 266 18 
rect 268 17 269 18 
<< labels >>
rlabel pdiffusion 31 498 32 499  0 t = 1
rlabel pdiffusion 34 498 35 499  0 t = 2
rlabel pdiffusion 31 503 32 504  0 t = 3
rlabel pdiffusion 34 503 35 504  0 t = 4
rlabel pdiffusion 30 498 36 504 0 cell no = 44
<< m1 >>
rect 31 498 32 499 
rect 34 498 35 499 
rect 31 503 32 504 
rect 34 503 35 504 
<< m2 >>
rect 31 498 32 499 
rect 34 498 35 499 
rect 31 503 32 504 
rect 34 503 35 504 
<< m2c >>
rect 31 498 32 499 
rect 34 498 35 499 
rect 31 503 32 504 
rect 34 503 35 504 
<< labels >>
rlabel pdiffusion 211 12 212 13  0 t = 1
rlabel pdiffusion 214 12 215 13  0 t = 2
rlabel pdiffusion 211 17 212 18  0 t = 3
rlabel pdiffusion 214 17 215 18  0 t = 4
rlabel pdiffusion 210 12 216 18 0 cell no = 45
<< m1 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2 >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< m2c >>
rect 211 12 212 13 
rect 214 12 215 13 
rect 211 17 212 18 
rect 214 17 215 18 
<< labels >>
rlabel pdiffusion 121 480 122 481  0 t = 1
rlabel pdiffusion 124 480 125 481  0 t = 2
rlabel pdiffusion 121 485 122 486  0 t = 3
rlabel pdiffusion 124 485 125 486  0 t = 4
rlabel pdiffusion 120 480 126 486 0 cell no = 46
<< m1 >>
rect 121 480 122 481 
rect 124 480 125 481 
rect 121 485 122 486 
rect 124 485 125 486 
<< m2 >>
rect 121 480 122 481 
rect 124 480 125 481 
rect 121 485 122 486 
rect 124 485 125 486 
<< m2c >>
rect 121 480 122 481 
rect 124 480 125 481 
rect 121 485 122 486 
rect 124 485 125 486 
<< labels >>
rlabel pdiffusion 175 30 176 31  0 t = 1
rlabel pdiffusion 178 30 179 31  0 t = 2
rlabel pdiffusion 175 35 176 36  0 t = 3
rlabel pdiffusion 178 35 179 36  0 t = 4
rlabel pdiffusion 174 30 180 36 0 cell no = 47
<< m1 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2 >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< m2c >>
rect 175 30 176 31 
rect 178 30 179 31 
rect 175 35 176 36 
rect 178 35 179 36 
<< labels >>
rlabel pdiffusion 283 48 284 49  0 t = 1
rlabel pdiffusion 286 48 287 49  0 t = 2
rlabel pdiffusion 283 53 284 54  0 t = 3
rlabel pdiffusion 286 53 287 54  0 t = 4
rlabel pdiffusion 282 48 288 54 0 cell no = 48
<< m1 >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< m2 >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< m2c >>
rect 283 48 284 49 
rect 286 48 287 49 
rect 283 53 284 54 
rect 286 53 287 54 
<< labels >>
rlabel pdiffusion 409 84 410 85  0 t = 1
rlabel pdiffusion 412 84 413 85  0 t = 2
rlabel pdiffusion 409 89 410 90  0 t = 3
rlabel pdiffusion 412 89 413 90  0 t = 4
rlabel pdiffusion 408 84 414 90 0 cell no = 49
<< m1 >>
rect 409 84 410 85 
rect 412 84 413 85 
rect 409 89 410 90 
rect 412 89 413 90 
<< m2 >>
rect 409 84 410 85 
rect 412 84 413 85 
rect 409 89 410 90 
rect 412 89 413 90 
<< m2c >>
rect 409 84 410 85 
rect 412 84 413 85 
rect 409 89 410 90 
rect 412 89 413 90 
<< labels >>
rlabel pdiffusion 211 228 212 229  0 t = 1
rlabel pdiffusion 214 228 215 229  0 t = 2
rlabel pdiffusion 211 233 212 234  0 t = 3
rlabel pdiffusion 214 233 215 234  0 t = 4
rlabel pdiffusion 210 228 216 234 0 cell no = 50
<< m1 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2 >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< m2c >>
rect 211 228 212 229 
rect 214 228 215 229 
rect 211 233 212 234 
rect 214 233 215 234 
<< labels >>
rlabel pdiffusion 229 12 230 13  0 t = 1
rlabel pdiffusion 232 12 233 13  0 t = 2
rlabel pdiffusion 229 17 230 18  0 t = 3
rlabel pdiffusion 232 17 233 18  0 t = 4
rlabel pdiffusion 228 12 234 18 0 cell no = 51
<< m1 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2 >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< m2c >>
rect 229 12 230 13 
rect 232 12 233 13 
rect 229 17 230 18 
rect 232 17 233 18 
<< labels >>
rlabel pdiffusion 283 12 284 13  0 t = 1
rlabel pdiffusion 286 12 287 13  0 t = 2
rlabel pdiffusion 283 17 284 18  0 t = 3
rlabel pdiffusion 286 17 287 18  0 t = 4
rlabel pdiffusion 282 12 288 18 0 cell no = 52
<< m1 >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< m2 >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< m2c >>
rect 283 12 284 13 
rect 286 12 287 13 
rect 283 17 284 18 
rect 286 17 287 18 
<< labels >>
rlabel pdiffusion 319 300 320 301  0 t = 1
rlabel pdiffusion 322 300 323 301  0 t = 2
rlabel pdiffusion 319 305 320 306  0 t = 3
rlabel pdiffusion 322 305 323 306  0 t = 4
rlabel pdiffusion 318 300 324 306 0 cell no = 53
<< m1 >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< m2 >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< m2c >>
rect 319 300 320 301 
rect 322 300 323 301 
rect 319 305 320 306 
rect 322 305 323 306 
<< labels >>
rlabel pdiffusion 481 48 482 49  0 t = 1
rlabel pdiffusion 484 48 485 49  0 t = 2
rlabel pdiffusion 481 53 482 54  0 t = 3
rlabel pdiffusion 484 53 485 54  0 t = 4
rlabel pdiffusion 480 48 486 54 0 cell no = 54
<< m1 >>
rect 481 48 482 49 
rect 484 48 485 49 
rect 481 53 482 54 
rect 484 53 485 54 
<< m2 >>
rect 481 48 482 49 
rect 484 48 485 49 
rect 481 53 482 54 
rect 484 53 485 54 
<< m2c >>
rect 481 48 482 49 
rect 484 48 485 49 
rect 481 53 482 54 
rect 484 53 485 54 
<< labels >>
rlabel pdiffusion 373 84 374 85  0 t = 1
rlabel pdiffusion 376 84 377 85  0 t = 2
rlabel pdiffusion 373 89 374 90  0 t = 3
rlabel pdiffusion 376 89 377 90  0 t = 4
rlabel pdiffusion 372 84 378 90 0 cell no = 55
<< m1 >>
rect 373 84 374 85 
rect 376 84 377 85 
rect 373 89 374 90 
rect 376 89 377 90 
<< m2 >>
rect 373 84 374 85 
rect 376 84 377 85 
rect 373 89 374 90 
rect 376 89 377 90 
<< m2c >>
rect 373 84 374 85 
rect 376 84 377 85 
rect 373 89 374 90 
rect 376 89 377 90 
<< labels >>
rlabel pdiffusion 445 336 446 337  0 t = 1
rlabel pdiffusion 448 336 449 337  0 t = 2
rlabel pdiffusion 445 341 446 342  0 t = 3
rlabel pdiffusion 448 341 449 342  0 t = 4
rlabel pdiffusion 444 336 450 342 0 cell no = 56
<< m1 >>
rect 445 336 446 337 
rect 448 336 449 337 
rect 445 341 446 342 
rect 448 341 449 342 
<< m2 >>
rect 445 336 446 337 
rect 448 336 449 337 
rect 445 341 446 342 
rect 448 341 449 342 
<< m2c >>
rect 445 336 446 337 
rect 448 336 449 337 
rect 445 341 446 342 
rect 448 341 449 342 
<< labels >>
rlabel pdiffusion 445 120 446 121  0 t = 1
rlabel pdiffusion 448 120 449 121  0 t = 2
rlabel pdiffusion 445 125 446 126  0 t = 3
rlabel pdiffusion 448 125 449 126  0 t = 4
rlabel pdiffusion 444 120 450 126 0 cell no = 57
<< m1 >>
rect 445 120 446 121 
rect 448 120 449 121 
rect 445 125 446 126 
rect 448 125 449 126 
<< m2 >>
rect 445 120 446 121 
rect 448 120 449 121 
rect 445 125 446 126 
rect 448 125 449 126 
<< m2c >>
rect 445 120 446 121 
rect 448 120 449 121 
rect 445 125 446 126 
rect 448 125 449 126 
<< labels >>
rlabel pdiffusion 265 372 266 373  0 t = 1
rlabel pdiffusion 268 372 269 373  0 t = 2
rlabel pdiffusion 265 377 266 378  0 t = 3
rlabel pdiffusion 268 377 269 378  0 t = 4
rlabel pdiffusion 264 372 270 378 0 cell no = 58
<< m1 >>
rect 265 372 266 373 
rect 268 372 269 373 
rect 265 377 266 378 
rect 268 377 269 378 
<< m2 >>
rect 265 372 266 373 
rect 268 372 269 373 
rect 265 377 266 378 
rect 268 377 269 378 
<< m2c >>
rect 265 372 266 373 
rect 268 372 269 373 
rect 265 377 266 378 
rect 268 377 269 378 
<< labels >>
rlabel pdiffusion 67 318 68 319  0 t = 1
rlabel pdiffusion 70 318 71 319  0 t = 2
rlabel pdiffusion 67 323 68 324  0 t = 3
rlabel pdiffusion 70 323 71 324  0 t = 4
rlabel pdiffusion 66 318 72 324 0 cell no = 59
<< m1 >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< m2 >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< m2c >>
rect 67 318 68 319 
rect 70 318 71 319 
rect 67 323 68 324 
rect 70 323 71 324 
<< labels >>
rlabel pdiffusion 517 48 518 49  0 t = 1
rlabel pdiffusion 520 48 521 49  0 t = 2
rlabel pdiffusion 517 53 518 54  0 t = 3
rlabel pdiffusion 520 53 521 54  0 t = 4
rlabel pdiffusion 516 48 522 54 0 cell no = 60
<< m1 >>
rect 517 48 518 49 
rect 520 48 521 49 
rect 517 53 518 54 
rect 520 53 521 54 
<< m2 >>
rect 517 48 518 49 
rect 520 48 521 49 
rect 517 53 518 54 
rect 520 53 521 54 
<< m2c >>
rect 517 48 518 49 
rect 520 48 521 49 
rect 517 53 518 54 
rect 520 53 521 54 
<< labels >>
rlabel pdiffusion 517 480 518 481  0 t = 1
rlabel pdiffusion 520 480 521 481  0 t = 2
rlabel pdiffusion 517 485 518 486  0 t = 3
rlabel pdiffusion 520 485 521 486  0 t = 4
rlabel pdiffusion 516 480 522 486 0 cell no = 61
<< m1 >>
rect 517 480 518 481 
rect 520 480 521 481 
rect 517 485 518 486 
rect 520 485 521 486 
<< m2 >>
rect 517 480 518 481 
rect 520 480 521 481 
rect 517 485 518 486 
rect 520 485 521 486 
<< m2c >>
rect 517 480 518 481 
rect 520 480 521 481 
rect 517 485 518 486 
rect 520 485 521 486 
<< labels >>
rlabel pdiffusion 139 210 140 211  0 t = 1
rlabel pdiffusion 142 210 143 211  0 t = 2
rlabel pdiffusion 139 215 140 216  0 t = 3
rlabel pdiffusion 142 215 143 216  0 t = 4
rlabel pdiffusion 138 210 144 216 0 cell no = 62
<< m1 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2 >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< m2c >>
rect 139 210 140 211 
rect 142 210 143 211 
rect 139 215 140 216 
rect 142 215 143 216 
<< labels >>
rlabel pdiffusion 373 120 374 121  0 t = 1
rlabel pdiffusion 376 120 377 121  0 t = 2
rlabel pdiffusion 373 125 374 126  0 t = 3
rlabel pdiffusion 376 125 377 126  0 t = 4
rlabel pdiffusion 372 120 378 126 0 cell no = 63
<< m1 >>
rect 373 120 374 121 
rect 376 120 377 121 
rect 373 125 374 126 
rect 376 125 377 126 
<< m2 >>
rect 373 120 374 121 
rect 376 120 377 121 
rect 373 125 374 126 
rect 376 125 377 126 
<< m2c >>
rect 373 120 374 121 
rect 376 120 377 121 
rect 373 125 374 126 
rect 376 125 377 126 
<< labels >>
rlabel pdiffusion 265 192 266 193  0 t = 1
rlabel pdiffusion 268 192 269 193  0 t = 2
rlabel pdiffusion 265 197 266 198  0 t = 3
rlabel pdiffusion 268 197 269 198  0 t = 4
rlabel pdiffusion 264 192 270 198 0 cell no = 64
<< m1 >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< m2 >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< m2c >>
rect 265 192 266 193 
rect 268 192 269 193 
rect 265 197 266 198 
rect 268 197 269 198 
<< labels >>
rlabel pdiffusion 121 48 122 49  0 t = 1
rlabel pdiffusion 124 48 125 49  0 t = 2
rlabel pdiffusion 121 53 122 54  0 t = 3
rlabel pdiffusion 124 53 125 54  0 t = 4
rlabel pdiffusion 120 48 126 54 0 cell no = 65
<< m1 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2 >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< m2c >>
rect 121 48 122 49 
rect 124 48 125 49 
rect 121 53 122 54 
rect 124 53 125 54 
<< labels >>
rlabel pdiffusion 121 228 122 229  0 t = 1
rlabel pdiffusion 124 228 125 229  0 t = 2
rlabel pdiffusion 121 233 122 234  0 t = 3
rlabel pdiffusion 124 233 125 234  0 t = 4
rlabel pdiffusion 120 228 126 234 0 cell no = 66
<< m1 >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< m2 >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< m2c >>
rect 121 228 122 229 
rect 124 228 125 229 
rect 121 233 122 234 
rect 124 233 125 234 
<< labels >>
rlabel pdiffusion 211 318 212 319  0 t = 1
rlabel pdiffusion 214 318 215 319  0 t = 2
rlabel pdiffusion 211 323 212 324  0 t = 3
rlabel pdiffusion 214 323 215 324  0 t = 4
rlabel pdiffusion 210 318 216 324 0 cell no = 67
<< m1 >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< m2 >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< m2c >>
rect 211 318 212 319 
rect 214 318 215 319 
rect 211 323 212 324 
rect 214 323 215 324 
<< labels >>
rlabel pdiffusion 211 48 212 49  0 t = 1
rlabel pdiffusion 214 48 215 49  0 t = 2
rlabel pdiffusion 211 53 212 54  0 t = 3
rlabel pdiffusion 214 53 215 54  0 t = 4
rlabel pdiffusion 210 48 216 54 0 cell no = 68
<< m1 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2 >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< m2c >>
rect 211 48 212 49 
rect 214 48 215 49 
rect 211 53 212 54 
rect 214 53 215 54 
<< labels >>
rlabel pdiffusion 103 84 104 85  0 t = 1
rlabel pdiffusion 106 84 107 85  0 t = 2
rlabel pdiffusion 103 89 104 90  0 t = 3
rlabel pdiffusion 106 89 107 90  0 t = 4
rlabel pdiffusion 102 84 108 90 0 cell no = 69
<< m1 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2 >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< m2c >>
rect 103 84 104 85 
rect 106 84 107 85 
rect 103 89 104 90 
rect 106 89 107 90 
<< labels >>
rlabel pdiffusion 85 66 86 67  0 t = 1
rlabel pdiffusion 88 66 89 67  0 t = 2
rlabel pdiffusion 85 71 86 72  0 t = 3
rlabel pdiffusion 88 71 89 72  0 t = 4
rlabel pdiffusion 84 66 90 72 0 cell no = 70
<< m1 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2 >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< m2c >>
rect 85 66 86 67 
rect 88 66 89 67 
rect 85 71 86 72 
rect 88 71 89 72 
<< labels >>
rlabel pdiffusion 427 138 428 139  0 t = 1
rlabel pdiffusion 430 138 431 139  0 t = 2
rlabel pdiffusion 427 143 428 144  0 t = 3
rlabel pdiffusion 430 143 431 144  0 t = 4
rlabel pdiffusion 426 138 432 144 0 cell no = 71
<< m1 >>
rect 427 138 428 139 
rect 430 138 431 139 
rect 427 143 428 144 
rect 430 143 431 144 
<< m2 >>
rect 427 138 428 139 
rect 430 138 431 139 
rect 427 143 428 144 
rect 430 143 431 144 
<< m2c >>
rect 427 138 428 139 
rect 430 138 431 139 
rect 427 143 428 144 
rect 430 143 431 144 
<< labels >>
rlabel pdiffusion 337 174 338 175  0 t = 1
rlabel pdiffusion 340 174 341 175  0 t = 2
rlabel pdiffusion 337 179 338 180  0 t = 3
rlabel pdiffusion 340 179 341 180  0 t = 4
rlabel pdiffusion 336 174 342 180 0 cell no = 72
<< m1 >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< m2 >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< m2c >>
rect 337 174 338 175 
rect 340 174 341 175 
rect 337 179 338 180 
rect 340 179 341 180 
<< labels >>
rlabel pdiffusion 355 30 356 31  0 t = 1
rlabel pdiffusion 358 30 359 31  0 t = 2
rlabel pdiffusion 355 35 356 36  0 t = 3
rlabel pdiffusion 358 35 359 36  0 t = 4
rlabel pdiffusion 354 30 360 36 0 cell no = 73
<< m1 >>
rect 355 30 356 31 
rect 358 30 359 31 
rect 355 35 356 36 
rect 358 35 359 36 
<< m2 >>
rect 355 30 356 31 
rect 358 30 359 31 
rect 355 35 356 36 
rect 358 35 359 36 
<< m2c >>
rect 355 30 356 31 
rect 358 30 359 31 
rect 355 35 356 36 
rect 358 35 359 36 
<< labels >>
rlabel pdiffusion 355 102 356 103  0 t = 1
rlabel pdiffusion 358 102 359 103  0 t = 2
rlabel pdiffusion 355 107 356 108  0 t = 3
rlabel pdiffusion 358 107 359 108  0 t = 4
rlabel pdiffusion 354 102 360 108 0 cell no = 74
<< m1 >>
rect 355 102 356 103 
rect 358 102 359 103 
rect 355 107 356 108 
rect 358 107 359 108 
<< m2 >>
rect 355 102 356 103 
rect 358 102 359 103 
rect 355 107 356 108 
rect 358 107 359 108 
<< m2c >>
rect 355 102 356 103 
rect 358 102 359 103 
rect 355 107 356 108 
rect 358 107 359 108 
<< labels >>
rlabel pdiffusion 265 30 266 31  0 t = 1
rlabel pdiffusion 268 30 269 31  0 t = 2
rlabel pdiffusion 265 35 266 36  0 t = 3
rlabel pdiffusion 268 35 269 36  0 t = 4
rlabel pdiffusion 264 30 270 36 0 cell no = 75
<< m1 >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< m2 >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< m2c >>
rect 265 30 266 31 
rect 268 30 269 31 
rect 265 35 266 36 
rect 268 35 269 36 
<< labels >>
rlabel pdiffusion 463 174 464 175  0 t = 1
rlabel pdiffusion 466 174 467 175  0 t = 2
rlabel pdiffusion 463 179 464 180  0 t = 3
rlabel pdiffusion 466 179 467 180  0 t = 4
rlabel pdiffusion 462 174 468 180 0 cell no = 76
<< m1 >>
rect 463 174 464 175 
rect 466 174 467 175 
rect 463 179 464 180 
rect 466 179 467 180 
<< m2 >>
rect 463 174 464 175 
rect 466 174 467 175 
rect 463 179 464 180 
rect 466 179 467 180 
<< m2c >>
rect 463 174 464 175 
rect 466 174 467 175 
rect 463 179 464 180 
rect 466 179 467 180 
<< labels >>
rlabel pdiffusion 409 192 410 193  0 t = 1
rlabel pdiffusion 412 192 413 193  0 t = 2
rlabel pdiffusion 409 197 410 198  0 t = 3
rlabel pdiffusion 412 197 413 198  0 t = 4
rlabel pdiffusion 408 192 414 198 0 cell no = 77
<< m1 >>
rect 409 192 410 193 
rect 412 192 413 193 
rect 409 197 410 198 
rect 412 197 413 198 
<< m2 >>
rect 409 192 410 193 
rect 412 192 413 193 
rect 409 197 410 198 
rect 412 197 413 198 
<< m2c >>
rect 409 192 410 193 
rect 412 192 413 193 
rect 409 197 410 198 
rect 412 197 413 198 
<< labels >>
rlabel pdiffusion 211 210 212 211  0 t = 1
rlabel pdiffusion 214 210 215 211  0 t = 2
rlabel pdiffusion 211 215 212 216  0 t = 3
rlabel pdiffusion 214 215 215 216  0 t = 4
rlabel pdiffusion 210 210 216 216 0 cell no = 78
<< m1 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2 >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< m2c >>
rect 211 210 212 211 
rect 214 210 215 211 
rect 211 215 212 216 
rect 214 215 215 216 
<< labels >>
rlabel pdiffusion 409 66 410 67  0 t = 1
rlabel pdiffusion 412 66 413 67  0 t = 2
rlabel pdiffusion 409 71 410 72  0 t = 3
rlabel pdiffusion 412 71 413 72  0 t = 4
rlabel pdiffusion 408 66 414 72 0 cell no = 79
<< m1 >>
rect 409 66 410 67 
rect 412 66 413 67 
rect 409 71 410 72 
rect 412 71 413 72 
<< m2 >>
rect 409 66 410 67 
rect 412 66 413 67 
rect 409 71 410 72 
rect 412 71 413 72 
<< m2c >>
rect 409 66 410 67 
rect 412 66 413 67 
rect 409 71 410 72 
rect 412 71 413 72 
<< labels >>
rlabel pdiffusion 229 336 230 337  0 t = 1
rlabel pdiffusion 232 336 233 337  0 t = 2
rlabel pdiffusion 229 341 230 342  0 t = 3
rlabel pdiffusion 232 341 233 342  0 t = 4
rlabel pdiffusion 228 336 234 342 0 cell no = 80
<< m1 >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< m2 >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< m2c >>
rect 229 336 230 337 
rect 232 336 233 337 
rect 229 341 230 342 
rect 232 341 233 342 
<< labels >>
rlabel pdiffusion 409 102 410 103  0 t = 1
rlabel pdiffusion 412 102 413 103  0 t = 2
rlabel pdiffusion 409 107 410 108  0 t = 3
rlabel pdiffusion 412 107 413 108  0 t = 4
rlabel pdiffusion 408 102 414 108 0 cell no = 81
<< m1 >>
rect 409 102 410 103 
rect 412 102 413 103 
rect 409 107 410 108 
rect 412 107 413 108 
<< m2 >>
rect 409 102 410 103 
rect 412 102 413 103 
rect 409 107 410 108 
rect 412 107 413 108 
<< m2c >>
rect 409 102 410 103 
rect 412 102 413 103 
rect 409 107 410 108 
rect 412 107 413 108 
<< labels >>
rlabel pdiffusion 139 120 140 121  0 t = 1
rlabel pdiffusion 142 120 143 121  0 t = 2
rlabel pdiffusion 139 125 140 126  0 t = 3
rlabel pdiffusion 142 125 143 126  0 t = 4
rlabel pdiffusion 138 120 144 126 0 cell no = 82
<< m1 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2 >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< m2c >>
rect 139 120 140 121 
rect 142 120 143 121 
rect 139 125 140 126 
rect 142 125 143 126 
<< labels >>
rlabel pdiffusion 427 156 428 157  0 t = 1
rlabel pdiffusion 430 156 431 157  0 t = 2
rlabel pdiffusion 427 161 428 162  0 t = 3
rlabel pdiffusion 430 161 431 162  0 t = 4
rlabel pdiffusion 426 156 432 162 0 cell no = 83
<< m1 >>
rect 427 156 428 157 
rect 430 156 431 157 
rect 427 161 428 162 
rect 430 161 431 162 
<< m2 >>
rect 427 156 428 157 
rect 430 156 431 157 
rect 427 161 428 162 
rect 430 161 431 162 
<< m2c >>
rect 427 156 428 157 
rect 430 156 431 157 
rect 427 161 428 162 
rect 430 161 431 162 
<< labels >>
rlabel pdiffusion 337 210 338 211  0 t = 1
rlabel pdiffusion 340 210 341 211  0 t = 2
rlabel pdiffusion 337 215 338 216  0 t = 3
rlabel pdiffusion 340 215 341 216  0 t = 4
rlabel pdiffusion 336 210 342 216 0 cell no = 84
<< m1 >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< m2 >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< m2c >>
rect 337 210 338 211 
rect 340 210 341 211 
rect 337 215 338 216 
rect 340 215 341 216 
<< labels >>
rlabel pdiffusion 283 30 284 31  0 t = 1
rlabel pdiffusion 286 30 287 31  0 t = 2
rlabel pdiffusion 283 35 284 36  0 t = 3
rlabel pdiffusion 286 35 287 36  0 t = 4
rlabel pdiffusion 282 30 288 36 0 cell no = 85
<< m1 >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< m2 >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< m2c >>
rect 283 30 284 31 
rect 286 30 287 31 
rect 283 35 284 36 
rect 286 35 287 36 
<< labels >>
rlabel pdiffusion 499 48 500 49  0 t = 1
rlabel pdiffusion 502 48 503 49  0 t = 2
rlabel pdiffusion 499 53 500 54  0 t = 3
rlabel pdiffusion 502 53 503 54  0 t = 4
rlabel pdiffusion 498 48 504 54 0 cell no = 86
<< m1 >>
rect 499 48 500 49 
rect 502 48 503 49 
rect 499 53 500 54 
rect 502 53 503 54 
<< m2 >>
rect 499 48 500 49 
rect 502 48 503 49 
rect 499 53 500 54 
rect 502 53 503 54 
<< m2c >>
rect 499 48 500 49 
rect 502 48 503 49 
rect 499 53 500 54 
rect 502 53 503 54 
<< labels >>
rlabel pdiffusion 481 282 482 283  0 t = 1
rlabel pdiffusion 484 282 485 283  0 t = 2
rlabel pdiffusion 481 287 482 288  0 t = 3
rlabel pdiffusion 484 287 485 288  0 t = 4
rlabel pdiffusion 480 282 486 288 0 cell no = 87
<< m1 >>
rect 481 282 482 283 
rect 484 282 485 283 
rect 481 287 482 288 
rect 484 287 485 288 
<< m2 >>
rect 481 282 482 283 
rect 484 282 485 283 
rect 481 287 482 288 
rect 484 287 485 288 
<< m2c >>
rect 481 282 482 283 
rect 484 282 485 283 
rect 481 287 482 288 
rect 484 287 485 288 
<< labels >>
rlabel pdiffusion 139 192 140 193  0 t = 1
rlabel pdiffusion 142 192 143 193  0 t = 2
rlabel pdiffusion 139 197 140 198  0 t = 3
rlabel pdiffusion 142 197 143 198  0 t = 4
rlabel pdiffusion 138 192 144 198 0 cell no = 88
<< m1 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2 >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< m2c >>
rect 139 192 140 193 
rect 142 192 143 193 
rect 139 197 140 198 
rect 142 197 143 198 
<< labels >>
rlabel pdiffusion 175 300 176 301  0 t = 1
rlabel pdiffusion 178 300 179 301  0 t = 2
rlabel pdiffusion 175 305 176 306  0 t = 3
rlabel pdiffusion 178 305 179 306  0 t = 4
rlabel pdiffusion 174 300 180 306 0 cell no = 89
<< m1 >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< m2 >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< m2c >>
rect 175 300 176 301 
rect 178 300 179 301 
rect 175 305 176 306 
rect 178 305 179 306 
<< labels >>
rlabel pdiffusion 139 156 140 157  0 t = 1
rlabel pdiffusion 142 156 143 157  0 t = 2
rlabel pdiffusion 139 161 140 162  0 t = 3
rlabel pdiffusion 142 161 143 162  0 t = 4
rlabel pdiffusion 138 156 144 162 0 cell no = 90
<< m1 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2 >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< m2c >>
rect 139 156 140 157 
rect 142 156 143 157 
rect 139 161 140 162 
rect 142 161 143 162 
<< labels >>
rlabel pdiffusion 67 30 68 31  0 t = 1
rlabel pdiffusion 70 30 71 31  0 t = 2
rlabel pdiffusion 67 35 68 36  0 t = 3
rlabel pdiffusion 70 35 71 36  0 t = 4
rlabel pdiffusion 66 30 72 36 0 cell no = 91
<< m1 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2 >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< m2c >>
rect 67 30 68 31 
rect 70 30 71 31 
rect 67 35 68 36 
rect 70 35 71 36 
<< labels >>
rlabel pdiffusion 31 66 32 67  0 t = 1
rlabel pdiffusion 34 66 35 67  0 t = 2
rlabel pdiffusion 31 71 32 72  0 t = 3
rlabel pdiffusion 34 71 35 72  0 t = 4
rlabel pdiffusion 30 66 36 72 0 cell no = 92
<< m1 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2 >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< m2c >>
rect 31 66 32 67 
rect 34 66 35 67 
rect 31 71 32 72 
rect 34 71 35 72 
<< labels >>
rlabel pdiffusion 31 156 32 157  0 t = 1
rlabel pdiffusion 34 156 35 157  0 t = 2
rlabel pdiffusion 31 161 32 162  0 t = 3
rlabel pdiffusion 34 161 35 162  0 t = 4
rlabel pdiffusion 30 156 36 162 0 cell no = 93
<< m1 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2 >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< m2c >>
rect 31 156 32 157 
rect 34 156 35 157 
rect 31 161 32 162 
rect 34 161 35 162 
<< labels >>
rlabel pdiffusion 157 156 158 157  0 t = 1
rlabel pdiffusion 160 156 161 157  0 t = 2
rlabel pdiffusion 157 161 158 162  0 t = 3
rlabel pdiffusion 160 161 161 162  0 t = 4
rlabel pdiffusion 156 156 162 162 0 cell no = 94
<< m1 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2 >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< m2c >>
rect 157 156 158 157 
rect 160 156 161 157 
rect 157 161 158 162 
rect 160 161 161 162 
<< labels >>
rlabel pdiffusion 49 318 50 319  0 t = 1
rlabel pdiffusion 52 318 53 319  0 t = 2
rlabel pdiffusion 49 323 50 324  0 t = 3
rlabel pdiffusion 52 323 53 324  0 t = 4
rlabel pdiffusion 48 318 54 324 0 cell no = 95
<< m1 >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< m2 >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< m2c >>
rect 49 318 50 319 
rect 52 318 53 319 
rect 49 323 50 324 
rect 52 323 53 324 
<< labels >>
rlabel pdiffusion 193 48 194 49  0 t = 1
rlabel pdiffusion 196 48 197 49  0 t = 2
rlabel pdiffusion 193 53 194 54  0 t = 3
rlabel pdiffusion 196 53 197 54  0 t = 4
rlabel pdiffusion 192 48 198 54 0 cell no = 96
<< m1 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2 >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< m2c >>
rect 193 48 194 49 
rect 196 48 197 49 
rect 193 53 194 54 
rect 196 53 197 54 
<< labels >>
rlabel pdiffusion 337 48 338 49  0 t = 1
rlabel pdiffusion 340 48 341 49  0 t = 2
rlabel pdiffusion 337 53 338 54  0 t = 3
rlabel pdiffusion 340 53 341 54  0 t = 4
rlabel pdiffusion 336 48 342 54 0 cell no = 97
<< m1 >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< m2 >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< m2c >>
rect 337 48 338 49 
rect 340 48 341 49 
rect 337 53 338 54 
rect 340 53 341 54 
<< labels >>
rlabel pdiffusion 265 426 266 427  0 t = 1
rlabel pdiffusion 268 426 269 427  0 t = 2
rlabel pdiffusion 265 431 266 432  0 t = 3
rlabel pdiffusion 268 431 269 432  0 t = 4
rlabel pdiffusion 264 426 270 432 0 cell no = 98
<< m1 >>
rect 265 426 266 427 
rect 268 426 269 427 
rect 265 431 266 432 
rect 268 431 269 432 
<< m2 >>
rect 265 426 266 427 
rect 268 426 269 427 
rect 265 431 266 432 
rect 268 431 269 432 
<< m2c >>
rect 265 426 266 427 
rect 268 426 269 427 
rect 265 431 266 432 
rect 268 431 269 432 
<< labels >>
rlabel pdiffusion 247 282 248 283  0 t = 1
rlabel pdiffusion 250 282 251 283  0 t = 2
rlabel pdiffusion 247 287 248 288  0 t = 3
rlabel pdiffusion 250 287 251 288  0 t = 4
rlabel pdiffusion 246 282 252 288 0 cell no = 99
<< m1 >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< m2 >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< m2c >>
rect 247 282 248 283 
rect 250 282 251 283 
rect 247 287 248 288 
rect 250 287 251 288 
<< labels >>
rlabel pdiffusion 121 138 122 139  0 t = 1
rlabel pdiffusion 124 138 125 139  0 t = 2
rlabel pdiffusion 121 143 122 144  0 t = 3
rlabel pdiffusion 124 143 125 144  0 t = 4
rlabel pdiffusion 120 138 126 144 0 cell no = 100
<< m1 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2 >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< m2c >>
rect 121 138 122 139 
rect 124 138 125 139 
rect 121 143 122 144 
rect 124 143 125 144 
<< labels >>
rlabel pdiffusion 211 30 212 31  0 t = 1
rlabel pdiffusion 214 30 215 31  0 t = 2
rlabel pdiffusion 211 35 212 36  0 t = 3
rlabel pdiffusion 214 35 215 36  0 t = 4
rlabel pdiffusion 210 30 216 36 0 cell no = 101
<< m1 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2 >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< m2c >>
rect 211 30 212 31 
rect 214 30 215 31 
rect 211 35 212 36 
rect 214 35 215 36 
<< labels >>
rlabel pdiffusion 265 66 266 67  0 t = 1
rlabel pdiffusion 268 66 269 67  0 t = 2
rlabel pdiffusion 265 71 266 72  0 t = 3
rlabel pdiffusion 268 71 269 72  0 t = 4
rlabel pdiffusion 264 66 270 72 0 cell no = 102
<< m1 >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< m2 >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< m2c >>
rect 265 66 266 67 
rect 268 66 269 67 
rect 265 71 266 72 
rect 268 71 269 72 
<< labels >>
rlabel pdiffusion 319 120 320 121  0 t = 1
rlabel pdiffusion 322 120 323 121  0 t = 2
rlabel pdiffusion 319 125 320 126  0 t = 3
rlabel pdiffusion 322 125 323 126  0 t = 4
rlabel pdiffusion 318 120 324 126 0 cell no = 103
<< m1 >>
rect 319 120 320 121 
rect 322 120 323 121 
rect 319 125 320 126 
rect 322 125 323 126 
<< m2 >>
rect 319 120 320 121 
rect 322 120 323 121 
rect 319 125 320 126 
rect 322 125 323 126 
<< m2c >>
rect 319 120 320 121 
rect 322 120 323 121 
rect 319 125 320 126 
rect 322 125 323 126 
<< labels >>
rlabel pdiffusion 265 48 266 49  0 t = 1
rlabel pdiffusion 268 48 269 49  0 t = 2
rlabel pdiffusion 265 53 266 54  0 t = 3
rlabel pdiffusion 268 53 269 54  0 t = 4
rlabel pdiffusion 264 48 270 54 0 cell no = 104
<< m1 >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< m2 >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< m2c >>
rect 265 48 266 49 
rect 268 48 269 49 
rect 265 53 266 54 
rect 268 53 269 54 
<< labels >>
rlabel pdiffusion 283 120 284 121  0 t = 1
rlabel pdiffusion 286 120 287 121  0 t = 2
rlabel pdiffusion 283 125 284 126  0 t = 3
rlabel pdiffusion 286 125 287 126  0 t = 4
rlabel pdiffusion 282 120 288 126 0 cell no = 105
<< m1 >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< m2 >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< m2c >>
rect 283 120 284 121 
rect 286 120 287 121 
rect 283 125 284 126 
rect 286 125 287 126 
<< labels >>
rlabel pdiffusion 247 192 248 193  0 t = 1
rlabel pdiffusion 250 192 251 193  0 t = 2
rlabel pdiffusion 247 197 248 198  0 t = 3
rlabel pdiffusion 250 197 251 198  0 t = 4
rlabel pdiffusion 246 192 252 198 0 cell no = 106
<< m1 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2 >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< m2c >>
rect 247 192 248 193 
rect 250 192 251 193 
rect 247 197 248 198 
rect 250 197 251 198 
<< labels >>
rlabel pdiffusion 481 354 482 355  0 t = 1
rlabel pdiffusion 484 354 485 355  0 t = 2
rlabel pdiffusion 481 359 482 360  0 t = 3
rlabel pdiffusion 484 359 485 360  0 t = 4
rlabel pdiffusion 480 354 486 360 0 cell no = 107
<< m1 >>
rect 481 354 482 355 
rect 484 354 485 355 
rect 481 359 482 360 
rect 484 359 485 360 
<< m2 >>
rect 481 354 482 355 
rect 484 354 485 355 
rect 481 359 482 360 
rect 484 359 485 360 
<< m2c >>
rect 481 354 482 355 
rect 484 354 485 355 
rect 481 359 482 360 
rect 484 359 485 360 
<< labels >>
rlabel pdiffusion 337 120 338 121  0 t = 1
rlabel pdiffusion 340 120 341 121  0 t = 2
rlabel pdiffusion 337 125 338 126  0 t = 3
rlabel pdiffusion 340 125 341 126  0 t = 4
rlabel pdiffusion 336 120 342 126 0 cell no = 108
<< m1 >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< m2 >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< m2c >>
rect 337 120 338 121 
rect 340 120 341 121 
rect 337 125 338 126 
rect 340 125 341 126 
<< labels >>
rlabel pdiffusion 391 48 392 49  0 t = 1
rlabel pdiffusion 394 48 395 49  0 t = 2
rlabel pdiffusion 391 53 392 54  0 t = 3
rlabel pdiffusion 394 53 395 54  0 t = 4
rlabel pdiffusion 390 48 396 54 0 cell no = 109
<< m1 >>
rect 391 48 392 49 
rect 394 48 395 49 
rect 391 53 392 54 
rect 394 53 395 54 
<< m2 >>
rect 391 48 392 49 
rect 394 48 395 49 
rect 391 53 392 54 
rect 394 53 395 54 
<< m2c >>
rect 391 48 392 49 
rect 394 48 395 49 
rect 391 53 392 54 
rect 394 53 395 54 
<< labels >>
rlabel pdiffusion 337 246 338 247  0 t = 1
rlabel pdiffusion 340 246 341 247  0 t = 2
rlabel pdiffusion 337 251 338 252  0 t = 3
rlabel pdiffusion 340 251 341 252  0 t = 4
rlabel pdiffusion 336 246 342 252 0 cell no = 110
<< m1 >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< m2 >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< m2c >>
rect 337 246 338 247 
rect 340 246 341 247 
rect 337 251 338 252 
rect 340 251 341 252 
<< labels >>
rlabel pdiffusion 391 174 392 175  0 t = 1
rlabel pdiffusion 394 174 395 175  0 t = 2
rlabel pdiffusion 391 179 392 180  0 t = 3
rlabel pdiffusion 394 179 395 180  0 t = 4
rlabel pdiffusion 390 174 396 180 0 cell no = 111
<< m1 >>
rect 391 174 392 175 
rect 394 174 395 175 
rect 391 179 392 180 
rect 394 179 395 180 
<< m2 >>
rect 391 174 392 175 
rect 394 174 395 175 
rect 391 179 392 180 
rect 394 179 395 180 
<< m2c >>
rect 391 174 392 175 
rect 394 174 395 175 
rect 391 179 392 180 
rect 394 179 395 180 
<< labels >>
rlabel pdiffusion 517 210 518 211  0 t = 1
rlabel pdiffusion 520 210 521 211  0 t = 2
rlabel pdiffusion 517 215 518 216  0 t = 3
rlabel pdiffusion 520 215 521 216  0 t = 4
rlabel pdiffusion 516 210 522 216 0 cell no = 112
<< m1 >>
rect 517 210 518 211 
rect 520 210 521 211 
rect 517 215 518 216 
rect 520 215 521 216 
<< m2 >>
rect 517 210 518 211 
rect 520 210 521 211 
rect 517 215 518 216 
rect 520 215 521 216 
<< m2c >>
rect 517 210 518 211 
rect 520 210 521 211 
rect 517 215 518 216 
rect 520 215 521 216 
<< labels >>
rlabel pdiffusion 229 48 230 49  0 t = 1
rlabel pdiffusion 232 48 233 49  0 t = 2
rlabel pdiffusion 229 53 230 54  0 t = 3
rlabel pdiffusion 232 53 233 54  0 t = 4
rlabel pdiffusion 228 48 234 54 0 cell no = 113
<< m1 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2 >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< m2c >>
rect 229 48 230 49 
rect 232 48 233 49 
rect 229 53 230 54 
rect 232 53 233 54 
<< labels >>
rlabel pdiffusion 463 120 464 121  0 t = 1
rlabel pdiffusion 466 120 467 121  0 t = 2
rlabel pdiffusion 463 125 464 126  0 t = 3
rlabel pdiffusion 466 125 467 126  0 t = 4
rlabel pdiffusion 462 120 468 126 0 cell no = 114
<< m1 >>
rect 463 120 464 121 
rect 466 120 467 121 
rect 463 125 464 126 
rect 466 125 467 126 
<< m2 >>
rect 463 120 464 121 
rect 466 120 467 121 
rect 463 125 464 126 
rect 466 125 467 126 
<< m2c >>
rect 463 120 464 121 
rect 466 120 467 121 
rect 463 125 464 126 
rect 466 125 467 126 
<< labels >>
rlabel pdiffusion 445 156 446 157  0 t = 1
rlabel pdiffusion 448 156 449 157  0 t = 2
rlabel pdiffusion 445 161 446 162  0 t = 3
rlabel pdiffusion 448 161 449 162  0 t = 4
rlabel pdiffusion 444 156 450 162 0 cell no = 115
<< m1 >>
rect 445 156 446 157 
rect 448 156 449 157 
rect 445 161 446 162 
rect 448 161 449 162 
<< m2 >>
rect 445 156 446 157 
rect 448 156 449 157 
rect 445 161 446 162 
rect 448 161 449 162 
<< m2c >>
rect 445 156 446 157 
rect 448 156 449 157 
rect 445 161 446 162 
rect 448 161 449 162 
<< labels >>
rlabel pdiffusion 13 102 14 103  0 t = 1
rlabel pdiffusion 16 102 17 103  0 t = 2
rlabel pdiffusion 13 107 14 108  0 t = 3
rlabel pdiffusion 16 107 17 108  0 t = 4
rlabel pdiffusion 12 102 18 108 0 cell no = 116
<< m1 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2 >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< m2c >>
rect 13 102 14 103 
rect 16 102 17 103 
rect 13 107 14 108 
rect 16 107 17 108 
<< labels >>
rlabel pdiffusion 229 120 230 121  0 t = 1
rlabel pdiffusion 232 120 233 121  0 t = 2
rlabel pdiffusion 229 125 230 126  0 t = 3
rlabel pdiffusion 232 125 233 126  0 t = 4
rlabel pdiffusion 228 120 234 126 0 cell no = 117
<< m1 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2 >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< m2c >>
rect 229 120 230 121 
rect 232 120 233 121 
rect 229 125 230 126 
rect 232 125 233 126 
<< labels >>
rlabel pdiffusion 67 12 68 13  0 t = 1
rlabel pdiffusion 70 12 71 13  0 t = 2
rlabel pdiffusion 67 17 68 18  0 t = 3
rlabel pdiffusion 70 17 71 18  0 t = 4
rlabel pdiffusion 66 12 72 18 0 cell no = 118
<< m1 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2 >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< m2c >>
rect 67 12 68 13 
rect 70 12 71 13 
rect 67 17 68 18 
rect 70 17 71 18 
<< labels >>
rlabel pdiffusion 13 66 14 67  0 t = 1
rlabel pdiffusion 16 66 17 67  0 t = 2
rlabel pdiffusion 13 71 14 72  0 t = 3
rlabel pdiffusion 16 71 17 72  0 t = 4
rlabel pdiffusion 12 66 18 72 0 cell no = 119
<< m1 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2 >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< m2c >>
rect 13 66 14 67 
rect 16 66 17 67 
rect 13 71 14 72 
rect 16 71 17 72 
<< labels >>
rlabel pdiffusion 121 66 122 67  0 t = 1
rlabel pdiffusion 124 66 125 67  0 t = 2
rlabel pdiffusion 121 71 122 72  0 t = 3
rlabel pdiffusion 124 71 125 72  0 t = 4
rlabel pdiffusion 120 66 126 72 0 cell no = 120
<< m1 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2 >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< m2c >>
rect 121 66 122 67 
rect 124 66 125 67 
rect 121 71 122 72 
rect 124 71 125 72 
<< labels >>
rlabel pdiffusion 103 48 104 49  0 t = 1
rlabel pdiffusion 106 48 107 49  0 t = 2
rlabel pdiffusion 103 53 104 54  0 t = 3
rlabel pdiffusion 106 53 107 54  0 t = 4
rlabel pdiffusion 102 48 108 54 0 cell no = 121
<< m1 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2 >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< m2c >>
rect 103 48 104 49 
rect 106 48 107 49 
rect 103 53 104 54 
rect 106 53 107 54 
<< labels >>
rlabel pdiffusion 193 390 194 391  0 t = 1
rlabel pdiffusion 196 390 197 391  0 t = 2
rlabel pdiffusion 193 395 194 396  0 t = 3
rlabel pdiffusion 196 395 197 396  0 t = 4
rlabel pdiffusion 192 390 198 396 0 cell no = 122
<< m1 >>
rect 193 390 194 391 
rect 196 390 197 391 
rect 193 395 194 396 
rect 196 395 197 396 
<< m2 >>
rect 193 390 194 391 
rect 196 390 197 391 
rect 193 395 194 396 
rect 196 395 197 396 
<< m2c >>
rect 193 390 194 391 
rect 196 390 197 391 
rect 193 395 194 396 
rect 196 395 197 396 
<< labels >>
rlabel pdiffusion 13 48 14 49  0 t = 1
rlabel pdiffusion 16 48 17 49  0 t = 2
rlabel pdiffusion 13 53 14 54  0 t = 3
rlabel pdiffusion 16 53 17 54  0 t = 4
rlabel pdiffusion 12 48 18 54 0 cell no = 123
<< m1 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2 >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< m2c >>
rect 13 48 14 49 
rect 16 48 17 49 
rect 13 53 14 54 
rect 16 53 17 54 
<< labels >>
rlabel pdiffusion 193 84 194 85  0 t = 1
rlabel pdiffusion 196 84 197 85  0 t = 2
rlabel pdiffusion 193 89 194 90  0 t = 3
rlabel pdiffusion 196 89 197 90  0 t = 4
rlabel pdiffusion 192 84 198 90 0 cell no = 124
<< m1 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2 >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< m2c >>
rect 193 84 194 85 
rect 196 84 197 85 
rect 193 89 194 90 
rect 196 89 197 90 
<< labels >>
rlabel pdiffusion 301 48 302 49  0 t = 1
rlabel pdiffusion 304 48 305 49  0 t = 2
rlabel pdiffusion 301 53 302 54  0 t = 3
rlabel pdiffusion 304 53 305 54  0 t = 4
rlabel pdiffusion 300 48 306 54 0 cell no = 125
<< m1 >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< m2 >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< m2c >>
rect 301 48 302 49 
rect 304 48 305 49 
rect 301 53 302 54 
rect 304 53 305 54 
<< labels >>
rlabel pdiffusion 175 84 176 85  0 t = 1
rlabel pdiffusion 178 84 179 85  0 t = 2
rlabel pdiffusion 175 89 176 90  0 t = 3
rlabel pdiffusion 178 89 179 90  0 t = 4
rlabel pdiffusion 174 84 180 90 0 cell no = 126
<< m1 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2 >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< m2c >>
rect 175 84 176 85 
rect 178 84 179 85 
rect 175 89 176 90 
rect 178 89 179 90 
<< labels >>
rlabel pdiffusion 247 66 248 67  0 t = 1
rlabel pdiffusion 250 66 251 67  0 t = 2
rlabel pdiffusion 247 71 248 72  0 t = 3
rlabel pdiffusion 250 71 251 72  0 t = 4
rlabel pdiffusion 246 66 252 72 0 cell no = 127
<< m1 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2 >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< m2c >>
rect 247 66 248 67 
rect 250 66 251 67 
rect 247 71 248 72 
rect 250 71 251 72 
<< labels >>
rlabel pdiffusion 301 138 302 139  0 t = 1
rlabel pdiffusion 304 138 305 139  0 t = 2
rlabel pdiffusion 301 143 302 144  0 t = 3
rlabel pdiffusion 304 143 305 144  0 t = 4
rlabel pdiffusion 300 138 306 144 0 cell no = 128
<< m1 >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< m2 >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< m2c >>
rect 301 138 302 139 
rect 304 138 305 139 
rect 301 143 302 144 
rect 304 143 305 144 
<< labels >>
rlabel pdiffusion 85 30 86 31  0 t = 1
rlabel pdiffusion 88 30 89 31  0 t = 2
rlabel pdiffusion 85 35 86 36  0 t = 3
rlabel pdiffusion 88 35 89 36  0 t = 4
rlabel pdiffusion 84 30 90 36 0 cell no = 129
<< m1 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2 >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< m2c >>
rect 85 30 86 31 
rect 88 30 89 31 
rect 85 35 86 36 
rect 88 35 89 36 
<< labels >>
rlabel pdiffusion 193 120 194 121  0 t = 1
rlabel pdiffusion 196 120 197 121  0 t = 2
rlabel pdiffusion 193 125 194 126  0 t = 3
rlabel pdiffusion 196 125 197 126  0 t = 4
rlabel pdiffusion 192 120 198 126 0 cell no = 130
<< m1 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2 >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< m2c >>
rect 193 120 194 121 
rect 196 120 197 121 
rect 193 125 194 126 
rect 196 125 197 126 
<< labels >>
rlabel pdiffusion 301 120 302 121  0 t = 1
rlabel pdiffusion 304 120 305 121  0 t = 2
rlabel pdiffusion 301 125 302 126  0 t = 3
rlabel pdiffusion 304 125 305 126  0 t = 4
rlabel pdiffusion 300 120 306 126 0 cell no = 131
<< m1 >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< m2 >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< m2c >>
rect 301 120 302 121 
rect 304 120 305 121 
rect 301 125 302 126 
rect 304 125 305 126 
<< labels >>
rlabel pdiffusion 175 66 176 67  0 t = 1
rlabel pdiffusion 178 66 179 67  0 t = 2
rlabel pdiffusion 175 71 176 72  0 t = 3
rlabel pdiffusion 178 71 179 72  0 t = 4
rlabel pdiffusion 174 66 180 72 0 cell no = 132
<< m1 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2 >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< m2c >>
rect 175 66 176 67 
rect 178 66 179 67 
rect 175 71 176 72 
rect 178 71 179 72 
<< labels >>
rlabel pdiffusion 193 318 194 319  0 t = 1
rlabel pdiffusion 196 318 197 319  0 t = 2
rlabel pdiffusion 193 323 194 324  0 t = 3
rlabel pdiffusion 196 323 197 324  0 t = 4
rlabel pdiffusion 192 318 198 324 0 cell no = 133
<< m1 >>
rect 193 318 194 319 
rect 196 318 197 319 
rect 193 323 194 324 
rect 196 323 197 324 
<< m2 >>
rect 193 318 194 319 
rect 196 318 197 319 
rect 193 323 194 324 
rect 196 323 197 324 
<< m2c >>
rect 193 318 194 319 
rect 196 318 197 319 
rect 193 323 194 324 
rect 196 323 197 324 
<< labels >>
rlabel pdiffusion 301 12 302 13  0 t = 1
rlabel pdiffusion 304 12 305 13  0 t = 2
rlabel pdiffusion 301 17 302 18  0 t = 3
rlabel pdiffusion 304 17 305 18  0 t = 4
rlabel pdiffusion 300 12 306 18 0 cell no = 134
<< m1 >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< m2 >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< m2c >>
rect 301 12 302 13 
rect 304 12 305 13 
rect 301 17 302 18 
rect 304 17 305 18 
<< labels >>
rlabel pdiffusion 499 138 500 139  0 t = 1
rlabel pdiffusion 502 138 503 139  0 t = 2
rlabel pdiffusion 499 143 500 144  0 t = 3
rlabel pdiffusion 502 143 503 144  0 t = 4
rlabel pdiffusion 498 138 504 144 0 cell no = 135
<< m1 >>
rect 499 138 500 139 
rect 502 138 503 139 
rect 499 143 500 144 
rect 502 143 503 144 
<< m2 >>
rect 499 138 500 139 
rect 502 138 503 139 
rect 499 143 500 144 
rect 502 143 503 144 
<< m2c >>
rect 499 138 500 139 
rect 502 138 503 139 
rect 499 143 500 144 
rect 502 143 503 144 
<< labels >>
rlabel pdiffusion 517 156 518 157  0 t = 1
rlabel pdiffusion 520 156 521 157  0 t = 2
rlabel pdiffusion 517 161 518 162  0 t = 3
rlabel pdiffusion 520 161 521 162  0 t = 4
rlabel pdiffusion 516 156 522 162 0 cell no = 136
<< m1 >>
rect 517 156 518 157 
rect 520 156 521 157 
rect 517 161 518 162 
rect 520 161 521 162 
<< m2 >>
rect 517 156 518 157 
rect 520 156 521 157 
rect 517 161 518 162 
rect 520 161 521 162 
<< m2c >>
rect 517 156 518 157 
rect 520 156 521 157 
rect 517 161 518 162 
rect 520 161 521 162 
<< labels >>
rlabel pdiffusion 175 480 176 481  0 t = 1
rlabel pdiffusion 178 480 179 481  0 t = 2
rlabel pdiffusion 175 485 176 486  0 t = 3
rlabel pdiffusion 178 485 179 486  0 t = 4
rlabel pdiffusion 174 480 180 486 0 cell no = 137
<< m1 >>
rect 175 480 176 481 
rect 178 480 179 481 
rect 175 485 176 486 
rect 178 485 179 486 
<< m2 >>
rect 175 480 176 481 
rect 178 480 179 481 
rect 175 485 176 486 
rect 178 485 179 486 
<< m2c >>
rect 175 480 176 481 
rect 178 480 179 481 
rect 175 485 176 486 
rect 178 485 179 486 
<< labels >>
rlabel pdiffusion 373 210 374 211  0 t = 1
rlabel pdiffusion 376 210 377 211  0 t = 2
rlabel pdiffusion 373 215 374 216  0 t = 3
rlabel pdiffusion 376 215 377 216  0 t = 4
rlabel pdiffusion 372 210 378 216 0 cell no = 138
<< m1 >>
rect 373 210 374 211 
rect 376 210 377 211 
rect 373 215 374 216 
rect 376 215 377 216 
<< m2 >>
rect 373 210 374 211 
rect 376 210 377 211 
rect 373 215 374 216 
rect 376 215 377 216 
<< m2c >>
rect 373 210 374 211 
rect 376 210 377 211 
rect 373 215 374 216 
rect 376 215 377 216 
<< labels >>
rlabel pdiffusion 247 174 248 175  0 t = 1
rlabel pdiffusion 250 174 251 175  0 t = 2
rlabel pdiffusion 247 179 248 180  0 t = 3
rlabel pdiffusion 250 179 251 180  0 t = 4
rlabel pdiffusion 246 174 252 180 0 cell no = 139
<< m1 >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< m2 >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< m2c >>
rect 247 174 248 175 
rect 250 174 251 175 
rect 247 179 248 180 
rect 250 179 251 180 
<< labels >>
rlabel pdiffusion 49 48 50 49  0 t = 1
rlabel pdiffusion 52 48 53 49  0 t = 2
rlabel pdiffusion 49 53 50 54  0 t = 3
rlabel pdiffusion 52 53 53 54  0 t = 4
rlabel pdiffusion 48 48 54 54 0 cell no = 140
<< m1 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2 >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< m2c >>
rect 49 48 50 49 
rect 52 48 53 49 
rect 49 53 50 54 
rect 52 53 53 54 
<< labels >>
rlabel pdiffusion 481 66 482 67  0 t = 1
rlabel pdiffusion 484 66 485 67  0 t = 2
rlabel pdiffusion 481 71 482 72  0 t = 3
rlabel pdiffusion 484 71 485 72  0 t = 4
rlabel pdiffusion 480 66 486 72 0 cell no = 141
<< m1 >>
rect 481 66 482 67 
rect 484 66 485 67 
rect 481 71 482 72 
rect 484 71 485 72 
<< m2 >>
rect 481 66 482 67 
rect 484 66 485 67 
rect 481 71 482 72 
rect 484 71 485 72 
<< m2c >>
rect 481 66 482 67 
rect 484 66 485 67 
rect 481 71 482 72 
rect 484 71 485 72 
<< labels >>
rlabel pdiffusion 13 354 14 355  0 t = 1
rlabel pdiffusion 16 354 17 355  0 t = 2
rlabel pdiffusion 13 359 14 360  0 t = 3
rlabel pdiffusion 16 359 17 360  0 t = 4
rlabel pdiffusion 12 354 18 360 0 cell no = 142
<< m1 >>
rect 13 354 14 355 
rect 16 354 17 355 
rect 13 359 14 360 
rect 16 359 17 360 
<< m2 >>
rect 13 354 14 355 
rect 16 354 17 355 
rect 13 359 14 360 
rect 16 359 17 360 
<< m2c >>
rect 13 354 14 355 
rect 16 354 17 355 
rect 13 359 14 360 
rect 16 359 17 360 
<< labels >>
rlabel pdiffusion 229 264 230 265  0 t = 1
rlabel pdiffusion 232 264 233 265  0 t = 2
rlabel pdiffusion 229 269 230 270  0 t = 3
rlabel pdiffusion 232 269 233 270  0 t = 4
rlabel pdiffusion 228 264 234 270 0 cell no = 143
<< m1 >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< m2 >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< m2c >>
rect 229 264 230 265 
rect 232 264 233 265 
rect 229 269 230 270 
rect 232 269 233 270 
<< labels >>
rlabel pdiffusion 337 66 338 67  0 t = 1
rlabel pdiffusion 340 66 341 67  0 t = 2
rlabel pdiffusion 337 71 338 72  0 t = 3
rlabel pdiffusion 340 71 341 72  0 t = 4
rlabel pdiffusion 336 66 342 72 0 cell no = 144
<< m1 >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< m2 >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< m2c >>
rect 337 66 338 67 
rect 340 66 341 67 
rect 337 71 338 72 
rect 340 71 341 72 
<< labels >>
rlabel pdiffusion 121 408 122 409  0 t = 1
rlabel pdiffusion 124 408 125 409  0 t = 2
rlabel pdiffusion 121 413 122 414  0 t = 3
rlabel pdiffusion 124 413 125 414  0 t = 4
rlabel pdiffusion 120 408 126 414 0 cell no = 145
<< m1 >>
rect 121 408 122 409 
rect 124 408 125 409 
rect 121 413 122 414 
rect 124 413 125 414 
<< m2 >>
rect 121 408 122 409 
rect 124 408 125 409 
rect 121 413 122 414 
rect 124 413 125 414 
<< m2c >>
rect 121 408 122 409 
rect 124 408 125 409 
rect 121 413 122 414 
rect 124 413 125 414 
<< labels >>
rlabel pdiffusion 247 300 248 301  0 t = 1
rlabel pdiffusion 250 300 251 301  0 t = 2
rlabel pdiffusion 247 305 248 306  0 t = 3
rlabel pdiffusion 250 305 251 306  0 t = 4
rlabel pdiffusion 246 300 252 306 0 cell no = 146
<< m1 >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< m2 >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< m2c >>
rect 247 300 248 301 
rect 250 300 251 301 
rect 247 305 248 306 
rect 250 305 251 306 
<< labels >>
rlabel pdiffusion 283 480 284 481  0 t = 1
rlabel pdiffusion 286 480 287 481  0 t = 2
rlabel pdiffusion 283 485 284 486  0 t = 3
rlabel pdiffusion 286 485 287 486  0 t = 4
rlabel pdiffusion 282 480 288 486 0 cell no = 147
<< m1 >>
rect 283 480 284 481 
rect 286 480 287 481 
rect 283 485 284 486 
rect 286 485 287 486 
<< m2 >>
rect 283 480 284 481 
rect 286 480 287 481 
rect 283 485 284 486 
rect 286 485 287 486 
<< m2c >>
rect 283 480 284 481 
rect 286 480 287 481 
rect 283 485 284 486 
rect 286 485 287 486 
<< labels >>
rlabel pdiffusion 31 102 32 103  0 t = 1
rlabel pdiffusion 34 102 35 103  0 t = 2
rlabel pdiffusion 31 107 32 108  0 t = 3
rlabel pdiffusion 34 107 35 108  0 t = 4
rlabel pdiffusion 30 102 36 108 0 cell no = 148
<< m1 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2 >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< m2c >>
rect 31 102 32 103 
rect 34 102 35 103 
rect 31 107 32 108 
rect 34 107 35 108 
<< labels >>
rlabel pdiffusion 175 336 176 337  0 t = 1
rlabel pdiffusion 178 336 179 337  0 t = 2
rlabel pdiffusion 175 341 176 342  0 t = 3
rlabel pdiffusion 178 341 179 342  0 t = 4
rlabel pdiffusion 174 336 180 342 0 cell no = 149
<< m1 >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< m2 >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< m2c >>
rect 175 336 176 337 
rect 178 336 179 337 
rect 175 341 176 342 
rect 178 341 179 342 
<< labels >>
rlabel pdiffusion 85 192 86 193  0 t = 1
rlabel pdiffusion 88 192 89 193  0 t = 2
rlabel pdiffusion 85 197 86 198  0 t = 3
rlabel pdiffusion 88 197 89 198  0 t = 4
rlabel pdiffusion 84 192 90 198 0 cell no = 150
<< m1 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2 >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< m2c >>
rect 85 192 86 193 
rect 88 192 89 193 
rect 85 197 86 198 
rect 88 197 89 198 
<< labels >>
rlabel pdiffusion 229 156 230 157  0 t = 1
rlabel pdiffusion 232 156 233 157  0 t = 2
rlabel pdiffusion 229 161 230 162  0 t = 3
rlabel pdiffusion 232 161 233 162  0 t = 4
rlabel pdiffusion 228 156 234 162 0 cell no = 151
<< m1 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2 >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< m2c >>
rect 229 156 230 157 
rect 232 156 233 157 
rect 229 161 230 162 
rect 232 161 233 162 
<< labels >>
rlabel pdiffusion 391 228 392 229  0 t = 1
rlabel pdiffusion 394 228 395 229  0 t = 2
rlabel pdiffusion 391 233 392 234  0 t = 3
rlabel pdiffusion 394 233 395 234  0 t = 4
rlabel pdiffusion 390 228 396 234 0 cell no = 152
<< m1 >>
rect 391 228 392 229 
rect 394 228 395 229 
rect 391 233 392 234 
rect 394 233 395 234 
<< m2 >>
rect 391 228 392 229 
rect 394 228 395 229 
rect 391 233 392 234 
rect 394 233 395 234 
<< m2c >>
rect 391 228 392 229 
rect 394 228 395 229 
rect 391 233 392 234 
rect 394 233 395 234 
<< labels >>
rlabel pdiffusion 103 138 104 139  0 t = 1
rlabel pdiffusion 106 138 107 139  0 t = 2
rlabel pdiffusion 103 143 104 144  0 t = 3
rlabel pdiffusion 106 143 107 144  0 t = 4
rlabel pdiffusion 102 138 108 144 0 cell no = 153
<< m1 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2 >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< m2c >>
rect 103 138 104 139 
rect 106 138 107 139 
rect 103 143 104 144 
rect 106 143 107 144 
<< labels >>
rlabel pdiffusion 175 48 176 49  0 t = 1
rlabel pdiffusion 178 48 179 49  0 t = 2
rlabel pdiffusion 175 53 176 54  0 t = 3
rlabel pdiffusion 178 53 179 54  0 t = 4
rlabel pdiffusion 174 48 180 54 0 cell no = 154
<< m1 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2 >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< m2c >>
rect 175 48 176 49 
rect 178 48 179 49 
rect 175 53 176 54 
rect 178 53 179 54 
<< labels >>
rlabel pdiffusion 481 84 482 85  0 t = 1
rlabel pdiffusion 484 84 485 85  0 t = 2
rlabel pdiffusion 481 89 482 90  0 t = 3
rlabel pdiffusion 484 89 485 90  0 t = 4
rlabel pdiffusion 480 84 486 90 0 cell no = 155
<< m1 >>
rect 481 84 482 85 
rect 484 84 485 85 
rect 481 89 482 90 
rect 484 89 485 90 
<< m2 >>
rect 481 84 482 85 
rect 484 84 485 85 
rect 481 89 482 90 
rect 484 89 485 90 
<< m2c >>
rect 481 84 482 85 
rect 484 84 485 85 
rect 481 89 482 90 
rect 484 89 485 90 
<< labels >>
rlabel pdiffusion 373 66 374 67  0 t = 1
rlabel pdiffusion 376 66 377 67  0 t = 2
rlabel pdiffusion 373 71 374 72  0 t = 3
rlabel pdiffusion 376 71 377 72  0 t = 4
rlabel pdiffusion 372 66 378 72 0 cell no = 156
<< m1 >>
rect 373 66 374 67 
rect 376 66 377 67 
rect 373 71 374 72 
rect 376 71 377 72 
<< m2 >>
rect 373 66 374 67 
rect 376 66 377 67 
rect 373 71 374 72 
rect 376 71 377 72 
<< m2c >>
rect 373 66 374 67 
rect 376 66 377 67 
rect 373 71 374 72 
rect 376 71 377 72 
<< labels >>
rlabel pdiffusion 211 282 212 283  0 t = 1
rlabel pdiffusion 214 282 215 283  0 t = 2
rlabel pdiffusion 211 287 212 288  0 t = 3
rlabel pdiffusion 214 287 215 288  0 t = 4
rlabel pdiffusion 210 282 216 288 0 cell no = 157
<< m1 >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< m2 >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< m2c >>
rect 211 282 212 283 
rect 214 282 215 283 
rect 211 287 212 288 
rect 214 287 215 288 
<< labels >>
rlabel pdiffusion 31 48 32 49  0 t = 1
rlabel pdiffusion 34 48 35 49  0 t = 2
rlabel pdiffusion 31 53 32 54  0 t = 3
rlabel pdiffusion 34 53 35 54  0 t = 4
rlabel pdiffusion 30 48 36 54 0 cell no = 158
<< m1 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2 >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< m2c >>
rect 31 48 32 49 
rect 34 48 35 49 
rect 31 53 32 54 
rect 34 53 35 54 
<< labels >>
rlabel pdiffusion 193 282 194 283  0 t = 1
rlabel pdiffusion 196 282 197 283  0 t = 2
rlabel pdiffusion 193 287 194 288  0 t = 3
rlabel pdiffusion 196 287 197 288  0 t = 4
rlabel pdiffusion 192 282 198 288 0 cell no = 159
<< m1 >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< m2 >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< m2c >>
rect 193 282 194 283 
rect 196 282 197 283 
rect 193 287 194 288 
rect 196 287 197 288 
<< labels >>
rlabel pdiffusion 481 30 482 31  0 t = 1
rlabel pdiffusion 484 30 485 31  0 t = 2
rlabel pdiffusion 481 35 482 36  0 t = 3
rlabel pdiffusion 484 35 485 36  0 t = 4
rlabel pdiffusion 480 30 486 36 0 cell no = 160
<< m1 >>
rect 481 30 482 31 
rect 484 30 485 31 
rect 481 35 482 36 
rect 484 35 485 36 
<< m2 >>
rect 481 30 482 31 
rect 484 30 485 31 
rect 481 35 482 36 
rect 484 35 485 36 
<< m2c >>
rect 481 30 482 31 
rect 484 30 485 31 
rect 481 35 482 36 
rect 484 35 485 36 
<< labels >>
rlabel pdiffusion 157 174 158 175  0 t = 1
rlabel pdiffusion 160 174 161 175  0 t = 2
rlabel pdiffusion 157 179 158 180  0 t = 3
rlabel pdiffusion 160 179 161 180  0 t = 4
rlabel pdiffusion 156 174 162 180 0 cell no = 161
<< m1 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2 >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< m2c >>
rect 157 174 158 175 
rect 160 174 161 175 
rect 157 179 158 180 
rect 160 179 161 180 
<< labels >>
rlabel pdiffusion 373 156 374 157  0 t = 1
rlabel pdiffusion 376 156 377 157  0 t = 2
rlabel pdiffusion 373 161 374 162  0 t = 3
rlabel pdiffusion 376 161 377 162  0 t = 4
rlabel pdiffusion 372 156 378 162 0 cell no = 162
<< m1 >>
rect 373 156 374 157 
rect 376 156 377 157 
rect 373 161 374 162 
rect 376 161 377 162 
<< m2 >>
rect 373 156 374 157 
rect 376 156 377 157 
rect 373 161 374 162 
rect 376 161 377 162 
<< m2c >>
rect 373 156 374 157 
rect 376 156 377 157 
rect 373 161 374 162 
rect 376 161 377 162 
<< labels >>
rlabel pdiffusion 373 408 374 409  0 t = 1
rlabel pdiffusion 376 408 377 409  0 t = 2
rlabel pdiffusion 373 413 374 414  0 t = 3
rlabel pdiffusion 376 413 377 414  0 t = 4
rlabel pdiffusion 372 408 378 414 0 cell no = 163
<< m1 >>
rect 373 408 374 409 
rect 376 408 377 409 
rect 373 413 374 414 
rect 376 413 377 414 
<< m2 >>
rect 373 408 374 409 
rect 376 408 377 409 
rect 373 413 374 414 
rect 376 413 377 414 
<< m2c >>
rect 373 408 374 409 
rect 376 408 377 409 
rect 373 413 374 414 
rect 376 413 377 414 
<< labels >>
rlabel pdiffusion 337 102 338 103  0 t = 1
rlabel pdiffusion 340 102 341 103  0 t = 2
rlabel pdiffusion 337 107 338 108  0 t = 3
rlabel pdiffusion 340 107 341 108  0 t = 4
rlabel pdiffusion 336 102 342 108 0 cell no = 164
<< m1 >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< m2 >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< m2c >>
rect 337 102 338 103 
rect 340 102 341 103 
rect 337 107 338 108 
rect 340 107 341 108 
<< labels >>
rlabel pdiffusion 319 30 320 31  0 t = 1
rlabel pdiffusion 322 30 323 31  0 t = 2
rlabel pdiffusion 319 35 320 36  0 t = 3
rlabel pdiffusion 322 35 323 36  0 t = 4
rlabel pdiffusion 318 30 324 36 0 cell no = 165
<< m1 >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< m2 >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< m2c >>
rect 319 30 320 31 
rect 322 30 323 31 
rect 319 35 320 36 
rect 322 35 323 36 
<< labels >>
rlabel pdiffusion 391 264 392 265  0 t = 1
rlabel pdiffusion 394 264 395 265  0 t = 2
rlabel pdiffusion 391 269 392 270  0 t = 3
rlabel pdiffusion 394 269 395 270  0 t = 4
rlabel pdiffusion 390 264 396 270 0 cell no = 166
<< m1 >>
rect 391 264 392 265 
rect 394 264 395 265 
rect 391 269 392 270 
rect 394 269 395 270 
<< m2 >>
rect 391 264 392 265 
rect 394 264 395 265 
rect 391 269 392 270 
rect 394 269 395 270 
<< m2c >>
rect 391 264 392 265 
rect 394 264 395 265 
rect 391 269 392 270 
rect 394 269 395 270 
<< labels >>
rlabel pdiffusion 517 66 518 67  0 t = 1
rlabel pdiffusion 520 66 521 67  0 t = 2
rlabel pdiffusion 517 71 518 72  0 t = 3
rlabel pdiffusion 520 71 521 72  0 t = 4
rlabel pdiffusion 516 66 522 72 0 cell no = 167
<< m1 >>
rect 517 66 518 67 
rect 520 66 521 67 
rect 517 71 518 72 
rect 520 71 521 72 
<< m2 >>
rect 517 66 518 67 
rect 520 66 521 67 
rect 517 71 518 72 
rect 520 71 521 72 
<< m2c >>
rect 517 66 518 67 
rect 520 66 521 67 
rect 517 71 518 72 
rect 520 71 521 72 
<< labels >>
rlabel pdiffusion 499 12 500 13  0 t = 1
rlabel pdiffusion 502 12 503 13  0 t = 2
rlabel pdiffusion 499 17 500 18  0 t = 3
rlabel pdiffusion 502 17 503 18  0 t = 4
rlabel pdiffusion 498 12 504 18 0 cell no = 168
<< m1 >>
rect 499 12 500 13 
rect 502 12 503 13 
rect 499 17 500 18 
rect 502 17 503 18 
<< m2 >>
rect 499 12 500 13 
rect 502 12 503 13 
rect 499 17 500 18 
rect 502 17 503 18 
<< m2c >>
rect 499 12 500 13 
rect 502 12 503 13 
rect 499 17 500 18 
rect 502 17 503 18 
<< labels >>
rlabel pdiffusion 355 120 356 121  0 t = 1
rlabel pdiffusion 358 120 359 121  0 t = 2
rlabel pdiffusion 355 125 356 126  0 t = 3
rlabel pdiffusion 358 125 359 126  0 t = 4
rlabel pdiffusion 354 120 360 126 0 cell no = 169
<< m1 >>
rect 355 120 356 121 
rect 358 120 359 121 
rect 355 125 356 126 
rect 358 125 359 126 
<< m2 >>
rect 355 120 356 121 
rect 358 120 359 121 
rect 355 125 356 126 
rect 358 125 359 126 
<< m2c >>
rect 355 120 356 121 
rect 358 120 359 121 
rect 355 125 356 126 
rect 358 125 359 126 
<< labels >>
rlabel pdiffusion 463 12 464 13  0 t = 1
rlabel pdiffusion 466 12 467 13  0 t = 2
rlabel pdiffusion 463 17 464 18  0 t = 3
rlabel pdiffusion 466 17 467 18  0 t = 4
rlabel pdiffusion 462 12 468 18 0 cell no = 170
<< m1 >>
rect 463 12 464 13 
rect 466 12 467 13 
rect 463 17 464 18 
rect 466 17 467 18 
<< m2 >>
rect 463 12 464 13 
rect 466 12 467 13 
rect 463 17 464 18 
rect 466 17 467 18 
<< m2c >>
rect 463 12 464 13 
rect 466 12 467 13 
rect 463 17 464 18 
rect 466 17 467 18 
<< labels >>
rlabel pdiffusion 193 444 194 445  0 t = 1
rlabel pdiffusion 196 444 197 445  0 t = 2
rlabel pdiffusion 193 449 194 450  0 t = 3
rlabel pdiffusion 196 449 197 450  0 t = 4
rlabel pdiffusion 192 444 198 450 0 cell no = 171
<< m1 >>
rect 193 444 194 445 
rect 196 444 197 445 
rect 193 449 194 450 
rect 196 449 197 450 
<< m2 >>
rect 193 444 194 445 
rect 196 444 197 445 
rect 193 449 194 450 
rect 196 449 197 450 
<< m2c >>
rect 193 444 194 445 
rect 196 444 197 445 
rect 193 449 194 450 
rect 196 449 197 450 
<< labels >>
rlabel pdiffusion 481 12 482 13  0 t = 1
rlabel pdiffusion 484 12 485 13  0 t = 2
rlabel pdiffusion 481 17 482 18  0 t = 3
rlabel pdiffusion 484 17 485 18  0 t = 4
rlabel pdiffusion 480 12 486 18 0 cell no = 172
<< m1 >>
rect 481 12 482 13 
rect 484 12 485 13 
rect 481 17 482 18 
rect 484 17 485 18 
<< m2 >>
rect 481 12 482 13 
rect 484 12 485 13 
rect 481 17 482 18 
rect 484 17 485 18 
<< m2c >>
rect 481 12 482 13 
rect 484 12 485 13 
rect 481 17 482 18 
rect 484 17 485 18 
<< labels >>
rlabel pdiffusion 445 138 446 139  0 t = 1
rlabel pdiffusion 448 138 449 139  0 t = 2
rlabel pdiffusion 445 143 446 144  0 t = 3
rlabel pdiffusion 448 143 449 144  0 t = 4
rlabel pdiffusion 444 138 450 144 0 cell no = 173
<< m1 >>
rect 445 138 446 139 
rect 448 138 449 139 
rect 445 143 446 144 
rect 448 143 449 144 
<< m2 >>
rect 445 138 446 139 
rect 448 138 449 139 
rect 445 143 446 144 
rect 448 143 449 144 
<< m2c >>
rect 445 138 446 139 
rect 448 138 449 139 
rect 445 143 446 144 
rect 448 143 449 144 
<< labels >>
rlabel pdiffusion 355 12 356 13  0 t = 1
rlabel pdiffusion 358 12 359 13  0 t = 2
rlabel pdiffusion 355 17 356 18  0 t = 3
rlabel pdiffusion 358 17 359 18  0 t = 4
rlabel pdiffusion 354 12 360 18 0 cell no = 174
<< m1 >>
rect 355 12 356 13 
rect 358 12 359 13 
rect 355 17 356 18 
rect 358 17 359 18 
<< m2 >>
rect 355 12 356 13 
rect 358 12 359 13 
rect 355 17 356 18 
rect 358 17 359 18 
<< m2c >>
rect 355 12 356 13 
rect 358 12 359 13 
rect 355 17 356 18 
rect 358 17 359 18 
<< labels >>
rlabel pdiffusion 67 66 68 67  0 t = 1
rlabel pdiffusion 70 66 71 67  0 t = 2
rlabel pdiffusion 67 71 68 72  0 t = 3
rlabel pdiffusion 70 71 71 72  0 t = 4
rlabel pdiffusion 66 66 72 72 0 cell no = 175
<< m1 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2 >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< m2c >>
rect 67 66 68 67 
rect 70 66 71 67 
rect 67 71 68 72 
rect 70 71 71 72 
<< labels >>
rlabel pdiffusion 85 174 86 175  0 t = 1
rlabel pdiffusion 88 174 89 175  0 t = 2
rlabel pdiffusion 85 179 86 180  0 t = 3
rlabel pdiffusion 88 179 89 180  0 t = 4
rlabel pdiffusion 84 174 90 180 0 cell no = 176
<< m1 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2 >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< m2c >>
rect 85 174 86 175 
rect 88 174 89 175 
rect 85 179 86 180 
rect 88 179 89 180 
<< labels >>
rlabel pdiffusion 85 84 86 85  0 t = 1
rlabel pdiffusion 88 84 89 85  0 t = 2
rlabel pdiffusion 85 89 86 90  0 t = 3
rlabel pdiffusion 88 89 89 90  0 t = 4
rlabel pdiffusion 84 84 90 90 0 cell no = 177
<< m1 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2 >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< m2c >>
rect 85 84 86 85 
rect 88 84 89 85 
rect 85 89 86 90 
rect 88 89 89 90 
<< labels >>
rlabel pdiffusion 157 48 158 49  0 t = 1
rlabel pdiffusion 160 48 161 49  0 t = 2
rlabel pdiffusion 157 53 158 54  0 t = 3
rlabel pdiffusion 160 53 161 54  0 t = 4
rlabel pdiffusion 156 48 162 54 0 cell no = 178
<< m1 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2 >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< m2c >>
rect 157 48 158 49 
rect 160 48 161 49 
rect 157 53 158 54 
rect 160 53 161 54 
<< labels >>
rlabel pdiffusion 301 102 302 103  0 t = 1
rlabel pdiffusion 304 102 305 103  0 t = 2
rlabel pdiffusion 301 107 302 108  0 t = 3
rlabel pdiffusion 304 107 305 108  0 t = 4
rlabel pdiffusion 300 102 306 108 0 cell no = 179
<< m1 >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< m2 >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< m2c >>
rect 301 102 302 103 
rect 304 102 305 103 
rect 301 107 302 108 
rect 304 107 305 108 
<< labels >>
rlabel pdiffusion 247 138 248 139  0 t = 1
rlabel pdiffusion 250 138 251 139  0 t = 2
rlabel pdiffusion 247 143 248 144  0 t = 3
rlabel pdiffusion 250 143 251 144  0 t = 4
rlabel pdiffusion 246 138 252 144 0 cell no = 180
<< m1 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2 >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< m2c >>
rect 247 138 248 139 
rect 250 138 251 139 
rect 247 143 248 144 
rect 250 143 251 144 
<< labels >>
rlabel pdiffusion 139 48 140 49  0 t = 1
rlabel pdiffusion 142 48 143 49  0 t = 2
rlabel pdiffusion 139 53 140 54  0 t = 3
rlabel pdiffusion 142 53 143 54  0 t = 4
rlabel pdiffusion 138 48 144 54 0 cell no = 181
<< m1 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2 >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< m2c >>
rect 139 48 140 49 
rect 142 48 143 49 
rect 139 53 140 54 
rect 142 53 143 54 
<< labels >>
rlabel pdiffusion 103 102 104 103  0 t = 1
rlabel pdiffusion 106 102 107 103  0 t = 2
rlabel pdiffusion 103 107 104 108  0 t = 3
rlabel pdiffusion 106 107 107 108  0 t = 4
rlabel pdiffusion 102 102 108 108 0 cell no = 182
<< m1 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2 >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< m2c >>
rect 103 102 104 103 
rect 106 102 107 103 
rect 103 107 104 108 
rect 106 107 107 108 
<< labels >>
rlabel pdiffusion 193 12 194 13  0 t = 1
rlabel pdiffusion 196 12 197 13  0 t = 2
rlabel pdiffusion 193 17 194 18  0 t = 3
rlabel pdiffusion 196 17 197 18  0 t = 4
rlabel pdiffusion 192 12 198 18 0 cell no = 183
<< m1 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2 >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< m2c >>
rect 193 12 194 13 
rect 196 12 197 13 
rect 193 17 194 18 
rect 196 17 197 18 
<< labels >>
rlabel pdiffusion 157 336 158 337  0 t = 1
rlabel pdiffusion 160 336 161 337  0 t = 2
rlabel pdiffusion 157 341 158 342  0 t = 3
rlabel pdiffusion 160 341 161 342  0 t = 4
rlabel pdiffusion 156 336 162 342 0 cell no = 184
<< m1 >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< m2 >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< m2c >>
rect 157 336 158 337 
rect 160 336 161 337 
rect 157 341 158 342 
rect 160 341 161 342 
<< labels >>
rlabel pdiffusion 427 426 428 427  0 t = 1
rlabel pdiffusion 430 426 431 427  0 t = 2
rlabel pdiffusion 427 431 428 432  0 t = 3
rlabel pdiffusion 430 431 431 432  0 t = 4
rlabel pdiffusion 426 426 432 432 0 cell no = 185
<< m1 >>
rect 427 426 428 427 
rect 430 426 431 427 
rect 427 431 428 432 
rect 430 431 431 432 
<< m2 >>
rect 427 426 428 427 
rect 430 426 431 427 
rect 427 431 428 432 
rect 430 431 431 432 
<< m2c >>
rect 427 426 428 427 
rect 430 426 431 427 
rect 427 431 428 432 
rect 430 431 431 432 
<< labels >>
rlabel pdiffusion 67 84 68 85  0 t = 1
rlabel pdiffusion 70 84 71 85  0 t = 2
rlabel pdiffusion 67 89 68 90  0 t = 3
rlabel pdiffusion 70 89 71 90  0 t = 4
rlabel pdiffusion 66 84 72 90 0 cell no = 186
<< m1 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2 >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< m2c >>
rect 67 84 68 85 
rect 70 84 71 85 
rect 67 89 68 90 
rect 70 89 71 90 
<< labels >>
rlabel pdiffusion 13 264 14 265  0 t = 1
rlabel pdiffusion 16 264 17 265  0 t = 2
rlabel pdiffusion 13 269 14 270  0 t = 3
rlabel pdiffusion 16 269 17 270  0 t = 4
rlabel pdiffusion 12 264 18 270 0 cell no = 187
<< m1 >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< m2 >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< m2c >>
rect 13 264 14 265 
rect 16 264 17 265 
rect 13 269 14 270 
rect 16 269 17 270 
<< labels >>
rlabel pdiffusion 355 192 356 193  0 t = 1
rlabel pdiffusion 358 192 359 193  0 t = 2
rlabel pdiffusion 355 197 356 198  0 t = 3
rlabel pdiffusion 358 197 359 198  0 t = 4
rlabel pdiffusion 354 192 360 198 0 cell no = 188
<< m1 >>
rect 355 192 356 193 
rect 358 192 359 193 
rect 355 197 356 198 
rect 358 197 359 198 
<< m2 >>
rect 355 192 356 193 
rect 358 192 359 193 
rect 355 197 356 198 
rect 358 197 359 198 
<< m2c >>
rect 355 192 356 193 
rect 358 192 359 193 
rect 355 197 356 198 
rect 358 197 359 198 
<< labels >>
rlabel pdiffusion 67 102 68 103  0 t = 1
rlabel pdiffusion 70 102 71 103  0 t = 2
rlabel pdiffusion 67 107 68 108  0 t = 3
rlabel pdiffusion 70 107 71 108  0 t = 4
rlabel pdiffusion 66 102 72 108 0 cell no = 189
<< m1 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2 >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< m2c >>
rect 67 102 68 103 
rect 70 102 71 103 
rect 67 107 68 108 
rect 70 107 71 108 
<< labels >>
rlabel pdiffusion 283 138 284 139  0 t = 1
rlabel pdiffusion 286 138 287 139  0 t = 2
rlabel pdiffusion 283 143 284 144  0 t = 3
rlabel pdiffusion 286 143 287 144  0 t = 4
rlabel pdiffusion 282 138 288 144 0 cell no = 190
<< m1 >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< m2 >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< m2c >>
rect 283 138 284 139 
rect 286 138 287 139 
rect 283 143 284 144 
rect 286 143 287 144 
<< labels >>
rlabel pdiffusion 265 210 266 211  0 t = 1
rlabel pdiffusion 268 210 269 211  0 t = 2
rlabel pdiffusion 265 215 266 216  0 t = 3
rlabel pdiffusion 268 215 269 216  0 t = 4
rlabel pdiffusion 264 210 270 216 0 cell no = 191
<< m1 >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< m2 >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< m2c >>
rect 265 210 266 211 
rect 268 210 269 211 
rect 265 215 266 216 
rect 268 215 269 216 
<< labels >>
rlabel pdiffusion 517 282 518 283  0 t = 1
rlabel pdiffusion 520 282 521 283  0 t = 2
rlabel pdiffusion 517 287 518 288  0 t = 3
rlabel pdiffusion 520 287 521 288  0 t = 4
rlabel pdiffusion 516 282 522 288 0 cell no = 192
<< m1 >>
rect 517 282 518 283 
rect 520 282 521 283 
rect 517 287 518 288 
rect 520 287 521 288 
<< m2 >>
rect 517 282 518 283 
rect 520 282 521 283 
rect 517 287 518 288 
rect 520 287 521 288 
<< m2c >>
rect 517 282 518 283 
rect 520 282 521 283 
rect 517 287 518 288 
rect 520 287 521 288 
<< labels >>
rlabel pdiffusion 121 372 122 373  0 t = 1
rlabel pdiffusion 124 372 125 373  0 t = 2
rlabel pdiffusion 121 377 122 378  0 t = 3
rlabel pdiffusion 124 377 125 378  0 t = 4
rlabel pdiffusion 120 372 126 378 0 cell no = 193
<< m1 >>
rect 121 372 122 373 
rect 124 372 125 373 
rect 121 377 122 378 
rect 124 377 125 378 
<< m2 >>
rect 121 372 122 373 
rect 124 372 125 373 
rect 121 377 122 378 
rect 124 377 125 378 
<< m2c >>
rect 121 372 122 373 
rect 124 372 125 373 
rect 121 377 122 378 
rect 124 377 125 378 
<< labels >>
rlabel pdiffusion 283 156 284 157  0 t = 1
rlabel pdiffusion 286 156 287 157  0 t = 2
rlabel pdiffusion 283 161 284 162  0 t = 3
rlabel pdiffusion 286 161 287 162  0 t = 4
rlabel pdiffusion 282 156 288 162 0 cell no = 194
<< m1 >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< m2 >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< m2c >>
rect 283 156 284 157 
rect 286 156 287 157 
rect 283 161 284 162 
rect 286 161 287 162 
<< labels >>
rlabel pdiffusion 373 48 374 49  0 t = 1
rlabel pdiffusion 376 48 377 49  0 t = 2
rlabel pdiffusion 373 53 374 54  0 t = 3
rlabel pdiffusion 376 53 377 54  0 t = 4
rlabel pdiffusion 372 48 378 54 0 cell no = 195
<< m1 >>
rect 373 48 374 49 
rect 376 48 377 49 
rect 373 53 374 54 
rect 376 53 377 54 
<< m2 >>
rect 373 48 374 49 
rect 376 48 377 49 
rect 373 53 374 54 
rect 376 53 377 54 
<< m2c >>
rect 373 48 374 49 
rect 376 48 377 49 
rect 373 53 374 54 
rect 376 53 377 54 
<< labels >>
rlabel pdiffusion 481 246 482 247  0 t = 1
rlabel pdiffusion 484 246 485 247  0 t = 2
rlabel pdiffusion 481 251 482 252  0 t = 3
rlabel pdiffusion 484 251 485 252  0 t = 4
rlabel pdiffusion 480 246 486 252 0 cell no = 196
<< m1 >>
rect 481 246 482 247 
rect 484 246 485 247 
rect 481 251 482 252 
rect 484 251 485 252 
<< m2 >>
rect 481 246 482 247 
rect 484 246 485 247 
rect 481 251 482 252 
rect 484 251 485 252 
<< m2c >>
rect 481 246 482 247 
rect 484 246 485 247 
rect 481 251 482 252 
rect 484 251 485 252 
<< labels >>
rlabel pdiffusion 517 102 518 103  0 t = 1
rlabel pdiffusion 520 102 521 103  0 t = 2
rlabel pdiffusion 517 107 518 108  0 t = 3
rlabel pdiffusion 520 107 521 108  0 t = 4
rlabel pdiffusion 516 102 522 108 0 cell no = 197
<< m1 >>
rect 517 102 518 103 
rect 520 102 521 103 
rect 517 107 518 108 
rect 520 107 521 108 
<< m2 >>
rect 517 102 518 103 
rect 520 102 521 103 
rect 517 107 518 108 
rect 520 107 521 108 
<< m2c >>
rect 517 102 518 103 
rect 520 102 521 103 
rect 517 107 518 108 
rect 520 107 521 108 
<< labels >>
rlabel pdiffusion 427 246 428 247  0 t = 1
rlabel pdiffusion 430 246 431 247  0 t = 2
rlabel pdiffusion 427 251 428 252  0 t = 3
rlabel pdiffusion 430 251 431 252  0 t = 4
rlabel pdiffusion 426 246 432 252 0 cell no = 198
<< m1 >>
rect 427 246 428 247 
rect 430 246 431 247 
rect 427 251 428 252 
rect 430 251 431 252 
<< m2 >>
rect 427 246 428 247 
rect 430 246 431 247 
rect 427 251 428 252 
rect 430 251 431 252 
<< m2c >>
rect 427 246 428 247 
rect 430 246 431 247 
rect 427 251 428 252 
rect 430 251 431 252 
<< labels >>
rlabel pdiffusion 517 120 518 121  0 t = 1
rlabel pdiffusion 520 120 521 121  0 t = 2
rlabel pdiffusion 517 125 518 126  0 t = 3
rlabel pdiffusion 520 125 521 126  0 t = 4
rlabel pdiffusion 516 120 522 126 0 cell no = 199
<< m1 >>
rect 517 120 518 121 
rect 520 120 521 121 
rect 517 125 518 126 
rect 520 125 521 126 
<< m2 >>
rect 517 120 518 121 
rect 520 120 521 121 
rect 517 125 518 126 
rect 520 125 521 126 
<< m2c >>
rect 517 120 518 121 
rect 520 120 521 121 
rect 517 125 518 126 
rect 520 125 521 126 
<< labels >>
rlabel pdiffusion 463 48 464 49  0 t = 1
rlabel pdiffusion 466 48 467 49  0 t = 2
rlabel pdiffusion 463 53 464 54  0 t = 3
rlabel pdiffusion 466 53 467 54  0 t = 4
rlabel pdiffusion 462 48 468 54 0 cell no = 200
<< m1 >>
rect 463 48 464 49 
rect 466 48 467 49 
rect 463 53 464 54 
rect 466 53 467 54 
<< m2 >>
rect 463 48 464 49 
rect 466 48 467 49 
rect 463 53 464 54 
rect 466 53 467 54 
<< m2c >>
rect 463 48 464 49 
rect 466 48 467 49 
rect 463 53 464 54 
rect 466 53 467 54 
<< labels >>
rlabel pdiffusion 463 156 464 157  0 t = 1
rlabel pdiffusion 466 156 467 157  0 t = 2
rlabel pdiffusion 463 161 464 162  0 t = 3
rlabel pdiffusion 466 161 467 162  0 t = 4
rlabel pdiffusion 462 156 468 162 0 cell no = 201
<< m1 >>
rect 463 156 464 157 
rect 466 156 467 157 
rect 463 161 464 162 
rect 466 161 467 162 
<< m2 >>
rect 463 156 464 157 
rect 466 156 467 157 
rect 463 161 464 162 
rect 466 161 467 162 
<< m2c >>
rect 463 156 464 157 
rect 466 156 467 157 
rect 463 161 464 162 
rect 466 161 467 162 
<< labels >>
rlabel pdiffusion 499 192 500 193  0 t = 1
rlabel pdiffusion 502 192 503 193  0 t = 2
rlabel pdiffusion 499 197 500 198  0 t = 3
rlabel pdiffusion 502 197 503 198  0 t = 4
rlabel pdiffusion 498 192 504 198 0 cell no = 202
<< m1 >>
rect 499 192 500 193 
rect 502 192 503 193 
rect 499 197 500 198 
rect 502 197 503 198 
<< m2 >>
rect 499 192 500 193 
rect 502 192 503 193 
rect 499 197 500 198 
rect 502 197 503 198 
<< m2c >>
rect 499 192 500 193 
rect 502 192 503 193 
rect 499 197 500 198 
rect 502 197 503 198 
<< labels >>
rlabel pdiffusion 445 300 446 301  0 t = 1
rlabel pdiffusion 448 300 449 301  0 t = 2
rlabel pdiffusion 445 305 446 306  0 t = 3
rlabel pdiffusion 448 305 449 306  0 t = 4
rlabel pdiffusion 444 300 450 306 0 cell no = 203
<< m1 >>
rect 445 300 446 301 
rect 448 300 449 301 
rect 445 305 446 306 
rect 448 305 449 306 
<< m2 >>
rect 445 300 446 301 
rect 448 300 449 301 
rect 445 305 446 306 
rect 448 305 449 306 
<< m2c >>
rect 445 300 446 301 
rect 448 300 449 301 
rect 445 305 446 306 
rect 448 305 449 306 
<< labels >>
rlabel pdiffusion 121 156 122 157  0 t = 1
rlabel pdiffusion 124 156 125 157  0 t = 2
rlabel pdiffusion 121 161 122 162  0 t = 3
rlabel pdiffusion 124 161 125 162  0 t = 4
rlabel pdiffusion 120 156 126 162 0 cell no = 204
<< m1 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2 >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< m2c >>
rect 121 156 122 157 
rect 124 156 125 157 
rect 121 161 122 162 
rect 124 161 125 162 
<< labels >>
rlabel pdiffusion 13 138 14 139  0 t = 1
rlabel pdiffusion 16 138 17 139  0 t = 2
rlabel pdiffusion 13 143 14 144  0 t = 3
rlabel pdiffusion 16 143 17 144  0 t = 4
rlabel pdiffusion 12 138 18 144 0 cell no = 205
<< m1 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2 >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< m2c >>
rect 13 138 14 139 
rect 16 138 17 139 
rect 13 143 14 144 
rect 16 143 17 144 
<< labels >>
rlabel pdiffusion 103 12 104 13  0 t = 1
rlabel pdiffusion 106 12 107 13  0 t = 2
rlabel pdiffusion 103 17 104 18  0 t = 3
rlabel pdiffusion 106 17 107 18  0 t = 4
rlabel pdiffusion 102 12 108 18 0 cell no = 206
<< m1 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2 >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< m2c >>
rect 103 12 104 13 
rect 106 12 107 13 
rect 103 17 104 18 
rect 106 17 107 18 
<< labels >>
rlabel pdiffusion 229 30 230 31  0 t = 1
rlabel pdiffusion 232 30 233 31  0 t = 2
rlabel pdiffusion 229 35 230 36  0 t = 3
rlabel pdiffusion 232 35 233 36  0 t = 4
rlabel pdiffusion 228 30 234 36 0 cell no = 207
<< m1 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2 >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< m2c >>
rect 229 30 230 31 
rect 232 30 233 31 
rect 229 35 230 36 
rect 232 35 233 36 
<< labels >>
rlabel pdiffusion 319 246 320 247  0 t = 1
rlabel pdiffusion 322 246 323 247  0 t = 2
rlabel pdiffusion 319 251 320 252  0 t = 3
rlabel pdiffusion 322 251 323 252  0 t = 4
rlabel pdiffusion 318 246 324 252 0 cell no = 208
<< m1 >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< m2 >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< m2c >>
rect 319 246 320 247 
rect 322 246 323 247 
rect 319 251 320 252 
rect 322 251 323 252 
<< labels >>
rlabel pdiffusion 49 192 50 193  0 t = 1
rlabel pdiffusion 52 192 53 193  0 t = 2
rlabel pdiffusion 49 197 50 198  0 t = 3
rlabel pdiffusion 52 197 53 198  0 t = 4
rlabel pdiffusion 48 192 54 198 0 cell no = 209
<< m1 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2 >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< m2c >>
rect 49 192 50 193 
rect 52 192 53 193 
rect 49 197 50 198 
rect 52 197 53 198 
<< labels >>
rlabel pdiffusion 121 318 122 319  0 t = 1
rlabel pdiffusion 124 318 125 319  0 t = 2
rlabel pdiffusion 121 323 122 324  0 t = 3
rlabel pdiffusion 124 323 125 324  0 t = 4
rlabel pdiffusion 120 318 126 324 0 cell no = 210
<< m1 >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< m2 >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< m2c >>
rect 121 318 122 319 
rect 124 318 125 319 
rect 121 323 122 324 
rect 124 323 125 324 
<< labels >>
rlabel pdiffusion 121 84 122 85  0 t = 1
rlabel pdiffusion 124 84 125 85  0 t = 2
rlabel pdiffusion 121 89 122 90  0 t = 3
rlabel pdiffusion 124 89 125 90  0 t = 4
rlabel pdiffusion 120 84 126 90 0 cell no = 211
<< m1 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2 >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< m2c >>
rect 121 84 122 85 
rect 124 84 125 85 
rect 121 89 122 90 
rect 124 89 125 90 
<< labels >>
rlabel pdiffusion 229 516 230 517  0 t = 1
rlabel pdiffusion 232 516 233 517  0 t = 2
rlabel pdiffusion 229 521 230 522  0 t = 3
rlabel pdiffusion 232 521 233 522  0 t = 4
rlabel pdiffusion 228 516 234 522 0 cell no = 212
<< m1 >>
rect 229 516 230 517 
rect 232 516 233 517 
rect 229 521 230 522 
rect 232 521 233 522 
<< m2 >>
rect 229 516 230 517 
rect 232 516 233 517 
rect 229 521 230 522 
rect 232 521 233 522 
<< m2c >>
rect 229 516 230 517 
rect 232 516 233 517 
rect 229 521 230 522 
rect 232 521 233 522 
<< labels >>
rlabel pdiffusion 427 102 428 103  0 t = 1
rlabel pdiffusion 430 102 431 103  0 t = 2
rlabel pdiffusion 427 107 428 108  0 t = 3
rlabel pdiffusion 430 107 431 108  0 t = 4
rlabel pdiffusion 426 102 432 108 0 cell no = 213
<< m1 >>
rect 427 102 428 103 
rect 430 102 431 103 
rect 427 107 428 108 
rect 430 107 431 108 
<< m2 >>
rect 427 102 428 103 
rect 430 102 431 103 
rect 427 107 428 108 
rect 430 107 431 108 
<< m2c >>
rect 427 102 428 103 
rect 430 102 431 103 
rect 427 107 428 108 
rect 430 107 431 108 
<< labels >>
rlabel pdiffusion 247 354 248 355  0 t = 1
rlabel pdiffusion 250 354 251 355  0 t = 2
rlabel pdiffusion 247 359 248 360  0 t = 3
rlabel pdiffusion 250 359 251 360  0 t = 4
rlabel pdiffusion 246 354 252 360 0 cell no = 214
<< m1 >>
rect 247 354 248 355 
rect 250 354 251 355 
rect 247 359 248 360 
rect 250 359 251 360 
<< m2 >>
rect 247 354 248 355 
rect 250 354 251 355 
rect 247 359 248 360 
rect 250 359 251 360 
<< m2c >>
rect 247 354 248 355 
rect 250 354 251 355 
rect 247 359 248 360 
rect 250 359 251 360 
<< labels >>
rlabel pdiffusion 211 102 212 103  0 t = 1
rlabel pdiffusion 214 102 215 103  0 t = 2
rlabel pdiffusion 211 107 212 108  0 t = 3
rlabel pdiffusion 214 107 215 108  0 t = 4
rlabel pdiffusion 210 102 216 108 0 cell no = 215
<< m1 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2 >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< m2c >>
rect 211 102 212 103 
rect 214 102 215 103 
rect 211 107 212 108 
rect 214 107 215 108 
<< labels >>
rlabel pdiffusion 139 462 140 463  0 t = 1
rlabel pdiffusion 142 462 143 463  0 t = 2
rlabel pdiffusion 139 467 140 468  0 t = 3
rlabel pdiffusion 142 467 143 468  0 t = 4
rlabel pdiffusion 138 462 144 468 0 cell no = 216
<< m1 >>
rect 139 462 140 463 
rect 142 462 143 463 
rect 139 467 140 468 
rect 142 467 143 468 
<< m2 >>
rect 139 462 140 463 
rect 142 462 143 463 
rect 139 467 140 468 
rect 142 467 143 468 
<< m2c >>
rect 139 462 140 463 
rect 142 462 143 463 
rect 139 467 140 468 
rect 142 467 143 468 
<< labels >>
rlabel pdiffusion 193 300 194 301  0 t = 1
rlabel pdiffusion 196 300 197 301  0 t = 2
rlabel pdiffusion 193 305 194 306  0 t = 3
rlabel pdiffusion 196 305 197 306  0 t = 4
rlabel pdiffusion 192 300 198 306 0 cell no = 217
<< m1 >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< m2 >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< m2c >>
rect 193 300 194 301 
rect 196 300 197 301 
rect 193 305 194 306 
rect 196 305 197 306 
<< labels >>
rlabel pdiffusion 67 228 68 229  0 t = 1
rlabel pdiffusion 70 228 71 229  0 t = 2
rlabel pdiffusion 67 233 68 234  0 t = 3
rlabel pdiffusion 70 233 71 234  0 t = 4
rlabel pdiffusion 66 228 72 234 0 cell no = 218
<< m1 >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< m2 >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< m2c >>
rect 67 228 68 229 
rect 70 228 71 229 
rect 67 233 68 234 
rect 70 233 71 234 
<< labels >>
rlabel pdiffusion 121 12 122 13  0 t = 1
rlabel pdiffusion 124 12 125 13  0 t = 2
rlabel pdiffusion 121 17 122 18  0 t = 3
rlabel pdiffusion 124 17 125 18  0 t = 4
rlabel pdiffusion 120 12 126 18 0 cell no = 219
<< m1 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2 >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< m2c >>
rect 121 12 122 13 
rect 124 12 125 13 
rect 121 17 122 18 
rect 124 17 125 18 
<< labels >>
rlabel pdiffusion 301 66 302 67  0 t = 1
rlabel pdiffusion 304 66 305 67  0 t = 2
rlabel pdiffusion 301 71 302 72  0 t = 3
rlabel pdiffusion 304 71 305 72  0 t = 4
rlabel pdiffusion 300 66 306 72 0 cell no = 220
<< m1 >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< m2 >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< m2c >>
rect 301 66 302 67 
rect 304 66 305 67 
rect 301 71 302 72 
rect 304 71 305 72 
<< labels >>
rlabel pdiffusion 175 138 176 139  0 t = 1
rlabel pdiffusion 178 138 179 139  0 t = 2
rlabel pdiffusion 175 143 176 144  0 t = 3
rlabel pdiffusion 178 143 179 144  0 t = 4
rlabel pdiffusion 174 138 180 144 0 cell no = 221
<< m1 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2 >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< m2c >>
rect 175 138 176 139 
rect 178 138 179 139 
rect 175 143 176 144 
rect 178 143 179 144 
<< labels >>
rlabel pdiffusion 445 102 446 103  0 t = 1
rlabel pdiffusion 448 102 449 103  0 t = 2
rlabel pdiffusion 445 107 446 108  0 t = 3
rlabel pdiffusion 448 107 449 108  0 t = 4
rlabel pdiffusion 444 102 450 108 0 cell no = 222
<< m1 >>
rect 445 102 446 103 
rect 448 102 449 103 
rect 445 107 446 108 
rect 448 107 449 108 
<< m2 >>
rect 445 102 446 103 
rect 448 102 449 103 
rect 445 107 446 108 
rect 448 107 449 108 
<< m2c >>
rect 445 102 446 103 
rect 448 102 449 103 
rect 445 107 446 108 
rect 448 107 449 108 
<< labels >>
rlabel pdiffusion 481 192 482 193  0 t = 1
rlabel pdiffusion 484 192 485 193  0 t = 2
rlabel pdiffusion 481 197 482 198  0 t = 3
rlabel pdiffusion 484 197 485 198  0 t = 4
rlabel pdiffusion 480 192 486 198 0 cell no = 223
<< m1 >>
rect 481 192 482 193 
rect 484 192 485 193 
rect 481 197 482 198 
rect 484 197 485 198 
<< m2 >>
rect 481 192 482 193 
rect 484 192 485 193 
rect 481 197 482 198 
rect 484 197 485 198 
<< m2c >>
rect 481 192 482 193 
rect 484 192 485 193 
rect 481 197 482 198 
rect 484 197 485 198 
<< labels >>
rlabel pdiffusion 427 84 428 85  0 t = 1
rlabel pdiffusion 430 84 431 85  0 t = 2
rlabel pdiffusion 427 89 428 90  0 t = 3
rlabel pdiffusion 430 89 431 90  0 t = 4
rlabel pdiffusion 426 84 432 90 0 cell no = 224
<< m1 >>
rect 427 84 428 85 
rect 430 84 431 85 
rect 427 89 428 90 
rect 430 89 431 90 
<< m2 >>
rect 427 84 428 85 
rect 430 84 431 85 
rect 427 89 428 90 
rect 430 89 431 90 
<< m2c >>
rect 427 84 428 85 
rect 430 84 431 85 
rect 427 89 428 90 
rect 430 89 431 90 
<< labels >>
rlabel pdiffusion 463 30 464 31  0 t = 1
rlabel pdiffusion 466 30 467 31  0 t = 2
rlabel pdiffusion 463 35 464 36  0 t = 3
rlabel pdiffusion 466 35 467 36  0 t = 4
rlabel pdiffusion 462 30 468 36 0 cell no = 225
<< m1 >>
rect 463 30 464 31 
rect 466 30 467 31 
rect 463 35 464 36 
rect 466 35 467 36 
<< m2 >>
rect 463 30 464 31 
rect 466 30 467 31 
rect 463 35 464 36 
rect 466 35 467 36 
<< m2c >>
rect 463 30 464 31 
rect 466 30 467 31 
rect 463 35 464 36 
rect 466 35 467 36 
<< labels >>
rlabel pdiffusion 247 84 248 85  0 t = 1
rlabel pdiffusion 250 84 251 85  0 t = 2
rlabel pdiffusion 247 89 248 90  0 t = 3
rlabel pdiffusion 250 89 251 90  0 t = 4
rlabel pdiffusion 246 84 252 90 0 cell no = 226
<< m1 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2 >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< m2c >>
rect 247 84 248 85 
rect 250 84 251 85 
rect 247 89 248 90 
rect 250 89 251 90 
<< labels >>
rlabel pdiffusion 355 210 356 211  0 t = 1
rlabel pdiffusion 358 210 359 211  0 t = 2
rlabel pdiffusion 355 215 356 216  0 t = 3
rlabel pdiffusion 358 215 359 216  0 t = 4
rlabel pdiffusion 354 210 360 216 0 cell no = 227
<< m1 >>
rect 355 210 356 211 
rect 358 210 359 211 
rect 355 215 356 216 
rect 358 215 359 216 
<< m2 >>
rect 355 210 356 211 
rect 358 210 359 211 
rect 355 215 356 216 
rect 358 215 359 216 
<< m2c >>
rect 355 210 356 211 
rect 358 210 359 211 
rect 355 215 356 216 
rect 358 215 359 216 
<< labels >>
rlabel pdiffusion 193 264 194 265  0 t = 1
rlabel pdiffusion 196 264 197 265  0 t = 2
rlabel pdiffusion 193 269 194 270  0 t = 3
rlabel pdiffusion 196 269 197 270  0 t = 4
rlabel pdiffusion 192 264 198 270 0 cell no = 228
<< m1 >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< m2 >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< m2c >>
rect 193 264 194 265 
rect 196 264 197 265 
rect 193 269 194 270 
rect 196 269 197 270 
<< labels >>
rlabel pdiffusion 481 228 482 229  0 t = 1
rlabel pdiffusion 484 228 485 229  0 t = 2
rlabel pdiffusion 481 233 482 234  0 t = 3
rlabel pdiffusion 484 233 485 234  0 t = 4
rlabel pdiffusion 480 228 486 234 0 cell no = 229
<< m1 >>
rect 481 228 482 229 
rect 484 228 485 229 
rect 481 233 482 234 
rect 484 233 485 234 
<< m2 >>
rect 481 228 482 229 
rect 484 228 485 229 
rect 481 233 482 234 
rect 484 233 485 234 
<< m2c >>
rect 481 228 482 229 
rect 484 228 485 229 
rect 481 233 482 234 
rect 484 233 485 234 
<< labels >>
rlabel pdiffusion 427 66 428 67  0 t = 1
rlabel pdiffusion 430 66 431 67  0 t = 2
rlabel pdiffusion 427 71 428 72  0 t = 3
rlabel pdiffusion 430 71 431 72  0 t = 4
rlabel pdiffusion 426 66 432 72 0 cell no = 230
<< m1 >>
rect 427 66 428 67 
rect 430 66 431 67 
rect 427 71 428 72 
rect 430 71 431 72 
<< m2 >>
rect 427 66 428 67 
rect 430 66 431 67 
rect 427 71 428 72 
rect 430 71 431 72 
<< m2c >>
rect 427 66 428 67 
rect 430 66 431 67 
rect 427 71 428 72 
rect 430 71 431 72 
<< labels >>
rlabel pdiffusion 427 30 428 31  0 t = 1
rlabel pdiffusion 430 30 431 31  0 t = 2
rlabel pdiffusion 427 35 428 36  0 t = 3
rlabel pdiffusion 430 35 431 36  0 t = 4
rlabel pdiffusion 426 30 432 36 0 cell no = 231
<< m1 >>
rect 427 30 428 31 
rect 430 30 431 31 
rect 427 35 428 36 
rect 430 35 431 36 
<< m2 >>
rect 427 30 428 31 
rect 430 30 431 31 
rect 427 35 428 36 
rect 430 35 431 36 
<< m2c >>
rect 427 30 428 31 
rect 430 30 431 31 
rect 427 35 428 36 
rect 430 35 431 36 
<< labels >>
rlabel pdiffusion 517 12 518 13  0 t = 1
rlabel pdiffusion 520 12 521 13  0 t = 2
rlabel pdiffusion 517 17 518 18  0 t = 3
rlabel pdiffusion 520 17 521 18  0 t = 4
rlabel pdiffusion 516 12 522 18 0 cell no = 232
<< m1 >>
rect 517 12 518 13 
rect 520 12 521 13 
rect 517 17 518 18 
rect 520 17 521 18 
<< m2 >>
rect 517 12 518 13 
rect 520 12 521 13 
rect 517 17 518 18 
rect 520 17 521 18 
<< m2c >>
rect 517 12 518 13 
rect 520 12 521 13 
rect 517 17 518 18 
rect 520 17 521 18 
<< labels >>
rlabel pdiffusion 67 192 68 193  0 t = 1
rlabel pdiffusion 70 192 71 193  0 t = 2
rlabel pdiffusion 67 197 68 198  0 t = 3
rlabel pdiffusion 70 197 71 198  0 t = 4
rlabel pdiffusion 66 192 72 198 0 cell no = 233
<< m1 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2 >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< m2c >>
rect 67 192 68 193 
rect 70 192 71 193 
rect 67 197 68 198 
rect 70 197 71 198 
<< labels >>
rlabel pdiffusion 13 228 14 229  0 t = 1
rlabel pdiffusion 16 228 17 229  0 t = 2
rlabel pdiffusion 13 233 14 234  0 t = 3
rlabel pdiffusion 16 233 17 234  0 t = 4
rlabel pdiffusion 12 228 18 234 0 cell no = 234
<< m1 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2 >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< m2c >>
rect 13 228 14 229 
rect 16 228 17 229 
rect 13 233 14 234 
rect 16 233 17 234 
<< labels >>
rlabel pdiffusion 121 246 122 247  0 t = 1
rlabel pdiffusion 124 246 125 247  0 t = 2
rlabel pdiffusion 121 251 122 252  0 t = 3
rlabel pdiffusion 124 251 125 252  0 t = 4
rlabel pdiffusion 120 246 126 252 0 cell no = 235
<< m1 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2 >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< m2c >>
rect 121 246 122 247 
rect 124 246 125 247 
rect 121 251 122 252 
rect 124 251 125 252 
<< labels >>
rlabel pdiffusion 175 120 176 121  0 t = 1
rlabel pdiffusion 178 120 179 121  0 t = 2
rlabel pdiffusion 175 125 176 126  0 t = 3
rlabel pdiffusion 178 125 179 126  0 t = 4
rlabel pdiffusion 174 120 180 126 0 cell no = 236
<< m1 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2 >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< m2c >>
rect 175 120 176 121 
rect 178 120 179 121 
rect 175 125 176 126 
rect 178 125 179 126 
<< labels >>
rlabel pdiffusion 31 246 32 247  0 t = 1
rlabel pdiffusion 34 246 35 247  0 t = 2
rlabel pdiffusion 31 251 32 252  0 t = 3
rlabel pdiffusion 34 251 35 252  0 t = 4
rlabel pdiffusion 30 246 36 252 0 cell no = 237
<< m1 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2 >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< m2c >>
rect 31 246 32 247 
rect 34 246 35 247 
rect 31 251 32 252 
rect 34 251 35 252 
<< labels >>
rlabel pdiffusion 49 246 50 247  0 t = 1
rlabel pdiffusion 52 246 53 247  0 t = 2
rlabel pdiffusion 49 251 50 252  0 t = 3
rlabel pdiffusion 52 251 53 252  0 t = 4
rlabel pdiffusion 48 246 54 252 0 cell no = 238
<< m1 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2 >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< m2c >>
rect 49 246 50 247 
rect 52 246 53 247 
rect 49 251 50 252 
rect 52 251 53 252 
<< labels >>
rlabel pdiffusion 157 192 158 193  0 t = 1
rlabel pdiffusion 160 192 161 193  0 t = 2
rlabel pdiffusion 157 197 158 198  0 t = 3
rlabel pdiffusion 160 197 161 198  0 t = 4
rlabel pdiffusion 156 192 162 198 0 cell no = 239
<< m1 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2 >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< m2c >>
rect 157 192 158 193 
rect 160 192 161 193 
rect 157 197 158 198 
rect 160 197 161 198 
<< labels >>
rlabel pdiffusion 49 174 50 175  0 t = 1
rlabel pdiffusion 52 174 53 175  0 t = 2
rlabel pdiffusion 49 179 50 180  0 t = 3
rlabel pdiffusion 52 179 53 180  0 t = 4
rlabel pdiffusion 48 174 54 180 0 cell no = 240
<< m1 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2 >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< m2c >>
rect 49 174 50 175 
rect 52 174 53 175 
rect 49 179 50 180 
rect 52 179 53 180 
<< labels >>
rlabel pdiffusion 49 66 50 67  0 t = 1
rlabel pdiffusion 52 66 53 67  0 t = 2
rlabel pdiffusion 49 71 50 72  0 t = 3
rlabel pdiffusion 52 71 53 72  0 t = 4
rlabel pdiffusion 48 66 54 72 0 cell no = 241
<< m1 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2 >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< m2c >>
rect 49 66 50 67 
rect 52 66 53 67 
rect 49 71 50 72 
rect 52 71 53 72 
<< labels >>
rlabel pdiffusion 193 102 194 103  0 t = 1
rlabel pdiffusion 196 102 197 103  0 t = 2
rlabel pdiffusion 193 107 194 108  0 t = 3
rlabel pdiffusion 196 107 197 108  0 t = 4
rlabel pdiffusion 192 102 198 108 0 cell no = 242
<< m1 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2 >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< m2c >>
rect 193 102 194 103 
rect 196 102 197 103 
rect 193 107 194 108 
rect 196 107 197 108 
<< labels >>
rlabel pdiffusion 355 66 356 67  0 t = 1
rlabel pdiffusion 358 66 359 67  0 t = 2
rlabel pdiffusion 355 71 356 72  0 t = 3
rlabel pdiffusion 358 71 359 72  0 t = 4
rlabel pdiffusion 354 66 360 72 0 cell no = 243
<< m1 >>
rect 355 66 356 67 
rect 358 66 359 67 
rect 355 71 356 72 
rect 358 71 359 72 
<< m2 >>
rect 355 66 356 67 
rect 358 66 359 67 
rect 355 71 356 72 
rect 358 71 359 72 
<< m2c >>
rect 355 66 356 67 
rect 358 66 359 67 
rect 355 71 356 72 
rect 358 71 359 72 
<< labels >>
rlabel pdiffusion 463 228 464 229  0 t = 1
rlabel pdiffusion 466 228 467 229  0 t = 2
rlabel pdiffusion 463 233 464 234  0 t = 3
rlabel pdiffusion 466 233 467 234  0 t = 4
rlabel pdiffusion 462 228 468 234 0 cell no = 244
<< m1 >>
rect 463 228 464 229 
rect 466 228 467 229 
rect 463 233 464 234 
rect 466 233 467 234 
<< m2 >>
rect 463 228 464 229 
rect 466 228 467 229 
rect 463 233 464 234 
rect 466 233 467 234 
<< m2c >>
rect 463 228 464 229 
rect 466 228 467 229 
rect 463 233 464 234 
rect 466 233 467 234 
<< labels >>
rlabel pdiffusion 337 30 338 31  0 t = 1
rlabel pdiffusion 340 30 341 31  0 t = 2
rlabel pdiffusion 337 35 338 36  0 t = 3
rlabel pdiffusion 340 35 341 36  0 t = 4
rlabel pdiffusion 336 30 342 36 0 cell no = 245
<< m1 >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< m2 >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< m2c >>
rect 337 30 338 31 
rect 340 30 341 31 
rect 337 35 338 36 
rect 340 35 341 36 
<< labels >>
rlabel pdiffusion 445 444 446 445  0 t = 1
rlabel pdiffusion 448 444 449 445  0 t = 2
rlabel pdiffusion 445 449 446 450  0 t = 3
rlabel pdiffusion 448 449 449 450  0 t = 4
rlabel pdiffusion 444 444 450 450 0 cell no = 246
<< m1 >>
rect 445 444 446 445 
rect 448 444 449 445 
rect 445 449 446 450 
rect 448 449 449 450 
<< m2 >>
rect 445 444 446 445 
rect 448 444 449 445 
rect 445 449 446 450 
rect 448 449 449 450 
<< m2c >>
rect 445 444 446 445 
rect 448 444 449 445 
rect 445 449 446 450 
rect 448 449 449 450 
<< labels >>
rlabel pdiffusion 355 300 356 301  0 t = 1
rlabel pdiffusion 358 300 359 301  0 t = 2
rlabel pdiffusion 355 305 356 306  0 t = 3
rlabel pdiffusion 358 305 359 306  0 t = 4
rlabel pdiffusion 354 300 360 306 0 cell no = 247
<< m1 >>
rect 355 300 356 301 
rect 358 300 359 301 
rect 355 305 356 306 
rect 358 305 359 306 
<< m2 >>
rect 355 300 356 301 
rect 358 300 359 301 
rect 355 305 356 306 
rect 358 305 359 306 
<< m2c >>
rect 355 300 356 301 
rect 358 300 359 301 
rect 355 305 356 306 
rect 358 305 359 306 
<< labels >>
rlabel pdiffusion 139 30 140 31  0 t = 1
rlabel pdiffusion 142 30 143 31  0 t = 2
rlabel pdiffusion 139 35 140 36  0 t = 3
rlabel pdiffusion 142 35 143 36  0 t = 4
rlabel pdiffusion 138 30 144 36 0 cell no = 248
<< m1 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2 >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< m2c >>
rect 139 30 140 31 
rect 142 30 143 31 
rect 139 35 140 36 
rect 142 35 143 36 
<< labels >>
rlabel pdiffusion 265 84 266 85  0 t = 1
rlabel pdiffusion 268 84 269 85  0 t = 2
rlabel pdiffusion 265 89 266 90  0 t = 3
rlabel pdiffusion 268 89 269 90  0 t = 4
rlabel pdiffusion 264 84 270 90 0 cell no = 249
<< m1 >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< m2 >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< m2c >>
rect 265 84 266 85 
rect 268 84 269 85 
rect 265 89 266 90 
rect 268 89 269 90 
<< labels >>
rlabel pdiffusion 229 84 230 85  0 t = 1
rlabel pdiffusion 232 84 233 85  0 t = 2
rlabel pdiffusion 229 89 230 90  0 t = 3
rlabel pdiffusion 232 89 233 90  0 t = 4
rlabel pdiffusion 228 84 234 90 0 cell no = 250
<< m1 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2 >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< m2c >>
rect 229 84 230 85 
rect 232 84 233 85 
rect 229 89 230 90 
rect 232 89 233 90 
<< labels >>
rlabel pdiffusion 301 30 302 31  0 t = 1
rlabel pdiffusion 304 30 305 31  0 t = 2
rlabel pdiffusion 301 35 302 36  0 t = 3
rlabel pdiffusion 304 35 305 36  0 t = 4
rlabel pdiffusion 300 30 306 36 0 cell no = 251
<< m1 >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< m2 >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< m2c >>
rect 301 30 302 31 
rect 304 30 305 31 
rect 301 35 302 36 
rect 304 35 305 36 
<< labels >>
rlabel pdiffusion 67 174 68 175  0 t = 1
rlabel pdiffusion 70 174 71 175  0 t = 2
rlabel pdiffusion 67 179 68 180  0 t = 3
rlabel pdiffusion 70 179 71 180  0 t = 4
rlabel pdiffusion 66 174 72 180 0 cell no = 252
<< m1 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2 >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< m2c >>
rect 67 174 68 175 
rect 70 174 71 175 
rect 67 179 68 180 
rect 70 179 71 180 
<< labels >>
rlabel pdiffusion 373 138 374 139  0 t = 1
rlabel pdiffusion 376 138 377 139  0 t = 2
rlabel pdiffusion 373 143 374 144  0 t = 3
rlabel pdiffusion 376 143 377 144  0 t = 4
rlabel pdiffusion 372 138 378 144 0 cell no = 253
<< m1 >>
rect 373 138 374 139 
rect 376 138 377 139 
rect 373 143 374 144 
rect 376 143 377 144 
<< m2 >>
rect 373 138 374 139 
rect 376 138 377 139 
rect 373 143 374 144 
rect 376 143 377 144 
<< m2c >>
rect 373 138 374 139 
rect 376 138 377 139 
rect 373 143 374 144 
rect 376 143 377 144 
<< labels >>
rlabel pdiffusion 499 66 500 67  0 t = 1
rlabel pdiffusion 502 66 503 67  0 t = 2
rlabel pdiffusion 499 71 500 72  0 t = 3
rlabel pdiffusion 502 71 503 72  0 t = 4
rlabel pdiffusion 498 66 504 72 0 cell no = 254
<< m1 >>
rect 499 66 500 67 
rect 502 66 503 67 
rect 499 71 500 72 
rect 502 71 503 72 
<< m2 >>
rect 499 66 500 67 
rect 502 66 503 67 
rect 499 71 500 72 
rect 502 71 503 72 
<< m2c >>
rect 499 66 500 67 
rect 502 66 503 67 
rect 499 71 500 72 
rect 502 71 503 72 
<< labels >>
rlabel pdiffusion 337 84 338 85  0 t = 1
rlabel pdiffusion 340 84 341 85  0 t = 2
rlabel pdiffusion 337 89 338 90  0 t = 3
rlabel pdiffusion 340 89 341 90  0 t = 4
rlabel pdiffusion 336 84 342 90 0 cell no = 255
<< m1 >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< m2 >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< m2c >>
rect 337 84 338 85 
rect 340 84 341 85 
rect 337 89 338 90 
rect 340 89 341 90 
<< labels >>
rlabel pdiffusion 391 210 392 211  0 t = 1
rlabel pdiffusion 394 210 395 211  0 t = 2
rlabel pdiffusion 391 215 392 216  0 t = 3
rlabel pdiffusion 394 215 395 216  0 t = 4
rlabel pdiffusion 390 210 396 216 0 cell no = 256
<< m1 >>
rect 391 210 392 211 
rect 394 210 395 211 
rect 391 215 392 216 
rect 394 215 395 216 
<< m2 >>
rect 391 210 392 211 
rect 394 210 395 211 
rect 391 215 392 216 
rect 394 215 395 216 
<< m2c >>
rect 391 210 392 211 
rect 394 210 395 211 
rect 391 215 392 216 
rect 394 215 395 216 
<< labels >>
rlabel pdiffusion 463 138 464 139  0 t = 1
rlabel pdiffusion 466 138 467 139  0 t = 2
rlabel pdiffusion 463 143 464 144  0 t = 3
rlabel pdiffusion 466 143 467 144  0 t = 4
rlabel pdiffusion 462 138 468 144 0 cell no = 257
<< m1 >>
rect 463 138 464 139 
rect 466 138 467 139 
rect 463 143 464 144 
rect 466 143 467 144 
<< m2 >>
rect 463 138 464 139 
rect 466 138 467 139 
rect 463 143 464 144 
rect 466 143 467 144 
<< m2c >>
rect 463 138 464 139 
rect 466 138 467 139 
rect 463 143 464 144 
rect 466 143 467 144 
<< labels >>
rlabel pdiffusion 481 210 482 211  0 t = 1
rlabel pdiffusion 484 210 485 211  0 t = 2
rlabel pdiffusion 481 215 482 216  0 t = 3
rlabel pdiffusion 484 215 485 216  0 t = 4
rlabel pdiffusion 480 210 486 216 0 cell no = 258
<< m1 >>
rect 481 210 482 211 
rect 484 210 485 211 
rect 481 215 482 216 
rect 484 215 485 216 
<< m2 >>
rect 481 210 482 211 
rect 484 210 485 211 
rect 481 215 482 216 
rect 484 215 485 216 
<< m2c >>
rect 481 210 482 211 
rect 484 210 485 211 
rect 481 215 482 216 
rect 484 215 485 216 
<< labels >>
rlabel pdiffusion 301 84 302 85  0 t = 1
rlabel pdiffusion 304 84 305 85  0 t = 2
rlabel pdiffusion 301 89 302 90  0 t = 3
rlabel pdiffusion 304 89 305 90  0 t = 4
rlabel pdiffusion 300 84 306 90 0 cell no = 259
<< m1 >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< m2 >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< m2c >>
rect 301 84 302 85 
rect 304 84 305 85 
rect 301 89 302 90 
rect 304 89 305 90 
<< labels >>
rlabel pdiffusion 481 156 482 157  0 t = 1
rlabel pdiffusion 484 156 485 157  0 t = 2
rlabel pdiffusion 481 161 482 162  0 t = 3
rlabel pdiffusion 484 161 485 162  0 t = 4
rlabel pdiffusion 480 156 486 162 0 cell no = 260
<< m1 >>
rect 481 156 482 157 
rect 484 156 485 157 
rect 481 161 482 162 
rect 484 161 485 162 
<< m2 >>
rect 481 156 482 157 
rect 484 156 485 157 
rect 481 161 482 162 
rect 484 161 485 162 
<< m2c >>
rect 481 156 482 157 
rect 484 156 485 157 
rect 481 161 482 162 
rect 484 161 485 162 
<< labels >>
rlabel pdiffusion 463 66 464 67  0 t = 1
rlabel pdiffusion 466 66 467 67  0 t = 2
rlabel pdiffusion 463 71 464 72  0 t = 3
rlabel pdiffusion 466 71 467 72  0 t = 4
rlabel pdiffusion 462 66 468 72 0 cell no = 261
<< m1 >>
rect 463 66 464 67 
rect 466 66 467 67 
rect 463 71 464 72 
rect 466 71 467 72 
<< m2 >>
rect 463 66 464 67 
rect 466 66 467 67 
rect 463 71 464 72 
rect 466 71 467 72 
<< m2c >>
rect 463 66 464 67 
rect 466 66 467 67 
rect 463 71 464 72 
rect 466 71 467 72 
<< labels >>
rlabel pdiffusion 427 300 428 301  0 t = 1
rlabel pdiffusion 430 300 431 301  0 t = 2
rlabel pdiffusion 427 305 428 306  0 t = 3
rlabel pdiffusion 430 305 431 306  0 t = 4
rlabel pdiffusion 426 300 432 306 0 cell no = 262
<< m1 >>
rect 427 300 428 301 
rect 430 300 431 301 
rect 427 305 428 306 
rect 430 305 431 306 
<< m2 >>
rect 427 300 428 301 
rect 430 300 431 301 
rect 427 305 428 306 
rect 430 305 431 306 
<< m2c >>
rect 427 300 428 301 
rect 430 300 431 301 
rect 427 305 428 306 
rect 430 305 431 306 
<< labels >>
rlabel pdiffusion 193 498 194 499  0 t = 1
rlabel pdiffusion 196 498 197 499  0 t = 2
rlabel pdiffusion 193 503 194 504  0 t = 3
rlabel pdiffusion 196 503 197 504  0 t = 4
rlabel pdiffusion 192 498 198 504 0 cell no = 263
<< m1 >>
rect 193 498 194 499 
rect 196 498 197 499 
rect 193 503 194 504 
rect 196 503 197 504 
<< m2 >>
rect 193 498 194 499 
rect 196 498 197 499 
rect 193 503 194 504 
rect 196 503 197 504 
<< m2c >>
rect 193 498 194 499 
rect 196 498 197 499 
rect 193 503 194 504 
rect 196 503 197 504 
<< labels >>
rlabel pdiffusion 31 336 32 337  0 t = 1
rlabel pdiffusion 34 336 35 337  0 t = 2
rlabel pdiffusion 31 341 32 342  0 t = 3
rlabel pdiffusion 34 341 35 342  0 t = 4
rlabel pdiffusion 30 336 36 342 0 cell no = 264
<< m1 >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< m2 >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< m2c >>
rect 31 336 32 337 
rect 34 336 35 337 
rect 31 341 32 342 
rect 34 341 35 342 
<< labels >>
rlabel pdiffusion 13 480 14 481  0 t = 1
rlabel pdiffusion 16 480 17 481  0 t = 2
rlabel pdiffusion 13 485 14 486  0 t = 3
rlabel pdiffusion 16 485 17 486  0 t = 4
rlabel pdiffusion 12 480 18 486 0 cell no = 265
<< m1 >>
rect 13 480 14 481 
rect 16 480 17 481 
rect 13 485 14 486 
rect 16 485 17 486 
<< m2 >>
rect 13 480 14 481 
rect 16 480 17 481 
rect 13 485 14 486 
rect 16 485 17 486 
<< m2c >>
rect 13 480 14 481 
rect 16 480 17 481 
rect 13 485 14 486 
rect 16 485 17 486 
<< labels >>
rlabel pdiffusion 103 372 104 373  0 t = 1
rlabel pdiffusion 106 372 107 373  0 t = 2
rlabel pdiffusion 103 377 104 378  0 t = 3
rlabel pdiffusion 106 377 107 378  0 t = 4
rlabel pdiffusion 102 372 108 378 0 cell no = 266
<< m1 >>
rect 103 372 104 373 
rect 106 372 107 373 
rect 103 377 104 378 
rect 106 377 107 378 
<< m2 >>
rect 103 372 104 373 
rect 106 372 107 373 
rect 103 377 104 378 
rect 106 377 107 378 
<< m2c >>
rect 103 372 104 373 
rect 106 372 107 373 
rect 103 377 104 378 
rect 106 377 107 378 
<< labels >>
rlabel pdiffusion 211 138 212 139  0 t = 1
rlabel pdiffusion 214 138 215 139  0 t = 2
rlabel pdiffusion 211 143 212 144  0 t = 3
rlabel pdiffusion 214 143 215 144  0 t = 4
rlabel pdiffusion 210 138 216 144 0 cell no = 267
<< m1 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2 >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< m2c >>
rect 211 138 212 139 
rect 214 138 215 139 
rect 211 143 212 144 
rect 214 143 215 144 
<< labels >>
rlabel pdiffusion 49 120 50 121  0 t = 1
rlabel pdiffusion 52 120 53 121  0 t = 2
rlabel pdiffusion 49 125 50 126  0 t = 3
rlabel pdiffusion 52 125 53 126  0 t = 4
rlabel pdiffusion 48 120 54 126 0 cell no = 268
<< m1 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2 >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< m2c >>
rect 49 120 50 121 
rect 52 120 53 121 
rect 49 125 50 126 
rect 52 125 53 126 
<< labels >>
rlabel pdiffusion 31 228 32 229  0 t = 1
rlabel pdiffusion 34 228 35 229  0 t = 2
rlabel pdiffusion 31 233 32 234  0 t = 3
rlabel pdiffusion 34 233 35 234  0 t = 4
rlabel pdiffusion 30 228 36 234 0 cell no = 269
<< m1 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2 >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< m2c >>
rect 31 228 32 229 
rect 34 228 35 229 
rect 31 233 32 234 
rect 34 233 35 234 
<< labels >>
rlabel pdiffusion 409 354 410 355  0 t = 1
rlabel pdiffusion 412 354 413 355  0 t = 2
rlabel pdiffusion 409 359 410 360  0 t = 3
rlabel pdiffusion 412 359 413 360  0 t = 4
rlabel pdiffusion 408 354 414 360 0 cell no = 270
<< m1 >>
rect 409 354 410 355 
rect 412 354 413 355 
rect 409 359 410 360 
rect 412 359 413 360 
<< m2 >>
rect 409 354 410 355 
rect 412 354 413 355 
rect 409 359 410 360 
rect 412 359 413 360 
<< m2c >>
rect 409 354 410 355 
rect 412 354 413 355 
rect 409 359 410 360 
rect 412 359 413 360 
<< labels >>
rlabel pdiffusion 391 246 392 247  0 t = 1
rlabel pdiffusion 394 246 395 247  0 t = 2
rlabel pdiffusion 391 251 392 252  0 t = 3
rlabel pdiffusion 394 251 395 252  0 t = 4
rlabel pdiffusion 390 246 396 252 0 cell no = 271
<< m1 >>
rect 391 246 392 247 
rect 394 246 395 247 
rect 391 251 392 252 
rect 394 251 395 252 
<< m2 >>
rect 391 246 392 247 
rect 394 246 395 247 
rect 391 251 392 252 
rect 394 251 395 252 
<< m2c >>
rect 391 246 392 247 
rect 394 246 395 247 
rect 391 251 392 252 
rect 394 251 395 252 
<< labels >>
rlabel pdiffusion 193 174 194 175  0 t = 1
rlabel pdiffusion 196 174 197 175  0 t = 2
rlabel pdiffusion 193 179 194 180  0 t = 3
rlabel pdiffusion 196 179 197 180  0 t = 4
rlabel pdiffusion 192 174 198 180 0 cell no = 272
<< m1 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2 >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< m2c >>
rect 193 174 194 175 
rect 196 174 197 175 
rect 193 179 194 180 
rect 196 179 197 180 
<< labels >>
rlabel pdiffusion 319 390 320 391  0 t = 1
rlabel pdiffusion 322 390 323 391  0 t = 2
rlabel pdiffusion 319 395 320 396  0 t = 3
rlabel pdiffusion 322 395 323 396  0 t = 4
rlabel pdiffusion 318 390 324 396 0 cell no = 273
<< m1 >>
rect 319 390 320 391 
rect 322 390 323 391 
rect 319 395 320 396 
rect 322 395 323 396 
<< m2 >>
rect 319 390 320 391 
rect 322 390 323 391 
rect 319 395 320 396 
rect 322 395 323 396 
<< m2c >>
rect 319 390 320 391 
rect 322 390 323 391 
rect 319 395 320 396 
rect 322 395 323 396 
<< labels >>
rlabel pdiffusion 67 372 68 373  0 t = 1
rlabel pdiffusion 70 372 71 373  0 t = 2
rlabel pdiffusion 67 377 68 378  0 t = 3
rlabel pdiffusion 70 377 71 378  0 t = 4
rlabel pdiffusion 66 372 72 378 0 cell no = 274
<< m1 >>
rect 67 372 68 373 
rect 70 372 71 373 
rect 67 377 68 378 
rect 70 377 71 378 
<< m2 >>
rect 67 372 68 373 
rect 70 372 71 373 
rect 67 377 68 378 
rect 70 377 71 378 
<< m2c >>
rect 67 372 68 373 
rect 70 372 71 373 
rect 67 377 68 378 
rect 70 377 71 378 
<< labels >>
rlabel pdiffusion 301 156 302 157  0 t = 1
rlabel pdiffusion 304 156 305 157  0 t = 2
rlabel pdiffusion 301 161 302 162  0 t = 3
rlabel pdiffusion 304 161 305 162  0 t = 4
rlabel pdiffusion 300 156 306 162 0 cell no = 275
<< m1 >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< m2 >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< m2c >>
rect 301 156 302 157 
rect 304 156 305 157 
rect 301 161 302 162 
rect 304 161 305 162 
<< labels >>
rlabel pdiffusion 157 84 158 85  0 t = 1
rlabel pdiffusion 160 84 161 85  0 t = 2
rlabel pdiffusion 157 89 158 90  0 t = 3
rlabel pdiffusion 160 89 161 90  0 t = 4
rlabel pdiffusion 156 84 162 90 0 cell no = 276
<< m1 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2 >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< m2c >>
rect 157 84 158 85 
rect 160 84 161 85 
rect 157 89 158 90 
rect 160 89 161 90 
<< labels >>
rlabel pdiffusion 247 210 248 211  0 t = 1
rlabel pdiffusion 250 210 251 211  0 t = 2
rlabel pdiffusion 247 215 248 216  0 t = 3
rlabel pdiffusion 250 215 251 216  0 t = 4
rlabel pdiffusion 246 210 252 216 0 cell no = 277
<< m1 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2 >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< m2c >>
rect 247 210 248 211 
rect 250 210 251 211 
rect 247 215 248 216 
rect 250 215 251 216 
<< labels >>
rlabel pdiffusion 337 336 338 337  0 t = 1
rlabel pdiffusion 340 336 341 337  0 t = 2
rlabel pdiffusion 337 341 338 342  0 t = 3
rlabel pdiffusion 340 341 341 342  0 t = 4
rlabel pdiffusion 336 336 342 342 0 cell no = 278
<< m1 >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< m2 >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< m2c >>
rect 337 336 338 337 
rect 340 336 341 337 
rect 337 341 338 342 
rect 340 341 341 342 
<< labels >>
rlabel pdiffusion 319 66 320 67  0 t = 1
rlabel pdiffusion 322 66 323 67  0 t = 2
rlabel pdiffusion 319 71 320 72  0 t = 3
rlabel pdiffusion 322 71 323 72  0 t = 4
rlabel pdiffusion 318 66 324 72 0 cell no = 279
<< m1 >>
rect 319 66 320 67 
rect 322 66 323 67 
rect 319 71 320 72 
rect 322 71 323 72 
<< m2 >>
rect 319 66 320 67 
rect 322 66 323 67 
rect 319 71 320 72 
rect 322 71 323 72 
<< m2c >>
rect 319 66 320 67 
rect 322 66 323 67 
rect 319 71 320 72 
rect 322 71 323 72 
<< labels >>
rlabel pdiffusion 445 354 446 355  0 t = 1
rlabel pdiffusion 448 354 449 355  0 t = 2
rlabel pdiffusion 445 359 446 360  0 t = 3
rlabel pdiffusion 448 359 449 360  0 t = 4
rlabel pdiffusion 444 354 450 360 0 cell no = 280
<< m1 >>
rect 445 354 446 355 
rect 448 354 449 355 
rect 445 359 446 360 
rect 448 359 449 360 
<< m2 >>
rect 445 354 446 355 
rect 448 354 449 355 
rect 445 359 446 360 
rect 448 359 449 360 
<< m2c >>
rect 445 354 446 355 
rect 448 354 449 355 
rect 445 359 446 360 
rect 448 359 449 360 
<< labels >>
rlabel pdiffusion 463 84 464 85  0 t = 1
rlabel pdiffusion 466 84 467 85  0 t = 2
rlabel pdiffusion 463 89 464 90  0 t = 3
rlabel pdiffusion 466 89 467 90  0 t = 4
rlabel pdiffusion 462 84 468 90 0 cell no = 281
<< m1 >>
rect 463 84 464 85 
rect 466 84 467 85 
rect 463 89 464 90 
rect 466 89 467 90 
<< m2 >>
rect 463 84 464 85 
rect 466 84 467 85 
rect 463 89 464 90 
rect 466 89 467 90 
<< m2c >>
rect 463 84 464 85 
rect 466 84 467 85 
rect 463 89 464 90 
rect 466 89 467 90 
<< labels >>
rlabel pdiffusion 283 264 284 265  0 t = 1
rlabel pdiffusion 286 264 287 265  0 t = 2
rlabel pdiffusion 283 269 284 270  0 t = 3
rlabel pdiffusion 286 269 287 270  0 t = 4
rlabel pdiffusion 282 264 288 270 0 cell no = 282
<< m1 >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< m2 >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< m2c >>
rect 283 264 284 265 
rect 286 264 287 265 
rect 283 269 284 270 
rect 286 269 287 270 
<< labels >>
rlabel pdiffusion 319 174 320 175  0 t = 1
rlabel pdiffusion 322 174 323 175  0 t = 2
rlabel pdiffusion 319 179 320 180  0 t = 3
rlabel pdiffusion 322 179 323 180  0 t = 4
rlabel pdiffusion 318 174 324 180 0 cell no = 283
<< m1 >>
rect 319 174 320 175 
rect 322 174 323 175 
rect 319 179 320 180 
rect 322 179 323 180 
<< m2 >>
rect 319 174 320 175 
rect 322 174 323 175 
rect 319 179 320 180 
rect 322 179 323 180 
<< m2c >>
rect 319 174 320 175 
rect 322 174 323 175 
rect 319 179 320 180 
rect 322 179 323 180 
<< labels >>
rlabel pdiffusion 319 156 320 157  0 t = 1
rlabel pdiffusion 322 156 323 157  0 t = 2
rlabel pdiffusion 319 161 320 162  0 t = 3
rlabel pdiffusion 322 161 323 162  0 t = 4
rlabel pdiffusion 318 156 324 162 0 cell no = 284
<< m1 >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< m2 >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< m2c >>
rect 319 156 320 157 
rect 322 156 323 157 
rect 319 161 320 162 
rect 322 161 323 162 
<< labels >>
rlabel pdiffusion 499 174 500 175  0 t = 1
rlabel pdiffusion 502 174 503 175  0 t = 2
rlabel pdiffusion 499 179 500 180  0 t = 3
rlabel pdiffusion 502 179 503 180  0 t = 4
rlabel pdiffusion 498 174 504 180 0 cell no = 285
<< m1 >>
rect 499 174 500 175 
rect 502 174 503 175 
rect 499 179 500 180 
rect 502 179 503 180 
<< m2 >>
rect 499 174 500 175 
rect 502 174 503 175 
rect 499 179 500 180 
rect 502 179 503 180 
<< m2c >>
rect 499 174 500 175 
rect 502 174 503 175 
rect 499 179 500 180 
rect 502 179 503 180 
<< labels >>
rlabel pdiffusion 139 336 140 337  0 t = 1
rlabel pdiffusion 142 336 143 337  0 t = 2
rlabel pdiffusion 139 341 140 342  0 t = 3
rlabel pdiffusion 142 341 143 342  0 t = 4
rlabel pdiffusion 138 336 144 342 0 cell no = 286
<< m1 >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< m2 >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< m2c >>
rect 139 336 140 337 
rect 142 336 143 337 
rect 139 341 140 342 
rect 142 341 143 342 
<< labels >>
rlabel pdiffusion 409 174 410 175  0 t = 1
rlabel pdiffusion 412 174 413 175  0 t = 2
rlabel pdiffusion 409 179 410 180  0 t = 3
rlabel pdiffusion 412 179 413 180  0 t = 4
rlabel pdiffusion 408 174 414 180 0 cell no = 287
<< m1 >>
rect 409 174 410 175 
rect 412 174 413 175 
rect 409 179 410 180 
rect 412 179 413 180 
<< m2 >>
rect 409 174 410 175 
rect 412 174 413 175 
rect 409 179 410 180 
rect 412 179 413 180 
<< m2c >>
rect 409 174 410 175 
rect 412 174 413 175 
rect 409 179 410 180 
rect 412 179 413 180 
<< labels >>
rlabel pdiffusion 517 138 518 139  0 t = 1
rlabel pdiffusion 520 138 521 139  0 t = 2
rlabel pdiffusion 517 143 518 144  0 t = 3
rlabel pdiffusion 520 143 521 144  0 t = 4
rlabel pdiffusion 516 138 522 144 0 cell no = 288
<< m1 >>
rect 517 138 518 139 
rect 520 138 521 139 
rect 517 143 518 144 
rect 520 143 521 144 
<< m2 >>
rect 517 138 518 139 
rect 520 138 521 139 
rect 517 143 518 144 
rect 520 143 521 144 
<< m2c >>
rect 517 138 518 139 
rect 520 138 521 139 
rect 517 143 518 144 
rect 520 143 521 144 
<< labels >>
rlabel pdiffusion 175 264 176 265  0 t = 1
rlabel pdiffusion 178 264 179 265  0 t = 2
rlabel pdiffusion 175 269 176 270  0 t = 3
rlabel pdiffusion 178 269 179 270  0 t = 4
rlabel pdiffusion 174 264 180 270 0 cell no = 289
<< m1 >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< m2 >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< m2c >>
rect 175 264 176 265 
rect 178 264 179 265 
rect 175 269 176 270 
rect 178 269 179 270 
<< labels >>
rlabel pdiffusion 409 210 410 211  0 t = 1
rlabel pdiffusion 412 210 413 211  0 t = 2
rlabel pdiffusion 409 215 410 216  0 t = 3
rlabel pdiffusion 412 215 413 216  0 t = 4
rlabel pdiffusion 408 210 414 216 0 cell no = 290
<< m1 >>
rect 409 210 410 211 
rect 412 210 413 211 
rect 409 215 410 216 
rect 412 215 413 216 
<< m2 >>
rect 409 210 410 211 
rect 412 210 413 211 
rect 409 215 410 216 
rect 412 215 413 216 
<< m2c >>
rect 409 210 410 211 
rect 412 210 413 211 
rect 409 215 410 216 
rect 412 215 413 216 
<< labels >>
rlabel pdiffusion 103 282 104 283  0 t = 1
rlabel pdiffusion 106 282 107 283  0 t = 2
rlabel pdiffusion 103 287 104 288  0 t = 3
rlabel pdiffusion 106 287 107 288  0 t = 4
rlabel pdiffusion 102 282 108 288 0 cell no = 291
<< m1 >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< m2 >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< m2c >>
rect 103 282 104 283 
rect 106 282 107 283 
rect 103 287 104 288 
rect 106 287 107 288 
<< labels >>
rlabel pdiffusion 31 120 32 121  0 t = 1
rlabel pdiffusion 34 120 35 121  0 t = 2
rlabel pdiffusion 31 125 32 126  0 t = 3
rlabel pdiffusion 34 125 35 126  0 t = 4
rlabel pdiffusion 30 120 36 126 0 cell no = 292
<< m1 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2 >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< m2c >>
rect 31 120 32 121 
rect 34 120 35 121 
rect 31 125 32 126 
rect 34 125 35 126 
<< labels >>
rlabel pdiffusion 139 84 140 85  0 t = 1
rlabel pdiffusion 142 84 143 85  0 t = 2
rlabel pdiffusion 139 89 140 90  0 t = 3
rlabel pdiffusion 142 89 143 90  0 t = 4
rlabel pdiffusion 138 84 144 90 0 cell no = 293
<< m1 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2 >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< m2c >>
rect 139 84 140 85 
rect 142 84 143 85 
rect 139 89 140 90 
rect 142 89 143 90 
<< labels >>
rlabel pdiffusion 49 156 50 157  0 t = 1
rlabel pdiffusion 52 156 53 157  0 t = 2
rlabel pdiffusion 49 161 50 162  0 t = 3
rlabel pdiffusion 52 161 53 162  0 t = 4
rlabel pdiffusion 48 156 54 162 0 cell no = 294
<< m1 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2 >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< m2c >>
rect 49 156 50 157 
rect 52 156 53 157 
rect 49 161 50 162 
rect 52 161 53 162 
<< labels >>
rlabel pdiffusion 49 84 50 85  0 t = 1
rlabel pdiffusion 52 84 53 85  0 t = 2
rlabel pdiffusion 49 89 50 90  0 t = 3
rlabel pdiffusion 52 89 53 90  0 t = 4
rlabel pdiffusion 48 84 54 90 0 cell no = 295
<< m1 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2 >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< m2c >>
rect 49 84 50 85 
rect 52 84 53 85 
rect 49 89 50 90 
rect 52 89 53 90 
<< labels >>
rlabel pdiffusion 31 138 32 139  0 t = 1
rlabel pdiffusion 34 138 35 139  0 t = 2
rlabel pdiffusion 31 143 32 144  0 t = 3
rlabel pdiffusion 34 143 35 144  0 t = 4
rlabel pdiffusion 30 138 36 144 0 cell no = 296
<< m1 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2 >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< m2c >>
rect 31 138 32 139 
rect 34 138 35 139 
rect 31 143 32 144 
rect 34 143 35 144 
<< labels >>
rlabel pdiffusion 67 246 68 247  0 t = 1
rlabel pdiffusion 70 246 71 247  0 t = 2
rlabel pdiffusion 67 251 68 252  0 t = 3
rlabel pdiffusion 70 251 71 252  0 t = 4
rlabel pdiffusion 66 246 72 252 0 cell no = 297
<< m1 >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< m2 >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< m2c >>
rect 67 246 68 247 
rect 70 246 71 247 
rect 67 251 68 252 
rect 70 251 71 252 
<< labels >>
rlabel pdiffusion 67 426 68 427  0 t = 1
rlabel pdiffusion 70 426 71 427  0 t = 2
rlabel pdiffusion 67 431 68 432  0 t = 3
rlabel pdiffusion 70 431 71 432  0 t = 4
rlabel pdiffusion 66 426 72 432 0 cell no = 298
<< m1 >>
rect 67 426 68 427 
rect 70 426 71 427 
rect 67 431 68 432 
rect 70 431 71 432 
<< m2 >>
rect 67 426 68 427 
rect 70 426 71 427 
rect 67 431 68 432 
rect 70 431 71 432 
<< m2c >>
rect 67 426 68 427 
rect 70 426 71 427 
rect 67 431 68 432 
rect 70 431 71 432 
<< labels >>
rlabel pdiffusion 175 462 176 463  0 t = 1
rlabel pdiffusion 178 462 179 463  0 t = 2
rlabel pdiffusion 175 467 176 468  0 t = 3
rlabel pdiffusion 178 467 179 468  0 t = 4
rlabel pdiffusion 174 462 180 468 0 cell no = 299
<< m1 >>
rect 175 462 176 463 
rect 178 462 179 463 
rect 175 467 176 468 
rect 178 467 179 468 
<< m2 >>
rect 175 462 176 463 
rect 178 462 179 463 
rect 175 467 176 468 
rect 178 467 179 468 
<< m2c >>
rect 175 462 176 463 
rect 178 462 179 463 
rect 175 467 176 468 
rect 178 467 179 468 
<< labels >>
rlabel pdiffusion 301 246 302 247  0 t = 1
rlabel pdiffusion 304 246 305 247  0 t = 2
rlabel pdiffusion 301 251 302 252  0 t = 3
rlabel pdiffusion 304 251 305 252  0 t = 4
rlabel pdiffusion 300 246 306 252 0 cell no = 300
<< m1 >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< m2 >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< m2c >>
rect 301 246 302 247 
rect 304 246 305 247 
rect 301 251 302 252 
rect 304 251 305 252 
<< labels >>
rlabel pdiffusion 157 138 158 139  0 t = 1
rlabel pdiffusion 160 138 161 139  0 t = 2
rlabel pdiffusion 157 143 158 144  0 t = 3
rlabel pdiffusion 160 143 161 144  0 t = 4
rlabel pdiffusion 156 138 162 144 0 cell no = 301
<< m1 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2 >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< m2c >>
rect 157 138 158 139 
rect 160 138 161 139 
rect 157 143 158 144 
rect 160 143 161 144 
<< labels >>
rlabel pdiffusion 139 138 140 139  0 t = 1
rlabel pdiffusion 142 138 143 139  0 t = 2
rlabel pdiffusion 139 143 140 144  0 t = 3
rlabel pdiffusion 142 143 143 144  0 t = 4
rlabel pdiffusion 138 138 144 144 0 cell no = 302
<< m1 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2 >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< m2c >>
rect 139 138 140 139 
rect 142 138 143 139 
rect 139 143 140 144 
rect 142 143 143 144 
<< labels >>
rlabel pdiffusion 355 48 356 49  0 t = 1
rlabel pdiffusion 358 48 359 49  0 t = 2
rlabel pdiffusion 355 53 356 54  0 t = 3
rlabel pdiffusion 358 53 359 54  0 t = 4
rlabel pdiffusion 354 48 360 54 0 cell no = 303
<< m1 >>
rect 355 48 356 49 
rect 358 48 359 49 
rect 355 53 356 54 
rect 358 53 359 54 
<< m2 >>
rect 355 48 356 49 
rect 358 48 359 49 
rect 355 53 356 54 
rect 358 53 359 54 
<< m2c >>
rect 355 48 356 49 
rect 358 48 359 49 
rect 355 53 356 54 
rect 358 53 359 54 
<< labels >>
rlabel pdiffusion 193 228 194 229  0 t = 1
rlabel pdiffusion 196 228 197 229  0 t = 2
rlabel pdiffusion 193 233 194 234  0 t = 3
rlabel pdiffusion 196 233 197 234  0 t = 4
rlabel pdiffusion 192 228 198 234 0 cell no = 304
<< m1 >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< m2 >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< m2c >>
rect 193 228 194 229 
rect 196 228 197 229 
rect 193 233 194 234 
rect 196 233 197 234 
<< labels >>
rlabel pdiffusion 85 426 86 427  0 t = 1
rlabel pdiffusion 88 426 89 427  0 t = 2
rlabel pdiffusion 85 431 86 432  0 t = 3
rlabel pdiffusion 88 431 89 432  0 t = 4
rlabel pdiffusion 84 426 90 432 0 cell no = 305
<< m1 >>
rect 85 426 86 427 
rect 88 426 89 427 
rect 85 431 86 432 
rect 88 431 89 432 
<< m2 >>
rect 85 426 86 427 
rect 88 426 89 427 
rect 85 431 86 432 
rect 88 431 89 432 
<< m2c >>
rect 85 426 86 427 
rect 88 426 89 427 
rect 85 431 86 432 
rect 88 431 89 432 
<< labels >>
rlabel pdiffusion 265 156 266 157  0 t = 1
rlabel pdiffusion 268 156 269 157  0 t = 2
rlabel pdiffusion 265 161 266 162  0 t = 3
rlabel pdiffusion 268 161 269 162  0 t = 4
rlabel pdiffusion 264 156 270 162 0 cell no = 306
<< m1 >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< m2 >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< m2c >>
rect 265 156 266 157 
rect 268 156 269 157 
rect 265 161 266 162 
rect 268 161 269 162 
<< labels >>
rlabel pdiffusion 391 66 392 67  0 t = 1
rlabel pdiffusion 394 66 395 67  0 t = 2
rlabel pdiffusion 391 71 392 72  0 t = 3
rlabel pdiffusion 394 71 395 72  0 t = 4
rlabel pdiffusion 390 66 396 72 0 cell no = 307
<< m1 >>
rect 391 66 392 67 
rect 394 66 395 67 
rect 391 71 392 72 
rect 394 71 395 72 
<< m2 >>
rect 391 66 392 67 
rect 394 66 395 67 
rect 391 71 392 72 
rect 394 71 395 72 
<< m2c >>
rect 391 66 392 67 
rect 394 66 395 67 
rect 391 71 392 72 
rect 394 71 395 72 
<< labels >>
rlabel pdiffusion 319 228 320 229  0 t = 1
rlabel pdiffusion 322 228 323 229  0 t = 2
rlabel pdiffusion 319 233 320 234  0 t = 3
rlabel pdiffusion 322 233 323 234  0 t = 4
rlabel pdiffusion 318 228 324 234 0 cell no = 308
<< m1 >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< m2 >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< m2c >>
rect 319 228 320 229 
rect 322 228 323 229 
rect 319 233 320 234 
rect 322 233 323 234 
<< labels >>
rlabel pdiffusion 229 372 230 373  0 t = 1
rlabel pdiffusion 232 372 233 373  0 t = 2
rlabel pdiffusion 229 377 230 378  0 t = 3
rlabel pdiffusion 232 377 233 378  0 t = 4
rlabel pdiffusion 228 372 234 378 0 cell no = 309
<< m1 >>
rect 229 372 230 373 
rect 232 372 233 373 
rect 229 377 230 378 
rect 232 377 233 378 
<< m2 >>
rect 229 372 230 373 
rect 232 372 233 373 
rect 229 377 230 378 
rect 232 377 233 378 
<< m2c >>
rect 229 372 230 373 
rect 232 372 233 373 
rect 229 377 230 378 
rect 232 377 233 378 
<< labels >>
rlabel pdiffusion 13 12 14 13  0 t = 1
rlabel pdiffusion 16 12 17 13  0 t = 2
rlabel pdiffusion 13 17 14 18  0 t = 3
rlabel pdiffusion 16 17 17 18  0 t = 4
rlabel pdiffusion 12 12 18 18 0 cell no = 310
<< m1 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2 >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< m2c >>
rect 13 12 14 13 
rect 16 12 17 13 
rect 13 17 14 18 
rect 16 17 17 18 
<< labels >>
rlabel pdiffusion 337 426 338 427  0 t = 1
rlabel pdiffusion 340 426 341 427  0 t = 2
rlabel pdiffusion 337 431 338 432  0 t = 3
rlabel pdiffusion 340 431 341 432  0 t = 4
rlabel pdiffusion 336 426 342 432 0 cell no = 311
<< m1 >>
rect 337 426 338 427 
rect 340 426 341 427 
rect 337 431 338 432 
rect 340 431 341 432 
<< m2 >>
rect 337 426 338 427 
rect 340 426 341 427 
rect 337 431 338 432 
rect 340 431 341 432 
<< m2c >>
rect 337 426 338 427 
rect 340 426 341 427 
rect 337 431 338 432 
rect 340 431 341 432 
<< labels >>
rlabel pdiffusion 409 228 410 229  0 t = 1
rlabel pdiffusion 412 228 413 229  0 t = 2
rlabel pdiffusion 409 233 410 234  0 t = 3
rlabel pdiffusion 412 233 413 234  0 t = 4
rlabel pdiffusion 408 228 414 234 0 cell no = 312
<< m1 >>
rect 409 228 410 229 
rect 412 228 413 229 
rect 409 233 410 234 
rect 412 233 413 234 
<< m2 >>
rect 409 228 410 229 
rect 412 228 413 229 
rect 409 233 410 234 
rect 412 233 413 234 
<< m2c >>
rect 409 228 410 229 
rect 412 228 413 229 
rect 409 233 410 234 
rect 412 233 413 234 
<< labels >>
rlabel pdiffusion 481 336 482 337  0 t = 1
rlabel pdiffusion 484 336 485 337  0 t = 2
rlabel pdiffusion 481 341 482 342  0 t = 3
rlabel pdiffusion 484 341 485 342  0 t = 4
rlabel pdiffusion 480 336 486 342 0 cell no = 313
<< m1 >>
rect 481 336 482 337 
rect 484 336 485 337 
rect 481 341 482 342 
rect 484 341 485 342 
<< m2 >>
rect 481 336 482 337 
rect 484 336 485 337 
rect 481 341 482 342 
rect 484 341 485 342 
<< m2c >>
rect 481 336 482 337 
rect 484 336 485 337 
rect 481 341 482 342 
rect 484 341 485 342 
<< labels >>
rlabel pdiffusion 409 12 410 13  0 t = 1
rlabel pdiffusion 412 12 413 13  0 t = 2
rlabel pdiffusion 409 17 410 18  0 t = 3
rlabel pdiffusion 412 17 413 18  0 t = 4
rlabel pdiffusion 408 12 414 18 0 cell no = 314
<< m1 >>
rect 409 12 410 13 
rect 412 12 413 13 
rect 409 17 410 18 
rect 412 17 413 18 
<< m2 >>
rect 409 12 410 13 
rect 412 12 413 13 
rect 409 17 410 18 
rect 412 17 413 18 
<< m2c >>
rect 409 12 410 13 
rect 412 12 413 13 
rect 409 17 410 18 
rect 412 17 413 18 
<< labels >>
rlabel pdiffusion 247 102 248 103  0 t = 1
rlabel pdiffusion 250 102 251 103  0 t = 2
rlabel pdiffusion 247 107 248 108  0 t = 3
rlabel pdiffusion 250 107 251 108  0 t = 4
rlabel pdiffusion 246 102 252 108 0 cell no = 315
<< m1 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2 >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< m2c >>
rect 247 102 248 103 
rect 250 102 251 103 
rect 247 107 248 108 
rect 250 107 251 108 
<< labels >>
rlabel pdiffusion 427 228 428 229  0 t = 1
rlabel pdiffusion 430 228 431 229  0 t = 2
rlabel pdiffusion 427 233 428 234  0 t = 3
rlabel pdiffusion 430 233 431 234  0 t = 4
rlabel pdiffusion 426 228 432 234 0 cell no = 316
<< m1 >>
rect 427 228 428 229 
rect 430 228 431 229 
rect 427 233 428 234 
rect 430 233 431 234 
<< m2 >>
rect 427 228 428 229 
rect 430 228 431 229 
rect 427 233 428 234 
rect 430 233 431 234 
<< m2c >>
rect 427 228 428 229 
rect 430 228 431 229 
rect 427 233 428 234 
rect 430 233 431 234 
<< labels >>
rlabel pdiffusion 391 138 392 139  0 t = 1
rlabel pdiffusion 394 138 395 139  0 t = 2
rlabel pdiffusion 391 143 392 144  0 t = 3
rlabel pdiffusion 394 143 395 144  0 t = 4
rlabel pdiffusion 390 138 396 144 0 cell no = 317
<< m1 >>
rect 391 138 392 139 
rect 394 138 395 139 
rect 391 143 392 144 
rect 394 143 395 144 
<< m2 >>
rect 391 138 392 139 
rect 394 138 395 139 
rect 391 143 392 144 
rect 394 143 395 144 
<< m2c >>
rect 391 138 392 139 
rect 394 138 395 139 
rect 391 143 392 144 
rect 394 143 395 144 
<< labels >>
rlabel pdiffusion 517 192 518 193  0 t = 1
rlabel pdiffusion 520 192 521 193  0 t = 2
rlabel pdiffusion 517 197 518 198  0 t = 3
rlabel pdiffusion 520 197 521 198  0 t = 4
rlabel pdiffusion 516 192 522 198 0 cell no = 318
<< m1 >>
rect 517 192 518 193 
rect 520 192 521 193 
rect 517 197 518 198 
rect 520 197 521 198 
<< m2 >>
rect 517 192 518 193 
rect 520 192 521 193 
rect 517 197 518 198 
rect 520 197 521 198 
<< m2c >>
rect 517 192 518 193 
rect 520 192 521 193 
rect 517 197 518 198 
rect 520 197 521 198 
<< labels >>
rlabel pdiffusion 499 120 500 121  0 t = 1
rlabel pdiffusion 502 120 503 121  0 t = 2
rlabel pdiffusion 499 125 500 126  0 t = 3
rlabel pdiffusion 502 125 503 126  0 t = 4
rlabel pdiffusion 498 120 504 126 0 cell no = 319
<< m1 >>
rect 499 120 500 121 
rect 502 120 503 121 
rect 499 125 500 126 
rect 502 125 503 126 
<< m2 >>
rect 499 120 500 121 
rect 502 120 503 121 
rect 499 125 500 126 
rect 502 125 503 126 
<< m2c >>
rect 499 120 500 121 
rect 502 120 503 121 
rect 499 125 500 126 
rect 502 125 503 126 
<< labels >>
rlabel pdiffusion 13 156 14 157  0 t = 1
rlabel pdiffusion 16 156 17 157  0 t = 2
rlabel pdiffusion 13 161 14 162  0 t = 3
rlabel pdiffusion 16 161 17 162  0 t = 4
rlabel pdiffusion 12 156 18 162 0 cell no = 320
<< m1 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2 >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< m2c >>
rect 13 156 14 157 
rect 16 156 17 157 
rect 13 161 14 162 
rect 16 161 17 162 
<< labels >>
rlabel pdiffusion 139 66 140 67  0 t = 1
rlabel pdiffusion 142 66 143 67  0 t = 2
rlabel pdiffusion 139 71 140 72  0 t = 3
rlabel pdiffusion 142 71 143 72  0 t = 4
rlabel pdiffusion 138 66 144 72 0 cell no = 321
<< m1 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2 >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< m2c >>
rect 139 66 140 67 
rect 142 66 143 67 
rect 139 71 140 72 
rect 142 71 143 72 
<< labels >>
rlabel pdiffusion 139 174 140 175  0 t = 1
rlabel pdiffusion 142 174 143 175  0 t = 2
rlabel pdiffusion 139 179 140 180  0 t = 3
rlabel pdiffusion 142 179 143 180  0 t = 4
rlabel pdiffusion 138 174 144 180 0 cell no = 322
<< m1 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2 >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< m2c >>
rect 139 174 140 175 
rect 142 174 143 175 
rect 139 179 140 180 
rect 142 179 143 180 
<< labels >>
rlabel pdiffusion 319 264 320 265  0 t = 1
rlabel pdiffusion 322 264 323 265  0 t = 2
rlabel pdiffusion 319 269 320 270  0 t = 3
rlabel pdiffusion 322 269 323 270  0 t = 4
rlabel pdiffusion 318 264 324 270 0 cell no = 323
<< m1 >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< m2 >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< m2c >>
rect 319 264 320 265 
rect 322 264 323 265 
rect 319 269 320 270 
rect 322 269 323 270 
<< labels >>
rlabel pdiffusion 67 300 68 301  0 t = 1
rlabel pdiffusion 70 300 71 301  0 t = 2
rlabel pdiffusion 67 305 68 306  0 t = 3
rlabel pdiffusion 70 305 71 306  0 t = 4
rlabel pdiffusion 66 300 72 306 0 cell no = 324
<< m1 >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< m2 >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< m2c >>
rect 67 300 68 301 
rect 70 300 71 301 
rect 67 305 68 306 
rect 70 305 71 306 
<< labels >>
rlabel pdiffusion 409 498 410 499  0 t = 1
rlabel pdiffusion 412 498 413 499  0 t = 2
rlabel pdiffusion 409 503 410 504  0 t = 3
rlabel pdiffusion 412 503 413 504  0 t = 4
rlabel pdiffusion 408 498 414 504 0 cell no = 325
<< m1 >>
rect 409 498 410 499 
rect 412 498 413 499 
rect 409 503 410 504 
rect 412 503 413 504 
<< m2 >>
rect 409 498 410 499 
rect 412 498 413 499 
rect 409 503 410 504 
rect 412 503 413 504 
<< m2c >>
rect 409 498 410 499 
rect 412 498 413 499 
rect 409 503 410 504 
rect 412 503 413 504 
<< labels >>
rlabel pdiffusion 85 300 86 301  0 t = 1
rlabel pdiffusion 88 300 89 301  0 t = 2
rlabel pdiffusion 85 305 86 306  0 t = 3
rlabel pdiffusion 88 305 89 306  0 t = 4
rlabel pdiffusion 84 300 90 306 0 cell no = 326
<< m1 >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< m2 >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< m2c >>
rect 85 300 86 301 
rect 88 300 89 301 
rect 85 305 86 306 
rect 88 305 89 306 
<< labels >>
rlabel pdiffusion 229 210 230 211  0 t = 1
rlabel pdiffusion 232 210 233 211  0 t = 2
rlabel pdiffusion 229 215 230 216  0 t = 3
rlabel pdiffusion 232 215 233 216  0 t = 4
rlabel pdiffusion 228 210 234 216 0 cell no = 327
<< m1 >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< m2 >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< m2c >>
rect 229 210 230 211 
rect 232 210 233 211 
rect 229 215 230 216 
rect 232 215 233 216 
<< labels >>
rlabel pdiffusion 121 264 122 265  0 t = 1
rlabel pdiffusion 124 264 125 265  0 t = 2
rlabel pdiffusion 121 269 122 270  0 t = 3
rlabel pdiffusion 124 269 125 270  0 t = 4
rlabel pdiffusion 120 264 126 270 0 cell no = 328
<< m1 >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< m2 >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< m2c >>
rect 121 264 122 265 
rect 124 264 125 265 
rect 121 269 122 270 
rect 124 269 125 270 
<< labels >>
rlabel pdiffusion 319 444 320 445  0 t = 1
rlabel pdiffusion 322 444 323 445  0 t = 2
rlabel pdiffusion 319 449 320 450  0 t = 3
rlabel pdiffusion 322 449 323 450  0 t = 4
rlabel pdiffusion 318 444 324 450 0 cell no = 329
<< m1 >>
rect 319 444 320 445 
rect 322 444 323 445 
rect 319 449 320 450 
rect 322 449 323 450 
<< m2 >>
rect 319 444 320 445 
rect 322 444 323 445 
rect 319 449 320 450 
rect 322 449 323 450 
<< m2c >>
rect 319 444 320 445 
rect 322 444 323 445 
rect 319 449 320 450 
rect 322 449 323 450 
<< labels >>
rlabel pdiffusion 103 174 104 175  0 t = 1
rlabel pdiffusion 106 174 107 175  0 t = 2
rlabel pdiffusion 103 179 104 180  0 t = 3
rlabel pdiffusion 106 179 107 180  0 t = 4
rlabel pdiffusion 102 174 108 180 0 cell no = 330
<< m1 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2 >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< m2c >>
rect 103 174 104 175 
rect 106 174 107 175 
rect 103 179 104 180 
rect 106 179 107 180 
<< labels >>
rlabel pdiffusion 517 84 518 85  0 t = 1
rlabel pdiffusion 520 84 521 85  0 t = 2
rlabel pdiffusion 517 89 518 90  0 t = 3
rlabel pdiffusion 520 89 521 90  0 t = 4
rlabel pdiffusion 516 84 522 90 0 cell no = 331
<< m1 >>
rect 517 84 518 85 
rect 520 84 521 85 
rect 517 89 518 90 
rect 520 89 521 90 
<< m2 >>
rect 517 84 518 85 
rect 520 84 521 85 
rect 517 89 518 90 
rect 520 89 521 90 
<< m2c >>
rect 517 84 518 85 
rect 520 84 521 85 
rect 517 89 518 90 
rect 520 89 521 90 
<< labels >>
rlabel pdiffusion 373 102 374 103  0 t = 1
rlabel pdiffusion 376 102 377 103  0 t = 2
rlabel pdiffusion 373 107 374 108  0 t = 3
rlabel pdiffusion 376 107 377 108  0 t = 4
rlabel pdiffusion 372 102 378 108 0 cell no = 332
<< m1 >>
rect 373 102 374 103 
rect 376 102 377 103 
rect 373 107 374 108 
rect 376 107 377 108 
<< m2 >>
rect 373 102 374 103 
rect 376 102 377 103 
rect 373 107 374 108 
rect 376 107 377 108 
<< m2c >>
rect 373 102 374 103 
rect 376 102 377 103 
rect 373 107 374 108 
rect 376 107 377 108 
<< labels >>
rlabel pdiffusion 247 480 248 481  0 t = 1
rlabel pdiffusion 250 480 251 481  0 t = 2
rlabel pdiffusion 247 485 248 486  0 t = 3
rlabel pdiffusion 250 485 251 486  0 t = 4
rlabel pdiffusion 246 480 252 486 0 cell no = 333
<< m1 >>
rect 247 480 248 481 
rect 250 480 251 481 
rect 247 485 248 486 
rect 250 485 251 486 
<< m2 >>
rect 247 480 248 481 
rect 250 480 251 481 
rect 247 485 248 486 
rect 250 485 251 486 
<< m2c >>
rect 247 480 248 481 
rect 250 480 251 481 
rect 247 485 248 486 
rect 250 485 251 486 
<< labels >>
rlabel pdiffusion 391 102 392 103  0 t = 1
rlabel pdiffusion 394 102 395 103  0 t = 2
rlabel pdiffusion 391 107 392 108  0 t = 3
rlabel pdiffusion 394 107 395 108  0 t = 4
rlabel pdiffusion 390 102 396 108 0 cell no = 334
<< m1 >>
rect 391 102 392 103 
rect 394 102 395 103 
rect 391 107 392 108 
rect 394 107 395 108 
<< m2 >>
rect 391 102 392 103 
rect 394 102 395 103 
rect 391 107 392 108 
rect 394 107 395 108 
<< m2c >>
rect 391 102 392 103 
rect 394 102 395 103 
rect 391 107 392 108 
rect 394 107 395 108 
<< labels >>
rlabel pdiffusion 427 408 428 409  0 t = 1
rlabel pdiffusion 430 408 431 409  0 t = 2
rlabel pdiffusion 427 413 428 414  0 t = 3
rlabel pdiffusion 430 413 431 414  0 t = 4
rlabel pdiffusion 426 408 432 414 0 cell no = 335
<< m1 >>
rect 427 408 428 409 
rect 430 408 431 409 
rect 427 413 428 414 
rect 430 413 431 414 
<< m2 >>
rect 427 408 428 409 
rect 430 408 431 409 
rect 427 413 428 414 
rect 430 413 431 414 
<< m2c >>
rect 427 408 428 409 
rect 430 408 431 409 
rect 427 413 428 414 
rect 430 413 431 414 
<< labels >>
rlabel pdiffusion 265 174 266 175  0 t = 1
rlabel pdiffusion 268 174 269 175  0 t = 2
rlabel pdiffusion 265 179 266 180  0 t = 3
rlabel pdiffusion 268 179 269 180  0 t = 4
rlabel pdiffusion 264 174 270 180 0 cell no = 336
<< m1 >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< m2 >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< m2c >>
rect 265 174 266 175 
rect 268 174 269 175 
rect 265 179 266 180 
rect 268 179 269 180 
<< labels >>
rlabel pdiffusion 211 246 212 247  0 t = 1
rlabel pdiffusion 214 246 215 247  0 t = 2
rlabel pdiffusion 211 251 212 252  0 t = 3
rlabel pdiffusion 214 251 215 252  0 t = 4
rlabel pdiffusion 210 246 216 252 0 cell no = 337
<< m1 >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< m2 >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< m2c >>
rect 211 246 212 247 
rect 214 246 215 247 
rect 211 251 212 252 
rect 214 251 215 252 
<< labels >>
rlabel pdiffusion 121 30 122 31  0 t = 1
rlabel pdiffusion 124 30 125 31  0 t = 2
rlabel pdiffusion 121 35 122 36  0 t = 3
rlabel pdiffusion 124 35 125 36  0 t = 4
rlabel pdiffusion 120 30 126 36 0 cell no = 338
<< m1 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2 >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< m2c >>
rect 121 30 122 31 
rect 124 30 125 31 
rect 121 35 122 36 
rect 124 35 125 36 
<< labels >>
rlabel pdiffusion 265 228 266 229  0 t = 1
rlabel pdiffusion 268 228 269 229  0 t = 2
rlabel pdiffusion 265 233 266 234  0 t = 3
rlabel pdiffusion 268 233 269 234  0 t = 4
rlabel pdiffusion 264 228 270 234 0 cell no = 339
<< m1 >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< m2 >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< m2c >>
rect 265 228 266 229 
rect 268 228 269 229 
rect 265 233 266 234 
rect 268 233 269 234 
<< labels >>
rlabel pdiffusion 301 282 302 283  0 t = 1
rlabel pdiffusion 304 282 305 283  0 t = 2
rlabel pdiffusion 301 287 302 288  0 t = 3
rlabel pdiffusion 304 287 305 288  0 t = 4
rlabel pdiffusion 300 282 306 288 0 cell no = 340
<< m1 >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< m2 >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< m2c >>
rect 301 282 302 283 
rect 304 282 305 283 
rect 301 287 302 288 
rect 304 287 305 288 
<< labels >>
rlabel pdiffusion 517 336 518 337  0 t = 1
rlabel pdiffusion 520 336 521 337  0 t = 2
rlabel pdiffusion 517 341 518 342  0 t = 3
rlabel pdiffusion 520 341 521 342  0 t = 4
rlabel pdiffusion 516 336 522 342 0 cell no = 341
<< m1 >>
rect 517 336 518 337 
rect 520 336 521 337 
rect 517 341 518 342 
rect 520 341 521 342 
<< m2 >>
rect 517 336 518 337 
rect 520 336 521 337 
rect 517 341 518 342 
rect 520 341 521 342 
<< m2c >>
rect 517 336 518 337 
rect 520 336 521 337 
rect 517 341 518 342 
rect 520 341 521 342 
<< labels >>
rlabel pdiffusion 427 48 428 49  0 t = 1
rlabel pdiffusion 430 48 431 49  0 t = 2
rlabel pdiffusion 427 53 428 54  0 t = 3
rlabel pdiffusion 430 53 431 54  0 t = 4
rlabel pdiffusion 426 48 432 54 0 cell no = 342
<< m1 >>
rect 427 48 428 49 
rect 430 48 431 49 
rect 427 53 428 54 
rect 430 53 431 54 
<< m2 >>
rect 427 48 428 49 
rect 430 48 431 49 
rect 427 53 428 54 
rect 430 53 431 54 
<< m2c >>
rect 427 48 428 49 
rect 430 48 431 49 
rect 427 53 428 54 
rect 430 53 431 54 
<< labels >>
rlabel pdiffusion 499 264 500 265  0 t = 1
rlabel pdiffusion 502 264 503 265  0 t = 2
rlabel pdiffusion 499 269 500 270  0 t = 3
rlabel pdiffusion 502 269 503 270  0 t = 4
rlabel pdiffusion 498 264 504 270 0 cell no = 343
<< m1 >>
rect 499 264 500 265 
rect 502 264 503 265 
rect 499 269 500 270 
rect 502 269 503 270 
<< m2 >>
rect 499 264 500 265 
rect 502 264 503 265 
rect 499 269 500 270 
rect 502 269 503 270 
<< m2c >>
rect 499 264 500 265 
rect 502 264 503 265 
rect 499 269 500 270 
rect 502 269 503 270 
<< labels >>
rlabel pdiffusion 463 354 464 355  0 t = 1
rlabel pdiffusion 466 354 467 355  0 t = 2
rlabel pdiffusion 463 359 464 360  0 t = 3
rlabel pdiffusion 466 359 467 360  0 t = 4
rlabel pdiffusion 462 354 468 360 0 cell no = 344
<< m1 >>
rect 463 354 464 355 
rect 466 354 467 355 
rect 463 359 464 360 
rect 466 359 467 360 
<< m2 >>
rect 463 354 464 355 
rect 466 354 467 355 
rect 463 359 464 360 
rect 466 359 467 360 
<< m2c >>
rect 463 354 464 355 
rect 466 354 467 355 
rect 463 359 464 360 
rect 466 359 467 360 
<< labels >>
rlabel pdiffusion 157 282 158 283  0 t = 1
rlabel pdiffusion 160 282 161 283  0 t = 2
rlabel pdiffusion 157 287 158 288  0 t = 3
rlabel pdiffusion 160 287 161 288  0 t = 4
rlabel pdiffusion 156 282 162 288 0 cell no = 345
<< m1 >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< m2 >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< m2c >>
rect 157 282 158 283 
rect 160 282 161 283 
rect 157 287 158 288 
rect 160 287 161 288 
<< labels >>
rlabel pdiffusion 283 66 284 67  0 t = 1
rlabel pdiffusion 286 66 287 67  0 t = 2
rlabel pdiffusion 283 71 284 72  0 t = 3
rlabel pdiffusion 286 71 287 72  0 t = 4
rlabel pdiffusion 282 66 288 72 0 cell no = 346
<< m1 >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< m2 >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< m2c >>
rect 283 66 284 67 
rect 286 66 287 67 
rect 283 71 284 72 
rect 286 71 287 72 
<< labels >>
rlabel pdiffusion 499 210 500 211  0 t = 1
rlabel pdiffusion 502 210 503 211  0 t = 2
rlabel pdiffusion 499 215 500 216  0 t = 3
rlabel pdiffusion 502 215 503 216  0 t = 4
rlabel pdiffusion 498 210 504 216 0 cell no = 347
<< m1 >>
rect 499 210 500 211 
rect 502 210 503 211 
rect 499 215 500 216 
rect 502 215 503 216 
<< m2 >>
rect 499 210 500 211 
rect 502 210 503 211 
rect 499 215 500 216 
rect 502 215 503 216 
<< m2c >>
rect 499 210 500 211 
rect 502 210 503 211 
rect 499 215 500 216 
rect 502 215 503 216 
<< labels >>
rlabel pdiffusion 391 318 392 319  0 t = 1
rlabel pdiffusion 394 318 395 319  0 t = 2
rlabel pdiffusion 391 323 392 324  0 t = 3
rlabel pdiffusion 394 323 395 324  0 t = 4
rlabel pdiffusion 390 318 396 324 0 cell no = 348
<< m1 >>
rect 391 318 392 319 
rect 394 318 395 319 
rect 391 323 392 324 
rect 394 323 395 324 
<< m2 >>
rect 391 318 392 319 
rect 394 318 395 319 
rect 391 323 392 324 
rect 394 323 395 324 
<< m2c >>
rect 391 318 392 319 
rect 394 318 395 319 
rect 391 323 392 324 
rect 394 323 395 324 
<< labels >>
rlabel pdiffusion 13 282 14 283  0 t = 1
rlabel pdiffusion 16 282 17 283  0 t = 2
rlabel pdiffusion 13 287 14 288  0 t = 3
rlabel pdiffusion 16 287 17 288  0 t = 4
rlabel pdiffusion 12 282 18 288 0 cell no = 349
<< m1 >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< m2 >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< m2c >>
rect 13 282 14 283 
rect 16 282 17 283 
rect 13 287 14 288 
rect 16 287 17 288 
<< labels >>
rlabel pdiffusion 175 210 176 211  0 t = 1
rlabel pdiffusion 178 210 179 211  0 t = 2
rlabel pdiffusion 175 215 176 216  0 t = 3
rlabel pdiffusion 178 215 179 216  0 t = 4
rlabel pdiffusion 174 210 180 216 0 cell no = 350
<< m1 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2 >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< m2c >>
rect 175 210 176 211 
rect 178 210 179 211 
rect 175 215 176 216 
rect 178 215 179 216 
<< labels >>
rlabel pdiffusion 175 246 176 247  0 t = 1
rlabel pdiffusion 178 246 179 247  0 t = 2
rlabel pdiffusion 175 251 176 252  0 t = 3
rlabel pdiffusion 178 251 179 252  0 t = 4
rlabel pdiffusion 174 246 180 252 0 cell no = 351
<< m1 >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< m2 >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< m2c >>
rect 175 246 176 247 
rect 178 246 179 247 
rect 175 251 176 252 
rect 178 251 179 252 
<< labels >>
rlabel pdiffusion 211 84 212 85  0 t = 1
rlabel pdiffusion 214 84 215 85  0 t = 2
rlabel pdiffusion 211 89 212 90  0 t = 3
rlabel pdiffusion 214 89 215 90  0 t = 4
rlabel pdiffusion 210 84 216 90 0 cell no = 352
<< m1 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2 >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< m2c >>
rect 211 84 212 85 
rect 214 84 215 85 
rect 211 89 212 90 
rect 214 89 215 90 
<< labels >>
rlabel pdiffusion 13 300 14 301  0 t = 1
rlabel pdiffusion 16 300 17 301  0 t = 2
rlabel pdiffusion 13 305 14 306  0 t = 3
rlabel pdiffusion 16 305 17 306  0 t = 4
rlabel pdiffusion 12 300 18 306 0 cell no = 353
<< m1 >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< m2 >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< m2c >>
rect 13 300 14 301 
rect 16 300 17 301 
rect 13 305 14 306 
rect 16 305 17 306 
<< labels >>
rlabel pdiffusion 49 408 50 409  0 t = 1
rlabel pdiffusion 52 408 53 409  0 t = 2
rlabel pdiffusion 49 413 50 414  0 t = 3
rlabel pdiffusion 52 413 53 414  0 t = 4
rlabel pdiffusion 48 408 54 414 0 cell no = 354
<< m1 >>
rect 49 408 50 409 
rect 52 408 53 409 
rect 49 413 50 414 
rect 52 413 53 414 
<< m2 >>
rect 49 408 50 409 
rect 52 408 53 409 
rect 49 413 50 414 
rect 52 413 53 414 
<< m2c >>
rect 49 408 50 409 
rect 52 408 53 409 
rect 49 413 50 414 
rect 52 413 53 414 
<< labels >>
rlabel pdiffusion 49 336 50 337  0 t = 1
rlabel pdiffusion 52 336 53 337  0 t = 2
rlabel pdiffusion 49 341 50 342  0 t = 3
rlabel pdiffusion 52 341 53 342  0 t = 4
rlabel pdiffusion 48 336 54 342 0 cell no = 355
<< m1 >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< m2 >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< m2c >>
rect 49 336 50 337 
rect 52 336 53 337 
rect 49 341 50 342 
rect 52 341 53 342 
<< labels >>
rlabel pdiffusion 247 498 248 499  0 t = 1
rlabel pdiffusion 250 498 251 499  0 t = 2
rlabel pdiffusion 247 503 248 504  0 t = 3
rlabel pdiffusion 250 503 251 504  0 t = 4
rlabel pdiffusion 246 498 252 504 0 cell no = 356
<< m1 >>
rect 247 498 248 499 
rect 250 498 251 499 
rect 247 503 248 504 
rect 250 503 251 504 
<< m2 >>
rect 247 498 248 499 
rect 250 498 251 499 
rect 247 503 248 504 
rect 250 503 251 504 
<< m2c >>
rect 247 498 248 499 
rect 250 498 251 499 
rect 247 503 248 504 
rect 250 503 251 504 
<< labels >>
rlabel pdiffusion 175 426 176 427  0 t = 1
rlabel pdiffusion 178 426 179 427  0 t = 2
rlabel pdiffusion 175 431 176 432  0 t = 3
rlabel pdiffusion 178 431 179 432  0 t = 4
rlabel pdiffusion 174 426 180 432 0 cell no = 357
<< m1 >>
rect 175 426 176 427 
rect 178 426 179 427 
rect 175 431 176 432 
rect 178 431 179 432 
<< m2 >>
rect 175 426 176 427 
rect 178 426 179 427 
rect 175 431 176 432 
rect 178 431 179 432 
<< m2c >>
rect 175 426 176 427 
rect 178 426 179 427 
rect 175 431 176 432 
rect 178 431 179 432 
<< labels >>
rlabel pdiffusion 139 300 140 301  0 t = 1
rlabel pdiffusion 142 300 143 301  0 t = 2
rlabel pdiffusion 139 305 140 306  0 t = 3
rlabel pdiffusion 142 305 143 306  0 t = 4
rlabel pdiffusion 138 300 144 306 0 cell no = 358
<< m1 >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< m2 >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< m2c >>
rect 139 300 140 301 
rect 142 300 143 301 
rect 139 305 140 306 
rect 142 305 143 306 
<< labels >>
rlabel pdiffusion 247 228 248 229  0 t = 1
rlabel pdiffusion 250 228 251 229  0 t = 2
rlabel pdiffusion 247 233 248 234  0 t = 3
rlabel pdiffusion 250 233 251 234  0 t = 4
rlabel pdiffusion 246 228 252 234 0 cell no = 359
<< m1 >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< m2 >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< m2c >>
rect 247 228 248 229 
rect 250 228 251 229 
rect 247 233 248 234 
rect 250 233 251 234 
<< labels >>
rlabel pdiffusion 355 354 356 355  0 t = 1
rlabel pdiffusion 358 354 359 355  0 t = 2
rlabel pdiffusion 355 359 356 360  0 t = 3
rlabel pdiffusion 358 359 359 360  0 t = 4
rlabel pdiffusion 354 354 360 360 0 cell no = 360
<< m1 >>
rect 355 354 356 355 
rect 358 354 359 355 
rect 355 359 356 360 
rect 358 359 359 360 
<< m2 >>
rect 355 354 356 355 
rect 358 354 359 355 
rect 355 359 356 360 
rect 358 359 359 360 
<< m2c >>
rect 355 354 356 355 
rect 358 354 359 355 
rect 355 359 356 360 
rect 358 359 359 360 
<< labels >>
rlabel pdiffusion 409 372 410 373  0 t = 1
rlabel pdiffusion 412 372 413 373  0 t = 2
rlabel pdiffusion 409 377 410 378  0 t = 3
rlabel pdiffusion 412 377 413 378  0 t = 4
rlabel pdiffusion 408 372 414 378 0 cell no = 361
<< m1 >>
rect 409 372 410 373 
rect 412 372 413 373 
rect 409 377 410 378 
rect 412 377 413 378 
<< m2 >>
rect 409 372 410 373 
rect 412 372 413 373 
rect 409 377 410 378 
rect 412 377 413 378 
<< m2c >>
rect 409 372 410 373 
rect 412 372 413 373 
rect 409 377 410 378 
rect 412 377 413 378 
<< labels >>
rlabel pdiffusion 157 300 158 301  0 t = 1
rlabel pdiffusion 160 300 161 301  0 t = 2
rlabel pdiffusion 157 305 158 306  0 t = 3
rlabel pdiffusion 160 305 161 306  0 t = 4
rlabel pdiffusion 156 300 162 306 0 cell no = 362
<< m1 >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< m2 >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< m2c >>
rect 157 300 158 301 
rect 160 300 161 301 
rect 157 305 158 306 
rect 160 305 161 306 
<< labels >>
rlabel pdiffusion 229 138 230 139  0 t = 1
rlabel pdiffusion 232 138 233 139  0 t = 2
rlabel pdiffusion 229 143 230 144  0 t = 3
rlabel pdiffusion 232 143 233 144  0 t = 4
rlabel pdiffusion 228 138 234 144 0 cell no = 363
<< m1 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2 >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< m2c >>
rect 229 138 230 139 
rect 232 138 233 139 
rect 229 143 230 144 
rect 232 143 233 144 
<< labels >>
rlabel pdiffusion 445 210 446 211  0 t = 1
rlabel pdiffusion 448 210 449 211  0 t = 2
rlabel pdiffusion 445 215 446 216  0 t = 3
rlabel pdiffusion 448 215 449 216  0 t = 4
rlabel pdiffusion 444 210 450 216 0 cell no = 364
<< m1 >>
rect 445 210 446 211 
rect 448 210 449 211 
rect 445 215 446 216 
rect 448 215 449 216 
<< m2 >>
rect 445 210 446 211 
rect 448 210 449 211 
rect 445 215 446 216 
rect 448 215 449 216 
<< m2c >>
rect 445 210 446 211 
rect 448 210 449 211 
rect 445 215 446 216 
rect 448 215 449 216 
<< labels >>
rlabel pdiffusion 265 264 266 265  0 t = 1
rlabel pdiffusion 268 264 269 265  0 t = 2
rlabel pdiffusion 265 269 266 270  0 t = 3
rlabel pdiffusion 268 269 269 270  0 t = 4
rlabel pdiffusion 264 264 270 270 0 cell no = 365
<< m1 >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< m2 >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< m2c >>
rect 265 264 266 265 
rect 268 264 269 265 
rect 265 269 266 270 
rect 268 269 269 270 
<< labels >>
rlabel pdiffusion 517 444 518 445  0 t = 1
rlabel pdiffusion 520 444 521 445  0 t = 2
rlabel pdiffusion 517 449 518 450  0 t = 3
rlabel pdiffusion 520 449 521 450  0 t = 4
rlabel pdiffusion 516 444 522 450 0 cell no = 366
<< m1 >>
rect 517 444 518 445 
rect 520 444 521 445 
rect 517 449 518 450 
rect 520 449 521 450 
<< m2 >>
rect 517 444 518 445 
rect 520 444 521 445 
rect 517 449 518 450 
rect 520 449 521 450 
<< m2c >>
rect 517 444 518 445 
rect 520 444 521 445 
rect 517 449 518 450 
rect 520 449 521 450 
<< labels >>
rlabel pdiffusion 229 300 230 301  0 t = 1
rlabel pdiffusion 232 300 233 301  0 t = 2
rlabel pdiffusion 229 305 230 306  0 t = 3
rlabel pdiffusion 232 305 233 306  0 t = 4
rlabel pdiffusion 228 300 234 306 0 cell no = 367
<< m1 >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< m2 >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< m2c >>
rect 229 300 230 301 
rect 232 300 233 301 
rect 229 305 230 306 
rect 232 305 233 306 
<< labels >>
rlabel pdiffusion 409 318 410 319  0 t = 1
rlabel pdiffusion 412 318 413 319  0 t = 2
rlabel pdiffusion 409 323 410 324  0 t = 3
rlabel pdiffusion 412 323 413 324  0 t = 4
rlabel pdiffusion 408 318 414 324 0 cell no = 368
<< m1 >>
rect 409 318 410 319 
rect 412 318 413 319 
rect 409 323 410 324 
rect 412 323 413 324 
<< m2 >>
rect 409 318 410 319 
rect 412 318 413 319 
rect 409 323 410 324 
rect 412 323 413 324 
<< m2c >>
rect 409 318 410 319 
rect 412 318 413 319 
rect 409 323 410 324 
rect 412 323 413 324 
<< labels >>
rlabel pdiffusion 85 246 86 247  0 t = 1
rlabel pdiffusion 88 246 89 247  0 t = 2
rlabel pdiffusion 85 251 86 252  0 t = 3
rlabel pdiffusion 88 251 89 252  0 t = 4
rlabel pdiffusion 84 246 90 252 0 cell no = 369
<< m1 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2 >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< m2c >>
rect 85 246 86 247 
rect 88 246 89 247 
rect 85 251 86 252 
rect 88 251 89 252 
<< labels >>
rlabel pdiffusion 373 174 374 175  0 t = 1
rlabel pdiffusion 376 174 377 175  0 t = 2
rlabel pdiffusion 373 179 374 180  0 t = 3
rlabel pdiffusion 376 179 377 180  0 t = 4
rlabel pdiffusion 372 174 378 180 0 cell no = 370
<< m1 >>
rect 373 174 374 175 
rect 376 174 377 175 
rect 373 179 374 180 
rect 376 179 377 180 
<< m2 >>
rect 373 174 374 175 
rect 376 174 377 175 
rect 373 179 374 180 
rect 376 179 377 180 
<< m2c >>
rect 373 174 374 175 
rect 376 174 377 175 
rect 373 179 374 180 
rect 376 179 377 180 
<< labels >>
rlabel pdiffusion 13 372 14 373  0 t = 1
rlabel pdiffusion 16 372 17 373  0 t = 2
rlabel pdiffusion 13 377 14 378  0 t = 3
rlabel pdiffusion 16 377 17 378  0 t = 4
rlabel pdiffusion 12 372 18 378 0 cell no = 371
<< m1 >>
rect 13 372 14 373 
rect 16 372 17 373 
rect 13 377 14 378 
rect 16 377 17 378 
<< m2 >>
rect 13 372 14 373 
rect 16 372 17 373 
rect 13 377 14 378 
rect 16 377 17 378 
<< m2c >>
rect 13 372 14 373 
rect 16 372 17 373 
rect 13 377 14 378 
rect 16 377 17 378 
<< labels >>
rlabel pdiffusion 445 462 446 463  0 t = 1
rlabel pdiffusion 448 462 449 463  0 t = 2
rlabel pdiffusion 445 467 446 468  0 t = 3
rlabel pdiffusion 448 467 449 468  0 t = 4
rlabel pdiffusion 444 462 450 468 0 cell no = 372
<< m1 >>
rect 445 462 446 463 
rect 448 462 449 463 
rect 445 467 446 468 
rect 448 467 449 468 
<< m2 >>
rect 445 462 446 463 
rect 448 462 449 463 
rect 445 467 446 468 
rect 448 467 449 468 
<< m2c >>
rect 445 462 446 463 
rect 448 462 449 463 
rect 445 467 446 468 
rect 448 467 449 468 
<< labels >>
rlabel pdiffusion 499 102 500 103  0 t = 1
rlabel pdiffusion 502 102 503 103  0 t = 2
rlabel pdiffusion 499 107 500 108  0 t = 3
rlabel pdiffusion 502 107 503 108  0 t = 4
rlabel pdiffusion 498 102 504 108 0 cell no = 373
<< m1 >>
rect 499 102 500 103 
rect 502 102 503 103 
rect 499 107 500 108 
rect 502 107 503 108 
<< m2 >>
rect 499 102 500 103 
rect 502 102 503 103 
rect 499 107 500 108 
rect 502 107 503 108 
<< m2c >>
rect 499 102 500 103 
rect 502 102 503 103 
rect 499 107 500 108 
rect 502 107 503 108 
<< labels >>
rlabel pdiffusion 463 192 464 193  0 t = 1
rlabel pdiffusion 466 192 467 193  0 t = 2
rlabel pdiffusion 463 197 464 198  0 t = 3
rlabel pdiffusion 466 197 467 198  0 t = 4
rlabel pdiffusion 462 192 468 198 0 cell no = 374
<< m1 >>
rect 463 192 464 193 
rect 466 192 467 193 
rect 463 197 464 198 
rect 466 197 467 198 
<< m2 >>
rect 463 192 464 193 
rect 466 192 467 193 
rect 463 197 464 198 
rect 466 197 467 198 
<< m2c >>
rect 463 192 464 193 
rect 466 192 467 193 
rect 463 197 464 198 
rect 466 197 467 198 
<< labels >>
rlabel pdiffusion 13 30 14 31  0 t = 1
rlabel pdiffusion 16 30 17 31  0 t = 2
rlabel pdiffusion 13 35 14 36  0 t = 3
rlabel pdiffusion 16 35 17 36  0 t = 4
rlabel pdiffusion 12 30 18 36 0 cell no = 375
<< m1 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2 >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< m2c >>
rect 13 30 14 31 
rect 16 30 17 31 
rect 13 35 14 36 
rect 16 35 17 36 
<< labels >>
rlabel pdiffusion 463 210 464 211  0 t = 1
rlabel pdiffusion 466 210 467 211  0 t = 2
rlabel pdiffusion 463 215 464 216  0 t = 3
rlabel pdiffusion 466 215 467 216  0 t = 4
rlabel pdiffusion 462 210 468 216 0 cell no = 376
<< m1 >>
rect 463 210 464 211 
rect 466 210 467 211 
rect 463 215 464 216 
rect 466 215 467 216 
<< m2 >>
rect 463 210 464 211 
rect 466 210 467 211 
rect 463 215 464 216 
rect 466 215 467 216 
<< m2c >>
rect 463 210 464 211 
rect 466 210 467 211 
rect 463 215 464 216 
rect 466 215 467 216 
<< labels >>
rlabel pdiffusion 139 102 140 103  0 t = 1
rlabel pdiffusion 142 102 143 103  0 t = 2
rlabel pdiffusion 139 107 140 108  0 t = 3
rlabel pdiffusion 142 107 143 108  0 t = 4
rlabel pdiffusion 138 102 144 108 0 cell no = 377
<< m1 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2 >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< m2c >>
rect 139 102 140 103 
rect 142 102 143 103 
rect 139 107 140 108 
rect 142 107 143 108 
<< labels >>
rlabel pdiffusion 13 390 14 391  0 t = 1
rlabel pdiffusion 16 390 17 391  0 t = 2
rlabel pdiffusion 13 395 14 396  0 t = 3
rlabel pdiffusion 16 395 17 396  0 t = 4
rlabel pdiffusion 12 390 18 396 0 cell no = 378
<< m1 >>
rect 13 390 14 391 
rect 16 390 17 391 
rect 13 395 14 396 
rect 16 395 17 396 
<< m2 >>
rect 13 390 14 391 
rect 16 390 17 391 
rect 13 395 14 396 
rect 16 395 17 396 
<< m2c >>
rect 13 390 14 391 
rect 16 390 17 391 
rect 13 395 14 396 
rect 16 395 17 396 
<< labels >>
rlabel pdiffusion 31 210 32 211  0 t = 1
rlabel pdiffusion 34 210 35 211  0 t = 2
rlabel pdiffusion 31 215 32 216  0 t = 3
rlabel pdiffusion 34 215 35 216  0 t = 4
rlabel pdiffusion 30 210 36 216 0 cell no = 379
<< m1 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2 >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< m2c >>
rect 31 210 32 211 
rect 34 210 35 211 
rect 31 215 32 216 
rect 34 215 35 216 
<< labels >>
rlabel pdiffusion 49 480 50 481  0 t = 1
rlabel pdiffusion 52 480 53 481  0 t = 2
rlabel pdiffusion 49 485 50 486  0 t = 3
rlabel pdiffusion 52 485 53 486  0 t = 4
rlabel pdiffusion 48 480 54 486 0 cell no = 380
<< m1 >>
rect 49 480 50 481 
rect 52 480 53 481 
rect 49 485 50 486 
rect 52 485 53 486 
<< m2 >>
rect 49 480 50 481 
rect 52 480 53 481 
rect 49 485 50 486 
rect 52 485 53 486 
<< m2c >>
rect 49 480 50 481 
rect 52 480 53 481 
rect 49 485 50 486 
rect 52 485 53 486 
<< labels >>
rlabel pdiffusion 103 210 104 211  0 t = 1
rlabel pdiffusion 106 210 107 211  0 t = 2
rlabel pdiffusion 103 215 104 216  0 t = 3
rlabel pdiffusion 106 215 107 216  0 t = 4
rlabel pdiffusion 102 210 108 216 0 cell no = 381
<< m1 >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< m2 >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< m2c >>
rect 103 210 104 211 
rect 106 210 107 211 
rect 103 215 104 216 
rect 106 215 107 216 
<< labels >>
rlabel pdiffusion 121 174 122 175  0 t = 1
rlabel pdiffusion 124 174 125 175  0 t = 2
rlabel pdiffusion 121 179 122 180  0 t = 3
rlabel pdiffusion 124 179 125 180  0 t = 4
rlabel pdiffusion 120 174 126 180 0 cell no = 382
<< m1 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2 >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< m2c >>
rect 121 174 122 175 
rect 124 174 125 175 
rect 121 179 122 180 
rect 124 179 125 180 
<< labels >>
rlabel pdiffusion 391 84 392 85  0 t = 1
rlabel pdiffusion 394 84 395 85  0 t = 2
rlabel pdiffusion 391 89 392 90  0 t = 3
rlabel pdiffusion 394 89 395 90  0 t = 4
rlabel pdiffusion 390 84 396 90 0 cell no = 383
<< m1 >>
rect 391 84 392 85 
rect 394 84 395 85 
rect 391 89 392 90 
rect 394 89 395 90 
<< m2 >>
rect 391 84 392 85 
rect 394 84 395 85 
rect 391 89 392 90 
rect 394 89 395 90 
<< m2c >>
rect 391 84 392 85 
rect 394 84 395 85 
rect 391 89 392 90 
rect 394 89 395 90 
<< labels >>
rlabel pdiffusion 409 120 410 121  0 t = 1
rlabel pdiffusion 412 120 413 121  0 t = 2
rlabel pdiffusion 409 125 410 126  0 t = 3
rlabel pdiffusion 412 125 413 126  0 t = 4
rlabel pdiffusion 408 120 414 126 0 cell no = 384
<< m1 >>
rect 409 120 410 121 
rect 412 120 413 121 
rect 409 125 410 126 
rect 412 125 413 126 
<< m2 >>
rect 409 120 410 121 
rect 412 120 413 121 
rect 409 125 410 126 
rect 412 125 413 126 
<< m2c >>
rect 409 120 410 121 
rect 412 120 413 121 
rect 409 125 410 126 
rect 412 125 413 126 
<< labels >>
rlabel pdiffusion 49 210 50 211  0 t = 1
rlabel pdiffusion 52 210 53 211  0 t = 2
rlabel pdiffusion 49 215 50 216  0 t = 3
rlabel pdiffusion 52 215 53 216  0 t = 4
rlabel pdiffusion 48 210 54 216 0 cell no = 385
<< m1 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2 >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< m2c >>
rect 49 210 50 211 
rect 52 210 53 211 
rect 49 215 50 216 
rect 52 215 53 216 
<< labels >>
rlabel pdiffusion 319 210 320 211  0 t = 1
rlabel pdiffusion 322 210 323 211  0 t = 2
rlabel pdiffusion 319 215 320 216  0 t = 3
rlabel pdiffusion 322 215 323 216  0 t = 4
rlabel pdiffusion 318 210 324 216 0 cell no = 386
<< m1 >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< m2 >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< m2c >>
rect 319 210 320 211 
rect 322 210 323 211 
rect 319 215 320 216 
rect 322 215 323 216 
<< labels >>
rlabel pdiffusion 373 462 374 463  0 t = 1
rlabel pdiffusion 376 462 377 463  0 t = 2
rlabel pdiffusion 373 467 374 468  0 t = 3
rlabel pdiffusion 376 467 377 468  0 t = 4
rlabel pdiffusion 372 462 378 468 0 cell no = 387
<< m1 >>
rect 373 462 374 463 
rect 376 462 377 463 
rect 373 467 374 468 
rect 376 467 377 468 
<< m2 >>
rect 373 462 374 463 
rect 376 462 377 463 
rect 373 467 374 468 
rect 376 467 377 468 
<< m2c >>
rect 373 462 374 463 
rect 376 462 377 463 
rect 373 467 374 468 
rect 376 467 377 468 
<< labels >>
rlabel pdiffusion 445 12 446 13  0 t = 1
rlabel pdiffusion 448 12 449 13  0 t = 2
rlabel pdiffusion 445 17 446 18  0 t = 3
rlabel pdiffusion 448 17 449 18  0 t = 4
rlabel pdiffusion 444 12 450 18 0 cell no = 388
<< m1 >>
rect 445 12 446 13 
rect 448 12 449 13 
rect 445 17 446 18 
rect 448 17 449 18 
<< m2 >>
rect 445 12 446 13 
rect 448 12 449 13 
rect 445 17 446 18 
rect 448 17 449 18 
<< m2c >>
rect 445 12 446 13 
rect 448 12 449 13 
rect 445 17 446 18 
rect 448 17 449 18 
<< labels >>
rlabel pdiffusion 391 282 392 283  0 t = 1
rlabel pdiffusion 394 282 395 283  0 t = 2
rlabel pdiffusion 391 287 392 288  0 t = 3
rlabel pdiffusion 394 287 395 288  0 t = 4
rlabel pdiffusion 390 282 396 288 0 cell no = 389
<< m1 >>
rect 391 282 392 283 
rect 394 282 395 283 
rect 391 287 392 288 
rect 394 287 395 288 
<< m2 >>
rect 391 282 392 283 
rect 394 282 395 283 
rect 391 287 392 288 
rect 394 287 395 288 
<< m2c >>
rect 391 282 392 283 
rect 394 282 395 283 
rect 391 287 392 288 
rect 394 287 395 288 
<< labels >>
rlabel pdiffusion 463 102 464 103  0 t = 1
rlabel pdiffusion 466 102 467 103  0 t = 2
rlabel pdiffusion 463 107 464 108  0 t = 3
rlabel pdiffusion 466 107 467 108  0 t = 4
rlabel pdiffusion 462 102 468 108 0 cell no = 390
<< m1 >>
rect 463 102 464 103 
rect 466 102 467 103 
rect 463 107 464 108 
rect 466 107 467 108 
<< m2 >>
rect 463 102 464 103 
rect 466 102 467 103 
rect 463 107 464 108 
rect 466 107 467 108 
<< m2c >>
rect 463 102 464 103 
rect 466 102 467 103 
rect 463 107 464 108 
rect 466 107 467 108 
<< labels >>
rlabel pdiffusion 283 174 284 175  0 t = 1
rlabel pdiffusion 286 174 287 175  0 t = 2
rlabel pdiffusion 283 179 284 180  0 t = 3
rlabel pdiffusion 286 179 287 180  0 t = 4
rlabel pdiffusion 282 174 288 180 0 cell no = 391
<< m1 >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< m2 >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< m2c >>
rect 283 174 284 175 
rect 286 174 287 175 
rect 283 179 284 180 
rect 286 179 287 180 
<< labels >>
rlabel pdiffusion 49 12 50 13  0 t = 1
rlabel pdiffusion 52 12 53 13  0 t = 2
rlabel pdiffusion 49 17 50 18  0 t = 3
rlabel pdiffusion 52 17 53 18  0 t = 4
rlabel pdiffusion 48 12 54 18 0 cell no = 392
<< m1 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2 >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< m2c >>
rect 49 12 50 13 
rect 52 12 53 13 
rect 49 17 50 18 
rect 52 17 53 18 
<< labels >>
rlabel pdiffusion 67 120 68 121  0 t = 1
rlabel pdiffusion 70 120 71 121  0 t = 2
rlabel pdiffusion 67 125 68 126  0 t = 3
rlabel pdiffusion 70 125 71 126  0 t = 4
rlabel pdiffusion 66 120 72 126 0 cell no = 393
<< m1 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2 >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< m2c >>
rect 67 120 68 121 
rect 70 120 71 121 
rect 67 125 68 126 
rect 70 125 71 126 
<< labels >>
rlabel pdiffusion 211 300 212 301  0 t = 1
rlabel pdiffusion 214 300 215 301  0 t = 2
rlabel pdiffusion 211 305 212 306  0 t = 3
rlabel pdiffusion 214 305 215 306  0 t = 4
rlabel pdiffusion 210 300 216 306 0 cell no = 394
<< m1 >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< m2 >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< m2c >>
rect 211 300 212 301 
rect 214 300 215 301 
rect 211 305 212 306 
rect 214 305 215 306 
<< labels >>
rlabel pdiffusion 409 264 410 265  0 t = 1
rlabel pdiffusion 412 264 413 265  0 t = 2
rlabel pdiffusion 409 269 410 270  0 t = 3
rlabel pdiffusion 412 269 413 270  0 t = 4
rlabel pdiffusion 408 264 414 270 0 cell no = 395
<< m1 >>
rect 409 264 410 265 
rect 412 264 413 265 
rect 409 269 410 270 
rect 412 269 413 270 
<< m2 >>
rect 409 264 410 265 
rect 412 264 413 265 
rect 409 269 410 270 
rect 412 269 413 270 
<< m2c >>
rect 409 264 410 265 
rect 412 264 413 265 
rect 409 269 410 270 
rect 412 269 413 270 
<< labels >>
rlabel pdiffusion 175 318 176 319  0 t = 1
rlabel pdiffusion 178 318 179 319  0 t = 2
rlabel pdiffusion 175 323 176 324  0 t = 3
rlabel pdiffusion 178 323 179 324  0 t = 4
rlabel pdiffusion 174 318 180 324 0 cell no = 396
<< m1 >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< m2 >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< m2c >>
rect 175 318 176 319 
rect 178 318 179 319 
rect 175 323 176 324 
rect 178 323 179 324 
<< labels >>
rlabel pdiffusion 67 264 68 265  0 t = 1
rlabel pdiffusion 70 264 71 265  0 t = 2
rlabel pdiffusion 67 269 68 270  0 t = 3
rlabel pdiffusion 70 269 71 270  0 t = 4
rlabel pdiffusion 66 264 72 270 0 cell no = 397
<< m1 >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< m2 >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< m2c >>
rect 67 264 68 265 
rect 70 264 71 265 
rect 67 269 68 270 
rect 70 269 71 270 
<< labels >>
rlabel pdiffusion 157 210 158 211  0 t = 1
rlabel pdiffusion 160 210 161 211  0 t = 2
rlabel pdiffusion 157 215 158 216  0 t = 3
rlabel pdiffusion 160 215 161 216  0 t = 4
rlabel pdiffusion 156 210 162 216 0 cell no = 398
<< m1 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2 >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< m2c >>
rect 157 210 158 211 
rect 160 210 161 211 
rect 157 215 158 216 
rect 160 215 161 216 
<< labels >>
rlabel pdiffusion 355 228 356 229  0 t = 1
rlabel pdiffusion 358 228 359 229  0 t = 2
rlabel pdiffusion 355 233 356 234  0 t = 3
rlabel pdiffusion 358 233 359 234  0 t = 4
rlabel pdiffusion 354 228 360 234 0 cell no = 399
<< m1 >>
rect 355 228 356 229 
rect 358 228 359 229 
rect 355 233 356 234 
rect 358 233 359 234 
<< m2 >>
rect 355 228 356 229 
rect 358 228 359 229 
rect 355 233 356 234 
rect 358 233 359 234 
<< m2c >>
rect 355 228 356 229 
rect 358 228 359 229 
rect 355 233 356 234 
rect 358 233 359 234 
<< labels >>
rlabel pdiffusion 481 174 482 175  0 t = 1
rlabel pdiffusion 484 174 485 175  0 t = 2
rlabel pdiffusion 481 179 482 180  0 t = 3
rlabel pdiffusion 484 179 485 180  0 t = 4
rlabel pdiffusion 480 174 486 180 0 cell no = 400
<< m1 >>
rect 481 174 482 175 
rect 484 174 485 175 
rect 481 179 482 180 
rect 484 179 485 180 
<< m2 >>
rect 481 174 482 175 
rect 484 174 485 175 
rect 481 179 482 180 
rect 484 179 485 180 
<< m2c >>
rect 481 174 482 175 
rect 484 174 485 175 
rect 481 179 482 180 
rect 484 179 485 180 
<< labels >>
rlabel pdiffusion 517 246 518 247  0 t = 1
rlabel pdiffusion 520 246 521 247  0 t = 2
rlabel pdiffusion 517 251 518 252  0 t = 3
rlabel pdiffusion 520 251 521 252  0 t = 4
rlabel pdiffusion 516 246 522 252 0 cell no = 401
<< m1 >>
rect 517 246 518 247 
rect 520 246 521 247 
rect 517 251 518 252 
rect 520 251 521 252 
<< m2 >>
rect 517 246 518 247 
rect 520 246 521 247 
rect 517 251 518 252 
rect 520 251 521 252 
<< m2c >>
rect 517 246 518 247 
rect 520 246 521 247 
rect 517 251 518 252 
rect 520 251 521 252 
<< labels >>
rlabel pdiffusion 463 246 464 247  0 t = 1
rlabel pdiffusion 466 246 467 247  0 t = 2
rlabel pdiffusion 463 251 464 252  0 t = 3
rlabel pdiffusion 466 251 467 252  0 t = 4
rlabel pdiffusion 462 246 468 252 0 cell no = 402
<< m1 >>
rect 463 246 464 247 
rect 466 246 467 247 
rect 463 251 464 252 
rect 466 251 467 252 
<< m2 >>
rect 463 246 464 247 
rect 466 246 467 247 
rect 463 251 464 252 
rect 466 251 467 252 
<< m2c >>
rect 463 246 464 247 
rect 466 246 467 247 
rect 463 251 464 252 
rect 466 251 467 252 
<< labels >>
rlabel pdiffusion 265 120 266 121  0 t = 1
rlabel pdiffusion 268 120 269 121  0 t = 2
rlabel pdiffusion 265 125 266 126  0 t = 3
rlabel pdiffusion 268 125 269 126  0 t = 4
rlabel pdiffusion 264 120 270 126 0 cell no = 403
<< m1 >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< m2 >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< m2c >>
rect 265 120 266 121 
rect 268 120 269 121 
rect 265 125 266 126 
rect 268 125 269 126 
<< labels >>
rlabel pdiffusion 85 336 86 337  0 t = 1
rlabel pdiffusion 88 336 89 337  0 t = 2
rlabel pdiffusion 85 341 86 342  0 t = 3
rlabel pdiffusion 88 341 89 342  0 t = 4
rlabel pdiffusion 84 336 90 342 0 cell no = 404
<< m1 >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< m2 >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< m2c >>
rect 85 336 86 337 
rect 88 336 89 337 
rect 85 341 86 342 
rect 88 341 89 342 
<< labels >>
rlabel pdiffusion 427 174 428 175  0 t = 1
rlabel pdiffusion 430 174 431 175  0 t = 2
rlabel pdiffusion 427 179 428 180  0 t = 3
rlabel pdiffusion 430 179 431 180  0 t = 4
rlabel pdiffusion 426 174 432 180 0 cell no = 405
<< m1 >>
rect 427 174 428 175 
rect 430 174 431 175 
rect 427 179 428 180 
rect 430 179 431 180 
<< m2 >>
rect 427 174 428 175 
rect 430 174 431 175 
rect 427 179 428 180 
rect 430 179 431 180 
<< m2c >>
rect 427 174 428 175 
rect 430 174 431 175 
rect 427 179 428 180 
rect 430 179 431 180 
<< labels >>
rlabel pdiffusion 427 372 428 373  0 t = 1
rlabel pdiffusion 430 372 431 373  0 t = 2
rlabel pdiffusion 427 377 428 378  0 t = 3
rlabel pdiffusion 430 377 431 378  0 t = 4
rlabel pdiffusion 426 372 432 378 0 cell no = 406
<< m1 >>
rect 427 372 428 373 
rect 430 372 431 373 
rect 427 377 428 378 
rect 430 377 431 378 
<< m2 >>
rect 427 372 428 373 
rect 430 372 431 373 
rect 427 377 428 378 
rect 430 377 431 378 
<< m2c >>
rect 427 372 428 373 
rect 430 372 431 373 
rect 427 377 428 378 
rect 430 377 431 378 
<< labels >>
rlabel pdiffusion 85 156 86 157  0 t = 1
rlabel pdiffusion 88 156 89 157  0 t = 2
rlabel pdiffusion 85 161 86 162  0 t = 3
rlabel pdiffusion 88 161 89 162  0 t = 4
rlabel pdiffusion 84 156 90 162 0 cell no = 407
<< m1 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2 >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< m2c >>
rect 85 156 86 157 
rect 88 156 89 157 
rect 85 161 86 162 
rect 88 161 89 162 
<< labels >>
rlabel pdiffusion 31 354 32 355  0 t = 1
rlabel pdiffusion 34 354 35 355  0 t = 2
rlabel pdiffusion 31 359 32 360  0 t = 3
rlabel pdiffusion 34 359 35 360  0 t = 4
rlabel pdiffusion 30 354 36 360 0 cell no = 408
<< m1 >>
rect 31 354 32 355 
rect 34 354 35 355 
rect 31 359 32 360 
rect 34 359 35 360 
<< m2 >>
rect 31 354 32 355 
rect 34 354 35 355 
rect 31 359 32 360 
rect 34 359 35 360 
<< m2c >>
rect 31 354 32 355 
rect 34 354 35 355 
rect 31 359 32 360 
rect 34 359 35 360 
<< labels >>
rlabel pdiffusion 175 192 176 193  0 t = 1
rlabel pdiffusion 178 192 179 193  0 t = 2
rlabel pdiffusion 175 197 176 198  0 t = 3
rlabel pdiffusion 178 197 179 198  0 t = 4
rlabel pdiffusion 174 192 180 198 0 cell no = 409
<< m1 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2 >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< m2c >>
rect 175 192 176 193 
rect 178 192 179 193 
rect 175 197 176 198 
rect 178 197 179 198 
<< labels >>
rlabel pdiffusion 265 480 266 481  0 t = 1
rlabel pdiffusion 268 480 269 481  0 t = 2
rlabel pdiffusion 265 485 266 486  0 t = 3
rlabel pdiffusion 268 485 269 486  0 t = 4
rlabel pdiffusion 264 480 270 486 0 cell no = 410
<< m1 >>
rect 265 480 266 481 
rect 268 480 269 481 
rect 265 485 266 486 
rect 268 485 269 486 
<< m2 >>
rect 265 480 266 481 
rect 268 480 269 481 
rect 265 485 266 486 
rect 268 485 269 486 
<< m2c >>
rect 265 480 266 481 
rect 268 480 269 481 
rect 265 485 266 486 
rect 268 485 269 486 
<< labels >>
rlabel pdiffusion 211 264 212 265  0 t = 1
rlabel pdiffusion 214 264 215 265  0 t = 2
rlabel pdiffusion 211 269 212 270  0 t = 3
rlabel pdiffusion 214 269 215 270  0 t = 4
rlabel pdiffusion 210 264 216 270 0 cell no = 411
<< m1 >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< m2 >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< m2c >>
rect 211 264 212 265 
rect 214 264 215 265 
rect 211 269 212 270 
rect 214 269 215 270 
<< labels >>
rlabel pdiffusion 13 246 14 247  0 t = 1
rlabel pdiffusion 16 246 17 247  0 t = 2
rlabel pdiffusion 13 251 14 252  0 t = 3
rlabel pdiffusion 16 251 17 252  0 t = 4
rlabel pdiffusion 12 246 18 252 0 cell no = 412
<< m1 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2 >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< m2c >>
rect 13 246 14 247 
rect 16 246 17 247 
rect 13 251 14 252 
rect 16 251 17 252 
<< labels >>
rlabel pdiffusion 139 228 140 229  0 t = 1
rlabel pdiffusion 142 228 143 229  0 t = 2
rlabel pdiffusion 139 233 140 234  0 t = 3
rlabel pdiffusion 142 233 143 234  0 t = 4
rlabel pdiffusion 138 228 144 234 0 cell no = 413
<< m1 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2 >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< m2c >>
rect 139 228 140 229 
rect 142 228 143 229 
rect 139 233 140 234 
rect 142 233 143 234 
<< labels >>
rlabel pdiffusion 67 282 68 283  0 t = 1
rlabel pdiffusion 70 282 71 283  0 t = 2
rlabel pdiffusion 67 287 68 288  0 t = 3
rlabel pdiffusion 70 287 71 288  0 t = 4
rlabel pdiffusion 66 282 72 288 0 cell no = 414
<< m1 >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< m2 >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< m2c >>
rect 67 282 68 283 
rect 70 282 71 283 
rect 67 287 68 288 
rect 70 287 71 288 
<< labels >>
rlabel pdiffusion 175 12 176 13  0 t = 1
rlabel pdiffusion 178 12 179 13  0 t = 2
rlabel pdiffusion 175 17 176 18  0 t = 3
rlabel pdiffusion 178 17 179 18  0 t = 4
rlabel pdiffusion 174 12 180 18 0 cell no = 415
<< m1 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2 >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< m2c >>
rect 175 12 176 13 
rect 178 12 179 13 
rect 175 17 176 18 
rect 178 17 179 18 
<< labels >>
rlabel pdiffusion 31 192 32 193  0 t = 1
rlabel pdiffusion 34 192 35 193  0 t = 2
rlabel pdiffusion 31 197 32 198  0 t = 3
rlabel pdiffusion 34 197 35 198  0 t = 4
rlabel pdiffusion 30 192 36 198 0 cell no = 416
<< m1 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2 >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< m2c >>
rect 31 192 32 193 
rect 34 192 35 193 
rect 31 197 32 198 
rect 34 197 35 198 
<< labels >>
rlabel pdiffusion 67 354 68 355  0 t = 1
rlabel pdiffusion 70 354 71 355  0 t = 2
rlabel pdiffusion 67 359 68 360  0 t = 3
rlabel pdiffusion 70 359 71 360  0 t = 4
rlabel pdiffusion 66 354 72 360 0 cell no = 417
<< m1 >>
rect 67 354 68 355 
rect 70 354 71 355 
rect 67 359 68 360 
rect 70 359 71 360 
<< m2 >>
rect 67 354 68 355 
rect 70 354 71 355 
rect 67 359 68 360 
rect 70 359 71 360 
<< m2c >>
rect 67 354 68 355 
rect 70 354 71 355 
rect 67 359 68 360 
rect 70 359 71 360 
<< labels >>
rlabel pdiffusion 139 282 140 283  0 t = 1
rlabel pdiffusion 142 282 143 283  0 t = 2
rlabel pdiffusion 139 287 140 288  0 t = 3
rlabel pdiffusion 142 287 143 288  0 t = 4
rlabel pdiffusion 138 282 144 288 0 cell no = 418
<< m1 >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< m2 >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< m2c >>
rect 139 282 140 283 
rect 142 282 143 283 
rect 139 287 140 288 
rect 142 287 143 288 
<< labels >>
rlabel pdiffusion 31 12 32 13  0 t = 1
rlabel pdiffusion 34 12 35 13  0 t = 2
rlabel pdiffusion 31 17 32 18  0 t = 3
rlabel pdiffusion 34 17 35 18  0 t = 4
rlabel pdiffusion 30 12 36 18 0 cell no = 419
<< m1 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2 >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< m2c >>
rect 31 12 32 13 
rect 34 12 35 13 
rect 31 17 32 18 
rect 34 17 35 18 
<< labels >>
rlabel pdiffusion 193 156 194 157  0 t = 1
rlabel pdiffusion 196 156 197 157  0 t = 2
rlabel pdiffusion 193 161 194 162  0 t = 3
rlabel pdiffusion 196 161 197 162  0 t = 4
rlabel pdiffusion 192 156 198 162 0 cell no = 420
<< m1 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2 >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< m2c >>
rect 193 156 194 157 
rect 196 156 197 157 
rect 193 161 194 162 
rect 196 161 197 162 
<< labels >>
rlabel pdiffusion 337 282 338 283  0 t = 1
rlabel pdiffusion 340 282 341 283  0 t = 2
rlabel pdiffusion 337 287 338 288  0 t = 3
rlabel pdiffusion 340 287 341 288  0 t = 4
rlabel pdiffusion 336 282 342 288 0 cell no = 421
<< m1 >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< m2 >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< m2c >>
rect 337 282 338 283 
rect 340 282 341 283 
rect 337 287 338 288 
rect 340 287 341 288 
<< labels >>
rlabel pdiffusion 229 246 230 247  0 t = 1
rlabel pdiffusion 232 246 233 247  0 t = 2
rlabel pdiffusion 229 251 230 252  0 t = 3
rlabel pdiffusion 232 251 233 252  0 t = 4
rlabel pdiffusion 228 246 234 252 0 cell no = 422
<< m1 >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< m2 >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< m2c >>
rect 229 246 230 247 
rect 232 246 233 247 
rect 229 251 230 252 
rect 232 251 233 252 
<< labels >>
rlabel pdiffusion 373 192 374 193  0 t = 1
rlabel pdiffusion 376 192 377 193  0 t = 2
rlabel pdiffusion 373 197 374 198  0 t = 3
rlabel pdiffusion 376 197 377 198  0 t = 4
rlabel pdiffusion 372 192 378 198 0 cell no = 423
<< m1 >>
rect 373 192 374 193 
rect 376 192 377 193 
rect 373 197 374 198 
rect 376 197 377 198 
<< m2 >>
rect 373 192 374 193 
rect 376 192 377 193 
rect 373 197 374 198 
rect 376 197 377 198 
<< m2c >>
rect 373 192 374 193 
rect 376 192 377 193 
rect 373 197 374 198 
rect 376 197 377 198 
<< labels >>
rlabel pdiffusion 373 228 374 229  0 t = 1
rlabel pdiffusion 376 228 377 229  0 t = 2
rlabel pdiffusion 373 233 374 234  0 t = 3
rlabel pdiffusion 376 233 377 234  0 t = 4
rlabel pdiffusion 372 228 378 234 0 cell no = 424
<< m1 >>
rect 373 228 374 229 
rect 376 228 377 229 
rect 373 233 374 234 
rect 376 233 377 234 
<< m2 >>
rect 373 228 374 229 
rect 376 228 377 229 
rect 373 233 374 234 
rect 376 233 377 234 
<< m2c >>
rect 373 228 374 229 
rect 376 228 377 229 
rect 373 233 374 234 
rect 376 233 377 234 
<< labels >>
rlabel pdiffusion 391 336 392 337  0 t = 1
rlabel pdiffusion 394 336 395 337  0 t = 2
rlabel pdiffusion 391 341 392 342  0 t = 3
rlabel pdiffusion 394 341 395 342  0 t = 4
rlabel pdiffusion 390 336 396 342 0 cell no = 425
<< m1 >>
rect 391 336 392 337 
rect 394 336 395 337 
rect 391 341 392 342 
rect 394 341 395 342 
<< m2 >>
rect 391 336 392 337 
rect 394 336 395 337 
rect 391 341 392 342 
rect 394 341 395 342 
<< m2c >>
rect 391 336 392 337 
rect 394 336 395 337 
rect 391 341 392 342 
rect 394 341 395 342 
<< labels >>
rlabel pdiffusion 373 336 374 337  0 t = 1
rlabel pdiffusion 376 336 377 337  0 t = 2
rlabel pdiffusion 373 341 374 342  0 t = 3
rlabel pdiffusion 376 341 377 342  0 t = 4
rlabel pdiffusion 372 336 378 342 0 cell no = 426
<< m1 >>
rect 373 336 374 337 
rect 376 336 377 337 
rect 373 341 374 342 
rect 376 341 377 342 
<< m2 >>
rect 373 336 374 337 
rect 376 336 377 337 
rect 373 341 374 342 
rect 376 341 377 342 
<< m2c >>
rect 373 336 374 337 
rect 376 336 377 337 
rect 373 341 374 342 
rect 376 341 377 342 
<< labels >>
rlabel pdiffusion 49 426 50 427  0 t = 1
rlabel pdiffusion 52 426 53 427  0 t = 2
rlabel pdiffusion 49 431 50 432  0 t = 3
rlabel pdiffusion 52 431 53 432  0 t = 4
rlabel pdiffusion 48 426 54 432 0 cell no = 427
<< m1 >>
rect 49 426 50 427 
rect 52 426 53 427 
rect 49 431 50 432 
rect 52 431 53 432 
<< m2 >>
rect 49 426 50 427 
rect 52 426 53 427 
rect 49 431 50 432 
rect 52 431 53 432 
<< m2c >>
rect 49 426 50 427 
rect 52 426 53 427 
rect 49 431 50 432 
rect 52 431 53 432 
<< labels >>
rlabel pdiffusion 319 318 320 319  0 t = 1
rlabel pdiffusion 322 318 323 319  0 t = 2
rlabel pdiffusion 319 323 320 324  0 t = 3
rlabel pdiffusion 322 323 323 324  0 t = 4
rlabel pdiffusion 318 318 324 324 0 cell no = 428
<< m1 >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< m2 >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< m2c >>
rect 319 318 320 319 
rect 322 318 323 319 
rect 319 323 320 324 
rect 322 323 323 324 
<< labels >>
rlabel pdiffusion 31 282 32 283  0 t = 1
rlabel pdiffusion 34 282 35 283  0 t = 2
rlabel pdiffusion 31 287 32 288  0 t = 3
rlabel pdiffusion 34 287 35 288  0 t = 4
rlabel pdiffusion 30 282 36 288 0 cell no = 429
<< m1 >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< m2 >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< m2c >>
rect 31 282 32 283 
rect 34 282 35 283 
rect 31 287 32 288 
rect 34 287 35 288 
<< labels >>
rlabel pdiffusion 157 30 158 31  0 t = 1
rlabel pdiffusion 160 30 161 31  0 t = 2
rlabel pdiffusion 157 35 158 36  0 t = 3
rlabel pdiffusion 160 35 161 36  0 t = 4
rlabel pdiffusion 156 30 162 36 0 cell no = 430
<< m1 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2 >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< m2c >>
rect 157 30 158 31 
rect 160 30 161 31 
rect 157 35 158 36 
rect 160 35 161 36 
<< labels >>
rlabel pdiffusion 283 426 284 427  0 t = 1
rlabel pdiffusion 286 426 287 427  0 t = 2
rlabel pdiffusion 283 431 284 432  0 t = 3
rlabel pdiffusion 286 431 287 432  0 t = 4
rlabel pdiffusion 282 426 288 432 0 cell no = 431
<< m1 >>
rect 283 426 284 427 
rect 286 426 287 427 
rect 283 431 284 432 
rect 286 431 287 432 
<< m2 >>
rect 283 426 284 427 
rect 286 426 287 427 
rect 283 431 284 432 
rect 286 431 287 432 
<< m2c >>
rect 283 426 284 427 
rect 286 426 287 427 
rect 283 431 284 432 
rect 286 431 287 432 
<< labels >>
rlabel pdiffusion 229 318 230 319  0 t = 1
rlabel pdiffusion 232 318 233 319  0 t = 2
rlabel pdiffusion 229 323 230 324  0 t = 3
rlabel pdiffusion 232 323 233 324  0 t = 4
rlabel pdiffusion 228 318 234 324 0 cell no = 432
<< m1 >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< m2 >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< m2c >>
rect 229 318 230 319 
rect 232 318 233 319 
rect 229 323 230 324 
rect 232 323 233 324 
<< labels >>
rlabel pdiffusion 355 426 356 427  0 t = 1
rlabel pdiffusion 358 426 359 427  0 t = 2
rlabel pdiffusion 355 431 356 432  0 t = 3
rlabel pdiffusion 358 431 359 432  0 t = 4
rlabel pdiffusion 354 426 360 432 0 cell no = 433
<< m1 >>
rect 355 426 356 427 
rect 358 426 359 427 
rect 355 431 356 432 
rect 358 431 359 432 
<< m2 >>
rect 355 426 356 427 
rect 358 426 359 427 
rect 355 431 356 432 
rect 358 431 359 432 
<< m2c >>
rect 355 426 356 427 
rect 358 426 359 427 
rect 355 431 356 432 
rect 358 431 359 432 
<< labels >>
rlabel pdiffusion 211 66 212 67  0 t = 1
rlabel pdiffusion 214 66 215 67  0 t = 2
rlabel pdiffusion 211 71 212 72  0 t = 3
rlabel pdiffusion 214 71 215 72  0 t = 4
rlabel pdiffusion 210 66 216 72 0 cell no = 434
<< m1 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2 >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< m2c >>
rect 211 66 212 67 
rect 214 66 215 67 
rect 211 71 212 72 
rect 214 71 215 72 
<< labels >>
rlabel pdiffusion 49 300 50 301  0 t = 1
rlabel pdiffusion 52 300 53 301  0 t = 2
rlabel pdiffusion 49 305 50 306  0 t = 3
rlabel pdiffusion 52 305 53 306  0 t = 4
rlabel pdiffusion 48 300 54 306 0 cell no = 435
<< m1 >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< m2 >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< m2c >>
rect 49 300 50 301 
rect 52 300 53 301 
rect 49 305 50 306 
rect 52 305 53 306 
<< labels >>
rlabel pdiffusion 103 246 104 247  0 t = 1
rlabel pdiffusion 106 246 107 247  0 t = 2
rlabel pdiffusion 103 251 104 252  0 t = 3
rlabel pdiffusion 106 251 107 252  0 t = 4
rlabel pdiffusion 102 246 108 252 0 cell no = 436
<< m1 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2 >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< m2c >>
rect 103 246 104 247 
rect 106 246 107 247 
rect 103 251 104 252 
rect 106 251 107 252 
<< labels >>
rlabel pdiffusion 247 372 248 373  0 t = 1
rlabel pdiffusion 250 372 251 373  0 t = 2
rlabel pdiffusion 247 377 248 378  0 t = 3
rlabel pdiffusion 250 377 251 378  0 t = 4
rlabel pdiffusion 246 372 252 378 0 cell no = 437
<< m1 >>
rect 247 372 248 373 
rect 250 372 251 373 
rect 247 377 248 378 
rect 250 377 251 378 
<< m2 >>
rect 247 372 248 373 
rect 250 372 251 373 
rect 247 377 248 378 
rect 250 377 251 378 
<< m2c >>
rect 247 372 248 373 
rect 250 372 251 373 
rect 247 377 248 378 
rect 250 377 251 378 
<< labels >>
rlabel pdiffusion 31 390 32 391  0 t = 1
rlabel pdiffusion 34 390 35 391  0 t = 2
rlabel pdiffusion 31 395 32 396  0 t = 3
rlabel pdiffusion 34 395 35 396  0 t = 4
rlabel pdiffusion 30 390 36 396 0 cell no = 438
<< m1 >>
rect 31 390 32 391 
rect 34 390 35 391 
rect 31 395 32 396 
rect 34 395 35 396 
<< m2 >>
rect 31 390 32 391 
rect 34 390 35 391 
rect 31 395 32 396 
rect 34 395 35 396 
<< m2c >>
rect 31 390 32 391 
rect 34 390 35 391 
rect 31 395 32 396 
rect 34 395 35 396 
<< labels >>
rlabel pdiffusion 139 264 140 265  0 t = 1
rlabel pdiffusion 142 264 143 265  0 t = 2
rlabel pdiffusion 139 269 140 270  0 t = 3
rlabel pdiffusion 142 269 143 270  0 t = 4
rlabel pdiffusion 138 264 144 270 0 cell no = 439
<< m1 >>
rect 139 264 140 265 
rect 142 264 143 265 
rect 139 269 140 270 
rect 142 269 143 270 
<< m2 >>
rect 139 264 140 265 
rect 142 264 143 265 
rect 139 269 140 270 
rect 142 269 143 270 
<< m2c >>
rect 139 264 140 265 
rect 142 264 143 265 
rect 139 269 140 270 
rect 142 269 143 270 
<< labels >>
rlabel pdiffusion 31 408 32 409  0 t = 1
rlabel pdiffusion 34 408 35 409  0 t = 2
rlabel pdiffusion 31 413 32 414  0 t = 3
rlabel pdiffusion 34 413 35 414  0 t = 4
rlabel pdiffusion 30 408 36 414 0 cell no = 440
<< m1 >>
rect 31 408 32 409 
rect 34 408 35 409 
rect 31 413 32 414 
rect 34 413 35 414 
<< m2 >>
rect 31 408 32 409 
rect 34 408 35 409 
rect 31 413 32 414 
rect 34 413 35 414 
<< m2c >>
rect 31 408 32 409 
rect 34 408 35 409 
rect 31 413 32 414 
rect 34 413 35 414 
<< labels >>
rlabel pdiffusion 121 300 122 301  0 t = 1
rlabel pdiffusion 124 300 125 301  0 t = 2
rlabel pdiffusion 121 305 122 306  0 t = 3
rlabel pdiffusion 124 305 125 306  0 t = 4
rlabel pdiffusion 120 300 126 306 0 cell no = 441
<< m1 >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< m2 >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< m2c >>
rect 121 300 122 301 
rect 124 300 125 301 
rect 121 305 122 306 
rect 124 305 125 306 
<< labels >>
rlabel pdiffusion 67 156 68 157  0 t = 1
rlabel pdiffusion 70 156 71 157  0 t = 2
rlabel pdiffusion 67 161 68 162  0 t = 3
rlabel pdiffusion 70 161 71 162  0 t = 4
rlabel pdiffusion 66 156 72 162 0 cell no = 442
<< m1 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2 >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< m2c >>
rect 67 156 68 157 
rect 70 156 71 157 
rect 67 161 68 162 
rect 70 161 71 162 
<< labels >>
rlabel pdiffusion 301 174 302 175  0 t = 1
rlabel pdiffusion 304 174 305 175  0 t = 2
rlabel pdiffusion 301 179 302 180  0 t = 3
rlabel pdiffusion 304 179 305 180  0 t = 4
rlabel pdiffusion 300 174 306 180 0 cell no = 443
<< m1 >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< m2 >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< m2c >>
rect 301 174 302 175 
rect 304 174 305 175 
rect 301 179 302 180 
rect 304 179 305 180 
<< labels >>
rlabel pdiffusion 319 498 320 499  0 t = 1
rlabel pdiffusion 322 498 323 499  0 t = 2
rlabel pdiffusion 319 503 320 504  0 t = 3
rlabel pdiffusion 322 503 323 504  0 t = 4
rlabel pdiffusion 318 498 324 504 0 cell no = 444
<< m1 >>
rect 319 498 320 499 
rect 322 498 323 499 
rect 319 503 320 504 
rect 322 503 323 504 
<< m2 >>
rect 319 498 320 499 
rect 322 498 323 499 
rect 319 503 320 504 
rect 322 503 323 504 
<< m2c >>
rect 319 498 320 499 
rect 322 498 323 499 
rect 319 503 320 504 
rect 322 503 323 504 
<< labels >>
rlabel pdiffusion 319 372 320 373  0 t = 1
rlabel pdiffusion 322 372 323 373  0 t = 2
rlabel pdiffusion 319 377 320 378  0 t = 3
rlabel pdiffusion 322 377 323 378  0 t = 4
rlabel pdiffusion 318 372 324 378 0 cell no = 445
<< m1 >>
rect 319 372 320 373 
rect 322 372 323 373 
rect 319 377 320 378 
rect 322 377 323 378 
<< m2 >>
rect 319 372 320 373 
rect 322 372 323 373 
rect 319 377 320 378 
rect 322 377 323 378 
<< m2c >>
rect 319 372 320 373 
rect 322 372 323 373 
rect 319 377 320 378 
rect 322 377 323 378 
<< labels >>
rlabel pdiffusion 121 354 122 355  0 t = 1
rlabel pdiffusion 124 354 125 355  0 t = 2
rlabel pdiffusion 121 359 122 360  0 t = 3
rlabel pdiffusion 124 359 125 360  0 t = 4
rlabel pdiffusion 120 354 126 360 0 cell no = 446
<< m1 >>
rect 121 354 122 355 
rect 124 354 125 355 
rect 121 359 122 360 
rect 124 359 125 360 
<< m2 >>
rect 121 354 122 355 
rect 124 354 125 355 
rect 121 359 122 360 
rect 124 359 125 360 
<< m2c >>
rect 121 354 122 355 
rect 124 354 125 355 
rect 121 359 122 360 
rect 124 359 125 360 
<< labels >>
rlabel pdiffusion 211 426 212 427  0 t = 1
rlabel pdiffusion 214 426 215 427  0 t = 2
rlabel pdiffusion 211 431 212 432  0 t = 3
rlabel pdiffusion 214 431 215 432  0 t = 4
rlabel pdiffusion 210 426 216 432 0 cell no = 447
<< m1 >>
rect 211 426 212 427 
rect 214 426 215 427 
rect 211 431 212 432 
rect 214 431 215 432 
<< m2 >>
rect 211 426 212 427 
rect 214 426 215 427 
rect 211 431 212 432 
rect 214 431 215 432 
<< m2c >>
rect 211 426 212 427 
rect 214 426 215 427 
rect 211 431 212 432 
rect 214 431 215 432 
<< labels >>
rlabel pdiffusion 409 48 410 49  0 t = 1
rlabel pdiffusion 412 48 413 49  0 t = 2
rlabel pdiffusion 409 53 410 54  0 t = 3
rlabel pdiffusion 412 53 413 54  0 t = 4
rlabel pdiffusion 408 48 414 54 0 cell no = 448
<< m1 >>
rect 409 48 410 49 
rect 412 48 413 49 
rect 409 53 410 54 
rect 412 53 413 54 
<< m2 >>
rect 409 48 410 49 
rect 412 48 413 49 
rect 409 53 410 54 
rect 412 53 413 54 
<< m2c >>
rect 409 48 410 49 
rect 412 48 413 49 
rect 409 53 410 54 
rect 412 53 413 54 
<< labels >>
rlabel pdiffusion 337 192 338 193  0 t = 1
rlabel pdiffusion 340 192 341 193  0 t = 2
rlabel pdiffusion 337 197 338 198  0 t = 3
rlabel pdiffusion 340 197 341 198  0 t = 4
rlabel pdiffusion 336 192 342 198 0 cell no = 449
<< m1 >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< m2 >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< m2c >>
rect 337 192 338 193 
rect 340 192 341 193 
rect 337 197 338 198 
rect 340 197 341 198 
<< labels >>
rlabel pdiffusion 121 390 122 391  0 t = 1
rlabel pdiffusion 124 390 125 391  0 t = 2
rlabel pdiffusion 121 395 122 396  0 t = 3
rlabel pdiffusion 124 395 125 396  0 t = 4
rlabel pdiffusion 120 390 126 396 0 cell no = 450
<< m1 >>
rect 121 390 122 391 
rect 124 390 125 391 
rect 121 395 122 396 
rect 124 395 125 396 
<< m2 >>
rect 121 390 122 391 
rect 124 390 125 391 
rect 121 395 122 396 
rect 124 395 125 396 
<< m2c >>
rect 121 390 122 391 
rect 124 390 125 391 
rect 121 395 122 396 
rect 124 395 125 396 
<< labels >>
rlabel pdiffusion 31 30 32 31  0 t = 1
rlabel pdiffusion 34 30 35 31  0 t = 2
rlabel pdiffusion 31 35 32 36  0 t = 3
rlabel pdiffusion 34 35 35 36  0 t = 4
rlabel pdiffusion 30 30 36 36 0 cell no = 451
<< m1 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2 >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< m2c >>
rect 31 30 32 31 
rect 34 30 35 31 
rect 31 35 32 36 
rect 34 35 35 36 
<< labels >>
rlabel pdiffusion 247 444 248 445  0 t = 1
rlabel pdiffusion 250 444 251 445  0 t = 2
rlabel pdiffusion 247 449 248 450  0 t = 3
rlabel pdiffusion 250 449 251 450  0 t = 4
rlabel pdiffusion 246 444 252 450 0 cell no = 452
<< m1 >>
rect 247 444 248 445 
rect 250 444 251 445 
rect 247 449 248 450 
rect 250 449 251 450 
<< m2 >>
rect 247 444 248 445 
rect 250 444 251 445 
rect 247 449 248 450 
rect 250 449 251 450 
<< m2c >>
rect 247 444 248 445 
rect 250 444 251 445 
rect 247 449 248 450 
rect 250 449 251 450 
<< labels >>
rlabel pdiffusion 211 192 212 193  0 t = 1
rlabel pdiffusion 214 192 215 193  0 t = 2
rlabel pdiffusion 211 197 212 198  0 t = 3
rlabel pdiffusion 214 197 215 198  0 t = 4
rlabel pdiffusion 210 192 216 198 0 cell no = 453
<< m1 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2 >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< m2c >>
rect 211 192 212 193 
rect 214 192 215 193 
rect 211 197 212 198 
rect 214 197 215 198 
<< labels >>
rlabel pdiffusion 427 210 428 211  0 t = 1
rlabel pdiffusion 430 210 431 211  0 t = 2
rlabel pdiffusion 427 215 428 216  0 t = 3
rlabel pdiffusion 430 215 431 216  0 t = 4
rlabel pdiffusion 426 210 432 216 0 cell no = 454
<< m1 >>
rect 427 210 428 211 
rect 430 210 431 211 
rect 427 215 428 216 
rect 430 215 431 216 
<< m2 >>
rect 427 210 428 211 
rect 430 210 431 211 
rect 427 215 428 216 
rect 430 215 431 216 
<< m2c >>
rect 427 210 428 211 
rect 430 210 431 211 
rect 427 215 428 216 
rect 430 215 431 216 
<< labels >>
rlabel pdiffusion 175 102 176 103  0 t = 1
rlabel pdiffusion 178 102 179 103  0 t = 2
rlabel pdiffusion 175 107 176 108  0 t = 3
rlabel pdiffusion 178 107 179 108  0 t = 4
rlabel pdiffusion 174 102 180 108 0 cell no = 455
<< m1 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2 >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< m2c >>
rect 175 102 176 103 
rect 178 102 179 103 
rect 175 107 176 108 
rect 178 107 179 108 
<< labels >>
rlabel pdiffusion 373 264 374 265  0 t = 1
rlabel pdiffusion 376 264 377 265  0 t = 2
rlabel pdiffusion 373 269 374 270  0 t = 3
rlabel pdiffusion 376 269 377 270  0 t = 4
rlabel pdiffusion 372 264 378 270 0 cell no = 456
<< m1 >>
rect 373 264 374 265 
rect 376 264 377 265 
rect 373 269 374 270 
rect 376 269 377 270 
<< m2 >>
rect 373 264 374 265 
rect 376 264 377 265 
rect 373 269 374 270 
rect 376 269 377 270 
<< m2c >>
rect 373 264 374 265 
rect 376 264 377 265 
rect 373 269 374 270 
rect 376 269 377 270 
<< labels >>
rlabel pdiffusion 139 246 140 247  0 t = 1
rlabel pdiffusion 142 246 143 247  0 t = 2
rlabel pdiffusion 139 251 140 252  0 t = 3
rlabel pdiffusion 142 251 143 252  0 t = 4
rlabel pdiffusion 138 246 144 252 0 cell no = 457
<< m1 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2 >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< m2c >>
rect 139 246 140 247 
rect 142 246 143 247 
rect 139 251 140 252 
rect 142 251 143 252 
<< labels >>
rlabel pdiffusion 481 300 482 301  0 t = 1
rlabel pdiffusion 484 300 485 301  0 t = 2
rlabel pdiffusion 481 305 482 306  0 t = 3
rlabel pdiffusion 484 305 485 306  0 t = 4
rlabel pdiffusion 480 300 486 306 0 cell no = 458
<< m1 >>
rect 481 300 482 301 
rect 484 300 485 301 
rect 481 305 482 306 
rect 484 305 485 306 
<< m2 >>
rect 481 300 482 301 
rect 484 300 485 301 
rect 481 305 482 306 
rect 484 305 485 306 
<< m2c >>
rect 481 300 482 301 
rect 484 300 485 301 
rect 481 305 482 306 
rect 484 305 485 306 
<< labels >>
rlabel pdiffusion 463 318 464 319  0 t = 1
rlabel pdiffusion 466 318 467 319  0 t = 2
rlabel pdiffusion 463 323 464 324  0 t = 3
rlabel pdiffusion 466 323 467 324  0 t = 4
rlabel pdiffusion 462 318 468 324 0 cell no = 459
<< m1 >>
rect 463 318 464 319 
rect 466 318 467 319 
rect 463 323 464 324 
rect 466 323 467 324 
<< m2 >>
rect 463 318 464 319 
rect 466 318 467 319 
rect 463 323 464 324 
rect 466 323 467 324 
<< m2c >>
rect 463 318 464 319 
rect 466 318 467 319 
rect 463 323 464 324 
rect 466 323 467 324 
<< labels >>
rlabel pdiffusion 499 246 500 247  0 t = 1
rlabel pdiffusion 502 246 503 247  0 t = 2
rlabel pdiffusion 499 251 500 252  0 t = 3
rlabel pdiffusion 502 251 503 252  0 t = 4
rlabel pdiffusion 498 246 504 252 0 cell no = 460
<< m1 >>
rect 499 246 500 247 
rect 502 246 503 247 
rect 499 251 500 252 
rect 502 251 503 252 
<< m2 >>
rect 499 246 500 247 
rect 502 246 503 247 
rect 499 251 500 252 
rect 502 251 503 252 
<< m2c >>
rect 499 246 500 247 
rect 502 246 503 247 
rect 499 251 500 252 
rect 502 251 503 252 
<< labels >>
rlabel pdiffusion 463 372 464 373  0 t = 1
rlabel pdiffusion 466 372 467 373  0 t = 2
rlabel pdiffusion 463 377 464 378  0 t = 3
rlabel pdiffusion 466 377 467 378  0 t = 4
rlabel pdiffusion 462 372 468 378 0 cell no = 461
<< m1 >>
rect 463 372 464 373 
rect 466 372 467 373 
rect 463 377 464 378 
rect 466 377 467 378 
<< m2 >>
rect 463 372 464 373 
rect 466 372 467 373 
rect 463 377 464 378 
rect 466 377 467 378 
<< m2c >>
rect 463 372 464 373 
rect 466 372 467 373 
rect 463 377 464 378 
rect 466 377 467 378 
<< labels >>
rlabel pdiffusion 499 282 500 283  0 t = 1
rlabel pdiffusion 502 282 503 283  0 t = 2
rlabel pdiffusion 499 287 500 288  0 t = 3
rlabel pdiffusion 502 287 503 288  0 t = 4
rlabel pdiffusion 498 282 504 288 0 cell no = 462
<< m1 >>
rect 499 282 500 283 
rect 502 282 503 283 
rect 499 287 500 288 
rect 502 287 503 288 
<< m2 >>
rect 499 282 500 283 
rect 502 282 503 283 
rect 499 287 500 288 
rect 502 287 503 288 
<< m2c >>
rect 499 282 500 283 
rect 502 282 503 283 
rect 499 287 500 288 
rect 502 287 503 288 
<< labels >>
rlabel pdiffusion 499 318 500 319  0 t = 1
rlabel pdiffusion 502 318 503 319  0 t = 2
rlabel pdiffusion 499 323 500 324  0 t = 3
rlabel pdiffusion 502 323 503 324  0 t = 4
rlabel pdiffusion 498 318 504 324 0 cell no = 463
<< m1 >>
rect 499 318 500 319 
rect 502 318 503 319 
rect 499 323 500 324 
rect 502 323 503 324 
<< m2 >>
rect 499 318 500 319 
rect 502 318 503 319 
rect 499 323 500 324 
rect 502 323 503 324 
<< m2c >>
rect 499 318 500 319 
rect 502 318 503 319 
rect 499 323 500 324 
rect 502 323 503 324 
<< labels >>
rlabel pdiffusion 481 498 482 499  0 t = 1
rlabel pdiffusion 484 498 485 499  0 t = 2
rlabel pdiffusion 481 503 482 504  0 t = 3
rlabel pdiffusion 484 503 485 504  0 t = 4
rlabel pdiffusion 480 498 486 504 0 cell no = 464
<< m1 >>
rect 481 498 482 499 
rect 484 498 485 499 
rect 481 503 482 504 
rect 484 503 485 504 
<< m2 >>
rect 481 498 482 499 
rect 484 498 485 499 
rect 481 503 482 504 
rect 484 503 485 504 
<< m2c >>
rect 481 498 482 499 
rect 484 498 485 499 
rect 481 503 482 504 
rect 484 503 485 504 
<< labels >>
rlabel pdiffusion 85 102 86 103  0 t = 1
rlabel pdiffusion 88 102 89 103  0 t = 2
rlabel pdiffusion 85 107 86 108  0 t = 3
rlabel pdiffusion 88 107 89 108  0 t = 4
rlabel pdiffusion 84 102 90 108 0 cell no = 465
<< m1 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2 >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< m2c >>
rect 85 102 86 103 
rect 88 102 89 103 
rect 85 107 86 108 
rect 88 107 89 108 
<< labels >>
rlabel pdiffusion 103 300 104 301  0 t = 1
rlabel pdiffusion 106 300 107 301  0 t = 2
rlabel pdiffusion 103 305 104 306  0 t = 3
rlabel pdiffusion 106 305 107 306  0 t = 4
rlabel pdiffusion 102 300 108 306 0 cell no = 466
<< m1 >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< m2 >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< m2c >>
rect 103 300 104 301 
rect 106 300 107 301 
rect 103 305 104 306 
rect 106 305 107 306 
<< labels >>
rlabel pdiffusion 103 408 104 409  0 t = 1
rlabel pdiffusion 106 408 107 409  0 t = 2
rlabel pdiffusion 103 413 104 414  0 t = 3
rlabel pdiffusion 106 413 107 414  0 t = 4
rlabel pdiffusion 102 408 108 414 0 cell no = 467
<< m1 >>
rect 103 408 104 409 
rect 106 408 107 409 
rect 103 413 104 414 
rect 106 413 107 414 
<< m2 >>
rect 103 408 104 409 
rect 106 408 107 409 
rect 103 413 104 414 
rect 106 413 107 414 
<< m2c >>
rect 103 408 104 409 
rect 106 408 107 409 
rect 103 413 104 414 
rect 106 413 107 414 
<< labels >>
rlabel pdiffusion 85 228 86 229  0 t = 1
rlabel pdiffusion 88 228 89 229  0 t = 2
rlabel pdiffusion 85 233 86 234  0 t = 3
rlabel pdiffusion 88 233 89 234  0 t = 4
rlabel pdiffusion 84 228 90 234 0 cell no = 468
<< m1 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2 >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< m2c >>
rect 85 228 86 229 
rect 88 228 89 229 
rect 85 233 86 234 
rect 88 233 89 234 
<< labels >>
rlabel pdiffusion 67 462 68 463  0 t = 1
rlabel pdiffusion 70 462 71 463  0 t = 2
rlabel pdiffusion 67 467 68 468  0 t = 3
rlabel pdiffusion 70 467 71 468  0 t = 4
rlabel pdiffusion 66 462 72 468 0 cell no = 469
<< m1 >>
rect 67 462 68 463 
rect 70 462 71 463 
rect 67 467 68 468 
rect 70 467 71 468 
<< m2 >>
rect 67 462 68 463 
rect 70 462 71 463 
rect 67 467 68 468 
rect 70 467 71 468 
<< m2c >>
rect 67 462 68 463 
rect 70 462 71 463 
rect 67 467 68 468 
rect 70 467 71 468 
<< labels >>
rlabel pdiffusion 193 30 194 31  0 t = 1
rlabel pdiffusion 196 30 197 31  0 t = 2
rlabel pdiffusion 193 35 194 36  0 t = 3
rlabel pdiffusion 196 35 197 36  0 t = 4
rlabel pdiffusion 192 30 198 36 0 cell no = 470
<< m1 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2 >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< m2c >>
rect 193 30 194 31 
rect 196 30 197 31 
rect 193 35 194 36 
rect 196 35 197 36 
<< labels >>
rlabel pdiffusion 139 480 140 481  0 t = 1
rlabel pdiffusion 142 480 143 481  0 t = 2
rlabel pdiffusion 139 485 140 486  0 t = 3
rlabel pdiffusion 142 485 143 486  0 t = 4
rlabel pdiffusion 138 480 144 486 0 cell no = 471
<< m1 >>
rect 139 480 140 481 
rect 142 480 143 481 
rect 139 485 140 486 
rect 142 485 143 486 
<< m2 >>
rect 139 480 140 481 
rect 142 480 143 481 
rect 139 485 140 486 
rect 142 485 143 486 
<< m2c >>
rect 139 480 140 481 
rect 142 480 143 481 
rect 139 485 140 486 
rect 142 485 143 486 
<< labels >>
rlabel pdiffusion 139 318 140 319  0 t = 1
rlabel pdiffusion 142 318 143 319  0 t = 2
rlabel pdiffusion 139 323 140 324  0 t = 3
rlabel pdiffusion 142 323 143 324  0 t = 4
rlabel pdiffusion 138 318 144 324 0 cell no = 472
<< m1 >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< m2 >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< m2c >>
rect 139 318 140 319 
rect 142 318 143 319 
rect 139 323 140 324 
rect 142 323 143 324 
<< labels >>
rlabel pdiffusion 283 84 284 85  0 t = 1
rlabel pdiffusion 286 84 287 85  0 t = 2
rlabel pdiffusion 283 89 284 90  0 t = 3
rlabel pdiffusion 286 89 287 90  0 t = 4
rlabel pdiffusion 282 84 288 90 0 cell no = 473
<< m1 >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< m2 >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< m2c >>
rect 283 84 284 85 
rect 286 84 287 85 
rect 283 89 284 90 
rect 286 89 287 90 
<< labels >>
rlabel pdiffusion 175 282 176 283  0 t = 1
rlabel pdiffusion 178 282 179 283  0 t = 2
rlabel pdiffusion 175 287 176 288  0 t = 3
rlabel pdiffusion 178 287 179 288  0 t = 4
rlabel pdiffusion 174 282 180 288 0 cell no = 474
<< m1 >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< m2 >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< m2c >>
rect 175 282 176 283 
rect 178 282 179 283 
rect 175 287 176 288 
rect 178 287 179 288 
<< labels >>
rlabel pdiffusion 247 318 248 319  0 t = 1
rlabel pdiffusion 250 318 251 319  0 t = 2
rlabel pdiffusion 247 323 248 324  0 t = 3
rlabel pdiffusion 250 323 251 324  0 t = 4
rlabel pdiffusion 246 318 252 324 0 cell no = 475
<< m1 >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< m2 >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< m2c >>
rect 247 318 248 319 
rect 250 318 251 319 
rect 247 323 248 324 
rect 250 323 251 324 
<< labels >>
rlabel pdiffusion 301 318 302 319  0 t = 1
rlabel pdiffusion 304 318 305 319  0 t = 2
rlabel pdiffusion 301 323 302 324  0 t = 3
rlabel pdiffusion 304 323 305 324  0 t = 4
rlabel pdiffusion 300 318 306 324 0 cell no = 476
<< m1 >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< m2 >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< m2c >>
rect 301 318 302 319 
rect 304 318 305 319 
rect 301 323 302 324 
rect 304 323 305 324 
<< labels >>
rlabel pdiffusion 445 228 446 229  0 t = 1
rlabel pdiffusion 448 228 449 229  0 t = 2
rlabel pdiffusion 445 233 446 234  0 t = 3
rlabel pdiffusion 448 233 449 234  0 t = 4
rlabel pdiffusion 444 228 450 234 0 cell no = 477
<< m1 >>
rect 445 228 446 229 
rect 448 228 449 229 
rect 445 233 446 234 
rect 448 233 449 234 
<< m2 >>
rect 445 228 446 229 
rect 448 228 449 229 
rect 445 233 446 234 
rect 448 233 449 234 
<< m2c >>
rect 445 228 446 229 
rect 448 228 449 229 
rect 445 233 446 234 
rect 448 233 449 234 
<< labels >>
rlabel pdiffusion 211 174 212 175  0 t = 1
rlabel pdiffusion 214 174 215 175  0 t = 2
rlabel pdiffusion 211 179 212 180  0 t = 3
rlabel pdiffusion 214 179 215 180  0 t = 4
rlabel pdiffusion 210 174 216 180 0 cell no = 478
<< m1 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2 >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< m2c >>
rect 211 174 212 175 
rect 214 174 215 175 
rect 211 179 212 180 
rect 214 179 215 180 
<< labels >>
rlabel pdiffusion 175 228 176 229  0 t = 1
rlabel pdiffusion 178 228 179 229  0 t = 2
rlabel pdiffusion 175 233 176 234  0 t = 3
rlabel pdiffusion 178 233 179 234  0 t = 4
rlabel pdiffusion 174 228 180 234 0 cell no = 479
<< m1 >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< m2 >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< m2c >>
rect 175 228 176 229 
rect 178 228 179 229 
rect 175 233 176 234 
rect 178 233 179 234 
<< labels >>
rlabel pdiffusion 229 426 230 427  0 t = 1
rlabel pdiffusion 232 426 233 427  0 t = 2
rlabel pdiffusion 229 431 230 432  0 t = 3
rlabel pdiffusion 232 431 233 432  0 t = 4
rlabel pdiffusion 228 426 234 432 0 cell no = 480
<< m1 >>
rect 229 426 230 427 
rect 232 426 233 427 
rect 229 431 230 432 
rect 232 431 233 432 
<< m2 >>
rect 229 426 230 427 
rect 232 426 233 427 
rect 229 431 230 432 
rect 232 431 233 432 
<< m2c >>
rect 229 426 230 427 
rect 232 426 233 427 
rect 229 431 230 432 
rect 232 431 233 432 
<< labels >>
rlabel pdiffusion 409 300 410 301  0 t = 1
rlabel pdiffusion 412 300 413 301  0 t = 2
rlabel pdiffusion 409 305 410 306  0 t = 3
rlabel pdiffusion 412 305 413 306  0 t = 4
rlabel pdiffusion 408 300 414 306 0 cell no = 481
<< m1 >>
rect 409 300 410 301 
rect 412 300 413 301 
rect 409 305 410 306 
rect 412 305 413 306 
<< m2 >>
rect 409 300 410 301 
rect 412 300 413 301 
rect 409 305 410 306 
rect 412 305 413 306 
<< m2c >>
rect 409 300 410 301 
rect 412 300 413 301 
rect 409 305 410 306 
rect 412 305 413 306 
<< labels >>
rlabel pdiffusion 409 246 410 247  0 t = 1
rlabel pdiffusion 412 246 413 247  0 t = 2
rlabel pdiffusion 409 251 410 252  0 t = 3
rlabel pdiffusion 412 251 413 252  0 t = 4
rlabel pdiffusion 408 246 414 252 0 cell no = 482
<< m1 >>
rect 409 246 410 247 
rect 412 246 413 247 
rect 409 251 410 252 
rect 412 251 413 252 
<< m2 >>
rect 409 246 410 247 
rect 412 246 413 247 
rect 409 251 410 252 
rect 412 251 413 252 
<< m2c >>
rect 409 246 410 247 
rect 412 246 413 247 
rect 409 251 410 252 
rect 412 251 413 252 
<< labels >>
rlabel pdiffusion 499 300 500 301  0 t = 1
rlabel pdiffusion 502 300 503 301  0 t = 2
rlabel pdiffusion 499 305 500 306  0 t = 3
rlabel pdiffusion 502 305 503 306  0 t = 4
rlabel pdiffusion 498 300 504 306 0 cell no = 483
<< m1 >>
rect 499 300 500 301 
rect 502 300 503 301 
rect 499 305 500 306 
rect 502 305 503 306 
<< m2 >>
rect 499 300 500 301 
rect 502 300 503 301 
rect 499 305 500 306 
rect 502 305 503 306 
<< m2c >>
rect 499 300 500 301 
rect 502 300 503 301 
rect 499 305 500 306 
rect 502 305 503 306 
<< labels >>
rlabel pdiffusion 445 84 446 85  0 t = 1
rlabel pdiffusion 448 84 449 85  0 t = 2
rlabel pdiffusion 445 89 446 90  0 t = 3
rlabel pdiffusion 448 89 449 90  0 t = 4
rlabel pdiffusion 444 84 450 90 0 cell no = 484
<< m1 >>
rect 445 84 446 85 
rect 448 84 449 85 
rect 445 89 446 90 
rect 448 89 449 90 
<< m2 >>
rect 445 84 446 85 
rect 448 84 449 85 
rect 445 89 446 90 
rect 448 89 449 90 
<< m2c >>
rect 445 84 446 85 
rect 448 84 449 85 
rect 445 89 446 90 
rect 448 89 449 90 
<< labels >>
rlabel pdiffusion 463 408 464 409  0 t = 1
rlabel pdiffusion 466 408 467 409  0 t = 2
rlabel pdiffusion 463 413 464 414  0 t = 3
rlabel pdiffusion 466 413 467 414  0 t = 4
rlabel pdiffusion 462 408 468 414 0 cell no = 485
<< m1 >>
rect 463 408 464 409 
rect 466 408 467 409 
rect 463 413 464 414 
rect 466 413 467 414 
<< m2 >>
rect 463 408 464 409 
rect 466 408 467 409 
rect 463 413 464 414 
rect 466 413 467 414 
<< m2c >>
rect 463 408 464 409 
rect 466 408 467 409 
rect 463 413 464 414 
rect 466 413 467 414 
<< labels >>
rlabel pdiffusion 373 300 374 301  0 t = 1
rlabel pdiffusion 376 300 377 301  0 t = 2
rlabel pdiffusion 373 305 374 306  0 t = 3
rlabel pdiffusion 376 305 377 306  0 t = 4
rlabel pdiffusion 372 300 378 306 0 cell no = 486
<< m1 >>
rect 373 300 374 301 
rect 376 300 377 301 
rect 373 305 374 306 
rect 376 305 377 306 
<< m2 >>
rect 373 300 374 301 
rect 376 300 377 301 
rect 373 305 374 306 
rect 376 305 377 306 
<< m2c >>
rect 373 300 374 301 
rect 376 300 377 301 
rect 373 305 374 306 
rect 376 305 377 306 
<< labels >>
rlabel pdiffusion 463 336 464 337  0 t = 1
rlabel pdiffusion 466 336 467 337  0 t = 2
rlabel pdiffusion 463 341 464 342  0 t = 3
rlabel pdiffusion 466 341 467 342  0 t = 4
rlabel pdiffusion 462 336 468 342 0 cell no = 487
<< m1 >>
rect 463 336 464 337 
rect 466 336 467 337 
rect 463 341 464 342 
rect 466 341 467 342 
<< m2 >>
rect 463 336 464 337 
rect 466 336 467 337 
rect 463 341 464 342 
rect 466 341 467 342 
<< m2c >>
rect 463 336 464 337 
rect 466 336 467 337 
rect 463 341 464 342 
rect 466 341 467 342 
<< labels >>
rlabel pdiffusion 445 372 446 373  0 t = 1
rlabel pdiffusion 448 372 449 373  0 t = 2
rlabel pdiffusion 445 377 446 378  0 t = 3
rlabel pdiffusion 448 377 449 378  0 t = 4
rlabel pdiffusion 444 372 450 378 0 cell no = 488
<< m1 >>
rect 445 372 446 373 
rect 448 372 449 373 
rect 445 377 446 378 
rect 448 377 449 378 
<< m2 >>
rect 445 372 446 373 
rect 448 372 449 373 
rect 445 377 446 378 
rect 448 377 449 378 
<< m2c >>
rect 445 372 446 373 
rect 448 372 449 373 
rect 445 377 446 378 
rect 448 377 449 378 
<< labels >>
rlabel pdiffusion 445 246 446 247  0 t = 1
rlabel pdiffusion 448 246 449 247  0 t = 2
rlabel pdiffusion 445 251 446 252  0 t = 3
rlabel pdiffusion 448 251 449 252  0 t = 4
rlabel pdiffusion 444 246 450 252 0 cell no = 489
<< m1 >>
rect 445 246 446 247 
rect 448 246 449 247 
rect 445 251 446 252 
rect 448 251 449 252 
<< m2 >>
rect 445 246 446 247 
rect 448 246 449 247 
rect 445 251 446 252 
rect 448 251 449 252 
<< m2c >>
rect 445 246 446 247 
rect 448 246 449 247 
rect 445 251 446 252 
rect 448 251 449 252 
<< labels >>
rlabel pdiffusion 247 246 248 247  0 t = 1
rlabel pdiffusion 250 246 251 247  0 t = 2
rlabel pdiffusion 247 251 248 252  0 t = 3
rlabel pdiffusion 250 251 251 252  0 t = 4
rlabel pdiffusion 246 246 252 252 0 cell no = 490
<< m1 >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< m2 >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< m2c >>
rect 247 246 248 247 
rect 250 246 251 247 
rect 247 251 248 252 
rect 250 251 251 252 
<< labels >>
rlabel pdiffusion 409 156 410 157  0 t = 1
rlabel pdiffusion 412 156 413 157  0 t = 2
rlabel pdiffusion 409 161 410 162  0 t = 3
rlabel pdiffusion 412 161 413 162  0 t = 4
rlabel pdiffusion 408 156 414 162 0 cell no = 491
<< m1 >>
rect 409 156 410 157 
rect 412 156 413 157 
rect 409 161 410 162 
rect 412 161 413 162 
<< m2 >>
rect 409 156 410 157 
rect 412 156 413 157 
rect 409 161 410 162 
rect 412 161 413 162 
<< m2c >>
rect 409 156 410 157 
rect 412 156 413 157 
rect 409 161 410 162 
rect 412 161 413 162 
<< labels >>
rlabel pdiffusion 373 246 374 247  0 t = 1
rlabel pdiffusion 376 246 377 247  0 t = 2
rlabel pdiffusion 373 251 374 252  0 t = 3
rlabel pdiffusion 376 251 377 252  0 t = 4
rlabel pdiffusion 372 246 378 252 0 cell no = 492
<< m1 >>
rect 373 246 374 247 
rect 376 246 377 247 
rect 373 251 374 252 
rect 376 251 377 252 
<< m2 >>
rect 373 246 374 247 
rect 376 246 377 247 
rect 373 251 374 252 
rect 376 251 377 252 
<< m2c >>
rect 373 246 374 247 
rect 376 246 377 247 
rect 373 251 374 252 
rect 376 251 377 252 
<< labels >>
rlabel pdiffusion 301 390 302 391  0 t = 1
rlabel pdiffusion 304 390 305 391  0 t = 2
rlabel pdiffusion 301 395 302 396  0 t = 3
rlabel pdiffusion 304 395 305 396  0 t = 4
rlabel pdiffusion 300 390 306 396 0 cell no = 493
<< m1 >>
rect 301 390 302 391 
rect 304 390 305 391 
rect 301 395 302 396 
rect 304 395 305 396 
<< m2 >>
rect 301 390 302 391 
rect 304 390 305 391 
rect 301 395 302 396 
rect 304 395 305 396 
<< m2c >>
rect 301 390 302 391 
rect 304 390 305 391 
rect 301 395 302 396 
rect 304 395 305 396 
<< labels >>
rlabel pdiffusion 355 462 356 463  0 t = 1
rlabel pdiffusion 358 462 359 463  0 t = 2
rlabel pdiffusion 355 467 356 468  0 t = 3
rlabel pdiffusion 358 467 359 468  0 t = 4
rlabel pdiffusion 354 462 360 468 0 cell no = 494
<< m1 >>
rect 355 462 356 463 
rect 358 462 359 463 
rect 355 467 356 468 
rect 358 467 359 468 
<< m2 >>
rect 355 462 356 463 
rect 358 462 359 463 
rect 355 467 356 468 
rect 358 467 359 468 
<< m2c >>
rect 355 462 356 463 
rect 358 462 359 463 
rect 355 467 356 468 
rect 358 467 359 468 
<< labels >>
rlabel pdiffusion 121 282 122 283  0 t = 1
rlabel pdiffusion 124 282 125 283  0 t = 2
rlabel pdiffusion 121 287 122 288  0 t = 3
rlabel pdiffusion 124 287 125 288  0 t = 4
rlabel pdiffusion 120 282 126 288 0 cell no = 495
<< m1 >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< m2 >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< m2c >>
rect 121 282 122 283 
rect 124 282 125 283 
rect 121 287 122 288 
rect 124 287 125 288 
<< labels >>
rlabel pdiffusion 139 498 140 499  0 t = 1
rlabel pdiffusion 142 498 143 499  0 t = 2
rlabel pdiffusion 139 503 140 504  0 t = 3
rlabel pdiffusion 142 503 143 504  0 t = 4
rlabel pdiffusion 138 498 144 504 0 cell no = 496
<< m1 >>
rect 139 498 140 499 
rect 142 498 143 499 
rect 139 503 140 504 
rect 142 503 143 504 
<< m2 >>
rect 139 498 140 499 
rect 142 498 143 499 
rect 139 503 140 504 
rect 142 503 143 504 
<< m2c >>
rect 139 498 140 499 
rect 142 498 143 499 
rect 139 503 140 504 
rect 142 503 143 504 
<< labels >>
rlabel pdiffusion 49 462 50 463  0 t = 1
rlabel pdiffusion 52 462 53 463  0 t = 2
rlabel pdiffusion 49 467 50 468  0 t = 3
rlabel pdiffusion 52 467 53 468  0 t = 4
rlabel pdiffusion 48 462 54 468 0 cell no = 497
<< m1 >>
rect 49 462 50 463 
rect 52 462 53 463 
rect 49 467 50 468 
rect 52 467 53 468 
<< m2 >>
rect 49 462 50 463 
rect 52 462 53 463 
rect 49 467 50 468 
rect 52 467 53 468 
<< m2c >>
rect 49 462 50 463 
rect 52 462 53 463 
rect 49 467 50 468 
rect 52 467 53 468 
<< labels >>
rlabel pdiffusion 319 192 320 193  0 t = 1
rlabel pdiffusion 322 192 323 193  0 t = 2
rlabel pdiffusion 319 197 320 198  0 t = 3
rlabel pdiffusion 322 197 323 198  0 t = 4
rlabel pdiffusion 318 192 324 198 0 cell no = 498
<< m1 >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< m2 >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< m2c >>
rect 319 192 320 193 
rect 322 192 323 193 
rect 319 197 320 198 
rect 322 197 323 198 
<< labels >>
rlabel pdiffusion 13 462 14 463  0 t = 1
rlabel pdiffusion 16 462 17 463  0 t = 2
rlabel pdiffusion 13 467 14 468  0 t = 3
rlabel pdiffusion 16 467 17 468  0 t = 4
rlabel pdiffusion 12 462 18 468 0 cell no = 499
<< m1 >>
rect 13 462 14 463 
rect 16 462 17 463 
rect 13 467 14 468 
rect 16 467 17 468 
<< m2 >>
rect 13 462 14 463 
rect 16 462 17 463 
rect 13 467 14 468 
rect 16 467 17 468 
<< m2c >>
rect 13 462 14 463 
rect 16 462 17 463 
rect 13 467 14 468 
rect 16 467 17 468 
<< labels >>
rlabel pdiffusion 31 426 32 427  0 t = 1
rlabel pdiffusion 34 426 35 427  0 t = 2
rlabel pdiffusion 31 431 32 432  0 t = 3
rlabel pdiffusion 34 431 35 432  0 t = 4
rlabel pdiffusion 30 426 36 432 0 cell no = 500
<< m1 >>
rect 31 426 32 427 
rect 34 426 35 427 
rect 31 431 32 432 
rect 34 431 35 432 
<< m2 >>
rect 31 426 32 427 
rect 34 426 35 427 
rect 31 431 32 432 
rect 34 431 35 432 
<< m2c >>
rect 31 426 32 427 
rect 34 426 35 427 
rect 31 431 32 432 
rect 34 431 35 432 
<< labels >>
rlabel pdiffusion 85 318 86 319  0 t = 1
rlabel pdiffusion 88 318 89 319  0 t = 2
rlabel pdiffusion 85 323 86 324  0 t = 3
rlabel pdiffusion 88 323 89 324  0 t = 4
rlabel pdiffusion 84 318 90 324 0 cell no = 501
<< m1 >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< m2 >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< m2c >>
rect 85 318 86 319 
rect 88 318 89 319 
rect 85 323 86 324 
rect 88 323 89 324 
<< labels >>
rlabel pdiffusion 67 210 68 211  0 t = 1
rlabel pdiffusion 70 210 71 211  0 t = 2
rlabel pdiffusion 67 215 68 216  0 t = 3
rlabel pdiffusion 70 215 71 216  0 t = 4
rlabel pdiffusion 66 210 72 216 0 cell no = 502
<< m1 >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< m2 >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< m2c >>
rect 67 210 68 211 
rect 70 210 71 211 
rect 67 215 68 216 
rect 70 215 71 216 
<< labels >>
rlabel pdiffusion 157 372 158 373  0 t = 1
rlabel pdiffusion 160 372 161 373  0 t = 2
rlabel pdiffusion 157 377 158 378  0 t = 3
rlabel pdiffusion 160 377 161 378  0 t = 4
rlabel pdiffusion 156 372 162 378 0 cell no = 503
<< m1 >>
rect 157 372 158 373 
rect 160 372 161 373 
rect 157 377 158 378 
rect 160 377 161 378 
<< m2 >>
rect 157 372 158 373 
rect 160 372 161 373 
rect 157 377 158 378 
rect 160 377 161 378 
<< m2c >>
rect 157 372 158 373 
rect 160 372 161 373 
rect 157 377 158 378 
rect 160 377 161 378 
<< labels >>
rlabel pdiffusion 355 156 356 157  0 t = 1
rlabel pdiffusion 358 156 359 157  0 t = 2
rlabel pdiffusion 355 161 356 162  0 t = 3
rlabel pdiffusion 358 161 359 162  0 t = 4
rlabel pdiffusion 354 156 360 162 0 cell no = 504
<< m1 >>
rect 355 156 356 157 
rect 358 156 359 157 
rect 355 161 356 162 
rect 358 161 359 162 
<< m2 >>
rect 355 156 356 157 
rect 358 156 359 157 
rect 355 161 356 162 
rect 358 161 359 162 
<< m2c >>
rect 355 156 356 157 
rect 358 156 359 157 
rect 355 161 356 162 
rect 358 161 359 162 
<< labels >>
rlabel pdiffusion 13 318 14 319  0 t = 1
rlabel pdiffusion 16 318 17 319  0 t = 2
rlabel pdiffusion 13 323 14 324  0 t = 3
rlabel pdiffusion 16 323 17 324  0 t = 4
rlabel pdiffusion 12 318 18 324 0 cell no = 505
<< m1 >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< m2 >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< m2c >>
rect 13 318 14 319 
rect 16 318 17 319 
rect 13 323 14 324 
rect 16 323 17 324 
<< labels >>
rlabel pdiffusion 85 120 86 121  0 t = 1
rlabel pdiffusion 88 120 89 121  0 t = 2
rlabel pdiffusion 85 125 86 126  0 t = 3
rlabel pdiffusion 88 125 89 126  0 t = 4
rlabel pdiffusion 84 120 90 126 0 cell no = 506
<< m1 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2 >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< m2c >>
rect 85 120 86 121 
rect 88 120 89 121 
rect 85 125 86 126 
rect 88 125 89 126 
<< labels >>
rlabel pdiffusion 427 336 428 337  0 t = 1
rlabel pdiffusion 430 336 431 337  0 t = 2
rlabel pdiffusion 427 341 428 342  0 t = 3
rlabel pdiffusion 430 341 431 342  0 t = 4
rlabel pdiffusion 426 336 432 342 0 cell no = 507
<< m1 >>
rect 427 336 428 337 
rect 430 336 431 337 
rect 427 341 428 342 
rect 430 341 431 342 
<< m2 >>
rect 427 336 428 337 
rect 430 336 431 337 
rect 427 341 428 342 
rect 430 341 431 342 
<< m2c >>
rect 427 336 428 337 
rect 430 336 431 337 
rect 427 341 428 342 
rect 430 341 431 342 
<< labels >>
rlabel pdiffusion 373 282 374 283  0 t = 1
rlabel pdiffusion 376 282 377 283  0 t = 2
rlabel pdiffusion 373 287 374 288  0 t = 3
rlabel pdiffusion 376 287 377 288  0 t = 4
rlabel pdiffusion 372 282 378 288 0 cell no = 508
<< m1 >>
rect 373 282 374 283 
rect 376 282 377 283 
rect 373 287 374 288 
rect 376 287 377 288 
<< m2 >>
rect 373 282 374 283 
rect 376 282 377 283 
rect 373 287 374 288 
rect 376 287 377 288 
<< m2c >>
rect 373 282 374 283 
rect 376 282 377 283 
rect 373 287 374 288 
rect 376 287 377 288 
<< labels >>
rlabel pdiffusion 337 444 338 445  0 t = 1
rlabel pdiffusion 340 444 341 445  0 t = 2
rlabel pdiffusion 337 449 338 450  0 t = 3
rlabel pdiffusion 340 449 341 450  0 t = 4
rlabel pdiffusion 336 444 342 450 0 cell no = 509
<< m1 >>
rect 337 444 338 445 
rect 340 444 341 445 
rect 337 449 338 450 
rect 340 449 341 450 
<< m2 >>
rect 337 444 338 445 
rect 340 444 341 445 
rect 337 449 338 450 
rect 340 449 341 450 
<< m2c >>
rect 337 444 338 445 
rect 340 444 341 445 
rect 337 449 338 450 
rect 340 449 341 450 
<< labels >>
rlabel pdiffusion 463 264 464 265  0 t = 1
rlabel pdiffusion 466 264 467 265  0 t = 2
rlabel pdiffusion 463 269 464 270  0 t = 3
rlabel pdiffusion 466 269 467 270  0 t = 4
rlabel pdiffusion 462 264 468 270 0 cell no = 510
<< m1 >>
rect 463 264 464 265 
rect 466 264 467 265 
rect 463 269 464 270 
rect 466 269 467 270 
<< m2 >>
rect 463 264 464 265 
rect 466 264 467 265 
rect 463 269 464 270 
rect 466 269 467 270 
<< m2c >>
rect 463 264 464 265 
rect 466 264 467 265 
rect 463 269 464 270 
rect 466 269 467 270 
<< labels >>
rlabel pdiffusion 265 354 266 355  0 t = 1
rlabel pdiffusion 268 354 269 355  0 t = 2
rlabel pdiffusion 265 359 266 360  0 t = 3
rlabel pdiffusion 268 359 269 360  0 t = 4
rlabel pdiffusion 264 354 270 360 0 cell no = 511
<< m1 >>
rect 265 354 266 355 
rect 268 354 269 355 
rect 265 359 266 360 
rect 268 359 269 360 
<< m2 >>
rect 265 354 266 355 
rect 268 354 269 355 
rect 265 359 266 360 
rect 268 359 269 360 
<< m2c >>
rect 265 354 266 355 
rect 268 354 269 355 
rect 265 359 266 360 
rect 268 359 269 360 
<< labels >>
rlabel pdiffusion 103 120 104 121  0 t = 1
rlabel pdiffusion 106 120 107 121  0 t = 2
rlabel pdiffusion 103 125 104 126  0 t = 3
rlabel pdiffusion 106 125 107 126  0 t = 4
rlabel pdiffusion 102 120 108 126 0 cell no = 512
<< m1 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2 >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< m2c >>
rect 103 120 104 121 
rect 106 120 107 121 
rect 103 125 104 126 
rect 106 125 107 126 
<< labels >>
rlabel pdiffusion 229 228 230 229  0 t = 1
rlabel pdiffusion 232 228 233 229  0 t = 2
rlabel pdiffusion 229 233 230 234  0 t = 3
rlabel pdiffusion 232 233 233 234  0 t = 4
rlabel pdiffusion 228 228 234 234 0 cell no = 513
<< m1 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2 >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< m2c >>
rect 229 228 230 229 
rect 232 228 233 229 
rect 229 233 230 234 
rect 232 233 233 234 
<< labels >>
rlabel pdiffusion 193 408 194 409  0 t = 1
rlabel pdiffusion 196 408 197 409  0 t = 2
rlabel pdiffusion 193 413 194 414  0 t = 3
rlabel pdiffusion 196 413 197 414  0 t = 4
rlabel pdiffusion 192 408 198 414 0 cell no = 514
<< m1 >>
rect 193 408 194 409 
rect 196 408 197 409 
rect 193 413 194 414 
rect 196 413 197 414 
<< m2 >>
rect 193 408 194 409 
rect 196 408 197 409 
rect 193 413 194 414 
rect 196 413 197 414 
<< m2c >>
rect 193 408 194 409 
rect 196 408 197 409 
rect 193 413 194 414 
rect 196 413 197 414 
<< labels >>
rlabel pdiffusion 337 372 338 373  0 t = 1
rlabel pdiffusion 340 372 341 373  0 t = 2
rlabel pdiffusion 337 377 338 378  0 t = 3
rlabel pdiffusion 340 377 341 378  0 t = 4
rlabel pdiffusion 336 372 342 378 0 cell no = 515
<< m1 >>
rect 337 372 338 373 
rect 340 372 341 373 
rect 337 377 338 378 
rect 340 377 341 378 
<< m2 >>
rect 337 372 338 373 
rect 340 372 341 373 
rect 337 377 338 378 
rect 340 377 341 378 
<< m2c >>
rect 337 372 338 373 
rect 340 372 341 373 
rect 337 377 338 378 
rect 340 377 341 378 
<< labels >>
rlabel pdiffusion 517 264 518 265  0 t = 1
rlabel pdiffusion 520 264 521 265  0 t = 2
rlabel pdiffusion 517 269 518 270  0 t = 3
rlabel pdiffusion 520 269 521 270  0 t = 4
rlabel pdiffusion 516 264 522 270 0 cell no = 516
<< m1 >>
rect 517 264 518 265 
rect 520 264 521 265 
rect 517 269 518 270 
rect 520 269 521 270 
<< m2 >>
rect 517 264 518 265 
rect 520 264 521 265 
rect 517 269 518 270 
rect 520 269 521 270 
<< m2c >>
rect 517 264 518 265 
rect 520 264 521 265 
rect 517 269 518 270 
rect 520 269 521 270 
<< labels >>
rlabel pdiffusion 463 300 464 301  0 t = 1
rlabel pdiffusion 466 300 467 301  0 t = 2
rlabel pdiffusion 463 305 464 306  0 t = 3
rlabel pdiffusion 466 305 467 306  0 t = 4
rlabel pdiffusion 462 300 468 306 0 cell no = 517
<< m1 >>
rect 463 300 464 301 
rect 466 300 467 301 
rect 463 305 464 306 
rect 466 305 467 306 
<< m2 >>
rect 463 300 464 301 
rect 466 300 467 301 
rect 463 305 464 306 
rect 466 305 467 306 
<< m2c >>
rect 463 300 464 301 
rect 466 300 467 301 
rect 463 305 464 306 
rect 466 305 467 306 
<< labels >>
rlabel pdiffusion 499 408 500 409  0 t = 1
rlabel pdiffusion 502 408 503 409  0 t = 2
rlabel pdiffusion 499 413 500 414  0 t = 3
rlabel pdiffusion 502 413 503 414  0 t = 4
rlabel pdiffusion 498 408 504 414 0 cell no = 518
<< m1 >>
rect 499 408 500 409 
rect 502 408 503 409 
rect 499 413 500 414 
rect 502 413 503 414 
<< m2 >>
rect 499 408 500 409 
rect 502 408 503 409 
rect 499 413 500 414 
rect 502 413 503 414 
<< m2c >>
rect 499 408 500 409 
rect 502 408 503 409 
rect 499 413 500 414 
rect 502 413 503 414 
<< labels >>
rlabel pdiffusion 445 318 446 319  0 t = 1
rlabel pdiffusion 448 318 449 319  0 t = 2
rlabel pdiffusion 445 323 446 324  0 t = 3
rlabel pdiffusion 448 323 449 324  0 t = 4
rlabel pdiffusion 444 318 450 324 0 cell no = 519
<< m1 >>
rect 445 318 446 319 
rect 448 318 449 319 
rect 445 323 446 324 
rect 448 323 449 324 
<< m2 >>
rect 445 318 446 319 
rect 448 318 449 319 
rect 445 323 446 324 
rect 448 323 449 324 
<< m2c >>
rect 445 318 446 319 
rect 448 318 449 319 
rect 445 323 446 324 
rect 448 323 449 324 
<< labels >>
rlabel pdiffusion 445 264 446 265  0 t = 1
rlabel pdiffusion 448 264 449 265  0 t = 2
rlabel pdiffusion 445 269 446 270  0 t = 3
rlabel pdiffusion 448 269 449 270  0 t = 4
rlabel pdiffusion 444 264 450 270 0 cell no = 520
<< m1 >>
rect 445 264 446 265 
rect 448 264 449 265 
rect 445 269 446 270 
rect 448 269 449 270 
<< m2 >>
rect 445 264 446 265 
rect 448 264 449 265 
rect 445 269 446 270 
rect 448 269 449 270 
<< m2c >>
rect 445 264 446 265 
rect 448 264 449 265 
rect 445 269 446 270 
rect 448 269 449 270 
<< labels >>
rlabel pdiffusion 409 138 410 139  0 t = 1
rlabel pdiffusion 412 138 413 139  0 t = 2
rlabel pdiffusion 409 143 410 144  0 t = 3
rlabel pdiffusion 412 143 413 144  0 t = 4
rlabel pdiffusion 408 138 414 144 0 cell no = 521
<< m1 >>
rect 409 138 410 139 
rect 412 138 413 139 
rect 409 143 410 144 
rect 412 143 413 144 
<< m2 >>
rect 409 138 410 139 
rect 412 138 413 139 
rect 409 143 410 144 
rect 412 143 413 144 
<< m2c >>
rect 409 138 410 139 
rect 412 138 413 139 
rect 409 143 410 144 
rect 412 143 413 144 
<< labels >>
rlabel pdiffusion 463 282 464 283  0 t = 1
rlabel pdiffusion 466 282 467 283  0 t = 2
rlabel pdiffusion 463 287 464 288  0 t = 3
rlabel pdiffusion 466 287 467 288  0 t = 4
rlabel pdiffusion 462 282 468 288 0 cell no = 522
<< m1 >>
rect 463 282 464 283 
rect 466 282 467 283 
rect 463 287 464 288 
rect 466 287 467 288 
<< m2 >>
rect 463 282 464 283 
rect 466 282 467 283 
rect 463 287 464 288 
rect 466 287 467 288 
<< m2c >>
rect 463 282 464 283 
rect 466 282 467 283 
rect 463 287 464 288 
rect 466 287 467 288 
<< labels >>
rlabel pdiffusion 103 318 104 319  0 t = 1
rlabel pdiffusion 106 318 107 319  0 t = 2
rlabel pdiffusion 103 323 104 324  0 t = 3
rlabel pdiffusion 106 323 107 324  0 t = 4
rlabel pdiffusion 102 318 108 324 0 cell no = 523
<< m1 >>
rect 103 318 104 319 
rect 106 318 107 319 
rect 103 323 104 324 
rect 106 323 107 324 
<< m2 >>
rect 103 318 104 319 
rect 106 318 107 319 
rect 103 323 104 324 
rect 106 323 107 324 
<< m2c >>
rect 103 318 104 319 
rect 106 318 107 319 
rect 103 323 104 324 
rect 106 323 107 324 
<< labels >>
rlabel pdiffusion 85 444 86 445  0 t = 1
rlabel pdiffusion 88 444 89 445  0 t = 2
rlabel pdiffusion 85 449 86 450  0 t = 3
rlabel pdiffusion 88 449 89 450  0 t = 4
rlabel pdiffusion 84 444 90 450 0 cell no = 524
<< m1 >>
rect 85 444 86 445 
rect 88 444 89 445 
rect 85 449 86 450 
rect 88 449 89 450 
<< m2 >>
rect 85 444 86 445 
rect 88 444 89 445 
rect 85 449 86 450 
rect 88 449 89 450 
<< m2c >>
rect 85 444 86 445 
rect 88 444 89 445 
rect 85 449 86 450 
rect 88 449 89 450 
<< labels >>
rlabel pdiffusion 445 426 446 427  0 t = 1
rlabel pdiffusion 448 426 449 427  0 t = 2
rlabel pdiffusion 445 431 446 432  0 t = 3
rlabel pdiffusion 448 431 449 432  0 t = 4
rlabel pdiffusion 444 426 450 432 0 cell no = 525
<< m1 >>
rect 445 426 446 427 
rect 448 426 449 427 
rect 445 431 446 432 
rect 448 431 449 432 
<< m2 >>
rect 445 426 446 427 
rect 448 426 449 427 
rect 445 431 446 432 
rect 448 431 449 432 
<< m2c >>
rect 445 426 446 427 
rect 448 426 449 427 
rect 445 431 446 432 
rect 448 431 449 432 
<< labels >>
rlabel pdiffusion 229 174 230 175  0 t = 1
rlabel pdiffusion 232 174 233 175  0 t = 2
rlabel pdiffusion 229 179 230 180  0 t = 3
rlabel pdiffusion 232 179 233 180  0 t = 4
rlabel pdiffusion 228 174 234 180 0 cell no = 526
<< m1 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2 >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< m2c >>
rect 229 174 230 175 
rect 232 174 233 175 
rect 229 179 230 180 
rect 232 179 233 180 
<< labels >>
rlabel pdiffusion 319 516 320 517  0 t = 1
rlabel pdiffusion 322 516 323 517  0 t = 2
rlabel pdiffusion 319 521 320 522  0 t = 3
rlabel pdiffusion 322 521 323 522  0 t = 4
rlabel pdiffusion 318 516 324 522 0 cell no = 527
<< m1 >>
rect 319 516 320 517 
rect 322 516 323 517 
rect 319 521 320 522 
rect 322 521 323 522 
<< m2 >>
rect 319 516 320 517 
rect 322 516 323 517 
rect 319 521 320 522 
rect 322 521 323 522 
<< m2c >>
rect 319 516 320 517 
rect 322 516 323 517 
rect 319 521 320 522 
rect 322 521 323 522 
<< labels >>
rlabel pdiffusion 103 228 104 229  0 t = 1
rlabel pdiffusion 106 228 107 229  0 t = 2
rlabel pdiffusion 103 233 104 234  0 t = 3
rlabel pdiffusion 106 233 107 234  0 t = 4
rlabel pdiffusion 102 228 108 234 0 cell no = 528
<< m1 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2 >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< m2c >>
rect 103 228 104 229 
rect 106 228 107 229 
rect 103 233 104 234 
rect 106 233 107 234 
<< labels >>
rlabel pdiffusion 283 444 284 445  0 t = 1
rlabel pdiffusion 286 444 287 445  0 t = 2
rlabel pdiffusion 283 449 284 450  0 t = 3
rlabel pdiffusion 286 449 287 450  0 t = 4
rlabel pdiffusion 282 444 288 450 0 cell no = 529
<< m1 >>
rect 283 444 284 445 
rect 286 444 287 445 
rect 283 449 284 450 
rect 286 449 287 450 
<< m2 >>
rect 283 444 284 445 
rect 286 444 287 445 
rect 283 449 284 450 
rect 286 449 287 450 
<< m2c >>
rect 283 444 284 445 
rect 286 444 287 445 
rect 283 449 284 450 
rect 286 449 287 450 
<< labels >>
rlabel pdiffusion 103 480 104 481  0 t = 1
rlabel pdiffusion 106 480 107 481  0 t = 2
rlabel pdiffusion 103 485 104 486  0 t = 3
rlabel pdiffusion 106 485 107 486  0 t = 4
rlabel pdiffusion 102 480 108 486 0 cell no = 530
<< m1 >>
rect 103 480 104 481 
rect 106 480 107 481 
rect 103 485 104 486 
rect 106 485 107 486 
<< m2 >>
rect 103 480 104 481 
rect 106 480 107 481 
rect 103 485 104 486 
rect 106 485 107 486 
<< m2c >>
rect 103 480 104 481 
rect 106 480 107 481 
rect 103 485 104 486 
rect 106 485 107 486 
<< labels >>
rlabel pdiffusion 193 192 194 193  0 t = 1
rlabel pdiffusion 196 192 197 193  0 t = 2
rlabel pdiffusion 193 197 194 198  0 t = 3
rlabel pdiffusion 196 197 197 198  0 t = 4
rlabel pdiffusion 192 192 198 198 0 cell no = 531
<< m1 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2 >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< m2c >>
rect 193 192 194 193 
rect 196 192 197 193 
rect 193 197 194 198 
rect 196 197 197 198 
<< labels >>
rlabel pdiffusion 157 228 158 229  0 t = 1
rlabel pdiffusion 160 228 161 229  0 t = 2
rlabel pdiffusion 157 233 158 234  0 t = 3
rlabel pdiffusion 160 233 161 234  0 t = 4
rlabel pdiffusion 156 228 162 234 0 cell no = 532
<< m1 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2 >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< m2c >>
rect 157 228 158 229 
rect 160 228 161 229 
rect 157 233 158 234 
rect 160 233 161 234 
<< labels >>
rlabel pdiffusion 355 372 356 373  0 t = 1
rlabel pdiffusion 358 372 359 373  0 t = 2
rlabel pdiffusion 355 377 356 378  0 t = 3
rlabel pdiffusion 358 377 359 378  0 t = 4
rlabel pdiffusion 354 372 360 378 0 cell no = 533
<< m1 >>
rect 355 372 356 373 
rect 358 372 359 373 
rect 355 377 356 378 
rect 358 377 359 378 
<< m2 >>
rect 355 372 356 373 
rect 358 372 359 373 
rect 355 377 356 378 
rect 358 377 359 378 
<< m2c >>
rect 355 372 356 373 
rect 358 372 359 373 
rect 355 377 356 378 
rect 358 377 359 378 
<< labels >>
rlabel pdiffusion 121 426 122 427  0 t = 1
rlabel pdiffusion 124 426 125 427  0 t = 2
rlabel pdiffusion 121 431 122 432  0 t = 3
rlabel pdiffusion 124 431 125 432  0 t = 4
rlabel pdiffusion 120 426 126 432 0 cell no = 534
<< m1 >>
rect 121 426 122 427 
rect 124 426 125 427 
rect 121 431 122 432 
rect 124 431 125 432 
<< m2 >>
rect 121 426 122 427 
rect 124 426 125 427 
rect 121 431 122 432 
rect 124 431 125 432 
<< m2c >>
rect 121 426 122 427 
rect 124 426 125 427 
rect 121 431 122 432 
rect 124 431 125 432 
<< labels >>
rlabel pdiffusion 211 336 212 337  0 t = 1
rlabel pdiffusion 214 336 215 337  0 t = 2
rlabel pdiffusion 211 341 212 342  0 t = 3
rlabel pdiffusion 214 341 215 342  0 t = 4
rlabel pdiffusion 210 336 216 342 0 cell no = 535
<< m1 >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< m2 >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< m2c >>
rect 211 336 212 337 
rect 214 336 215 337 
rect 211 341 212 342 
rect 214 341 215 342 
<< labels >>
rlabel pdiffusion 337 354 338 355  0 t = 1
rlabel pdiffusion 340 354 341 355  0 t = 2
rlabel pdiffusion 337 359 338 360  0 t = 3
rlabel pdiffusion 340 359 341 360  0 t = 4
rlabel pdiffusion 336 354 342 360 0 cell no = 536
<< m1 >>
rect 337 354 338 355 
rect 340 354 341 355 
rect 337 359 338 360 
rect 340 359 341 360 
<< m2 >>
rect 337 354 338 355 
rect 340 354 341 355 
rect 337 359 338 360 
rect 340 359 341 360 
<< m2c >>
rect 337 354 338 355 
rect 340 354 341 355 
rect 337 359 338 360 
rect 340 359 341 360 
<< labels >>
rlabel pdiffusion 301 228 302 229  0 t = 1
rlabel pdiffusion 304 228 305 229  0 t = 2
rlabel pdiffusion 301 233 302 234  0 t = 3
rlabel pdiffusion 304 233 305 234  0 t = 4
rlabel pdiffusion 300 228 306 234 0 cell no = 537
<< m1 >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< m2 >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< m2c >>
rect 301 228 302 229 
rect 304 228 305 229 
rect 301 233 302 234 
rect 304 233 305 234 
<< labels >>
rlabel pdiffusion 427 444 428 445  0 t = 1
rlabel pdiffusion 430 444 431 445  0 t = 2
rlabel pdiffusion 427 449 428 450  0 t = 3
rlabel pdiffusion 430 449 431 450  0 t = 4
rlabel pdiffusion 426 444 432 450 0 cell no = 538
<< m1 >>
rect 427 444 428 445 
rect 430 444 431 445 
rect 427 449 428 450 
rect 430 449 431 450 
<< m2 >>
rect 427 444 428 445 
rect 430 444 431 445 
rect 427 449 428 450 
rect 430 449 431 450 
<< m2c >>
rect 427 444 428 445 
rect 430 444 431 445 
rect 427 449 428 450 
rect 430 449 431 450 
<< labels >>
rlabel pdiffusion 265 390 266 391  0 t = 1
rlabel pdiffusion 268 390 269 391  0 t = 2
rlabel pdiffusion 265 395 266 396  0 t = 3
rlabel pdiffusion 268 395 269 396  0 t = 4
rlabel pdiffusion 264 390 270 396 0 cell no = 539
<< m1 >>
rect 265 390 266 391 
rect 268 390 269 391 
rect 265 395 266 396 
rect 268 395 269 396 
<< m2 >>
rect 265 390 266 391 
rect 268 390 269 391 
rect 265 395 266 396 
rect 268 395 269 396 
<< m2c >>
rect 265 390 266 391 
rect 268 390 269 391 
rect 265 395 266 396 
rect 268 395 269 396 
<< labels >>
rlabel pdiffusion 373 480 374 481  0 t = 1
rlabel pdiffusion 376 480 377 481  0 t = 2
rlabel pdiffusion 373 485 374 486  0 t = 3
rlabel pdiffusion 376 485 377 486  0 t = 4
rlabel pdiffusion 372 480 378 486 0 cell no = 540
<< m1 >>
rect 373 480 374 481 
rect 376 480 377 481 
rect 373 485 374 486 
rect 376 485 377 486 
<< m2 >>
rect 373 480 374 481 
rect 376 480 377 481 
rect 373 485 374 486 
rect 376 485 377 486 
<< m2c >>
rect 373 480 374 481 
rect 376 480 377 481 
rect 373 485 374 486 
rect 376 485 377 486 
<< labels >>
rlabel pdiffusion 355 264 356 265  0 t = 1
rlabel pdiffusion 358 264 359 265  0 t = 2
rlabel pdiffusion 355 269 356 270  0 t = 3
rlabel pdiffusion 358 269 359 270  0 t = 4
rlabel pdiffusion 354 264 360 270 0 cell no = 541
<< m1 >>
rect 355 264 356 265 
rect 358 264 359 265 
rect 355 269 356 270 
rect 358 269 359 270 
<< m2 >>
rect 355 264 356 265 
rect 358 264 359 265 
rect 355 269 356 270 
rect 358 269 359 270 
<< m2c >>
rect 355 264 356 265 
rect 358 264 359 265 
rect 355 269 356 270 
rect 358 269 359 270 
<< labels >>
rlabel pdiffusion 283 354 284 355  0 t = 1
rlabel pdiffusion 286 354 287 355  0 t = 2
rlabel pdiffusion 283 359 284 360  0 t = 3
rlabel pdiffusion 286 359 287 360  0 t = 4
rlabel pdiffusion 282 354 288 360 0 cell no = 542
<< m1 >>
rect 283 354 284 355 
rect 286 354 287 355 
rect 283 359 284 360 
rect 286 359 287 360 
<< m2 >>
rect 283 354 284 355 
rect 286 354 287 355 
rect 283 359 284 360 
rect 286 359 287 360 
<< m2c >>
rect 283 354 284 355 
rect 286 354 287 355 
rect 283 359 284 360 
rect 286 359 287 360 
<< labels >>
rlabel pdiffusion 409 336 410 337  0 t = 1
rlabel pdiffusion 412 336 413 337  0 t = 2
rlabel pdiffusion 409 341 410 342  0 t = 3
rlabel pdiffusion 412 341 413 342  0 t = 4
rlabel pdiffusion 408 336 414 342 0 cell no = 543
<< m1 >>
rect 409 336 410 337 
rect 412 336 413 337 
rect 409 341 410 342 
rect 412 341 413 342 
<< m2 >>
rect 409 336 410 337 
rect 412 336 413 337 
rect 409 341 410 342 
rect 412 341 413 342 
<< m2c >>
rect 409 336 410 337 
rect 412 336 413 337 
rect 409 341 410 342 
rect 412 341 413 342 
<< labels >>
rlabel pdiffusion 445 282 446 283  0 t = 1
rlabel pdiffusion 448 282 449 283  0 t = 2
rlabel pdiffusion 445 287 446 288  0 t = 3
rlabel pdiffusion 448 287 449 288  0 t = 4
rlabel pdiffusion 444 282 450 288 0 cell no = 544
<< m1 >>
rect 445 282 446 283 
rect 448 282 449 283 
rect 445 287 446 288 
rect 448 287 449 288 
<< m2 >>
rect 445 282 446 283 
rect 448 282 449 283 
rect 445 287 446 288 
rect 448 287 449 288 
<< m2c >>
rect 445 282 446 283 
rect 448 282 449 283 
rect 445 287 446 288 
rect 448 287 449 288 
<< labels >>
rlabel pdiffusion 517 390 518 391  0 t = 1
rlabel pdiffusion 520 390 521 391  0 t = 2
rlabel pdiffusion 517 395 518 396  0 t = 3
rlabel pdiffusion 520 395 521 396  0 t = 4
rlabel pdiffusion 516 390 522 396 0 cell no = 545
<< m1 >>
rect 517 390 518 391 
rect 520 390 521 391 
rect 517 395 518 396 
rect 520 395 521 396 
<< m2 >>
rect 517 390 518 391 
rect 520 390 521 391 
rect 517 395 518 396 
rect 520 395 521 396 
<< m2c >>
rect 517 390 518 391 
rect 520 390 521 391 
rect 517 395 518 396 
rect 520 395 521 396 
<< labels >>
rlabel pdiffusion 373 354 374 355  0 t = 1
rlabel pdiffusion 376 354 377 355  0 t = 2
rlabel pdiffusion 373 359 374 360  0 t = 3
rlabel pdiffusion 376 359 377 360  0 t = 4
rlabel pdiffusion 372 354 378 360 0 cell no = 546
<< m1 >>
rect 373 354 374 355 
rect 376 354 377 355 
rect 373 359 374 360 
rect 376 359 377 360 
<< m2 >>
rect 373 354 374 355 
rect 376 354 377 355 
rect 373 359 374 360 
rect 376 359 377 360 
<< m2c >>
rect 373 354 374 355 
rect 376 354 377 355 
rect 373 359 374 360 
rect 376 359 377 360 
<< labels >>
rlabel pdiffusion 481 408 482 409  0 t = 1
rlabel pdiffusion 484 408 485 409  0 t = 2
rlabel pdiffusion 481 413 482 414  0 t = 3
rlabel pdiffusion 484 413 485 414  0 t = 4
rlabel pdiffusion 480 408 486 414 0 cell no = 547
<< m1 >>
rect 481 408 482 409 
rect 484 408 485 409 
rect 481 413 482 414 
rect 484 413 485 414 
<< m2 >>
rect 481 408 482 409 
rect 484 408 485 409 
rect 481 413 482 414 
rect 484 413 485 414 
<< m2c >>
rect 481 408 482 409 
rect 484 408 485 409 
rect 481 413 482 414 
rect 484 413 485 414 
<< labels >>
rlabel pdiffusion 229 498 230 499  0 t = 1
rlabel pdiffusion 232 498 233 499  0 t = 2
rlabel pdiffusion 229 503 230 504  0 t = 3
rlabel pdiffusion 232 503 233 504  0 t = 4
rlabel pdiffusion 228 498 234 504 0 cell no = 548
<< m1 >>
rect 229 498 230 499 
rect 232 498 233 499 
rect 229 503 230 504 
rect 232 503 233 504 
<< m2 >>
rect 229 498 230 499 
rect 232 498 233 499 
rect 229 503 230 504 
rect 232 503 233 504 
<< m2c >>
rect 229 498 230 499 
rect 232 498 233 499 
rect 229 503 230 504 
rect 232 503 233 504 
<< labels >>
rlabel pdiffusion 319 282 320 283  0 t = 1
rlabel pdiffusion 322 282 323 283  0 t = 2
rlabel pdiffusion 319 287 320 288  0 t = 3
rlabel pdiffusion 322 287 323 288  0 t = 4
rlabel pdiffusion 318 282 324 288 0 cell no = 549
<< m1 >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< m2 >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< m2c >>
rect 319 282 320 283 
rect 322 282 323 283 
rect 319 287 320 288 
rect 322 287 323 288 
<< labels >>
rlabel pdiffusion 355 282 356 283  0 t = 1
rlabel pdiffusion 358 282 359 283  0 t = 2
rlabel pdiffusion 355 287 356 288  0 t = 3
rlabel pdiffusion 358 287 359 288  0 t = 4
rlabel pdiffusion 354 282 360 288 0 cell no = 550
<< m1 >>
rect 355 282 356 283 
rect 358 282 359 283 
rect 355 287 356 288 
rect 358 287 359 288 
<< m2 >>
rect 355 282 356 283 
rect 358 282 359 283 
rect 355 287 356 288 
rect 358 287 359 288 
<< m2c >>
rect 355 282 356 283 
rect 358 282 359 283 
rect 355 287 356 288 
rect 358 287 359 288 
<< labels >>
rlabel pdiffusion 49 390 50 391  0 t = 1
rlabel pdiffusion 52 390 53 391  0 t = 2
rlabel pdiffusion 49 395 50 396  0 t = 3
rlabel pdiffusion 52 395 53 396  0 t = 4
rlabel pdiffusion 48 390 54 396 0 cell no = 551
<< m1 >>
rect 49 390 50 391 
rect 52 390 53 391 
rect 49 395 50 396 
rect 52 395 53 396 
<< m2 >>
rect 49 390 50 391 
rect 52 390 53 391 
rect 49 395 50 396 
rect 52 395 53 396 
<< m2c >>
rect 49 390 50 391 
rect 52 390 53 391 
rect 49 395 50 396 
rect 52 395 53 396 
<< labels >>
rlabel pdiffusion 175 354 176 355  0 t = 1
rlabel pdiffusion 178 354 179 355  0 t = 2
rlabel pdiffusion 175 359 176 360  0 t = 3
rlabel pdiffusion 178 359 179 360  0 t = 4
rlabel pdiffusion 174 354 180 360 0 cell no = 552
<< m1 >>
rect 175 354 176 355 
rect 178 354 179 355 
rect 175 359 176 360 
rect 178 359 179 360 
<< m2 >>
rect 175 354 176 355 
rect 178 354 179 355 
rect 175 359 176 360 
rect 178 359 179 360 
<< m2c >>
rect 175 354 176 355 
rect 178 354 179 355 
rect 175 359 176 360 
rect 178 359 179 360 
<< labels >>
rlabel pdiffusion 211 354 212 355  0 t = 1
rlabel pdiffusion 214 354 215 355  0 t = 2
rlabel pdiffusion 211 359 212 360  0 t = 3
rlabel pdiffusion 214 359 215 360  0 t = 4
rlabel pdiffusion 210 354 216 360 0 cell no = 553
<< m1 >>
rect 211 354 212 355 
rect 214 354 215 355 
rect 211 359 212 360 
rect 214 359 215 360 
<< m2 >>
rect 211 354 212 355 
rect 214 354 215 355 
rect 211 359 212 360 
rect 214 359 215 360 
<< m2c >>
rect 211 354 212 355 
rect 214 354 215 355 
rect 211 359 212 360 
rect 214 359 215 360 
<< labels >>
rlabel pdiffusion 85 264 86 265  0 t = 1
rlabel pdiffusion 88 264 89 265  0 t = 2
rlabel pdiffusion 85 269 86 270  0 t = 3
rlabel pdiffusion 88 269 89 270  0 t = 4
rlabel pdiffusion 84 264 90 270 0 cell no = 554
<< m1 >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< m2 >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< m2c >>
rect 85 264 86 265 
rect 88 264 89 265 
rect 85 269 86 270 
rect 88 269 89 270 
<< labels >>
rlabel pdiffusion 193 210 194 211  0 t = 1
rlabel pdiffusion 196 210 197 211  0 t = 2
rlabel pdiffusion 193 215 194 216  0 t = 3
rlabel pdiffusion 196 215 197 216  0 t = 4
rlabel pdiffusion 192 210 198 216 0 cell no = 555
<< m1 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2 >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< m2c >>
rect 193 210 194 211 
rect 196 210 197 211 
rect 193 215 194 216 
rect 196 215 197 216 
<< labels >>
rlabel pdiffusion 49 264 50 265  0 t = 1
rlabel pdiffusion 52 264 53 265  0 t = 2
rlabel pdiffusion 49 269 50 270  0 t = 3
rlabel pdiffusion 52 269 53 270  0 t = 4
rlabel pdiffusion 48 264 54 270 0 cell no = 556
<< m1 >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< m2 >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< m2c >>
rect 49 264 50 265 
rect 52 264 53 265 
rect 49 269 50 270 
rect 52 269 53 270 
<< labels >>
rlabel pdiffusion 265 246 266 247  0 t = 1
rlabel pdiffusion 268 246 269 247  0 t = 2
rlabel pdiffusion 265 251 266 252  0 t = 3
rlabel pdiffusion 268 251 269 252  0 t = 4
rlabel pdiffusion 264 246 270 252 0 cell no = 557
<< m1 >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< m2 >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< m2c >>
rect 265 246 266 247 
rect 268 246 269 247 
rect 265 251 266 252 
rect 268 251 269 252 
<< labels >>
rlabel pdiffusion 103 264 104 265  0 t = 1
rlabel pdiffusion 106 264 107 265  0 t = 2
rlabel pdiffusion 103 269 104 270  0 t = 3
rlabel pdiffusion 106 269 107 270  0 t = 4
rlabel pdiffusion 102 264 108 270 0 cell no = 558
<< m1 >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< m2 >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< m2c >>
rect 103 264 104 265 
rect 106 264 107 265 
rect 103 269 104 270 
rect 106 269 107 270 
<< labels >>
rlabel pdiffusion 121 192 122 193  0 t = 1
rlabel pdiffusion 124 192 125 193  0 t = 2
rlabel pdiffusion 121 197 122 198  0 t = 3
rlabel pdiffusion 124 197 125 198  0 t = 4
rlabel pdiffusion 120 192 126 198 0 cell no = 559
<< m1 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2 >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< m2c >>
rect 121 192 122 193 
rect 124 192 125 193 
rect 121 197 122 198 
rect 124 197 125 198 
<< labels >>
rlabel pdiffusion 427 354 428 355  0 t = 1
rlabel pdiffusion 430 354 431 355  0 t = 2
rlabel pdiffusion 427 359 428 360  0 t = 3
rlabel pdiffusion 430 359 431 360  0 t = 4
rlabel pdiffusion 426 354 432 360 0 cell no = 560
<< m1 >>
rect 427 354 428 355 
rect 430 354 431 355 
rect 427 359 428 360 
rect 430 359 431 360 
<< m2 >>
rect 427 354 428 355 
rect 430 354 431 355 
rect 427 359 428 360 
rect 430 359 431 360 
<< m2c >>
rect 427 354 428 355 
rect 430 354 431 355 
rect 427 359 428 360 
rect 430 359 431 360 
<< labels >>
rlabel pdiffusion 121 120 122 121  0 t = 1
rlabel pdiffusion 124 120 125 121  0 t = 2
rlabel pdiffusion 121 125 122 126  0 t = 3
rlabel pdiffusion 124 125 125 126  0 t = 4
rlabel pdiffusion 120 120 126 126 0 cell no = 561
<< m1 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2 >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< m2c >>
rect 121 120 122 121 
rect 124 120 125 121 
rect 121 125 122 126 
rect 124 125 125 126 
<< labels >>
rlabel pdiffusion 337 264 338 265  0 t = 1
rlabel pdiffusion 340 264 341 265  0 t = 2
rlabel pdiffusion 337 269 338 270  0 t = 3
rlabel pdiffusion 340 269 341 270  0 t = 4
rlabel pdiffusion 336 264 342 270 0 cell no = 562
<< m1 >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< m2 >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< m2c >>
rect 337 264 338 265 
rect 340 264 341 265 
rect 337 269 338 270 
rect 340 269 341 270 
<< labels >>
rlabel pdiffusion 139 390 140 391  0 t = 1
rlabel pdiffusion 142 390 143 391  0 t = 2
rlabel pdiffusion 139 395 140 396  0 t = 3
rlabel pdiffusion 142 395 143 396  0 t = 4
rlabel pdiffusion 138 390 144 396 0 cell no = 563
<< m1 >>
rect 139 390 140 391 
rect 142 390 143 391 
rect 139 395 140 396 
rect 142 395 143 396 
<< m2 >>
rect 139 390 140 391 
rect 142 390 143 391 
rect 139 395 140 396 
rect 142 395 143 396 
<< m2c >>
rect 139 390 140 391 
rect 142 390 143 391 
rect 139 395 140 396 
rect 142 395 143 396 
<< labels >>
rlabel pdiffusion 481 390 482 391  0 t = 1
rlabel pdiffusion 484 390 485 391  0 t = 2
rlabel pdiffusion 481 395 482 396  0 t = 3
rlabel pdiffusion 484 395 485 396  0 t = 4
rlabel pdiffusion 480 390 486 396 0 cell no = 564
<< m1 >>
rect 481 390 482 391 
rect 484 390 485 391 
rect 481 395 482 396 
rect 484 395 485 396 
<< m2 >>
rect 481 390 482 391 
rect 484 390 485 391 
rect 481 395 482 396 
rect 484 395 485 396 
<< m2c >>
rect 481 390 482 391 
rect 484 390 485 391 
rect 481 395 482 396 
rect 484 395 485 396 
<< labels >>
rlabel pdiffusion 247 408 248 409  0 t = 1
rlabel pdiffusion 250 408 251 409  0 t = 2
rlabel pdiffusion 247 413 248 414  0 t = 3
rlabel pdiffusion 250 413 251 414  0 t = 4
rlabel pdiffusion 246 408 252 414 0 cell no = 565
<< m1 >>
rect 247 408 248 409 
rect 250 408 251 409 
rect 247 413 248 414 
rect 250 413 251 414 
<< m2 >>
rect 247 408 248 409 
rect 250 408 251 409 
rect 247 413 248 414 
rect 250 413 251 414 
<< m2c >>
rect 247 408 248 409 
rect 250 408 251 409 
rect 247 413 248 414 
rect 250 413 251 414 
<< labels >>
rlabel pdiffusion 337 408 338 409  0 t = 1
rlabel pdiffusion 340 408 341 409  0 t = 2
rlabel pdiffusion 337 413 338 414  0 t = 3
rlabel pdiffusion 340 413 341 414  0 t = 4
rlabel pdiffusion 336 408 342 414 0 cell no = 566
<< m1 >>
rect 337 408 338 409 
rect 340 408 341 409 
rect 337 413 338 414 
rect 340 413 341 414 
<< m2 >>
rect 337 408 338 409 
rect 340 408 341 409 
rect 337 413 338 414 
rect 340 413 341 414 
<< m2c >>
rect 337 408 338 409 
rect 340 408 341 409 
rect 337 413 338 414 
rect 340 413 341 414 
<< labels >>
rlabel pdiffusion 301 300 302 301  0 t = 1
rlabel pdiffusion 304 300 305 301  0 t = 2
rlabel pdiffusion 301 305 302 306  0 t = 3
rlabel pdiffusion 304 305 305 306  0 t = 4
rlabel pdiffusion 300 300 306 306 0 cell no = 567
<< m1 >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< m2 >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< m2c >>
rect 301 300 302 301 
rect 304 300 305 301 
rect 301 305 302 306 
rect 304 305 305 306 
<< labels >>
rlabel pdiffusion 265 138 266 139  0 t = 1
rlabel pdiffusion 268 138 269 139  0 t = 2
rlabel pdiffusion 265 143 266 144  0 t = 3
rlabel pdiffusion 268 143 269 144  0 t = 4
rlabel pdiffusion 264 138 270 144 0 cell no = 568
<< m1 >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< m2 >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< m2c >>
rect 265 138 266 139 
rect 268 138 269 139 
rect 265 143 266 144 
rect 268 143 269 144 
<< labels >>
rlabel pdiffusion 229 390 230 391  0 t = 1
rlabel pdiffusion 232 390 233 391  0 t = 2
rlabel pdiffusion 229 395 230 396  0 t = 3
rlabel pdiffusion 232 395 233 396  0 t = 4
rlabel pdiffusion 228 390 234 396 0 cell no = 569
<< m1 >>
rect 229 390 230 391 
rect 232 390 233 391 
rect 229 395 230 396 
rect 232 395 233 396 
<< m2 >>
rect 229 390 230 391 
rect 232 390 233 391 
rect 229 395 230 396 
rect 232 395 233 396 
<< m2c >>
rect 229 390 230 391 
rect 232 390 233 391 
rect 229 395 230 396 
rect 232 395 233 396 
<< labels >>
rlabel pdiffusion 355 336 356 337  0 t = 1
rlabel pdiffusion 358 336 359 337  0 t = 2
rlabel pdiffusion 355 341 356 342  0 t = 3
rlabel pdiffusion 358 341 359 342  0 t = 4
rlabel pdiffusion 354 336 360 342 0 cell no = 570
<< m1 >>
rect 355 336 356 337 
rect 358 336 359 337 
rect 355 341 356 342 
rect 358 341 359 342 
<< m2 >>
rect 355 336 356 337 
rect 358 336 359 337 
rect 355 341 356 342 
rect 358 341 359 342 
<< m2c >>
rect 355 336 356 337 
rect 358 336 359 337 
rect 355 341 356 342 
rect 358 341 359 342 
<< labels >>
rlabel pdiffusion 301 408 302 409  0 t = 1
rlabel pdiffusion 304 408 305 409  0 t = 2
rlabel pdiffusion 301 413 302 414  0 t = 3
rlabel pdiffusion 304 413 305 414  0 t = 4
rlabel pdiffusion 300 408 306 414 0 cell no = 571
<< m1 >>
rect 301 408 302 409 
rect 304 408 305 409 
rect 301 413 302 414 
rect 304 413 305 414 
<< m2 >>
rect 301 408 302 409 
rect 304 408 305 409 
rect 301 413 302 414 
rect 304 413 305 414 
<< m2c >>
rect 301 408 302 409 
rect 304 408 305 409 
rect 301 413 302 414 
rect 304 413 305 414 
<< labels >>
rlabel pdiffusion 85 372 86 373  0 t = 1
rlabel pdiffusion 88 372 89 373  0 t = 2
rlabel pdiffusion 85 377 86 378  0 t = 3
rlabel pdiffusion 88 377 89 378  0 t = 4
rlabel pdiffusion 84 372 90 378 0 cell no = 572
<< m1 >>
rect 85 372 86 373 
rect 88 372 89 373 
rect 85 377 86 378 
rect 88 377 89 378 
<< m2 >>
rect 85 372 86 373 
rect 88 372 89 373 
rect 85 377 86 378 
rect 88 377 89 378 
<< m2c >>
rect 85 372 86 373 
rect 88 372 89 373 
rect 85 377 86 378 
rect 88 377 89 378 
<< labels >>
rlabel pdiffusion 427 192 428 193  0 t = 1
rlabel pdiffusion 430 192 431 193  0 t = 2
rlabel pdiffusion 427 197 428 198  0 t = 3
rlabel pdiffusion 430 197 431 198  0 t = 4
rlabel pdiffusion 426 192 432 198 0 cell no = 573
<< m1 >>
rect 427 192 428 193 
rect 430 192 431 193 
rect 427 197 428 198 
rect 430 197 431 198 
<< m2 >>
rect 427 192 428 193 
rect 430 192 431 193 
rect 427 197 428 198 
rect 430 197 431 198 
<< m2c >>
rect 427 192 428 193 
rect 430 192 431 193 
rect 427 197 428 198 
rect 430 197 431 198 
<< labels >>
rlabel pdiffusion 391 498 392 499  0 t = 1
rlabel pdiffusion 394 498 395 499  0 t = 2
rlabel pdiffusion 391 503 392 504  0 t = 3
rlabel pdiffusion 394 503 395 504  0 t = 4
rlabel pdiffusion 390 498 396 504 0 cell no = 574
<< m1 >>
rect 391 498 392 499 
rect 394 498 395 499 
rect 391 503 392 504 
rect 394 503 395 504 
<< m2 >>
rect 391 498 392 499 
rect 394 498 395 499 
rect 391 503 392 504 
rect 394 503 395 504 
<< m2c >>
rect 391 498 392 499 
rect 394 498 395 499 
rect 391 503 392 504 
rect 394 503 395 504 
<< labels >>
rlabel pdiffusion 517 462 518 463  0 t = 1
rlabel pdiffusion 520 462 521 463  0 t = 2
rlabel pdiffusion 517 467 518 468  0 t = 3
rlabel pdiffusion 520 467 521 468  0 t = 4
rlabel pdiffusion 516 462 522 468 0 cell no = 575
<< m1 >>
rect 517 462 518 463 
rect 520 462 521 463 
rect 517 467 518 468 
rect 520 467 521 468 
<< m2 >>
rect 517 462 518 463 
rect 520 462 521 463 
rect 517 467 518 468 
rect 520 467 521 468 
<< m2c >>
rect 517 462 518 463 
rect 520 462 521 463 
rect 517 467 518 468 
rect 520 467 521 468 
<< labels >>
rlabel pdiffusion 481 444 482 445  0 t = 1
rlabel pdiffusion 484 444 485 445  0 t = 2
rlabel pdiffusion 481 449 482 450  0 t = 3
rlabel pdiffusion 484 449 485 450  0 t = 4
rlabel pdiffusion 480 444 486 450 0 cell no = 576
<< m1 >>
rect 481 444 482 445 
rect 484 444 485 445 
rect 481 449 482 450 
rect 484 449 485 450 
<< m2 >>
rect 481 444 482 445 
rect 484 444 485 445 
rect 481 449 482 450 
rect 484 449 485 450 
<< m2c >>
rect 481 444 482 445 
rect 484 444 485 445 
rect 481 449 482 450 
rect 484 449 485 450 
<< labels >>
rlabel pdiffusion 445 390 446 391  0 t = 1
rlabel pdiffusion 448 390 449 391  0 t = 2
rlabel pdiffusion 445 395 446 396  0 t = 3
rlabel pdiffusion 448 395 449 396  0 t = 4
rlabel pdiffusion 444 390 450 396 0 cell no = 577
<< m1 >>
rect 445 390 446 391 
rect 448 390 449 391 
rect 445 395 446 396 
rect 448 395 449 396 
<< m2 >>
rect 445 390 446 391 
rect 448 390 449 391 
rect 445 395 446 396 
rect 448 395 449 396 
<< m2c >>
rect 445 390 446 391 
rect 448 390 449 391 
rect 445 395 446 396 
rect 448 395 449 396 
<< labels >>
rlabel pdiffusion 427 390 428 391  0 t = 1
rlabel pdiffusion 430 390 431 391  0 t = 2
rlabel pdiffusion 427 395 428 396  0 t = 3
rlabel pdiffusion 430 395 431 396  0 t = 4
rlabel pdiffusion 426 390 432 396 0 cell no = 578
<< m1 >>
rect 427 390 428 391 
rect 430 390 431 391 
rect 427 395 428 396 
rect 430 395 431 396 
<< m2 >>
rect 427 390 428 391 
rect 430 390 431 391 
rect 427 395 428 396 
rect 430 395 431 396 
<< m2c >>
rect 427 390 428 391 
rect 430 390 431 391 
rect 427 395 428 396 
rect 430 395 431 396 
<< labels >>
rlabel pdiffusion 445 408 446 409  0 t = 1
rlabel pdiffusion 448 408 449 409  0 t = 2
rlabel pdiffusion 445 413 446 414  0 t = 3
rlabel pdiffusion 448 413 449 414  0 t = 4
rlabel pdiffusion 444 408 450 414 0 cell no = 579
<< m1 >>
rect 445 408 446 409 
rect 448 408 449 409 
rect 445 413 446 414 
rect 448 413 449 414 
<< m2 >>
rect 445 408 446 409 
rect 448 408 449 409 
rect 445 413 446 414 
rect 448 413 449 414 
<< m2c >>
rect 445 408 446 409 
rect 448 408 449 409 
rect 445 413 446 414 
rect 448 413 449 414 
<< labels >>
rlabel pdiffusion 463 390 464 391  0 t = 1
rlabel pdiffusion 466 390 467 391  0 t = 2
rlabel pdiffusion 463 395 464 396  0 t = 3
rlabel pdiffusion 466 395 467 396  0 t = 4
rlabel pdiffusion 462 390 468 396 0 cell no = 580
<< m1 >>
rect 463 390 464 391 
rect 466 390 467 391 
rect 463 395 464 396 
rect 466 395 467 396 
<< m2 >>
rect 463 390 464 391 
rect 466 390 467 391 
rect 463 395 464 396 
rect 466 395 467 396 
<< m2c >>
rect 463 390 464 391 
rect 466 390 467 391 
rect 463 395 464 396 
rect 466 395 467 396 
<< labels >>
rlabel pdiffusion 85 408 86 409  0 t = 1
rlabel pdiffusion 88 408 89 409  0 t = 2
rlabel pdiffusion 85 413 86 414  0 t = 3
rlabel pdiffusion 88 413 89 414  0 t = 4
rlabel pdiffusion 84 408 90 414 0 cell no = 581
<< m1 >>
rect 85 408 86 409 
rect 88 408 89 409 
rect 85 413 86 414 
rect 88 413 89 414 
<< m2 >>
rect 85 408 86 409 
rect 88 408 89 409 
rect 85 413 86 414 
rect 88 413 89 414 
<< m2c >>
rect 85 408 86 409 
rect 88 408 89 409 
rect 85 413 86 414 
rect 88 413 89 414 
<< labels >>
rlabel pdiffusion 85 480 86 481  0 t = 1
rlabel pdiffusion 88 480 89 481  0 t = 2
rlabel pdiffusion 85 485 86 486  0 t = 3
rlabel pdiffusion 88 485 89 486  0 t = 4
rlabel pdiffusion 84 480 90 486 0 cell no = 582
<< m1 >>
rect 85 480 86 481 
rect 88 480 89 481 
rect 85 485 86 486 
rect 88 485 89 486 
<< m2 >>
rect 85 480 86 481 
rect 88 480 89 481 
rect 85 485 86 486 
rect 88 485 89 486 
<< m2c >>
rect 85 480 86 481 
rect 88 480 89 481 
rect 85 485 86 486 
rect 88 485 89 486 
<< labels >>
rlabel pdiffusion 391 156 392 157  0 t = 1
rlabel pdiffusion 394 156 395 157  0 t = 2
rlabel pdiffusion 391 161 392 162  0 t = 3
rlabel pdiffusion 394 161 395 162  0 t = 4
rlabel pdiffusion 390 156 396 162 0 cell no = 583
<< m1 >>
rect 391 156 392 157 
rect 394 156 395 157 
rect 391 161 392 162 
rect 394 161 395 162 
<< m2 >>
rect 391 156 392 157 
rect 394 156 395 157 
rect 391 161 392 162 
rect 394 161 395 162 
<< m2c >>
rect 391 156 392 157 
rect 394 156 395 157 
rect 391 161 392 162 
rect 394 161 395 162 
<< labels >>
rlabel pdiffusion 265 516 266 517  0 t = 1
rlabel pdiffusion 268 516 269 517  0 t = 2
rlabel pdiffusion 265 521 266 522  0 t = 3
rlabel pdiffusion 268 521 269 522  0 t = 4
rlabel pdiffusion 264 516 270 522 0 cell no = 584
<< m1 >>
rect 265 516 266 517 
rect 268 516 269 517 
rect 265 521 266 522 
rect 268 521 269 522 
<< m2 >>
rect 265 516 266 517 
rect 268 516 269 517 
rect 265 521 266 522 
rect 268 521 269 522 
<< m2c >>
rect 265 516 266 517 
rect 268 516 269 517 
rect 265 521 266 522 
rect 268 521 269 522 
<< labels >>
rlabel pdiffusion 49 354 50 355  0 t = 1
rlabel pdiffusion 52 354 53 355  0 t = 2
rlabel pdiffusion 49 359 50 360  0 t = 3
rlabel pdiffusion 52 359 53 360  0 t = 4
rlabel pdiffusion 48 354 54 360 0 cell no = 585
<< m1 >>
rect 49 354 50 355 
rect 52 354 53 355 
rect 49 359 50 360 
rect 52 359 53 360 
<< m2 >>
rect 49 354 50 355 
rect 52 354 53 355 
rect 49 359 50 360 
rect 52 359 53 360 
<< m2c >>
rect 49 354 50 355 
rect 52 354 53 355 
rect 49 359 50 360 
rect 52 359 53 360 
<< labels >>
rlabel pdiffusion 499 228 500 229  0 t = 1
rlabel pdiffusion 502 228 503 229  0 t = 2
rlabel pdiffusion 499 233 500 234  0 t = 3
rlabel pdiffusion 502 233 503 234  0 t = 4
rlabel pdiffusion 498 228 504 234 0 cell no = 586
<< m1 >>
rect 499 228 500 229 
rect 502 228 503 229 
rect 499 233 500 234 
rect 502 233 503 234 
<< m2 >>
rect 499 228 500 229 
rect 502 228 503 229 
rect 499 233 500 234 
rect 502 233 503 234 
<< m2c >>
rect 499 228 500 229 
rect 502 228 503 229 
rect 499 233 500 234 
rect 502 233 503 234 
<< labels >>
rlabel pdiffusion 121 462 122 463  0 t = 1
rlabel pdiffusion 124 462 125 463  0 t = 2
rlabel pdiffusion 121 467 122 468  0 t = 3
rlabel pdiffusion 124 467 125 468  0 t = 4
rlabel pdiffusion 120 462 126 468 0 cell no = 587
<< m1 >>
rect 121 462 122 463 
rect 124 462 125 463 
rect 121 467 122 468 
rect 124 467 125 468 
<< m2 >>
rect 121 462 122 463 
rect 124 462 125 463 
rect 121 467 122 468 
rect 124 467 125 468 
<< m2c >>
rect 121 462 122 463 
rect 124 462 125 463 
rect 121 467 122 468 
rect 124 467 125 468 
<< labels >>
rlabel pdiffusion 13 408 14 409  0 t = 1
rlabel pdiffusion 16 408 17 409  0 t = 2
rlabel pdiffusion 13 413 14 414  0 t = 3
rlabel pdiffusion 16 413 17 414  0 t = 4
rlabel pdiffusion 12 408 18 414 0 cell no = 588
<< m1 >>
rect 13 408 14 409 
rect 16 408 17 409 
rect 13 413 14 414 
rect 16 413 17 414 
<< m2 >>
rect 13 408 14 409 
rect 16 408 17 409 
rect 13 413 14 414 
rect 16 413 17 414 
<< m2c >>
rect 13 408 14 409 
rect 16 408 17 409 
rect 13 413 14 414 
rect 16 413 17 414 
<< labels >>
rlabel pdiffusion 211 390 212 391  0 t = 1
rlabel pdiffusion 214 390 215 391  0 t = 2
rlabel pdiffusion 211 395 212 396  0 t = 3
rlabel pdiffusion 214 395 215 396  0 t = 4
rlabel pdiffusion 210 390 216 396 0 cell no = 589
<< m1 >>
rect 211 390 212 391 
rect 214 390 215 391 
rect 211 395 212 396 
rect 214 395 215 396 
<< m2 >>
rect 211 390 212 391 
rect 214 390 215 391 
rect 211 395 212 396 
rect 214 395 215 396 
<< m2c >>
rect 211 390 212 391 
rect 214 390 215 391 
rect 211 395 212 396 
rect 214 395 215 396 
<< labels >>
rlabel pdiffusion 67 516 68 517  0 t = 1
rlabel pdiffusion 70 516 71 517  0 t = 2
rlabel pdiffusion 67 521 68 522  0 t = 3
rlabel pdiffusion 70 521 71 522  0 t = 4
rlabel pdiffusion 66 516 72 522 0 cell no = 590
<< m1 >>
rect 67 516 68 517 
rect 70 516 71 517 
rect 67 521 68 522 
rect 70 521 71 522 
<< m2 >>
rect 67 516 68 517 
rect 70 516 71 517 
rect 67 521 68 522 
rect 70 521 71 522 
<< m2c >>
rect 67 516 68 517 
rect 70 516 71 517 
rect 67 521 68 522 
rect 70 521 71 522 
<< labels >>
rlabel pdiffusion 193 246 194 247  0 t = 1
rlabel pdiffusion 196 246 197 247  0 t = 2
rlabel pdiffusion 193 251 194 252  0 t = 3
rlabel pdiffusion 196 251 197 252  0 t = 4
rlabel pdiffusion 192 246 198 252 0 cell no = 591
<< m1 >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< m2 >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< m2c >>
rect 193 246 194 247 
rect 196 246 197 247 
rect 193 251 194 252 
rect 196 251 197 252 
<< labels >>
rlabel pdiffusion 427 318 428 319  0 t = 1
rlabel pdiffusion 430 318 431 319  0 t = 2
rlabel pdiffusion 427 323 428 324  0 t = 3
rlabel pdiffusion 430 323 431 324  0 t = 4
rlabel pdiffusion 426 318 432 324 0 cell no = 592
<< m1 >>
rect 427 318 428 319 
rect 430 318 431 319 
rect 427 323 428 324 
rect 430 323 431 324 
<< m2 >>
rect 427 318 428 319 
rect 430 318 431 319 
rect 427 323 428 324 
rect 430 323 431 324 
<< m2c >>
rect 427 318 428 319 
rect 430 318 431 319 
rect 427 323 428 324 
rect 430 323 431 324 
<< labels >>
rlabel pdiffusion 121 516 122 517  0 t = 1
rlabel pdiffusion 124 516 125 517  0 t = 2
rlabel pdiffusion 121 521 122 522  0 t = 3
rlabel pdiffusion 124 521 125 522  0 t = 4
rlabel pdiffusion 120 516 126 522 0 cell no = 593
<< m1 >>
rect 121 516 122 517 
rect 124 516 125 517 
rect 121 521 122 522 
rect 124 521 125 522 
<< m2 >>
rect 121 516 122 517 
rect 124 516 125 517 
rect 121 521 122 522 
rect 124 521 125 522 
<< m2c >>
rect 121 516 122 517 
rect 124 516 125 517 
rect 121 521 122 522 
rect 124 521 125 522 
<< labels >>
rlabel pdiffusion 265 462 266 463  0 t = 1
rlabel pdiffusion 268 462 269 463  0 t = 2
rlabel pdiffusion 265 467 266 468  0 t = 3
rlabel pdiffusion 268 467 269 468  0 t = 4
rlabel pdiffusion 264 462 270 468 0 cell no = 594
<< m1 >>
rect 265 462 266 463 
rect 268 462 269 463 
rect 265 467 266 468 
rect 268 467 269 468 
<< m2 >>
rect 265 462 266 463 
rect 268 462 269 463 
rect 265 467 266 468 
rect 268 467 269 468 
<< m2c >>
rect 265 462 266 463 
rect 268 462 269 463 
rect 265 467 266 468 
rect 268 467 269 468 
<< labels >>
rlabel pdiffusion 301 264 302 265  0 t = 1
rlabel pdiffusion 304 264 305 265  0 t = 2
rlabel pdiffusion 301 269 302 270  0 t = 3
rlabel pdiffusion 304 269 305 270  0 t = 4
rlabel pdiffusion 300 264 306 270 0 cell no = 595
<< m1 >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< m2 >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< m2c >>
rect 301 264 302 265 
rect 304 264 305 265 
rect 301 269 302 270 
rect 304 269 305 270 
<< labels >>
rlabel pdiffusion 319 426 320 427  0 t = 1
rlabel pdiffusion 322 426 323 427  0 t = 2
rlabel pdiffusion 319 431 320 432  0 t = 3
rlabel pdiffusion 322 431 323 432  0 t = 4
rlabel pdiffusion 318 426 324 432 0 cell no = 596
<< m1 >>
rect 319 426 320 427 
rect 322 426 323 427 
rect 319 431 320 432 
rect 322 431 323 432 
<< m2 >>
rect 319 426 320 427 
rect 322 426 323 427 
rect 319 431 320 432 
rect 322 431 323 432 
<< m2c >>
rect 319 426 320 427 
rect 322 426 323 427 
rect 319 431 320 432 
rect 322 431 323 432 
<< labels >>
rlabel pdiffusion 13 120 14 121  0 t = 1
rlabel pdiffusion 16 120 17 121  0 t = 2
rlabel pdiffusion 13 125 14 126  0 t = 3
rlabel pdiffusion 16 125 17 126  0 t = 4
rlabel pdiffusion 12 120 18 126 0 cell no = 597
<< m1 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2 >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< m2c >>
rect 13 120 14 121 
rect 16 120 17 121 
rect 13 125 14 126 
rect 16 125 17 126 
<< labels >>
rlabel pdiffusion 175 174 176 175  0 t = 1
rlabel pdiffusion 178 174 179 175  0 t = 2
rlabel pdiffusion 175 179 176 180  0 t = 3
rlabel pdiffusion 178 179 179 180  0 t = 4
rlabel pdiffusion 174 174 180 180 0 cell no = 598
<< m1 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2 >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< m2c >>
rect 175 174 176 175 
rect 178 174 179 175 
rect 175 179 176 180 
rect 178 179 179 180 
<< labels >>
rlabel pdiffusion 319 354 320 355  0 t = 1
rlabel pdiffusion 322 354 323 355  0 t = 2
rlabel pdiffusion 319 359 320 360  0 t = 3
rlabel pdiffusion 322 359 323 360  0 t = 4
rlabel pdiffusion 318 354 324 360 0 cell no = 599
<< m1 >>
rect 319 354 320 355 
rect 322 354 323 355 
rect 319 359 320 360 
rect 322 359 323 360 
<< m2 >>
rect 319 354 320 355 
rect 322 354 323 355 
rect 319 359 320 360 
rect 322 359 323 360 
<< m2c >>
rect 319 354 320 355 
rect 322 354 323 355 
rect 319 359 320 360 
rect 322 359 323 360 
<< labels >>
rlabel pdiffusion 121 336 122 337  0 t = 1
rlabel pdiffusion 124 336 125 337  0 t = 2
rlabel pdiffusion 121 341 122 342  0 t = 3
rlabel pdiffusion 124 341 125 342  0 t = 4
rlabel pdiffusion 120 336 126 342 0 cell no = 600
<< m1 >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< m2 >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< m2c >>
rect 121 336 122 337 
rect 124 336 125 337 
rect 121 341 122 342 
rect 124 341 125 342 
<< labels >>
rlabel pdiffusion 409 282 410 283  0 t = 1
rlabel pdiffusion 412 282 413 283  0 t = 2
rlabel pdiffusion 409 287 410 288  0 t = 3
rlabel pdiffusion 412 287 413 288  0 t = 4
rlabel pdiffusion 408 282 414 288 0 cell no = 601
<< m1 >>
rect 409 282 410 283 
rect 412 282 413 283 
rect 409 287 410 288 
rect 412 287 413 288 
<< m2 >>
rect 409 282 410 283 
rect 412 282 413 283 
rect 409 287 410 288 
rect 412 287 413 288 
<< m2c >>
rect 409 282 410 283 
rect 412 282 413 283 
rect 409 287 410 288 
rect 412 287 413 288 
<< labels >>
rlabel pdiffusion 193 354 194 355  0 t = 1
rlabel pdiffusion 196 354 197 355  0 t = 2
rlabel pdiffusion 193 359 194 360  0 t = 3
rlabel pdiffusion 196 359 197 360  0 t = 4
rlabel pdiffusion 192 354 198 360 0 cell no = 602
<< m1 >>
rect 193 354 194 355 
rect 196 354 197 355 
rect 193 359 194 360 
rect 196 359 197 360 
<< m2 >>
rect 193 354 194 355 
rect 196 354 197 355 
rect 193 359 194 360 
rect 196 359 197 360 
<< m2c >>
rect 193 354 194 355 
rect 196 354 197 355 
rect 193 359 194 360 
rect 196 359 197 360 
<< labels >>
rlabel pdiffusion 427 480 428 481  0 t = 1
rlabel pdiffusion 430 480 431 481  0 t = 2
rlabel pdiffusion 427 485 428 486  0 t = 3
rlabel pdiffusion 430 485 431 486  0 t = 4
rlabel pdiffusion 426 480 432 486 0 cell no = 603
<< m1 >>
rect 427 480 428 481 
rect 430 480 431 481 
rect 427 485 428 486 
rect 430 485 431 486 
<< m2 >>
rect 427 480 428 481 
rect 430 480 431 481 
rect 427 485 428 486 
rect 430 485 431 486 
<< m2c >>
rect 427 480 428 481 
rect 430 480 431 481 
rect 427 485 428 486 
rect 430 485 431 486 
<< labels >>
rlabel pdiffusion 409 408 410 409  0 t = 1
rlabel pdiffusion 412 408 413 409  0 t = 2
rlabel pdiffusion 409 413 410 414  0 t = 3
rlabel pdiffusion 412 413 413 414  0 t = 4
rlabel pdiffusion 408 408 414 414 0 cell no = 604
<< m1 >>
rect 409 408 410 409 
rect 412 408 413 409 
rect 409 413 410 414 
rect 412 413 413 414 
<< m2 >>
rect 409 408 410 409 
rect 412 408 413 409 
rect 409 413 410 414 
rect 412 413 413 414 
<< m2c >>
rect 409 408 410 409 
rect 412 408 413 409 
rect 409 413 410 414 
rect 412 413 413 414 
<< labels >>
rlabel pdiffusion 517 372 518 373  0 t = 1
rlabel pdiffusion 520 372 521 373  0 t = 2
rlabel pdiffusion 517 377 518 378  0 t = 3
rlabel pdiffusion 520 377 521 378  0 t = 4
rlabel pdiffusion 516 372 522 378 0 cell no = 605
<< m1 >>
rect 517 372 518 373 
rect 520 372 521 373 
rect 517 377 518 378 
rect 520 377 521 378 
<< m2 >>
rect 517 372 518 373 
rect 520 372 521 373 
rect 517 377 518 378 
rect 520 377 521 378 
<< m2c >>
rect 517 372 518 373 
rect 520 372 521 373 
rect 517 377 518 378 
rect 520 377 521 378 
<< labels >>
rlabel pdiffusion 499 336 500 337  0 t = 1
rlabel pdiffusion 502 336 503 337  0 t = 2
rlabel pdiffusion 499 341 500 342  0 t = 3
rlabel pdiffusion 502 341 503 342  0 t = 4
rlabel pdiffusion 498 336 504 342 0 cell no = 606
<< m1 >>
rect 499 336 500 337 
rect 502 336 503 337 
rect 499 341 500 342 
rect 502 341 503 342 
<< m2 >>
rect 499 336 500 337 
rect 502 336 503 337 
rect 499 341 500 342 
rect 502 341 503 342 
<< m2c >>
rect 499 336 500 337 
rect 502 336 503 337 
rect 499 341 500 342 
rect 502 341 503 342 
<< labels >>
rlabel pdiffusion 319 336 320 337  0 t = 1
rlabel pdiffusion 322 336 323 337  0 t = 2
rlabel pdiffusion 319 341 320 342  0 t = 3
rlabel pdiffusion 322 341 323 342  0 t = 4
rlabel pdiffusion 318 336 324 342 0 cell no = 607
<< m1 >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< m2 >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< m2c >>
rect 319 336 320 337 
rect 322 336 323 337 
rect 319 341 320 342 
rect 322 341 323 342 
<< labels >>
rlabel pdiffusion 373 318 374 319  0 t = 1
rlabel pdiffusion 376 318 377 319  0 t = 2
rlabel pdiffusion 373 323 374 324  0 t = 3
rlabel pdiffusion 376 323 377 324  0 t = 4
rlabel pdiffusion 372 318 378 324 0 cell no = 608
<< m1 >>
rect 373 318 374 319 
rect 376 318 377 319 
rect 373 323 374 324 
rect 376 323 377 324 
<< m2 >>
rect 373 318 374 319 
rect 376 318 377 319 
rect 373 323 374 324 
rect 376 323 377 324 
<< m2c >>
rect 373 318 374 319 
rect 376 318 377 319 
rect 373 323 374 324 
rect 376 323 377 324 
<< labels >>
rlabel pdiffusion 517 408 518 409  0 t = 1
rlabel pdiffusion 520 408 521 409  0 t = 2
rlabel pdiffusion 517 413 518 414  0 t = 3
rlabel pdiffusion 520 413 521 414  0 t = 4
rlabel pdiffusion 516 408 522 414 0 cell no = 609
<< m1 >>
rect 517 408 518 409 
rect 520 408 521 409 
rect 517 413 518 414 
rect 520 413 521 414 
<< m2 >>
rect 517 408 518 409 
rect 520 408 521 409 
rect 517 413 518 414 
rect 520 413 521 414 
<< m2c >>
rect 517 408 518 409 
rect 520 408 521 409 
rect 517 413 518 414 
rect 520 413 521 414 
<< labels >>
rlabel pdiffusion 517 30 518 31  0 t = 1
rlabel pdiffusion 520 30 521 31  0 t = 2
rlabel pdiffusion 517 35 518 36  0 t = 3
rlabel pdiffusion 520 35 521 36  0 t = 4
rlabel pdiffusion 516 30 522 36 0 cell no = 610
<< m1 >>
rect 517 30 518 31 
rect 520 30 521 31 
rect 517 35 518 36 
rect 520 35 521 36 
<< m2 >>
rect 517 30 518 31 
rect 520 30 521 31 
rect 517 35 518 36 
rect 520 35 521 36 
<< m2c >>
rect 517 30 518 31 
rect 520 30 521 31 
rect 517 35 518 36 
rect 520 35 521 36 
<< labels >>
rlabel pdiffusion 283 210 284 211  0 t = 1
rlabel pdiffusion 286 210 287 211  0 t = 2
rlabel pdiffusion 283 215 284 216  0 t = 3
rlabel pdiffusion 286 215 287 216  0 t = 4
rlabel pdiffusion 282 210 288 216 0 cell no = 611
<< m1 >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< m2 >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< m2c >>
rect 283 210 284 211 
rect 286 210 287 211 
rect 283 215 284 216 
rect 286 215 287 216 
<< labels >>
rlabel pdiffusion 103 426 104 427  0 t = 1
rlabel pdiffusion 106 426 107 427  0 t = 2
rlabel pdiffusion 103 431 104 432  0 t = 3
rlabel pdiffusion 106 431 107 432  0 t = 4
rlabel pdiffusion 102 426 108 432 0 cell no = 612
<< m1 >>
rect 103 426 104 427 
rect 106 426 107 427 
rect 103 431 104 432 
rect 106 431 107 432 
<< m2 >>
rect 103 426 104 427 
rect 106 426 107 427 
rect 103 431 104 432 
rect 106 431 107 432 
<< m2c >>
rect 103 426 104 427 
rect 106 426 107 427 
rect 103 431 104 432 
rect 106 431 107 432 
<< labels >>
rlabel pdiffusion 337 228 338 229  0 t = 1
rlabel pdiffusion 340 228 341 229  0 t = 2
rlabel pdiffusion 337 233 338 234  0 t = 3
rlabel pdiffusion 340 233 341 234  0 t = 4
rlabel pdiffusion 336 228 342 234 0 cell no = 613
<< m1 >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< m2 >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< m2c >>
rect 337 228 338 229 
rect 340 228 341 229 
rect 337 233 338 234 
rect 340 233 341 234 
<< labels >>
rlabel pdiffusion 265 282 266 283  0 t = 1
rlabel pdiffusion 268 282 269 283  0 t = 2
rlabel pdiffusion 265 287 266 288  0 t = 3
rlabel pdiffusion 268 287 269 288  0 t = 4
rlabel pdiffusion 264 282 270 288 0 cell no = 614
<< m1 >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< m2 >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< m2c >>
rect 265 282 266 283 
rect 268 282 269 283 
rect 265 287 266 288 
rect 268 287 269 288 
<< labels >>
rlabel pdiffusion 175 408 176 409  0 t = 1
rlabel pdiffusion 178 408 179 409  0 t = 2
rlabel pdiffusion 175 413 176 414  0 t = 3
rlabel pdiffusion 178 413 179 414  0 t = 4
rlabel pdiffusion 174 408 180 414 0 cell no = 615
<< m1 >>
rect 175 408 176 409 
rect 178 408 179 409 
rect 175 413 176 414 
rect 178 413 179 414 
<< m2 >>
rect 175 408 176 409 
rect 178 408 179 409 
rect 175 413 176 414 
rect 178 413 179 414 
<< m2c >>
rect 175 408 176 409 
rect 178 408 179 409 
rect 175 413 176 414 
rect 178 413 179 414 
<< labels >>
rlabel pdiffusion 283 192 284 193  0 t = 1
rlabel pdiffusion 286 192 287 193  0 t = 2
rlabel pdiffusion 283 197 284 198  0 t = 3
rlabel pdiffusion 286 197 287 198  0 t = 4
rlabel pdiffusion 282 192 288 198 0 cell no = 616
<< m1 >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< m2 >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< m2c >>
rect 283 192 284 193 
rect 286 192 287 193 
rect 283 197 284 198 
rect 286 197 287 198 
<< labels >>
rlabel pdiffusion 139 516 140 517  0 t = 1
rlabel pdiffusion 142 516 143 517  0 t = 2
rlabel pdiffusion 139 521 140 522  0 t = 3
rlabel pdiffusion 142 521 143 522  0 t = 4
rlabel pdiffusion 138 516 144 522 0 cell no = 617
<< m1 >>
rect 139 516 140 517 
rect 142 516 143 517 
rect 139 521 140 522 
rect 142 521 143 522 
<< m2 >>
rect 139 516 140 517 
rect 142 516 143 517 
rect 139 521 140 522 
rect 142 521 143 522 
<< m2c >>
rect 139 516 140 517 
rect 142 516 143 517 
rect 139 521 140 522 
rect 142 521 143 522 
<< labels >>
rlabel pdiffusion 391 444 392 445  0 t = 1
rlabel pdiffusion 394 444 395 445  0 t = 2
rlabel pdiffusion 391 449 392 450  0 t = 3
rlabel pdiffusion 394 449 395 450  0 t = 4
rlabel pdiffusion 390 444 396 450 0 cell no = 618
<< m1 >>
rect 391 444 392 445 
rect 394 444 395 445 
rect 391 449 392 450 
rect 394 449 395 450 
<< m2 >>
rect 391 444 392 445 
rect 394 444 395 445 
rect 391 449 392 450 
rect 394 449 395 450 
<< m2c >>
rect 391 444 392 445 
rect 394 444 395 445 
rect 391 449 392 450 
rect 394 449 395 450 
<< labels >>
rlabel pdiffusion 373 30 374 31  0 t = 1
rlabel pdiffusion 376 30 377 31  0 t = 2
rlabel pdiffusion 373 35 374 36  0 t = 3
rlabel pdiffusion 376 35 377 36  0 t = 4
rlabel pdiffusion 372 30 378 36 0 cell no = 619
<< m1 >>
rect 373 30 374 31 
rect 376 30 377 31 
rect 373 35 374 36 
rect 376 35 377 36 
<< m2 >>
rect 373 30 374 31 
rect 376 30 377 31 
rect 373 35 374 36 
rect 376 35 377 36 
<< m2c >>
rect 373 30 374 31 
rect 376 30 377 31 
rect 373 35 374 36 
rect 376 35 377 36 
<< labels >>
rlabel pdiffusion 13 336 14 337  0 t = 1
rlabel pdiffusion 16 336 17 337  0 t = 2
rlabel pdiffusion 13 341 14 342  0 t = 3
rlabel pdiffusion 16 341 17 342  0 t = 4
rlabel pdiffusion 12 336 18 342 0 cell no = 620
<< m1 >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< m2 >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< m2c >>
rect 13 336 14 337 
rect 16 336 17 337 
rect 13 341 14 342 
rect 16 341 17 342 
<< labels >>
rlabel pdiffusion 175 516 176 517  0 t = 1
rlabel pdiffusion 178 516 179 517  0 t = 2
rlabel pdiffusion 175 521 176 522  0 t = 3
rlabel pdiffusion 178 521 179 522  0 t = 4
rlabel pdiffusion 174 516 180 522 0 cell no = 621
<< m1 >>
rect 175 516 176 517 
rect 178 516 179 517 
rect 175 521 176 522 
rect 178 521 179 522 
<< m2 >>
rect 175 516 176 517 
rect 178 516 179 517 
rect 175 521 176 522 
rect 178 521 179 522 
<< m2c >>
rect 175 516 176 517 
rect 178 516 179 517 
rect 175 521 176 522 
rect 178 521 179 522 
<< labels >>
rlabel pdiffusion 391 372 392 373  0 t = 1
rlabel pdiffusion 394 372 395 373  0 t = 2
rlabel pdiffusion 391 377 392 378  0 t = 3
rlabel pdiffusion 394 377 395 378  0 t = 4
rlabel pdiffusion 390 372 396 378 0 cell no = 622
<< m1 >>
rect 391 372 392 373 
rect 394 372 395 373 
rect 391 377 392 378 
rect 394 377 395 378 
<< m2 >>
rect 391 372 392 373 
rect 394 372 395 373 
rect 391 377 392 378 
rect 394 377 395 378 
<< m2c >>
rect 391 372 392 373 
rect 394 372 395 373 
rect 391 377 392 378 
rect 394 377 395 378 
<< labels >>
rlabel pdiffusion 157 426 158 427  0 t = 1
rlabel pdiffusion 160 426 161 427  0 t = 2
rlabel pdiffusion 157 431 158 432  0 t = 3
rlabel pdiffusion 160 431 161 432  0 t = 4
rlabel pdiffusion 156 426 162 432 0 cell no = 623
<< m1 >>
rect 157 426 158 427 
rect 160 426 161 427 
rect 157 431 158 432 
rect 160 431 161 432 
<< m2 >>
rect 157 426 158 427 
rect 160 426 161 427 
rect 157 431 158 432 
rect 160 431 161 432 
<< m2c >>
rect 157 426 158 427 
rect 160 426 161 427 
rect 157 431 158 432 
rect 160 431 161 432 
<< labels >>
rlabel pdiffusion 211 462 212 463  0 t = 1
rlabel pdiffusion 214 462 215 463  0 t = 2
rlabel pdiffusion 211 467 212 468  0 t = 3
rlabel pdiffusion 214 467 215 468  0 t = 4
rlabel pdiffusion 210 462 216 468 0 cell no = 624
<< m1 >>
rect 211 462 212 463 
rect 214 462 215 463 
rect 211 467 212 468 
rect 214 467 215 468 
<< m2 >>
rect 211 462 212 463 
rect 214 462 215 463 
rect 211 467 212 468 
rect 214 467 215 468 
<< m2c >>
rect 211 462 212 463 
rect 214 462 215 463 
rect 211 467 212 468 
rect 214 467 215 468 
<< labels >>
rlabel pdiffusion 337 390 338 391  0 t = 1
rlabel pdiffusion 340 390 341 391  0 t = 2
rlabel pdiffusion 337 395 338 396  0 t = 3
rlabel pdiffusion 340 395 341 396  0 t = 4
rlabel pdiffusion 336 390 342 396 0 cell no = 625
<< m1 >>
rect 337 390 338 391 
rect 340 390 341 391 
rect 337 395 338 396 
rect 340 395 341 396 
<< m2 >>
rect 337 390 338 391 
rect 340 390 341 391 
rect 337 395 338 396 
rect 340 395 341 396 
<< m2c >>
rect 337 390 338 391 
rect 340 390 341 391 
rect 337 395 338 396 
rect 340 395 341 396 
<< labels >>
rlabel pdiffusion 211 444 212 445  0 t = 1
rlabel pdiffusion 214 444 215 445  0 t = 2
rlabel pdiffusion 211 449 212 450  0 t = 3
rlabel pdiffusion 214 449 215 450  0 t = 4
rlabel pdiffusion 210 444 216 450 0 cell no = 626
<< m1 >>
rect 211 444 212 445 
rect 214 444 215 445 
rect 211 449 212 450 
rect 214 449 215 450 
<< m2 >>
rect 211 444 212 445 
rect 214 444 215 445 
rect 211 449 212 450 
rect 214 449 215 450 
<< m2c >>
rect 211 444 212 445 
rect 214 444 215 445 
rect 211 449 212 450 
rect 214 449 215 450 
<< labels >>
rlabel pdiffusion 283 408 284 409  0 t = 1
rlabel pdiffusion 286 408 287 409  0 t = 2
rlabel pdiffusion 283 413 284 414  0 t = 3
rlabel pdiffusion 286 413 287 414  0 t = 4
rlabel pdiffusion 282 408 288 414 0 cell no = 627
<< m1 >>
rect 283 408 284 409 
rect 286 408 287 409 
rect 283 413 284 414 
rect 286 413 287 414 
<< m2 >>
rect 283 408 284 409 
rect 286 408 287 409 
rect 283 413 284 414 
rect 286 413 287 414 
<< m2c >>
rect 283 408 284 409 
rect 286 408 287 409 
rect 283 413 284 414 
rect 286 413 287 414 
<< labels >>
rlabel pdiffusion 103 354 104 355  0 t = 1
rlabel pdiffusion 106 354 107 355  0 t = 2
rlabel pdiffusion 103 359 104 360  0 t = 3
rlabel pdiffusion 106 359 107 360  0 t = 4
rlabel pdiffusion 102 354 108 360 0 cell no = 628
<< m1 >>
rect 103 354 104 355 
rect 106 354 107 355 
rect 103 359 104 360 
rect 106 359 107 360 
<< m2 >>
rect 103 354 104 355 
rect 106 354 107 355 
rect 103 359 104 360 
rect 106 359 107 360 
<< m2c >>
rect 103 354 104 355 
rect 106 354 107 355 
rect 103 359 104 360 
rect 106 359 107 360 
<< labels >>
rlabel pdiffusion 301 336 302 337  0 t = 1
rlabel pdiffusion 304 336 305 337  0 t = 2
rlabel pdiffusion 301 341 302 342  0 t = 3
rlabel pdiffusion 304 341 305 342  0 t = 4
rlabel pdiffusion 300 336 306 342 0 cell no = 629
<< m1 >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< m2 >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< m2c >>
rect 301 336 302 337 
rect 304 336 305 337 
rect 301 341 302 342 
rect 304 341 305 342 
<< labels >>
rlabel pdiffusion 373 444 374 445  0 t = 1
rlabel pdiffusion 376 444 377 445  0 t = 2
rlabel pdiffusion 373 449 374 450  0 t = 3
rlabel pdiffusion 376 449 377 450  0 t = 4
rlabel pdiffusion 372 444 378 450 0 cell no = 630
<< m1 >>
rect 373 444 374 445 
rect 376 444 377 445 
rect 373 449 374 450 
rect 376 449 377 450 
<< m2 >>
rect 373 444 374 445 
rect 376 444 377 445 
rect 373 449 374 450 
rect 376 449 377 450 
<< m2c >>
rect 373 444 374 445 
rect 376 444 377 445 
rect 373 449 374 450 
rect 376 449 377 450 
<< labels >>
rlabel pdiffusion 337 498 338 499  0 t = 1
rlabel pdiffusion 340 498 341 499  0 t = 2
rlabel pdiffusion 337 503 338 504  0 t = 3
rlabel pdiffusion 340 503 341 504  0 t = 4
rlabel pdiffusion 336 498 342 504 0 cell no = 631
<< m1 >>
rect 337 498 338 499 
rect 340 498 341 499 
rect 337 503 338 504 
rect 340 503 341 504 
<< m2 >>
rect 337 498 338 499 
rect 340 498 341 499 
rect 337 503 338 504 
rect 340 503 341 504 
<< m2c >>
rect 337 498 338 499 
rect 340 498 341 499 
rect 337 503 338 504 
rect 340 503 341 504 
<< labels >>
rlabel pdiffusion 103 192 104 193  0 t = 1
rlabel pdiffusion 106 192 107 193  0 t = 2
rlabel pdiffusion 103 197 104 198  0 t = 3
rlabel pdiffusion 106 197 107 198  0 t = 4
rlabel pdiffusion 102 192 108 198 0 cell no = 632
<< m1 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2 >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< m2c >>
rect 103 192 104 193 
rect 106 192 107 193 
rect 103 197 104 198 
rect 106 197 107 198 
<< labels >>
rlabel pdiffusion 391 408 392 409  0 t = 1
rlabel pdiffusion 394 408 395 409  0 t = 2
rlabel pdiffusion 391 413 392 414  0 t = 3
rlabel pdiffusion 394 413 395 414  0 t = 4
rlabel pdiffusion 390 408 396 414 0 cell no = 633
<< m1 >>
rect 391 408 392 409 
rect 394 408 395 409 
rect 391 413 392 414 
rect 394 413 395 414 
<< m2 >>
rect 391 408 392 409 
rect 394 408 395 409 
rect 391 413 392 414 
rect 394 413 395 414 
<< m2c >>
rect 391 408 392 409 
rect 394 408 395 409 
rect 391 413 392 414 
rect 394 413 395 414 
<< labels >>
rlabel pdiffusion 517 354 518 355  0 t = 1
rlabel pdiffusion 520 354 521 355  0 t = 2
rlabel pdiffusion 517 359 518 360  0 t = 3
rlabel pdiffusion 520 359 521 360  0 t = 4
rlabel pdiffusion 516 354 522 360 0 cell no = 634
<< m1 >>
rect 517 354 518 355 
rect 520 354 521 355 
rect 517 359 518 360 
rect 520 359 521 360 
<< m2 >>
rect 517 354 518 355 
rect 520 354 521 355 
rect 517 359 518 360 
rect 520 359 521 360 
<< m2c >>
rect 517 354 518 355 
rect 520 354 521 355 
rect 517 359 518 360 
rect 520 359 521 360 
<< labels >>
rlabel pdiffusion 481 462 482 463  0 t = 1
rlabel pdiffusion 484 462 485 463  0 t = 2
rlabel pdiffusion 481 467 482 468  0 t = 3
rlabel pdiffusion 484 467 485 468  0 t = 4
rlabel pdiffusion 480 462 486 468 0 cell no = 635
<< m1 >>
rect 481 462 482 463 
rect 484 462 485 463 
rect 481 467 482 468 
rect 484 467 485 468 
<< m2 >>
rect 481 462 482 463 
rect 484 462 485 463 
rect 481 467 482 468 
rect 484 467 485 468 
<< m2c >>
rect 481 462 482 463 
rect 484 462 485 463 
rect 481 467 482 468 
rect 484 467 485 468 
<< labels >>
rlabel pdiffusion 301 426 302 427  0 t = 1
rlabel pdiffusion 304 426 305 427  0 t = 2
rlabel pdiffusion 301 431 302 432  0 t = 3
rlabel pdiffusion 304 431 305 432  0 t = 4
rlabel pdiffusion 300 426 306 432 0 cell no = 636
<< m1 >>
rect 301 426 302 427 
rect 304 426 305 427 
rect 301 431 302 432 
rect 304 431 305 432 
<< m2 >>
rect 301 426 302 427 
rect 304 426 305 427 
rect 301 431 302 432 
rect 304 431 305 432 
<< m2c >>
rect 301 426 302 427 
rect 304 426 305 427 
rect 301 431 302 432 
rect 304 431 305 432 
<< labels >>
rlabel pdiffusion 481 516 482 517  0 t = 1
rlabel pdiffusion 484 516 485 517  0 t = 2
rlabel pdiffusion 481 521 482 522  0 t = 3
rlabel pdiffusion 484 521 485 522  0 t = 4
rlabel pdiffusion 480 516 486 522 0 cell no = 637
<< m1 >>
rect 481 516 482 517 
rect 484 516 485 517 
rect 481 521 482 522 
rect 484 521 485 522 
<< m2 >>
rect 481 516 482 517 
rect 484 516 485 517 
rect 481 521 482 522 
rect 484 521 485 522 
<< m2c >>
rect 481 516 482 517 
rect 484 516 485 517 
rect 481 521 482 522 
rect 484 521 485 522 
<< labels >>
rlabel pdiffusion 247 264 248 265  0 t = 1
rlabel pdiffusion 250 264 251 265  0 t = 2
rlabel pdiffusion 247 269 248 270  0 t = 3
rlabel pdiffusion 250 269 251 270  0 t = 4
rlabel pdiffusion 246 264 252 270 0 cell no = 638
<< m1 >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< m2 >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< m2c >>
rect 247 264 248 265 
rect 250 264 251 265 
rect 247 269 248 270 
rect 250 269 251 270 
<< labels >>
rlabel pdiffusion 85 354 86 355  0 t = 1
rlabel pdiffusion 88 354 89 355  0 t = 2
rlabel pdiffusion 85 359 86 360  0 t = 3
rlabel pdiffusion 88 359 89 360  0 t = 4
rlabel pdiffusion 84 354 90 360 0 cell no = 639
<< m1 >>
rect 85 354 86 355 
rect 88 354 89 355 
rect 85 359 86 360 
rect 88 359 89 360 
<< m2 >>
rect 85 354 86 355 
rect 88 354 89 355 
rect 85 359 86 360 
rect 88 359 89 360 
<< m2c >>
rect 85 354 86 355 
rect 88 354 89 355 
rect 85 359 86 360 
rect 88 359 89 360 
<< labels >>
rlabel pdiffusion 67 138 68 139  0 t = 1
rlabel pdiffusion 70 138 71 139  0 t = 2
rlabel pdiffusion 67 143 68 144  0 t = 3
rlabel pdiffusion 70 143 71 144  0 t = 4
rlabel pdiffusion 66 138 72 144 0 cell no = 640
<< m1 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2 >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< m2c >>
rect 67 138 68 139 
rect 70 138 71 139 
rect 67 143 68 144 
rect 70 143 71 144 
<< labels >>
rlabel pdiffusion 355 390 356 391  0 t = 1
rlabel pdiffusion 358 390 359 391  0 t = 2
rlabel pdiffusion 355 395 356 396  0 t = 3
rlabel pdiffusion 358 395 359 396  0 t = 4
rlabel pdiffusion 354 390 360 396 0 cell no = 641
<< m1 >>
rect 355 390 356 391 
rect 358 390 359 391 
rect 355 395 356 396 
rect 358 395 359 396 
<< m2 >>
rect 355 390 356 391 
rect 358 390 359 391 
rect 355 395 356 396 
rect 358 395 359 396 
<< m2c >>
rect 355 390 356 391 
rect 358 390 359 391 
rect 355 395 356 396 
rect 358 395 359 396 
<< labels >>
rlabel pdiffusion 391 354 392 355  0 t = 1
rlabel pdiffusion 394 354 395 355  0 t = 2
rlabel pdiffusion 391 359 392 360  0 t = 3
rlabel pdiffusion 394 359 395 360  0 t = 4
rlabel pdiffusion 390 354 396 360 0 cell no = 642
<< m1 >>
rect 391 354 392 355 
rect 394 354 395 355 
rect 391 359 392 360 
rect 394 359 395 360 
<< m2 >>
rect 391 354 392 355 
rect 394 354 395 355 
rect 391 359 392 360 
rect 394 359 395 360 
<< m2c >>
rect 391 354 392 355 
rect 394 354 395 355 
rect 391 359 392 360 
rect 394 359 395 360 
<< labels >>
rlabel pdiffusion 157 246 158 247  0 t = 1
rlabel pdiffusion 160 246 161 247  0 t = 2
rlabel pdiffusion 157 251 158 252  0 t = 3
rlabel pdiffusion 160 251 161 252  0 t = 4
rlabel pdiffusion 156 246 162 252 0 cell no = 643
<< m1 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2 >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< m2c >>
rect 157 246 158 247 
rect 160 246 161 247 
rect 157 251 158 252 
rect 160 251 161 252 
<< labels >>
rlabel pdiffusion 67 336 68 337  0 t = 1
rlabel pdiffusion 70 336 71 337  0 t = 2
rlabel pdiffusion 67 341 68 342  0 t = 3
rlabel pdiffusion 70 341 71 342  0 t = 4
rlabel pdiffusion 66 336 72 342 0 cell no = 644
<< m1 >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< m2 >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< m2c >>
rect 67 336 68 337 
rect 70 336 71 337 
rect 67 341 68 342 
rect 70 341 71 342 
<< labels >>
rlabel pdiffusion 319 102 320 103  0 t = 1
rlabel pdiffusion 322 102 323 103  0 t = 2
rlabel pdiffusion 319 107 320 108  0 t = 3
rlabel pdiffusion 322 107 323 108  0 t = 4
rlabel pdiffusion 318 102 324 108 0 cell no = 645
<< m1 >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< m2 >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< m2c >>
rect 319 102 320 103 
rect 322 102 323 103 
rect 319 107 320 108 
rect 322 107 323 108 
<< labels >>
rlabel pdiffusion 85 48 86 49  0 t = 1
rlabel pdiffusion 88 48 89 49  0 t = 2
rlabel pdiffusion 85 53 86 54  0 t = 3
rlabel pdiffusion 88 53 89 54  0 t = 4
rlabel pdiffusion 84 48 90 54 0 cell no = 646
<< m1 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2 >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< m2c >>
rect 85 48 86 49 
rect 88 48 89 49 
rect 85 53 86 54 
rect 88 53 89 54 
<< labels >>
rlabel pdiffusion 265 300 266 301  0 t = 1
rlabel pdiffusion 268 300 269 301  0 t = 2
rlabel pdiffusion 265 305 266 306  0 t = 3
rlabel pdiffusion 268 305 269 306  0 t = 4
rlabel pdiffusion 264 300 270 306 0 cell no = 647
<< m1 >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< m2 >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< m2c >>
rect 265 300 266 301 
rect 268 300 269 301 
rect 265 305 266 306 
rect 268 305 269 306 
<< labels >>
rlabel pdiffusion 67 408 68 409  0 t = 1
rlabel pdiffusion 70 408 71 409  0 t = 2
rlabel pdiffusion 67 413 68 414  0 t = 3
rlabel pdiffusion 70 413 71 414  0 t = 4
rlabel pdiffusion 66 408 72 414 0 cell no = 648
<< m1 >>
rect 67 408 68 409 
rect 70 408 71 409 
rect 67 413 68 414 
rect 70 413 71 414 
<< m2 >>
rect 67 408 68 409 
rect 70 408 71 409 
rect 67 413 68 414 
rect 70 413 71 414 
<< m2c >>
rect 67 408 68 409 
rect 70 408 71 409 
rect 67 413 68 414 
rect 70 413 71 414 
<< labels >>
rlabel pdiffusion 229 480 230 481  0 t = 1
rlabel pdiffusion 232 480 233 481  0 t = 2
rlabel pdiffusion 229 485 230 486  0 t = 3
rlabel pdiffusion 232 485 233 486  0 t = 4
rlabel pdiffusion 228 480 234 486 0 cell no = 649
<< m1 >>
rect 229 480 230 481 
rect 232 480 233 481 
rect 229 485 230 486 
rect 232 485 233 486 
<< m2 >>
rect 229 480 230 481 
rect 232 480 233 481 
rect 229 485 230 486 
rect 232 485 233 486 
<< m2c >>
rect 229 480 230 481 
rect 232 480 233 481 
rect 229 485 230 486 
rect 232 485 233 486 
<< labels >>
rlabel pdiffusion 283 228 284 229  0 t = 1
rlabel pdiffusion 286 228 287 229  0 t = 2
rlabel pdiffusion 283 233 284 234  0 t = 3
rlabel pdiffusion 286 233 287 234  0 t = 4
rlabel pdiffusion 282 228 288 234 0 cell no = 650
<< m1 >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< m2 >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< m2c >>
rect 283 228 284 229 
rect 286 228 287 229 
rect 283 233 284 234 
rect 286 233 287 234 
<< labels >>
rlabel pdiffusion 265 408 266 409  0 t = 1
rlabel pdiffusion 268 408 269 409  0 t = 2
rlabel pdiffusion 265 413 266 414  0 t = 3
rlabel pdiffusion 268 413 269 414  0 t = 4
rlabel pdiffusion 264 408 270 414 0 cell no = 651
<< m1 >>
rect 265 408 266 409 
rect 268 408 269 409 
rect 265 413 266 414 
rect 268 413 269 414 
<< m2 >>
rect 265 408 266 409 
rect 268 408 269 409 
rect 265 413 266 414 
rect 268 413 269 414 
<< m2c >>
rect 265 408 266 409 
rect 268 408 269 409 
rect 265 413 266 414 
rect 268 413 269 414 
<< labels >>
rlabel pdiffusion 337 318 338 319  0 t = 1
rlabel pdiffusion 340 318 341 319  0 t = 2
rlabel pdiffusion 337 323 338 324  0 t = 3
rlabel pdiffusion 340 323 341 324  0 t = 4
rlabel pdiffusion 336 318 342 324 0 cell no = 652
<< m1 >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< m2 >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< m2c >>
rect 337 318 338 319 
rect 340 318 341 319 
rect 337 323 338 324 
rect 340 323 341 324 
<< labels >>
rlabel pdiffusion 355 516 356 517  0 t = 1
rlabel pdiffusion 358 516 359 517  0 t = 2
rlabel pdiffusion 355 521 356 522  0 t = 3
rlabel pdiffusion 358 521 359 522  0 t = 4
rlabel pdiffusion 354 516 360 522 0 cell no = 653
<< m1 >>
rect 355 516 356 517 
rect 358 516 359 517 
rect 355 521 356 522 
rect 358 521 359 522 
<< m2 >>
rect 355 516 356 517 
rect 358 516 359 517 
rect 355 521 356 522 
rect 358 521 359 522 
<< m2c >>
rect 355 516 356 517 
rect 358 516 359 517 
rect 355 521 356 522 
rect 358 521 359 522 
<< labels >>
rlabel pdiffusion 463 426 464 427  0 t = 1
rlabel pdiffusion 466 426 467 427  0 t = 2
rlabel pdiffusion 463 431 464 432  0 t = 3
rlabel pdiffusion 466 431 467 432  0 t = 4
rlabel pdiffusion 462 426 468 432 0 cell no = 654
<< m1 >>
rect 463 426 464 427 
rect 466 426 467 427 
rect 463 431 464 432 
rect 466 431 467 432 
<< m2 >>
rect 463 426 464 427 
rect 466 426 467 427 
rect 463 431 464 432 
rect 466 431 467 432 
<< m2c >>
rect 463 426 464 427 
rect 466 426 467 427 
rect 463 431 464 432 
rect 466 431 467 432 
<< labels >>
rlabel pdiffusion 193 462 194 463  0 t = 1
rlabel pdiffusion 196 462 197 463  0 t = 2
rlabel pdiffusion 193 467 194 468  0 t = 3
rlabel pdiffusion 196 467 197 468  0 t = 4
rlabel pdiffusion 192 462 198 468 0 cell no = 655
<< m1 >>
rect 193 462 194 463 
rect 196 462 197 463 
rect 193 467 194 468 
rect 196 467 197 468 
<< m2 >>
rect 193 462 194 463 
rect 196 462 197 463 
rect 193 467 194 468 
rect 196 467 197 468 
<< m2c >>
rect 193 462 194 463 
rect 196 462 197 463 
rect 193 467 194 468 
rect 196 467 197 468 
<< labels >>
rlabel pdiffusion 67 390 68 391  0 t = 1
rlabel pdiffusion 70 390 71 391  0 t = 2
rlabel pdiffusion 67 395 68 396  0 t = 3
rlabel pdiffusion 70 395 71 396  0 t = 4
rlabel pdiffusion 66 390 72 396 0 cell no = 656
<< m1 >>
rect 67 390 68 391 
rect 70 390 71 391 
rect 67 395 68 396 
rect 70 395 71 396 
<< m2 >>
rect 67 390 68 391 
rect 70 390 71 391 
rect 67 395 68 396 
rect 70 395 71 396 
<< m2c >>
rect 67 390 68 391 
rect 70 390 71 391 
rect 67 395 68 396 
rect 70 395 71 396 
<< labels >>
rlabel pdiffusion 481 426 482 427  0 t = 1
rlabel pdiffusion 484 426 485 427  0 t = 2
rlabel pdiffusion 481 431 482 432  0 t = 3
rlabel pdiffusion 484 431 485 432  0 t = 4
rlabel pdiffusion 480 426 486 432 0 cell no = 657
<< m1 >>
rect 481 426 482 427 
rect 484 426 485 427 
rect 481 431 482 432 
rect 484 431 485 432 
<< m2 >>
rect 481 426 482 427 
rect 484 426 485 427 
rect 481 431 482 432 
rect 484 431 485 432 
<< m2c >>
rect 481 426 482 427 
rect 484 426 485 427 
rect 481 431 482 432 
rect 484 431 485 432 
<< labels >>
rlabel pdiffusion 301 210 302 211  0 t = 1
rlabel pdiffusion 304 210 305 211  0 t = 2
rlabel pdiffusion 301 215 302 216  0 t = 3
rlabel pdiffusion 304 215 305 216  0 t = 4
rlabel pdiffusion 300 210 306 216 0 cell no = 658
<< m1 >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< m2 >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< m2c >>
rect 301 210 302 211 
rect 304 210 305 211 
rect 301 215 302 216 
rect 304 215 305 216 
<< labels >>
rlabel pdiffusion 517 318 518 319  0 t = 1
rlabel pdiffusion 520 318 521 319  0 t = 2
rlabel pdiffusion 517 323 518 324  0 t = 3
rlabel pdiffusion 520 323 521 324  0 t = 4
rlabel pdiffusion 516 318 522 324 0 cell no = 659
<< m1 >>
rect 517 318 518 319 
rect 520 318 521 319 
rect 517 323 518 324 
rect 520 323 521 324 
<< m2 >>
rect 517 318 518 319 
rect 520 318 521 319 
rect 517 323 518 324 
rect 520 323 521 324 
<< m2c >>
rect 517 318 518 319 
rect 520 318 521 319 
rect 517 323 518 324 
rect 520 323 521 324 
<< labels >>
rlabel pdiffusion 211 372 212 373  0 t = 1
rlabel pdiffusion 214 372 215 373  0 t = 2
rlabel pdiffusion 211 377 212 378  0 t = 3
rlabel pdiffusion 214 377 215 378  0 t = 4
rlabel pdiffusion 210 372 216 378 0 cell no = 660
<< m1 >>
rect 211 372 212 373 
rect 214 372 215 373 
rect 211 377 212 378 
rect 214 377 215 378 
<< m2 >>
rect 211 372 212 373 
rect 214 372 215 373 
rect 211 377 212 378 
rect 214 377 215 378 
<< m2c >>
rect 211 372 212 373 
rect 214 372 215 373 
rect 211 377 212 378 
rect 214 377 215 378 
<< labels >>
rlabel pdiffusion 31 174 32 175  0 t = 1
rlabel pdiffusion 34 174 35 175  0 t = 2
rlabel pdiffusion 31 179 32 180  0 t = 3
rlabel pdiffusion 34 179 35 180  0 t = 4
rlabel pdiffusion 30 174 36 180 0 cell no = 661
<< m1 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2 >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< m2c >>
rect 31 174 32 175 
rect 34 174 35 175 
rect 31 179 32 180 
rect 34 179 35 180 
<< labels >>
rlabel pdiffusion 391 516 392 517  0 t = 1
rlabel pdiffusion 394 516 395 517  0 t = 2
rlabel pdiffusion 391 521 392 522  0 t = 3
rlabel pdiffusion 394 521 395 522  0 t = 4
rlabel pdiffusion 390 516 396 522 0 cell no = 662
<< m1 >>
rect 391 516 392 517 
rect 394 516 395 517 
rect 391 521 392 522 
rect 394 521 395 522 
<< m2 >>
rect 391 516 392 517 
rect 394 516 395 517 
rect 391 521 392 522 
rect 394 521 395 522 
<< m2c >>
rect 391 516 392 517 
rect 394 516 395 517 
rect 391 521 392 522 
rect 394 521 395 522 
<< labels >>
rlabel pdiffusion 373 372 374 373  0 t = 1
rlabel pdiffusion 376 372 377 373  0 t = 2
rlabel pdiffusion 373 377 374 378  0 t = 3
rlabel pdiffusion 376 377 377 378  0 t = 4
rlabel pdiffusion 372 372 378 378 0 cell no = 663
<< m1 >>
rect 373 372 374 373 
rect 376 372 377 373 
rect 373 377 374 378 
rect 376 377 377 378 
<< m2 >>
rect 373 372 374 373 
rect 376 372 377 373 
rect 373 377 374 378 
rect 376 377 377 378 
<< m2c >>
rect 373 372 374 373 
rect 376 372 377 373 
rect 373 377 374 378 
rect 376 377 377 378 
<< labels >>
rlabel pdiffusion 229 408 230 409  0 t = 1
rlabel pdiffusion 232 408 233 409  0 t = 2
rlabel pdiffusion 229 413 230 414  0 t = 3
rlabel pdiffusion 232 413 233 414  0 t = 4
rlabel pdiffusion 228 408 234 414 0 cell no = 664
<< m1 >>
rect 229 408 230 409 
rect 232 408 233 409 
rect 229 413 230 414 
rect 232 413 233 414 
<< m2 >>
rect 229 408 230 409 
rect 232 408 233 409 
rect 229 413 230 414 
rect 232 413 233 414 
<< m2c >>
rect 229 408 230 409 
rect 232 408 233 409 
rect 229 413 230 414 
rect 232 413 233 414 
<< labels >>
rlabel pdiffusion 229 66 230 67  0 t = 1
rlabel pdiffusion 232 66 233 67  0 t = 2
rlabel pdiffusion 229 71 230 72  0 t = 3
rlabel pdiffusion 232 71 233 72  0 t = 4
rlabel pdiffusion 228 66 234 72 0 cell no = 665
<< m1 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2 >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< m2c >>
rect 229 66 230 67 
rect 232 66 233 67 
rect 229 71 230 72 
rect 232 71 233 72 
<< labels >>
rlabel pdiffusion 391 426 392 427  0 t = 1
rlabel pdiffusion 394 426 395 427  0 t = 2
rlabel pdiffusion 391 431 392 432  0 t = 3
rlabel pdiffusion 394 431 395 432  0 t = 4
rlabel pdiffusion 390 426 396 432 0 cell no = 666
<< m1 >>
rect 391 426 392 427 
rect 394 426 395 427 
rect 391 431 392 432 
rect 394 431 395 432 
<< m2 >>
rect 391 426 392 427 
rect 394 426 395 427 
rect 391 431 392 432 
rect 394 431 395 432 
<< m2c >>
rect 391 426 392 427 
rect 394 426 395 427 
rect 391 431 392 432 
rect 394 431 395 432 
<< labels >>
rlabel pdiffusion 517 516 518 517  0 t = 1
rlabel pdiffusion 520 516 521 517  0 t = 2
rlabel pdiffusion 517 521 518 522  0 t = 3
rlabel pdiffusion 520 521 521 522  0 t = 4
rlabel pdiffusion 516 516 522 522 0 cell no = 667
<< m1 >>
rect 517 516 518 517 
rect 520 516 521 517 
rect 517 521 518 522 
rect 520 521 521 522 
<< m2 >>
rect 517 516 518 517 
rect 520 516 521 517 
rect 517 521 518 522 
rect 520 521 521 522 
<< m2c >>
rect 517 516 518 517 
rect 520 516 521 517 
rect 517 521 518 522 
rect 520 521 521 522 
<< labels >>
rlabel pdiffusion 301 192 302 193  0 t = 1
rlabel pdiffusion 304 192 305 193  0 t = 2
rlabel pdiffusion 301 197 302 198  0 t = 3
rlabel pdiffusion 304 197 305 198  0 t = 4
rlabel pdiffusion 300 192 306 198 0 cell no = 668
<< m1 >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< m2 >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< m2c >>
rect 301 192 302 193 
rect 304 192 305 193 
rect 301 197 302 198 
rect 304 197 305 198 
<< labels >>
rlabel pdiffusion 49 372 50 373  0 t = 1
rlabel pdiffusion 52 372 53 373  0 t = 2
rlabel pdiffusion 49 377 50 378  0 t = 3
rlabel pdiffusion 52 377 53 378  0 t = 4
rlabel pdiffusion 48 372 54 378 0 cell no = 669
<< m1 >>
rect 49 372 50 373 
rect 52 372 53 373 
rect 49 377 50 378 
rect 52 377 53 378 
<< m2 >>
rect 49 372 50 373 
rect 52 372 53 373 
rect 49 377 50 378 
rect 52 377 53 378 
<< m2c >>
rect 49 372 50 373 
rect 52 372 53 373 
rect 49 377 50 378 
rect 52 377 53 378 
<< labels >>
rlabel pdiffusion 139 408 140 409  0 t = 1
rlabel pdiffusion 142 408 143 409  0 t = 2
rlabel pdiffusion 139 413 140 414  0 t = 3
rlabel pdiffusion 142 413 143 414  0 t = 4
rlabel pdiffusion 138 408 144 414 0 cell no = 670
<< m1 >>
rect 139 408 140 409 
rect 142 408 143 409 
rect 139 413 140 414 
rect 142 413 143 414 
<< m2 >>
rect 139 408 140 409 
rect 142 408 143 409 
rect 139 413 140 414 
rect 142 413 143 414 
<< m2c >>
rect 139 408 140 409 
rect 142 408 143 409 
rect 139 413 140 414 
rect 142 413 143 414 
<< labels >>
rlabel pdiffusion 247 336 248 337  0 t = 1
rlabel pdiffusion 250 336 251 337  0 t = 2
rlabel pdiffusion 247 341 248 342  0 t = 3
rlabel pdiffusion 250 341 251 342  0 t = 4
rlabel pdiffusion 246 336 252 342 0 cell no = 671
<< m1 >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< m2 >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< m2c >>
rect 247 336 248 337 
rect 250 336 251 337 
rect 247 341 248 342 
rect 250 341 251 342 
<< labels >>
rlabel pdiffusion 13 426 14 427  0 t = 1
rlabel pdiffusion 16 426 17 427  0 t = 2
rlabel pdiffusion 13 431 14 432  0 t = 3
rlabel pdiffusion 16 431 17 432  0 t = 4
rlabel pdiffusion 12 426 18 432 0 cell no = 672
<< m1 >>
rect 13 426 14 427 
rect 16 426 17 427 
rect 13 431 14 432 
rect 16 431 17 432 
<< m2 >>
rect 13 426 14 427 
rect 16 426 17 427 
rect 13 431 14 432 
rect 16 431 17 432 
<< m2c >>
rect 13 426 14 427 
rect 16 426 17 427 
rect 13 431 14 432 
rect 16 431 17 432 
<< labels >>
rlabel pdiffusion 31 444 32 445  0 t = 1
rlabel pdiffusion 34 444 35 445  0 t = 2
rlabel pdiffusion 31 449 32 450  0 t = 3
rlabel pdiffusion 34 449 35 450  0 t = 4
rlabel pdiffusion 30 444 36 450 0 cell no = 673
<< m1 >>
rect 31 444 32 445 
rect 34 444 35 445 
rect 31 449 32 450 
rect 34 449 35 450 
<< m2 >>
rect 31 444 32 445 
rect 34 444 35 445 
rect 31 449 32 450 
rect 34 449 35 450 
<< m2c >>
rect 31 444 32 445 
rect 34 444 35 445 
rect 31 449 32 450 
rect 34 449 35 450 
<< labels >>
rlabel pdiffusion 229 282 230 283  0 t = 1
rlabel pdiffusion 232 282 233 283  0 t = 2
rlabel pdiffusion 229 287 230 288  0 t = 3
rlabel pdiffusion 232 287 233 288  0 t = 4
rlabel pdiffusion 228 282 234 288 0 cell no = 674
<< m1 >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< m2 >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< m2c >>
rect 229 282 230 283 
rect 232 282 233 283 
rect 229 287 230 288 
rect 232 287 233 288 
<< labels >>
rlabel pdiffusion 103 498 104 499  0 t = 1
rlabel pdiffusion 106 498 107 499  0 t = 2
rlabel pdiffusion 103 503 104 504  0 t = 3
rlabel pdiffusion 106 503 107 504  0 t = 4
rlabel pdiffusion 102 498 108 504 0 cell no = 675
<< m1 >>
rect 103 498 104 499 
rect 106 498 107 499 
rect 103 503 104 504 
rect 106 503 107 504 
<< m2 >>
rect 103 498 104 499 
rect 106 498 107 499 
rect 103 503 104 504 
rect 106 503 107 504 
<< m2c >>
rect 103 498 104 499 
rect 106 498 107 499 
rect 103 503 104 504 
rect 106 503 107 504 
<< labels >>
rlabel pdiffusion 31 372 32 373  0 t = 1
rlabel pdiffusion 34 372 35 373  0 t = 2
rlabel pdiffusion 31 377 32 378  0 t = 3
rlabel pdiffusion 34 377 35 378  0 t = 4
rlabel pdiffusion 30 372 36 378 0 cell no = 676
<< m1 >>
rect 31 372 32 373 
rect 34 372 35 373 
rect 31 377 32 378 
rect 34 377 35 378 
<< m2 >>
rect 31 372 32 373 
rect 34 372 35 373 
rect 31 377 32 378 
rect 34 377 35 378 
<< m2c >>
rect 31 372 32 373 
rect 34 372 35 373 
rect 31 377 32 378 
rect 34 377 35 378 
<< labels >>
rlabel pdiffusion 85 462 86 463  0 t = 1
rlabel pdiffusion 88 462 89 463  0 t = 2
rlabel pdiffusion 85 467 86 468  0 t = 3
rlabel pdiffusion 88 467 89 468  0 t = 4
rlabel pdiffusion 84 462 90 468 0 cell no = 677
<< m1 >>
rect 85 462 86 463 
rect 88 462 89 463 
rect 85 467 86 468 
rect 88 467 89 468 
<< m2 >>
rect 85 462 86 463 
rect 88 462 89 463 
rect 85 467 86 468 
rect 88 467 89 468 
<< m2c >>
rect 85 462 86 463 
rect 88 462 89 463 
rect 85 467 86 468 
rect 88 467 89 468 
<< labels >>
rlabel pdiffusion 229 462 230 463  0 t = 1
rlabel pdiffusion 232 462 233 463  0 t = 2
rlabel pdiffusion 229 467 230 468  0 t = 3
rlabel pdiffusion 232 467 233 468  0 t = 4
rlabel pdiffusion 228 462 234 468 0 cell no = 678
<< m1 >>
rect 229 462 230 463 
rect 232 462 233 463 
rect 229 467 230 468 
rect 232 467 233 468 
<< m2 >>
rect 229 462 230 463 
rect 232 462 233 463 
rect 229 467 230 468 
rect 232 467 233 468 
<< m2c >>
rect 229 462 230 463 
rect 232 462 233 463 
rect 229 467 230 468 
rect 232 467 233 468 
<< labels >>
rlabel pdiffusion 301 516 302 517  0 t = 1
rlabel pdiffusion 304 516 305 517  0 t = 2
rlabel pdiffusion 301 521 302 522  0 t = 3
rlabel pdiffusion 304 521 305 522  0 t = 4
rlabel pdiffusion 300 516 306 522 0 cell no = 679
<< m1 >>
rect 301 516 302 517 
rect 304 516 305 517 
rect 301 521 302 522 
rect 304 521 305 522 
<< m2 >>
rect 301 516 302 517 
rect 304 516 305 517 
rect 301 521 302 522 
rect 304 521 305 522 
<< m2c >>
rect 301 516 302 517 
rect 304 516 305 517 
rect 301 521 302 522 
rect 304 521 305 522 
<< labels >>
rlabel pdiffusion 211 498 212 499  0 t = 1
rlabel pdiffusion 214 498 215 499  0 t = 2
rlabel pdiffusion 211 503 212 504  0 t = 3
rlabel pdiffusion 214 503 215 504  0 t = 4
rlabel pdiffusion 210 498 216 504 0 cell no = 680
<< m1 >>
rect 211 498 212 499 
rect 214 498 215 499 
rect 211 503 212 504 
rect 214 503 215 504 
<< m2 >>
rect 211 498 212 499 
rect 214 498 215 499 
rect 211 503 212 504 
rect 214 503 215 504 
<< m2c >>
rect 211 498 212 499 
rect 214 498 215 499 
rect 211 503 212 504 
rect 214 503 215 504 
<< labels >>
rlabel pdiffusion 283 390 284 391  0 t = 1
rlabel pdiffusion 286 390 287 391  0 t = 2
rlabel pdiffusion 283 395 284 396  0 t = 3
rlabel pdiffusion 286 395 287 396  0 t = 4
rlabel pdiffusion 282 390 288 396 0 cell no = 681
<< m1 >>
rect 283 390 284 391 
rect 286 390 287 391 
rect 283 395 284 396 
rect 286 395 287 396 
<< m2 >>
rect 283 390 284 391 
rect 286 390 287 391 
rect 283 395 284 396 
rect 286 395 287 396 
<< m2c >>
rect 283 390 284 391 
rect 286 390 287 391 
rect 283 395 284 396 
rect 286 395 287 396 
<< labels >>
rlabel pdiffusion 301 372 302 373  0 t = 1
rlabel pdiffusion 304 372 305 373  0 t = 2
rlabel pdiffusion 301 377 302 378  0 t = 3
rlabel pdiffusion 304 377 305 378  0 t = 4
rlabel pdiffusion 300 372 306 378 0 cell no = 682
<< m1 >>
rect 301 372 302 373 
rect 304 372 305 373 
rect 301 377 302 378 
rect 304 377 305 378 
<< m2 >>
rect 301 372 302 373 
rect 304 372 305 373 
rect 301 377 302 378 
rect 304 377 305 378 
<< m2c >>
rect 301 372 302 373 
rect 304 372 305 373 
rect 301 377 302 378 
rect 304 377 305 378 
<< labels >>
rlabel pdiffusion 247 390 248 391  0 t = 1
rlabel pdiffusion 250 390 251 391  0 t = 2
rlabel pdiffusion 247 395 248 396  0 t = 3
rlabel pdiffusion 250 395 251 396  0 t = 4
rlabel pdiffusion 246 390 252 396 0 cell no = 683
<< m1 >>
rect 247 390 248 391 
rect 250 390 251 391 
rect 247 395 248 396 
rect 250 395 251 396 
<< m2 >>
rect 247 390 248 391 
rect 250 390 251 391 
rect 247 395 248 396 
rect 250 395 251 396 
<< m2c >>
rect 247 390 248 391 
rect 250 390 251 391 
rect 247 395 248 396 
rect 250 395 251 396 
<< labels >>
rlabel pdiffusion 301 462 302 463  0 t = 1
rlabel pdiffusion 304 462 305 463  0 t = 2
rlabel pdiffusion 301 467 302 468  0 t = 3
rlabel pdiffusion 304 467 305 468  0 t = 4
rlabel pdiffusion 300 462 306 468 0 cell no = 684
<< m1 >>
rect 301 462 302 463 
rect 304 462 305 463 
rect 301 467 302 468 
rect 304 467 305 468 
<< m2 >>
rect 301 462 302 463 
rect 304 462 305 463 
rect 301 467 302 468 
rect 304 467 305 468 
<< m2c >>
rect 301 462 302 463 
rect 304 462 305 463 
rect 301 467 302 468 
rect 304 467 305 468 
<< labels >>
rlabel pdiffusion 283 318 284 319  0 t = 1
rlabel pdiffusion 286 318 287 319  0 t = 2
rlabel pdiffusion 283 323 284 324  0 t = 3
rlabel pdiffusion 286 323 287 324  0 t = 4
rlabel pdiffusion 282 318 288 324 0 cell no = 685
<< m1 >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< m2 >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< m2c >>
rect 283 318 284 319 
rect 286 318 287 319 
rect 283 323 284 324 
rect 286 323 287 324 
<< labels >>
rlabel pdiffusion 373 498 374 499  0 t = 1
rlabel pdiffusion 376 498 377 499  0 t = 2
rlabel pdiffusion 373 503 374 504  0 t = 3
rlabel pdiffusion 376 503 377 504  0 t = 4
rlabel pdiffusion 372 498 378 504 0 cell no = 686
<< m1 >>
rect 373 498 374 499 
rect 376 498 377 499 
rect 373 503 374 504 
rect 376 503 377 504 
<< m2 >>
rect 373 498 374 499 
rect 376 498 377 499 
rect 373 503 374 504 
rect 376 503 377 504 
<< m2c >>
rect 373 498 374 499 
rect 376 498 377 499 
rect 373 503 374 504 
rect 376 503 377 504 
<< labels >>
rlabel pdiffusion 373 426 374 427  0 t = 1
rlabel pdiffusion 376 426 377 427  0 t = 2
rlabel pdiffusion 373 431 374 432  0 t = 3
rlabel pdiffusion 376 431 377 432  0 t = 4
rlabel pdiffusion 372 426 378 432 0 cell no = 687
<< m1 >>
rect 373 426 374 427 
rect 376 426 377 427 
rect 373 431 374 432 
rect 376 431 377 432 
<< m2 >>
rect 373 426 374 427 
rect 376 426 377 427 
rect 373 431 374 432 
rect 376 431 377 432 
<< m2c >>
rect 373 426 374 427 
rect 376 426 377 427 
rect 373 431 374 432 
rect 376 431 377 432 
<< labels >>
rlabel pdiffusion 427 264 428 265  0 t = 1
rlabel pdiffusion 430 264 431 265  0 t = 2
rlabel pdiffusion 427 269 428 270  0 t = 3
rlabel pdiffusion 430 269 431 270  0 t = 4
rlabel pdiffusion 426 264 432 270 0 cell no = 688
<< m1 >>
rect 427 264 428 265 
rect 430 264 431 265 
rect 427 269 428 270 
rect 430 269 431 270 
<< m2 >>
rect 427 264 428 265 
rect 430 264 431 265 
rect 427 269 428 270 
rect 430 269 431 270 
<< m2c >>
rect 427 264 428 265 
rect 430 264 431 265 
rect 427 269 428 270 
rect 430 269 431 270 
<< labels >>
rlabel pdiffusion 391 480 392 481  0 t = 1
rlabel pdiffusion 394 480 395 481  0 t = 2
rlabel pdiffusion 391 485 392 486  0 t = 3
rlabel pdiffusion 394 485 395 486  0 t = 4
rlabel pdiffusion 390 480 396 486 0 cell no = 689
<< m1 >>
rect 391 480 392 481 
rect 394 480 395 481 
rect 391 485 392 486 
rect 394 485 395 486 
<< m2 >>
rect 391 480 392 481 
rect 394 480 395 481 
rect 391 485 392 486 
rect 394 485 395 486 
<< m2c >>
rect 391 480 392 481 
rect 394 480 395 481 
rect 391 485 392 486 
rect 394 485 395 486 
<< labels >>
rlabel pdiffusion 157 390 158 391  0 t = 1
rlabel pdiffusion 160 390 161 391  0 t = 2
rlabel pdiffusion 157 395 158 396  0 t = 3
rlabel pdiffusion 160 395 161 396  0 t = 4
rlabel pdiffusion 156 390 162 396 0 cell no = 690
<< m1 >>
rect 157 390 158 391 
rect 160 390 161 391 
rect 157 395 158 396 
rect 160 395 161 396 
<< m2 >>
rect 157 390 158 391 
rect 160 390 161 391 
rect 157 395 158 396 
rect 160 395 161 396 
<< m2c >>
rect 157 390 158 391 
rect 160 390 161 391 
rect 157 395 158 396 
rect 160 395 161 396 
<< labels >>
rlabel pdiffusion 409 426 410 427  0 t = 1
rlabel pdiffusion 412 426 413 427  0 t = 2
rlabel pdiffusion 409 431 410 432  0 t = 3
rlabel pdiffusion 412 431 413 432  0 t = 4
rlabel pdiffusion 408 426 414 432 0 cell no = 691
<< m1 >>
rect 409 426 410 427 
rect 412 426 413 427 
rect 409 431 410 432 
rect 412 431 413 432 
<< m2 >>
rect 409 426 410 427 
rect 412 426 413 427 
rect 409 431 410 432 
rect 412 431 413 432 
<< m2c >>
rect 409 426 410 427 
rect 412 426 413 427 
rect 409 431 410 432 
rect 412 431 413 432 
<< labels >>
rlabel pdiffusion 499 516 500 517  0 t = 1
rlabel pdiffusion 502 516 503 517  0 t = 2
rlabel pdiffusion 499 521 500 522  0 t = 3
rlabel pdiffusion 502 521 503 522  0 t = 4
rlabel pdiffusion 498 516 504 522 0 cell no = 692
<< m1 >>
rect 499 516 500 517 
rect 502 516 503 517 
rect 499 521 500 522 
rect 502 521 503 522 
<< m2 >>
rect 499 516 500 517 
rect 502 516 503 517 
rect 499 521 500 522 
rect 502 521 503 522 
<< m2c >>
rect 499 516 500 517 
rect 502 516 503 517 
rect 499 521 500 522 
rect 502 521 503 522 
<< labels >>
rlabel pdiffusion 445 498 446 499  0 t = 1
rlabel pdiffusion 448 498 449 499  0 t = 2
rlabel pdiffusion 445 503 446 504  0 t = 3
rlabel pdiffusion 448 503 449 504  0 t = 4
rlabel pdiffusion 444 498 450 504 0 cell no = 693
<< m1 >>
rect 445 498 446 499 
rect 448 498 449 499 
rect 445 503 446 504 
rect 448 503 449 504 
<< m2 >>
rect 445 498 446 499 
rect 448 498 449 499 
rect 445 503 446 504 
rect 448 503 449 504 
<< m2c >>
rect 445 498 446 499 
rect 448 498 449 499 
rect 445 503 446 504 
rect 448 503 449 504 
<< labels >>
rlabel pdiffusion 463 480 464 481  0 t = 1
rlabel pdiffusion 466 480 467 481  0 t = 2
rlabel pdiffusion 463 485 464 486  0 t = 3
rlabel pdiffusion 466 485 467 486  0 t = 4
rlabel pdiffusion 462 480 468 486 0 cell no = 694
<< m1 >>
rect 463 480 464 481 
rect 466 480 467 481 
rect 463 485 464 486 
rect 466 485 467 486 
<< m2 >>
rect 463 480 464 481 
rect 466 480 467 481 
rect 463 485 464 486 
rect 466 485 467 486 
<< m2c >>
rect 463 480 464 481 
rect 466 480 467 481 
rect 463 485 464 486 
rect 466 485 467 486 
<< labels >>
rlabel pdiffusion 499 354 500 355  0 t = 1
rlabel pdiffusion 502 354 503 355  0 t = 2
rlabel pdiffusion 499 359 500 360  0 t = 3
rlabel pdiffusion 502 359 503 360  0 t = 4
rlabel pdiffusion 498 354 504 360 0 cell no = 695
<< m1 >>
rect 499 354 500 355 
rect 502 354 503 355 
rect 499 359 500 360 
rect 502 359 503 360 
<< m2 >>
rect 499 354 500 355 
rect 502 354 503 355 
rect 499 359 500 360 
rect 502 359 503 360 
<< m2c >>
rect 499 354 500 355 
rect 502 354 503 355 
rect 499 359 500 360 
rect 502 359 503 360 
<< labels >>
rlabel pdiffusion 499 372 500 373  0 t = 1
rlabel pdiffusion 502 372 503 373  0 t = 2
rlabel pdiffusion 499 377 500 378  0 t = 3
rlabel pdiffusion 502 377 503 378  0 t = 4
rlabel pdiffusion 498 372 504 378 0 cell no = 696
<< m1 >>
rect 499 372 500 373 
rect 502 372 503 373 
rect 499 377 500 378 
rect 502 377 503 378 
<< m2 >>
rect 499 372 500 373 
rect 502 372 503 373 
rect 499 377 500 378 
rect 502 377 503 378 
<< m2c >>
rect 499 372 500 373 
rect 502 372 503 373 
rect 499 377 500 378 
rect 502 377 503 378 
<< labels >>
rlabel pdiffusion 13 210 14 211  0 t = 1
rlabel pdiffusion 16 210 17 211  0 t = 2
rlabel pdiffusion 13 215 14 216  0 t = 3
rlabel pdiffusion 16 215 17 216  0 t = 4
rlabel pdiffusion 12 210 18 216 0 cell no = 697
<< m1 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2 >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< m2c >>
rect 13 210 14 211 
rect 16 210 17 211 
rect 13 215 14 216 
rect 16 215 17 216 
<< labels >>
rlabel pdiffusion 85 390 86 391  0 t = 1
rlabel pdiffusion 88 390 89 391  0 t = 2
rlabel pdiffusion 85 395 86 396  0 t = 3
rlabel pdiffusion 88 395 89 396  0 t = 4
rlabel pdiffusion 84 390 90 396 0 cell no = 698
<< m1 >>
rect 85 390 86 391 
rect 88 390 89 391 
rect 85 395 86 396 
rect 88 395 89 396 
<< m2 >>
rect 85 390 86 391 
rect 88 390 89 391 
rect 85 395 86 396 
rect 88 395 89 396 
<< m2c >>
rect 85 390 86 391 
rect 88 390 89 391 
rect 85 395 86 396 
rect 88 395 89 396 
<< labels >>
rlabel pdiffusion 67 480 68 481  0 t = 1
rlabel pdiffusion 70 480 71 481  0 t = 2
rlabel pdiffusion 67 485 68 486  0 t = 3
rlabel pdiffusion 70 485 71 486  0 t = 4
rlabel pdiffusion 66 480 72 486 0 cell no = 699
<< m1 >>
rect 67 480 68 481 
rect 70 480 71 481 
rect 67 485 68 486 
rect 70 485 71 486 
<< m2 >>
rect 67 480 68 481 
rect 70 480 71 481 
rect 67 485 68 486 
rect 70 485 71 486 
<< m2c >>
rect 67 480 68 481 
rect 70 480 71 481 
rect 67 485 68 486 
rect 70 485 71 486 
<< labels >>
rlabel pdiffusion 139 354 140 355  0 t = 1
rlabel pdiffusion 142 354 143 355  0 t = 2
rlabel pdiffusion 139 359 140 360  0 t = 3
rlabel pdiffusion 142 359 143 360  0 t = 4
rlabel pdiffusion 138 354 144 360 0 cell no = 700
<< m1 >>
rect 139 354 140 355 
rect 142 354 143 355 
rect 139 359 140 360 
rect 142 359 143 360 
<< m2 >>
rect 139 354 140 355 
rect 142 354 143 355 
rect 139 359 140 360 
rect 142 359 143 360 
<< m2c >>
rect 139 354 140 355 
rect 142 354 143 355 
rect 139 359 140 360 
rect 142 359 143 360 
<< labels >>
rlabel pdiffusion 157 264 158 265  0 t = 1
rlabel pdiffusion 160 264 161 265  0 t = 2
rlabel pdiffusion 157 269 158 270  0 t = 3
rlabel pdiffusion 160 269 161 270  0 t = 4
rlabel pdiffusion 156 264 162 270 0 cell no = 701
<< m1 >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< m2 >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< m2c >>
rect 157 264 158 265 
rect 160 264 161 265 
rect 157 269 158 270 
rect 160 269 161 270 
<< labels >>
rlabel pdiffusion 157 480 158 481  0 t = 1
rlabel pdiffusion 160 480 161 481  0 t = 2
rlabel pdiffusion 157 485 158 486  0 t = 3
rlabel pdiffusion 160 485 161 486  0 t = 4
rlabel pdiffusion 156 480 162 486 0 cell no = 702
<< m1 >>
rect 157 480 158 481 
rect 160 480 161 481 
rect 157 485 158 486 
rect 160 485 161 486 
<< m2 >>
rect 157 480 158 481 
rect 160 480 161 481 
rect 157 485 158 486 
rect 160 485 161 486 
<< m2c >>
rect 157 480 158 481 
rect 160 480 161 481 
rect 157 485 158 486 
rect 160 485 161 486 
<< labels >>
rlabel pdiffusion 103 390 104 391  0 t = 1
rlabel pdiffusion 106 390 107 391  0 t = 2
rlabel pdiffusion 103 395 104 396  0 t = 3
rlabel pdiffusion 106 395 107 396  0 t = 4
rlabel pdiffusion 102 390 108 396 0 cell no = 703
<< m1 >>
rect 103 390 104 391 
rect 106 390 107 391 
rect 103 395 104 396 
rect 106 395 107 396 
<< m2 >>
rect 103 390 104 391 
rect 106 390 107 391 
rect 103 395 104 396 
rect 106 395 107 396 
<< m2c >>
rect 103 390 104 391 
rect 106 390 107 391 
rect 103 395 104 396 
rect 106 395 107 396 
<< labels >>
rlabel pdiffusion 13 498 14 499  0 t = 1
rlabel pdiffusion 16 498 17 499  0 t = 2
rlabel pdiffusion 13 503 14 504  0 t = 3
rlabel pdiffusion 16 503 17 504  0 t = 4
rlabel pdiffusion 12 498 18 504 0 cell no = 704
<< m1 >>
rect 13 498 14 499 
rect 16 498 17 499 
rect 13 503 14 504 
rect 16 503 17 504 
<< m2 >>
rect 13 498 14 499 
rect 16 498 17 499 
rect 13 503 14 504 
rect 16 503 17 504 
<< m2c >>
rect 13 498 14 499 
rect 16 498 17 499 
rect 13 503 14 504 
rect 16 503 17 504 
<< labels >>
rlabel pdiffusion 157 444 158 445  0 t = 1
rlabel pdiffusion 160 444 161 445  0 t = 2
rlabel pdiffusion 157 449 158 450  0 t = 3
rlabel pdiffusion 160 449 161 450  0 t = 4
rlabel pdiffusion 156 444 162 450 0 cell no = 705
<< m1 >>
rect 157 444 158 445 
rect 160 444 161 445 
rect 157 449 158 450 
rect 160 449 161 450 
<< m2 >>
rect 157 444 158 445 
rect 160 444 161 445 
rect 157 449 158 450 
rect 160 449 161 450 
<< m2c >>
rect 157 444 158 445 
rect 160 444 161 445 
rect 157 449 158 450 
rect 160 449 161 450 
<< labels >>
rlabel pdiffusion 121 444 122 445  0 t = 1
rlabel pdiffusion 124 444 125 445  0 t = 2
rlabel pdiffusion 121 449 122 450  0 t = 3
rlabel pdiffusion 124 449 125 450  0 t = 4
rlabel pdiffusion 120 444 126 450 0 cell no = 706
<< m1 >>
rect 121 444 122 445 
rect 124 444 125 445 
rect 121 449 122 450 
rect 124 449 125 450 
<< m2 >>
rect 121 444 122 445 
rect 124 444 125 445 
rect 121 449 122 450 
rect 124 449 125 450 
<< m2c >>
rect 121 444 122 445 
rect 124 444 125 445 
rect 121 449 122 450 
rect 124 449 125 450 
<< labels >>
rlabel pdiffusion 229 444 230 445  0 t = 1
rlabel pdiffusion 232 444 233 445  0 t = 2
rlabel pdiffusion 229 449 230 450  0 t = 3
rlabel pdiffusion 232 449 233 450  0 t = 4
rlabel pdiffusion 228 444 234 450 0 cell no = 707
<< m1 >>
rect 229 444 230 445 
rect 232 444 233 445 
rect 229 449 230 450 
rect 232 449 233 450 
<< m2 >>
rect 229 444 230 445 
rect 232 444 233 445 
rect 229 449 230 450 
rect 232 449 233 450 
<< m2c >>
rect 229 444 230 445 
rect 232 444 233 445 
rect 229 449 230 450 
rect 232 449 233 450 
<< labels >>
rlabel pdiffusion 85 516 86 517  0 t = 1
rlabel pdiffusion 88 516 89 517  0 t = 2
rlabel pdiffusion 85 521 86 522  0 t = 3
rlabel pdiffusion 88 521 89 522  0 t = 4
rlabel pdiffusion 84 516 90 522 0 cell no = 708
<< m1 >>
rect 85 516 86 517 
rect 88 516 89 517 
rect 85 521 86 522 
rect 88 521 89 522 
<< m2 >>
rect 85 516 86 517 
rect 88 516 89 517 
rect 85 521 86 522 
rect 88 521 89 522 
<< m2c >>
rect 85 516 86 517 
rect 88 516 89 517 
rect 85 521 86 522 
rect 88 521 89 522 
<< labels >>
rlabel pdiffusion 157 354 158 355  0 t = 1
rlabel pdiffusion 160 354 161 355  0 t = 2
rlabel pdiffusion 157 359 158 360  0 t = 3
rlabel pdiffusion 160 359 161 360  0 t = 4
rlabel pdiffusion 156 354 162 360 0 cell no = 709
<< m1 >>
rect 157 354 158 355 
rect 160 354 161 355 
rect 157 359 158 360 
rect 160 359 161 360 
<< m2 >>
rect 157 354 158 355 
rect 160 354 161 355 
rect 157 359 158 360 
rect 160 359 161 360 
<< m2c >>
rect 157 354 158 355 
rect 160 354 161 355 
rect 157 359 158 360 
rect 160 359 161 360 
<< labels >>
rlabel pdiffusion 211 480 212 481  0 t = 1
rlabel pdiffusion 214 480 215 481  0 t = 2
rlabel pdiffusion 211 485 212 486  0 t = 3
rlabel pdiffusion 214 485 215 486  0 t = 4
rlabel pdiffusion 210 480 216 486 0 cell no = 710
<< m1 >>
rect 211 480 212 481 
rect 214 480 215 481 
rect 211 485 212 486 
rect 214 485 215 486 
<< m2 >>
rect 211 480 212 481 
rect 214 480 215 481 
rect 211 485 212 486 
rect 214 485 215 486 
<< m2c >>
rect 211 480 212 481 
rect 214 480 215 481 
rect 211 485 212 486 
rect 214 485 215 486 
<< labels >>
rlabel pdiffusion 193 480 194 481  0 t = 1
rlabel pdiffusion 196 480 197 481  0 t = 2
rlabel pdiffusion 193 485 194 486  0 t = 3
rlabel pdiffusion 196 485 197 486  0 t = 4
rlabel pdiffusion 192 480 198 486 0 cell no = 711
<< m1 >>
rect 193 480 194 481 
rect 196 480 197 481 
rect 193 485 194 486 
rect 196 485 197 486 
<< m2 >>
rect 193 480 194 481 
rect 196 480 197 481 
rect 193 485 194 486 
rect 196 485 197 486 
<< m2c >>
rect 193 480 194 481 
rect 196 480 197 481 
rect 193 485 194 486 
rect 196 485 197 486 
<< labels >>
rlabel pdiffusion 373 516 374 517  0 t = 1
rlabel pdiffusion 376 516 377 517  0 t = 2
rlabel pdiffusion 373 521 374 522  0 t = 3
rlabel pdiffusion 376 521 377 522  0 t = 4
rlabel pdiffusion 372 516 378 522 0 cell no = 712
<< m1 >>
rect 373 516 374 517 
rect 376 516 377 517 
rect 373 521 374 522 
rect 376 521 377 522 
<< m2 >>
rect 373 516 374 517 
rect 376 516 377 517 
rect 373 521 374 522 
rect 376 521 377 522 
<< m2c >>
rect 373 516 374 517 
rect 376 516 377 517 
rect 373 521 374 522 
rect 376 521 377 522 
<< labels >>
rlabel pdiffusion 319 480 320 481  0 t = 1
rlabel pdiffusion 322 480 323 481  0 t = 2
rlabel pdiffusion 319 485 320 486  0 t = 3
rlabel pdiffusion 322 485 323 486  0 t = 4
rlabel pdiffusion 318 480 324 486 0 cell no = 713
<< m1 >>
rect 319 480 320 481 
rect 322 480 323 481 
rect 319 485 320 486 
rect 322 485 323 486 
<< m2 >>
rect 319 480 320 481 
rect 322 480 323 481 
rect 319 485 320 486 
rect 322 485 323 486 
<< m2c >>
rect 319 480 320 481 
rect 322 480 323 481 
rect 319 485 320 486 
rect 322 485 323 486 
<< labels >>
rlabel pdiffusion 49 282 50 283  0 t = 1
rlabel pdiffusion 52 282 53 283  0 t = 2
rlabel pdiffusion 49 287 50 288  0 t = 3
rlabel pdiffusion 52 287 53 288  0 t = 4
rlabel pdiffusion 48 282 54 288 0 cell no = 714
<< m1 >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< m2 >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< m2c >>
rect 49 282 50 283 
rect 52 282 53 283 
rect 49 287 50 288 
rect 52 287 53 288 
<< labels >>
rlabel pdiffusion 211 120 212 121  0 t = 1
rlabel pdiffusion 214 120 215 121  0 t = 2
rlabel pdiffusion 211 125 212 126  0 t = 3
rlabel pdiffusion 214 125 215 126  0 t = 4
rlabel pdiffusion 210 120 216 126 0 cell no = 715
<< m1 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2 >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< m2c >>
rect 211 120 212 121 
rect 214 120 215 121 
rect 211 125 212 126 
rect 214 125 215 126 
<< labels >>
rlabel pdiffusion 499 444 500 445  0 t = 1
rlabel pdiffusion 502 444 503 445  0 t = 2
rlabel pdiffusion 499 449 500 450  0 t = 3
rlabel pdiffusion 502 449 503 450  0 t = 4
rlabel pdiffusion 498 444 504 450 0 cell no = 716
<< m1 >>
rect 499 444 500 445 
rect 502 444 503 445 
rect 499 449 500 450 
rect 502 449 503 450 
<< m2 >>
rect 499 444 500 445 
rect 502 444 503 445 
rect 499 449 500 450 
rect 502 449 503 450 
<< m2c >>
rect 499 444 500 445 
rect 502 444 503 445 
rect 499 449 500 450 
rect 502 449 503 450 
<< labels >>
rlabel pdiffusion 319 408 320 409  0 t = 1
rlabel pdiffusion 322 408 323 409  0 t = 2
rlabel pdiffusion 319 413 320 414  0 t = 3
rlabel pdiffusion 322 413 323 414  0 t = 4
rlabel pdiffusion 318 408 324 414 0 cell no = 717
<< m1 >>
rect 319 408 320 409 
rect 322 408 323 409 
rect 319 413 320 414 
rect 322 413 323 414 
<< m2 >>
rect 319 408 320 409 
rect 322 408 323 409 
rect 319 413 320 414 
rect 322 413 323 414 
<< m2c >>
rect 319 408 320 409 
rect 322 408 323 409 
rect 319 413 320 414 
rect 322 413 323 414 
<< labels >>
rlabel pdiffusion 499 426 500 427  0 t = 1
rlabel pdiffusion 502 426 503 427  0 t = 2
rlabel pdiffusion 499 431 500 432  0 t = 3
rlabel pdiffusion 502 431 503 432  0 t = 4
rlabel pdiffusion 498 426 504 432 0 cell no = 718
<< m1 >>
rect 499 426 500 427 
rect 502 426 503 427 
rect 499 431 500 432 
rect 502 431 503 432 
<< m2 >>
rect 499 426 500 427 
rect 502 426 503 427 
rect 499 431 500 432 
rect 502 431 503 432 
<< m2c >>
rect 499 426 500 427 
rect 502 426 503 427 
rect 499 431 500 432 
rect 502 431 503 432 
<< labels >>
rlabel pdiffusion 427 282 428 283  0 t = 1
rlabel pdiffusion 430 282 431 283  0 t = 2
rlabel pdiffusion 427 287 428 288  0 t = 3
rlabel pdiffusion 430 287 431 288  0 t = 4
rlabel pdiffusion 426 282 432 288 0 cell no = 719
<< m1 >>
rect 427 282 428 283 
rect 430 282 431 283 
rect 427 287 428 288 
rect 430 287 431 288 
<< m2 >>
rect 427 282 428 283 
rect 430 282 431 283 
rect 427 287 428 288 
rect 430 287 431 288 
<< m2c >>
rect 427 282 428 283 
rect 430 282 431 283 
rect 427 287 428 288 
rect 430 287 431 288 
<< labels >>
rlabel pdiffusion 175 390 176 391  0 t = 1
rlabel pdiffusion 178 390 179 391  0 t = 2
rlabel pdiffusion 175 395 176 396  0 t = 3
rlabel pdiffusion 178 395 179 396  0 t = 4
rlabel pdiffusion 174 390 180 396 0 cell no = 720
<< m1 >>
rect 175 390 176 391 
rect 178 390 179 391 
rect 175 395 176 396 
rect 178 395 179 396 
<< m2 >>
rect 175 390 176 391 
rect 178 390 179 391 
rect 175 395 176 396 
rect 178 395 179 396 
<< m2c >>
rect 175 390 176 391 
rect 178 390 179 391 
rect 175 395 176 396 
rect 178 395 179 396 
<< labels >>
rlabel pdiffusion 463 516 464 517  0 t = 1
rlabel pdiffusion 466 516 467 517  0 t = 2
rlabel pdiffusion 463 521 464 522  0 t = 3
rlabel pdiffusion 466 521 467 522  0 t = 4
rlabel pdiffusion 462 516 468 522 0 cell no = 721
<< m1 >>
rect 463 516 464 517 
rect 466 516 467 517 
rect 463 521 464 522 
rect 466 521 467 522 
<< m2 >>
rect 463 516 464 517 
rect 466 516 467 517 
rect 463 521 464 522 
rect 466 521 467 522 
<< m2c >>
rect 463 516 464 517 
rect 466 516 467 517 
rect 463 521 464 522 
rect 466 521 467 522 
<< labels >>
rlabel pdiffusion 499 480 500 481  0 t = 1
rlabel pdiffusion 502 480 503 481  0 t = 2
rlabel pdiffusion 499 485 500 486  0 t = 3
rlabel pdiffusion 502 485 503 486  0 t = 4
rlabel pdiffusion 498 480 504 486 0 cell no = 722
<< m1 >>
rect 499 480 500 481 
rect 502 480 503 481 
rect 499 485 500 486 
rect 502 485 503 486 
<< m2 >>
rect 499 480 500 481 
rect 502 480 503 481 
rect 499 485 500 486 
rect 502 485 503 486 
<< m2c >>
rect 499 480 500 481 
rect 502 480 503 481 
rect 499 485 500 486 
rect 502 485 503 486 
<< labels >>
rlabel pdiffusion 211 156 212 157  0 t = 1
rlabel pdiffusion 214 156 215 157  0 t = 2
rlabel pdiffusion 211 161 212 162  0 t = 3
rlabel pdiffusion 214 161 215 162  0 t = 4
rlabel pdiffusion 210 156 216 162 0 cell no = 723
<< m1 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2 >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< m2c >>
rect 211 156 212 157 
rect 214 156 215 157 
rect 211 161 212 162 
rect 214 161 215 162 
<< labels >>
rlabel pdiffusion 499 390 500 391  0 t = 1
rlabel pdiffusion 502 390 503 391  0 t = 2
rlabel pdiffusion 499 395 500 396  0 t = 3
rlabel pdiffusion 502 395 503 396  0 t = 4
rlabel pdiffusion 498 390 504 396 0 cell no = 724
<< m1 >>
rect 499 390 500 391 
rect 502 390 503 391 
rect 499 395 500 396 
rect 502 395 503 396 
<< m2 >>
rect 499 390 500 391 
rect 502 390 503 391 
rect 499 395 500 396 
rect 502 395 503 396 
<< m2c >>
rect 499 390 500 391 
rect 502 390 503 391 
rect 499 395 500 396 
rect 502 395 503 396 
<< labels >>
rlabel pdiffusion 445 516 446 517  0 t = 1
rlabel pdiffusion 448 516 449 517  0 t = 2
rlabel pdiffusion 445 521 446 522  0 t = 3
rlabel pdiffusion 448 521 449 522  0 t = 4
rlabel pdiffusion 444 516 450 522 0 cell no = 725
<< m1 >>
rect 445 516 446 517 
rect 448 516 449 517 
rect 445 521 446 522 
rect 448 521 449 522 
<< m2 >>
rect 445 516 446 517 
rect 448 516 449 517 
rect 445 521 446 522 
rect 448 521 449 522 
<< m2c >>
rect 445 516 446 517 
rect 448 516 449 517 
rect 445 521 446 522 
rect 448 521 449 522 
<< labels >>
rlabel pdiffusion 175 372 176 373  0 t = 1
rlabel pdiffusion 178 372 179 373  0 t = 2
rlabel pdiffusion 175 377 176 378  0 t = 3
rlabel pdiffusion 178 377 179 378  0 t = 4
rlabel pdiffusion 174 372 180 378 0 cell no = 726
<< m1 >>
rect 175 372 176 373 
rect 178 372 179 373 
rect 175 377 176 378 
rect 178 377 179 378 
<< m2 >>
rect 175 372 176 373 
rect 178 372 179 373 
rect 175 377 176 378 
rect 178 377 179 378 
<< m2c >>
rect 175 372 176 373 
rect 178 372 179 373 
rect 175 377 176 378 
rect 178 377 179 378 
<< labels >>
rlabel pdiffusion 103 462 104 463  0 t = 1
rlabel pdiffusion 106 462 107 463  0 t = 2
rlabel pdiffusion 103 467 104 468  0 t = 3
rlabel pdiffusion 106 467 107 468  0 t = 4
rlabel pdiffusion 102 462 108 468 0 cell no = 727
<< m1 >>
rect 103 462 104 463 
rect 106 462 107 463 
rect 103 467 104 468 
rect 106 467 107 468 
<< m2 >>
rect 103 462 104 463 
rect 106 462 107 463 
rect 103 467 104 468 
rect 106 467 107 468 
<< m2c >>
rect 103 462 104 463 
rect 106 462 107 463 
rect 103 467 104 468 
rect 106 467 107 468 
<< labels >>
rlabel pdiffusion 247 156 248 157  0 t = 1
rlabel pdiffusion 250 156 251 157  0 t = 2
rlabel pdiffusion 247 161 248 162  0 t = 3
rlabel pdiffusion 250 161 251 162  0 t = 4
rlabel pdiffusion 246 156 252 162 0 cell no = 728
<< m1 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2 >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< m2c >>
rect 247 156 248 157 
rect 250 156 251 157 
rect 247 161 248 162 
rect 250 161 251 162 
<< labels >>
rlabel pdiffusion 193 336 194 337  0 t = 1
rlabel pdiffusion 196 336 197 337  0 t = 2
rlabel pdiffusion 193 341 194 342  0 t = 3
rlabel pdiffusion 196 341 197 342  0 t = 4
rlabel pdiffusion 192 336 198 342 0 cell no = 729
<< m1 >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< m2 >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< m2c >>
rect 193 336 194 337 
rect 196 336 197 337 
rect 193 341 194 342 
rect 196 341 197 342 
<< labels >>
rlabel pdiffusion 49 444 50 445  0 t = 1
rlabel pdiffusion 52 444 53 445  0 t = 2
rlabel pdiffusion 49 449 50 450  0 t = 3
rlabel pdiffusion 52 449 53 450  0 t = 4
rlabel pdiffusion 48 444 54 450 0 cell no = 730
<< m1 >>
rect 49 444 50 445 
rect 52 444 53 445 
rect 49 449 50 450 
rect 52 449 53 450 
<< m2 >>
rect 49 444 50 445 
rect 52 444 53 445 
rect 49 449 50 450 
rect 52 449 53 450 
<< m2c >>
rect 49 444 50 445 
rect 52 444 53 445 
rect 49 449 50 450 
rect 52 449 53 450 
<< labels >>
rlabel pdiffusion 67 444 68 445  0 t = 1
rlabel pdiffusion 70 444 71 445  0 t = 2
rlabel pdiffusion 67 449 68 450  0 t = 3
rlabel pdiffusion 70 449 71 450  0 t = 4
rlabel pdiffusion 66 444 72 450 0 cell no = 731
<< m1 >>
rect 67 444 68 445 
rect 70 444 71 445 
rect 67 449 68 450 
rect 70 449 71 450 
<< m2 >>
rect 67 444 68 445 
rect 70 444 71 445 
rect 67 449 68 450 
rect 70 449 71 450 
<< m2c >>
rect 67 444 68 445 
rect 70 444 71 445 
rect 67 449 68 450 
rect 70 449 71 450 
<< labels >>
rlabel pdiffusion 157 120 158 121  0 t = 1
rlabel pdiffusion 160 120 161 121  0 t = 2
rlabel pdiffusion 157 125 158 126  0 t = 3
rlabel pdiffusion 160 125 161 126  0 t = 4
rlabel pdiffusion 156 120 162 126 0 cell no = 732
<< m1 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2 >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< m2c >>
rect 157 120 158 121 
rect 160 120 161 121 
rect 157 125 158 126 
rect 160 125 161 126 
<< labels >>
rlabel pdiffusion 175 444 176 445  0 t = 1
rlabel pdiffusion 178 444 179 445  0 t = 2
rlabel pdiffusion 175 449 176 450  0 t = 3
rlabel pdiffusion 178 449 179 450  0 t = 4
rlabel pdiffusion 174 444 180 450 0 cell no = 733
<< m1 >>
rect 175 444 176 445 
rect 178 444 179 445 
rect 175 449 176 450 
rect 178 449 179 450 
<< m2 >>
rect 175 444 176 445 
rect 178 444 179 445 
rect 175 449 176 450 
rect 178 449 179 450 
<< m2c >>
rect 175 444 176 445 
rect 178 444 179 445 
rect 175 449 176 450 
rect 178 449 179 450 
<< labels >>
rlabel pdiffusion 157 462 158 463  0 t = 1
rlabel pdiffusion 160 462 161 463  0 t = 2
rlabel pdiffusion 157 467 158 468  0 t = 3
rlabel pdiffusion 160 467 161 468  0 t = 4
rlabel pdiffusion 156 462 162 468 0 cell no = 734
<< m1 >>
rect 157 462 158 463 
rect 160 462 161 463 
rect 157 467 158 468 
rect 160 467 161 468 
<< m2 >>
rect 157 462 158 463 
rect 160 462 161 463 
rect 157 467 158 468 
rect 160 467 161 468 
<< m2c >>
rect 157 462 158 463 
rect 160 462 161 463 
rect 157 467 158 468 
rect 160 467 161 468 
<< labels >>
rlabel pdiffusion 265 444 266 445  0 t = 1
rlabel pdiffusion 268 444 269 445  0 t = 2
rlabel pdiffusion 265 449 266 450  0 t = 3
rlabel pdiffusion 268 449 269 450  0 t = 4
rlabel pdiffusion 264 444 270 450 0 cell no = 735
<< m1 >>
rect 265 444 266 445 
rect 268 444 269 445 
rect 265 449 266 450 
rect 268 449 269 450 
<< m2 >>
rect 265 444 266 445 
rect 268 444 269 445 
rect 265 449 266 450 
rect 268 449 269 450 
<< m2c >>
rect 265 444 266 445 
rect 268 444 269 445 
rect 265 449 266 450 
rect 268 449 269 450 
<< labels >>
rlabel pdiffusion 301 444 302 445  0 t = 1
rlabel pdiffusion 304 444 305 445  0 t = 2
rlabel pdiffusion 301 449 302 450  0 t = 3
rlabel pdiffusion 304 449 305 450  0 t = 4
rlabel pdiffusion 300 444 306 450 0 cell no = 736
<< m1 >>
rect 301 444 302 445 
rect 304 444 305 445 
rect 301 449 302 450 
rect 304 449 305 450 
<< m2 >>
rect 301 444 302 445 
rect 304 444 305 445 
rect 301 449 302 450 
rect 304 449 305 450 
<< m2c >>
rect 301 444 302 445 
rect 304 444 305 445 
rect 301 449 302 450 
rect 304 449 305 450 
<< labels >>
rlabel pdiffusion 265 336 266 337  0 t = 1
rlabel pdiffusion 268 336 269 337  0 t = 2
rlabel pdiffusion 265 341 266 342  0 t = 3
rlabel pdiffusion 268 341 269 342  0 t = 4
rlabel pdiffusion 264 336 270 342 0 cell no = 737
<< m1 >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< m2 >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< m2c >>
rect 265 336 266 337 
rect 268 336 269 337 
rect 265 341 266 342 
rect 268 341 269 342 
<< labels >>
rlabel pdiffusion 373 390 374 391  0 t = 1
rlabel pdiffusion 376 390 377 391  0 t = 2
rlabel pdiffusion 373 395 374 396  0 t = 3
rlabel pdiffusion 376 395 377 396  0 t = 4
rlabel pdiffusion 372 390 378 396 0 cell no = 738
<< m1 >>
rect 373 390 374 391 
rect 376 390 377 391 
rect 373 395 374 396 
rect 376 395 377 396 
<< m2 >>
rect 373 390 374 391 
rect 376 390 377 391 
rect 373 395 374 396 
rect 376 395 377 396 
<< m2c >>
rect 373 390 374 391 
rect 376 390 377 391 
rect 373 395 374 396 
rect 376 395 377 396 
<< labels >>
rlabel pdiffusion 283 372 284 373  0 t = 1
rlabel pdiffusion 286 372 287 373  0 t = 2
rlabel pdiffusion 283 377 284 378  0 t = 3
rlabel pdiffusion 286 377 287 378  0 t = 4
rlabel pdiffusion 282 372 288 378 0 cell no = 739
<< m1 >>
rect 283 372 284 373 
rect 286 372 287 373 
rect 283 377 284 378 
rect 286 377 287 378 
<< m2 >>
rect 283 372 284 373 
rect 286 372 287 373 
rect 283 377 284 378 
rect 286 377 287 378 
<< m2c >>
rect 283 372 284 373 
rect 286 372 287 373 
rect 283 377 284 378 
rect 286 377 287 378 
<< labels >>
rlabel pdiffusion 301 480 302 481  0 t = 1
rlabel pdiffusion 304 480 305 481  0 t = 2
rlabel pdiffusion 301 485 302 486  0 t = 3
rlabel pdiffusion 304 485 305 486  0 t = 4
rlabel pdiffusion 300 480 306 486 0 cell no = 740
<< m1 >>
rect 301 480 302 481 
rect 304 480 305 481 
rect 301 485 302 486 
rect 304 485 305 486 
<< m2 >>
rect 301 480 302 481 
rect 304 480 305 481 
rect 301 485 302 486 
rect 304 485 305 486 
<< m2c >>
rect 301 480 302 481 
rect 304 480 305 481 
rect 301 485 302 486 
rect 304 485 305 486 
<< labels >>
rlabel pdiffusion 139 426 140 427  0 t = 1
rlabel pdiffusion 142 426 143 427  0 t = 2
rlabel pdiffusion 139 431 140 432  0 t = 3
rlabel pdiffusion 142 431 143 432  0 t = 4
rlabel pdiffusion 138 426 144 432 0 cell no = 741
<< m1 >>
rect 139 426 140 427 
rect 142 426 143 427 
rect 139 431 140 432 
rect 142 431 143 432 
<< m2 >>
rect 139 426 140 427 
rect 142 426 143 427 
rect 139 431 140 432 
rect 142 431 143 432 
<< m2c >>
rect 139 426 140 427 
rect 142 426 143 427 
rect 139 431 140 432 
rect 142 431 143 432 
<< labels >>
rlabel pdiffusion 337 516 338 517  0 t = 1
rlabel pdiffusion 340 516 341 517  0 t = 2
rlabel pdiffusion 337 521 338 522  0 t = 3
rlabel pdiffusion 340 521 341 522  0 t = 4
rlabel pdiffusion 336 516 342 522 0 cell no = 742
<< m1 >>
rect 337 516 338 517 
rect 340 516 341 517 
rect 337 521 338 522 
rect 340 521 341 522 
<< m2 >>
rect 337 516 338 517 
rect 340 516 341 517 
rect 337 521 338 522 
rect 340 521 341 522 
<< m2c >>
rect 337 516 338 517 
rect 340 516 341 517 
rect 337 521 338 522 
rect 340 521 341 522 
<< labels >>
rlabel pdiffusion 427 516 428 517  0 t = 1
rlabel pdiffusion 430 516 431 517  0 t = 2
rlabel pdiffusion 427 521 428 522  0 t = 3
rlabel pdiffusion 430 521 431 522  0 t = 4
rlabel pdiffusion 426 516 432 522 0 cell no = 743
<< m1 >>
rect 427 516 428 517 
rect 430 516 431 517 
rect 427 521 428 522 
rect 430 521 431 522 
<< m2 >>
rect 427 516 428 517 
rect 430 516 431 517 
rect 427 521 428 522 
rect 430 521 431 522 
<< m2c >>
rect 427 516 428 517 
rect 430 516 431 517 
rect 427 521 428 522 
rect 430 521 431 522 
<< labels >>
rlabel pdiffusion 355 444 356 445  0 t = 1
rlabel pdiffusion 358 444 359 445  0 t = 2
rlabel pdiffusion 355 449 356 450  0 t = 3
rlabel pdiffusion 358 449 359 450  0 t = 4
rlabel pdiffusion 354 444 360 450 0 cell no = 744
<< m1 >>
rect 355 444 356 445 
rect 358 444 359 445 
rect 355 449 356 450 
rect 358 449 359 450 
<< m2 >>
rect 355 444 356 445 
rect 358 444 359 445 
rect 355 449 356 450 
rect 358 449 359 450 
<< m2c >>
rect 355 444 356 445 
rect 358 444 359 445 
rect 355 449 356 450 
rect 358 449 359 450 
<< labels >>
rlabel pdiffusion 481 264 482 265  0 t = 1
rlabel pdiffusion 484 264 485 265  0 t = 2
rlabel pdiffusion 481 269 482 270  0 t = 3
rlabel pdiffusion 484 269 485 270  0 t = 4
rlabel pdiffusion 480 264 486 270 0 cell no = 745
<< m1 >>
rect 481 264 482 265 
rect 484 264 485 265 
rect 481 269 482 270 
rect 484 269 485 270 
<< m2 >>
rect 481 264 482 265 
rect 484 264 485 265 
rect 481 269 482 270 
rect 484 269 485 270 
<< m2c >>
rect 481 264 482 265 
rect 484 264 485 265 
rect 481 269 482 270 
rect 484 269 485 270 
<< labels >>
rlabel pdiffusion 337 480 338 481  0 t = 1
rlabel pdiffusion 340 480 341 481  0 t = 2
rlabel pdiffusion 337 485 338 486  0 t = 3
rlabel pdiffusion 340 485 341 486  0 t = 4
rlabel pdiffusion 336 480 342 486 0 cell no = 746
<< m1 >>
rect 337 480 338 481 
rect 340 480 341 481 
rect 337 485 338 486 
rect 340 485 341 486 
<< m2 >>
rect 337 480 338 481 
rect 340 480 341 481 
rect 337 485 338 486 
rect 340 485 341 486 
<< m2c >>
rect 337 480 338 481 
rect 340 480 341 481 
rect 337 485 338 486 
rect 340 485 341 486 
<< labels >>
rlabel pdiffusion 265 498 266 499  0 t = 1
rlabel pdiffusion 268 498 269 499  0 t = 2
rlabel pdiffusion 265 503 266 504  0 t = 3
rlabel pdiffusion 268 503 269 504  0 t = 4
rlabel pdiffusion 264 498 270 504 0 cell no = 747
<< m1 >>
rect 265 498 266 499 
rect 268 498 269 499 
rect 265 503 266 504 
rect 268 503 269 504 
<< m2 >>
rect 265 498 266 499 
rect 268 498 269 499 
rect 265 503 266 504 
rect 268 503 269 504 
<< m2c >>
rect 265 498 266 499 
rect 268 498 269 499 
rect 265 503 266 504 
rect 268 503 269 504 
<< labels >>
rlabel pdiffusion 355 498 356 499  0 t = 1
rlabel pdiffusion 358 498 359 499  0 t = 2
rlabel pdiffusion 355 503 356 504  0 t = 3
rlabel pdiffusion 358 503 359 504  0 t = 4
rlabel pdiffusion 354 498 360 504 0 cell no = 748
<< m1 >>
rect 355 498 356 499 
rect 358 498 359 499 
rect 355 503 356 504 
rect 358 503 359 504 
<< m2 >>
rect 355 498 356 499 
rect 358 498 359 499 
rect 355 503 356 504 
rect 358 503 359 504 
<< m2c >>
rect 355 498 356 499 
rect 358 498 359 499 
rect 355 503 356 504 
rect 358 503 359 504 
<< labels >>
rlabel pdiffusion 499 498 500 499  0 t = 1
rlabel pdiffusion 502 498 503 499  0 t = 2
rlabel pdiffusion 499 503 500 504  0 t = 3
rlabel pdiffusion 502 503 503 504  0 t = 4
rlabel pdiffusion 498 498 504 504 0 cell no = 749
<< m1 >>
rect 499 498 500 499 
rect 502 498 503 499 
rect 499 503 500 504 
rect 502 503 503 504 
<< m2 >>
rect 499 498 500 499 
rect 502 498 503 499 
rect 499 503 500 504 
rect 502 503 503 504 
<< m2c >>
rect 499 498 500 499 
rect 502 498 503 499 
rect 499 503 500 504 
rect 502 503 503 504 
<< labels >>
rlabel pdiffusion 409 462 410 463  0 t = 1
rlabel pdiffusion 412 462 413 463  0 t = 2
rlabel pdiffusion 409 467 410 468  0 t = 3
rlabel pdiffusion 412 467 413 468  0 t = 4
rlabel pdiffusion 408 462 414 468 0 cell no = 750
<< m1 >>
rect 409 462 410 463 
rect 412 462 413 463 
rect 409 467 410 468 
rect 412 467 413 468 
<< m2 >>
rect 409 462 410 463 
rect 412 462 413 463 
rect 409 467 410 468 
rect 412 467 413 468 
<< m2c >>
rect 409 462 410 463 
rect 412 462 413 463 
rect 409 467 410 468 
rect 412 467 413 468 
<< labels >>
rlabel pdiffusion 463 444 464 445  0 t = 1
rlabel pdiffusion 466 444 467 445  0 t = 2
rlabel pdiffusion 463 449 464 450  0 t = 3
rlabel pdiffusion 466 449 467 450  0 t = 4
rlabel pdiffusion 462 444 468 450 0 cell no = 751
<< m1 >>
rect 463 444 464 445 
rect 466 444 467 445 
rect 463 449 464 450 
rect 466 449 467 450 
<< m2 >>
rect 463 444 464 445 
rect 466 444 467 445 
rect 463 449 464 450 
rect 466 449 467 450 
<< m2c >>
rect 463 444 464 445 
rect 466 444 467 445 
rect 463 449 464 450 
rect 466 449 467 450 
<< labels >>
rlabel pdiffusion 409 480 410 481  0 t = 1
rlabel pdiffusion 412 480 413 481  0 t = 2
rlabel pdiffusion 409 485 410 486  0 t = 3
rlabel pdiffusion 412 485 413 486  0 t = 4
rlabel pdiffusion 408 480 414 486 0 cell no = 752
<< m1 >>
rect 409 480 410 481 
rect 412 480 413 481 
rect 409 485 410 486 
rect 412 485 413 486 
<< m2 >>
rect 409 480 410 481 
rect 412 480 413 481 
rect 409 485 410 486 
rect 412 485 413 486 
<< m2c >>
rect 409 480 410 481 
rect 412 480 413 481 
rect 409 485 410 486 
rect 412 485 413 486 
<< labels >>
rlabel pdiffusion 517 498 518 499  0 t = 1
rlabel pdiffusion 520 498 521 499  0 t = 2
rlabel pdiffusion 517 503 518 504  0 t = 3
rlabel pdiffusion 520 503 521 504  0 t = 4
rlabel pdiffusion 516 498 522 504 0 cell no = 753
<< m1 >>
rect 517 498 518 499 
rect 520 498 521 499 
rect 517 503 518 504 
rect 520 503 521 504 
<< m2 >>
rect 517 498 518 499 
rect 520 498 521 499 
rect 517 503 518 504 
rect 520 503 521 504 
<< m2c >>
rect 517 498 518 499 
rect 520 498 521 499 
rect 517 503 518 504 
rect 520 503 521 504 
<< labels >>
rlabel pdiffusion 409 444 410 445  0 t = 1
rlabel pdiffusion 412 444 413 445  0 t = 2
rlabel pdiffusion 409 449 410 450  0 t = 3
rlabel pdiffusion 412 449 413 450  0 t = 4
rlabel pdiffusion 408 444 414 450 0 cell no = 754
<< m1 >>
rect 409 444 410 445 
rect 412 444 413 445 
rect 409 449 410 450 
rect 412 449 413 450 
<< m2 >>
rect 409 444 410 445 
rect 412 444 413 445 
rect 409 449 410 450 
rect 412 449 413 450 
<< m2c >>
rect 409 444 410 445 
rect 412 444 413 445 
rect 409 449 410 450 
rect 412 449 413 450 
<< labels >>
rlabel pdiffusion 49 498 50 499  0 t = 1
rlabel pdiffusion 52 498 53 499  0 t = 2
rlabel pdiffusion 49 503 50 504  0 t = 3
rlabel pdiffusion 52 503 53 504  0 t = 4
rlabel pdiffusion 48 498 54 504 0 cell no = 755
<< m1 >>
rect 49 498 50 499 
rect 52 498 53 499 
rect 49 503 50 504 
rect 52 503 53 504 
<< m2 >>
rect 49 498 50 499 
rect 52 498 53 499 
rect 49 503 50 504 
rect 52 503 53 504 
<< m2c >>
rect 49 498 50 499 
rect 52 498 53 499 
rect 49 503 50 504 
rect 52 503 53 504 
<< labels >>
rlabel pdiffusion 391 300 392 301  0 t = 1
rlabel pdiffusion 394 300 395 301  0 t = 2
rlabel pdiffusion 391 305 392 306  0 t = 3
rlabel pdiffusion 394 305 395 306  0 t = 4
rlabel pdiffusion 390 300 396 306 0 cell no = 756
<< m1 >>
rect 391 300 392 301 
rect 394 300 395 301 
rect 391 305 392 306 
rect 394 305 395 306 
<< m2 >>
rect 391 300 392 301 
rect 394 300 395 301 
rect 391 305 392 306 
rect 394 305 395 306 
<< m2c >>
rect 391 300 392 301 
rect 394 300 395 301 
rect 391 305 392 306 
rect 394 305 395 306 
<< labels >>
rlabel pdiffusion 193 426 194 427  0 t = 1
rlabel pdiffusion 196 426 197 427  0 t = 2
rlabel pdiffusion 193 431 194 432  0 t = 3
rlabel pdiffusion 196 431 197 432  0 t = 4
rlabel pdiffusion 192 426 198 432 0 cell no = 757
<< m1 >>
rect 193 426 194 427 
rect 196 426 197 427 
rect 193 431 194 432 
rect 196 431 197 432 
<< m2 >>
rect 193 426 194 427 
rect 196 426 197 427 
rect 193 431 194 432 
rect 196 431 197 432 
<< m2c >>
rect 193 426 194 427 
rect 196 426 197 427 
rect 193 431 194 432 
rect 196 431 197 432 
<< labels >>
rlabel pdiffusion 121 498 122 499  0 t = 1
rlabel pdiffusion 124 498 125 499  0 t = 2
rlabel pdiffusion 121 503 122 504  0 t = 3
rlabel pdiffusion 124 503 125 504  0 t = 4
rlabel pdiffusion 120 498 126 504 0 cell no = 758
<< m1 >>
rect 121 498 122 499 
rect 124 498 125 499 
rect 121 503 122 504 
rect 124 503 125 504 
<< m2 >>
rect 121 498 122 499 
rect 124 498 125 499 
rect 121 503 122 504 
rect 124 503 125 504 
<< m2c >>
rect 121 498 122 499 
rect 124 498 125 499 
rect 121 503 122 504 
rect 124 503 125 504 
<< labels >>
rlabel pdiffusion 67 498 68 499  0 t = 1
rlabel pdiffusion 70 498 71 499  0 t = 2
rlabel pdiffusion 67 503 68 504  0 t = 3
rlabel pdiffusion 70 503 71 504  0 t = 4
rlabel pdiffusion 66 498 72 504 0 cell no = 759
<< m1 >>
rect 67 498 68 499 
rect 70 498 71 499 
rect 67 503 68 504 
rect 70 503 71 504 
<< m2 >>
rect 67 498 68 499 
rect 70 498 71 499 
rect 67 503 68 504 
rect 70 503 71 504 
<< m2c >>
rect 67 498 68 499 
rect 70 498 71 499 
rect 67 503 68 504 
rect 70 503 71 504 
<< labels >>
rlabel pdiffusion 247 462 248 463  0 t = 1
rlabel pdiffusion 250 462 251 463  0 t = 2
rlabel pdiffusion 247 467 248 468  0 t = 3
rlabel pdiffusion 250 467 251 468  0 t = 4
rlabel pdiffusion 246 462 252 468 0 cell no = 760
<< m1 >>
rect 247 462 248 463 
rect 250 462 251 463 
rect 247 467 248 468 
rect 250 467 251 468 
<< m2 >>
rect 247 462 248 463 
rect 250 462 251 463 
rect 247 467 248 468 
rect 250 467 251 468 
<< m2c >>
rect 247 462 248 463 
rect 250 462 251 463 
rect 247 467 248 468 
rect 250 467 251 468 
<< labels >>
rlabel pdiffusion 31 318 32 319  0 t = 1
rlabel pdiffusion 34 318 35 319  0 t = 2
rlabel pdiffusion 31 323 32 324  0 t = 3
rlabel pdiffusion 34 323 35 324  0 t = 4
rlabel pdiffusion 30 318 36 324 0 cell no = 761
<< m1 >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< m2 >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< m2c >>
rect 31 318 32 319 
rect 34 318 35 319 
rect 31 323 32 324 
rect 34 323 35 324 
<< labels >>
rlabel pdiffusion 157 516 158 517  0 t = 1
rlabel pdiffusion 160 516 161 517  0 t = 2
rlabel pdiffusion 157 521 158 522  0 t = 3
rlabel pdiffusion 160 521 161 522  0 t = 4
rlabel pdiffusion 156 516 162 522 0 cell no = 762
<< m1 >>
rect 157 516 158 517 
rect 160 516 161 517 
rect 157 521 158 522 
rect 160 521 161 522 
<< m2 >>
rect 157 516 158 517 
rect 160 516 161 517 
rect 157 521 158 522 
rect 160 521 161 522 
<< m2c >>
rect 157 516 158 517 
rect 160 516 161 517 
rect 157 521 158 522 
rect 160 521 161 522 
<< labels >>
rlabel pdiffusion 283 498 284 499  0 t = 1
rlabel pdiffusion 286 498 287 499  0 t = 2
rlabel pdiffusion 283 503 284 504  0 t = 3
rlabel pdiffusion 286 503 287 504  0 t = 4
rlabel pdiffusion 282 498 288 504 0 cell no = 763
<< m1 >>
rect 283 498 284 499 
rect 286 498 287 499 
rect 283 503 284 504 
rect 286 503 287 504 
<< m2 >>
rect 283 498 284 499 
rect 286 498 287 499 
rect 283 503 284 504 
rect 286 503 287 504 
<< m2c >>
rect 283 498 284 499 
rect 286 498 287 499 
rect 283 503 284 504 
rect 286 503 287 504 
<< labels >>
rlabel pdiffusion 337 300 338 301  0 t = 1
rlabel pdiffusion 340 300 341 301  0 t = 2
rlabel pdiffusion 337 305 338 306  0 t = 3
rlabel pdiffusion 340 305 341 306  0 t = 4
rlabel pdiffusion 336 300 342 306 0 cell no = 764
<< m1 >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< m2 >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< m2c >>
rect 337 300 338 301 
rect 340 300 341 301 
rect 337 305 338 306 
rect 340 305 341 306 
<< labels >>
rlabel pdiffusion 283 300 284 301  0 t = 1
rlabel pdiffusion 286 300 287 301  0 t = 2
rlabel pdiffusion 283 305 284 306  0 t = 3
rlabel pdiffusion 286 305 287 306  0 t = 4
rlabel pdiffusion 282 300 288 306 0 cell no = 765
<< m1 >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< m2 >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< m2c >>
rect 283 300 284 301 
rect 286 300 287 301 
rect 283 305 284 306 
rect 286 305 287 306 
<< labels >>
rlabel pdiffusion 139 372 140 373  0 t = 1
rlabel pdiffusion 142 372 143 373  0 t = 2
rlabel pdiffusion 139 377 140 378  0 t = 3
rlabel pdiffusion 142 377 143 378  0 t = 4
rlabel pdiffusion 138 372 144 378 0 cell no = 766
<< m1 >>
rect 139 372 140 373 
rect 142 372 143 373 
rect 139 377 140 378 
rect 142 377 143 378 
<< m2 >>
rect 139 372 140 373 
rect 142 372 143 373 
rect 139 377 140 378 
rect 142 377 143 378 
<< m2c >>
rect 139 372 140 373 
rect 142 372 143 373 
rect 139 377 140 378 
rect 142 377 143 378 
<< labels >>
rlabel pdiffusion 193 66 194 67  0 t = 1
rlabel pdiffusion 196 66 197 67  0 t = 2
rlabel pdiffusion 193 71 194 72  0 t = 3
rlabel pdiffusion 196 71 197 72  0 t = 4
rlabel pdiffusion 192 66 198 72 0 cell no = 767
<< m1 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2 >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< m2c >>
rect 193 66 194 67 
rect 196 66 197 67 
rect 193 71 194 72 
rect 196 71 197 72 
<< labels >>
rlabel pdiffusion 211 408 212 409  0 t = 1
rlabel pdiffusion 214 408 215 409  0 t = 2
rlabel pdiffusion 211 413 212 414  0 t = 3
rlabel pdiffusion 214 413 215 414  0 t = 4
rlabel pdiffusion 210 408 216 414 0 cell no = 768
<< m1 >>
rect 211 408 212 409 
rect 214 408 215 409 
rect 211 413 212 414 
rect 214 413 215 414 
<< m2 >>
rect 211 408 212 409 
rect 214 408 215 409 
rect 211 413 212 414 
rect 214 413 215 414 
<< m2c >>
rect 211 408 212 409 
rect 214 408 215 409 
rect 211 413 212 414 
rect 214 413 215 414 
<< labels >>
rlabel pdiffusion 427 462 428 463  0 t = 1
rlabel pdiffusion 430 462 431 463  0 t = 2
rlabel pdiffusion 427 467 428 468  0 t = 3
rlabel pdiffusion 430 467 431 468  0 t = 4
rlabel pdiffusion 426 462 432 468 0 cell no = 769
<< m1 >>
rect 427 462 428 463 
rect 430 462 431 463 
rect 427 467 428 468 
rect 430 467 431 468 
<< m2 >>
rect 427 462 428 463 
rect 430 462 431 463 
rect 427 467 428 468 
rect 430 467 431 468 
<< m2c >>
rect 427 462 428 463 
rect 430 462 431 463 
rect 427 467 428 468 
rect 430 467 431 468 
<< labels >>
rlabel pdiffusion 445 192 446 193  0 t = 1
rlabel pdiffusion 448 192 449 193  0 t = 2
rlabel pdiffusion 445 197 446 198  0 t = 3
rlabel pdiffusion 448 197 449 198  0 t = 4
rlabel pdiffusion 444 192 450 198 0 cell no = 770
<< m1 >>
rect 445 192 446 193 
rect 448 192 449 193 
rect 445 197 446 198 
rect 448 197 449 198 
<< m2 >>
rect 445 192 446 193 
rect 448 192 449 193 
rect 445 197 446 198 
rect 448 197 449 198 
<< m2c >>
rect 445 192 446 193 
rect 448 192 449 193 
rect 445 197 446 198 
rect 448 197 449 198 
<< labels >>
rlabel pdiffusion 283 516 284 517  0 t = 1
rlabel pdiffusion 286 516 287 517  0 t = 2
rlabel pdiffusion 283 521 284 522  0 t = 3
rlabel pdiffusion 286 521 287 522  0 t = 4
rlabel pdiffusion 282 516 288 522 0 cell no = 771
<< m1 >>
rect 283 516 284 517 
rect 286 516 287 517 
rect 283 521 284 522 
rect 286 521 287 522 
<< m2 >>
rect 283 516 284 517 
rect 286 516 287 517 
rect 283 521 284 522 
rect 286 521 287 522 
<< m2c >>
rect 283 516 284 517 
rect 286 516 287 517 
rect 283 521 284 522 
rect 286 521 287 522 
<< labels >>
rlabel pdiffusion 319 462 320 463  0 t = 1
rlabel pdiffusion 322 462 323 463  0 t = 2
rlabel pdiffusion 319 467 320 468  0 t = 3
rlabel pdiffusion 322 467 323 468  0 t = 4
rlabel pdiffusion 318 462 324 468 0 cell no = 772
<< m1 >>
rect 319 462 320 463 
rect 322 462 323 463 
rect 319 467 320 468 
rect 322 467 323 468 
<< m2 >>
rect 319 462 320 463 
rect 322 462 323 463 
rect 319 467 320 468 
rect 322 467 323 468 
<< m2c >>
rect 319 462 320 463 
rect 322 462 323 463 
rect 319 467 320 468 
rect 322 467 323 468 
<< labels >>
rlabel pdiffusion 409 516 410 517  0 t = 1
rlabel pdiffusion 412 516 413 517  0 t = 2
rlabel pdiffusion 409 521 410 522  0 t = 3
rlabel pdiffusion 412 521 413 522  0 t = 4
rlabel pdiffusion 408 516 414 522 0 cell no = 773
<< m1 >>
rect 409 516 410 517 
rect 412 516 413 517 
rect 409 521 410 522 
rect 412 521 413 522 
<< m2 >>
rect 409 516 410 517 
rect 412 516 413 517 
rect 409 521 410 522 
rect 412 521 413 522 
<< m2c >>
rect 409 516 410 517 
rect 412 516 413 517 
rect 409 521 410 522 
rect 412 521 413 522 
<< labels >>
rlabel pdiffusion 463 462 464 463  0 t = 1
rlabel pdiffusion 466 462 467 463  0 t = 2
rlabel pdiffusion 463 467 464 468  0 t = 3
rlabel pdiffusion 466 467 467 468  0 t = 4
rlabel pdiffusion 462 462 468 468 0 cell no = 774
<< m1 >>
rect 463 462 464 463 
rect 466 462 467 463 
rect 463 467 464 468 
rect 466 467 467 468 
<< m2 >>
rect 463 462 464 463 
rect 466 462 467 463 
rect 463 467 464 468 
rect 466 467 467 468 
<< m2c >>
rect 463 462 464 463 
rect 466 462 467 463 
rect 463 467 464 468 
rect 466 467 467 468 
<< labels >>
rlabel pdiffusion 337 462 338 463  0 t = 1
rlabel pdiffusion 340 462 341 463  0 t = 2
rlabel pdiffusion 337 467 338 468  0 t = 3
rlabel pdiffusion 340 467 341 468  0 t = 4
rlabel pdiffusion 336 462 342 468 0 cell no = 775
<< m1 >>
rect 337 462 338 463 
rect 340 462 341 463 
rect 337 467 338 468 
rect 340 467 341 468 
<< m2 >>
rect 337 462 338 463 
rect 340 462 341 463 
rect 337 467 338 468 
rect 340 467 341 468 
<< m2c >>
rect 337 462 338 463 
rect 340 462 341 463 
rect 337 467 338 468 
rect 340 467 341 468 
<< labels >>
rlabel pdiffusion 391 462 392 463  0 t = 1
rlabel pdiffusion 394 462 395 463  0 t = 2
rlabel pdiffusion 391 467 392 468  0 t = 3
rlabel pdiffusion 394 467 395 468  0 t = 4
rlabel pdiffusion 390 462 396 468 0 cell no = 776
<< m1 >>
rect 391 462 392 463 
rect 394 462 395 463 
rect 391 467 392 468 
rect 394 467 395 468 
<< m2 >>
rect 391 462 392 463 
rect 394 462 395 463 
rect 391 467 392 468 
rect 394 467 395 468 
<< m2c >>
rect 391 462 392 463 
rect 394 462 395 463 
rect 391 467 392 468 
rect 394 467 395 468 
<< labels >>
rlabel pdiffusion 463 498 464 499  0 t = 1
rlabel pdiffusion 466 498 467 499  0 t = 2
rlabel pdiffusion 463 503 464 504  0 t = 3
rlabel pdiffusion 466 503 467 504  0 t = 4
rlabel pdiffusion 462 498 468 504 0 cell no = 777
<< m1 >>
rect 463 498 464 499 
rect 466 498 467 499 
rect 463 503 464 504 
rect 466 503 467 504 
<< m2 >>
rect 463 498 464 499 
rect 466 498 467 499 
rect 463 503 464 504 
rect 466 503 467 504 
<< m2c >>
rect 463 498 464 499 
rect 466 498 467 499 
rect 463 503 464 504 
rect 466 503 467 504 
<< labels >>
rlabel pdiffusion 517 426 518 427  0 t = 1
rlabel pdiffusion 520 426 521 427  0 t = 2
rlabel pdiffusion 517 431 518 432  0 t = 3
rlabel pdiffusion 520 431 521 432  0 t = 4
rlabel pdiffusion 516 426 522 432 0 cell no = 778
<< m1 >>
rect 517 426 518 427 
rect 520 426 521 427 
rect 517 431 518 432 
rect 520 431 521 432 
<< m2 >>
rect 517 426 518 427 
rect 520 426 521 427 
rect 517 431 518 432 
rect 520 431 521 432 
<< m2c >>
rect 517 426 518 427 
rect 520 426 521 427 
rect 517 431 518 432 
rect 520 431 521 432 
<< labels >>
rlabel pdiffusion 499 462 500 463  0 t = 1
rlabel pdiffusion 502 462 503 463  0 t = 2
rlabel pdiffusion 499 467 500 468  0 t = 3
rlabel pdiffusion 502 467 503 468  0 t = 4
rlabel pdiffusion 498 462 504 468 0 cell no = 779
<< m1 >>
rect 499 462 500 463 
rect 502 462 503 463 
rect 499 467 500 468 
rect 502 467 503 468 
<< m2 >>
rect 499 462 500 463 
rect 502 462 503 463 
rect 499 467 500 468 
rect 502 467 503 468 
<< m2c >>
rect 499 462 500 463 
rect 502 462 503 463 
rect 499 467 500 468 
rect 502 467 503 468 
<< labels >>
rlabel pdiffusion 265 318 266 319  0 t = 1
rlabel pdiffusion 268 318 269 319  0 t = 2
rlabel pdiffusion 265 323 266 324  0 t = 3
rlabel pdiffusion 268 323 269 324  0 t = 4
rlabel pdiffusion 264 318 270 324 0 cell no = 780
<< m1 >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< m2 >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< m2c >>
rect 265 318 266 319 
rect 268 318 269 319 
rect 265 323 266 324 
rect 268 323 269 324 
<< labels >>
rlabel pdiffusion 481 480 482 481  0 t = 1
rlabel pdiffusion 484 480 485 481  0 t = 2
rlabel pdiffusion 481 485 482 486  0 t = 3
rlabel pdiffusion 484 485 485 486  0 t = 4
rlabel pdiffusion 480 480 486 486 0 cell no = 781
<< m1 >>
rect 481 480 482 481 
rect 484 480 485 481 
rect 481 485 482 486 
rect 484 485 485 486 
<< m2 >>
rect 481 480 482 481 
rect 484 480 485 481 
rect 481 485 482 486 
rect 484 485 485 486 
<< m2c >>
rect 481 480 482 481 
rect 484 480 485 481 
rect 481 485 482 486 
rect 484 485 485 486 
<< labels >>
rlabel pdiffusion 445 480 446 481  0 t = 1
rlabel pdiffusion 448 480 449 481  0 t = 2
rlabel pdiffusion 445 485 446 486  0 t = 3
rlabel pdiffusion 448 485 449 486  0 t = 4
rlabel pdiffusion 444 480 450 486 0 cell no = 782
<< m1 >>
rect 445 480 446 481 
rect 448 480 449 481 
rect 445 485 446 486 
rect 448 485 449 486 
<< m2 >>
rect 445 480 446 481 
rect 448 480 449 481 
rect 445 485 446 486 
rect 448 485 449 486 
<< m2c >>
rect 445 480 446 481 
rect 448 480 449 481 
rect 445 485 446 486 
rect 448 485 449 486 
<< labels >>
rlabel pdiffusion 229 354 230 355  0 t = 1
rlabel pdiffusion 232 354 233 355  0 t = 2
rlabel pdiffusion 229 359 230 360  0 t = 3
rlabel pdiffusion 232 359 233 360  0 t = 4
rlabel pdiffusion 228 354 234 360 0 cell no = 783
<< m1 >>
rect 229 354 230 355 
rect 232 354 233 355 
rect 229 359 230 360 
rect 232 359 233 360 
<< m2 >>
rect 229 354 230 355 
rect 232 354 233 355 
rect 229 359 230 360 
rect 232 359 233 360 
<< m2c >>
rect 229 354 230 355 
rect 232 354 233 355 
rect 229 359 230 360 
rect 232 359 233 360 
<< labels >>
rlabel pdiffusion 31 516 32 517  0 t = 1
rlabel pdiffusion 34 516 35 517  0 t = 2
rlabel pdiffusion 31 521 32 522  0 t = 3
rlabel pdiffusion 34 521 35 522  0 t = 4
rlabel pdiffusion 30 516 36 522 0 cell no = 784
<< m1 >>
rect 31 516 32 517 
rect 34 516 35 517 
rect 31 521 32 522 
rect 34 521 35 522 
<< m2 >>
rect 31 516 32 517 
rect 34 516 35 517 
rect 31 521 32 522 
rect 34 521 35 522 
<< m2c >>
rect 31 516 32 517 
rect 34 516 35 517 
rect 31 521 32 522 
rect 34 521 35 522 
<< labels >>
rlabel pdiffusion 103 444 104 445  0 t = 1
rlabel pdiffusion 106 444 107 445  0 t = 2
rlabel pdiffusion 103 449 104 450  0 t = 3
rlabel pdiffusion 106 449 107 450  0 t = 4
rlabel pdiffusion 102 444 108 450 0 cell no = 785
<< m1 >>
rect 103 444 104 445 
rect 106 444 107 445 
rect 103 449 104 450 
rect 106 449 107 450 
<< m2 >>
rect 103 444 104 445 
rect 106 444 107 445 
rect 103 449 104 450 
rect 106 449 107 450 
<< m2c >>
rect 103 444 104 445 
rect 106 444 107 445 
rect 103 449 104 450 
rect 106 449 107 450 
<< labels >>
rlabel pdiffusion 31 480 32 481  0 t = 1
rlabel pdiffusion 34 480 35 481  0 t = 2
rlabel pdiffusion 31 485 32 486  0 t = 3
rlabel pdiffusion 34 485 35 486  0 t = 4
rlabel pdiffusion 30 480 36 486 0 cell no = 786
<< m1 >>
rect 31 480 32 481 
rect 34 480 35 481 
rect 31 485 32 486 
rect 34 485 35 486 
<< m2 >>
rect 31 480 32 481 
rect 34 480 35 481 
rect 31 485 32 486 
rect 34 485 35 486 
<< m2c >>
rect 31 480 32 481 
rect 34 480 35 481 
rect 31 485 32 486 
rect 34 485 35 486 
<< labels >>
rlabel pdiffusion 175 156 176 157  0 t = 1
rlabel pdiffusion 178 156 179 157  0 t = 2
rlabel pdiffusion 175 161 176 162  0 t = 3
rlabel pdiffusion 178 161 179 162  0 t = 4
rlabel pdiffusion 174 156 180 162 0 cell no = 787
<< m1 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2 >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< m2c >>
rect 175 156 176 157 
rect 178 156 179 157 
rect 175 161 176 162 
rect 178 161 179 162 
<< labels >>
rlabel pdiffusion 85 498 86 499  0 t = 1
rlabel pdiffusion 88 498 89 499  0 t = 2
rlabel pdiffusion 85 503 86 504  0 t = 3
rlabel pdiffusion 88 503 89 504  0 t = 4
rlabel pdiffusion 84 498 90 504 0 cell no = 788
<< m1 >>
rect 85 498 86 499 
rect 88 498 89 499 
rect 85 503 86 504 
rect 88 503 89 504 
<< m2 >>
rect 85 498 86 499 
rect 88 498 89 499 
rect 85 503 86 504 
rect 88 503 89 504 
<< m2c >>
rect 85 498 86 499 
rect 88 498 89 499 
rect 85 503 86 504 
rect 88 503 89 504 
<< labels >>
rlabel pdiffusion 31 300 32 301  0 t = 1
rlabel pdiffusion 34 300 35 301  0 t = 2
rlabel pdiffusion 31 305 32 306  0 t = 3
rlabel pdiffusion 34 305 35 306  0 t = 4
rlabel pdiffusion 30 300 36 306 0 cell no = 789
<< m1 >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< m2 >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< m2c >>
rect 31 300 32 301 
rect 34 300 35 301 
rect 31 305 32 306 
rect 34 305 35 306 
<< labels >>
rlabel pdiffusion 193 516 194 517  0 t = 1
rlabel pdiffusion 196 516 197 517  0 t = 2
rlabel pdiffusion 193 521 194 522  0 t = 3
rlabel pdiffusion 196 521 197 522  0 t = 4
rlabel pdiffusion 192 516 198 522 0 cell no = 790
<< m1 >>
rect 193 516 194 517 
rect 196 516 197 517 
rect 193 521 194 522 
rect 196 521 197 522 
<< m2 >>
rect 193 516 194 517 
rect 196 516 197 517 
rect 193 521 194 522 
rect 196 521 197 522 
<< m2c >>
rect 193 516 194 517 
rect 196 516 197 517 
rect 193 521 194 522 
rect 196 521 197 522 
<< labels >>
rlabel pdiffusion 49 516 50 517  0 t = 1
rlabel pdiffusion 52 516 53 517  0 t = 2
rlabel pdiffusion 49 521 50 522  0 t = 3
rlabel pdiffusion 52 521 53 522  0 t = 4
rlabel pdiffusion 48 516 54 522 0 cell no = 791
<< m1 >>
rect 49 516 50 517 
rect 52 516 53 517 
rect 49 521 50 522 
rect 52 521 53 522 
<< m2 >>
rect 49 516 50 517 
rect 52 516 53 517 
rect 49 521 50 522 
rect 52 521 53 522 
<< m2c >>
rect 49 516 50 517 
rect 52 516 53 517 
rect 49 521 50 522 
rect 52 521 53 522 
<< labels >>
rlabel pdiffusion 355 480 356 481  0 t = 1
rlabel pdiffusion 358 480 359 481  0 t = 2
rlabel pdiffusion 355 485 356 486  0 t = 3
rlabel pdiffusion 358 485 359 486  0 t = 4
rlabel pdiffusion 354 480 360 486 0 cell no = 792
<< m1 >>
rect 355 480 356 481 
rect 358 480 359 481 
rect 355 485 356 486 
rect 358 485 359 486 
<< m2 >>
rect 355 480 356 481 
rect 358 480 359 481 
rect 355 485 356 486 
rect 358 485 359 486 
<< m2c >>
rect 355 480 356 481 
rect 358 480 359 481 
rect 355 485 356 486 
rect 358 485 359 486 
<< labels >>
rlabel pdiffusion 13 444 14 445  0 t = 1
rlabel pdiffusion 16 444 17 445  0 t = 2
rlabel pdiffusion 13 449 14 450  0 t = 3
rlabel pdiffusion 16 449 17 450  0 t = 4
rlabel pdiffusion 12 444 18 450 0 cell no = 793
<< m1 >>
rect 13 444 14 445 
rect 16 444 17 445 
rect 13 449 14 450 
rect 16 449 17 450 
<< m2 >>
rect 13 444 14 445 
rect 16 444 17 445 
rect 13 449 14 450 
rect 16 449 17 450 
<< m2c >>
rect 13 444 14 445 
rect 16 444 17 445 
rect 13 449 14 450 
rect 16 449 17 450 
<< labels >>
rlabel pdiffusion 247 516 248 517  0 t = 1
rlabel pdiffusion 250 516 251 517  0 t = 2
rlabel pdiffusion 247 521 248 522  0 t = 3
rlabel pdiffusion 250 521 251 522  0 t = 4
rlabel pdiffusion 246 516 252 522 0 cell no = 794
<< m1 >>
rect 247 516 248 517 
rect 250 516 251 517 
rect 247 521 248 522 
rect 250 521 251 522 
<< m2 >>
rect 247 516 248 517 
rect 250 516 251 517 
rect 247 521 248 522 
rect 250 521 251 522 
<< m2c >>
rect 247 516 248 517 
rect 250 516 251 517 
rect 247 521 248 522 
rect 250 521 251 522 
<< labels >>
rlabel pdiffusion 247 426 248 427  0 t = 1
rlabel pdiffusion 250 426 251 427  0 t = 2
rlabel pdiffusion 247 431 248 432  0 t = 3
rlabel pdiffusion 250 431 251 432  0 t = 4
rlabel pdiffusion 246 426 252 432 0 cell no = 795
<< m1 >>
rect 247 426 248 427 
rect 250 426 251 427 
rect 247 431 248 432 
rect 250 431 251 432 
<< m2 >>
rect 247 426 248 427 
rect 250 426 251 427 
rect 247 431 248 432 
rect 250 431 251 432 
<< m2c >>
rect 247 426 248 427 
rect 250 426 251 427 
rect 247 431 248 432 
rect 250 431 251 432 
<< labels >>
rlabel pdiffusion 85 210 86 211  0 t = 1
rlabel pdiffusion 88 210 89 211  0 t = 2
rlabel pdiffusion 85 215 86 216  0 t = 3
rlabel pdiffusion 88 215 89 216  0 t = 4
rlabel pdiffusion 84 210 90 216 0 cell no = 796
<< m1 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2 >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< m2c >>
rect 85 210 86 211 
rect 88 210 89 211 
rect 85 215 86 216 
rect 88 215 89 216 
<< labels >>
rlabel pdiffusion 175 498 176 499  0 t = 1
rlabel pdiffusion 178 498 179 499  0 t = 2
rlabel pdiffusion 175 503 176 504  0 t = 3
rlabel pdiffusion 178 503 179 504  0 t = 4
rlabel pdiffusion 174 498 180 504 0 cell no = 797
<< m1 >>
rect 175 498 176 499 
rect 178 498 179 499 
rect 175 503 176 504 
rect 178 503 179 504 
<< m2 >>
rect 175 498 176 499 
rect 178 498 179 499 
rect 175 503 176 504 
rect 178 503 179 504 
<< m2c >>
rect 175 498 176 499 
rect 178 498 179 499 
rect 175 503 176 504 
rect 178 503 179 504 
<< labels >>
rlabel pdiffusion 283 462 284 463  0 t = 1
rlabel pdiffusion 286 462 287 463  0 t = 2
rlabel pdiffusion 283 467 284 468  0 t = 3
rlabel pdiffusion 286 467 287 468  0 t = 4
rlabel pdiffusion 282 462 288 468 0 cell no = 798
<< m1 >>
rect 283 462 284 463 
rect 286 462 287 463 
rect 283 467 284 468 
rect 286 467 287 468 
<< m2 >>
rect 283 462 284 463 
rect 286 462 287 463 
rect 283 467 284 468 
rect 286 467 287 468 
<< m2c >>
rect 283 462 284 463 
rect 286 462 287 463 
rect 283 467 284 468 
rect 286 467 287 468 
<< labels >>
rlabel pdiffusion 481 318 482 319  0 t = 1
rlabel pdiffusion 484 318 485 319  0 t = 2
rlabel pdiffusion 481 323 482 324  0 t = 3
rlabel pdiffusion 484 323 485 324  0 t = 4
rlabel pdiffusion 480 318 486 324 0 cell no = 799
<< m1 >>
rect 481 318 482 319 
rect 484 318 485 319 
rect 481 323 482 324 
rect 484 323 485 324 
<< m2 >>
rect 481 318 482 319 
rect 484 318 485 319 
rect 481 323 482 324 
rect 484 323 485 324 
<< m2c >>
rect 481 318 482 319 
rect 484 318 485 319 
rect 481 323 482 324 
rect 484 323 485 324 
<< labels >>
rlabel pdiffusion 409 390 410 391  0 t = 1
rlabel pdiffusion 412 390 413 391  0 t = 2
rlabel pdiffusion 409 395 410 396  0 t = 3
rlabel pdiffusion 412 395 413 396  0 t = 4
rlabel pdiffusion 408 390 414 396 0 cell no = 800
<< m1 >>
rect 409 390 410 391 
rect 412 390 413 391 
rect 409 395 410 396 
rect 412 395 413 396 
<< m2 >>
rect 409 390 410 391 
rect 412 390 413 391 
rect 409 395 410 396 
rect 412 395 413 396 
<< m2c >>
rect 409 390 410 391 
rect 412 390 413 391 
rect 409 395 410 396 
rect 412 395 413 396 
<< end >> 
